// Benchmark "x3.blif" written by ABC on Fri Feb 25 15:12:41 2022

module x3  ( 
    b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y,
    z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, r0, s0,
    t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1,
    l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2,
    d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2,
    v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3,
    n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4,
    f4, g4, h4,
    i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4,
    a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5,
    s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6,
    k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7,
    c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7,
    u7, v7, w7, x7, y7, z7, a8, b8, c8  );
  input  b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v,
    w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0,
    r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1,
    j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2,
    b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2,
    t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3,
    l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4,
    d4, e4, f4, g4, h4;
  output i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4,
    z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5,
    r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6,
    j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7,
    b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7,
    t7, u7, v7, w7, x7, y7, z7, a8, b8, c8;
  wire new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n301_, new_n302_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n351_, new_n352_, new_n353_, new_n354_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n366_, new_n367_, new_n368_, new_n369_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n381_, new_n382_, new_n383_, new_n384_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n433_, new_n434_, new_n435_, new_n436_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n448_, new_n449_, new_n450_, new_n451_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n463_, new_n464_, new_n465_, new_n466_, new_n468_,
    new_n469_, new_n470_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n570_,
    new_n571_, new_n572_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1008_, new_n1010_, new_n1011_, new_n1012_, new_n1014_, new_n1015_,
    new_n1016_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1064_,
    new_n1065_, new_n1066_;
  assign i4 = ~x1 | a2;
  assign new_n236_ = ~d & ~e;
  assign new_n237_ = q2 & r2;
  assign new_n238_ = ~x1 & new_n237_;
  assign new_n239_ = i2 & new_n238_;
  assign new_n240_ = ~o0 & ~new_n239_;
  assign new_n241_ = new_n236_ & ~new_n240_;
  assign new_n242_ = ~c & new_n241_;
  assign j4 = y1 | new_n242_;
  assign new_n244_ = i0 & ~l2;
  assign new_n245_ = ~h0 & ~new_n244_;
  assign new_n246_ = ~i0 & ~l2;
  assign new_n247_ = n2 & ~new_n246_;
  assign new_n248_ = ~new_n245_ & new_n247_;
  assign new_n249_ = k0 & ~l2;
  assign new_n250_ = ~j0 & ~new_n249_;
  assign new_n251_ = ~k0 & ~l2;
  assign new_n252_ = ~n2 & ~new_n251_;
  assign new_n253_ = ~new_n250_ & new_n252_;
  assign new_n254_ = ~o2 & ~p2;
  assign new_n255_ = m2 & ~new_n253_;
  assign new_n256_ = new_n248_ & ~new_n255_;
  assign new_n257_ = m2 & new_n253_;
  assign new_n258_ = ~new_n256_ & ~new_n257_;
  assign new_n259_ = new_n254_ & ~new_n258_;
  assign new_n260_ = ~y1 & new_n259_;
  assign new_n261_ = ~j2 & ~k2;
  assign new_n262_ = ~a2 & new_n261_;
  assign new_n263_ = ~q2 & ~r2;
  assign new_n264_ = i2 & ~new_n263_;
  assign new_n265_ = ~y1 & ~a2;
  assign new_n266_ = z1 & r2;
  assign new_n267_ = ~z1 & r2;
  assign new_n268_ = c0 & ~new_n267_;
  assign new_n269_ = ~new_n266_ & ~new_n268_;
  assign new_n270_ = ~i2 & ~i3;
  assign new_n271_ = d0 & r2;
  assign new_n272_ = ~q2 & ~new_n271_;
  assign new_n273_ = ~new_n270_ & ~new_n272_;
  assign new_n274_ = ~i2 & i3;
  assign new_n275_ = ~new_n273_ & ~new_n274_;
  assign new_n276_ = ~r2 & i3;
  assign new_n277_ = new_n275_ & ~new_n276_;
  assign new_n278_ = i2 & ~new_n269_;
  assign new_n279_ = q2 & new_n278_;
  assign new_n280_ = ~j2 & ~new_n264_;
  assign new_n281_ = ~k2 & new_n280_;
  assign new_n282_ = ~new_n279_ & ~new_n281_;
  assign new_n283_ = ~new_n277_ & new_n282_;
  assign new_n284_ = ~y1 & a2;
  assign new_n285_ = ~e2 & f2;
  assign new_n286_ = d0 & new_n285_;
  assign new_n287_ = e2 & ~f2;
  assign new_n288_ = ~d0 & new_n287_;
  assign new_n289_ = ~new_n286_ & ~new_n288_;
  assign new_n290_ = new_n284_ & ~new_n289_;
  assign new_n291_ = m0 & new_n290_;
  assign new_n292_ = new_n259_ & new_n265_;
  assign new_n293_ = x1 & new_n292_;
  assign new_n294_ = ~new_n291_ & ~new_n293_;
  assign new_n295_ = new_n262_ & ~new_n264_;
  assign new_n296_ = new_n260_ & new_n295_;
  assign new_n297_ = new_n265_ & new_n283_;
  assign new_n298_ = ~x1 & new_n297_;
  assign new_n299_ = ~new_n296_ & ~new_n298_;
  assign k4 = ~new_n294_ | ~new_n299_;
  assign new_n301_ = g2 & h2;
  assign new_n302_ = ~c2 & ~new_n301_;
  assign l4 = ~n0 & ~new_n302_;
  assign new_n304_ = i & ~r;
  assign new_n305_ = r0 & ~new_n304_;
  assign new_n306_ = ~j & ~new_n305_;
  assign new_n307_ = ~r0 & ~new_n304_;
  assign new_n308_ = ~new_n306_ & ~new_n307_;
  assign m4 = ~y1 & new_n308_;
  assign new_n310_ = s0 & ~new_n304_;
  assign new_n311_ = ~k & ~new_n310_;
  assign new_n312_ = ~s0 & ~new_n304_;
  assign new_n313_ = ~new_n311_ & ~new_n312_;
  assign n4 = ~y1 & new_n313_;
  assign new_n315_ = t0 & ~new_n304_;
  assign new_n316_ = ~l & ~new_n315_;
  assign new_n317_ = ~t0 & ~new_n304_;
  assign new_n318_ = ~new_n316_ & ~new_n317_;
  assign o4 = ~y1 & new_n318_;
  assign new_n320_ = u0 & ~new_n304_;
  assign new_n321_ = ~m & ~new_n320_;
  assign new_n322_ = ~u0 & ~new_n304_;
  assign new_n323_ = ~new_n321_ & ~new_n322_;
  assign p4 = ~y1 & new_n323_;
  assign new_n325_ = v0 & ~new_n304_;
  assign new_n326_ = ~n & ~new_n325_;
  assign new_n327_ = ~v0 & ~new_n304_;
  assign new_n328_ = ~new_n326_ & ~new_n327_;
  assign q4 = ~y1 & new_n328_;
  assign new_n330_ = w0 & ~new_n304_;
  assign new_n331_ = ~o & ~new_n330_;
  assign new_n332_ = ~w0 & ~new_n304_;
  assign new_n333_ = ~new_n331_ & ~new_n332_;
  assign r4 = ~y1 & new_n333_;
  assign new_n335_ = x0 & ~new_n304_;
  assign new_n336_ = ~p & ~new_n335_;
  assign new_n337_ = ~x0 & ~new_n304_;
  assign new_n338_ = ~new_n336_ & ~new_n337_;
  assign s4 = ~y1 & new_n338_;
  assign new_n340_ = y0 & ~new_n304_;
  assign new_n341_ = ~q & ~new_n340_;
  assign new_n342_ = ~y0 & ~new_n304_;
  assign new_n343_ = ~new_n341_ & ~new_n342_;
  assign t4 = ~y1 & new_n343_;
  assign new_n345_ = i & r;
  assign new_n346_ = z0 & ~new_n345_;
  assign new_n347_ = ~j & ~new_n346_;
  assign new_n348_ = ~z0 & ~new_n345_;
  assign new_n349_ = ~new_n347_ & ~new_n348_;
  assign u4 = ~y1 & new_n349_;
  assign new_n351_ = a1 & ~new_n345_;
  assign new_n352_ = ~k & ~new_n351_;
  assign new_n353_ = ~a1 & ~new_n345_;
  assign new_n354_ = ~new_n352_ & ~new_n353_;
  assign v4 = ~y1 & new_n354_;
  assign new_n356_ = b1 & ~new_n345_;
  assign new_n357_ = ~l & ~new_n356_;
  assign new_n358_ = ~b1 & ~new_n345_;
  assign new_n359_ = ~new_n357_ & ~new_n358_;
  assign w4 = ~y1 & new_n359_;
  assign new_n361_ = c1 & ~new_n345_;
  assign new_n362_ = ~m & ~new_n361_;
  assign new_n363_ = ~c1 & ~new_n345_;
  assign new_n364_ = ~new_n362_ & ~new_n363_;
  assign x4 = ~y1 & new_n364_;
  assign new_n366_ = d1 & ~new_n345_;
  assign new_n367_ = ~n & ~new_n366_;
  assign new_n368_ = ~d1 & ~new_n345_;
  assign new_n369_ = ~new_n367_ & ~new_n368_;
  assign y4 = ~y1 & new_n369_;
  assign new_n371_ = e1 & ~new_n345_;
  assign new_n372_ = ~o & ~new_n371_;
  assign new_n373_ = ~e1 & ~new_n345_;
  assign new_n374_ = ~new_n372_ & ~new_n373_;
  assign z4 = ~y1 & new_n374_;
  assign new_n376_ = f1 & ~new_n345_;
  assign new_n377_ = ~p & ~new_n376_;
  assign new_n378_ = ~f1 & ~new_n345_;
  assign new_n379_ = ~new_n377_ & ~new_n378_;
  assign a5 = ~y1 & new_n379_;
  assign new_n381_ = g1 & ~new_n345_;
  assign new_n382_ = ~q & ~new_n381_;
  assign new_n383_ = ~g1 & ~new_n345_;
  assign new_n384_ = ~new_n382_ & ~new_n383_;
  assign b5 = ~y1 & new_n384_;
  assign new_n386_ = s & ~b0;
  assign new_n387_ = h1 & ~new_n386_;
  assign new_n388_ = ~t & ~new_n387_;
  assign new_n389_ = ~h1 & ~new_n386_;
  assign new_n390_ = ~new_n388_ & ~new_n389_;
  assign c5 = ~y1 & new_n390_;
  assign new_n392_ = i1 & ~new_n386_;
  assign new_n393_ = ~u & ~new_n392_;
  assign new_n394_ = ~i1 & ~new_n386_;
  assign new_n395_ = ~new_n393_ & ~new_n394_;
  assign d5 = ~y1 & new_n395_;
  assign new_n397_ = j1 & ~new_n386_;
  assign new_n398_ = ~v & ~new_n397_;
  assign new_n399_ = ~j1 & ~new_n386_;
  assign new_n400_ = ~new_n398_ & ~new_n399_;
  assign e5 = ~y1 & new_n400_;
  assign new_n402_ = k1 & ~new_n386_;
  assign new_n403_ = ~w & ~new_n402_;
  assign new_n404_ = ~k1 & ~new_n386_;
  assign new_n405_ = ~new_n403_ & ~new_n404_;
  assign f5 = ~y1 & new_n405_;
  assign new_n407_ = l1 & ~new_n386_;
  assign new_n408_ = ~x & ~new_n407_;
  assign new_n409_ = ~l1 & ~new_n386_;
  assign new_n410_ = ~new_n408_ & ~new_n409_;
  assign g5 = ~y1 & new_n410_;
  assign new_n412_ = m1 & ~new_n386_;
  assign new_n413_ = ~y & ~new_n412_;
  assign new_n414_ = ~m1 & ~new_n386_;
  assign new_n415_ = ~new_n413_ & ~new_n414_;
  assign h5 = ~y1 & new_n415_;
  assign new_n417_ = n1 & ~new_n386_;
  assign new_n418_ = ~z & ~new_n417_;
  assign new_n419_ = ~n1 & ~new_n386_;
  assign new_n420_ = ~new_n418_ & ~new_n419_;
  assign i5 = ~y1 & new_n420_;
  assign new_n422_ = o1 & ~new_n386_;
  assign new_n423_ = ~a0 & ~new_n422_;
  assign new_n424_ = ~o1 & ~new_n386_;
  assign new_n425_ = ~new_n423_ & ~new_n424_;
  assign j5 = ~y1 & new_n425_;
  assign new_n427_ = s & b0;
  assign new_n428_ = p1 & ~new_n427_;
  assign new_n429_ = ~t & ~new_n428_;
  assign new_n430_ = ~p1 & ~new_n427_;
  assign new_n431_ = ~new_n429_ & ~new_n430_;
  assign k5 = ~y1 & new_n431_;
  assign new_n433_ = q1 & ~new_n427_;
  assign new_n434_ = ~u & ~new_n433_;
  assign new_n435_ = ~q1 & ~new_n427_;
  assign new_n436_ = ~new_n434_ & ~new_n435_;
  assign l5 = ~y1 & new_n436_;
  assign new_n438_ = r1 & ~new_n427_;
  assign new_n439_ = ~v & ~new_n438_;
  assign new_n440_ = ~r1 & ~new_n427_;
  assign new_n441_ = ~new_n439_ & ~new_n440_;
  assign m5 = ~y1 & new_n441_;
  assign new_n443_ = s1 & ~new_n427_;
  assign new_n444_ = ~w & ~new_n443_;
  assign new_n445_ = ~s1 & ~new_n427_;
  assign new_n446_ = ~new_n444_ & ~new_n445_;
  assign n5 = ~y1 & new_n446_;
  assign new_n448_ = t1 & ~new_n427_;
  assign new_n449_ = ~x & ~new_n448_;
  assign new_n450_ = ~t1 & ~new_n427_;
  assign new_n451_ = ~new_n449_ & ~new_n450_;
  assign o5 = ~y1 & new_n451_;
  assign new_n453_ = u1 & ~new_n427_;
  assign new_n454_ = ~y & ~new_n453_;
  assign new_n455_ = ~u1 & ~new_n427_;
  assign new_n456_ = ~new_n454_ & ~new_n455_;
  assign p5 = ~y1 & new_n456_;
  assign new_n458_ = v1 & ~new_n427_;
  assign new_n459_ = ~z & ~new_n458_;
  assign new_n460_ = ~v1 & ~new_n427_;
  assign new_n461_ = ~new_n459_ & ~new_n460_;
  assign q5 = ~y1 & new_n461_;
  assign new_n463_ = w1 & ~new_n427_;
  assign new_n464_ = ~a0 & ~new_n463_;
  assign new_n465_ = ~w1 & ~new_n427_;
  assign new_n466_ = ~new_n464_ & ~new_n465_;
  assign r5 = ~y1 & new_n466_;
  assign new_n468_ = ~e & x1;
  assign new_n469_ = ~c & new_n468_;
  assign new_n470_ = ~d & new_n469_;
  assign s5 = y1 | new_n470_;
  assign t5 = n0 | new_n239_;
  assign new_n473_ = ~y1 & ~z1;
  assign new_n474_ = ~c0 & q2;
  assign new_n475_ = ~new_n271_ & ~new_n474_;
  assign new_n476_ = i2 & ~new_n475_;
  assign new_n477_ = ~i2 & ~new_n261_;
  assign new_n478_ = i3 & new_n477_;
  assign new_n479_ = ~new_n476_ & ~new_n478_;
  assign new_n480_ = new_n261_ & ~new_n264_;
  assign new_n481_ = new_n259_ & new_n480_;
  assign new_n482_ = ~new_n261_ & new_n276_;
  assign new_n483_ = ~q2 & new_n482_;
  assign new_n484_ = ~new_n481_ & ~new_n483_;
  assign new_n485_ = new_n479_ & new_n484_;
  assign new_n486_ = ~r2 & ~i3;
  assign new_n487_ = c0 & q2;
  assign new_n488_ = ~d0 & r2;
  assign new_n489_ = ~new_n487_ & ~new_n488_;
  assign new_n490_ = i2 & ~new_n489_;
  assign new_n491_ = ~x1 & ~new_n490_;
  assign new_n492_ = ~i3 & new_n477_;
  assign new_n493_ = new_n491_ & ~new_n492_;
  assign new_n494_ = ~new_n259_ & new_n480_;
  assign new_n495_ = ~new_n261_ & new_n486_;
  assign new_n496_ = ~q2 & new_n495_;
  assign new_n497_ = ~new_n494_ & ~new_n496_;
  assign new_n498_ = new_n493_ & new_n497_;
  assign new_n499_ = ~y1 & i2;
  assign new_n500_ = ~x1 & new_n499_;
  assign new_n501_ = new_n237_ & new_n500_;
  assign new_n502_ = new_n473_ & ~new_n485_;
  assign new_n503_ = ~x1 & new_n502_;
  assign new_n504_ = ~y1 & ~new_n498_;
  assign new_n505_ = z1 & new_n504_;
  assign new_n506_ = ~new_n503_ & ~new_n505_;
  assign u5 = new_n501_ | ~new_n506_;
  assign new_n508_ = ~i0 & ~j0;
  assign new_n509_ = l0 & d2;
  assign new_n510_ = ~k0 & new_n509_;
  assign new_n511_ = j0 & ~f4;
  assign new_n512_ = ~k0 & ~g4;
  assign new_n513_ = k0 & g4;
  assign new_n514_ = ~new_n512_ & ~new_n513_;
  assign new_n515_ = ~new_n511_ & ~new_n514_;
  assign new_n516_ = i0 & ~e4;
  assign new_n517_ = ~j0 & f4;
  assign new_n518_ = ~new_n516_ & ~new_n517_;
  assign new_n519_ = new_n515_ & new_n518_;
  assign new_n520_ = h0 & d4;
  assign new_n521_ = ~i0 & e4;
  assign new_n522_ = ~new_n520_ & ~new_n521_;
  assign new_n523_ = new_n519_ & new_n522_;
  assign new_n524_ = ~h0 & ~d4;
  assign new_n525_ = c4 & ~new_n524_;
  assign new_n526_ = new_n523_ & new_n525_;
  assign new_n527_ = a4 & b4;
  assign new_n528_ = new_n526_ & new_n527_;
  assign new_n529_ = y3 & z3;
  assign new_n530_ = new_n528_ & new_n529_;
  assign new_n531_ = h4 & new_n530_;
  assign new_n532_ = e2 & f2;
  assign new_n533_ = a2 & ~new_n532_;
  assign new_n534_ = ~new_n531_ & ~new_n533_;
  assign new_n535_ = new_n508_ & new_n510_;
  assign new_n536_ = ~h0 & new_n535_;
  assign new_n537_ = new_n534_ & ~new_n536_;
  assign v5 = ~y1 & ~new_n537_;
  assign new_n539_ = ~f4 & ~g4;
  assign new_n540_ = b2 & y3;
  assign new_n541_ = new_n539_ & new_n540_;
  assign new_n542_ = z3 & new_n527_;
  assign new_n543_ = d4 & ~e4;
  assign new_n544_ = c4 & new_n543_;
  assign new_n545_ = z3 & a4;
  assign new_n546_ = y3 & new_n545_;
  assign new_n547_ = c4 & d4;
  assign new_n548_ = b4 & new_n547_;
  assign new_n549_ = ~e4 & new_n539_;
  assign new_n550_ = new_n546_ & new_n548_;
  assign new_n551_ = new_n549_ & new_n550_;
  assign new_n552_ = ~l0 & ~n0;
  assign new_n553_ = ~b2 & ~new_n551_;
  assign new_n554_ = new_n542_ & new_n544_;
  assign new_n555_ = new_n541_ & new_n554_;
  assign new_n556_ = ~new_n553_ & ~new_n555_;
  assign w5 = new_n552_ & new_n556_;
  assign new_n558_ = ~l0 & new_n548_;
  assign new_n559_ = new_n549_ & new_n558_;
  assign new_n560_ = b2 & ~c2;
  assign new_n561_ = ~n0 & new_n560_;
  assign new_n562_ = ~n0 & c2;
  assign new_n563_ = new_n541_ & new_n542_;
  assign new_n564_ = new_n544_ & new_n563_;
  assign new_n565_ = new_n546_ & new_n561_;
  assign new_n566_ = new_n559_ & new_n565_;
  assign new_n567_ = new_n562_ & ~new_n564_;
  assign new_n568_ = ~l0 & new_n567_;
  assign x5 = new_n566_ | new_n568_;
  assign new_n570_ = ~l0 & ~d2;
  assign new_n571_ = ~n0 & ~new_n570_;
  assign new_n572_ = b & new_n571_;
  assign y5 = ~new_n301_ & new_n572_;
  assign new_n574_ = ~a2 & e2;
  assign new_n575_ = ~new_n531_ & ~new_n536_;
  assign new_n576_ = ~a2 & new_n575_;
  assign new_n577_ = new_n574_ & new_n575_;
  assign new_n578_ = ~e2 & ~new_n576_;
  assign new_n579_ = ~new_n577_ & ~new_n578_;
  assign z5 = ~n0 & ~new_n579_;
  assign new_n581_ = ~a2 & f2;
  assign new_n582_ = ~a2 & ~new_n531_;
  assign new_n583_ = ~new_n536_ & new_n582_;
  assign new_n584_ = ~n0 & new_n285_;
  assign new_n585_ = new_n575_ & new_n581_;
  assign new_n586_ = new_n287_ & ~new_n583_;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = ~n0 & ~new_n587_;
  assign a6 = new_n584_ | new_n588_;
  assign b6 = ~n0 & h2;
  assign c6 = l0 & ~n0;
  assign new_n592_ = g0 & new_n254_;
  assign new_n593_ = ~m2 & ~new_n592_;
  assign new_n594_ = l2 & new_n593_;
  assign new_n595_ = n2 & new_n594_;
  assign new_n596_ = j2 & ~p2;
  assign new_n597_ = o2 & ~new_n596_;
  assign new_n598_ = new_n595_ & ~new_n597_;
  assign new_n599_ = ~x1 & new_n598_;
  assign new_n600_ = ~i2 & ~new_n599_;
  assign d6 = ~y1 & ~new_n600_;
  assign new_n602_ = ~j2 & o2;
  assign new_n603_ = ~m2 & ~new_n602_;
  assign new_n604_ = l2 & new_n603_;
  assign new_n605_ = ~e0 & ~f0;
  assign new_n606_ = ~o2 & new_n605_;
  assign new_n607_ = n2 & ~new_n606_;
  assign new_n608_ = new_n604_ & new_n607_;
  assign new_n609_ = ~g0 & ~o2;
  assign new_n610_ = new_n608_ & ~new_n609_;
  assign new_n611_ = ~p2 & new_n610_;
  assign new_n612_ = ~j2 & ~new_n611_;
  assign new_n613_ = j2 & new_n611_;
  assign new_n614_ = ~x1 & new_n613_;
  assign new_n615_ = ~new_n612_ & ~new_n614_;
  assign new_n616_ = ~y1 & new_n615_;
  assign new_n617_ = x1 & ~j2;
  assign e6 = new_n616_ & ~new_n617_;
  assign new_n619_ = ~f0 & g0;
  assign new_n620_ = ~e0 & new_n619_;
  assign new_n621_ = ~m2 & n2;
  assign new_n622_ = l2 & new_n621_;
  assign new_n623_ = ~p2 & ~new_n620_;
  assign new_n624_ = new_n622_ & ~new_n623_;
  assign new_n625_ = ~o2 & new_n624_;
  assign new_n626_ = ~k2 & ~new_n625_;
  assign new_n627_ = k2 & new_n625_;
  assign new_n628_ = ~x1 & new_n627_;
  assign new_n629_ = ~new_n626_ & ~new_n628_;
  assign new_n630_ = ~y1 & new_n629_;
  assign new_n631_ = x1 & ~k2;
  assign f6 = new_n630_ & ~new_n631_;
  assign new_n633_ = ~c & ~d;
  assign new_n634_ = new_n468_ & new_n633_;
  assign new_n635_ = ~c & new_n236_;
  assign new_n636_ = x1 & ~l2;
  assign new_n637_ = new_n635_ & new_n636_;
  assign new_n638_ = l2 & ~new_n634_;
  assign new_n639_ = ~new_n637_ & ~new_n638_;
  assign g6 = ~y1 & new_n639_;
  assign new_n641_ = x1 & ~m2;
  assign new_n642_ = ~e & new_n641_;
  assign new_n643_ = ~c & new_n642_;
  assign new_n644_ = ~d & new_n643_;
  assign new_n645_ = ~y1 & ~new_n644_;
  assign new_n646_ = m2 & ~new_n634_;
  assign new_n647_ = l2 & ~new_n646_;
  assign new_n648_ = m2 & ~new_n638_;
  assign new_n649_ = ~new_n647_ & ~new_n648_;
  assign h6 = new_n645_ & ~new_n649_;
  assign new_n651_ = m2 & n2;
  assign new_n652_ = l2 & m2;
  assign new_n653_ = ~new_n470_ & new_n652_;
  assign new_n654_ = ~n2 & ~new_n653_;
  assign new_n655_ = ~new_n634_ & new_n651_;
  assign new_n656_ = l2 & new_n655_;
  assign new_n657_ = ~new_n654_ & ~new_n656_;
  assign i6 = ~y1 & new_n657_;
  assign new_n659_ = n2 & o2;
  assign new_n660_ = m2 & new_n659_;
  assign new_n661_ = l2 & new_n651_;
  assign new_n662_ = ~new_n470_ & new_n661_;
  assign new_n663_ = ~o2 & ~new_n662_;
  assign new_n664_ = ~new_n634_ & new_n660_;
  assign new_n665_ = l2 & new_n664_;
  assign new_n666_ = ~new_n663_ & ~new_n665_;
  assign j6 = ~y1 & new_n666_;
  assign new_n668_ = o2 & p2;
  assign new_n669_ = n2 & new_n668_;
  assign new_n670_ = l2 & ~new_n470_;
  assign new_n671_ = new_n660_ & new_n670_;
  assign new_n672_ = ~p2 & ~new_n671_;
  assign new_n673_ = ~new_n634_ & new_n669_;
  assign new_n674_ = new_n652_ & new_n673_;
  assign new_n675_ = ~new_n672_ & ~new_n674_;
  assign k6 = ~y1 & new_n675_;
  assign new_n677_ = ~i2 & ~new_n598_;
  assign new_n678_ = ~x1 & ~new_n677_;
  assign new_n679_ = ~q2 & ~new_n678_;
  assign new_n680_ = ~y1 & ~new_n679_;
  assign new_n681_ = q2 & new_n678_;
  assign l6 = new_n680_ & ~new_n681_;
  assign new_n683_ = ~r2 & ~new_n681_;
  assign new_n684_ = new_n237_ & ~new_n677_;
  assign new_n685_ = ~x1 & new_n684_;
  assign new_n686_ = ~new_n683_ & ~new_n685_;
  assign m6 = ~y1 & new_n686_;
  assign new_n688_ = ~f & ~s2;
  assign new_n689_ = ~h & ~t2;
  assign new_n690_ = f & new_n689_;
  assign new_n691_ = ~new_n688_ & ~new_n690_;
  assign new_n692_ = ~y1 & new_n691_;
  assign new_n693_ = h & ~s2;
  assign n6 = new_n692_ & ~new_n693_;
  assign new_n695_ = ~f & ~t2;
  assign new_n696_ = ~h & ~u2;
  assign new_n697_ = f & new_n696_;
  assign new_n698_ = ~new_n695_ & ~new_n697_;
  assign new_n699_ = ~y1 & new_n698_;
  assign new_n700_ = h & ~t2;
  assign o6 = new_n699_ & ~new_n700_;
  assign new_n702_ = ~f & ~u2;
  assign new_n703_ = ~h & ~v2;
  assign new_n704_ = f & new_n703_;
  assign new_n705_ = ~new_n702_ & ~new_n704_;
  assign new_n706_ = ~y1 & new_n705_;
  assign new_n707_ = h & ~u2;
  assign p6 = new_n706_ & ~new_n707_;
  assign new_n709_ = ~f & ~v2;
  assign new_n710_ = ~h & ~w2;
  assign new_n711_ = f & new_n710_;
  assign new_n712_ = ~new_n709_ & ~new_n711_;
  assign new_n713_ = ~y1 & new_n712_;
  assign new_n714_ = h & ~v2;
  assign q6 = new_n713_ & ~new_n714_;
  assign new_n716_ = ~f & ~w2;
  assign new_n717_ = ~h & ~x2;
  assign new_n718_ = f & new_n717_;
  assign new_n719_ = ~new_n716_ & ~new_n718_;
  assign new_n720_ = ~y1 & new_n719_;
  assign new_n721_ = h & ~w2;
  assign r6 = new_n720_ & ~new_n721_;
  assign new_n723_ = ~f & ~x2;
  assign new_n724_ = ~h & ~y2;
  assign new_n725_ = f & new_n724_;
  assign new_n726_ = ~new_n723_ & ~new_n725_;
  assign new_n727_ = ~y1 & new_n726_;
  assign new_n728_ = h & ~x2;
  assign s6 = new_n727_ & ~new_n728_;
  assign new_n730_ = ~f & ~y2;
  assign new_n731_ = ~h & ~z2;
  assign new_n732_ = f & new_n731_;
  assign new_n733_ = ~new_n730_ & ~new_n732_;
  assign new_n734_ = ~y1 & new_n733_;
  assign new_n735_ = h & ~y2;
  assign t6 = new_n734_ & ~new_n735_;
  assign new_n737_ = ~g & ~h;
  assign new_n738_ = f & new_n737_;
  assign new_n739_ = ~f & ~z2;
  assign new_n740_ = ~new_n738_ & ~new_n739_;
  assign new_n741_ = ~y1 & new_n740_;
  assign new_n742_ = h & ~z2;
  assign u6 = new_n741_ & ~new_n742_;
  assign new_n744_ = ~f & ~a3;
  assign new_n745_ = h & ~b3;
  assign new_n746_ = f & new_n745_;
  assign new_n747_ = ~new_n744_ & ~new_n746_;
  assign new_n748_ = ~y1 & new_n747_;
  assign new_n749_ = ~h & ~a3;
  assign v6 = new_n748_ & ~new_n749_;
  assign new_n751_ = ~f & ~b3;
  assign new_n752_ = h & ~c3;
  assign new_n753_ = f & new_n752_;
  assign new_n754_ = ~new_n751_ & ~new_n753_;
  assign new_n755_ = ~y1 & new_n754_;
  assign new_n756_ = ~h & ~b3;
  assign w6 = new_n755_ & ~new_n756_;
  assign new_n758_ = ~f & ~c3;
  assign new_n759_ = h & ~d3;
  assign new_n760_ = f & new_n759_;
  assign new_n761_ = ~new_n758_ & ~new_n760_;
  assign new_n762_ = ~y1 & new_n761_;
  assign new_n763_ = ~h & ~c3;
  assign x6 = new_n762_ & ~new_n763_;
  assign new_n765_ = ~f & ~d3;
  assign new_n766_ = h & ~e3;
  assign new_n767_ = f & new_n766_;
  assign new_n768_ = ~new_n765_ & ~new_n767_;
  assign new_n769_ = ~y1 & new_n768_;
  assign new_n770_ = ~h & ~d3;
  assign y6 = new_n769_ & ~new_n770_;
  assign new_n772_ = ~f & ~e3;
  assign new_n773_ = h & ~f3;
  assign new_n774_ = f & new_n773_;
  assign new_n775_ = ~new_n772_ & ~new_n774_;
  assign new_n776_ = ~y1 & new_n775_;
  assign new_n777_ = ~h & ~e3;
  assign z6 = new_n776_ & ~new_n777_;
  assign new_n779_ = ~f & ~f3;
  assign new_n780_ = h & ~g3;
  assign new_n781_ = f & new_n780_;
  assign new_n782_ = ~new_n779_ & ~new_n781_;
  assign new_n783_ = ~y1 & new_n782_;
  assign new_n784_ = ~h & ~f3;
  assign a7 = new_n783_ & ~new_n784_;
  assign new_n786_ = ~f & ~g3;
  assign new_n787_ = h & ~h3;
  assign new_n788_ = f & new_n787_;
  assign new_n789_ = ~new_n786_ & ~new_n788_;
  assign new_n790_ = ~y1 & new_n789_;
  assign new_n791_ = ~h & ~g3;
  assign b7 = new_n790_ & ~new_n791_;
  assign new_n793_ = ~f & ~h3;
  assign new_n794_ = ~g & h;
  assign new_n795_ = f & new_n794_;
  assign new_n796_ = ~new_n793_ & ~new_n795_;
  assign new_n797_ = ~y1 & new_n796_;
  assign new_n798_ = ~h & ~h3;
  assign c7 = new_n797_ & ~new_n798_;
  assign new_n800_ = ~x1 & ~new_n261_;
  assign new_n801_ = i3 & ~new_n800_;
  assign new_n802_ = j3 & new_n800_;
  assign new_n803_ = ~new_n801_ & ~new_n802_;
  assign new_n804_ = c & new_n236_;
  assign new_n805_ = ~s2 & new_n804_;
  assign new_n806_ = ~e & ~r0;
  assign new_n807_ = d & new_n806_;
  assign new_n808_ = e & ~h1;
  assign new_n809_ = ~new_n807_ & ~new_n808_;
  assign new_n810_ = ~new_n805_ & new_n809_;
  assign new_n811_ = new_n236_ & new_n803_;
  assign new_n812_ = ~c & new_n811_;
  assign new_n813_ = new_n810_ & ~new_n812_;
  assign d7 = ~y1 & new_n813_;
  assign new_n815_ = j3 & ~new_n800_;
  assign new_n816_ = k3 & new_n800_;
  assign new_n817_ = ~new_n815_ & ~new_n816_;
  assign new_n818_ = ~t2 & new_n804_;
  assign new_n819_ = ~e & ~s0;
  assign new_n820_ = d & new_n819_;
  assign new_n821_ = e & ~i1;
  assign new_n822_ = ~new_n820_ & ~new_n821_;
  assign new_n823_ = ~new_n818_ & new_n822_;
  assign new_n824_ = new_n236_ & new_n817_;
  assign new_n825_ = ~c & new_n824_;
  assign new_n826_ = new_n823_ & ~new_n825_;
  assign e7 = ~y1 & new_n826_;
  assign new_n828_ = k3 & ~new_n800_;
  assign new_n829_ = l3 & new_n800_;
  assign new_n830_ = ~new_n828_ & ~new_n829_;
  assign new_n831_ = ~u2 & new_n804_;
  assign new_n832_ = ~e & ~t0;
  assign new_n833_ = d & new_n832_;
  assign new_n834_ = e & ~j1;
  assign new_n835_ = ~new_n833_ & ~new_n834_;
  assign new_n836_ = ~new_n831_ & new_n835_;
  assign new_n837_ = new_n236_ & new_n830_;
  assign new_n838_ = ~c & new_n837_;
  assign new_n839_ = new_n836_ & ~new_n838_;
  assign f7 = ~y1 & new_n839_;
  assign new_n841_ = l3 & ~new_n800_;
  assign new_n842_ = m3 & new_n800_;
  assign new_n843_ = ~new_n841_ & ~new_n842_;
  assign new_n844_ = ~v2 & new_n804_;
  assign new_n845_ = ~e & ~u0;
  assign new_n846_ = d & new_n845_;
  assign new_n847_ = e & ~k1;
  assign new_n848_ = ~new_n846_ & ~new_n847_;
  assign new_n849_ = ~new_n844_ & new_n848_;
  assign new_n850_ = new_n236_ & new_n843_;
  assign new_n851_ = ~c & new_n850_;
  assign new_n852_ = new_n849_ & ~new_n851_;
  assign g7 = ~y1 & new_n852_;
  assign new_n854_ = m3 & ~new_n800_;
  assign new_n855_ = n3 & new_n800_;
  assign new_n856_ = ~new_n854_ & ~new_n855_;
  assign new_n857_ = ~w2 & new_n804_;
  assign new_n858_ = ~e & ~v0;
  assign new_n859_ = d & new_n858_;
  assign new_n860_ = e & ~l1;
  assign new_n861_ = ~new_n859_ & ~new_n860_;
  assign new_n862_ = ~new_n857_ & new_n861_;
  assign new_n863_ = new_n236_ & new_n856_;
  assign new_n864_ = ~c & new_n863_;
  assign new_n865_ = new_n862_ & ~new_n864_;
  assign h7 = ~y1 & new_n865_;
  assign new_n867_ = n3 & ~new_n800_;
  assign new_n868_ = o3 & new_n800_;
  assign new_n869_ = ~new_n867_ & ~new_n868_;
  assign new_n870_ = ~x2 & new_n804_;
  assign new_n871_ = ~e & ~w0;
  assign new_n872_ = d & new_n871_;
  assign new_n873_ = e & ~m1;
  assign new_n874_ = ~new_n872_ & ~new_n873_;
  assign new_n875_ = ~new_n870_ & new_n874_;
  assign new_n876_ = new_n236_ & new_n869_;
  assign new_n877_ = ~c & new_n876_;
  assign new_n878_ = new_n875_ & ~new_n877_;
  assign i7 = ~y1 & new_n878_;
  assign new_n880_ = o3 & ~new_n800_;
  assign new_n881_ = p3 & new_n800_;
  assign new_n882_ = ~new_n880_ & ~new_n881_;
  assign new_n883_ = ~y2 & new_n804_;
  assign new_n884_ = ~e & ~x0;
  assign new_n885_ = d & new_n884_;
  assign new_n886_ = e & ~n1;
  assign new_n887_ = ~new_n885_ & ~new_n886_;
  assign new_n888_ = ~new_n883_ & new_n887_;
  assign new_n889_ = new_n236_ & new_n882_;
  assign new_n890_ = ~c & new_n889_;
  assign new_n891_ = new_n888_ & ~new_n890_;
  assign j7 = ~y1 & new_n891_;
  assign new_n893_ = p3 & ~new_n800_;
  assign new_n894_ = q3 & new_n800_;
  assign new_n895_ = ~new_n893_ & ~new_n894_;
  assign new_n896_ = ~z2 & new_n804_;
  assign new_n897_ = ~e & ~y0;
  assign new_n898_ = d & new_n897_;
  assign new_n899_ = e & ~o1;
  assign new_n900_ = ~new_n898_ & ~new_n899_;
  assign new_n901_ = ~new_n896_ & new_n900_;
  assign new_n902_ = new_n236_ & new_n895_;
  assign new_n903_ = ~c & new_n902_;
  assign new_n904_ = new_n901_ & ~new_n903_;
  assign k7 = ~y1 & new_n904_;
  assign new_n906_ = q3 & ~new_n800_;
  assign new_n907_ = r3 & new_n800_;
  assign new_n908_ = ~new_n906_ & ~new_n907_;
  assign new_n909_ = ~a3 & new_n804_;
  assign new_n910_ = ~e & ~z0;
  assign new_n911_ = d & new_n910_;
  assign new_n912_ = e & ~p1;
  assign new_n913_ = ~new_n911_ & ~new_n912_;
  assign new_n914_ = ~new_n909_ & new_n913_;
  assign new_n915_ = new_n236_ & new_n908_;
  assign new_n916_ = ~c & new_n915_;
  assign new_n917_ = new_n914_ & ~new_n916_;
  assign l7 = ~y1 & new_n917_;
  assign new_n919_ = r3 & ~new_n800_;
  assign new_n920_ = s3 & new_n800_;
  assign new_n921_ = ~new_n919_ & ~new_n920_;
  assign new_n922_ = ~b3 & new_n804_;
  assign new_n923_ = ~e & ~a1;
  assign new_n924_ = d & new_n923_;
  assign new_n925_ = e & ~q1;
  assign new_n926_ = ~new_n924_ & ~new_n925_;
  assign new_n927_ = ~new_n922_ & new_n926_;
  assign new_n928_ = new_n236_ & new_n921_;
  assign new_n929_ = ~c & new_n928_;
  assign new_n930_ = new_n927_ & ~new_n929_;
  assign m7 = ~y1 & new_n930_;
  assign new_n932_ = s3 & ~new_n800_;
  assign new_n933_ = t3 & new_n800_;
  assign new_n934_ = ~new_n932_ & ~new_n933_;
  assign new_n935_ = ~c3 & new_n804_;
  assign new_n936_ = ~e & ~b1;
  assign new_n937_ = d & new_n936_;
  assign new_n938_ = e & ~r1;
  assign new_n939_ = ~new_n937_ & ~new_n938_;
  assign new_n940_ = ~new_n935_ & new_n939_;
  assign new_n941_ = new_n236_ & new_n934_;
  assign new_n942_ = ~c & new_n941_;
  assign new_n943_ = new_n940_ & ~new_n942_;
  assign n7 = ~y1 & new_n943_;
  assign new_n945_ = t3 & ~new_n800_;
  assign new_n946_ = u3 & new_n800_;
  assign new_n947_ = ~new_n945_ & ~new_n946_;
  assign new_n948_ = ~d3 & new_n804_;
  assign new_n949_ = ~e & ~c1;
  assign new_n950_ = d & new_n949_;
  assign new_n951_ = e & ~s1;
  assign new_n952_ = ~new_n950_ & ~new_n951_;
  assign new_n953_ = ~new_n948_ & new_n952_;
  assign new_n954_ = new_n236_ & new_n947_;
  assign new_n955_ = ~c & new_n954_;
  assign new_n956_ = new_n953_ & ~new_n955_;
  assign o7 = ~y1 & new_n956_;
  assign new_n958_ = u3 & ~new_n800_;
  assign new_n959_ = v3 & new_n800_;
  assign new_n960_ = ~new_n958_ & ~new_n959_;
  assign new_n961_ = ~e3 & new_n804_;
  assign new_n962_ = ~e & ~d1;
  assign new_n963_ = d & new_n962_;
  assign new_n964_ = e & ~t1;
  assign new_n965_ = ~new_n963_ & ~new_n964_;
  assign new_n966_ = ~new_n961_ & new_n965_;
  assign new_n967_ = new_n236_ & new_n960_;
  assign new_n968_ = ~c & new_n967_;
  assign new_n969_ = new_n966_ & ~new_n968_;
  assign p7 = ~y1 & new_n969_;
  assign new_n971_ = v3 & ~new_n800_;
  assign new_n972_ = w3 & new_n800_;
  assign new_n973_ = ~new_n971_ & ~new_n972_;
  assign new_n974_ = ~f3 & new_n804_;
  assign new_n975_ = ~e & ~e1;
  assign new_n976_ = d & new_n975_;
  assign new_n977_ = e & ~u1;
  assign new_n978_ = ~new_n976_ & ~new_n977_;
  assign new_n979_ = ~new_n974_ & new_n978_;
  assign new_n980_ = new_n236_ & new_n973_;
  assign new_n981_ = ~c & new_n980_;
  assign new_n982_ = new_n979_ & ~new_n981_;
  assign q7 = ~y1 & new_n982_;
  assign new_n984_ = w3 & ~new_n800_;
  assign new_n985_ = x3 & new_n800_;
  assign new_n986_ = ~new_n984_ & ~new_n985_;
  assign new_n987_ = ~g3 & new_n804_;
  assign new_n988_ = ~e & ~f1;
  assign new_n989_ = d & new_n988_;
  assign new_n990_ = e & ~v1;
  assign new_n991_ = ~new_n989_ & ~new_n990_;
  assign new_n992_ = ~new_n987_ & new_n991_;
  assign new_n993_ = new_n236_ & new_n986_;
  assign new_n994_ = ~c & new_n993_;
  assign new_n995_ = new_n992_ & ~new_n994_;
  assign r7 = ~y1 & new_n995_;
  assign new_n997_ = x3 & ~new_n800_;
  assign new_n998_ = ~h3 & new_n804_;
  assign new_n999_ = ~e & ~g1;
  assign new_n1000_ = d & new_n999_;
  assign new_n1001_ = e & ~w1;
  assign new_n1002_ = ~new_n1000_ & ~new_n1001_;
  assign new_n1003_ = ~new_n998_ & new_n1002_;
  assign new_n1004_ = new_n236_ & ~new_n997_;
  assign new_n1005_ = ~c & new_n1004_;
  assign new_n1006_ = new_n1003_ & ~new_n1005_;
  assign s7 = ~y1 & new_n1006_;
  assign new_n1008_ = ~n0 & ~y3;
  assign t7 = ~l0 & new_n1008_;
  assign new_n1010_ = ~n0 & ~new_n529_;
  assign new_n1011_ = ~l0 & new_n1010_;
  assign new_n1012_ = ~y3 & ~z3;
  assign u7 = new_n1011_ & ~new_n1012_;
  assign new_n1014_ = ~n0 & ~new_n546_;
  assign new_n1015_ = ~l0 & new_n1014_;
  assign new_n1016_ = ~a4 & ~new_n529_;
  assign v7 = new_n1015_ & ~new_n1016_;
  assign new_n1018_ = ~b4 & ~new_n546_;
  assign new_n1019_ = y3 & new_n527_;
  assign new_n1020_ = z3 & new_n1019_;
  assign new_n1021_ = ~new_n1018_ & ~new_n1020_;
  assign w7 = new_n552_ & new_n1021_;
  assign new_n1023_ = b4 & c4;
  assign new_n1024_ = a4 & new_n1023_;
  assign new_n1025_ = new_n527_ & new_n529_;
  assign new_n1026_ = ~c4 & ~new_n1025_;
  assign new_n1027_ = y3 & new_n1024_;
  assign new_n1028_ = z3 & new_n1027_;
  assign new_n1029_ = ~new_n1026_ & ~new_n1028_;
  assign x7 = new_n552_ & new_n1029_;
  assign new_n1031_ = new_n529_ & new_n1024_;
  assign new_n1032_ = ~d4 & ~new_n1031_;
  assign new_n1033_ = new_n545_ & new_n548_;
  assign new_n1034_ = y3 & new_n1033_;
  assign new_n1035_ = ~new_n1032_ & ~new_n1034_;
  assign y7 = new_n552_ & new_n1035_;
  assign new_n1037_ = ~d4 & e4;
  assign new_n1038_ = c4 & new_n1037_;
  assign new_n1039_ = c4 & ~d4;
  assign new_n1040_ = b4 & new_n1039_;
  assign new_n1041_ = new_n546_ & new_n1040_;
  assign new_n1042_ = ~e4 & ~new_n1041_;
  assign new_n1043_ = new_n542_ & new_n1038_;
  assign new_n1044_ = y3 & new_n1043_;
  assign new_n1045_ = ~new_n1042_ & ~new_n1044_;
  assign z7 = new_n552_ & new_n1045_;
  assign new_n1047_ = e4 & f4;
  assign new_n1048_ = ~d4 & new_n1047_;
  assign new_n1049_ = y3 & new_n542_;
  assign new_n1050_ = new_n1038_ & new_n1049_;
  assign new_n1051_ = ~f4 & ~new_n1050_;
  assign new_n1052_ = new_n1024_ & new_n1048_;
  assign new_n1053_ = new_n529_ & new_n1052_;
  assign new_n1054_ = ~new_n1051_ & ~new_n1053_;
  assign a8 = new_n552_ & new_n1054_;
  assign new_n1056_ = f4 & g4;
  assign new_n1057_ = e4 & new_n1056_;
  assign new_n1058_ = new_n1031_ & new_n1048_;
  assign new_n1059_ = ~g4 & ~new_n1058_;
  assign new_n1060_ = new_n1040_ & new_n1057_;
  assign new_n1061_ = new_n546_ & new_n1060_;
  assign new_n1062_ = ~new_n1059_ & ~new_n1061_;
  assign b8 = new_n552_ & new_n1062_;
  assign new_n1064_ = ~n0 & ~new_n301_;
  assign new_n1065_ = b & new_n1064_;
  assign new_n1066_ = ~h4 & ~new_n509_;
  assign c8 = new_n1065_ & ~new_n1066_;
endmodule


