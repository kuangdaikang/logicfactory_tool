// Benchmark "log2" written by ABC on Thu Sep 14 20:18:57 2023

module log2 ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] ;
  wire new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n120_, new_n121_, new_n122_, new_n123_,
    new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_,
    new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_,
    new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1883_, new_n1884_, new_n1885_,
    new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_,
    new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_,
    new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_,
    new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_,
    new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_,
    new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_,
    new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_,
    new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_,
    new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_,
    new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_,
    new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_,
    new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_,
    new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_,
    new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_,
    new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_,
    new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_,
    new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_,
    new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_,
    new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_,
    new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_,
    new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_,
    new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_,
    new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_,
    new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_,
    new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_,
    new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_,
    new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_,
    new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_,
    new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_,
    new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_,
    new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_,
    new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_,
    new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2576_, new_n2577_,
    new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_,
    new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_,
    new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_,
    new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_,
    new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_,
    new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_,
    new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_,
    new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_,
    new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_,
    new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_,
    new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_,
    new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_,
    new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_,
    new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_,
    new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_,
    new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_,
    new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_,
    new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_,
    new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_,
    new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_,
    new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_,
    new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_,
    new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_,
    new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_,
    new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_,
    new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_,
    new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_,
    new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_,
    new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_,
    new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_,
    new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_,
    new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_,
    new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_,
    new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_,
    new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_,
    new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_,
    new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_,
    new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_,
    new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_,
    new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_,
    new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_,
    new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_,
    new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_,
    new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_,
    new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_,
    new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_,
    new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_,
    new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_,
    new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_,
    new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_,
    new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_,
    new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_,
    new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_,
    new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_,
    new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_,
    new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_,
    new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_,
    new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_,
    new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_,
    new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_,
    new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_,
    new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_,
    new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_,
    new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_,
    new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_,
    new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_,
    new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_,
    new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_,
    new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_,
    new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_,
    new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_,
    new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_,
    new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_,
    new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_,
    new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_,
    new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_,
    new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_,
    new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_,
    new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_,
    new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_,
    new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_,
    new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_,
    new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_,
    new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_,
    new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_,
    new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_,
    new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_,
    new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_,
    new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_,
    new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_,
    new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_,
    new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_,
    new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_,
    new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_,
    new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_,
    new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_,
    new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_,
    new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_,
    new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_,
    new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_,
    new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_,
    new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_,
    new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_,
    new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_,
    new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_,
    new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_,
    new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_,
    new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_,
    new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_,
    new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_,
    new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_,
    new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_,
    new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_,
    new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_,
    new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_,
    new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_,
    new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_,
    new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_,
    new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_,
    new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_,
    new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_,
    new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_,
    new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_,
    new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_,
    new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_,
    new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_,
    new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_,
    new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_,
    new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_,
    new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_,
    new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_,
    new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_,
    new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_,
    new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_,
    new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_,
    new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_,
    new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_,
    new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_,
    new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_,
    new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_,
    new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_,
    new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_,
    new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_,
    new_n4264_, new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_,
    new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_,
    new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_,
    new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_,
    new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_,
    new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_,
    new_n4312_, new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_,
    new_n4318_, new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_,
    new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_,
    new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_,
    new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_,
    new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_,
    new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_,
    new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_,
    new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_,
    new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_,
    new_n4372_, new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_,
    new_n4378_, new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_,
    new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_,
    new_n4390_, new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_,
    new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_,
    new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_,
    new_n4408_, new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_,
    new_n4414_, new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_,
    new_n4420_, new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_,
    new_n4426_, new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_,
    new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_,
    new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_,
    new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_,
    new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_,
    new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_,
    new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_,
    new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_,
    new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_,
    new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_,
    new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4491_,
    new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_, new_n4497_,
    new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_, new_n4503_,
    new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_, new_n4509_,
    new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_, new_n4515_,
    new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_, new_n4521_,
    new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_, new_n4527_,
    new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_, new_n4533_,
    new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_, new_n4539_,
    new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_,
    new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_,
    new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_,
    new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_,
    new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_,
    new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_,
    new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_,
    new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_,
    new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_,
    new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_,
    new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_,
    new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_,
    new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_,
    new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_,
    new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_,
    new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_,
    new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_,
    new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_,
    new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_,
    new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_,
    new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_,
    new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_,
    new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_,
    new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_,
    new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_,
    new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_,
    new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_,
    new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_,
    new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_,
    new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_,
    new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_,
    new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_,
    new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_,
    new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_,
    new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_,
    new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_,
    new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_,
    new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_,
    new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_,
    new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_,
    new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_,
    new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_,
    new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_,
    new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_,
    new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_,
    new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_,
    new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_,
    new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_,
    new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_,
    new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_,
    new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_,
    new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_,
    new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_,
    new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_,
    new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_,
    new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_,
    new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_,
    new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_,
    new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_,
    new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_,
    new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_,
    new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_,
    new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_,
    new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_,
    new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_,
    new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_,
    new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_,
    new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_,
    new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_,
    new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_,
    new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_,
    new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_,
    new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_,
    new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_,
    new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_,
    new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_,
    new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_,
    new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_,
    new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_,
    new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_,
    new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_,
    new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_,
    new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_,
    new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_,
    new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_,
    new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_,
    new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_,
    new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_,
    new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_,
    new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_,
    new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_,
    new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_,
    new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_,
    new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_,
    new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_,
    new_n5290_, new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_,
    new_n5296_, new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_,
    new_n5302_, new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_,
    new_n5308_, new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_,
    new_n5314_, new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_,
    new_n5320_, new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_,
    new_n5326_, new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_,
    new_n5332_, new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_,
    new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_,
    new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_,
    new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_,
    new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_,
    new_n5362_, new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_,
    new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_,
    new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_,
    new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_,
    new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_,
    new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_,
    new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_,
    new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_,
    new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_,
    new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_,
    new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_,
    new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_,
    new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_,
    new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_,
    new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_,
    new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_,
    new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_,
    new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_,
    new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_,
    new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_,
    new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_,
    new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_,
    new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_,
    new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_,
    new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_,
    new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_,
    new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_,
    new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_,
    new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_,
    new_n5536_, new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_,
    new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_,
    new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_,
    new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_,
    new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_,
    new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_,
    new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_,
    new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_,
    new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_,
    new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_,
    new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_,
    new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_,
    new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_,
    new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_,
    new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_,
    new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_,
    new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_,
    new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_,
    new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_,
    new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_,
    new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_,
    new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_,
    new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_,
    new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_,
    new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_,
    new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_,
    new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_,
    new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_,
    new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_,
    new_n5710_, new_n5711_, new_n5712_, new_n5714_, new_n5715_, new_n5716_,
    new_n5717_, new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_,
    new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_,
    new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_,
    new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_,
    new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_,
    new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_,
    new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_,
    new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_,
    new_n5765_, new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_,
    new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_,
    new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_,
    new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_,
    new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_,
    new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_,
    new_n5801_, new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_,
    new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_,
    new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_,
    new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_,
    new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_,
    new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_,
    new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_,
    new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_,
    new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_,
    new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_,
    new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_,
    new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_,
    new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_,
    new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_,
    new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_,
    new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_,
    new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_,
    new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_,
    new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_,
    new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_,
    new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_,
    new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_,
    new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_,
    new_n5939_, new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_,
    new_n5945_, new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_,
    new_n5951_, new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_,
    new_n5957_, new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_,
    new_n5963_, new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_,
    new_n5969_, new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_,
    new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_,
    new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_,
    new_n5987_, new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_,
    new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_,
    new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_,
    new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_,
    new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_,
    new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_,
    new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_,
    new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_,
    new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_,
    new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_,
    new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_,
    new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_,
    new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_,
    new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_,
    new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_,
    new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_,
    new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_,
    new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_,
    new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_,
    new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_,
    new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_,
    new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_,
    new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_,
    new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_,
    new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_,
    new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_,
    new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_,
    new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_,
    new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_,
    new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_,
    new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_,
    new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_,
    new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_,
    new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_,
    new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_,
    new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_,
    new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_,
    new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_,
    new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_,
    new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_,
    new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_,
    new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_,
    new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_,
    new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_,
    new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_,
    new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_,
    new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_,
    new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_,
    new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_,
    new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_,
    new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_,
    new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_,
    new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_,
    new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_,
    new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_,
    new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_,
    new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_,
    new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_,
    new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_,
    new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_,
    new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_,
    new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_,
    new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_,
    new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_,
    new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_,
    new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_,
    new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_,
    new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_,
    new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_,
    new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_,
    new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_,
    new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_,
    new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_,
    new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_,
    new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_,
    new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_,
    new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_,
    new_n6455_, new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_,
    new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_,
    new_n6467_, new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_,
    new_n6473_, new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_,
    new_n6479_, new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_,
    new_n6485_, new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_,
    new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_,
    new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_,
    new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_,
    new_n6509_, new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_,
    new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_,
    new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_,
    new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_,
    new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_,
    new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_,
    new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_,
    new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_,
    new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_,
    new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_,
    new_n6569_, new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_,
    new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_,
    new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_,
    new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_,
    new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_,
    new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_,
    new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_,
    new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_,
    new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_,
    new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_,
    new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_,
    new_n6635_, new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_,
    new_n6641_, new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_,
    new_n6647_, new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_,
    new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_,
    new_n6659_, new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_,
    new_n6665_, new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_,
    new_n6671_, new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_,
    new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_,
    new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_,
    new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_,
    new_n6695_, new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_,
    new_n6701_, new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_,
    new_n6707_, new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_,
    new_n6713_, new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_,
    new_n6719_, new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_,
    new_n6725_, new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_,
    new_n6731_, new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_,
    new_n6737_, new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_,
    new_n6743_, new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_,
    new_n6749_, new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_,
    new_n6755_, new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_,
    new_n6761_, new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_,
    new_n6767_, new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_,
    new_n6773_, new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_,
    new_n6779_, new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_,
    new_n6785_, new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_,
    new_n6791_, new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_,
    new_n6797_, new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_,
    new_n6803_, new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_,
    new_n6809_, new_n6810_, new_n6811_, new_n6812_, new_n6813_, new_n6814_,
    new_n6815_, new_n6816_, new_n6817_, new_n6818_, new_n6819_, new_n6820_,
    new_n6821_, new_n6822_, new_n6823_, new_n6824_, new_n6825_, new_n6826_,
    new_n6827_, new_n6828_, new_n6829_, new_n6830_, new_n6831_, new_n6832_,
    new_n6833_, new_n6834_, new_n6835_, new_n6836_, new_n6837_, new_n6838_,
    new_n6839_, new_n6840_, new_n6841_, new_n6842_, new_n6843_, new_n6844_,
    new_n6845_, new_n6846_, new_n6847_, new_n6848_, new_n6849_, new_n6850_,
    new_n6851_, new_n6852_, new_n6853_, new_n6854_, new_n6855_, new_n6856_,
    new_n6857_, new_n6858_, new_n6859_, new_n6860_, new_n6861_, new_n6862_,
    new_n6863_, new_n6864_, new_n6865_, new_n6866_, new_n6867_, new_n6868_,
    new_n6869_, new_n6870_, new_n6871_, new_n6872_, new_n6873_, new_n6874_,
    new_n6875_, new_n6876_, new_n6877_, new_n6878_, new_n6879_, new_n6880_,
    new_n6881_, new_n6882_, new_n6883_, new_n6884_, new_n6885_, new_n6886_,
    new_n6887_, new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_,
    new_n6893_, new_n6894_, new_n6895_, new_n6896_, new_n6897_, new_n6898_,
    new_n6899_, new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_,
    new_n6905_, new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_,
    new_n6911_, new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_,
    new_n6917_, new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_,
    new_n6923_, new_n6924_, new_n6925_, new_n6926_, new_n6927_, new_n6928_,
    new_n6929_, new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_,
    new_n6935_, new_n6936_, new_n6937_, new_n6938_, new_n6939_, new_n6940_,
    new_n6941_, new_n6942_, new_n6943_, new_n6944_, new_n6945_, new_n6946_,
    new_n6947_, new_n6948_, new_n6949_, new_n6950_, new_n6951_, new_n6952_,
    new_n6953_, new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_,
    new_n6959_, new_n6960_, new_n6961_, new_n6962_, new_n6963_, new_n6964_,
    new_n6965_, new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_,
    new_n6971_, new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_,
    new_n6977_, new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_,
    new_n6983_, new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_,
    new_n6989_, new_n6990_, new_n6991_, new_n6992_, new_n6993_, new_n6994_,
    new_n6995_, new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_,
    new_n7001_, new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_,
    new_n7007_, new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_,
    new_n7013_, new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_,
    new_n7019_, new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_,
    new_n7025_, new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_,
    new_n7031_, new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7038_,
    new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_,
    new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_,
    new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_,
    new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_,
    new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_,
    new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_,
    new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_,
    new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_,
    new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_,
    new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_,
    new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_,
    new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_,
    new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_,
    new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_,
    new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_,
    new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_,
    new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_,
    new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_,
    new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_,
    new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_,
    new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_,
    new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_,
    new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_,
    new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_,
    new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_,
    new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_,
    new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_,
    new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_,
    new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_,
    new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_,
    new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_,
    new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_,
    new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_,
    new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_,
    new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_,
    new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_,
    new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_,
    new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_,
    new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_,
    new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_,
    new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_,
    new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_,
    new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_,
    new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_,
    new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_,
    new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_,
    new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_,
    new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_,
    new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_,
    new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_,
    new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_,
    new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_,
    new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_,
    new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_,
    new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_,
    new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_,
    new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_,
    new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_,
    new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_,
    new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_,
    new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_,
    new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_,
    new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_,
    new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_,
    new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_,
    new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_,
    new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_,
    new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_,
    new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_,
    new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_,
    new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_,
    new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_,
    new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_,
    new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_,
    new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_,
    new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_,
    new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_,
    new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_,
    new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_,
    new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_,
    new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_,
    new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_,
    new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_,
    new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_,
    new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_,
    new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_,
    new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_,
    new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_,
    new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_,
    new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_,
    new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_,
    new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_,
    new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_,
    new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_,
    new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_,
    new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_,
    new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_,
    new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_,
    new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_,
    new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_,
    new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_,
    new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_,
    new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_,
    new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_,
    new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_,
    new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_,
    new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7735_, new_n7736_,
    new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_,
    new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_,
    new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_,
    new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_,
    new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_,
    new_n7767_, new_n7768_, new_n7769_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_,
    new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_,
    new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_,
    new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_,
    new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_,
    new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_,
    new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_,
    new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_,
    new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_,
    new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_,
    new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_,
    new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_,
    new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_,
    new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_,
    new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_,
    new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_,
    new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_,
    new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_,
    new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_,
    new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_,
    new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_,
    new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_,
    new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_,
    new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_,
    new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_,
    new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_,
    new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_,
    new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_,
    new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_,
    new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_,
    new_n8032_, new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_,
    new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_,
    new_n8044_, new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_,
    new_n8050_, new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_,
    new_n8056_, new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_,
    new_n8062_, new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_,
    new_n8068_, new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_,
    new_n8074_, new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_,
    new_n8080_, new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_,
    new_n8086_, new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_,
    new_n8092_, new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_,
    new_n8098_, new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_,
    new_n8104_, new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_,
    new_n8110_, new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_,
    new_n8116_, new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_,
    new_n8122_, new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_,
    new_n8128_, new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_,
    new_n8134_, new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_,
    new_n8140_, new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_,
    new_n8146_, new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_,
    new_n8152_, new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_,
    new_n8158_, new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_,
    new_n8164_, new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_,
    new_n8170_, new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_,
    new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_,
    new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_,
    new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_,
    new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_,
    new_n8200_, new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_,
    new_n8206_, new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_,
    new_n8212_, new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_,
    new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_,
    new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_,
    new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_,
    new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_,
    new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_,
    new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_,
    new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_,
    new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_,
    new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_,
    new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_,
    new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_,
    new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_,
    new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_,
    new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_,
    new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_,
    new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_,
    new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_,
    new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_,
    new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_,
    new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_,
    new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_,
    new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_,
    new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_,
    new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_,
    new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_,
    new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_,
    new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_,
    new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_,
    new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_,
    new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_,
    new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_,
    new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_,
    new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_,
    new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_,
    new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_,
    new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_,
    new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_,
    new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_,
    new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_,
    new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_,
    new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_,
    new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_,
    new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_,
    new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_,
    new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_,
    new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_,
    new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_,
    new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_,
    new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_,
    new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_,
    new_n8525_, new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_,
    new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_,
    new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_,
    new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_,
    new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_,
    new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_,
    new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_,
    new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_,
    new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_,
    new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_,
    new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_,
    new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_,
    new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_,
    new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_,
    new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_,
    new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_,
    new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_,
    new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_,
    new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_,
    new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_,
    new_n8645_, new_n8646_, new_n8648_, new_n8649_, new_n8650_, new_n8651_,
    new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_,
    new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_,
    new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_,
    new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_,
    new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_,
    new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_,
    new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_,
    new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_,
    new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_,
    new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_,
    new_n8737_, new_n8738_, new_n8740_, new_n8741_, new_n8742_, new_n8743_,
    new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_,
    new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_,
    new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_,
    new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_, new_n8767_,
    new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_,
    new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_,
    new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_,
    new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_,
    new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_,
    new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_,
    new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_,
    new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_, new_n8821_,
    new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_,
    new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_,
    new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_,
    new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_,
    new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_,
    new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_,
    new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_,
    new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_,
    new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_,
    new_n9182_, new_n9183_, new_n9184_, new_n9186_, new_n9187_, new_n9188_,
    new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_,
    new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_,
    new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_,
    new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_,
    new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_,
    new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_,
    new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_,
    new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_,
    new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_,
    new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_,
    new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_,
    new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9261_,
    new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_,
    new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_,
    new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_,
    new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_,
    new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_,
    new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_,
    new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_,
    new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_,
    new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_,
    new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_,
    new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_,
    new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_,
    new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_,
    new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_,
    new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_,
    new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_,
    new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_,
    new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_,
    new_n9382_, new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_,
    new_n9388_, new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_,
    new_n9394_, new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_,
    new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_,
    new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_,
    new_n9412_, new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_,
    new_n9418_, new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_,
    new_n9424_, new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_,
    new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_,
    new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_,
    new_n9442_, new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_,
    new_n9448_, new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_,
    new_n9454_, new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_,
    new_n9460_, new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_,
    new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_,
    new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_,
    new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_,
    new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_,
    new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_,
    new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_,
    new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_,
    new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_, new_n9513_,
    new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_,
    new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_, new_n9525_,
    new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_, new_n9531_,
    new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_,
    new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_, new_n9543_,
    new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_, new_n9549_,
    new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_, new_n9555_,
    new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_, new_n9561_,
    new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_, new_n9567_,
    new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_, new_n9573_,
    new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_, new_n9579_,
    new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_, new_n9585_,
    new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_, new_n9591_,
    new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_, new_n9597_,
    new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_, new_n9603_,
    new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_,
    new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_,
    new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_,
    new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_,
    new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_,
    new_n9634_, new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_,
    new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_,
    new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_,
    new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_,
    new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_,
    new_n9664_, new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_,
    new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_,
    new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_,
    new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_,
    new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_,
    new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_,
    new_n9700_, new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_,
    new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_,
    new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_,
    new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_,
    new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_,
    new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_,
    new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_,
    new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_,
    new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_,
    new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_,
    new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_,
    new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_,
    new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_,
    new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_,
    new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_,
    new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_,
    new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_,
    new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_,
    new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_,
    new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_,
    new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_,
    new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_,
    new_n9832_, new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_,
    new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_,
    new_n9844_, new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_,
    new_n9850_, new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_,
    new_n9856_, new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_,
    new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_,
    new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_,
    new_n9874_, new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_,
    new_n9880_, new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_,
    new_n9886_, new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_,
    new_n9892_, new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_,
    new_n9898_, new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_,
    new_n9904_, new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_,
    new_n9910_, new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_,
    new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_,
    new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_,
    new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_,
    new_n9934_, new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_,
    new_n9940_, new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_,
    new_n9946_, new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_,
    new_n9952_, new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_,
    new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_,
    new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_,
    new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_,
    new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_,
    new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_,
    new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_,
    new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10350_, new_n10351_, new_n10352_, new_n10353_, new_n10354_,
    new_n10355_, new_n10356_, new_n10357_, new_n10358_, new_n10359_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10367_, new_n10368_, new_n10369_,
    new_n10370_, new_n10371_, new_n10372_, new_n10373_, new_n10374_,
    new_n10375_, new_n10376_, new_n10377_, new_n10378_, new_n10379_,
    new_n10380_, new_n10381_, new_n10382_, new_n10383_, new_n10384_,
    new_n10385_, new_n10386_, new_n10387_, new_n10388_, new_n10389_,
    new_n10390_, new_n10391_, new_n10392_, new_n10393_, new_n10394_,
    new_n10395_, new_n10396_, new_n10397_, new_n10398_, new_n10399_,
    new_n10400_, new_n10401_, new_n10402_, new_n10403_, new_n10404_,
    new_n10405_, new_n10406_, new_n10407_, new_n10408_, new_n10409_,
    new_n10410_, new_n10411_, new_n10412_, new_n10413_, new_n10414_,
    new_n10415_, new_n10416_, new_n10417_, new_n10418_, new_n10419_,
    new_n10420_, new_n10421_, new_n10422_, new_n10423_, new_n10424_,
    new_n10425_, new_n10426_, new_n10427_, new_n10428_, new_n10429_,
    new_n10430_, new_n10431_, new_n10432_, new_n10433_, new_n10434_,
    new_n10435_, new_n10436_, new_n10437_, new_n10438_, new_n10439_,
    new_n10440_, new_n10441_, new_n10442_, new_n10443_, new_n10444_,
    new_n10445_, new_n10446_, new_n10447_, new_n10448_, new_n10449_,
    new_n10450_, new_n10451_, new_n10452_, new_n10453_, new_n10454_,
    new_n10455_, new_n10456_, new_n10457_, new_n10458_, new_n10459_,
    new_n10460_, new_n10461_, new_n10462_, new_n10463_, new_n10464_,
    new_n10465_, new_n10466_, new_n10467_, new_n10468_, new_n10469_,
    new_n10470_, new_n10471_, new_n10472_, new_n10473_, new_n10474_,
    new_n10475_, new_n10476_, new_n10477_, new_n10478_, new_n10479_,
    new_n10480_, new_n10481_, new_n10482_, new_n10483_, new_n10484_,
    new_n10485_, new_n10486_, new_n10487_, new_n10488_, new_n10489_,
    new_n10490_, new_n10491_, new_n10492_, new_n10493_, new_n10494_,
    new_n10495_, new_n10496_, new_n10497_, new_n10498_, new_n10499_,
    new_n10500_, new_n10501_, new_n10502_, new_n10503_, new_n10504_,
    new_n10505_, new_n10506_, new_n10507_, new_n10508_, new_n10509_,
    new_n10510_, new_n10511_, new_n10512_, new_n10513_, new_n10514_,
    new_n10515_, new_n10516_, new_n10517_, new_n10518_, new_n10519_,
    new_n10520_, new_n10521_, new_n10522_, new_n10523_, new_n10524_,
    new_n10525_, new_n10526_, new_n10527_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10567_, new_n10568_, new_n10569_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10613_, new_n10614_,
    new_n10615_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10627_, new_n10628_, new_n10629_,
    new_n10630_, new_n10631_, new_n10632_, new_n10633_, new_n10634_,
    new_n10635_, new_n10636_, new_n10637_, new_n10638_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10645_, new_n10646_, new_n10647_, new_n10648_, new_n10649_,
    new_n10650_, new_n10651_, new_n10652_, new_n10653_, new_n10654_,
    new_n10655_, new_n10656_, new_n10657_, new_n10658_, new_n10659_,
    new_n10660_, new_n10661_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10728_, new_n10729_,
    new_n10730_, new_n10731_, new_n10732_, new_n10733_, new_n10734_,
    new_n10735_, new_n10736_, new_n10737_, new_n10738_, new_n10739_,
    new_n10740_, new_n10741_, new_n10742_, new_n10743_, new_n10744_,
    new_n10745_, new_n10746_, new_n10747_, new_n10748_, new_n10749_,
    new_n10750_, new_n10751_, new_n10752_, new_n10753_, new_n10754_,
    new_n10755_, new_n10756_, new_n10757_, new_n10758_, new_n10759_,
    new_n10760_, new_n10761_, new_n10762_, new_n10763_, new_n10764_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10817_, new_n10818_, new_n10819_,
    new_n10820_, new_n10821_, new_n10822_, new_n10823_, new_n10824_,
    new_n10825_, new_n10826_, new_n10827_, new_n10828_, new_n10829_,
    new_n10830_, new_n10831_, new_n10832_, new_n10833_, new_n10834_,
    new_n10835_, new_n10836_, new_n10837_, new_n10838_, new_n10839_,
    new_n10840_, new_n10841_, new_n10842_, new_n10843_, new_n10844_,
    new_n10845_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11262_, new_n11263_, new_n11264_, new_n11265_, new_n11266_,
    new_n11267_, new_n11268_, new_n11269_, new_n11270_, new_n11271_,
    new_n11272_, new_n11273_, new_n11274_, new_n11275_, new_n11276_,
    new_n11277_, new_n11278_, new_n11279_, new_n11280_, new_n11281_,
    new_n11282_, new_n11283_, new_n11284_, new_n11285_, new_n11286_,
    new_n11287_, new_n11288_, new_n11289_, new_n11290_, new_n11291_,
    new_n11292_, new_n11293_, new_n11294_, new_n11295_, new_n11296_,
    new_n11297_, new_n11298_, new_n11299_, new_n11300_, new_n11301_,
    new_n11302_, new_n11303_, new_n11304_, new_n11305_, new_n11306_,
    new_n11307_, new_n11308_, new_n11309_, new_n11310_, new_n11311_,
    new_n11312_, new_n11313_, new_n11314_, new_n11315_, new_n11316_,
    new_n11317_, new_n11318_, new_n11319_, new_n11320_, new_n11321_,
    new_n11322_, new_n11323_, new_n11324_, new_n11325_, new_n11326_,
    new_n11327_, new_n11328_, new_n11329_, new_n11330_, new_n11331_,
    new_n11332_, new_n11333_, new_n11334_, new_n11335_, new_n11336_,
    new_n11337_, new_n11338_, new_n11339_, new_n11340_, new_n11341_,
    new_n11342_, new_n11343_, new_n11344_, new_n11345_, new_n11346_,
    new_n11347_, new_n11348_, new_n11349_, new_n11350_, new_n11351_,
    new_n11352_, new_n11353_, new_n11354_, new_n11355_, new_n11356_,
    new_n11357_, new_n11358_, new_n11359_, new_n11360_, new_n11361_,
    new_n11362_, new_n11363_, new_n11364_, new_n11365_, new_n11366_,
    new_n11367_, new_n11368_, new_n11369_, new_n11370_, new_n11371_,
    new_n11372_, new_n11373_, new_n11374_, new_n11375_, new_n11376_,
    new_n11377_, new_n11378_, new_n11379_, new_n11380_, new_n11381_,
    new_n11382_, new_n11383_, new_n11384_, new_n11385_, new_n11386_,
    new_n11387_, new_n11388_, new_n11389_, new_n11390_, new_n11391_,
    new_n11392_, new_n11393_, new_n11394_, new_n11395_, new_n11396_,
    new_n11397_, new_n11398_, new_n11399_, new_n11400_, new_n11401_,
    new_n11402_, new_n11403_, new_n11404_, new_n11405_, new_n11406_,
    new_n11407_, new_n11408_, new_n11409_, new_n11410_, new_n11411_,
    new_n11412_, new_n11413_, new_n11414_, new_n11415_, new_n11416_,
    new_n11417_, new_n11418_, new_n11419_, new_n11420_, new_n11421_,
    new_n11422_, new_n11423_, new_n11424_, new_n11425_, new_n11426_,
    new_n11427_, new_n11428_, new_n11429_, new_n11430_, new_n11431_,
    new_n11432_, new_n11433_, new_n11434_, new_n11435_, new_n11436_,
    new_n11437_, new_n11438_, new_n11439_, new_n11440_, new_n11441_,
    new_n11442_, new_n11443_, new_n11444_, new_n11445_, new_n11446_,
    new_n11447_, new_n11448_, new_n11449_, new_n11450_, new_n11451_,
    new_n11452_, new_n11453_, new_n11454_, new_n11455_, new_n11456_,
    new_n11457_, new_n11458_, new_n11459_, new_n11460_, new_n11461_,
    new_n11462_, new_n11463_, new_n11464_, new_n11465_, new_n11466_,
    new_n11467_, new_n11468_, new_n11469_, new_n11470_, new_n11471_,
    new_n11472_, new_n11473_, new_n11474_, new_n11475_, new_n11476_,
    new_n11477_, new_n11478_, new_n11479_, new_n11480_, new_n11481_,
    new_n11482_, new_n11483_, new_n11484_, new_n11485_, new_n11486_,
    new_n11487_, new_n11488_, new_n11489_, new_n11490_, new_n11491_,
    new_n11492_, new_n11493_, new_n11494_, new_n11495_, new_n11496_,
    new_n11497_, new_n11498_, new_n11499_, new_n11500_, new_n11501_,
    new_n11502_, new_n11503_, new_n11504_, new_n11505_, new_n11506_,
    new_n11507_, new_n11508_, new_n11509_, new_n11510_, new_n11511_,
    new_n11512_, new_n11513_, new_n11514_, new_n11515_, new_n11516_,
    new_n11517_, new_n11518_, new_n11519_, new_n11520_, new_n11521_,
    new_n11522_, new_n11523_, new_n11524_, new_n11525_, new_n11526_,
    new_n11527_, new_n11528_, new_n11529_, new_n11530_, new_n11531_,
    new_n11532_, new_n11533_, new_n11534_, new_n11535_, new_n11536_,
    new_n11537_, new_n11538_, new_n11539_, new_n11540_, new_n11541_,
    new_n11542_, new_n11543_, new_n11544_, new_n11545_, new_n11546_,
    new_n11547_, new_n11548_, new_n11549_, new_n11550_, new_n11551_,
    new_n11552_, new_n11553_, new_n11554_, new_n11555_, new_n11556_,
    new_n11557_, new_n11558_, new_n11559_, new_n11560_, new_n11561_,
    new_n11562_, new_n11563_, new_n11564_, new_n11565_, new_n11566_,
    new_n11567_, new_n11568_, new_n11569_, new_n11570_, new_n11571_,
    new_n11572_, new_n11573_, new_n11574_, new_n11575_, new_n11576_,
    new_n11577_, new_n11578_, new_n11579_, new_n11580_, new_n11581_,
    new_n11582_, new_n11583_, new_n11584_, new_n11585_, new_n11586_,
    new_n11587_, new_n11588_, new_n11589_, new_n11590_, new_n11591_,
    new_n11592_, new_n11593_, new_n11594_, new_n11595_, new_n11596_,
    new_n11597_, new_n11598_, new_n11599_, new_n11600_, new_n11601_,
    new_n11602_, new_n11603_, new_n11604_, new_n11605_, new_n11606_,
    new_n11607_, new_n11608_, new_n11609_, new_n11610_, new_n11611_,
    new_n11612_, new_n11613_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11618_, new_n11619_, new_n11620_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11645_, new_n11646_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11652_, new_n11653_, new_n11654_, new_n11655_, new_n11656_,
    new_n11657_, new_n11658_, new_n11659_, new_n11660_, new_n11661_,
    new_n11662_, new_n11663_, new_n11664_, new_n11665_, new_n11666_,
    new_n11667_, new_n11668_, new_n11669_, new_n11670_, new_n11671_,
    new_n11672_, new_n11673_, new_n11674_, new_n11675_, new_n11676_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11682_, new_n11683_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11712_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11721_,
    new_n11722_, new_n11723_, new_n11724_, new_n11725_, new_n11726_,
    new_n11727_, new_n11728_, new_n11729_, new_n11730_, new_n11731_,
    new_n11732_, new_n11733_, new_n11734_, new_n11735_, new_n11736_,
    new_n11737_, new_n11738_, new_n11739_, new_n11740_, new_n11741_,
    new_n11742_, new_n11743_, new_n11744_, new_n11745_, new_n11746_,
    new_n11747_, new_n11748_, new_n11749_, new_n11750_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11761_,
    new_n11762_, new_n11763_, new_n11764_, new_n11765_, new_n11766_,
    new_n11767_, new_n11768_, new_n11769_, new_n11770_, new_n11771_,
    new_n11772_, new_n11773_, new_n11774_, new_n11775_, new_n11776_,
    new_n11777_, new_n11778_, new_n11779_, new_n11780_, new_n11781_,
    new_n11782_, new_n11783_, new_n11784_, new_n11785_, new_n11786_,
    new_n11787_, new_n11788_, new_n11789_, new_n11790_, new_n11791_,
    new_n11792_, new_n11793_, new_n11794_, new_n11795_, new_n11796_,
    new_n11797_, new_n11798_, new_n11799_, new_n11800_, new_n11801_,
    new_n11802_, new_n11803_, new_n11804_, new_n11805_, new_n11806_,
    new_n11807_, new_n11808_, new_n11809_, new_n11810_, new_n11811_,
    new_n11812_, new_n11813_, new_n11814_, new_n11815_, new_n11816_,
    new_n11817_, new_n11818_, new_n11819_, new_n11820_, new_n11821_,
    new_n11822_, new_n11823_, new_n11824_, new_n11825_, new_n11826_,
    new_n11827_, new_n11828_, new_n11829_, new_n11830_, new_n11831_,
    new_n11832_, new_n11833_, new_n11834_, new_n11835_, new_n11836_,
    new_n11837_, new_n11838_, new_n11839_, new_n11840_, new_n11841_,
    new_n11842_, new_n11843_, new_n11844_, new_n11845_, new_n11846_,
    new_n11847_, new_n11848_, new_n11849_, new_n11850_, new_n11851_,
    new_n11852_, new_n11853_, new_n11854_, new_n11855_, new_n11856_,
    new_n11857_, new_n11858_, new_n11859_, new_n11860_, new_n11861_,
    new_n11862_, new_n11863_, new_n11864_, new_n11865_, new_n11866_,
    new_n11867_, new_n11868_, new_n11869_, new_n11870_, new_n11871_,
    new_n11872_, new_n11873_, new_n11874_, new_n11875_, new_n11876_,
    new_n11877_, new_n11878_, new_n11879_, new_n11880_, new_n11881_,
    new_n11882_, new_n11883_, new_n11884_, new_n11885_, new_n11886_,
    new_n11887_, new_n11888_, new_n11889_, new_n11890_, new_n11891_,
    new_n11892_, new_n11893_, new_n11894_, new_n11895_, new_n11896_,
    new_n11897_, new_n11898_, new_n11899_, new_n11900_, new_n11901_,
    new_n11902_, new_n11903_, new_n11904_, new_n11905_, new_n11906_,
    new_n11907_, new_n11908_, new_n11909_, new_n11910_, new_n11911_,
    new_n11912_, new_n11913_, new_n11914_, new_n11915_, new_n11916_,
    new_n11917_, new_n11918_, new_n11919_, new_n11920_, new_n11921_,
    new_n11922_, new_n11923_, new_n11924_, new_n11925_, new_n11926_,
    new_n11927_, new_n11928_, new_n11929_, new_n11930_, new_n11931_,
    new_n11932_, new_n11933_, new_n11934_, new_n11935_, new_n11936_,
    new_n11937_, new_n11938_, new_n11939_, new_n11940_, new_n11941_,
    new_n11942_, new_n11943_, new_n11944_, new_n11945_, new_n11946_,
    new_n11947_, new_n11948_, new_n11949_, new_n11950_, new_n11951_,
    new_n11952_, new_n11953_, new_n11954_, new_n11955_, new_n11956_,
    new_n11957_, new_n11958_, new_n11959_, new_n11960_, new_n11961_,
    new_n11962_, new_n11963_, new_n11964_, new_n11965_, new_n11966_,
    new_n11967_, new_n11968_, new_n11969_, new_n11970_, new_n11971_,
    new_n11972_, new_n11973_, new_n11974_, new_n11975_, new_n11976_,
    new_n11977_, new_n11978_, new_n11979_, new_n11980_, new_n11981_,
    new_n11982_, new_n11983_, new_n11984_, new_n11985_, new_n11986_,
    new_n11987_, new_n11988_, new_n11989_, new_n11990_, new_n11991_,
    new_n11992_, new_n11993_, new_n11994_, new_n11995_, new_n11996_,
    new_n11997_, new_n11998_, new_n11999_, new_n12000_, new_n12001_,
    new_n12002_, new_n12003_, new_n12004_, new_n12005_, new_n12006_,
    new_n12007_, new_n12008_, new_n12009_, new_n12010_, new_n12011_,
    new_n12012_, new_n12013_, new_n12014_, new_n12015_, new_n12016_,
    new_n12017_, new_n12018_, new_n12019_, new_n12020_, new_n12021_,
    new_n12022_, new_n12023_, new_n12024_, new_n12025_, new_n12026_,
    new_n12027_, new_n12028_, new_n12029_, new_n12030_, new_n12031_,
    new_n12032_, new_n12033_, new_n12034_, new_n12035_, new_n12036_,
    new_n12037_, new_n12038_, new_n12039_, new_n12040_, new_n12041_,
    new_n12042_, new_n12043_, new_n12044_, new_n12045_, new_n12046_,
    new_n12047_, new_n12048_, new_n12049_, new_n12050_, new_n12051_,
    new_n12052_, new_n12053_, new_n12054_, new_n12055_, new_n12056_,
    new_n12057_, new_n12058_, new_n12059_, new_n12060_, new_n12061_,
    new_n12062_, new_n12063_, new_n12064_, new_n12065_, new_n12066_,
    new_n12067_, new_n12068_, new_n12069_, new_n12070_, new_n12071_,
    new_n12072_, new_n12073_, new_n12074_, new_n12075_, new_n12076_,
    new_n12077_, new_n12078_, new_n12079_, new_n12080_, new_n12081_,
    new_n12082_, new_n12083_, new_n12084_, new_n12085_, new_n12086_,
    new_n12087_, new_n12088_, new_n12089_, new_n12090_, new_n12091_,
    new_n12092_, new_n12093_, new_n12094_, new_n12095_, new_n12096_,
    new_n12097_, new_n12098_, new_n12099_, new_n12100_, new_n12101_,
    new_n12102_, new_n12104_, new_n12105_, new_n12106_, new_n12108_,
    new_n12109_, new_n12110_, new_n12111_, new_n12112_, new_n12113_,
    new_n12114_, new_n12115_, new_n12116_, new_n12117_, new_n12118_,
    new_n12119_, new_n12120_, new_n12121_, new_n12122_, new_n12123_,
    new_n12124_, new_n12125_, new_n12126_, new_n12127_, new_n12128_,
    new_n12129_, new_n12130_, new_n12131_, new_n12132_, new_n12133_,
    new_n12134_, new_n12135_, new_n12136_, new_n12137_, new_n12138_,
    new_n12139_, new_n12140_, new_n12141_, new_n12142_, new_n12143_,
    new_n12144_, new_n12145_, new_n12146_, new_n12147_, new_n12148_,
    new_n12149_, new_n12150_, new_n12151_, new_n12152_, new_n12153_,
    new_n12154_, new_n12155_, new_n12156_, new_n12157_, new_n12158_,
    new_n12159_, new_n12160_, new_n12161_, new_n12162_, new_n12163_,
    new_n12164_, new_n12165_, new_n12166_, new_n12167_, new_n12168_,
    new_n12169_, new_n12170_, new_n12171_, new_n12172_, new_n12173_,
    new_n12174_, new_n12175_, new_n12176_, new_n12177_, new_n12178_,
    new_n12179_, new_n12180_, new_n12181_, new_n12182_, new_n12183_,
    new_n12184_, new_n12185_, new_n12186_, new_n12187_, new_n12188_,
    new_n12189_, new_n12190_, new_n12191_, new_n12192_, new_n12193_,
    new_n12194_, new_n12195_, new_n12196_, new_n12197_, new_n12198_,
    new_n12199_, new_n12200_, new_n12201_, new_n12202_, new_n12203_,
    new_n12204_, new_n12205_, new_n12206_, new_n12207_, new_n12208_,
    new_n12209_, new_n12210_, new_n12211_, new_n12212_, new_n12213_,
    new_n12214_, new_n12215_, new_n12216_, new_n12217_, new_n12218_,
    new_n12219_, new_n12220_, new_n12221_, new_n12222_, new_n12223_,
    new_n12224_, new_n12225_, new_n12226_, new_n12227_, new_n12228_,
    new_n12229_, new_n12230_, new_n12231_, new_n12232_, new_n12233_,
    new_n12234_, new_n12235_, new_n12236_, new_n12237_, new_n12238_,
    new_n12239_, new_n12240_, new_n12241_, new_n12242_, new_n12243_,
    new_n12244_, new_n12245_, new_n12246_, new_n12247_, new_n12248_,
    new_n12249_, new_n12250_, new_n12251_, new_n12252_, new_n12253_,
    new_n12254_, new_n12255_, new_n12256_, new_n12257_, new_n12258_,
    new_n12259_, new_n12260_, new_n12261_, new_n12262_, new_n12263_,
    new_n12264_, new_n12265_, new_n12266_, new_n12267_, new_n12268_,
    new_n12269_, new_n12270_, new_n12271_, new_n12272_, new_n12273_,
    new_n12274_, new_n12275_, new_n12276_, new_n12277_, new_n12278_,
    new_n12279_, new_n12280_, new_n12281_, new_n12282_, new_n12283_,
    new_n12284_, new_n12285_, new_n12286_, new_n12287_, new_n12288_,
    new_n12289_, new_n12290_, new_n12291_, new_n12292_, new_n12293_,
    new_n12294_, new_n12295_, new_n12296_, new_n12297_, new_n12298_,
    new_n12299_, new_n12300_, new_n12301_, new_n12302_, new_n12303_,
    new_n12304_, new_n12305_, new_n12306_, new_n12307_, new_n12308_,
    new_n12309_, new_n12310_, new_n12311_, new_n12312_, new_n12313_,
    new_n12314_, new_n12315_, new_n12316_, new_n12317_, new_n12318_,
    new_n12319_, new_n12320_, new_n12321_, new_n12322_, new_n12323_,
    new_n12324_, new_n12325_, new_n12326_, new_n12327_, new_n12328_,
    new_n12329_, new_n12330_, new_n12331_, new_n12332_, new_n12333_,
    new_n12334_, new_n12335_, new_n12336_, new_n12337_, new_n12338_,
    new_n12339_, new_n12340_, new_n12341_, new_n12342_, new_n12343_,
    new_n12344_, new_n12345_, new_n12346_, new_n12347_, new_n12348_,
    new_n12349_, new_n12350_, new_n12351_, new_n12352_, new_n12353_,
    new_n12354_, new_n12355_, new_n12356_, new_n12357_, new_n12358_,
    new_n12359_, new_n12360_, new_n12361_, new_n12362_, new_n12363_,
    new_n12364_, new_n12365_, new_n12366_, new_n12367_, new_n12368_,
    new_n12369_, new_n12370_, new_n12371_, new_n12372_, new_n12373_,
    new_n12374_, new_n12375_, new_n12376_, new_n12377_, new_n12378_,
    new_n12379_, new_n12380_, new_n12381_, new_n12382_, new_n12383_,
    new_n12384_, new_n12385_, new_n12386_, new_n12387_, new_n12388_,
    new_n12389_, new_n12390_, new_n12391_, new_n12392_, new_n12393_,
    new_n12394_, new_n12395_, new_n12396_, new_n12397_, new_n12398_,
    new_n12399_, new_n12400_, new_n12401_, new_n12402_, new_n12403_,
    new_n12404_, new_n12405_, new_n12406_, new_n12407_, new_n12408_,
    new_n12409_, new_n12410_, new_n12411_, new_n12412_, new_n12413_,
    new_n12414_, new_n12415_, new_n12416_, new_n12417_, new_n12418_,
    new_n12419_, new_n12420_, new_n12421_, new_n12422_, new_n12423_,
    new_n12424_, new_n12425_, new_n12426_, new_n12427_, new_n12428_,
    new_n12429_, new_n12430_, new_n12431_, new_n12432_, new_n12433_,
    new_n12434_, new_n12435_, new_n12436_, new_n12437_, new_n12438_,
    new_n12439_, new_n12440_, new_n12441_, new_n12442_, new_n12443_,
    new_n12444_, new_n12445_, new_n12446_, new_n12447_, new_n12448_,
    new_n12449_, new_n12450_, new_n12451_, new_n12452_, new_n12453_,
    new_n12454_, new_n12455_, new_n12456_, new_n12457_, new_n12458_,
    new_n12459_, new_n12460_, new_n12461_, new_n12462_, new_n12463_,
    new_n12464_, new_n12465_, new_n12466_, new_n12467_, new_n12468_,
    new_n12469_, new_n12470_, new_n12471_, new_n12472_, new_n12473_,
    new_n12474_, new_n12475_, new_n12476_, new_n12477_, new_n12478_,
    new_n12479_, new_n12480_, new_n12481_, new_n12482_, new_n12483_,
    new_n12484_, new_n12485_, new_n12486_, new_n12487_, new_n12488_,
    new_n12489_, new_n12490_, new_n12491_, new_n12492_, new_n12493_,
    new_n12494_, new_n12495_, new_n12496_, new_n12497_, new_n12498_,
    new_n12499_, new_n12500_, new_n12501_, new_n12502_, new_n12503_,
    new_n12504_, new_n12505_, new_n12506_, new_n12507_, new_n12508_,
    new_n12509_, new_n12510_, new_n12511_, new_n12512_, new_n12513_,
    new_n12514_, new_n12515_, new_n12516_, new_n12517_, new_n12518_,
    new_n12519_, new_n12520_, new_n12521_, new_n12522_, new_n12523_,
    new_n12524_, new_n12525_, new_n12526_, new_n12527_, new_n12528_,
    new_n12529_, new_n12530_, new_n12531_, new_n12532_, new_n12533_,
    new_n12534_, new_n12535_, new_n12536_, new_n12537_, new_n12538_,
    new_n12539_, new_n12540_, new_n12541_, new_n12542_, new_n12543_,
    new_n12544_, new_n12545_, new_n12546_, new_n12547_, new_n12548_,
    new_n12549_, new_n12550_, new_n12551_, new_n12552_, new_n12553_,
    new_n12554_, new_n12555_, new_n12556_, new_n12557_, new_n12558_,
    new_n12559_, new_n12560_, new_n12561_, new_n12562_, new_n12563_,
    new_n12564_, new_n12565_, new_n12566_, new_n12567_, new_n12568_,
    new_n12569_, new_n12570_, new_n12571_, new_n12572_, new_n12573_,
    new_n12574_, new_n12575_, new_n12576_, new_n12577_, new_n12578_,
    new_n12579_, new_n12580_, new_n12581_, new_n12582_, new_n12583_,
    new_n12584_, new_n12585_, new_n12586_, new_n12587_, new_n12588_,
    new_n12589_, new_n12590_, new_n12591_, new_n12592_, new_n12593_,
    new_n12594_, new_n12595_, new_n12596_, new_n12597_, new_n12598_,
    new_n12599_, new_n12600_, new_n12601_, new_n12602_, new_n12603_,
    new_n12604_, new_n12605_, new_n12606_, new_n12607_, new_n12608_,
    new_n12609_, new_n12611_, new_n12612_, new_n12613_, new_n12614_,
    new_n12615_, new_n12616_, new_n12617_, new_n12618_, new_n12619_,
    new_n12620_, new_n12621_, new_n12622_, new_n12623_, new_n12624_,
    new_n12625_, new_n12626_, new_n12627_, new_n12628_, new_n12629_,
    new_n12630_, new_n12631_, new_n12632_, new_n12633_, new_n12634_,
    new_n12635_, new_n12636_, new_n12637_, new_n12638_, new_n12639_,
    new_n12640_, new_n12641_, new_n12642_, new_n12643_, new_n12644_,
    new_n12645_, new_n12646_, new_n12647_, new_n12648_, new_n12649_,
    new_n12650_, new_n12651_, new_n12652_, new_n12653_, new_n12654_,
    new_n12655_, new_n12656_, new_n12657_, new_n12658_, new_n12659_,
    new_n12660_, new_n12661_, new_n12662_, new_n12663_, new_n12664_,
    new_n12665_, new_n12666_, new_n12667_, new_n12668_, new_n12669_,
    new_n12670_, new_n12671_, new_n12672_, new_n12673_, new_n12674_,
    new_n12675_, new_n12676_, new_n12677_, new_n12678_, new_n12679_,
    new_n12680_, new_n12681_, new_n12682_, new_n12683_, new_n12684_,
    new_n12685_, new_n12686_, new_n12687_, new_n12688_, new_n12689_,
    new_n12690_, new_n12691_, new_n12692_, new_n12693_, new_n12694_,
    new_n12695_, new_n12696_, new_n12697_, new_n12698_, new_n12699_,
    new_n12700_, new_n12701_, new_n12702_, new_n12703_, new_n12704_,
    new_n12705_, new_n12706_, new_n12707_, new_n12708_, new_n12709_,
    new_n12710_, new_n12711_, new_n12712_, new_n12713_, new_n12714_,
    new_n12715_, new_n12716_, new_n12717_, new_n12718_, new_n12719_,
    new_n12720_, new_n12721_, new_n12722_, new_n12723_, new_n12724_,
    new_n12725_, new_n12726_, new_n12727_, new_n12728_, new_n12729_,
    new_n12730_, new_n12731_, new_n12732_, new_n12733_, new_n12734_,
    new_n12735_, new_n12736_, new_n12737_, new_n12738_, new_n12739_,
    new_n12740_, new_n12741_, new_n12742_, new_n12743_, new_n12744_,
    new_n12745_, new_n12746_, new_n12747_, new_n12748_, new_n12749_,
    new_n12750_, new_n12751_, new_n12752_, new_n12753_, new_n12754_,
    new_n12755_, new_n12756_, new_n12757_, new_n12758_, new_n12759_,
    new_n12760_, new_n12761_, new_n12762_, new_n12763_, new_n12764_,
    new_n12765_, new_n12766_, new_n12767_, new_n12768_, new_n12769_,
    new_n12770_, new_n12771_, new_n12772_, new_n12773_, new_n12774_,
    new_n12775_, new_n12776_, new_n12777_, new_n12778_, new_n12779_,
    new_n12780_, new_n12781_, new_n12782_, new_n12783_, new_n12784_,
    new_n12785_, new_n12786_, new_n12787_, new_n12788_, new_n12789_,
    new_n12790_, new_n12791_, new_n12792_, new_n12793_, new_n12794_,
    new_n12795_, new_n12796_, new_n12797_, new_n12798_, new_n12799_,
    new_n12800_, new_n12801_, new_n12802_, new_n12803_, new_n12804_,
    new_n12805_, new_n12806_, new_n12807_, new_n12808_, new_n12809_,
    new_n12810_, new_n12811_, new_n12812_, new_n12813_, new_n12814_,
    new_n12815_, new_n12816_, new_n12817_, new_n12818_, new_n12819_,
    new_n12820_, new_n12821_, new_n12822_, new_n12823_, new_n12824_,
    new_n12825_, new_n12826_, new_n12827_, new_n12828_, new_n12829_,
    new_n12830_, new_n12831_, new_n12832_, new_n12833_, new_n12834_,
    new_n12835_, new_n12836_, new_n12837_, new_n12838_, new_n12839_,
    new_n12840_, new_n12841_, new_n12842_, new_n12843_, new_n12844_,
    new_n12845_, new_n12846_, new_n12847_, new_n12848_, new_n12849_,
    new_n12850_, new_n12851_, new_n12852_, new_n12853_, new_n12854_,
    new_n12855_, new_n12856_, new_n12857_, new_n12858_, new_n12859_,
    new_n12860_, new_n12861_, new_n12862_, new_n12863_, new_n12864_,
    new_n12865_, new_n12866_, new_n12867_, new_n12868_, new_n12869_,
    new_n12870_, new_n12871_, new_n12872_, new_n12873_, new_n12874_,
    new_n12875_, new_n12876_, new_n12877_, new_n12878_, new_n12879_,
    new_n12880_, new_n12881_, new_n12882_, new_n12883_, new_n12884_,
    new_n12885_, new_n12886_, new_n12887_, new_n12888_, new_n12889_,
    new_n12890_, new_n12891_, new_n12892_, new_n12893_, new_n12894_,
    new_n12895_, new_n12896_, new_n12897_, new_n12898_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13006_, new_n13007_, new_n13008_, new_n13009_,
    new_n13010_, new_n13011_, new_n13012_, new_n13013_, new_n13014_,
    new_n13015_, new_n13016_, new_n13017_, new_n13018_, new_n13019_,
    new_n13020_, new_n13021_, new_n13022_, new_n13023_, new_n13024_,
    new_n13025_, new_n13026_, new_n13027_, new_n13028_, new_n13029_,
    new_n13030_, new_n13031_, new_n13032_, new_n13033_, new_n13034_,
    new_n13035_, new_n13036_, new_n13037_, new_n13038_, new_n13039_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13046_, new_n13047_, new_n13048_, new_n13049_,
    new_n13050_, new_n13051_, new_n13052_, new_n13053_, new_n13054_,
    new_n13055_, new_n13056_, new_n13057_, new_n13058_, new_n13059_,
    new_n13060_, new_n13061_, new_n13062_, new_n13063_, new_n13064_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13069_,
    new_n13070_, new_n13071_, new_n13072_, new_n13073_, new_n13074_,
    new_n13075_, new_n13076_, new_n13077_, new_n13078_, new_n13079_,
    new_n13080_, new_n13081_, new_n13082_, new_n13083_, new_n13084_,
    new_n13085_, new_n13086_, new_n13087_, new_n13088_, new_n13089_,
    new_n13090_, new_n13091_, new_n13092_, new_n13093_, new_n13094_,
    new_n13095_, new_n13096_, new_n13097_, new_n13098_, new_n13099_,
    new_n13100_, new_n13101_, new_n13102_, new_n13103_, new_n13104_,
    new_n13105_, new_n13106_, new_n13107_, new_n13108_, new_n13109_,
    new_n13110_, new_n13111_, new_n13112_, new_n13113_, new_n13114_,
    new_n13115_, new_n13116_, new_n13117_, new_n13118_, new_n13119_,
    new_n13120_, new_n13121_, new_n13122_, new_n13123_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13222_, new_n13223_, new_n13224_, new_n13225_, new_n13226_,
    new_n13227_, new_n13228_, new_n13229_, new_n13230_, new_n13231_,
    new_n13232_, new_n13233_, new_n13234_, new_n13235_, new_n13236_,
    new_n13237_, new_n13238_, new_n13239_, new_n13240_, new_n13241_,
    new_n13242_, new_n13243_, new_n13244_, new_n13245_, new_n13246_,
    new_n13247_, new_n13248_, new_n13249_, new_n13250_, new_n13251_,
    new_n13252_, new_n13253_, new_n13254_, new_n13255_, new_n13256_,
    new_n13257_, new_n13258_, new_n13259_, new_n13260_, new_n13261_,
    new_n13262_, new_n13263_, new_n13264_, new_n13265_, new_n13266_,
    new_n13267_, new_n13268_, new_n13269_, new_n13270_, new_n13271_,
    new_n13272_, new_n13273_, new_n13274_, new_n13275_, new_n13276_,
    new_n13277_, new_n13278_, new_n13279_, new_n13280_, new_n13281_,
    new_n13282_, new_n13283_, new_n13284_, new_n13285_, new_n13286_,
    new_n13287_, new_n13288_, new_n13289_, new_n13290_, new_n13291_,
    new_n13292_, new_n13293_, new_n13294_, new_n13295_, new_n13296_,
    new_n13297_, new_n13298_, new_n13299_, new_n13300_, new_n13301_,
    new_n13302_, new_n13303_, new_n13304_, new_n13306_, new_n13307_,
    new_n13308_, new_n13309_, new_n13310_, new_n13311_, new_n13312_,
    new_n13313_, new_n13314_, new_n13315_, new_n13316_, new_n13317_,
    new_n13318_, new_n13319_, new_n13320_, new_n13321_, new_n13322_,
    new_n13323_, new_n13324_, new_n13325_, new_n13326_, new_n13327_,
    new_n13328_, new_n13329_, new_n13330_, new_n13331_, new_n13332_,
    new_n13333_, new_n13334_, new_n13335_, new_n13336_, new_n13337_,
    new_n13338_, new_n13339_, new_n13340_, new_n13341_, new_n13342_,
    new_n13343_, new_n13344_, new_n13345_, new_n13346_, new_n13347_,
    new_n13348_, new_n13349_, new_n13350_, new_n13351_, new_n13352_,
    new_n13353_, new_n13354_, new_n13355_, new_n13356_, new_n13357_,
    new_n13358_, new_n13359_, new_n13360_, new_n13361_, new_n13362_,
    new_n13363_, new_n13364_, new_n13365_, new_n13366_, new_n13367_,
    new_n13368_, new_n13369_, new_n13370_, new_n13371_, new_n13372_,
    new_n13373_, new_n13374_, new_n13375_, new_n13376_, new_n13377_,
    new_n13378_, new_n13379_, new_n13380_, new_n13381_, new_n13382_,
    new_n13383_, new_n13384_, new_n13385_, new_n13386_, new_n13387_,
    new_n13388_, new_n13389_, new_n13390_, new_n13391_, new_n13392_,
    new_n13393_, new_n13394_, new_n13395_, new_n13396_, new_n13397_,
    new_n13398_, new_n13399_, new_n13400_, new_n13401_, new_n13402_,
    new_n13403_, new_n13405_, new_n13406_, new_n13407_, new_n13408_,
    new_n13410_, new_n13411_, new_n13413_, new_n13414_, new_n13416_,
    new_n13417_, new_n13418_, new_n13419_, new_n13420_, new_n13421_,
    new_n13422_, new_n13423_, new_n13424_, new_n13425_, new_n13426_,
    new_n13427_, new_n13428_, new_n13429_, new_n13430_, new_n13431_,
    new_n13432_, new_n13433_, new_n13434_, new_n13435_, new_n13436_,
    new_n13437_, new_n13438_, new_n13439_, new_n13440_, new_n13441_,
    new_n13442_, new_n13443_, new_n13444_, new_n13445_, new_n13446_,
    new_n13447_, new_n13448_, new_n13449_, new_n13450_, new_n13451_,
    new_n13452_, new_n13453_, new_n13454_, new_n13455_, new_n13456_,
    new_n13457_, new_n13458_, new_n13459_, new_n13460_, new_n13461_,
    new_n13462_, new_n13463_, new_n13464_, new_n13465_, new_n13466_,
    new_n13467_, new_n13468_, new_n13469_, new_n13470_, new_n13471_,
    new_n13472_, new_n13473_, new_n13474_, new_n13475_, new_n13476_,
    new_n13477_, new_n13478_, new_n13479_, new_n13480_, new_n13481_,
    new_n13482_, new_n13483_, new_n13484_, new_n13485_, new_n13486_,
    new_n13487_, new_n13488_, new_n13489_, new_n13490_, new_n13491_,
    new_n13492_, new_n13493_, new_n13494_, new_n13495_, new_n13496_,
    new_n13497_, new_n13498_, new_n13499_, new_n13500_, new_n13501_,
    new_n13502_, new_n13503_, new_n13504_, new_n13505_, new_n13506_,
    new_n13507_, new_n13508_, new_n13509_, new_n13510_, new_n13511_,
    new_n13512_, new_n13513_, new_n13514_, new_n13515_, new_n13516_,
    new_n13517_, new_n13518_, new_n13519_, new_n13520_, new_n13521_,
    new_n13522_, new_n13523_, new_n13524_, new_n13525_, new_n13526_,
    new_n13527_, new_n13528_, new_n13529_, new_n13530_, new_n13531_,
    new_n13532_, new_n13533_, new_n13534_, new_n13535_, new_n13536_,
    new_n13537_, new_n13538_, new_n13539_, new_n13540_, new_n13541_,
    new_n13542_, new_n13543_, new_n13544_, new_n13545_, new_n13546_,
    new_n13547_, new_n13548_, new_n13549_, new_n13550_, new_n13551_,
    new_n13552_, new_n13553_, new_n13554_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13596_,
    new_n13597_, new_n13598_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13605_, new_n13606_,
    new_n13607_, new_n13608_, new_n13609_, new_n13610_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13637_, new_n13638_, new_n13639_, new_n13640_, new_n13641_,
    new_n13642_, new_n13643_, new_n13644_, new_n13645_, new_n13646_,
    new_n13647_, new_n13648_, new_n13649_, new_n13650_, new_n13651_,
    new_n13652_, new_n13653_, new_n13654_, new_n13655_, new_n13656_,
    new_n13657_, new_n13658_, new_n13659_, new_n13660_, new_n13661_,
    new_n13662_, new_n13663_, new_n13664_, new_n13665_, new_n13666_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13744_, new_n13745_, new_n13746_,
    new_n13747_, new_n13748_, new_n13749_, new_n13750_, new_n13751_,
    new_n13752_, new_n13753_, new_n13754_, new_n13755_, new_n13756_,
    new_n13757_, new_n13758_, new_n13759_, new_n13760_, new_n13761_,
    new_n13762_, new_n13763_, new_n13764_, new_n13765_, new_n13766_,
    new_n13767_, new_n13768_, new_n13769_, new_n13770_, new_n13771_,
    new_n13772_, new_n13773_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13785_, new_n13786_,
    new_n13787_, new_n13788_, new_n13789_, new_n13790_, new_n13791_,
    new_n13792_, new_n13793_, new_n13794_, new_n13795_, new_n13796_,
    new_n13797_, new_n13798_, new_n13799_, new_n13800_, new_n13801_,
    new_n13802_, new_n13803_, new_n13804_, new_n13805_, new_n13806_,
    new_n13807_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13814_, new_n13815_, new_n13816_,
    new_n13817_, new_n13818_, new_n13819_, new_n13820_, new_n13821_,
    new_n13822_, new_n13823_, new_n13824_, new_n13825_, new_n13826_,
    new_n13827_, new_n13828_, new_n13829_, new_n13830_, new_n13831_,
    new_n13832_, new_n13833_, new_n13834_, new_n13835_, new_n13836_,
    new_n13837_, new_n13838_, new_n13839_, new_n13840_, new_n13841_,
    new_n13842_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13847_, new_n13848_, new_n13849_, new_n13850_, new_n13851_,
    new_n13852_, new_n13853_, new_n13854_, new_n13855_, new_n13856_,
    new_n13857_, new_n13858_, new_n13859_, new_n13860_, new_n13861_,
    new_n13862_, new_n13863_, new_n13864_, new_n13865_, new_n13866_,
    new_n13867_, new_n13868_, new_n13869_, new_n13870_, new_n13871_,
    new_n13872_, new_n13873_, new_n13874_, new_n13875_, new_n13876_,
    new_n13877_, new_n13878_, new_n13879_, new_n13880_, new_n13881_,
    new_n13882_, new_n13883_, new_n13884_, new_n13885_, new_n13886_,
    new_n13887_, new_n13888_, new_n13889_, new_n13890_, new_n13891_,
    new_n13892_, new_n13893_, new_n13894_, new_n13895_, new_n13896_,
    new_n13897_, new_n13898_, new_n13899_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13951_,
    new_n13952_, new_n13953_, new_n13954_, new_n13955_, new_n13956_,
    new_n13957_, new_n13958_, new_n13959_, new_n13960_, new_n13961_,
    new_n13962_, new_n13963_, new_n13964_, new_n13965_, new_n13966_,
    new_n13967_, new_n13968_, new_n13969_, new_n13970_, new_n13971_,
    new_n13972_, new_n13973_, new_n13974_, new_n13975_, new_n13976_,
    new_n13977_, new_n13978_, new_n13979_, new_n13980_, new_n13981_,
    new_n13982_, new_n13983_, new_n13984_, new_n13985_, new_n13986_,
    new_n13987_, new_n13988_, new_n13989_, new_n13990_, new_n13991_,
    new_n13992_, new_n13993_, new_n13994_, new_n13995_, new_n13996_,
    new_n13997_, new_n13998_, new_n13999_, new_n14000_, new_n14001_,
    new_n14002_, new_n14003_, new_n14004_, new_n14005_, new_n14006_,
    new_n14007_, new_n14008_, new_n14009_, new_n14010_, new_n14011_,
    new_n14012_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14020_, new_n14021_,
    new_n14022_, new_n14023_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14124_, new_n14125_, new_n14126_,
    new_n14127_, new_n14128_, new_n14129_, new_n14130_, new_n14131_,
    new_n14132_, new_n14133_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14139_, new_n14140_, new_n14141_,
    new_n14142_, new_n14143_, new_n14144_, new_n14145_, new_n14146_,
    new_n14147_, new_n14148_, new_n14149_, new_n14150_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14157_, new_n14158_, new_n14159_, new_n14160_, new_n14161_,
    new_n14162_, new_n14163_, new_n14164_, new_n14165_, new_n14166_,
    new_n14167_, new_n14168_, new_n14169_, new_n14170_, new_n14171_,
    new_n14172_, new_n14173_, new_n14174_, new_n14175_, new_n14176_,
    new_n14177_, new_n14178_, new_n14179_, new_n14180_, new_n14181_,
    new_n14182_, new_n14183_, new_n14184_, new_n14185_, new_n14186_,
    new_n14187_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14192_, new_n14193_, new_n14194_, new_n14195_, new_n14196_,
    new_n14197_, new_n14198_, new_n14199_, new_n14200_, new_n14201_,
    new_n14202_, new_n14203_, new_n14204_, new_n14205_, new_n14206_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14211_,
    new_n14212_, new_n14213_, new_n14214_, new_n14215_, new_n14216_,
    new_n14217_, new_n14218_, new_n14219_, new_n14220_, new_n14221_,
    new_n14222_, new_n14223_, new_n14224_, new_n14225_, new_n14226_,
    new_n14227_, new_n14228_, new_n14229_, new_n14230_, new_n14231_,
    new_n14232_, new_n14233_, new_n14234_, new_n14235_, new_n14236_,
    new_n14237_, new_n14238_, new_n14239_, new_n14240_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14252_, new_n14253_, new_n14254_, new_n14255_, new_n14256_,
    new_n14257_, new_n14258_, new_n14259_, new_n14260_, new_n14261_,
    new_n14262_, new_n14263_, new_n14264_, new_n14265_, new_n14266_,
    new_n14267_, new_n14268_, new_n14269_, new_n14270_, new_n14271_,
    new_n14272_, new_n14273_, new_n14274_, new_n14275_, new_n14276_,
    new_n14277_, new_n14278_, new_n14279_, new_n14280_, new_n14281_,
    new_n14282_, new_n14283_, new_n14284_, new_n14285_, new_n14286_,
    new_n14287_, new_n14288_, new_n14289_, new_n14290_, new_n14291_,
    new_n14292_, new_n14293_, new_n14294_, new_n14295_, new_n14296_,
    new_n14297_, new_n14298_, new_n14299_, new_n14300_, new_n14301_,
    new_n14302_, new_n14303_, new_n14304_, new_n14305_, new_n14306_,
    new_n14307_, new_n14308_, new_n14309_, new_n14310_, new_n14311_,
    new_n14312_, new_n14313_, new_n14314_, new_n14315_, new_n14316_,
    new_n14317_, new_n14318_, new_n14319_, new_n14320_, new_n14321_,
    new_n14322_, new_n14323_, new_n14324_, new_n14325_, new_n14326_,
    new_n14327_, new_n14328_, new_n14329_, new_n14330_, new_n14331_,
    new_n14332_, new_n14333_, new_n14334_, new_n14335_, new_n14336_,
    new_n14337_, new_n14338_, new_n14339_, new_n14340_, new_n14341_,
    new_n14342_, new_n14343_, new_n14344_, new_n14345_, new_n14346_,
    new_n14347_, new_n14348_, new_n14349_, new_n14350_, new_n14351_,
    new_n14352_, new_n14353_, new_n14354_, new_n14355_, new_n14356_,
    new_n14357_, new_n14358_, new_n14359_, new_n14360_, new_n14361_,
    new_n14362_, new_n14363_, new_n14364_, new_n14365_, new_n14366_,
    new_n14367_, new_n14368_, new_n14369_, new_n14370_, new_n14371_,
    new_n14372_, new_n14373_, new_n14374_, new_n14375_, new_n14376_,
    new_n14377_, new_n14378_, new_n14379_, new_n14380_, new_n14381_,
    new_n14382_, new_n14383_, new_n14384_, new_n14385_, new_n14386_,
    new_n14387_, new_n14388_, new_n14389_, new_n14390_, new_n14391_,
    new_n14392_, new_n14393_, new_n14394_, new_n14395_, new_n14396_,
    new_n14397_, new_n14398_, new_n14399_, new_n14400_, new_n14401_,
    new_n14402_, new_n14403_, new_n14404_, new_n14405_, new_n14406_,
    new_n14407_, new_n14408_, new_n14409_, new_n14410_, new_n14411_,
    new_n14412_, new_n14413_, new_n14414_, new_n14415_, new_n14416_,
    new_n14417_, new_n14418_, new_n14419_, new_n14420_, new_n14421_,
    new_n14422_, new_n14423_, new_n14425_, new_n14426_, new_n14427_,
    new_n14428_, new_n14429_, new_n14430_, new_n14431_, new_n14432_,
    new_n14433_, new_n14434_, new_n14435_, new_n14436_, new_n14437_,
    new_n14438_, new_n14439_, new_n14440_, new_n14441_, new_n14442_,
    new_n14443_, new_n14444_, new_n14445_, new_n14446_, new_n14447_,
    new_n14448_, new_n14449_, new_n14450_, new_n14451_, new_n14452_,
    new_n14453_, new_n14454_, new_n14455_, new_n14456_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14465_, new_n14466_, new_n14467_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14474_, new_n14475_, new_n14476_, new_n14477_,
    new_n14478_, new_n14479_, new_n14480_, new_n14481_, new_n14482_,
    new_n14483_, new_n14484_, new_n14485_, new_n14486_, new_n14487_,
    new_n14488_, new_n14489_, new_n14490_, new_n14491_, new_n14492_,
    new_n14493_, new_n14494_, new_n14495_, new_n14496_, new_n14497_,
    new_n14498_, new_n14499_, new_n14500_, new_n14501_, new_n14502_,
    new_n14503_, new_n14504_, new_n14505_, new_n14506_, new_n14507_,
    new_n14508_, new_n14509_, new_n14510_, new_n14511_, new_n14512_,
    new_n14513_, new_n14514_, new_n14515_, new_n14516_, new_n14517_,
    new_n14518_, new_n14519_, new_n14520_, new_n14521_, new_n14522_,
    new_n14523_, new_n14524_, new_n14525_, new_n14526_, new_n14527_,
    new_n14528_, new_n14529_, new_n14530_, new_n14531_, new_n14532_,
    new_n14533_, new_n14534_, new_n14535_, new_n14536_, new_n14537_,
    new_n14538_, new_n14539_, new_n14540_, new_n14541_, new_n14542_,
    new_n14543_, new_n14544_, new_n14545_, new_n14546_, new_n14547_,
    new_n14548_, new_n14549_, new_n14550_, new_n14551_, new_n14552_,
    new_n14553_, new_n14554_, new_n14555_, new_n14556_, new_n14557_,
    new_n14558_, new_n14559_, new_n14560_, new_n14561_, new_n14562_,
    new_n14563_, new_n14564_, new_n14565_, new_n14566_, new_n14567_,
    new_n14568_, new_n14569_, new_n14570_, new_n14571_, new_n14572_,
    new_n14573_, new_n14574_, new_n14575_, new_n14576_, new_n14577_,
    new_n14578_, new_n14579_, new_n14580_, new_n14581_, new_n14582_,
    new_n14583_, new_n14584_, new_n14585_, new_n14586_, new_n14587_,
    new_n14588_, new_n14589_, new_n14590_, new_n14591_, new_n14592_,
    new_n14593_, new_n14594_, new_n14595_, new_n14596_, new_n14597_,
    new_n14598_, new_n14599_, new_n14600_, new_n14601_, new_n14602_,
    new_n14603_, new_n14604_, new_n14605_, new_n14606_, new_n14607_,
    new_n14608_, new_n14609_, new_n14610_, new_n14611_, new_n14612_,
    new_n14614_, new_n14615_, new_n14616_, new_n14617_, new_n14618_,
    new_n14619_, new_n14620_, new_n14621_, new_n14622_, new_n14623_,
    new_n14624_, new_n14625_, new_n14626_, new_n14627_, new_n14628_,
    new_n14629_, new_n14630_, new_n14631_, new_n14632_, new_n14633_,
    new_n14634_, new_n14635_, new_n14636_, new_n14637_, new_n14638_,
    new_n14639_, new_n14640_, new_n14641_, new_n14642_, new_n14643_,
    new_n14644_, new_n14645_, new_n14646_, new_n14647_, new_n14648_,
    new_n14649_, new_n14650_, new_n14651_, new_n14652_, new_n14653_,
    new_n14654_, new_n14655_, new_n14656_, new_n14657_, new_n14658_,
    new_n14659_, new_n14660_, new_n14661_, new_n14662_, new_n14663_,
    new_n14664_, new_n14665_, new_n14666_, new_n14667_, new_n14668_,
    new_n14669_, new_n14670_, new_n14671_, new_n14672_, new_n14673_,
    new_n14674_, new_n14675_, new_n14676_, new_n14677_, new_n14678_,
    new_n14679_, new_n14680_, new_n14681_, new_n14682_, new_n14683_,
    new_n14684_, new_n14685_, new_n14686_, new_n14687_, new_n14688_,
    new_n14689_, new_n14690_, new_n14691_, new_n14692_, new_n14693_,
    new_n14694_, new_n14695_, new_n14696_, new_n14697_, new_n14698_,
    new_n14699_, new_n14700_, new_n14701_, new_n14702_, new_n14703_,
    new_n14704_, new_n14705_, new_n14706_, new_n14707_, new_n14708_,
    new_n14710_, new_n14711_, new_n14712_, new_n14713_, new_n14714_,
    new_n14715_, new_n14716_, new_n14717_, new_n14718_, new_n14719_,
    new_n14720_, new_n14721_, new_n14722_, new_n14723_, new_n14724_,
    new_n14725_, new_n14726_, new_n14727_, new_n14728_, new_n14729_,
    new_n14730_, new_n14731_, new_n14732_, new_n14733_, new_n14734_,
    new_n14735_, new_n14736_, new_n14737_, new_n14738_, new_n14739_,
    new_n14740_, new_n14741_, new_n14742_, new_n14743_, new_n14744_,
    new_n14745_, new_n14746_, new_n14747_, new_n14748_, new_n14749_,
    new_n14750_, new_n14751_, new_n14752_, new_n14753_, new_n14754_,
    new_n14755_, new_n14756_, new_n14757_, new_n14758_, new_n14759_,
    new_n14760_, new_n14761_, new_n14762_, new_n14763_, new_n14764_,
    new_n14765_, new_n14766_, new_n14767_, new_n14768_, new_n14769_,
    new_n14770_, new_n14771_, new_n14772_, new_n14773_, new_n14774_,
    new_n14775_, new_n14776_, new_n14777_, new_n14778_, new_n14779_,
    new_n14780_, new_n14781_, new_n14782_, new_n14783_, new_n14784_,
    new_n14785_, new_n14786_, new_n14787_, new_n14788_, new_n14789_,
    new_n14790_, new_n14791_, new_n14792_, new_n14793_, new_n14794_,
    new_n14795_, new_n14796_, new_n14797_, new_n14798_, new_n14799_,
    new_n14800_, new_n14801_, new_n14802_, new_n14803_, new_n14804_,
    new_n14805_, new_n14806_, new_n14807_, new_n14808_, new_n14809_,
    new_n14810_, new_n14811_, new_n14812_, new_n14813_, new_n14814_,
    new_n14815_, new_n14816_, new_n14817_, new_n14818_, new_n14819_,
    new_n14820_, new_n14821_, new_n14822_, new_n14823_, new_n14824_,
    new_n14825_, new_n14826_, new_n14827_, new_n14828_, new_n14829_,
    new_n14830_, new_n14831_, new_n14832_, new_n14833_, new_n14834_,
    new_n14835_, new_n14836_, new_n14837_, new_n14838_, new_n14839_,
    new_n14840_, new_n14841_, new_n14842_, new_n14843_, new_n14844_,
    new_n14845_, new_n14846_, new_n14847_, new_n14848_, new_n14849_,
    new_n14850_, new_n14851_, new_n14852_, new_n14853_, new_n14854_,
    new_n14855_, new_n14856_, new_n14857_, new_n14858_, new_n14859_,
    new_n14860_, new_n14861_, new_n14862_, new_n14863_, new_n14864_,
    new_n14865_, new_n14866_, new_n14867_, new_n14868_, new_n14869_,
    new_n14870_, new_n14871_, new_n14872_, new_n14873_, new_n14874_,
    new_n14875_, new_n14876_, new_n14877_, new_n14878_, new_n14879_,
    new_n14880_, new_n14881_, new_n14882_, new_n14883_, new_n14884_,
    new_n14885_, new_n14886_, new_n14887_, new_n14888_, new_n14889_,
    new_n14890_, new_n14891_, new_n14892_, new_n14893_, new_n14894_,
    new_n14895_, new_n14896_, new_n14897_, new_n14898_, new_n14899_,
    new_n14900_, new_n14901_, new_n14902_, new_n14903_, new_n14904_,
    new_n14905_, new_n14906_, new_n14907_, new_n14909_, new_n14910_,
    new_n14911_, new_n14912_, new_n14913_, new_n14914_, new_n14915_,
    new_n14916_, new_n14917_, new_n14918_, new_n14919_, new_n14920_,
    new_n14921_, new_n14922_, new_n14923_, new_n14924_, new_n14925_,
    new_n14926_, new_n14927_, new_n14928_, new_n14929_, new_n14930_,
    new_n14931_, new_n14932_, new_n14933_, new_n14934_, new_n14935_,
    new_n14936_, new_n14937_, new_n14938_, new_n14939_, new_n14940_,
    new_n14941_, new_n14942_, new_n14943_, new_n14944_, new_n14945_,
    new_n14946_, new_n14947_, new_n14948_, new_n14949_, new_n14950_,
    new_n14951_, new_n14952_, new_n14953_, new_n14954_, new_n14955_,
    new_n14956_, new_n14957_, new_n14958_, new_n14959_, new_n14960_,
    new_n14961_, new_n14962_, new_n14963_, new_n14964_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14976_, new_n14977_, new_n14978_, new_n14979_, new_n14980_,
    new_n14981_, new_n14982_, new_n14983_, new_n14984_, new_n14985_,
    new_n14986_, new_n14987_, new_n14988_, new_n14989_, new_n14990_,
    new_n14991_, new_n14992_, new_n14993_, new_n14994_, new_n14995_,
    new_n14996_, new_n14997_, new_n14998_, new_n14999_, new_n15000_,
    new_n15001_, new_n15002_, new_n15003_, new_n15004_, new_n15005_,
    new_n15006_, new_n15007_, new_n15008_, new_n15009_, new_n15010_,
    new_n15011_, new_n15012_, new_n15013_, new_n15014_, new_n15015_,
    new_n15016_, new_n15017_, new_n15018_, new_n15019_, new_n15020_,
    new_n15021_, new_n15022_, new_n15023_, new_n15024_, new_n15025_,
    new_n15026_, new_n15027_, new_n15028_, new_n15029_, new_n15030_,
    new_n15031_, new_n15032_, new_n15033_, new_n15034_, new_n15035_,
    new_n15036_, new_n15037_, new_n15038_, new_n15039_, new_n15040_,
    new_n15041_, new_n15042_, new_n15043_, new_n15044_, new_n15045_,
    new_n15046_, new_n15047_, new_n15048_, new_n15049_, new_n15050_,
    new_n15051_, new_n15052_, new_n15053_, new_n15054_, new_n15055_,
    new_n15056_, new_n15057_, new_n15058_, new_n15059_, new_n15060_,
    new_n15061_, new_n15062_, new_n15063_, new_n15064_, new_n15065_,
    new_n15066_, new_n15067_, new_n15068_, new_n15069_, new_n15070_,
    new_n15071_, new_n15072_, new_n15073_, new_n15074_, new_n15075_,
    new_n15076_, new_n15077_, new_n15078_, new_n15079_, new_n15080_,
    new_n15081_, new_n15082_, new_n15083_, new_n15084_, new_n15085_,
    new_n15086_, new_n15087_, new_n15088_, new_n15089_, new_n15090_,
    new_n15091_, new_n15092_, new_n15093_, new_n15094_, new_n15095_,
    new_n15096_, new_n15097_, new_n15098_, new_n15099_, new_n15100_,
    new_n15101_, new_n15102_, new_n15103_, new_n15104_, new_n15105_,
    new_n15106_, new_n15107_, new_n15108_, new_n15109_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15115_,
    new_n15116_, new_n15117_, new_n15118_, new_n15119_, new_n15120_,
    new_n15121_, new_n15122_, new_n15123_, new_n15124_, new_n15125_,
    new_n15126_, new_n15127_, new_n15128_, new_n15129_, new_n15130_,
    new_n15131_, new_n15132_, new_n15133_, new_n15134_, new_n15135_,
    new_n15136_, new_n15137_, new_n15138_, new_n15139_, new_n15140_,
    new_n15141_, new_n15142_, new_n15143_, new_n15144_, new_n15145_,
    new_n15147_, new_n15148_, new_n15149_, new_n15150_, new_n15151_,
    new_n15152_, new_n15153_, new_n15154_, new_n15155_, new_n15156_,
    new_n15157_, new_n15158_, new_n15159_, new_n15160_, new_n15161_,
    new_n15162_, new_n15163_, new_n15164_, new_n15165_, new_n15166_,
    new_n15167_, new_n15168_, new_n15169_, new_n15170_, new_n15171_,
    new_n15172_, new_n15173_, new_n15174_, new_n15175_, new_n15176_,
    new_n15177_, new_n15178_, new_n15180_, new_n15181_, new_n15182_,
    new_n15183_, new_n15184_, new_n15185_, new_n15186_, new_n15187_,
    new_n15188_, new_n15189_, new_n15190_, new_n15191_, new_n15192_,
    new_n15193_, new_n15194_, new_n15195_, new_n15196_, new_n15197_,
    new_n15198_, new_n15199_, new_n15200_, new_n15201_, new_n15202_,
    new_n15203_, new_n15204_, new_n15205_, new_n15206_, new_n15207_,
    new_n15208_, new_n15209_, new_n15210_, new_n15211_, new_n15212_,
    new_n15213_, new_n15214_, new_n15215_, new_n15216_, new_n15217_,
    new_n15218_, new_n15219_, new_n15220_, new_n15221_, new_n15222_,
    new_n15223_, new_n15224_, new_n15225_, new_n15226_, new_n15227_,
    new_n15228_, new_n15229_, new_n15230_, new_n15231_, new_n15232_,
    new_n15233_, new_n15234_, new_n15235_, new_n15236_, new_n15237_,
    new_n15238_, new_n15239_, new_n15240_, new_n15241_, new_n15242_,
    new_n15243_, new_n15244_, new_n15245_, new_n15246_, new_n15247_,
    new_n15248_, new_n15249_, new_n15250_, new_n15251_, new_n15252_,
    new_n15253_, new_n15254_, new_n15255_, new_n15256_, new_n15257_,
    new_n15258_, new_n15259_, new_n15260_, new_n15261_, new_n15262_,
    new_n15263_, new_n15264_, new_n15265_, new_n15266_, new_n15267_,
    new_n15268_, new_n15269_, new_n15270_, new_n15271_, new_n15272_,
    new_n15273_, new_n15274_, new_n15275_, new_n15276_, new_n15277_,
    new_n15278_, new_n15279_, new_n15280_, new_n15281_, new_n15282_,
    new_n15283_, new_n15284_, new_n15285_, new_n15286_, new_n15287_,
    new_n15288_, new_n15289_, new_n15290_, new_n15291_, new_n15292_,
    new_n15293_, new_n15294_, new_n15295_, new_n15296_, new_n15297_,
    new_n15298_, new_n15299_, new_n15300_, new_n15301_, new_n15302_,
    new_n15303_, new_n15304_, new_n15305_, new_n15306_, new_n15307_,
    new_n15308_, new_n15309_, new_n15310_, new_n15311_, new_n15312_,
    new_n15313_, new_n15314_, new_n15315_, new_n15316_, new_n15317_,
    new_n15318_, new_n15319_, new_n15320_, new_n15321_, new_n15322_,
    new_n15323_, new_n15324_, new_n15325_, new_n15327_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15334_,
    new_n15336_, new_n15337_, new_n15338_, new_n15339_, new_n15340_,
    new_n15341_, new_n15342_, new_n15343_, new_n15344_, new_n15345_,
    new_n15346_, new_n15347_, new_n15348_, new_n15349_, new_n15350_,
    new_n15351_, new_n15352_, new_n15353_, new_n15354_, new_n15355_,
    new_n15356_, new_n15357_, new_n15358_, new_n15359_, new_n15360_,
    new_n15361_, new_n15362_, new_n15363_, new_n15364_, new_n15365_,
    new_n15366_, new_n15367_, new_n15368_, new_n15369_, new_n15370_,
    new_n15371_, new_n15372_, new_n15373_, new_n15374_, new_n15375_,
    new_n15376_, new_n15378_, new_n15379_, new_n15380_, new_n15381_,
    new_n15382_, new_n15383_, new_n15384_, new_n15385_, new_n15386_,
    new_n15387_, new_n15388_, new_n15389_, new_n15390_, new_n15391_,
    new_n15392_, new_n15393_, new_n15394_, new_n15395_, new_n15396_,
    new_n15397_, new_n15398_, new_n15399_, new_n15400_, new_n15401_,
    new_n15402_, new_n15403_, new_n15404_, new_n15405_, new_n15406_,
    new_n15407_, new_n15408_, new_n15409_, new_n15410_, new_n15411_,
    new_n15412_, new_n15413_, new_n15414_, new_n15415_, new_n15416_,
    new_n15417_, new_n15418_, new_n15419_, new_n15420_, new_n15421_,
    new_n15422_, new_n15423_, new_n15424_, new_n15425_, new_n15426_,
    new_n15427_, new_n15428_, new_n15429_, new_n15430_, new_n15431_,
    new_n15432_, new_n15433_, new_n15435_, new_n15436_, new_n15437_,
    new_n15438_, new_n15439_, new_n15440_, new_n15441_, new_n15442_,
    new_n15443_, new_n15444_, new_n15445_, new_n15446_, new_n15447_,
    new_n15448_, new_n15449_, new_n15450_, new_n15451_, new_n15452_,
    new_n15453_, new_n15454_, new_n15455_, new_n15456_, new_n15457_,
    new_n15458_, new_n15459_, new_n15460_, new_n15461_, new_n15462_,
    new_n15463_, new_n15464_, new_n15465_, new_n15466_, new_n15467_,
    new_n15468_, new_n15469_, new_n15470_, new_n15471_, new_n15472_,
    new_n15473_, new_n15474_, new_n15475_, new_n15476_, new_n15477_,
    new_n15478_, new_n15479_, new_n15480_, new_n15481_, new_n15482_,
    new_n15483_, new_n15484_, new_n15485_, new_n15486_, new_n15487_,
    new_n15488_, new_n15489_, new_n15490_, new_n15491_, new_n15492_,
    new_n15493_, new_n15494_, new_n15495_, new_n15496_, new_n15497_,
    new_n15498_, new_n15499_, new_n15500_, new_n15501_, new_n15502_,
    new_n15503_, new_n15504_, new_n15505_, new_n15506_, new_n15507_,
    new_n15508_, new_n15509_, new_n15510_, new_n15511_, new_n15512_,
    new_n15513_, new_n15514_, new_n15515_, new_n15516_, new_n15517_,
    new_n15518_, new_n15519_, new_n15520_, new_n15521_, new_n15522_,
    new_n15523_, new_n15524_, new_n15525_, new_n15526_, new_n15527_,
    new_n15528_, new_n15529_, new_n15530_, new_n15531_, new_n15532_,
    new_n15534_, new_n15535_, new_n15536_, new_n15537_, new_n15538_,
    new_n15539_, new_n15540_, new_n15541_, new_n15542_, new_n15543_,
    new_n15544_, new_n15545_, new_n15546_, new_n15547_, new_n15548_,
    new_n15549_, new_n15550_, new_n15551_, new_n15552_, new_n15553_,
    new_n15554_, new_n15555_, new_n15556_, new_n15557_, new_n15558_,
    new_n15559_, new_n15560_, new_n15561_, new_n15562_, new_n15563_,
    new_n15564_, new_n15565_, new_n15566_, new_n15567_, new_n15568_,
    new_n15569_, new_n15570_, new_n15571_, new_n15572_, new_n15573_,
    new_n15574_, new_n15575_, new_n15576_, new_n15577_, new_n15578_,
    new_n15579_, new_n15580_, new_n15581_, new_n15582_, new_n15583_,
    new_n15584_, new_n15585_, new_n15586_, new_n15587_, new_n15588_,
    new_n15589_, new_n15590_, new_n15591_, new_n15592_, new_n15593_,
    new_n15594_, new_n15595_, new_n15596_, new_n15597_, new_n15598_,
    new_n15599_, new_n15600_, new_n15601_, new_n15602_, new_n15603_,
    new_n15604_, new_n15605_, new_n15606_, new_n15607_, new_n15608_,
    new_n15609_, new_n15610_, new_n15611_, new_n15612_, new_n15613_,
    new_n15614_, new_n15615_, new_n15616_, new_n15617_, new_n15618_,
    new_n15619_, new_n15620_, new_n15621_, new_n15622_, new_n15623_,
    new_n15624_, new_n15625_, new_n15626_, new_n15627_, new_n15628_,
    new_n15629_, new_n15630_, new_n15631_, new_n15632_, new_n15633_,
    new_n15634_, new_n15635_, new_n15636_, new_n15637_, new_n15638_,
    new_n15639_, new_n15640_, new_n15641_, new_n15642_, new_n15643_,
    new_n15644_, new_n15645_, new_n15646_, new_n15647_, new_n15648_,
    new_n15649_, new_n15650_, new_n15651_, new_n15652_, new_n15653_,
    new_n15654_, new_n15655_, new_n15656_, new_n15657_, new_n15658_,
    new_n15659_, new_n15660_, new_n15661_, new_n15662_, new_n15663_,
    new_n15664_, new_n15665_, new_n15666_, new_n15667_, new_n15668_,
    new_n15669_, new_n15670_, new_n15671_, new_n15672_, new_n15673_,
    new_n15674_, new_n15675_, new_n15676_, new_n15677_, new_n15678_,
    new_n15679_, new_n15680_, new_n15681_, new_n15682_, new_n15683_,
    new_n15684_, new_n15685_, new_n15686_, new_n15687_, new_n15688_,
    new_n15689_, new_n15690_, new_n15691_, new_n15692_, new_n15693_,
    new_n15694_, new_n15695_, new_n15696_, new_n15697_, new_n15698_,
    new_n15699_, new_n15700_, new_n15701_, new_n15702_, new_n15703_,
    new_n15704_, new_n15705_, new_n15706_, new_n15707_, new_n15708_,
    new_n15709_, new_n15710_, new_n15711_, new_n15712_, new_n15713_,
    new_n15714_, new_n15715_, new_n15716_, new_n15718_, new_n15719_,
    new_n15720_, new_n15721_, new_n15722_, new_n15723_, new_n15724_,
    new_n15725_, new_n15726_, new_n15727_, new_n15728_, new_n15729_,
    new_n15730_, new_n15731_, new_n15732_, new_n15733_, new_n15734_,
    new_n15735_, new_n15736_, new_n15737_, new_n15738_, new_n15739_,
    new_n15740_, new_n15741_, new_n15742_, new_n15743_, new_n15744_,
    new_n15745_, new_n15746_, new_n15747_, new_n15748_, new_n15749_,
    new_n15750_, new_n15751_, new_n15752_, new_n15753_, new_n15754_,
    new_n15755_, new_n15756_, new_n15757_, new_n15758_, new_n15759_,
    new_n15760_, new_n15761_, new_n15762_, new_n15763_, new_n15764_,
    new_n15765_, new_n15766_, new_n15767_, new_n15768_, new_n15769_,
    new_n15770_, new_n15771_, new_n15772_, new_n15773_, new_n15774_,
    new_n15775_, new_n15776_, new_n15777_, new_n15778_, new_n15779_,
    new_n15780_, new_n15781_, new_n15782_, new_n15783_, new_n15784_,
    new_n15785_, new_n15786_, new_n15787_, new_n15788_, new_n15789_,
    new_n15790_, new_n15791_, new_n15792_, new_n15793_, new_n15794_,
    new_n15795_, new_n15796_, new_n15797_, new_n15798_, new_n15799_,
    new_n15800_, new_n15801_, new_n15802_, new_n15803_, new_n15804_,
    new_n15805_, new_n15806_, new_n15807_, new_n15808_, new_n15809_,
    new_n15810_, new_n15811_, new_n15812_, new_n15813_, new_n15814_,
    new_n15815_, new_n15816_, new_n15817_, new_n15818_, new_n15819_,
    new_n15820_, new_n15821_, new_n15822_, new_n15823_, new_n15824_,
    new_n15825_, new_n15826_, new_n15827_, new_n15828_, new_n15829_,
    new_n15830_, new_n15831_, new_n15832_, new_n15833_, new_n15834_,
    new_n15835_, new_n15836_, new_n15837_, new_n15838_, new_n15839_,
    new_n15840_, new_n15841_, new_n15842_, new_n15843_, new_n15844_,
    new_n15845_, new_n15846_, new_n15847_, new_n15848_, new_n15849_,
    new_n15850_, new_n15851_, new_n15852_, new_n15853_, new_n15854_,
    new_n15855_, new_n15856_, new_n15857_, new_n15858_, new_n15859_,
    new_n15860_, new_n15861_, new_n15862_, new_n15863_, new_n15864_,
    new_n15865_, new_n15866_, new_n15867_, new_n15868_, new_n15869_,
    new_n15870_, new_n15871_, new_n15872_, new_n15873_, new_n15874_,
    new_n15875_, new_n15876_, new_n15877_, new_n15878_, new_n15879_,
    new_n15880_, new_n15881_, new_n15882_, new_n15883_, new_n15884_,
    new_n15885_, new_n15886_, new_n15887_, new_n15888_, new_n15889_,
    new_n15890_, new_n15891_, new_n15892_, new_n15893_, new_n15894_,
    new_n15895_, new_n15896_, new_n15898_, new_n15899_, new_n15900_,
    new_n15901_, new_n15902_, new_n15903_, new_n15904_, new_n15905_,
    new_n15906_, new_n15907_, new_n15908_, new_n15909_, new_n15910_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15916_, new_n15917_, new_n15918_, new_n15919_, new_n15920_,
    new_n15921_, new_n15922_, new_n15923_, new_n15924_, new_n15925_,
    new_n15926_, new_n15927_, new_n15928_, new_n15929_, new_n15930_,
    new_n15931_, new_n15932_, new_n15933_, new_n15934_, new_n15935_,
    new_n15936_, new_n15937_, new_n15938_, new_n15939_, new_n15940_,
    new_n15941_, new_n15942_, new_n15943_, new_n15944_, new_n15945_,
    new_n15946_, new_n15947_, new_n15948_, new_n15949_, new_n15950_,
    new_n15951_, new_n15952_, new_n15953_, new_n15954_, new_n15955_,
    new_n15956_, new_n15957_, new_n15958_, new_n15959_, new_n15960_,
    new_n15961_, new_n15962_, new_n15963_, new_n15964_, new_n15965_,
    new_n15966_, new_n15967_, new_n15968_, new_n15969_, new_n15970_,
    new_n15971_, new_n15972_, new_n15973_, new_n15974_, new_n15975_,
    new_n15976_, new_n15977_, new_n15978_, new_n15979_, new_n15980_,
    new_n15981_, new_n15982_, new_n15983_, new_n15984_, new_n15985_,
    new_n15986_, new_n15987_, new_n15988_, new_n15989_, new_n15990_,
    new_n15991_, new_n15992_, new_n15993_, new_n15994_, new_n15995_,
    new_n15996_, new_n15997_, new_n15998_, new_n15999_, new_n16000_,
    new_n16001_, new_n16002_, new_n16003_, new_n16004_, new_n16005_,
    new_n16006_, new_n16007_, new_n16008_, new_n16009_, new_n16010_,
    new_n16011_, new_n16012_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16031_, new_n16032_, new_n16033_, new_n16034_, new_n16035_,
    new_n16036_, new_n16037_, new_n16038_, new_n16039_, new_n16040_,
    new_n16041_, new_n16042_, new_n16043_, new_n16044_, new_n16045_,
    new_n16046_, new_n16047_, new_n16048_, new_n16049_, new_n16050_,
    new_n16051_, new_n16052_, new_n16053_, new_n16054_, new_n16055_,
    new_n16056_, new_n16057_, new_n16058_, new_n16059_, new_n16060_,
    new_n16061_, new_n16062_, new_n16063_, new_n16064_, new_n16065_,
    new_n16066_, new_n16067_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16072_, new_n16073_, new_n16074_, new_n16075_,
    new_n16076_, new_n16077_, new_n16078_, new_n16079_, new_n16080_,
    new_n16081_, new_n16082_, new_n16083_, new_n16084_, new_n16085_,
    new_n16086_, new_n16087_, new_n16088_, new_n16089_, new_n16090_,
    new_n16091_, new_n16092_, new_n16093_, new_n16094_, new_n16095_,
    new_n16096_, new_n16097_, new_n16098_, new_n16099_, new_n16100_,
    new_n16102_, new_n16103_, new_n16104_, new_n16105_, new_n16106_,
    new_n16107_, new_n16108_, new_n16109_, new_n16110_, new_n16111_,
    new_n16112_, new_n16113_, new_n16114_, new_n16115_, new_n16116_,
    new_n16117_, new_n16118_, new_n16119_, new_n16120_, new_n16121_,
    new_n16122_, new_n16123_, new_n16124_, new_n16125_, new_n16126_,
    new_n16127_, new_n16128_, new_n16129_, new_n16130_, new_n16131_,
    new_n16132_, new_n16133_, new_n16134_, new_n16135_, new_n16136_,
    new_n16137_, new_n16138_, new_n16139_, new_n16140_, new_n16141_,
    new_n16142_, new_n16143_, new_n16144_, new_n16145_, new_n16146_,
    new_n16147_, new_n16148_, new_n16149_, new_n16150_, new_n16151_,
    new_n16152_, new_n16153_, new_n16154_, new_n16155_, new_n16156_,
    new_n16157_, new_n16158_, new_n16159_, new_n16160_, new_n16161_,
    new_n16162_, new_n16163_, new_n16164_, new_n16165_, new_n16166_,
    new_n16167_, new_n16168_, new_n16169_, new_n16170_, new_n16171_,
    new_n16172_, new_n16173_, new_n16174_, new_n16175_, new_n16176_,
    new_n16177_, new_n16178_, new_n16179_, new_n16180_, new_n16181_,
    new_n16182_, new_n16183_, new_n16184_, new_n16185_, new_n16186_,
    new_n16187_, new_n16188_, new_n16189_, new_n16190_, new_n16191_,
    new_n16192_, new_n16193_, new_n16194_, new_n16195_, new_n16196_,
    new_n16197_, new_n16198_, new_n16199_, new_n16200_, new_n16201_,
    new_n16202_, new_n16203_, new_n16204_, new_n16205_, new_n16206_,
    new_n16207_, new_n16208_, new_n16209_, new_n16210_, new_n16211_,
    new_n16212_, new_n16213_, new_n16214_, new_n16215_, new_n16216_,
    new_n16217_, new_n16218_, new_n16219_, new_n16220_, new_n16221_,
    new_n16222_, new_n16223_, new_n16224_, new_n16225_, new_n16226_,
    new_n16227_, new_n16228_, new_n16229_, new_n16230_, new_n16231_,
    new_n16232_, new_n16233_, new_n16234_, new_n16235_, new_n16236_,
    new_n16237_, new_n16238_, new_n16239_, new_n16240_, new_n16241_,
    new_n16242_, new_n16243_, new_n16244_, new_n16245_, new_n16246_,
    new_n16247_, new_n16248_, new_n16249_, new_n16250_, new_n16251_,
    new_n16252_, new_n16253_, new_n16254_, new_n16255_, new_n16256_,
    new_n16257_, new_n16258_, new_n16259_, new_n16260_, new_n16261_,
    new_n16262_, new_n16263_, new_n16264_, new_n16265_, new_n16266_,
    new_n16267_, new_n16268_, new_n16269_, new_n16270_, new_n16271_,
    new_n16272_, new_n16273_, new_n16274_, new_n16275_, new_n16276_,
    new_n16277_, new_n16278_, new_n16279_, new_n16280_, new_n16281_,
    new_n16282_, new_n16283_, new_n16284_, new_n16285_, new_n16286_,
    new_n16287_, new_n16288_, new_n16289_, new_n16290_, new_n16291_,
    new_n16292_, new_n16293_, new_n16294_, new_n16295_, new_n16296_,
    new_n16297_, new_n16298_, new_n16299_, new_n16300_, new_n16301_,
    new_n16302_, new_n16303_, new_n16304_, new_n16305_, new_n16306_,
    new_n16307_, new_n16309_, new_n16310_, new_n16311_, new_n16312_,
    new_n16313_, new_n16314_, new_n16315_, new_n16316_, new_n16317_,
    new_n16318_, new_n16319_, new_n16320_, new_n16321_, new_n16322_,
    new_n16323_, new_n16324_, new_n16325_, new_n16326_, new_n16327_,
    new_n16328_, new_n16329_, new_n16330_, new_n16331_, new_n16332_,
    new_n16333_, new_n16334_, new_n16335_, new_n16336_, new_n16337_,
    new_n16338_, new_n16339_, new_n16340_, new_n16341_, new_n16342_,
    new_n16343_, new_n16344_, new_n16345_, new_n16346_, new_n16347_,
    new_n16348_, new_n16349_, new_n16350_, new_n16351_, new_n16352_,
    new_n16353_, new_n16354_, new_n16355_, new_n16356_, new_n16357_,
    new_n16358_, new_n16359_, new_n16360_, new_n16361_, new_n16362_,
    new_n16363_, new_n16364_, new_n16365_, new_n16366_, new_n16367_,
    new_n16368_, new_n16369_, new_n16370_, new_n16371_, new_n16372_,
    new_n16373_, new_n16374_, new_n16375_, new_n16376_, new_n16377_,
    new_n16378_, new_n16379_, new_n16380_, new_n16381_, new_n16382_,
    new_n16383_, new_n16384_, new_n16385_, new_n16386_, new_n16387_,
    new_n16388_, new_n16389_, new_n16390_, new_n16391_, new_n16392_,
    new_n16393_, new_n16394_, new_n16395_, new_n16396_, new_n16397_,
    new_n16398_, new_n16399_, new_n16400_, new_n16401_, new_n16402_,
    new_n16403_, new_n16404_, new_n16405_, new_n16406_, new_n16407_,
    new_n16408_, new_n16409_, new_n16410_, new_n16411_, new_n16412_,
    new_n16413_, new_n16414_, new_n16415_, new_n16416_, new_n16417_,
    new_n16418_, new_n16419_, new_n16420_, new_n16421_, new_n16422_,
    new_n16423_, new_n16424_, new_n16425_, new_n16426_, new_n16427_,
    new_n16428_, new_n16429_, new_n16430_, new_n16431_, new_n16432_,
    new_n16433_, new_n16434_, new_n16435_, new_n16436_, new_n16437_,
    new_n16438_, new_n16439_, new_n16440_, new_n16441_, new_n16442_,
    new_n16443_, new_n16444_, new_n16445_, new_n16446_, new_n16447_,
    new_n16448_, new_n16449_, new_n16450_, new_n16451_, new_n16452_,
    new_n16453_, new_n16454_, new_n16455_, new_n16456_, new_n16457_,
    new_n16458_, new_n16459_, new_n16460_, new_n16461_, new_n16462_,
    new_n16463_, new_n16464_, new_n16465_, new_n16466_, new_n16467_,
    new_n16468_, new_n16469_, new_n16470_, new_n16471_, new_n16472_,
    new_n16473_, new_n16474_, new_n16475_, new_n16476_, new_n16477_,
    new_n16478_, new_n16479_, new_n16480_, new_n16481_, new_n16482_,
    new_n16483_, new_n16484_, new_n16485_, new_n16486_, new_n16487_,
    new_n16488_, new_n16489_, new_n16490_, new_n16491_, new_n16492_,
    new_n16493_, new_n16494_, new_n16495_, new_n16496_, new_n16497_,
    new_n16498_, new_n16499_, new_n16500_, new_n16501_, new_n16502_,
    new_n16503_, new_n16504_, new_n16505_, new_n16506_, new_n16507_,
    new_n16508_, new_n16510_, new_n16511_, new_n16512_, new_n16513_,
    new_n16514_, new_n16515_, new_n16516_, new_n16517_, new_n16518_,
    new_n16519_, new_n16520_, new_n16521_, new_n16522_, new_n16523_,
    new_n16524_, new_n16525_, new_n16526_, new_n16527_, new_n16528_,
    new_n16529_, new_n16530_, new_n16531_, new_n16532_, new_n16533_,
    new_n16534_, new_n16535_, new_n16536_, new_n16537_, new_n16538_,
    new_n16539_, new_n16540_, new_n16541_, new_n16542_, new_n16543_,
    new_n16544_, new_n16545_, new_n16546_, new_n16547_, new_n16548_,
    new_n16549_, new_n16550_, new_n16551_, new_n16552_, new_n16553_,
    new_n16554_, new_n16555_, new_n16556_, new_n16557_, new_n16558_,
    new_n16559_, new_n16560_, new_n16561_, new_n16562_, new_n16563_,
    new_n16564_, new_n16565_, new_n16566_, new_n16567_, new_n16568_,
    new_n16569_, new_n16570_, new_n16571_, new_n16572_, new_n16573_,
    new_n16574_, new_n16575_, new_n16576_, new_n16577_, new_n16578_,
    new_n16579_, new_n16580_, new_n16581_, new_n16582_, new_n16583_,
    new_n16584_, new_n16585_, new_n16586_, new_n16587_, new_n16588_,
    new_n16589_, new_n16590_, new_n16591_, new_n16592_, new_n16593_,
    new_n16594_, new_n16595_, new_n16596_, new_n16597_, new_n16598_,
    new_n16599_, new_n16600_, new_n16601_, new_n16602_, new_n16603_,
    new_n16604_, new_n16605_, new_n16606_, new_n16607_, new_n16608_,
    new_n16609_, new_n16610_, new_n16611_, new_n16612_, new_n16613_,
    new_n16614_, new_n16615_, new_n16616_, new_n16617_, new_n16618_,
    new_n16619_, new_n16620_, new_n16621_, new_n16622_, new_n16623_,
    new_n16624_, new_n16625_, new_n16626_, new_n16627_, new_n16628_,
    new_n16629_, new_n16630_, new_n16631_, new_n16632_, new_n16633_,
    new_n16634_, new_n16635_, new_n16636_, new_n16637_, new_n16638_,
    new_n16639_, new_n16640_, new_n16641_, new_n16642_, new_n16643_,
    new_n16644_, new_n16645_, new_n16646_, new_n16647_, new_n16648_,
    new_n16649_, new_n16650_, new_n16651_, new_n16652_, new_n16653_,
    new_n16654_, new_n16655_, new_n16656_, new_n16657_, new_n16658_,
    new_n16659_, new_n16660_, new_n16661_, new_n16662_, new_n16663_,
    new_n16664_, new_n16665_, new_n16666_, new_n16667_, new_n16668_,
    new_n16669_, new_n16670_, new_n16671_, new_n16672_, new_n16673_,
    new_n16674_, new_n16675_, new_n16676_, new_n16677_, new_n16678_,
    new_n16679_, new_n16680_, new_n16681_, new_n16682_, new_n16683_,
    new_n16684_, new_n16685_, new_n16686_, new_n16687_, new_n16688_,
    new_n16689_, new_n16690_, new_n16691_, new_n16692_, new_n16693_,
    new_n16694_, new_n16695_, new_n16696_, new_n16697_, new_n16698_,
    new_n16699_, new_n16700_, new_n16701_, new_n16702_, new_n16703_,
    new_n16704_, new_n16705_, new_n16706_, new_n16707_, new_n16708_,
    new_n16709_, new_n16710_, new_n16711_, new_n16712_, new_n16714_,
    new_n16715_, new_n16716_, new_n16717_, new_n16718_, new_n16719_,
    new_n16720_, new_n16721_, new_n16722_, new_n16723_, new_n16724_,
    new_n16725_, new_n16726_, new_n16727_, new_n16728_, new_n16729_,
    new_n16730_, new_n16731_, new_n16732_, new_n16733_, new_n16734_,
    new_n16735_, new_n16736_, new_n16737_, new_n16738_, new_n16739_,
    new_n16740_, new_n16741_, new_n16742_, new_n16743_, new_n16744_,
    new_n16745_, new_n16746_, new_n16747_, new_n16748_, new_n16749_,
    new_n16750_, new_n16751_, new_n16752_, new_n16753_, new_n16754_,
    new_n16755_, new_n16756_, new_n16757_, new_n16758_, new_n16759_,
    new_n16760_, new_n16761_, new_n16762_, new_n16763_, new_n16764_,
    new_n16765_, new_n16766_, new_n16767_, new_n16768_, new_n16769_,
    new_n16770_, new_n16771_, new_n16772_, new_n16773_, new_n16774_,
    new_n16775_, new_n16776_, new_n16777_, new_n16778_, new_n16779_,
    new_n16780_, new_n16781_, new_n16782_, new_n16783_, new_n16784_,
    new_n16785_, new_n16786_, new_n16787_, new_n16788_, new_n16789_,
    new_n16790_, new_n16791_, new_n16792_, new_n16793_, new_n16794_,
    new_n16795_, new_n16796_, new_n16797_, new_n16798_, new_n16799_,
    new_n16800_, new_n16801_, new_n16802_, new_n16803_, new_n16804_,
    new_n16805_, new_n16806_, new_n16807_, new_n16808_, new_n16809_,
    new_n16810_, new_n16811_, new_n16812_, new_n16813_, new_n16814_,
    new_n16815_, new_n16816_, new_n16817_, new_n16818_, new_n16819_,
    new_n16820_, new_n16821_, new_n16822_, new_n16823_, new_n16824_,
    new_n16825_, new_n16826_, new_n16827_, new_n16828_, new_n16829_,
    new_n16830_, new_n16831_, new_n16832_, new_n16833_, new_n16834_,
    new_n16835_, new_n16836_, new_n16837_, new_n16838_, new_n16839_,
    new_n16840_, new_n16841_, new_n16842_, new_n16843_, new_n16844_,
    new_n16845_, new_n16846_, new_n16847_, new_n16848_, new_n16849_,
    new_n16850_, new_n16851_, new_n16852_, new_n16853_, new_n16854_,
    new_n16855_, new_n16856_, new_n16857_, new_n16858_, new_n16859_,
    new_n16860_, new_n16861_, new_n16863_, new_n16864_, new_n16865_,
    new_n16866_, new_n16867_, new_n16868_, new_n16869_, new_n16870_,
    new_n16871_, new_n16872_, new_n16873_, new_n16874_, new_n16875_,
    new_n16876_, new_n16877_, new_n16878_, new_n16879_, new_n16880_,
    new_n16881_, new_n16882_, new_n16883_, new_n16884_, new_n16885_,
    new_n16886_, new_n16887_, new_n16888_, new_n16889_, new_n16890_,
    new_n16891_, new_n16892_, new_n16893_, new_n16894_, new_n16895_,
    new_n16896_, new_n16897_, new_n16898_, new_n16899_, new_n16900_,
    new_n16901_, new_n16902_, new_n16903_, new_n16904_, new_n16905_,
    new_n16906_, new_n16907_, new_n16908_, new_n16909_, new_n16910_,
    new_n16911_, new_n16912_, new_n16913_, new_n16914_, new_n16915_,
    new_n16916_, new_n16917_, new_n16918_, new_n16919_, new_n16920_,
    new_n16921_, new_n16922_, new_n16923_, new_n16924_, new_n16925_,
    new_n16926_, new_n16927_, new_n16928_, new_n16929_, new_n16930_,
    new_n16931_, new_n16932_, new_n16933_, new_n16934_, new_n16935_,
    new_n16936_, new_n16937_, new_n16938_, new_n16939_, new_n16940_,
    new_n16942_, new_n16943_, new_n16944_, new_n16945_, new_n16946_,
    new_n16947_, new_n16948_, new_n16949_, new_n16950_, new_n16951_,
    new_n16952_, new_n16953_, new_n16954_, new_n16955_, new_n16956_,
    new_n16957_, new_n16958_, new_n16959_, new_n16960_, new_n16961_,
    new_n16962_, new_n16963_, new_n16964_, new_n16965_, new_n16966_,
    new_n16967_, new_n16968_, new_n16969_, new_n16970_, new_n16971_,
    new_n16972_, new_n16973_, new_n16974_, new_n16975_, new_n16976_,
    new_n16977_, new_n16978_, new_n16979_, new_n16980_, new_n16981_,
    new_n16982_, new_n16983_, new_n16984_, new_n16985_, new_n16986_,
    new_n16987_, new_n16988_, new_n16989_, new_n16990_, new_n16991_,
    new_n16992_, new_n16993_, new_n16994_, new_n16995_, new_n16996_,
    new_n16997_, new_n16998_, new_n16999_, new_n17000_, new_n17001_,
    new_n17002_, new_n17003_, new_n17004_, new_n17005_, new_n17006_,
    new_n17007_, new_n17008_, new_n17009_, new_n17010_, new_n17012_,
    new_n17013_, new_n17014_, new_n17015_, new_n17016_, new_n17017_,
    new_n17018_, new_n17019_, new_n17020_, new_n17021_, new_n17022_,
    new_n17023_, new_n17024_, new_n17025_, new_n17026_, new_n17027_,
    new_n17028_, new_n17029_, new_n17030_, new_n17031_, new_n17032_,
    new_n17033_, new_n17034_, new_n17035_, new_n17036_, new_n17037_,
    new_n17038_, new_n17039_, new_n17040_, new_n17041_, new_n17042_,
    new_n17043_, new_n17044_, new_n17045_, new_n17046_, new_n17047_,
    new_n17048_, new_n17049_, new_n17050_, new_n17051_, new_n17052_,
    new_n17053_, new_n17054_, new_n17055_, new_n17056_, new_n17057_,
    new_n17058_, new_n17059_, new_n17060_, new_n17061_, new_n17062_,
    new_n17063_, new_n17064_, new_n17065_, new_n17066_, new_n17067_,
    new_n17068_, new_n17069_, new_n17070_, new_n17071_, new_n17072_,
    new_n17073_, new_n17074_, new_n17075_, new_n17076_, new_n17077_,
    new_n17078_, new_n17079_, new_n17080_, new_n17081_, new_n17082_,
    new_n17083_, new_n17084_, new_n17085_, new_n17086_, new_n17087_,
    new_n17088_, new_n17089_, new_n17090_, new_n17091_, new_n17092_,
    new_n17093_, new_n17094_, new_n17095_, new_n17096_, new_n17097_,
    new_n17098_, new_n17099_, new_n17100_, new_n17101_, new_n17102_,
    new_n17103_, new_n17104_, new_n17105_, new_n17106_, new_n17107_,
    new_n17108_, new_n17109_, new_n17110_, new_n17111_, new_n17112_,
    new_n17113_, new_n17114_, new_n17115_, new_n17116_, new_n17117_,
    new_n17118_, new_n17119_, new_n17120_, new_n17121_, new_n17122_,
    new_n17123_, new_n17124_, new_n17125_, new_n17126_, new_n17127_,
    new_n17128_, new_n17129_, new_n17130_, new_n17131_, new_n17132_,
    new_n17133_, new_n17134_, new_n17135_, new_n17136_, new_n17137_,
    new_n17138_, new_n17139_, new_n17140_, new_n17141_, new_n17142_,
    new_n17143_, new_n17144_, new_n17145_, new_n17146_, new_n17147_,
    new_n17148_, new_n17149_, new_n17150_, new_n17151_, new_n17152_,
    new_n17153_, new_n17154_, new_n17155_, new_n17156_, new_n17157_,
    new_n17158_, new_n17159_, new_n17160_, new_n17161_, new_n17162_,
    new_n17163_, new_n17164_, new_n17165_, new_n17166_, new_n17167_,
    new_n17168_, new_n17169_, new_n17170_, new_n17171_, new_n17172_,
    new_n17173_, new_n17174_, new_n17175_, new_n17176_, new_n17177_,
    new_n17178_, new_n17179_, new_n17180_, new_n17181_, new_n17182_,
    new_n17184_, new_n17185_, new_n17186_, new_n17187_, new_n17188_,
    new_n17189_, new_n17190_, new_n17191_, new_n17192_, new_n17193_,
    new_n17194_, new_n17195_, new_n17196_, new_n17197_, new_n17198_,
    new_n17199_, new_n17200_, new_n17201_, new_n17202_, new_n17203_,
    new_n17204_, new_n17205_, new_n17206_, new_n17207_, new_n17208_,
    new_n17209_, new_n17210_, new_n17211_, new_n17212_, new_n17213_,
    new_n17214_, new_n17215_, new_n17216_, new_n17217_, new_n17218_,
    new_n17219_, new_n17220_, new_n17221_, new_n17222_, new_n17223_,
    new_n17224_, new_n17225_, new_n17226_, new_n17227_, new_n17228_,
    new_n17229_, new_n17230_, new_n17231_, new_n17232_, new_n17233_,
    new_n17234_, new_n17235_, new_n17236_, new_n17237_, new_n17238_,
    new_n17239_, new_n17240_, new_n17241_, new_n17242_, new_n17243_,
    new_n17244_, new_n17245_, new_n17246_, new_n17247_, new_n17248_,
    new_n17249_, new_n17250_, new_n17251_, new_n17252_, new_n17253_,
    new_n17254_, new_n17255_, new_n17256_, new_n17257_, new_n17258_,
    new_n17259_, new_n17260_, new_n17261_, new_n17262_, new_n17263_,
    new_n17264_, new_n17265_, new_n17266_, new_n17267_, new_n17268_,
    new_n17269_, new_n17270_, new_n17271_, new_n17272_, new_n17273_,
    new_n17274_, new_n17275_, new_n17276_, new_n17277_, new_n17278_,
    new_n17279_, new_n17280_, new_n17281_, new_n17282_, new_n17283_,
    new_n17284_, new_n17285_, new_n17286_, new_n17287_, new_n17288_,
    new_n17289_, new_n17290_, new_n17291_, new_n17292_, new_n17293_,
    new_n17294_, new_n17295_, new_n17296_, new_n17297_, new_n17298_,
    new_n17299_, new_n17300_, new_n17301_, new_n17302_, new_n17303_,
    new_n17304_, new_n17305_, new_n17306_, new_n17307_, new_n17308_,
    new_n17309_, new_n17310_, new_n17312_, new_n17313_, new_n17314_,
    new_n17315_, new_n17316_, new_n17317_, new_n17318_, new_n17319_,
    new_n17320_, new_n17321_, new_n17322_, new_n17323_, new_n17324_,
    new_n17325_, new_n17326_, new_n17327_, new_n17328_, new_n17329_,
    new_n17330_, new_n17331_, new_n17332_, new_n17333_, new_n17334_,
    new_n17335_, new_n17336_, new_n17337_, new_n17338_, new_n17339_,
    new_n17340_, new_n17341_, new_n17342_, new_n17343_, new_n17344_,
    new_n17345_, new_n17346_, new_n17347_, new_n17348_, new_n17349_,
    new_n17350_, new_n17351_, new_n17352_, new_n17353_, new_n17354_,
    new_n17355_, new_n17356_, new_n17357_, new_n17358_, new_n17359_,
    new_n17360_, new_n17361_, new_n17362_, new_n17363_, new_n17364_,
    new_n17365_, new_n17366_, new_n17367_, new_n17368_, new_n17369_,
    new_n17370_, new_n17371_, new_n17372_, new_n17373_, new_n17374_,
    new_n17375_, new_n17376_, new_n17377_, new_n17378_, new_n17379_,
    new_n17380_, new_n17381_, new_n17382_, new_n17383_, new_n17384_,
    new_n17385_, new_n17386_, new_n17387_, new_n17388_, new_n17389_,
    new_n17390_, new_n17391_, new_n17392_, new_n17393_, new_n17394_,
    new_n17395_, new_n17396_, new_n17397_, new_n17398_, new_n17399_,
    new_n17400_, new_n17401_, new_n17402_, new_n17403_, new_n17404_,
    new_n17405_, new_n17406_, new_n17408_, new_n17409_, new_n17410_,
    new_n17411_, new_n17412_, new_n17413_, new_n17414_, new_n17415_,
    new_n17416_, new_n17417_, new_n17418_, new_n17419_, new_n17420_,
    new_n17421_, new_n17422_, new_n17423_, new_n17424_, new_n17425_,
    new_n17426_, new_n17427_, new_n17428_, new_n17429_, new_n17430_,
    new_n17431_, new_n17432_, new_n17433_, new_n17434_, new_n17435_,
    new_n17436_, new_n17437_, new_n17438_, new_n17439_, new_n17440_,
    new_n17441_, new_n17442_, new_n17443_, new_n17444_, new_n17445_,
    new_n17446_, new_n17447_, new_n17448_, new_n17449_, new_n17450_,
    new_n17451_, new_n17452_, new_n17453_, new_n17454_, new_n17455_,
    new_n17456_, new_n17457_, new_n17458_, new_n17459_, new_n17460_,
    new_n17461_, new_n17462_, new_n17463_, new_n17464_, new_n17465_,
    new_n17466_, new_n17467_, new_n17468_, new_n17469_, new_n17470_,
    new_n17471_, new_n17472_, new_n17473_, new_n17474_, new_n17475_,
    new_n17476_, new_n17477_, new_n17478_, new_n17479_, new_n17480_,
    new_n17481_, new_n17482_, new_n17483_, new_n17484_, new_n17485_,
    new_n17486_, new_n17487_, new_n17488_, new_n17489_, new_n17490_,
    new_n17491_, new_n17492_, new_n17493_, new_n17494_, new_n17495_,
    new_n17496_, new_n17497_, new_n17498_, new_n17499_, new_n17500_,
    new_n17501_, new_n17502_, new_n17503_, new_n17504_, new_n17505_,
    new_n17506_, new_n17507_, new_n17508_, new_n17509_, new_n17511_,
    new_n17512_, new_n17513_, new_n17514_, new_n17515_, new_n17516_,
    new_n17517_, new_n17518_, new_n17519_, new_n17520_, new_n17521_,
    new_n17522_, new_n17523_, new_n17524_, new_n17525_, new_n17526_,
    new_n17527_, new_n17528_, new_n17529_, new_n17530_, new_n17531_,
    new_n17532_, new_n17533_, new_n17534_, new_n17535_, new_n17536_,
    new_n17537_, new_n17538_, new_n17539_, new_n17540_, new_n17541_,
    new_n17542_, new_n17543_, new_n17544_, new_n17545_, new_n17546_,
    new_n17547_, new_n17548_, new_n17549_, new_n17550_, new_n17551_,
    new_n17552_, new_n17553_, new_n17554_, new_n17555_, new_n17556_,
    new_n17557_, new_n17558_, new_n17559_, new_n17560_, new_n17561_,
    new_n17562_, new_n17563_, new_n17564_, new_n17565_, new_n17566_,
    new_n17567_, new_n17568_, new_n17569_, new_n17570_, new_n17571_,
    new_n17572_, new_n17573_, new_n17574_, new_n17575_, new_n17576_,
    new_n17577_, new_n17578_, new_n17579_, new_n17580_, new_n17581_,
    new_n17582_, new_n17583_, new_n17584_, new_n17585_, new_n17586_,
    new_n17587_, new_n17588_, new_n17589_, new_n17590_, new_n17591_,
    new_n17592_, new_n17593_, new_n17594_, new_n17595_, new_n17596_,
    new_n17597_, new_n17598_, new_n17599_, new_n17600_, new_n17601_,
    new_n17602_, new_n17603_, new_n17604_, new_n17605_, new_n17606_,
    new_n17607_, new_n17608_, new_n17609_, new_n17610_, new_n17611_,
    new_n17612_, new_n17613_, new_n17614_, new_n17615_, new_n17616_,
    new_n17617_, new_n17618_, new_n17619_, new_n17620_, new_n17621_,
    new_n17622_, new_n17623_, new_n17624_, new_n17625_, new_n17626_,
    new_n17628_, new_n17629_, new_n17630_, new_n17631_, new_n17632_,
    new_n17633_, new_n17634_, new_n17635_, new_n17636_, new_n17637_,
    new_n17638_, new_n17639_, new_n17640_, new_n17641_, new_n17642_,
    new_n17643_, new_n17644_, new_n17645_, new_n17646_, new_n17647_,
    new_n17648_, new_n17649_, new_n17650_, new_n17651_, new_n17652_,
    new_n17653_, new_n17654_, new_n17655_, new_n17656_, new_n17657_,
    new_n17658_, new_n17659_, new_n17660_, new_n17661_, new_n17662_,
    new_n17663_, new_n17664_, new_n17665_, new_n17666_, new_n17667_,
    new_n17668_, new_n17669_, new_n17670_, new_n17671_, new_n17672_,
    new_n17673_, new_n17674_, new_n17675_, new_n17676_, new_n17677_,
    new_n17678_, new_n17679_, new_n17680_, new_n17681_, new_n17682_,
    new_n17683_, new_n17684_, new_n17685_, new_n17686_, new_n17687_,
    new_n17688_, new_n17689_, new_n17690_, new_n17691_, new_n17692_,
    new_n17693_, new_n17694_, new_n17695_, new_n17696_, new_n17697_,
    new_n17698_, new_n17699_, new_n17700_, new_n17701_, new_n17702_,
    new_n17703_, new_n17704_, new_n17705_, new_n17706_, new_n17707_,
    new_n17708_, new_n17709_, new_n17710_, new_n17712_, new_n17713_,
    new_n17714_, new_n17715_, new_n17716_, new_n17717_, new_n17718_,
    new_n17719_, new_n17720_, new_n17721_, new_n17722_, new_n17723_,
    new_n17724_, new_n17725_, new_n17726_, new_n17727_, new_n17728_,
    new_n17729_, new_n17730_, new_n17731_, new_n17732_, new_n17733_,
    new_n17734_, new_n17735_, new_n17736_, new_n17737_, new_n17738_,
    new_n17739_, new_n17740_, new_n17741_, new_n17742_, new_n17743_,
    new_n17744_, new_n17745_, new_n17746_, new_n17747_, new_n17748_,
    new_n17749_, new_n17750_, new_n17751_, new_n17752_, new_n17753_,
    new_n17754_, new_n17755_, new_n17756_, new_n17757_, new_n17758_,
    new_n17759_, new_n17760_, new_n17761_, new_n17762_, new_n17763_,
    new_n17764_, new_n17765_, new_n17766_, new_n17767_, new_n17768_,
    new_n17769_, new_n17770_, new_n17771_, new_n17772_, new_n17773_,
    new_n17774_, new_n17775_, new_n17776_, new_n17777_, new_n17778_,
    new_n17779_, new_n17780_, new_n17781_, new_n17782_, new_n17783_,
    new_n17784_, new_n17785_, new_n17786_, new_n17787_, new_n17788_,
    new_n17789_, new_n17790_, new_n17791_, new_n17792_, new_n17793_,
    new_n17794_, new_n17795_, new_n17796_, new_n17797_, new_n17798_,
    new_n17799_, new_n17800_, new_n17801_, new_n17803_, new_n17804_,
    new_n17805_, new_n17806_, new_n17807_, new_n17808_, new_n17809_,
    new_n17810_, new_n17811_, new_n17812_, new_n17813_, new_n17814_,
    new_n17815_, new_n17816_, new_n17817_, new_n17818_, new_n17819_,
    new_n17820_, new_n17821_, new_n17822_, new_n17823_, new_n17824_,
    new_n17825_, new_n17826_, new_n17827_, new_n17828_, new_n17829_,
    new_n17830_, new_n17831_, new_n17832_, new_n17833_, new_n17834_,
    new_n17835_, new_n17836_, new_n17837_, new_n17838_, new_n17839_,
    new_n17840_, new_n17841_, new_n17842_, new_n17843_, new_n17844_,
    new_n17845_, new_n17846_, new_n17847_, new_n17848_, new_n17849_,
    new_n17850_, new_n17851_, new_n17852_, new_n17853_, new_n17854_,
    new_n17855_, new_n17856_, new_n17857_, new_n17858_, new_n17859_,
    new_n17860_, new_n17861_, new_n17862_, new_n17863_, new_n17864_,
    new_n17865_, new_n17866_, new_n17867_, new_n17868_, new_n17869_,
    new_n17870_, new_n17871_, new_n17872_, new_n17873_, new_n17874_,
    new_n17875_, new_n17876_, new_n17877_, new_n17878_, new_n17879_,
    new_n17880_, new_n17881_, new_n17882_, new_n17883_, new_n17884_,
    new_n17885_, new_n17886_, new_n17887_, new_n17888_, new_n17889_,
    new_n17890_, new_n17891_, new_n17892_, new_n17893_, new_n17894_,
    new_n17895_, new_n17896_, new_n17897_, new_n17898_, new_n17899_,
    new_n17900_, new_n17901_, new_n17903_, new_n17904_, new_n17905_,
    new_n17906_, new_n17907_, new_n17908_, new_n17909_, new_n17910_,
    new_n17911_, new_n17912_, new_n17913_, new_n17914_, new_n17915_,
    new_n17916_, new_n17917_, new_n17918_, new_n17919_, new_n17920_,
    new_n17921_, new_n17922_, new_n17923_, new_n17924_, new_n17925_,
    new_n17926_, new_n17927_, new_n17928_, new_n17929_, new_n17930_,
    new_n17931_, new_n17932_, new_n17933_, new_n17934_, new_n17935_,
    new_n17936_, new_n17937_, new_n17938_, new_n17939_, new_n17940_,
    new_n17941_, new_n17942_, new_n17943_, new_n17944_, new_n17945_,
    new_n17946_, new_n17947_, new_n17948_, new_n17949_, new_n17950_,
    new_n17951_, new_n17952_, new_n17953_, new_n17954_, new_n17955_,
    new_n17956_, new_n17957_, new_n17958_, new_n17959_, new_n17960_,
    new_n17961_, new_n17962_, new_n17963_, new_n17964_, new_n17965_,
    new_n17966_, new_n17967_, new_n17968_, new_n17969_, new_n17970_,
    new_n17971_, new_n17972_, new_n17973_, new_n17975_, new_n17976_,
    new_n17977_, new_n17978_, new_n17979_, new_n17980_, new_n17981_,
    new_n17982_, new_n17983_, new_n17984_, new_n17985_, new_n17986_,
    new_n17987_, new_n17988_, new_n17989_, new_n17990_, new_n17991_,
    new_n17992_, new_n17993_, new_n17994_, new_n17995_, new_n17996_,
    new_n17997_, new_n17998_, new_n17999_, new_n18000_, new_n18001_,
    new_n18002_, new_n18003_, new_n18004_, new_n18005_, new_n18006_,
    new_n18007_, new_n18008_, new_n18009_, new_n18010_, new_n18011_,
    new_n18012_, new_n18013_, new_n18014_, new_n18015_, new_n18016_,
    new_n18017_, new_n18018_, new_n18019_, new_n18020_, new_n18021_,
    new_n18022_, new_n18023_, new_n18024_, new_n18025_, new_n18026_,
    new_n18027_, new_n18028_, new_n18029_, new_n18030_, new_n18031_,
    new_n18032_, new_n18033_, new_n18034_, new_n18035_, new_n18036_,
    new_n18037_, new_n18038_, new_n18039_, new_n18040_, new_n18041_,
    new_n18042_, new_n18043_, new_n18045_, new_n18046_, new_n18047_,
    new_n18048_, new_n18049_, new_n18050_, new_n18051_, new_n18052_,
    new_n18053_, new_n18054_, new_n18055_, new_n18056_, new_n18057_,
    new_n18058_, new_n18059_, new_n18060_, new_n18061_, new_n18062_,
    new_n18063_, new_n18064_, new_n18065_, new_n18066_, new_n18067_,
    new_n18068_, new_n18069_, new_n18070_, new_n18071_, new_n18072_,
    new_n18073_, new_n18074_, new_n18075_, new_n18076_, new_n18077_,
    new_n18078_, new_n18079_, new_n18080_, new_n18081_, new_n18082_,
    new_n18083_, new_n18084_, new_n18085_, new_n18086_, new_n18087_,
    new_n18088_, new_n18089_, new_n18090_, new_n18091_, new_n18092_,
    new_n18093_, new_n18094_, new_n18095_, new_n18096_, new_n18097_,
    new_n18098_, new_n18099_, new_n18100_, new_n18101_, new_n18102_,
    new_n18103_, new_n18104_, new_n18105_, new_n18106_, new_n18107_,
    new_n18108_, new_n18109_, new_n18110_, new_n18111_, new_n18112_,
    new_n18113_, new_n18114_, new_n18115_, new_n18116_, new_n18117_,
    new_n18118_, new_n18119_, new_n18120_, new_n18121_, new_n18122_,
    new_n18123_, new_n18124_, new_n18125_, new_n18126_, new_n18127_,
    new_n18128_, new_n18129_, new_n18130_, new_n18131_, new_n18132_,
    new_n18133_, new_n18134_, new_n18136_, new_n18137_, new_n18138_,
    new_n18139_, new_n18140_, new_n18141_, new_n18142_, new_n18143_,
    new_n18144_, new_n18145_, new_n18146_, new_n18147_, new_n18148_,
    new_n18149_, new_n18150_, new_n18151_, new_n18152_, new_n18153_,
    new_n18154_, new_n18155_, new_n18156_, new_n18157_, new_n18158_,
    new_n18159_, new_n18160_, new_n18161_, new_n18162_, new_n18163_,
    new_n18164_, new_n18165_, new_n18166_, new_n18167_, new_n18168_,
    new_n18169_, new_n18170_, new_n18171_, new_n18172_, new_n18173_,
    new_n18174_, new_n18175_, new_n18176_, new_n18177_, new_n18178_,
    new_n18179_, new_n18180_, new_n18181_, new_n18182_, new_n18183_,
    new_n18184_, new_n18185_, new_n18186_, new_n18187_, new_n18188_,
    new_n18189_, new_n18190_, new_n18191_, new_n18192_, new_n18193_,
    new_n18194_, new_n18195_, new_n18196_, new_n18197_, new_n18198_,
    new_n18199_, new_n18200_, new_n18201_, new_n18202_, new_n18203_,
    new_n18204_, new_n18206_, new_n18207_, new_n18208_, new_n18209_,
    new_n18210_, new_n18211_, new_n18212_, new_n18213_, new_n18214_,
    new_n18215_, new_n18216_, new_n18217_, new_n18218_, new_n18219_,
    new_n18220_, new_n18221_, new_n18222_, new_n18223_, new_n18224_,
    new_n18225_, new_n18226_, new_n18227_, new_n18228_, new_n18229_,
    new_n18230_, new_n18231_, new_n18232_, new_n18233_, new_n18234_,
    new_n18235_, new_n18236_, new_n18237_, new_n18238_, new_n18239_,
    new_n18240_, new_n18241_, new_n18242_, new_n18243_, new_n18244_,
    new_n18245_, new_n18246_, new_n18247_, new_n18248_, new_n18249_,
    new_n18250_, new_n18251_, new_n18252_, new_n18253_, new_n18254_,
    new_n18255_, new_n18256_, new_n18257_, new_n18258_, new_n18259_,
    new_n18260_, new_n18261_, new_n18262_, new_n18263_, new_n18264_,
    new_n18265_, new_n18266_, new_n18267_, new_n18268_, new_n18270_,
    new_n18271_, new_n18272_, new_n18273_, new_n18274_, new_n18275_,
    new_n18276_, new_n18277_, new_n18278_, new_n18279_, new_n18280_,
    new_n18281_, new_n18282_, new_n18283_, new_n18284_, new_n18285_,
    new_n18286_, new_n18287_, new_n18288_, new_n18289_, new_n18290_,
    new_n18291_, new_n18292_, new_n18293_, new_n18294_, new_n18295_,
    new_n18296_, new_n18297_, new_n18298_, new_n18299_, new_n18300_,
    new_n18301_, new_n18302_, new_n18303_, new_n18304_, new_n18305_,
    new_n18306_, new_n18307_, new_n18308_, new_n18309_, new_n18310_,
    new_n18311_, new_n18312_, new_n18313_, new_n18314_, new_n18315_,
    new_n18316_, new_n18317_, new_n18318_, new_n18319_, new_n18320_,
    new_n18321_, new_n18322_, new_n18323_, new_n18324_, new_n18325_,
    new_n18326_, new_n18327_, new_n18328_, new_n18329_, new_n18330_,
    new_n18331_, new_n18332_, new_n18333_, new_n18334_, new_n18335_,
    new_n18336_, new_n18337_, new_n18339_, new_n18340_, new_n18341_,
    new_n18342_, new_n18343_, new_n18344_, new_n18345_, new_n18346_,
    new_n18347_, new_n18348_, new_n18349_, new_n18350_, new_n18351_,
    new_n18352_, new_n18353_, new_n18354_, new_n18355_, new_n18356_,
    new_n18357_, new_n18358_, new_n18359_, new_n18360_, new_n18361_,
    new_n18362_, new_n18363_, new_n18364_, new_n18365_, new_n18366_,
    new_n18367_, new_n18368_, new_n18369_, new_n18370_, new_n18371_,
    new_n18372_, new_n18373_, new_n18374_, new_n18375_, new_n18376_,
    new_n18377_, new_n18378_, new_n18379_, new_n18380_, new_n18381_,
    new_n18382_, new_n18383_, new_n18384_, new_n18385_, new_n18386_,
    new_n18387_, new_n18388_, new_n18389_, new_n18390_, new_n18391_,
    new_n18392_, new_n18394_, new_n18395_, new_n18396_, new_n18397_,
    new_n18398_, new_n18399_, new_n18400_, new_n18401_, new_n18402_,
    new_n18403_, new_n18404_, new_n18405_, new_n18406_, new_n18407_,
    new_n18408_, new_n18409_, new_n18410_, new_n18411_, new_n18412_,
    new_n18413_, new_n18414_, new_n18415_, new_n18416_, new_n18417_,
    new_n18418_, new_n18419_, new_n18420_, new_n18421_, new_n18422_,
    new_n18423_, new_n18424_, new_n18425_, new_n18426_, new_n18427_,
    new_n18428_, new_n18429_, new_n18430_, new_n18431_, new_n18432_,
    new_n18433_, new_n18434_, new_n18435_, new_n18436_, new_n18437_,
    new_n18438_, new_n18440_, new_n18441_, new_n18442_, new_n18443_,
    new_n18444_, new_n18445_, new_n18446_, new_n18447_, new_n18448_,
    new_n18449_, new_n18450_, new_n18451_, new_n18452_, new_n18453_,
    new_n18454_, new_n18455_, new_n18456_, new_n18457_, new_n18458_,
    new_n18459_, new_n18460_, new_n18461_, new_n18462_, new_n18463_,
    new_n18464_, new_n18465_, new_n18466_, new_n18467_, new_n18468_,
    new_n18469_, new_n18470_, new_n18471_, new_n18472_, new_n18473_,
    new_n18474_, new_n18475_, new_n18476_, new_n18477_, new_n18478_,
    new_n18479_, new_n18480_, new_n18481_, new_n18482_, new_n18483_,
    new_n18484_, new_n18485_, new_n18486_, new_n18487_, new_n18488_,
    new_n18489_, new_n18490_, new_n18492_, new_n18493_, new_n18494_,
    new_n18495_, new_n18496_, new_n18497_, new_n18498_, new_n18499_,
    new_n18500_, new_n18501_, new_n18502_, new_n18503_, new_n18504_,
    new_n18505_, new_n18506_, new_n18507_, new_n18508_, new_n18509_,
    new_n18510_, new_n18511_, new_n18512_, new_n18513_, new_n18514_,
    new_n18515_, new_n18516_, new_n18517_, new_n18518_, new_n18519_,
    new_n18520_, new_n18521_, new_n18522_, new_n18523_, new_n18524_,
    new_n18525_, new_n18526_, new_n18527_;
  INV_X1     g00000(.I(\a[26] ), .ZN(new_n65_));
  INV_X1     g00001(.I(\a[25] ), .ZN(new_n66_));
  NOR2_X1    g00002(.A1(new_n66_), .A2(\a[23] ), .ZN(new_n67_));
  INV_X1     g00003(.I(\a[23] ), .ZN(new_n68_));
  NOR2_X1    g00004(.A1(new_n68_), .A2(\a[25] ), .ZN(new_n69_));
  NOR2_X1    g00005(.A1(new_n67_), .A2(new_n69_), .ZN(new_n70_));
  NOR3_X1    g00006(.A1(new_n70_), .A2(\a[24] ), .A3(new_n65_), .ZN(new_n71_));
  INV_X1     g00007(.I(\a[29] ), .ZN(new_n72_));
  INV_X1     g00008(.I(\a[27] ), .ZN(new_n73_));
  NOR2_X1    g00009(.A1(new_n73_), .A2(\a[29] ), .ZN(new_n74_));
  NOR2_X1    g00010(.A1(new_n72_), .A2(\a[27] ), .ZN(new_n75_));
  INV_X1     g00011(.I(\a[28] ), .ZN(new_n76_));
  NOR2_X1    g00012(.A1(new_n76_), .A2(\a[26] ), .ZN(new_n77_));
  NOR2_X1    g00013(.A1(new_n65_), .A2(\a[28] ), .ZN(new_n78_));
  OAI22_X1   g00014(.A1(new_n74_), .A2(new_n75_), .B1(new_n77_), .B2(new_n78_), .ZN(new_n79_));
  NOR2_X1    g00015(.A1(new_n79_), .A2(new_n72_), .ZN(new_n80_));
  XOR2_X1    g00016(.A1(\a[29] ), .A2(\a[30] ), .Z(new_n81_));
  NAND2_X1   g00017(.A1(new_n81_), .A2(\a[31] ), .ZN(new_n82_));
  INV_X1     g00018(.I(\a[31] ), .ZN(new_n83_));
  INV_X1     g00019(.I(\a[30] ), .ZN(new_n84_));
  NOR2_X1    g00020(.A1(new_n72_), .A2(new_n84_), .ZN(new_n85_));
  INV_X1     g00021(.I(new_n85_), .ZN(new_n86_));
  NOR2_X1    g00022(.A1(new_n86_), .A2(new_n83_), .ZN(new_n87_));
  INV_X1     g00023(.I(new_n87_), .ZN(new_n88_));
  NOR2_X1    g00024(.A1(new_n88_), .A2(new_n82_), .ZN(new_n89_));
  INV_X1     g00025(.I(\a[20] ), .ZN(new_n90_));
  NOR3_X1    g00026(.A1(new_n83_), .A2(\a[29] ), .A3(\a[30] ), .ZN(new_n91_));
  AOI21_X1   g00027(.A1(new_n83_), .A2(new_n85_), .B(new_n91_), .ZN(new_n92_));
  NOR2_X1    g00028(.A1(new_n82_), .A2(new_n92_), .ZN(new_n93_));
  INV_X1     g00029(.I(new_n93_), .ZN(new_n94_));
  NOR2_X1    g00030(.A1(new_n94_), .A2(new_n90_), .ZN(new_n95_));
  NOR2_X1    g00031(.A1(new_n89_), .A2(new_n80_), .ZN(new_n96_));
  NAND2_X1   g00032(.A1(new_n72_), .A2(\a[27] ), .ZN(new_n97_));
  NAND2_X1   g00033(.A1(new_n73_), .A2(\a[29] ), .ZN(new_n98_));
  NAND2_X1   g00034(.A1(new_n65_), .A2(\a[28] ), .ZN(new_n99_));
  NAND2_X1   g00035(.A1(new_n76_), .A2(\a[26] ), .ZN(new_n100_));
  AOI22_X1   g00036(.A1(new_n97_), .A2(new_n98_), .B1(new_n99_), .B2(new_n100_), .ZN(new_n101_));
  NAND2_X1   g00037(.A1(new_n101_), .A2(\a[29] ), .ZN(new_n102_));
  INV_X1     g00038(.I(new_n89_), .ZN(new_n103_));
  NOR2_X1    g00039(.A1(new_n95_), .A2(new_n102_), .ZN(new_n104_));
  NOR2_X1    g00040(.A1(new_n104_), .A2(new_n103_), .ZN(new_n105_));
  NAND2_X1   g00041(.A1(new_n104_), .A2(new_n103_), .ZN(new_n106_));
  INV_X1     g00042(.I(new_n106_), .ZN(new_n107_));
  NOR2_X1    g00043(.A1(new_n107_), .A2(new_n105_), .ZN(new_n108_));
  NOR2_X1    g00044(.A1(new_n108_), .A2(new_n102_), .ZN(new_n109_));
  NOR2_X1    g00045(.A1(new_n109_), .A2(new_n96_), .ZN(new_n110_));
  NOR2_X1    g00046(.A1(new_n110_), .A2(new_n71_), .ZN(new_n111_));
  NAND2_X1   g00047(.A1(new_n65_), .A2(\a[24] ), .ZN(new_n112_));
  INV_X1     g00048(.I(\a[24] ), .ZN(new_n113_));
  NAND2_X1   g00049(.A1(new_n113_), .A2(\a[26] ), .ZN(new_n114_));
  NAND2_X1   g00050(.A1(new_n68_), .A2(\a[25] ), .ZN(new_n115_));
  NAND2_X1   g00051(.A1(new_n66_), .A2(\a[23] ), .ZN(new_n116_));
  AOI22_X1   g00052(.A1(new_n112_), .A2(new_n114_), .B1(new_n115_), .B2(new_n116_), .ZN(new_n117_));
  NAND2_X1   g00053(.A1(new_n117_), .A2(\a[26] ), .ZN(new_n118_));
  XOR2_X1    g00054(.A1(new_n108_), .A2(new_n80_), .Z(new_n119_));
  NOR2_X1    g00055(.A1(new_n119_), .A2(new_n118_), .ZN(new_n120_));
  NOR2_X1    g00056(.A1(new_n120_), .A2(new_n111_), .ZN(new_n121_));
  XOR2_X1    g00057(.A1(new_n95_), .A2(new_n80_), .Z(new_n122_));
  INV_X1     g00058(.I(new_n122_), .ZN(new_n123_));
  NOR2_X1    g00059(.A1(new_n93_), .A2(\a[17] ), .ZN(new_n124_));
  INV_X1     g00060(.I(new_n124_), .ZN(new_n125_));
  INV_X1     g00061(.I(\a[17] ), .ZN(new_n126_));
  NOR2_X1    g00062(.A1(new_n94_), .A2(new_n126_), .ZN(new_n127_));
  AOI21_X1   g00063(.A1(new_n89_), .A2(new_n125_), .B(new_n127_), .ZN(new_n128_));
  INV_X1     g00064(.I(new_n128_), .ZN(new_n129_));
  NOR2_X1    g00065(.A1(new_n129_), .A2(new_n80_), .ZN(new_n130_));
  NOR2_X1    g00066(.A1(new_n130_), .A2(new_n93_), .ZN(new_n131_));
  NOR2_X1    g00067(.A1(new_n128_), .A2(new_n102_), .ZN(new_n132_));
  NOR2_X1    g00068(.A1(new_n131_), .A2(new_n132_), .ZN(new_n133_));
  XOR2_X1    g00069(.A1(new_n93_), .A2(new_n90_), .Z(new_n134_));
  AOI21_X1   g00070(.A1(new_n133_), .A2(new_n94_), .B(new_n134_), .ZN(new_n135_));
  NAND2_X1   g00071(.A1(new_n133_), .A2(new_n94_), .ZN(new_n136_));
  INV_X1     g00072(.I(new_n134_), .ZN(new_n137_));
  NOR2_X1    g00073(.A1(new_n136_), .A2(new_n137_), .ZN(new_n138_));
  NOR2_X1    g00074(.A1(new_n138_), .A2(new_n80_), .ZN(new_n139_));
  NOR2_X1    g00075(.A1(new_n139_), .A2(new_n135_), .ZN(new_n140_));
  NOR2_X1    g00076(.A1(new_n140_), .A2(new_n123_), .ZN(new_n141_));
  NAND2_X1   g00077(.A1(new_n140_), .A2(new_n123_), .ZN(new_n142_));
  AOI21_X1   g00078(.A1(new_n118_), .A2(new_n142_), .B(new_n141_), .ZN(new_n143_));
  NOR2_X1    g00079(.A1(new_n143_), .A2(new_n121_), .ZN(new_n144_));
  AOI21_X1   g00080(.A1(new_n143_), .A2(new_n121_), .B(new_n68_), .ZN(new_n145_));
  INV_X1     g00081(.I(new_n96_), .ZN(new_n146_));
  AOI21_X1   g00082(.A1(new_n118_), .A2(new_n146_), .B(new_n109_), .ZN(new_n147_));
  NOR2_X1    g00083(.A1(new_n89_), .A2(\a[23] ), .ZN(new_n148_));
  NOR2_X1    g00084(.A1(new_n103_), .A2(new_n68_), .ZN(new_n149_));
  NOR2_X1    g00085(.A1(new_n149_), .A2(new_n148_), .ZN(new_n150_));
  INV_X1     g00086(.I(new_n150_), .ZN(new_n151_));
  NOR2_X1    g00087(.A1(new_n151_), .A2(new_n80_), .ZN(new_n152_));
  NOR2_X1    g00088(.A1(new_n150_), .A2(new_n102_), .ZN(new_n153_));
  NOR2_X1    g00089(.A1(new_n152_), .A2(new_n153_), .ZN(new_n154_));
  NOR2_X1    g00090(.A1(new_n154_), .A2(new_n107_), .ZN(new_n155_));
  NOR4_X1    g00091(.A1(new_n95_), .A2(new_n68_), .A3(new_n102_), .A4(new_n89_), .ZN(new_n156_));
  NOR2_X1    g00092(.A1(new_n155_), .A2(new_n156_), .ZN(new_n157_));
  XOR2_X1    g00093(.A1(new_n157_), .A2(new_n71_), .Z(new_n158_));
  NOR2_X1    g00094(.A1(new_n158_), .A2(new_n147_), .ZN(new_n159_));
  INV_X1     g00095(.I(new_n147_), .ZN(new_n160_));
  NOR3_X1    g00096(.A1(new_n155_), .A2(new_n71_), .A3(new_n156_), .ZN(new_n161_));
  NOR2_X1    g00097(.A1(new_n157_), .A2(new_n118_), .ZN(new_n162_));
  NOR2_X1    g00098(.A1(new_n162_), .A2(new_n161_), .ZN(new_n163_));
  NOR2_X1    g00099(.A1(new_n163_), .A2(new_n160_), .ZN(new_n164_));
  NOR2_X1    g00100(.A1(new_n159_), .A2(new_n164_), .ZN(new_n165_));
  NOR3_X1    g00101(.A1(new_n145_), .A2(new_n144_), .A3(new_n165_), .ZN(new_n166_));
  NOR2_X1    g00102(.A1(new_n161_), .A2(new_n147_), .ZN(new_n167_));
  NOR2_X1    g00103(.A1(new_n153_), .A2(new_n107_), .ZN(new_n168_));
  NOR2_X1    g00104(.A1(new_n168_), .A2(new_n152_), .ZN(new_n169_));
  NOR2_X1    g00105(.A1(new_n149_), .A2(new_n93_), .ZN(new_n170_));
  INV_X1     g00106(.I(new_n149_), .ZN(new_n171_));
  NOR2_X1    g00107(.A1(new_n171_), .A2(new_n94_), .ZN(new_n172_));
  OAI21_X1   g00108(.A1(new_n172_), .A2(new_n170_), .B(new_n102_), .ZN(new_n173_));
  NOR2_X1    g00109(.A1(new_n149_), .A2(new_n94_), .ZN(new_n174_));
  NOR2_X1    g00110(.A1(new_n171_), .A2(new_n93_), .ZN(new_n175_));
  OAI21_X1   g00111(.A1(new_n175_), .A2(new_n174_), .B(new_n80_), .ZN(new_n176_));
  NAND2_X1   g00112(.A1(new_n173_), .A2(new_n176_), .ZN(new_n177_));
  XNOR2_X1   g00113(.A1(new_n177_), .A2(new_n169_), .ZN(new_n178_));
  NOR2_X1    g00114(.A1(new_n178_), .A2(new_n118_), .ZN(new_n179_));
  NOR2_X1    g00115(.A1(new_n177_), .A2(new_n169_), .ZN(new_n180_));
  INV_X1     g00116(.I(new_n180_), .ZN(new_n181_));
  NAND2_X1   g00117(.A1(new_n177_), .A2(new_n169_), .ZN(new_n182_));
  AOI21_X1   g00118(.A1(new_n181_), .A2(new_n182_), .B(new_n71_), .ZN(new_n183_));
  OAI22_X1   g00119(.A1(new_n179_), .A2(new_n183_), .B1(new_n162_), .B2(new_n167_), .ZN(new_n184_));
  INV_X1     g00120(.I(\a[22] ), .ZN(new_n185_));
  NOR2_X1    g00121(.A1(new_n185_), .A2(\a[20] ), .ZN(new_n186_));
  NOR2_X1    g00122(.A1(new_n90_), .A2(\a[22] ), .ZN(new_n187_));
  NOR2_X1    g00123(.A1(new_n186_), .A2(new_n187_), .ZN(new_n188_));
  NOR3_X1    g00124(.A1(new_n188_), .A2(\a[21] ), .A3(new_n68_), .ZN(new_n189_));
  XOR2_X1    g00125(.A1(new_n133_), .A2(new_n93_), .Z(new_n190_));
  NOR2_X1    g00126(.A1(new_n190_), .A2(new_n102_), .ZN(new_n191_));
  INV_X1     g00127(.I(new_n191_), .ZN(new_n192_));
  NAND2_X1   g00128(.A1(new_n190_), .A2(new_n102_), .ZN(new_n193_));
  AOI21_X1   g00129(.A1(new_n192_), .A2(new_n193_), .B(new_n118_), .ZN(new_n194_));
  XOR2_X1    g00130(.A1(new_n190_), .A2(new_n80_), .Z(new_n195_));
  NOR2_X1    g00131(.A1(new_n195_), .A2(new_n71_), .ZN(new_n196_));
  NOR2_X1    g00132(.A1(new_n129_), .A2(new_n102_), .ZN(new_n197_));
  NOR2_X1    g00133(.A1(new_n128_), .A2(new_n80_), .ZN(new_n198_));
  OAI21_X1   g00134(.A1(new_n197_), .A2(new_n198_), .B(new_n94_), .ZN(new_n199_));
  OAI21_X1   g00135(.A1(new_n130_), .A2(new_n132_), .B(new_n93_), .ZN(new_n200_));
  NAND2_X1   g00136(.A1(new_n199_), .A2(new_n200_), .ZN(new_n201_));
  INV_X1     g00137(.I(new_n201_), .ZN(new_n202_));
  NOR2_X1    g00138(.A1(new_n89_), .A2(new_n94_), .ZN(new_n203_));
  NOR2_X1    g00139(.A1(new_n203_), .A2(new_n102_), .ZN(new_n204_));
  NOR2_X1    g00140(.A1(new_n103_), .A2(new_n93_), .ZN(new_n205_));
  NOR2_X1    g00141(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1     g00142(.I(new_n206_), .ZN(new_n207_));
  NOR2_X1    g00143(.A1(new_n94_), .A2(\a[17] ), .ZN(new_n208_));
  NOR2_X1    g00144(.A1(new_n93_), .A2(new_n126_), .ZN(new_n209_));
  OAI21_X1   g00145(.A1(new_n208_), .A2(new_n209_), .B(new_n89_), .ZN(new_n210_));
  OAI21_X1   g00146(.A1(new_n127_), .A2(new_n124_), .B(new_n103_), .ZN(new_n211_));
  NAND2_X1   g00147(.A1(new_n211_), .A2(new_n210_), .ZN(new_n212_));
  INV_X1     g00148(.I(new_n212_), .ZN(new_n213_));
  NOR2_X1    g00149(.A1(new_n213_), .A2(new_n102_), .ZN(new_n214_));
  INV_X1     g00150(.I(new_n214_), .ZN(new_n215_));
  NOR2_X1    g00151(.A1(new_n212_), .A2(new_n80_), .ZN(new_n216_));
  AOI21_X1   g00152(.A1(new_n215_), .A2(new_n207_), .B(new_n216_), .ZN(new_n217_));
  INV_X1     g00153(.I(new_n217_), .ZN(new_n218_));
  NOR2_X1    g00154(.A1(new_n218_), .A2(new_n202_), .ZN(new_n219_));
  INV_X1     g00155(.I(new_n219_), .ZN(new_n220_));
  NOR2_X1    g00156(.A1(new_n217_), .A2(new_n201_), .ZN(new_n221_));
  AOI21_X1   g00157(.A1(new_n220_), .A2(new_n118_), .B(new_n221_), .ZN(new_n222_));
  INV_X1     g00158(.I(new_n222_), .ZN(new_n223_));
  NOR3_X1    g00159(.A1(new_n196_), .A2(new_n194_), .A3(new_n223_), .ZN(new_n224_));
  NOR2_X1    g00160(.A1(new_n224_), .A2(new_n189_), .ZN(new_n225_));
  NOR2_X1    g00161(.A1(new_n196_), .A2(new_n194_), .ZN(new_n226_));
  NOR2_X1    g00162(.A1(new_n226_), .A2(new_n222_), .ZN(new_n227_));
  NOR2_X1    g00163(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1   g00164(.A1(new_n118_), .A2(new_n191_), .B(new_n193_), .ZN(new_n229_));
  INV_X1     g00165(.I(new_n229_), .ZN(new_n230_));
  XOR2_X1    g00166(.A1(new_n136_), .A2(new_n134_), .Z(new_n231_));
  OAI21_X1   g00167(.A1(new_n138_), .A2(new_n135_), .B(new_n80_), .ZN(new_n232_));
  OAI21_X1   g00168(.A1(new_n231_), .A2(new_n80_), .B(new_n232_), .ZN(new_n233_));
  NOR2_X1    g00169(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1     g00170(.I(new_n234_), .ZN(new_n235_));
  NAND2_X1   g00171(.A1(new_n230_), .A2(new_n233_), .ZN(new_n236_));
  AOI21_X1   g00172(.A1(new_n235_), .A2(new_n236_), .B(new_n71_), .ZN(new_n237_));
  XOR2_X1    g00173(.A1(new_n229_), .A2(new_n233_), .Z(new_n238_));
  NOR2_X1    g00174(.A1(new_n238_), .A2(new_n118_), .ZN(new_n239_));
  NOR3_X1    g00175(.A1(new_n237_), .A2(new_n239_), .A3(new_n189_), .ZN(new_n240_));
  NOR2_X1    g00176(.A1(new_n240_), .A2(new_n228_), .ZN(new_n241_));
  NAND2_X1   g00177(.A1(new_n68_), .A2(\a[21] ), .ZN(new_n242_));
  INV_X1     g00178(.I(\a[21] ), .ZN(new_n243_));
  NAND2_X1   g00179(.A1(new_n243_), .A2(\a[23] ), .ZN(new_n244_));
  NAND2_X1   g00180(.A1(new_n90_), .A2(\a[22] ), .ZN(new_n245_));
  NAND2_X1   g00181(.A1(new_n185_), .A2(\a[20] ), .ZN(new_n246_));
  AOI22_X1   g00182(.A1(new_n242_), .A2(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1   g00183(.A1(new_n247_), .A2(\a[23] ), .ZN(new_n248_));
  NOR2_X1    g00184(.A1(new_n237_), .A2(new_n239_), .ZN(new_n249_));
  NOR2_X1    g00185(.A1(new_n249_), .A2(new_n248_), .ZN(new_n250_));
  NOR2_X1    g00186(.A1(new_n241_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1    g00187(.A1(new_n140_), .A2(new_n122_), .Z(new_n252_));
  NOR2_X1    g00188(.A1(new_n252_), .A2(new_n71_), .ZN(new_n253_));
  INV_X1     g00189(.I(new_n141_), .ZN(new_n254_));
  AOI21_X1   g00190(.A1(new_n254_), .A2(new_n142_), .B(new_n118_), .ZN(new_n255_));
  NOR2_X1    g00191(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1   g00192(.A1(new_n236_), .A2(new_n118_), .ZN(new_n257_));
  NAND2_X1   g00193(.A1(new_n257_), .A2(new_n235_), .ZN(new_n258_));
  NOR2_X1    g00194(.A1(new_n258_), .A2(new_n189_), .ZN(new_n259_));
  INV_X1     g00195(.I(new_n259_), .ZN(new_n260_));
  NAND2_X1   g00196(.A1(new_n258_), .A2(new_n189_), .ZN(new_n261_));
  AOI21_X1   g00197(.A1(new_n260_), .A2(new_n261_), .B(new_n256_), .ZN(new_n262_));
  INV_X1     g00198(.I(new_n256_), .ZN(new_n263_));
  XOR2_X1    g00199(.A1(new_n258_), .A2(new_n248_), .Z(new_n264_));
  NOR2_X1    g00200(.A1(new_n264_), .A2(new_n263_), .ZN(new_n265_));
  NOR2_X1    g00201(.A1(new_n265_), .A2(new_n262_), .ZN(new_n266_));
  NOR2_X1    g00202(.A1(new_n266_), .A2(new_n251_), .ZN(new_n267_));
  INV_X1     g00203(.I(\a[18] ), .ZN(new_n268_));
  NAND2_X1   g00204(.A1(new_n126_), .A2(\a[19] ), .ZN(new_n269_));
  INV_X1     g00205(.I(\a[19] ), .ZN(new_n270_));
  NAND2_X1   g00206(.A1(new_n270_), .A2(\a[17] ), .ZN(new_n271_));
  NAND2_X1   g00207(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1   g00208(.A1(new_n272_), .A2(new_n268_), .A3(\a[20] ), .ZN(new_n273_));
  OAI21_X1   g00209(.A1(new_n205_), .A2(new_n203_), .B(new_n80_), .ZN(new_n274_));
  NOR2_X1    g00210(.A1(new_n89_), .A2(new_n93_), .ZN(new_n275_));
  NOR2_X1    g00211(.A1(new_n103_), .A2(new_n94_), .ZN(new_n276_));
  OAI21_X1   g00212(.A1(new_n276_), .A2(new_n275_), .B(new_n102_), .ZN(new_n277_));
  NAND2_X1   g00213(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1     g00214(.I(\a[14] ), .ZN(new_n279_));
  NOR2_X1    g00215(.A1(new_n103_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1    g00216(.A1(new_n280_), .A2(new_n94_), .ZN(new_n281_));
  INV_X1     g00217(.I(new_n281_), .ZN(new_n282_));
  NOR3_X1    g00218(.A1(new_n103_), .A2(new_n279_), .A3(new_n93_), .ZN(new_n283_));
  AOI21_X1   g00219(.A1(new_n282_), .A2(new_n102_), .B(new_n283_), .ZN(new_n284_));
  INV_X1     g00220(.I(new_n284_), .ZN(new_n285_));
  NOR2_X1    g00221(.A1(new_n285_), .A2(new_n278_), .ZN(new_n286_));
  INV_X1     g00222(.I(new_n278_), .ZN(new_n287_));
  NOR2_X1    g00223(.A1(new_n287_), .A2(new_n284_), .ZN(new_n288_));
  OAI21_X1   g00224(.A1(new_n286_), .A2(new_n288_), .B(new_n118_), .ZN(new_n289_));
  XOR2_X1    g00225(.A1(new_n284_), .A2(new_n278_), .Z(new_n290_));
  OAI21_X1   g00226(.A1(new_n118_), .A2(new_n290_), .B(new_n289_), .ZN(new_n291_));
  NOR2_X1    g00227(.A1(new_n93_), .A2(\a[11] ), .ZN(new_n292_));
  NOR2_X1    g00228(.A1(new_n292_), .A2(new_n94_), .ZN(new_n293_));
  INV_X1     g00229(.I(\a[11] ), .ZN(new_n294_));
  NOR2_X1    g00230(.A1(new_n94_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1    g00231(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1     g00232(.I(new_n296_), .ZN(new_n297_));
  NOR2_X1    g00233(.A1(new_n297_), .A2(new_n103_), .ZN(new_n298_));
  NOR2_X1    g00234(.A1(new_n298_), .A2(new_n80_), .ZN(new_n299_));
  NOR2_X1    g00235(.A1(new_n296_), .A2(new_n89_), .ZN(new_n300_));
  NOR2_X1    g00236(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1   g00237(.A1(new_n301_), .A2(new_n103_), .ZN(new_n302_));
  XOR2_X1    g00238(.A1(new_n89_), .A2(new_n279_), .Z(new_n303_));
  INV_X1     g00239(.I(new_n303_), .ZN(new_n304_));
  NOR2_X1    g00240(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1   g00241(.A1(new_n302_), .A2(new_n304_), .ZN(new_n306_));
  OAI21_X1   g00242(.A1(new_n80_), .A2(new_n305_), .B(new_n306_), .ZN(new_n307_));
  NAND2_X1   g00243(.A1(new_n307_), .A2(new_n71_), .ZN(new_n308_));
  XOR2_X1    g00244(.A1(new_n280_), .A2(new_n93_), .Z(new_n309_));
  OAI21_X1   g00245(.A1(new_n281_), .A2(new_n283_), .B(new_n80_), .ZN(new_n310_));
  OAI21_X1   g00246(.A1(new_n309_), .A2(new_n80_), .B(new_n310_), .ZN(new_n311_));
  NOR2_X1    g00247(.A1(new_n307_), .A2(new_n71_), .ZN(new_n312_));
  OAI21_X1   g00248(.A1(new_n311_), .A2(new_n312_), .B(new_n308_), .ZN(new_n313_));
  NOR2_X1    g00249(.A1(new_n313_), .A2(new_n291_), .ZN(new_n314_));
  NAND2_X1   g00250(.A1(new_n313_), .A2(new_n291_), .ZN(new_n315_));
  INV_X1     g00251(.I(new_n315_), .ZN(new_n316_));
  OAI21_X1   g00252(.A1(new_n316_), .A2(new_n314_), .B(new_n189_), .ZN(new_n317_));
  XNOR2_X1   g00253(.A1(new_n313_), .A2(new_n291_), .ZN(new_n318_));
  OAI21_X1   g00254(.A1(new_n189_), .A2(new_n318_), .B(new_n317_), .ZN(new_n319_));
  XOR2_X1    g00255(.A1(new_n307_), .A2(new_n71_), .Z(new_n320_));
  NAND2_X1   g00256(.A1(new_n320_), .A2(new_n311_), .ZN(new_n321_));
  INV_X1     g00257(.I(new_n308_), .ZN(new_n322_));
  NOR2_X1    g00258(.A1(new_n322_), .A2(new_n312_), .ZN(new_n323_));
  OAI21_X1   g00259(.A1(new_n311_), .A2(new_n323_), .B(new_n321_), .ZN(new_n324_));
  XOR2_X1    g00260(.A1(new_n302_), .A2(new_n303_), .Z(new_n325_));
  NOR2_X1    g00261(.A1(new_n325_), .A2(new_n80_), .ZN(new_n326_));
  INV_X1     g00262(.I(new_n305_), .ZN(new_n327_));
  AOI21_X1   g00263(.A1(new_n327_), .A2(new_n306_), .B(new_n102_), .ZN(new_n328_));
  NOR2_X1    g00264(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  XOR2_X1    g00265(.A1(new_n301_), .A2(new_n89_), .Z(new_n330_));
  NOR2_X1    g00266(.A1(new_n330_), .A2(new_n102_), .ZN(new_n331_));
  INV_X1     g00267(.I(new_n331_), .ZN(new_n332_));
  NAND2_X1   g00268(.A1(new_n330_), .A2(new_n102_), .ZN(new_n333_));
  INV_X1     g00269(.I(new_n333_), .ZN(new_n334_));
  AOI21_X1   g00270(.A1(new_n71_), .A2(new_n332_), .B(new_n334_), .ZN(new_n335_));
  INV_X1     g00271(.I(new_n335_), .ZN(new_n336_));
  NOR2_X1    g00272(.A1(new_n336_), .A2(new_n329_), .ZN(new_n337_));
  INV_X1     g00273(.I(new_n337_), .ZN(new_n338_));
  NOR3_X1    g00274(.A1(new_n335_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n339_));
  AOI21_X1   g00275(.A1(new_n338_), .A2(new_n118_), .B(new_n339_), .ZN(new_n340_));
  INV_X1     g00276(.I(new_n340_), .ZN(new_n341_));
  NOR2_X1    g00277(.A1(new_n341_), .A2(new_n324_), .ZN(new_n342_));
  INV_X1     g00278(.I(new_n342_), .ZN(new_n343_));
  NAND2_X1   g00279(.A1(new_n341_), .A2(new_n324_), .ZN(new_n344_));
  INV_X1     g00280(.I(new_n344_), .ZN(new_n345_));
  AOI21_X1   g00281(.A1(new_n248_), .A2(new_n343_), .B(new_n345_), .ZN(new_n346_));
  INV_X1     g00282(.I(new_n346_), .ZN(new_n347_));
  NOR2_X1    g00283(.A1(new_n347_), .A2(new_n319_), .ZN(new_n348_));
  INV_X1     g00284(.I(new_n348_), .ZN(new_n349_));
  NAND2_X1   g00285(.A1(new_n347_), .A2(new_n319_), .ZN(new_n350_));
  INV_X1     g00286(.I(new_n350_), .ZN(new_n351_));
  AOI21_X1   g00287(.A1(new_n273_), .A2(new_n349_), .B(new_n351_), .ZN(new_n352_));
  NOR2_X1    g00288(.A1(new_n270_), .A2(\a[17] ), .ZN(new_n353_));
  NOR2_X1    g00289(.A1(new_n126_), .A2(\a[19] ), .ZN(new_n354_));
  NOR2_X1    g00290(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NOR3_X1    g00291(.A1(new_n355_), .A2(\a[18] ), .A3(new_n90_), .ZN(new_n356_));
  OAI21_X1   g00292(.A1(new_n248_), .A2(new_n314_), .B(new_n315_), .ZN(new_n357_));
  NOR2_X1    g00293(.A1(new_n286_), .A2(new_n71_), .ZN(new_n358_));
  NOR2_X1    g00294(.A1(new_n358_), .A2(new_n288_), .ZN(new_n359_));
  OAI21_X1   g00295(.A1(new_n214_), .A2(new_n216_), .B(new_n207_), .ZN(new_n360_));
  XOR2_X1    g00296(.A1(new_n212_), .A2(new_n102_), .Z(new_n361_));
  OAI21_X1   g00297(.A1(new_n207_), .A2(new_n361_), .B(new_n360_), .ZN(new_n362_));
  XOR2_X1    g00298(.A1(new_n359_), .A2(new_n362_), .Z(new_n363_));
  NOR2_X1    g00299(.A1(new_n363_), .A2(new_n71_), .ZN(new_n364_));
  INV_X1     g00300(.I(new_n359_), .ZN(new_n365_));
  NOR2_X1    g00301(.A1(new_n365_), .A2(new_n362_), .ZN(new_n366_));
  INV_X1     g00302(.I(new_n366_), .ZN(new_n367_));
  NAND2_X1   g00303(.A1(new_n365_), .A2(new_n362_), .ZN(new_n368_));
  AOI21_X1   g00304(.A1(new_n367_), .A2(new_n368_), .B(new_n118_), .ZN(new_n369_));
  NOR2_X1    g00305(.A1(new_n369_), .A2(new_n364_), .ZN(new_n370_));
  XNOR2_X1   g00306(.A1(new_n357_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1    g00307(.A1(new_n371_), .A2(new_n189_), .ZN(new_n372_));
  INV_X1     g00308(.I(new_n357_), .ZN(new_n373_));
  INV_X1     g00309(.I(new_n370_), .ZN(new_n374_));
  NOR2_X1    g00310(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NOR2_X1    g00311(.A1(new_n357_), .A2(new_n370_), .ZN(new_n376_));
  NOR2_X1    g00312(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NOR2_X1    g00313(.A1(new_n377_), .A2(new_n248_), .ZN(new_n378_));
  NOR2_X1    g00314(.A1(new_n378_), .A2(new_n372_), .ZN(new_n379_));
  NOR2_X1    g00315(.A1(new_n379_), .A2(new_n356_), .ZN(new_n380_));
  NAND2_X1   g00316(.A1(new_n379_), .A2(new_n356_), .ZN(new_n381_));
  OAI21_X1   g00317(.A1(new_n352_), .A2(new_n380_), .B(new_n381_), .ZN(new_n382_));
  INV_X1     g00318(.I(new_n382_), .ZN(new_n383_));
  AOI21_X1   g00319(.A1(new_n349_), .A2(new_n350_), .B(new_n356_), .ZN(new_n384_));
  XOR2_X1    g00320(.A1(new_n346_), .A2(new_n319_), .Z(new_n385_));
  NOR2_X1    g00321(.A1(new_n385_), .A2(new_n273_), .ZN(new_n386_));
  NOR2_X1    g00322(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  AOI21_X1   g00323(.A1(new_n343_), .A2(new_n344_), .B(new_n189_), .ZN(new_n388_));
  XOR2_X1    g00324(.A1(new_n340_), .A2(new_n324_), .Z(new_n389_));
  NOR2_X1    g00325(.A1(new_n389_), .A2(new_n248_), .ZN(new_n390_));
  NOR2_X1    g00326(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1     g00327(.I(new_n391_), .ZN(new_n392_));
  XOR2_X1    g00328(.A1(new_n335_), .A2(new_n329_), .Z(new_n393_));
  OAI21_X1   g00329(.A1(new_n337_), .A2(new_n339_), .B(new_n71_), .ZN(new_n394_));
  OAI21_X1   g00330(.A1(new_n71_), .A2(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1     g00331(.I(new_n395_), .ZN(new_n396_));
  AOI21_X1   g00332(.A1(new_n332_), .A2(new_n333_), .B(new_n118_), .ZN(new_n397_));
  XOR2_X1    g00333(.A1(new_n330_), .A2(new_n80_), .Z(new_n398_));
  NOR2_X1    g00334(.A1(new_n398_), .A2(new_n71_), .ZN(new_n399_));
  NOR2_X1    g00335(.A1(new_n297_), .A2(new_n89_), .ZN(new_n400_));
  NOR2_X1    g00336(.A1(new_n296_), .A2(new_n103_), .ZN(new_n401_));
  OAI21_X1   g00337(.A1(new_n400_), .A2(new_n401_), .B(new_n102_), .ZN(new_n402_));
  OAI21_X1   g00338(.A1(new_n298_), .A2(new_n300_), .B(new_n80_), .ZN(new_n403_));
  NAND2_X1   g00339(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1     g00340(.I(new_n404_), .ZN(new_n405_));
  NOR2_X1    g00341(.A1(new_n102_), .A2(\a[11] ), .ZN(new_n406_));
  INV_X1     g00342(.I(new_n406_), .ZN(new_n407_));
  NOR2_X1    g00343(.A1(new_n80_), .A2(new_n294_), .ZN(new_n408_));
  AOI21_X1   g00344(.A1(new_n207_), .A2(new_n407_), .B(new_n408_), .ZN(new_n409_));
  INV_X1     g00345(.I(new_n409_), .ZN(new_n410_));
  NOR2_X1    g00346(.A1(new_n405_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1     g00347(.I(new_n411_), .ZN(new_n412_));
  NOR2_X1    g00348(.A1(new_n404_), .A2(new_n409_), .ZN(new_n413_));
  AOI21_X1   g00349(.A1(new_n412_), .A2(new_n118_), .B(new_n413_), .ZN(new_n414_));
  INV_X1     g00350(.I(new_n414_), .ZN(new_n415_));
  NOR3_X1    g00351(.A1(new_n399_), .A2(new_n397_), .A3(new_n415_), .ZN(new_n416_));
  NOR2_X1    g00352(.A1(new_n399_), .A2(new_n397_), .ZN(new_n417_));
  NOR2_X1    g00353(.A1(new_n417_), .A2(new_n414_), .ZN(new_n418_));
  INV_X1     g00354(.I(new_n418_), .ZN(new_n419_));
  OAI21_X1   g00355(.A1(new_n189_), .A2(new_n416_), .B(new_n419_), .ZN(new_n420_));
  NOR2_X1    g00356(.A1(new_n396_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1     g00357(.I(new_n421_), .ZN(new_n422_));
  NAND2_X1   g00358(.A1(new_n396_), .A2(new_n420_), .ZN(new_n423_));
  INV_X1     g00359(.I(new_n423_), .ZN(new_n424_));
  AOI21_X1   g00360(.A1(new_n248_), .A2(new_n422_), .B(new_n424_), .ZN(new_n425_));
  INV_X1     g00361(.I(new_n425_), .ZN(new_n426_));
  NOR2_X1    g00362(.A1(new_n392_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1    g00363(.A1(new_n427_), .A2(new_n356_), .ZN(new_n428_));
  NOR2_X1    g00364(.A1(new_n391_), .A2(new_n425_), .ZN(new_n429_));
  NOR2_X1    g00365(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NOR2_X1    g00366(.A1(new_n387_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1   g00367(.A1(new_n387_), .A2(new_n430_), .B(new_n126_), .ZN(new_n432_));
  NOR2_X1    g00368(.A1(new_n432_), .A2(new_n431_), .ZN(new_n433_));
  XOR2_X1    g00369(.A1(new_n379_), .A2(new_n273_), .Z(new_n434_));
  INV_X1     g00370(.I(new_n381_), .ZN(new_n435_));
  OAI21_X1   g00371(.A1(new_n435_), .A2(new_n380_), .B(new_n352_), .ZN(new_n436_));
  OAI21_X1   g00372(.A1(new_n352_), .A2(new_n434_), .B(new_n436_), .ZN(new_n437_));
  NAND2_X1   g00373(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1     g00374(.I(\a[16] ), .ZN(new_n439_));
  NOR2_X1    g00375(.A1(new_n439_), .A2(\a[14] ), .ZN(new_n440_));
  NOR2_X1    g00376(.A1(new_n279_), .A2(\a[16] ), .ZN(new_n441_));
  NOR2_X1    g00377(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NOR3_X1    g00378(.A1(new_n442_), .A2(\a[15] ), .A3(new_n126_), .ZN(new_n443_));
  NOR2_X1    g00379(.A1(new_n418_), .A2(new_n416_), .ZN(new_n444_));
  NOR2_X1    g00380(.A1(new_n444_), .A2(new_n189_), .ZN(new_n445_));
  XOR2_X1    g00381(.A1(new_n417_), .A2(new_n415_), .Z(new_n446_));
  NOR2_X1    g00382(.A1(new_n446_), .A2(new_n248_), .ZN(new_n447_));
  OAI21_X1   g00383(.A1(new_n411_), .A2(new_n413_), .B(new_n118_), .ZN(new_n448_));
  XOR2_X1    g00384(.A1(new_n404_), .A2(new_n410_), .Z(new_n449_));
  OAI21_X1   g00385(.A1(new_n118_), .A2(new_n449_), .B(new_n448_), .ZN(new_n450_));
  INV_X1     g00386(.I(\a[2] ), .ZN(new_n451_));
  INV_X1     g00387(.I(\a[5] ), .ZN(new_n452_));
  NOR2_X1    g00388(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1   g00389(.A1(\a[8] ), .A2(new_n453_), .B(new_n93_), .ZN(new_n454_));
  AOI21_X1   g00390(.A1(new_n454_), .A2(new_n93_), .B(new_n80_), .ZN(new_n455_));
  NOR2_X1    g00391(.A1(new_n454_), .A2(new_n93_), .ZN(new_n456_));
  NOR2_X1    g00392(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1     g00393(.I(new_n457_), .ZN(new_n458_));
  NOR2_X1    g00394(.A1(new_n278_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1     g00395(.I(new_n459_), .ZN(new_n460_));
  NOR2_X1    g00396(.A1(new_n287_), .A2(new_n457_), .ZN(new_n461_));
  AOI21_X1   g00397(.A1(new_n118_), .A2(new_n460_), .B(new_n461_), .ZN(new_n462_));
  INV_X1     g00398(.I(new_n462_), .ZN(new_n463_));
  OAI21_X1   g00399(.A1(new_n406_), .A2(new_n408_), .B(new_n207_), .ZN(new_n464_));
  XOR2_X1    g00400(.A1(new_n102_), .A2(new_n294_), .Z(new_n465_));
  OAI21_X1   g00401(.A1(new_n207_), .A2(new_n465_), .B(new_n464_), .ZN(new_n466_));
  NOR2_X1    g00402(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1     g00403(.I(new_n467_), .ZN(new_n468_));
  INV_X1     g00404(.I(new_n466_), .ZN(new_n469_));
  NOR2_X1    g00405(.A1(new_n469_), .A2(new_n462_), .ZN(new_n470_));
  AOI21_X1   g00406(.A1(new_n468_), .A2(new_n118_), .B(new_n470_), .ZN(new_n471_));
  INV_X1     g00407(.I(new_n471_), .ZN(new_n472_));
  NOR2_X1    g00408(.A1(new_n472_), .A2(new_n189_), .ZN(new_n473_));
  INV_X1     g00409(.I(new_n473_), .ZN(new_n474_));
  NOR2_X1    g00410(.A1(new_n471_), .A2(new_n248_), .ZN(new_n475_));
  AOI21_X1   g00411(.A1(new_n474_), .A2(new_n450_), .B(new_n475_), .ZN(new_n476_));
  INV_X1     g00412(.I(new_n476_), .ZN(new_n477_));
  NOR3_X1    g00413(.A1(new_n447_), .A2(new_n445_), .A3(new_n477_), .ZN(new_n478_));
  NOR2_X1    g00414(.A1(new_n447_), .A2(new_n445_), .ZN(new_n479_));
  NOR2_X1    g00415(.A1(new_n479_), .A2(new_n476_), .ZN(new_n480_));
  OAI21_X1   g00416(.A1(new_n480_), .A2(new_n478_), .B(new_n356_), .ZN(new_n481_));
  XOR2_X1    g00417(.A1(new_n479_), .A2(new_n477_), .Z(new_n482_));
  OAI21_X1   g00418(.A1(new_n482_), .A2(new_n356_), .B(new_n481_), .ZN(new_n483_));
  OAI21_X1   g00419(.A1(new_n473_), .A2(new_n475_), .B(new_n450_), .ZN(new_n484_));
  INV_X1     g00420(.I(new_n450_), .ZN(new_n485_));
  XOR2_X1    g00421(.A1(new_n471_), .A2(new_n248_), .Z(new_n486_));
  NAND2_X1   g00422(.A1(new_n486_), .A2(new_n485_), .ZN(new_n487_));
  AND2_X2    g00423(.A1(new_n487_), .A2(new_n484_), .Z(new_n488_));
  INV_X1     g00424(.I(new_n488_), .ZN(new_n489_));
  XOR2_X1    g00425(.A1(new_n462_), .A2(new_n466_), .Z(new_n490_));
  OAI21_X1   g00426(.A1(new_n467_), .A2(new_n470_), .B(new_n71_), .ZN(new_n491_));
  OAI21_X1   g00427(.A1(new_n490_), .A2(new_n71_), .B(new_n491_), .ZN(new_n492_));
  OAI21_X1   g00428(.A1(new_n461_), .A2(new_n459_), .B(new_n118_), .ZN(new_n493_));
  XOR2_X1    g00429(.A1(new_n278_), .A2(new_n458_), .Z(new_n494_));
  NAND2_X1   g00430(.A1(new_n494_), .A2(new_n71_), .ZN(new_n495_));
  AND2_X2    g00431(.A1(new_n495_), .A2(new_n493_), .Z(new_n496_));
  INV_X1     g00432(.I(new_n496_), .ZN(new_n497_));
  INV_X1     g00433(.I(\a[8] ), .ZN(new_n498_));
  INV_X1     g00434(.I(new_n453_), .ZN(new_n499_));
  NOR3_X1    g00435(.A1(new_n93_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NOR2_X1    g00436(.A1(new_n500_), .A2(new_n80_), .ZN(new_n501_));
  NOR4_X1    g00437(.A1(new_n93_), .A2(new_n102_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n502_));
  NOR2_X1    g00438(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1     g00439(.I(new_n503_), .ZN(new_n504_));
  NAND2_X1   g00440(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n505_));
  INV_X1     g00441(.I(new_n505_), .ZN(new_n506_));
  NOR2_X1    g00442(.A1(new_n451_), .A2(new_n452_), .ZN(new_n507_));
  NOR2_X1    g00443(.A1(new_n80_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1    g00444(.A1(new_n451_), .A2(new_n452_), .ZN(new_n509_));
  NOR2_X1    g00445(.A1(new_n94_), .A2(\a[2] ), .ZN(new_n510_));
  NAND2_X1   g00446(.A1(new_n81_), .A2(new_n83_), .ZN(new_n511_));
  NOR2_X1    g00447(.A1(new_n82_), .A2(new_n511_), .ZN(new_n512_));
  NOR2_X1    g00448(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n513_));
  NOR2_X1    g00449(.A1(new_n453_), .A2(new_n513_), .ZN(new_n514_));
  OAI21_X1   g00450(.A1(new_n512_), .A2(new_n514_), .B(new_n510_), .ZN(new_n515_));
  NAND2_X1   g00451(.A1(new_n512_), .A2(new_n514_), .ZN(new_n516_));
  AOI21_X1   g00452(.A1(new_n515_), .A2(new_n516_), .B(new_n509_), .ZN(new_n517_));
  NOR2_X1    g00453(.A1(new_n517_), .A2(new_n508_), .ZN(new_n518_));
  NOR2_X1    g00454(.A1(new_n518_), .A2(new_n506_), .ZN(new_n519_));
  NOR2_X1    g00455(.A1(new_n93_), .A2(\a[8] ), .ZN(new_n520_));
  NOR2_X1    g00456(.A1(new_n94_), .A2(new_n498_), .ZN(new_n521_));
  OAI21_X1   g00457(.A1(new_n521_), .A2(new_n520_), .B(new_n506_), .ZN(new_n522_));
  NOR3_X1    g00458(.A1(new_n93_), .A2(new_n498_), .A3(new_n453_), .ZN(new_n523_));
  INV_X1     g00459(.I(new_n523_), .ZN(new_n524_));
  AND2_X2    g00460(.A1(new_n522_), .A2(new_n524_), .Z(new_n525_));
  INV_X1     g00461(.I(new_n525_), .ZN(new_n526_));
  NOR2_X1    g00462(.A1(new_n519_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1     g00463(.I(new_n527_), .ZN(new_n528_));
  NOR3_X1    g00464(.A1(new_n518_), .A2(new_n506_), .A3(new_n525_), .ZN(new_n529_));
  AOI21_X1   g00465(.A1(new_n528_), .A2(new_n102_), .B(new_n529_), .ZN(new_n530_));
  AND2_X2    g00466(.A1(new_n530_), .A2(new_n504_), .Z(new_n531_));
  NOR2_X1    g00467(.A1(new_n531_), .A2(new_n71_), .ZN(new_n532_));
  NOR2_X1    g00468(.A1(new_n530_), .A2(new_n504_), .ZN(new_n533_));
  NOR2_X1    g00469(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1     g00470(.I(new_n534_), .ZN(new_n535_));
  NOR2_X1    g00471(.A1(new_n535_), .A2(new_n497_), .ZN(new_n536_));
  INV_X1     g00472(.I(new_n536_), .ZN(new_n537_));
  NOR2_X1    g00473(.A1(new_n534_), .A2(new_n496_), .ZN(new_n538_));
  AOI21_X1   g00474(.A1(new_n537_), .A2(new_n189_), .B(new_n538_), .ZN(new_n539_));
  AND2_X2    g00475(.A1(new_n539_), .A2(new_n492_), .Z(new_n540_));
  NOR2_X1    g00476(.A1(new_n540_), .A2(new_n189_), .ZN(new_n541_));
  NOR2_X1    g00477(.A1(new_n539_), .A2(new_n492_), .ZN(new_n542_));
  NOR3_X1    g00478(.A1(new_n541_), .A2(new_n489_), .A3(new_n542_), .ZN(new_n543_));
  NOR2_X1    g00479(.A1(new_n541_), .A2(new_n542_), .ZN(new_n544_));
  NOR2_X1    g00480(.A1(new_n544_), .A2(new_n488_), .ZN(new_n545_));
  INV_X1     g00481(.I(new_n545_), .ZN(new_n546_));
  OAI21_X1   g00482(.A1(new_n356_), .A2(new_n543_), .B(new_n546_), .ZN(new_n547_));
  NOR2_X1    g00483(.A1(new_n547_), .A2(new_n483_), .ZN(new_n548_));
  NAND2_X1   g00484(.A1(new_n547_), .A2(new_n483_), .ZN(new_n549_));
  OAI21_X1   g00485(.A1(new_n443_), .A2(new_n548_), .B(new_n549_), .ZN(new_n550_));
  NOR2_X1    g00486(.A1(new_n478_), .A2(new_n273_), .ZN(new_n551_));
  NOR2_X1    g00487(.A1(new_n551_), .A2(new_n480_), .ZN(new_n552_));
  XOR2_X1    g00488(.A1(new_n420_), .A2(new_n395_), .Z(new_n553_));
  NOR2_X1    g00489(.A1(new_n553_), .A2(new_n189_), .ZN(new_n554_));
  AOI21_X1   g00490(.A1(new_n422_), .A2(new_n423_), .B(new_n248_), .ZN(new_n555_));
  NOR2_X1    g00491(.A1(new_n555_), .A2(new_n554_), .ZN(new_n556_));
  XNOR2_X1   g00492(.A1(new_n556_), .A2(new_n552_), .ZN(new_n557_));
  NAND2_X1   g00493(.A1(new_n557_), .A2(new_n273_), .ZN(new_n558_));
  INV_X1     g00494(.I(new_n556_), .ZN(new_n559_));
  NOR2_X1    g00495(.A1(new_n559_), .A2(new_n552_), .ZN(new_n560_));
  NAND2_X1   g00496(.A1(new_n559_), .A2(new_n552_), .ZN(new_n561_));
  INV_X1     g00497(.I(new_n561_), .ZN(new_n562_));
  OAI21_X1   g00498(.A1(new_n562_), .A2(new_n560_), .B(new_n356_), .ZN(new_n563_));
  NAND2_X1   g00499(.A1(new_n563_), .A2(new_n558_), .ZN(new_n564_));
  INV_X1     g00500(.I(new_n564_), .ZN(new_n565_));
  NOR2_X1    g00501(.A1(new_n565_), .A2(new_n443_), .ZN(new_n566_));
  INV_X1     g00502(.I(new_n566_), .ZN(new_n567_));
  INV_X1     g00503(.I(new_n443_), .ZN(new_n568_));
  NOR2_X1    g00504(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1   g00505(.A1(new_n567_), .A2(new_n550_), .B(new_n569_), .ZN(new_n570_));
  INV_X1     g00506(.I(new_n570_), .ZN(new_n571_));
  INV_X1     g00507(.I(new_n549_), .ZN(new_n572_));
  OAI21_X1   g00508(.A1(new_n572_), .A2(new_n548_), .B(new_n568_), .ZN(new_n573_));
  XNOR2_X1   g00509(.A1(new_n547_), .A2(new_n483_), .ZN(new_n574_));
  OAI21_X1   g00510(.A1(new_n568_), .A2(new_n574_), .B(new_n573_), .ZN(new_n575_));
  INV_X1     g00511(.I(new_n575_), .ZN(new_n576_));
  OAI21_X1   g00512(.A1(new_n545_), .A2(new_n543_), .B(new_n273_), .ZN(new_n577_));
  XOR2_X1    g00513(.A1(new_n544_), .A2(new_n489_), .Z(new_n578_));
  OAI21_X1   g00514(.A1(new_n578_), .A2(new_n273_), .B(new_n577_), .ZN(new_n579_));
  XOR2_X1    g00515(.A1(new_n539_), .A2(new_n492_), .Z(new_n580_));
  NAND2_X1   g00516(.A1(new_n580_), .A2(new_n248_), .ZN(new_n581_));
  OAI21_X1   g00517(.A1(new_n540_), .A2(new_n542_), .B(new_n189_), .ZN(new_n582_));
  NAND2_X1   g00518(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1     g00519(.I(new_n583_), .ZN(new_n584_));
  OAI21_X1   g00520(.A1(new_n536_), .A2(new_n538_), .B(new_n189_), .ZN(new_n585_));
  XOR2_X1    g00521(.A1(new_n534_), .A2(new_n497_), .Z(new_n586_));
  OAI21_X1   g00522(.A1(new_n189_), .A2(new_n586_), .B(new_n585_), .ZN(new_n587_));
  OAI21_X1   g00523(.A1(new_n531_), .A2(new_n533_), .B(new_n118_), .ZN(new_n588_));
  XOR2_X1    g00524(.A1(new_n530_), .A2(new_n503_), .Z(new_n589_));
  OAI21_X1   g00525(.A1(new_n118_), .A2(new_n589_), .B(new_n588_), .ZN(new_n590_));
  XOR2_X1    g00526(.A1(new_n519_), .A2(new_n525_), .Z(new_n591_));
  OAI21_X1   g00527(.A1(new_n527_), .A2(new_n529_), .B(new_n80_), .ZN(new_n592_));
  OAI21_X1   g00528(.A1(new_n591_), .A2(new_n80_), .B(new_n592_), .ZN(new_n593_));
  XOR2_X1    g00529(.A1(new_n518_), .A2(new_n505_), .Z(new_n594_));
  INV_X1     g00530(.I(new_n594_), .ZN(new_n595_));
  NOR2_X1    g00531(.A1(new_n595_), .A2(new_n102_), .ZN(new_n596_));
  INV_X1     g00532(.I(new_n596_), .ZN(new_n597_));
  NOR2_X1    g00533(.A1(new_n594_), .A2(new_n80_), .ZN(new_n598_));
  AOI21_X1   g00534(.A1(new_n597_), .A2(new_n71_), .B(new_n598_), .ZN(new_n599_));
  AND2_X2    g00535(.A1(new_n599_), .A2(new_n593_), .Z(new_n600_));
  NOR2_X1    g00536(.A1(new_n600_), .A2(new_n71_), .ZN(new_n601_));
  NOR2_X1    g00537(.A1(new_n599_), .A2(new_n593_), .ZN(new_n602_));
  NOR2_X1    g00538(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1     g00539(.I(new_n603_), .ZN(new_n604_));
  NOR2_X1    g00540(.A1(new_n604_), .A2(new_n590_), .ZN(new_n605_));
  INV_X1     g00541(.I(new_n605_), .ZN(new_n606_));
  NAND2_X1   g00542(.A1(new_n604_), .A2(new_n590_), .ZN(new_n607_));
  INV_X1     g00543(.I(new_n607_), .ZN(new_n608_));
  AOI21_X1   g00544(.A1(new_n248_), .A2(new_n606_), .B(new_n608_), .ZN(new_n609_));
  INV_X1     g00545(.I(new_n609_), .ZN(new_n610_));
  NOR2_X1    g00546(.A1(new_n610_), .A2(new_n587_), .ZN(new_n611_));
  INV_X1     g00547(.I(new_n611_), .ZN(new_n612_));
  INV_X1     g00548(.I(new_n587_), .ZN(new_n613_));
  NOR2_X1    g00549(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  AOI21_X1   g00550(.A1(new_n612_), .A2(new_n273_), .B(new_n614_), .ZN(new_n615_));
  INV_X1     g00551(.I(new_n615_), .ZN(new_n616_));
  NOR2_X1    g00552(.A1(new_n616_), .A2(new_n584_), .ZN(new_n617_));
  INV_X1     g00553(.I(new_n617_), .ZN(new_n618_));
  NOR2_X1    g00554(.A1(new_n615_), .A2(new_n583_), .ZN(new_n619_));
  AOI21_X1   g00555(.A1(new_n618_), .A2(new_n273_), .B(new_n619_), .ZN(new_n620_));
  INV_X1     g00556(.I(new_n620_), .ZN(new_n621_));
  NOR2_X1    g00557(.A1(new_n621_), .A2(new_n579_), .ZN(new_n622_));
  NOR2_X1    g00558(.A1(new_n622_), .A2(new_n443_), .ZN(new_n623_));
  INV_X1     g00559(.I(new_n579_), .ZN(new_n624_));
  NOR2_X1    g00560(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1    g00561(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1    g00562(.A1(new_n626_), .A2(new_n576_), .ZN(new_n627_));
  AOI21_X1   g00563(.A1(new_n626_), .A2(new_n576_), .B(new_n279_), .ZN(new_n628_));
  NOR2_X1    g00564(.A1(new_n628_), .A2(new_n627_), .ZN(new_n629_));
  INV_X1     g00565(.I(new_n629_), .ZN(new_n630_));
  INV_X1     g00566(.I(new_n550_), .ZN(new_n631_));
  XOR2_X1    g00567(.A1(new_n564_), .A2(new_n443_), .Z(new_n632_));
  OAI21_X1   g00568(.A1(new_n566_), .A2(new_n569_), .B(new_n631_), .ZN(new_n633_));
  OAI21_X1   g00569(.A1(new_n631_), .A2(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1     g00570(.I(new_n634_), .ZN(new_n635_));
  NOR2_X1    g00571(.A1(new_n630_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1   g00572(.A1(new_n636_), .A2(new_n571_), .ZN(new_n637_));
  XOR2_X1    g00573(.A1(\a[12] ), .A2(\a[14] ), .Z(new_n638_));
  NAND2_X1   g00574(.A1(new_n294_), .A2(\a[13] ), .ZN(new_n639_));
  INV_X1     g00575(.I(\a[13] ), .ZN(new_n640_));
  NAND2_X1   g00576(.A1(new_n640_), .A2(\a[11] ), .ZN(new_n641_));
  NAND2_X1   g00577(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1   g00578(.A1(new_n642_), .A2(new_n638_), .ZN(new_n643_));
  NOR2_X1    g00579(.A1(new_n643_), .A2(new_n279_), .ZN(new_n644_));
  OAI21_X1   g00580(.A1(new_n611_), .A2(new_n614_), .B(new_n273_), .ZN(new_n645_));
  XOR2_X1    g00581(.A1(new_n609_), .A2(new_n587_), .Z(new_n646_));
  OAI21_X1   g00582(.A1(new_n273_), .A2(new_n646_), .B(new_n645_), .ZN(new_n647_));
  AOI21_X1   g00583(.A1(new_n606_), .A2(new_n607_), .B(new_n189_), .ZN(new_n648_));
  XOR2_X1    g00584(.A1(new_n603_), .A2(new_n590_), .Z(new_n649_));
  NOR2_X1    g00585(.A1(new_n649_), .A2(new_n248_), .ZN(new_n650_));
  NOR2_X1    g00586(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  XOR2_X1    g00587(.A1(new_n599_), .A2(new_n593_), .Z(new_n652_));
  NAND2_X1   g00588(.A1(new_n652_), .A2(new_n118_), .ZN(new_n653_));
  OAI21_X1   g00589(.A1(new_n600_), .A2(new_n602_), .B(new_n71_), .ZN(new_n654_));
  NAND2_X1   g00590(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI21_X1   g00591(.A1(new_n596_), .A2(new_n598_), .B(new_n71_), .ZN(new_n656_));
  XOR2_X1    g00592(.A1(new_n594_), .A2(new_n102_), .Z(new_n657_));
  OAI21_X1   g00593(.A1(new_n71_), .A2(new_n657_), .B(new_n656_), .ZN(new_n658_));
  NOR2_X1    g00594(.A1(new_n451_), .A2(new_n452_), .ZN(new_n659_));
  OAI21_X1   g00595(.A1(new_n517_), .A2(new_n507_), .B(new_n80_), .ZN(new_n660_));
  OAI21_X1   g00596(.A1(new_n80_), .A2(new_n659_), .B(new_n660_), .ZN(new_n661_));
  INV_X1     g00597(.I(new_n661_), .ZN(new_n662_));
  XOR2_X1    g00598(.A1(new_n93_), .A2(\a[2] ), .Z(new_n663_));
  NOR2_X1    g00599(.A1(new_n663_), .A2(new_n80_), .ZN(new_n664_));
  NAND2_X1   g00600(.A1(new_n94_), .A2(new_n451_), .ZN(new_n665_));
  INV_X1     g00601(.I(new_n665_), .ZN(new_n666_));
  NOR2_X1    g00602(.A1(new_n666_), .A2(new_n89_), .ZN(new_n667_));
  INV_X1     g00603(.I(new_n667_), .ZN(new_n668_));
  NOR2_X1    g00604(.A1(new_n665_), .A2(new_n103_), .ZN(new_n669_));
  AOI21_X1   g00605(.A1(new_n668_), .A2(new_n664_), .B(new_n669_), .ZN(new_n670_));
  INV_X1     g00606(.I(new_n670_), .ZN(new_n671_));
  NAND2_X1   g00607(.A1(new_n94_), .A2(new_n451_), .ZN(new_n672_));
  NAND2_X1   g00608(.A1(new_n672_), .A2(new_n103_), .ZN(new_n673_));
  NOR2_X1    g00609(.A1(new_n672_), .A2(new_n103_), .ZN(new_n674_));
  AOI21_X1   g00610(.A1(new_n671_), .A2(new_n673_), .B(new_n674_), .ZN(new_n675_));
  XNOR2_X1   g00611(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n676_));
  INV_X1     g00612(.I(new_n676_), .ZN(new_n677_));
  NOR2_X1    g00613(.A1(new_n102_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1    g00614(.A1(new_n80_), .A2(new_n676_), .ZN(new_n679_));
  INV_X1     g00615(.I(new_n679_), .ZN(new_n680_));
  OAI21_X1   g00616(.A1(new_n675_), .A2(new_n678_), .B(new_n680_), .ZN(new_n681_));
  NOR2_X1    g00617(.A1(new_n681_), .A2(new_n662_), .ZN(new_n682_));
  INV_X1     g00618(.I(new_n682_), .ZN(new_n683_));
  NAND2_X1   g00619(.A1(new_n681_), .A2(new_n662_), .ZN(new_n684_));
  INV_X1     g00620(.I(new_n684_), .ZN(new_n685_));
  AOI21_X1   g00621(.A1(new_n118_), .A2(new_n683_), .B(new_n685_), .ZN(new_n686_));
  INV_X1     g00622(.I(new_n686_), .ZN(new_n687_));
  NOR2_X1    g00623(.A1(new_n687_), .A2(new_n658_), .ZN(new_n688_));
  INV_X1     g00624(.I(new_n688_), .ZN(new_n689_));
  INV_X1     g00625(.I(new_n658_), .ZN(new_n690_));
  NOR2_X1    g00626(.A1(new_n690_), .A2(new_n686_), .ZN(new_n691_));
  AOI21_X1   g00627(.A1(new_n689_), .A2(new_n248_), .B(new_n691_), .ZN(new_n692_));
  AND2_X2    g00628(.A1(new_n655_), .A2(new_n692_), .Z(new_n693_));
  NOR2_X1    g00629(.A1(new_n693_), .A2(new_n189_), .ZN(new_n694_));
  NOR2_X1    g00630(.A1(new_n655_), .A2(new_n692_), .ZN(new_n695_));
  NOR3_X1    g00631(.A1(new_n694_), .A2(new_n356_), .A3(new_n695_), .ZN(new_n696_));
  NOR2_X1    g00632(.A1(new_n651_), .A2(new_n696_), .ZN(new_n697_));
  NOR2_X1    g00633(.A1(new_n694_), .A2(new_n695_), .ZN(new_n698_));
  NOR2_X1    g00634(.A1(new_n698_), .A2(new_n273_), .ZN(new_n699_));
  NOR2_X1    g00635(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1     g00636(.I(new_n700_), .ZN(new_n701_));
  NOR2_X1    g00637(.A1(new_n647_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1     g00638(.I(new_n702_), .ZN(new_n703_));
  NAND2_X1   g00639(.A1(new_n647_), .A2(new_n701_), .ZN(new_n704_));
  AOI21_X1   g00640(.A1(new_n703_), .A2(new_n704_), .B(new_n568_), .ZN(new_n705_));
  XOR2_X1    g00641(.A1(new_n647_), .A2(new_n700_), .Z(new_n706_));
  NOR2_X1    g00642(.A1(new_n706_), .A2(new_n443_), .ZN(new_n707_));
  NOR2_X1    g00643(.A1(new_n707_), .A2(new_n705_), .ZN(new_n708_));
  INV_X1     g00644(.I(new_n708_), .ZN(new_n709_));
  NOR2_X1    g00645(.A1(new_n699_), .A2(new_n696_), .ZN(new_n710_));
  XOR2_X1    g00646(.A1(new_n698_), .A2(new_n273_), .Z(new_n711_));
  NAND2_X1   g00647(.A1(new_n711_), .A2(new_n651_), .ZN(new_n712_));
  OAI21_X1   g00648(.A1(new_n651_), .A2(new_n710_), .B(new_n712_), .ZN(new_n713_));
  XOR2_X1    g00649(.A1(new_n655_), .A2(new_n692_), .Z(new_n714_));
  NAND2_X1   g00650(.A1(new_n714_), .A2(new_n248_), .ZN(new_n715_));
  OAI21_X1   g00651(.A1(new_n693_), .A2(new_n695_), .B(new_n189_), .ZN(new_n716_));
  NAND2_X1   g00652(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1     g00653(.I(new_n717_), .ZN(new_n718_));
  OAI21_X1   g00654(.A1(new_n691_), .A2(new_n688_), .B(new_n248_), .ZN(new_n719_));
  XOR2_X1    g00655(.A1(new_n658_), .A2(new_n686_), .Z(new_n720_));
  OAI21_X1   g00656(.A1(new_n248_), .A2(new_n720_), .B(new_n719_), .ZN(new_n721_));
  AOI21_X1   g00657(.A1(new_n683_), .A2(new_n684_), .B(new_n71_), .ZN(new_n722_));
  XOR2_X1    g00658(.A1(new_n681_), .A2(new_n661_), .Z(new_n723_));
  NOR2_X1    g00659(.A1(new_n723_), .A2(new_n118_), .ZN(new_n724_));
  NAND3_X1   g00660(.A1(new_n89_), .A2(new_n94_), .A3(new_n451_), .ZN(new_n725_));
  XOR2_X1    g00661(.A1(new_n672_), .A2(new_n89_), .Z(new_n726_));
  OAI21_X1   g00662(.A1(new_n671_), .A2(new_n726_), .B(new_n725_), .ZN(new_n727_));
  NOR2_X1    g00663(.A1(new_n727_), .A2(new_n80_), .ZN(new_n728_));
  INV_X1     g00664(.I(new_n728_), .ZN(new_n729_));
  NAND2_X1   g00665(.A1(new_n727_), .A2(new_n80_), .ZN(new_n730_));
  INV_X1     g00666(.I(new_n730_), .ZN(new_n731_));
  AOI21_X1   g00667(.A1(new_n118_), .A2(new_n729_), .B(new_n731_), .ZN(new_n732_));
  NOR2_X1    g00668(.A1(new_n679_), .A2(new_n678_), .ZN(new_n733_));
  NOR2_X1    g00669(.A1(new_n675_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1     g00670(.I(new_n675_), .ZN(new_n735_));
  XOR2_X1    g00671(.A1(new_n102_), .A2(new_n676_), .Z(new_n736_));
  NOR2_X1    g00672(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NOR2_X1    g00673(.A1(new_n737_), .A2(new_n734_), .ZN(new_n738_));
  AND2_X2    g00674(.A1(new_n732_), .A2(new_n738_), .Z(new_n739_));
  NOR2_X1    g00675(.A1(new_n739_), .A2(new_n71_), .ZN(new_n740_));
  NOR2_X1    g00676(.A1(new_n732_), .A2(new_n738_), .ZN(new_n741_));
  NOR4_X1    g00677(.A1(new_n740_), .A2(new_n722_), .A3(new_n724_), .A4(new_n741_), .ZN(new_n742_));
  NOR2_X1    g00678(.A1(new_n742_), .A2(new_n189_), .ZN(new_n743_));
  NOR2_X1    g00679(.A1(new_n724_), .A2(new_n722_), .ZN(new_n744_));
  NOR2_X1    g00680(.A1(new_n740_), .A2(new_n741_), .ZN(new_n745_));
  NOR2_X1    g00681(.A1(new_n745_), .A2(new_n744_), .ZN(new_n746_));
  NOR2_X1    g00682(.A1(new_n743_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1     g00683(.I(new_n747_), .ZN(new_n748_));
  NOR2_X1    g00684(.A1(new_n748_), .A2(new_n721_), .ZN(new_n749_));
  INV_X1     g00685(.I(new_n749_), .ZN(new_n750_));
  INV_X1     g00686(.I(new_n721_), .ZN(new_n751_));
  NOR2_X1    g00687(.A1(new_n751_), .A2(new_n747_), .ZN(new_n752_));
  AOI21_X1   g00688(.A1(new_n750_), .A2(new_n356_), .B(new_n752_), .ZN(new_n753_));
  INV_X1     g00689(.I(new_n753_), .ZN(new_n754_));
  NOR2_X1    g00690(.A1(new_n754_), .A2(new_n718_), .ZN(new_n755_));
  INV_X1     g00691(.I(new_n755_), .ZN(new_n756_));
  NOR2_X1    g00692(.A1(new_n753_), .A2(new_n717_), .ZN(new_n757_));
  AOI21_X1   g00693(.A1(new_n756_), .A2(new_n273_), .B(new_n757_), .ZN(new_n758_));
  INV_X1     g00694(.I(new_n758_), .ZN(new_n759_));
  NOR2_X1    g00695(.A1(new_n759_), .A2(new_n713_), .ZN(new_n760_));
  NAND2_X1   g00696(.A1(new_n759_), .A2(new_n713_), .ZN(new_n761_));
  OAI21_X1   g00697(.A1(new_n443_), .A2(new_n760_), .B(new_n761_), .ZN(new_n762_));
  NOR2_X1    g00698(.A1(new_n709_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1   g00699(.A1(new_n709_), .A2(new_n762_), .ZN(new_n764_));
  OAI21_X1   g00700(.A1(new_n644_), .A2(new_n763_), .B(new_n764_), .ZN(new_n765_));
  INV_X1     g00701(.I(new_n765_), .ZN(new_n766_));
  OAI21_X1   g00702(.A1(new_n568_), .A2(new_n702_), .B(new_n704_), .ZN(new_n767_));
  XOR2_X1    g00703(.A1(new_n615_), .A2(new_n584_), .Z(new_n768_));
  OAI21_X1   g00704(.A1(new_n617_), .A2(new_n619_), .B(new_n356_), .ZN(new_n769_));
  OAI21_X1   g00705(.A1(new_n356_), .A2(new_n768_), .B(new_n769_), .ZN(new_n770_));
  XOR2_X1    g00706(.A1(new_n770_), .A2(new_n767_), .Z(new_n771_));
  NOR2_X1    g00707(.A1(new_n771_), .A2(new_n443_), .ZN(new_n772_));
  INV_X1     g00708(.I(new_n767_), .ZN(new_n773_));
  NOR2_X1    g00709(.A1(new_n770_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1     g00710(.I(new_n774_), .ZN(new_n775_));
  NAND2_X1   g00711(.A1(new_n770_), .A2(new_n773_), .ZN(new_n776_));
  AOI21_X1   g00712(.A1(new_n775_), .A2(new_n776_), .B(new_n568_), .ZN(new_n777_));
  NOR2_X1    g00713(.A1(new_n772_), .A2(new_n777_), .ZN(new_n778_));
  NOR2_X1    g00714(.A1(new_n778_), .A2(new_n644_), .ZN(new_n779_));
  NOR2_X1    g00715(.A1(new_n779_), .A2(new_n766_), .ZN(new_n780_));
  XNOR2_X1   g00716(.A1(\a[12] ), .A2(\a[14] ), .ZN(new_n781_));
  NOR2_X1    g00717(.A1(new_n640_), .A2(\a[11] ), .ZN(new_n782_));
  NOR2_X1    g00718(.A1(new_n294_), .A2(\a[13] ), .ZN(new_n783_));
  NOR2_X1    g00719(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1    g00720(.A1(new_n784_), .A2(new_n781_), .ZN(new_n785_));
  NAND2_X1   g00721(.A1(new_n785_), .A2(\a[14] ), .ZN(new_n786_));
  NOR3_X1    g00722(.A1(new_n772_), .A2(new_n786_), .A3(new_n777_), .ZN(new_n787_));
  OAI21_X1   g00723(.A1(new_n622_), .A2(new_n625_), .B(new_n568_), .ZN(new_n788_));
  XOR2_X1    g00724(.A1(new_n620_), .A2(new_n579_), .Z(new_n789_));
  OAI21_X1   g00725(.A1(new_n568_), .A2(new_n789_), .B(new_n788_), .ZN(new_n790_));
  NAND2_X1   g00726(.A1(new_n776_), .A2(new_n568_), .ZN(new_n791_));
  NAND2_X1   g00727(.A1(new_n791_), .A2(new_n775_), .ZN(new_n792_));
  XNOR2_X1   g00728(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  NOR2_X1    g00729(.A1(new_n793_), .A2(new_n786_), .ZN(new_n794_));
  NOR2_X1    g00730(.A1(new_n790_), .A2(new_n792_), .ZN(new_n795_));
  INV_X1     g00731(.I(new_n795_), .ZN(new_n796_));
  NAND2_X1   g00732(.A1(new_n790_), .A2(new_n792_), .ZN(new_n797_));
  AOI21_X1   g00733(.A1(new_n796_), .A2(new_n797_), .B(new_n644_), .ZN(new_n798_));
  OAI22_X1   g00734(.A1(new_n794_), .A2(new_n798_), .B1(new_n780_), .B2(new_n787_), .ZN(new_n799_));
  XNOR2_X1   g00735(.A1(\a[9] ), .A2(\a[11] ), .ZN(new_n800_));
  INV_X1     g00736(.I(\a[10] ), .ZN(new_n801_));
  NOR2_X1    g00737(.A1(new_n801_), .A2(\a[8] ), .ZN(new_n802_));
  NOR2_X1    g00738(.A1(new_n498_), .A2(\a[10] ), .ZN(new_n803_));
  NOR2_X1    g00739(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1    g00740(.A1(new_n804_), .A2(new_n800_), .ZN(new_n805_));
  NAND2_X1   g00741(.A1(new_n805_), .A2(\a[11] ), .ZN(new_n806_));
  OAI21_X1   g00742(.A1(new_n749_), .A2(new_n752_), .B(new_n356_), .ZN(new_n807_));
  XOR2_X1    g00743(.A1(new_n747_), .A2(new_n721_), .Z(new_n808_));
  OAI21_X1   g00744(.A1(new_n356_), .A2(new_n808_), .B(new_n807_), .ZN(new_n809_));
  OAI21_X1   g00745(.A1(new_n746_), .A2(new_n742_), .B(new_n248_), .ZN(new_n810_));
  XNOR2_X1   g00746(.A1(new_n745_), .A2(new_n744_), .ZN(new_n811_));
  OAI21_X1   g00747(.A1(new_n248_), .A2(new_n811_), .B(new_n810_), .ZN(new_n812_));
  XOR2_X1    g00748(.A1(new_n732_), .A2(new_n738_), .Z(new_n813_));
  NAND2_X1   g00749(.A1(new_n813_), .A2(new_n118_), .ZN(new_n814_));
  OAI21_X1   g00750(.A1(new_n739_), .A2(new_n741_), .B(new_n71_), .ZN(new_n815_));
  NAND2_X1   g00751(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1     g00752(.I(new_n816_), .ZN(new_n817_));
  AOI21_X1   g00753(.A1(new_n729_), .A2(new_n730_), .B(new_n71_), .ZN(new_n818_));
  XOR2_X1    g00754(.A1(new_n727_), .A2(new_n102_), .Z(new_n819_));
  NOR2_X1    g00755(.A1(new_n819_), .A2(new_n118_), .ZN(new_n820_));
  NOR2_X1    g00756(.A1(new_n820_), .A2(new_n818_), .ZN(new_n821_));
  INV_X1     g00757(.I(new_n821_), .ZN(new_n822_));
  OAI21_X1   g00758(.A1(new_n667_), .A2(new_n669_), .B(new_n664_), .ZN(new_n823_));
  INV_X1     g00759(.I(new_n823_), .ZN(new_n824_));
  XOR2_X1    g00760(.A1(new_n665_), .A2(new_n89_), .Z(new_n825_));
  NOR2_X1    g00761(.A1(new_n825_), .A2(new_n664_), .ZN(new_n826_));
  NOR2_X1    g00762(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1     g00763(.I(new_n827_), .ZN(new_n828_));
  NOR2_X1    g00764(.A1(new_n828_), .A2(new_n102_), .ZN(new_n829_));
  INV_X1     g00765(.I(new_n829_), .ZN(new_n830_));
  NOR2_X1    g00766(.A1(new_n827_), .A2(new_n80_), .ZN(new_n831_));
  AOI21_X1   g00767(.A1(new_n830_), .A2(new_n118_), .B(new_n831_), .ZN(new_n832_));
  INV_X1     g00768(.I(new_n832_), .ZN(new_n833_));
  NOR2_X1    g00769(.A1(new_n822_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1     g00770(.I(new_n834_), .ZN(new_n835_));
  NOR2_X1    g00771(.A1(new_n821_), .A2(new_n832_), .ZN(new_n836_));
  AOI21_X1   g00772(.A1(new_n835_), .A2(new_n189_), .B(new_n836_), .ZN(new_n837_));
  INV_X1     g00773(.I(new_n837_), .ZN(new_n838_));
  NOR2_X1    g00774(.A1(new_n838_), .A2(new_n817_), .ZN(new_n839_));
  INV_X1     g00775(.I(new_n839_), .ZN(new_n840_));
  NOR2_X1    g00776(.A1(new_n837_), .A2(new_n816_), .ZN(new_n841_));
  AOI21_X1   g00777(.A1(new_n840_), .A2(new_n248_), .B(new_n841_), .ZN(new_n842_));
  INV_X1     g00778(.I(new_n842_), .ZN(new_n843_));
  NOR2_X1    g00779(.A1(new_n843_), .A2(new_n812_), .ZN(new_n844_));
  NAND2_X1   g00780(.A1(new_n843_), .A2(new_n812_), .ZN(new_n845_));
  OAI21_X1   g00781(.A1(new_n356_), .A2(new_n844_), .B(new_n845_), .ZN(new_n846_));
  NOR2_X1    g00782(.A1(new_n846_), .A2(new_n809_), .ZN(new_n847_));
  NAND2_X1   g00783(.A1(new_n846_), .A2(new_n809_), .ZN(new_n848_));
  INV_X1     g00784(.I(new_n848_), .ZN(new_n849_));
  OAI21_X1   g00785(.A1(new_n849_), .A2(new_n847_), .B(new_n568_), .ZN(new_n850_));
  XNOR2_X1   g00786(.A1(new_n846_), .A2(new_n809_), .ZN(new_n851_));
  OAI21_X1   g00787(.A1(new_n568_), .A2(new_n851_), .B(new_n850_), .ZN(new_n852_));
  XNOR2_X1   g00788(.A1(new_n837_), .A2(new_n816_), .ZN(new_n853_));
  OAI21_X1   g00789(.A1(new_n839_), .A2(new_n841_), .B(new_n189_), .ZN(new_n854_));
  OAI21_X1   g00790(.A1(new_n189_), .A2(new_n853_), .B(new_n854_), .ZN(new_n855_));
  INV_X1     g00791(.I(new_n855_), .ZN(new_n856_));
  OAI21_X1   g00792(.A1(new_n834_), .A2(new_n836_), .B(new_n189_), .ZN(new_n857_));
  XOR2_X1    g00793(.A1(new_n821_), .A2(new_n833_), .Z(new_n858_));
  OAI21_X1   g00794(.A1(new_n189_), .A2(new_n858_), .B(new_n857_), .ZN(new_n859_));
  OAI21_X1   g00795(.A1(new_n829_), .A2(new_n831_), .B(new_n118_), .ZN(new_n860_));
  XOR2_X1    g00796(.A1(new_n827_), .A2(new_n80_), .Z(new_n861_));
  NAND2_X1   g00797(.A1(new_n861_), .A2(new_n71_), .ZN(new_n862_));
  XOR2_X1    g00798(.A1(\a[26] ), .A2(\a[27] ), .Z(new_n863_));
  NOR3_X1    g00799(.A1(new_n79_), .A2(new_n72_), .A3(new_n863_), .ZN(new_n864_));
  NAND4_X1   g00800(.A1(new_n80_), .A2(\a[31] ), .A3(new_n81_), .A4(new_n85_), .ZN(new_n865_));
  AOI21_X1   g00801(.A1(new_n865_), .A2(new_n94_), .B(new_n80_), .ZN(new_n866_));
  XOR2_X1    g00802(.A1(new_n663_), .A2(new_n80_), .Z(new_n867_));
  NOR2_X1    g00803(.A1(new_n867_), .A2(new_n118_), .ZN(new_n868_));
  INV_X1     g00804(.I(new_n868_), .ZN(new_n869_));
  NAND2_X1   g00805(.A1(new_n867_), .A2(new_n118_), .ZN(new_n870_));
  INV_X1     g00806(.I(new_n870_), .ZN(new_n871_));
  AOI21_X1   g00807(.A1(new_n866_), .A2(new_n869_), .B(new_n871_), .ZN(new_n872_));
  AOI21_X1   g00808(.A1(new_n862_), .A2(new_n860_), .B(new_n872_), .ZN(new_n873_));
  NAND2_X1   g00809(.A1(new_n862_), .A2(new_n860_), .ZN(new_n874_));
  INV_X1     g00810(.I(new_n872_), .ZN(new_n875_));
  NOR2_X1    g00811(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1    g00812(.A1(new_n876_), .A2(new_n68_), .ZN(new_n877_));
  NOR2_X1    g00813(.A1(new_n877_), .A2(new_n873_), .ZN(new_n878_));
  INV_X1     g00814(.I(new_n878_), .ZN(new_n879_));
  NOR2_X1    g00815(.A1(new_n859_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1     g00816(.I(new_n880_), .ZN(new_n881_));
  AND2_X2    g00817(.A1(new_n859_), .A2(new_n879_), .Z(new_n882_));
  AOI21_X1   g00818(.A1(new_n273_), .A2(new_n881_), .B(new_n882_), .ZN(new_n883_));
  INV_X1     g00819(.I(new_n883_), .ZN(new_n884_));
  NOR2_X1    g00820(.A1(new_n856_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1     g00821(.I(new_n885_), .ZN(new_n886_));
  NOR2_X1    g00822(.A1(new_n855_), .A2(new_n883_), .ZN(new_n887_));
  AOI21_X1   g00823(.A1(new_n886_), .A2(new_n273_), .B(new_n887_), .ZN(new_n888_));
  INV_X1     g00824(.I(new_n845_), .ZN(new_n889_));
  OAI21_X1   g00825(.A1(new_n889_), .A2(new_n844_), .B(new_n273_), .ZN(new_n890_));
  XOR2_X1    g00826(.A1(new_n842_), .A2(new_n812_), .Z(new_n891_));
  OAI21_X1   g00827(.A1(new_n273_), .A2(new_n891_), .B(new_n890_), .ZN(new_n892_));
  INV_X1     g00828(.I(new_n888_), .ZN(new_n893_));
  OAI21_X1   g00829(.A1(new_n443_), .A2(new_n893_), .B(new_n892_), .ZN(new_n894_));
  OAI21_X1   g00830(.A1(new_n568_), .A2(new_n888_), .B(new_n894_), .ZN(new_n895_));
  NOR2_X1    g00831(.A1(new_n895_), .A2(new_n852_), .ZN(new_n896_));
  NAND2_X1   g00832(.A1(new_n895_), .A2(new_n852_), .ZN(new_n897_));
  INV_X1     g00833(.I(new_n897_), .ZN(new_n898_));
  OAI21_X1   g00834(.A1(new_n898_), .A2(new_n896_), .B(new_n644_), .ZN(new_n899_));
  XNOR2_X1   g00835(.A1(new_n895_), .A2(new_n852_), .ZN(new_n900_));
  OAI21_X1   g00836(.A1(new_n644_), .A2(new_n900_), .B(new_n899_), .ZN(new_n901_));
  XOR2_X1    g00837(.A1(new_n888_), .A2(new_n568_), .Z(new_n902_));
  INV_X1     g00838(.I(new_n902_), .ZN(new_n903_));
  XOR2_X1    g00839(.A1(new_n888_), .A2(new_n443_), .Z(new_n904_));
  NOR2_X1    g00840(.A1(new_n904_), .A2(new_n892_), .ZN(new_n905_));
  AOI21_X1   g00841(.A1(new_n892_), .A2(new_n903_), .B(new_n905_), .ZN(new_n906_));
  INV_X1     g00842(.I(new_n906_), .ZN(new_n907_));
  XNOR2_X1   g00843(.A1(new_n855_), .A2(new_n883_), .ZN(new_n908_));
  OAI21_X1   g00844(.A1(new_n885_), .A2(new_n887_), .B(new_n356_), .ZN(new_n909_));
  OAI21_X1   g00845(.A1(new_n908_), .A2(new_n356_), .B(new_n909_), .ZN(new_n910_));
  INV_X1     g00846(.I(new_n910_), .ZN(new_n911_));
  OAI21_X1   g00847(.A1(new_n882_), .A2(new_n880_), .B(new_n273_), .ZN(new_n912_));
  XOR2_X1    g00848(.A1(new_n859_), .A2(new_n878_), .Z(new_n913_));
  OAI21_X1   g00849(.A1(new_n913_), .A2(new_n273_), .B(new_n912_), .ZN(new_n914_));
  XOR2_X1    g00850(.A1(new_n874_), .A2(new_n875_), .Z(new_n915_));
  XOR2_X1    g00851(.A1(new_n915_), .A2(new_n68_), .Z(new_n916_));
  INV_X1     g00852(.I(new_n916_), .ZN(new_n917_));
  XNOR2_X1   g00853(.A1(\a[26] ), .A2(\a[27] ), .ZN(new_n918_));
  NAND2_X1   g00854(.A1(new_n68_), .A2(\a[24] ), .ZN(new_n919_));
  NAND2_X1   g00855(.A1(new_n113_), .A2(\a[23] ), .ZN(new_n920_));
  NAND3_X1   g00856(.A1(new_n919_), .A2(new_n920_), .A3(\a[26] ), .ZN(new_n921_));
  AOI21_X1   g00857(.A1(new_n71_), .A2(new_n921_), .B(new_n918_), .ZN(new_n922_));
  NOR4_X1    g00858(.A1(new_n65_), .A2(new_n72_), .A3(\a[27] ), .A4(\a[28] ), .ZN(new_n923_));
  INV_X1     g00859(.I(new_n923_), .ZN(new_n924_));
  NAND3_X1   g00860(.A1(new_n79_), .A2(\a[29] ), .A3(new_n918_), .ZN(new_n925_));
  NAND2_X1   g00861(.A1(new_n925_), .A2(new_n924_), .ZN(new_n926_));
  AOI21_X1   g00862(.A1(new_n926_), .A2(new_n71_), .B(new_n922_), .ZN(new_n927_));
  NOR3_X1    g00863(.A1(new_n101_), .A2(new_n72_), .A3(new_n863_), .ZN(new_n928_));
  NOR3_X1    g00864(.A1(new_n928_), .A2(new_n71_), .A3(new_n923_), .ZN(new_n929_));
  NOR3_X1    g00865(.A1(new_n79_), .A2(new_n72_), .A3(new_n918_), .ZN(new_n930_));
  NAND2_X1   g00866(.A1(new_n930_), .A2(new_n118_), .ZN(new_n931_));
  OAI21_X1   g00867(.A1(new_n927_), .A2(new_n929_), .B(new_n931_), .ZN(new_n932_));
  NAND3_X1   g00868(.A1(new_n101_), .A2(\a[29] ), .A3(new_n863_), .ZN(new_n933_));
  NAND2_X1   g00869(.A1(new_n933_), .A2(new_n71_), .ZN(new_n934_));
  XNOR2_X1   g00870(.A1(\a[29] ), .A2(\a[30] ), .ZN(new_n935_));
  NAND4_X1   g00871(.A1(new_n101_), .A2(\a[29] ), .A3(new_n935_), .A4(new_n918_), .ZN(new_n936_));
  NOR4_X1    g00872(.A1(new_n76_), .A2(new_n72_), .A3(\a[26] ), .A4(\a[27] ), .ZN(new_n937_));
  INV_X1     g00873(.I(new_n937_), .ZN(new_n938_));
  XOR2_X1    g00874(.A1(\a[29] ), .A2(\a[30] ), .Z(new_n939_));
  AOI21_X1   g00875(.A1(new_n101_), .A2(\a[29] ), .B(new_n939_), .ZN(new_n940_));
  NOR2_X1    g00876(.A1(new_n77_), .A2(new_n78_), .ZN(new_n941_));
  NOR4_X1    g00877(.A1(new_n941_), .A2(new_n935_), .A3(\a[27] ), .A4(new_n72_), .ZN(new_n942_));
  OAI21_X1   g00878(.A1(new_n940_), .A2(new_n942_), .B(new_n938_), .ZN(new_n943_));
  AOI21_X1   g00879(.A1(new_n943_), .A2(new_n936_), .B(new_n118_), .ZN(new_n944_));
  AOI21_X1   g00880(.A1(new_n932_), .A2(new_n934_), .B(new_n944_), .ZN(new_n945_));
  INV_X1     g00881(.I(new_n936_), .ZN(new_n946_));
  OAI21_X1   g00882(.A1(new_n79_), .A2(new_n72_), .B(new_n935_), .ZN(new_n947_));
  NAND3_X1   g00883(.A1(new_n101_), .A2(\a[29] ), .A3(new_n939_), .ZN(new_n948_));
  AOI21_X1   g00884(.A1(new_n947_), .A2(new_n948_), .B(new_n937_), .ZN(new_n949_));
  NOR3_X1    g00885(.A1(new_n949_), .A2(new_n946_), .A3(new_n71_), .ZN(new_n950_));
  AOI21_X1   g00886(.A1(new_n864_), .A2(new_n939_), .B(new_n102_), .ZN(new_n951_));
  NOR2_X1    g00887(.A1(new_n80_), .A2(new_n935_), .ZN(new_n952_));
  NOR3_X1    g00888(.A1(new_n951_), .A2(new_n71_), .A3(new_n952_), .ZN(new_n953_));
  INV_X1     g00889(.I(new_n953_), .ZN(new_n954_));
  OAI21_X1   g00890(.A1(new_n945_), .A2(new_n950_), .B(new_n954_), .ZN(new_n955_));
  OAI21_X1   g00891(.A1(new_n935_), .A2(new_n938_), .B(new_n80_), .ZN(new_n956_));
  NAND2_X1   g00892(.A1(new_n102_), .A2(new_n939_), .ZN(new_n957_));
  AOI21_X1   g00893(.A1(new_n956_), .A2(new_n957_), .B(new_n118_), .ZN(new_n958_));
  INV_X1     g00894(.I(new_n958_), .ZN(new_n959_));
  XNOR2_X1   g00895(.A1(\a[29] ), .A2(\a[30] ), .ZN(new_n960_));
  NOR2_X1    g00896(.A1(new_n960_), .A2(new_n83_), .ZN(new_n961_));
  NOR2_X1    g00897(.A1(new_n960_), .A2(\a[31] ), .ZN(new_n962_));
  NOR3_X1    g00898(.A1(new_n80_), .A2(new_n961_), .A3(new_n962_), .ZN(new_n963_));
  INV_X1     g00899(.I(new_n963_), .ZN(new_n964_));
  NAND2_X1   g00900(.A1(new_n961_), .A2(new_n962_), .ZN(new_n965_));
  NOR2_X1    g00901(.A1(new_n965_), .A2(new_n80_), .ZN(new_n966_));
  NOR2_X1    g00902(.A1(new_n512_), .A2(new_n102_), .ZN(new_n967_));
  OAI22_X1   g00903(.A1(new_n966_), .A2(new_n967_), .B1(new_n80_), .B2(new_n939_), .ZN(new_n968_));
  AOI21_X1   g00904(.A1(new_n968_), .A2(new_n964_), .B(new_n118_), .ZN(new_n969_));
  AOI21_X1   g00905(.A1(new_n955_), .A2(new_n959_), .B(new_n969_), .ZN(new_n970_));
  NAND2_X1   g00906(.A1(new_n512_), .A2(new_n102_), .ZN(new_n971_));
  NAND2_X1   g00907(.A1(new_n965_), .A2(new_n80_), .ZN(new_n972_));
  AOI22_X1   g00908(.A1(new_n972_), .A2(new_n971_), .B1(new_n102_), .B2(new_n935_), .ZN(new_n973_));
  NOR3_X1    g00909(.A1(new_n973_), .A2(new_n71_), .A3(new_n963_), .ZN(new_n974_));
  NOR2_X1    g00910(.A1(new_n970_), .A2(new_n974_), .ZN(new_n975_));
  AOI21_X1   g00911(.A1(new_n965_), .A2(new_n939_), .B(new_n80_), .ZN(new_n976_));
  INV_X1     g00912(.I(new_n976_), .ZN(new_n977_));
  NOR2_X1    g00913(.A1(new_n977_), .A2(new_n118_), .ZN(new_n978_));
  NOR2_X1    g00914(.A1(new_n976_), .A2(new_n71_), .ZN(new_n979_));
  INV_X1     g00915(.I(new_n979_), .ZN(new_n980_));
  OAI21_X1   g00916(.A1(new_n975_), .A2(new_n978_), .B(new_n980_), .ZN(new_n981_));
  NOR4_X1    g00917(.A1(new_n80_), .A2(new_n88_), .A3(new_n82_), .A4(new_n511_), .ZN(new_n982_));
  OAI21_X1   g00918(.A1(new_n512_), .A2(new_n935_), .B(new_n102_), .ZN(new_n983_));
  INV_X1     g00919(.I(new_n983_), .ZN(new_n984_));
  NOR2_X1    g00920(.A1(new_n89_), .A2(new_n80_), .ZN(new_n985_));
  INV_X1     g00921(.I(new_n985_), .ZN(new_n986_));
  NAND2_X1   g00922(.A1(new_n89_), .A2(new_n80_), .ZN(new_n987_));
  AOI21_X1   g00923(.A1(new_n986_), .A2(new_n987_), .B(new_n984_), .ZN(new_n988_));
  NOR2_X1    g00924(.A1(new_n988_), .A2(new_n982_), .ZN(new_n989_));
  NOR2_X1    g00925(.A1(new_n989_), .A2(new_n118_), .ZN(new_n990_));
  INV_X1     g00926(.I(new_n990_), .ZN(new_n991_));
  INV_X1     g00927(.I(new_n989_), .ZN(new_n992_));
  NOR2_X1    g00928(.A1(new_n992_), .A2(new_n71_), .ZN(new_n993_));
  AOI21_X1   g00929(.A1(new_n981_), .A2(new_n991_), .B(new_n993_), .ZN(new_n994_));
  NOR2_X1    g00930(.A1(new_n865_), .A2(new_n80_), .ZN(new_n995_));
  NOR2_X1    g00931(.A1(new_n89_), .A2(new_n102_), .ZN(new_n996_));
  NOR2_X1    g00932(.A1(new_n995_), .A2(new_n996_), .ZN(new_n997_));
  NOR2_X1    g00933(.A1(new_n997_), .A2(new_n118_), .ZN(new_n998_));
  INV_X1     g00934(.I(new_n997_), .ZN(new_n999_));
  NOR2_X1    g00935(.A1(new_n999_), .A2(new_n71_), .ZN(new_n1000_));
  INV_X1     g00936(.I(new_n1000_), .ZN(new_n1001_));
  OAI21_X1   g00937(.A1(new_n994_), .A2(new_n998_), .B(new_n1001_), .ZN(new_n1002_));
  NAND2_X1   g00938(.A1(new_n1002_), .A2(new_n118_), .ZN(new_n1003_));
  XOR2_X1    g00939(.A1(new_n93_), .A2(new_n80_), .Z(new_n1004_));
  XOR2_X1    g00940(.A1(new_n1004_), .A2(new_n995_), .Z(new_n1005_));
  INV_X1     g00941(.I(new_n1005_), .ZN(new_n1006_));
  OAI21_X1   g00942(.A1(new_n1002_), .A2(new_n118_), .B(new_n1006_), .ZN(new_n1007_));
  NAND3_X1   g00943(.A1(new_n865_), .A2(new_n102_), .A3(new_n94_), .ZN(new_n1008_));
  AND2_X2    g00944(.A1(new_n1008_), .A2(new_n118_), .Z(new_n1009_));
  AOI21_X1   g00945(.A1(new_n1007_), .A2(new_n1003_), .B(new_n1009_), .ZN(new_n1010_));
  NOR2_X1    g00946(.A1(new_n1008_), .A2(new_n118_), .ZN(new_n1011_));
  NOR2_X1    g00947(.A1(new_n1010_), .A2(new_n1011_), .ZN(new_n1012_));
  INV_X1     g00948(.I(new_n866_), .ZN(new_n1013_));
  XOR2_X1    g00949(.A1(new_n867_), .A2(new_n71_), .Z(new_n1014_));
  NOR2_X1    g00950(.A1(new_n1014_), .A2(new_n1013_), .ZN(new_n1015_));
  AOI21_X1   g00951(.A1(new_n869_), .A2(new_n870_), .B(new_n866_), .ZN(new_n1016_));
  NOR2_X1    g00952(.A1(new_n1015_), .A2(new_n1016_), .ZN(new_n1017_));
  NOR2_X1    g00953(.A1(new_n1017_), .A2(new_n248_), .ZN(new_n1018_));
  INV_X1     g00954(.I(new_n1017_), .ZN(new_n1019_));
  NOR2_X1    g00955(.A1(new_n1019_), .A2(new_n189_), .ZN(new_n1020_));
  INV_X1     g00956(.I(new_n1020_), .ZN(new_n1021_));
  OAI21_X1   g00957(.A1(new_n1012_), .A2(new_n1018_), .B(new_n1021_), .ZN(new_n1022_));
  NOR2_X1    g00958(.A1(new_n917_), .A2(new_n1022_), .ZN(new_n1023_));
  INV_X1     g00959(.I(new_n1023_), .ZN(new_n1024_));
  NAND2_X1   g00960(.A1(new_n917_), .A2(new_n1022_), .ZN(new_n1025_));
  INV_X1     g00961(.I(new_n1025_), .ZN(new_n1026_));
  AOI21_X1   g00962(.A1(new_n273_), .A2(new_n1024_), .B(new_n1026_), .ZN(new_n1027_));
  INV_X1     g00963(.I(new_n1027_), .ZN(new_n1028_));
  NOR2_X1    g00964(.A1(new_n1028_), .A2(new_n914_), .ZN(new_n1029_));
  NOR2_X1    g00965(.A1(new_n1029_), .A2(new_n568_), .ZN(new_n1030_));
  INV_X1     g00966(.I(new_n914_), .ZN(new_n1031_));
  NOR2_X1    g00967(.A1(new_n1031_), .A2(new_n1027_), .ZN(new_n1032_));
  NOR2_X1    g00968(.A1(new_n1030_), .A2(new_n1032_), .ZN(new_n1033_));
  INV_X1     g00969(.I(new_n1033_), .ZN(new_n1034_));
  NOR2_X1    g00970(.A1(new_n911_), .A2(new_n1034_), .ZN(new_n1035_));
  INV_X1     g00971(.I(new_n1035_), .ZN(new_n1036_));
  NOR2_X1    g00972(.A1(new_n910_), .A2(new_n1033_), .ZN(new_n1037_));
  AOI21_X1   g00973(.A1(new_n1036_), .A2(new_n568_), .B(new_n1037_), .ZN(new_n1038_));
  INV_X1     g00974(.I(new_n1038_), .ZN(new_n1039_));
  NOR2_X1    g00975(.A1(new_n907_), .A2(new_n1039_), .ZN(new_n1040_));
  INV_X1     g00976(.I(new_n1040_), .ZN(new_n1041_));
  NOR2_X1    g00977(.A1(new_n906_), .A2(new_n1038_), .ZN(new_n1042_));
  AOI21_X1   g00978(.A1(new_n1041_), .A2(new_n786_), .B(new_n1042_), .ZN(new_n1043_));
  INV_X1     g00979(.I(new_n1043_), .ZN(new_n1044_));
  NOR2_X1    g00980(.A1(new_n1044_), .A2(new_n901_), .ZN(new_n1045_));
  INV_X1     g00981(.I(new_n1045_), .ZN(new_n1046_));
  NAND2_X1   g00982(.A1(new_n1044_), .A2(new_n901_), .ZN(new_n1047_));
  INV_X1     g00983(.I(new_n1047_), .ZN(new_n1048_));
  AOI21_X1   g00984(.A1(new_n806_), .A2(new_n1046_), .B(new_n1048_), .ZN(new_n1049_));
  OAI21_X1   g00985(.A1(new_n786_), .A2(new_n896_), .B(new_n897_), .ZN(new_n1050_));
  INV_X1     g00986(.I(new_n1050_), .ZN(new_n1051_));
  OAI21_X1   g00987(.A1(new_n443_), .A2(new_n847_), .B(new_n848_), .ZN(new_n1052_));
  XNOR2_X1   g00988(.A1(new_n753_), .A2(new_n717_), .ZN(new_n1053_));
  OAI21_X1   g00989(.A1(new_n755_), .A2(new_n757_), .B(new_n356_), .ZN(new_n1054_));
  OAI21_X1   g00990(.A1(new_n356_), .A2(new_n1053_), .B(new_n1054_), .ZN(new_n1055_));
  XOR2_X1    g00991(.A1(new_n1055_), .A2(new_n1052_), .Z(new_n1056_));
  NOR2_X1    g00992(.A1(new_n1056_), .A2(new_n443_), .ZN(new_n1057_));
  INV_X1     g00993(.I(new_n1052_), .ZN(new_n1058_));
  NOR2_X1    g00994(.A1(new_n1058_), .A2(new_n1055_), .ZN(new_n1059_));
  INV_X1     g00995(.I(new_n1059_), .ZN(new_n1060_));
  NAND2_X1   g00996(.A1(new_n1058_), .A2(new_n1055_), .ZN(new_n1061_));
  AOI21_X1   g00997(.A1(new_n1060_), .A2(new_n1061_), .B(new_n568_), .ZN(new_n1062_));
  NOR2_X1    g00998(.A1(new_n1062_), .A2(new_n1057_), .ZN(new_n1063_));
  INV_X1     g00999(.I(new_n1063_), .ZN(new_n1064_));
  NOR2_X1    g01000(.A1(new_n1051_), .A2(new_n1064_), .ZN(new_n1065_));
  NOR2_X1    g01001(.A1(new_n1050_), .A2(new_n1063_), .ZN(new_n1066_));
  NOR2_X1    g01002(.A1(new_n1065_), .A2(new_n1066_), .ZN(new_n1067_));
  NOR2_X1    g01003(.A1(new_n1067_), .A2(new_n644_), .ZN(new_n1068_));
  XNOR2_X1   g01004(.A1(new_n1050_), .A2(new_n1063_), .ZN(new_n1069_));
  NOR2_X1    g01005(.A1(new_n1069_), .A2(new_n786_), .ZN(new_n1070_));
  NOR2_X1    g01006(.A1(new_n1068_), .A2(new_n1070_), .ZN(new_n1071_));
  NOR2_X1    g01007(.A1(new_n1049_), .A2(new_n1071_), .ZN(new_n1072_));
  AOI21_X1   g01008(.A1(new_n1049_), .A2(new_n1071_), .B(\a[11] ), .ZN(new_n1073_));
  NOR2_X1    g01009(.A1(new_n1073_), .A2(new_n1072_), .ZN(new_n1074_));
  INV_X1     g01010(.I(\a[9] ), .ZN(new_n1075_));
  NOR2_X1    g01011(.A1(new_n1075_), .A2(\a[11] ), .ZN(new_n1076_));
  NOR2_X1    g01012(.A1(new_n294_), .A2(\a[9] ), .ZN(new_n1077_));
  OAI22_X1   g01013(.A1(new_n1076_), .A2(new_n1077_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n1078_));
  NOR2_X1    g01014(.A1(new_n1078_), .A2(new_n294_), .ZN(new_n1079_));
  INV_X1     g01015(.I(new_n760_), .ZN(new_n1080_));
  AOI21_X1   g01016(.A1(new_n1080_), .A2(new_n761_), .B(new_n443_), .ZN(new_n1081_));
  XOR2_X1    g01017(.A1(new_n713_), .A2(new_n758_), .Z(new_n1082_));
  NOR2_X1    g01018(.A1(new_n1082_), .A2(new_n568_), .ZN(new_n1083_));
  NAND2_X1   g01019(.A1(new_n1061_), .A2(new_n568_), .ZN(new_n1084_));
  NAND2_X1   g01020(.A1(new_n1084_), .A2(new_n1060_), .ZN(new_n1085_));
  NOR3_X1    g01021(.A1(new_n1085_), .A2(new_n1081_), .A3(new_n1083_), .ZN(new_n1086_));
  NOR2_X1    g01022(.A1(new_n1081_), .A2(new_n1083_), .ZN(new_n1087_));
  INV_X1     g01023(.I(new_n1085_), .ZN(new_n1088_));
  NOR2_X1    g01024(.A1(new_n1088_), .A2(new_n1087_), .ZN(new_n1089_));
  NOR2_X1    g01025(.A1(new_n1089_), .A2(new_n1086_), .ZN(new_n1090_));
  NOR2_X1    g01026(.A1(new_n1090_), .A2(new_n644_), .ZN(new_n1091_));
  XOR2_X1    g01027(.A1(new_n1087_), .A2(new_n1085_), .Z(new_n1092_));
  NOR2_X1    g01028(.A1(new_n1092_), .A2(new_n786_), .ZN(new_n1093_));
  NOR2_X1    g01029(.A1(new_n1093_), .A2(new_n1091_), .ZN(new_n1094_));
  INV_X1     g01030(.I(new_n1066_), .ZN(new_n1095_));
  AOI21_X1   g01031(.A1(new_n786_), .A2(new_n1095_), .B(new_n1065_), .ZN(new_n1096_));
  XOR2_X1    g01032(.A1(new_n1094_), .A2(new_n1096_), .Z(new_n1097_));
  INV_X1     g01033(.I(new_n1094_), .ZN(new_n1098_));
  INV_X1     g01034(.I(new_n1096_), .ZN(new_n1099_));
  NOR2_X1    g01035(.A1(new_n1098_), .A2(new_n1099_), .ZN(new_n1100_));
  NOR2_X1    g01036(.A1(new_n1094_), .A2(new_n1096_), .ZN(new_n1101_));
  NOR2_X1    g01037(.A1(new_n1100_), .A2(new_n1101_), .ZN(new_n1102_));
  NOR2_X1    g01038(.A1(new_n1102_), .A2(new_n1079_), .ZN(new_n1103_));
  AOI21_X1   g01039(.A1(new_n1097_), .A2(new_n1079_), .B(new_n1103_), .ZN(new_n1104_));
  NAND3_X1   g01040(.A1(new_n943_), .A2(new_n71_), .A3(new_n936_), .ZN(new_n1105_));
  OAI21_X1   g01041(.A1(new_n949_), .A2(new_n946_), .B(new_n118_), .ZN(new_n1106_));
  AOI22_X1   g01042(.A1(new_n932_), .A2(new_n934_), .B1(new_n1105_), .B2(new_n1106_), .ZN(new_n1107_));
  INV_X1     g01043(.I(new_n921_), .ZN(new_n1108_));
  OAI21_X1   g01044(.A1(new_n118_), .A2(new_n1108_), .B(new_n863_), .ZN(new_n1109_));
  OAI21_X1   g01045(.A1(new_n928_), .A2(new_n923_), .B(new_n71_), .ZN(new_n1110_));
  NAND2_X1   g01046(.A1(new_n1110_), .A2(new_n1109_), .ZN(new_n1111_));
  NAND3_X1   g01047(.A1(new_n925_), .A2(new_n118_), .A3(new_n924_), .ZN(new_n1112_));
  INV_X1     g01048(.I(new_n931_), .ZN(new_n1113_));
  AOI21_X1   g01049(.A1(new_n1111_), .A2(new_n1112_), .B(new_n1113_), .ZN(new_n1114_));
  INV_X1     g01050(.I(new_n934_), .ZN(new_n1115_));
  NOR2_X1    g01051(.A1(new_n950_), .A2(new_n944_), .ZN(new_n1116_));
  NOR3_X1    g01052(.A1(new_n1116_), .A2(new_n1114_), .A3(new_n1115_), .ZN(new_n1117_));
  NOR2_X1    g01053(.A1(new_n1117_), .A2(new_n1107_), .ZN(new_n1118_));
  NOR2_X1    g01054(.A1(new_n1118_), .A2(new_n248_), .ZN(new_n1119_));
  XNOR2_X1   g01055(.A1(\a[23] ), .A2(\a[24] ), .ZN(new_n1120_));
  XNOR2_X1   g01056(.A1(\a[20] ), .A2(\a[21] ), .ZN(new_n1121_));
  NAND2_X1   g01057(.A1(new_n1121_), .A2(\a[23] ), .ZN(new_n1122_));
  AOI21_X1   g01058(.A1(new_n189_), .A2(new_n1122_), .B(new_n1120_), .ZN(new_n1123_));
  NOR4_X1    g01059(.A1(new_n68_), .A2(new_n65_), .A3(\a[24] ), .A4(\a[25] ), .ZN(new_n1124_));
  INV_X1     g01060(.I(new_n1124_), .ZN(new_n1125_));
  NOR2_X1    g01061(.A1(new_n113_), .A2(\a[26] ), .ZN(new_n1126_));
  NOR2_X1    g01062(.A1(new_n65_), .A2(\a[24] ), .ZN(new_n1127_));
  OAI22_X1   g01063(.A1(new_n1126_), .A2(new_n1127_), .B1(new_n67_), .B2(new_n69_), .ZN(new_n1128_));
  NAND3_X1   g01064(.A1(new_n1128_), .A2(\a[26] ), .A3(new_n1120_), .ZN(new_n1129_));
  AOI21_X1   g01065(.A1(new_n1129_), .A2(new_n1125_), .B(new_n248_), .ZN(new_n1130_));
  NAND3_X1   g01066(.A1(new_n1129_), .A2(new_n248_), .A3(new_n1125_), .ZN(new_n1131_));
  OAI21_X1   g01067(.A1(new_n1130_), .A2(new_n1123_), .B(new_n1131_), .ZN(new_n1132_));
  NOR4_X1    g01068(.A1(new_n68_), .A2(new_n65_), .A3(\a[24] ), .A4(\a[25] ), .ZN(new_n1133_));
  INV_X1     g01069(.I(new_n1133_), .ZN(new_n1134_));
  NOR2_X1    g01070(.A1(new_n189_), .A2(new_n1134_), .ZN(new_n1135_));
  INV_X1     g01071(.I(new_n1135_), .ZN(new_n1136_));
  NOR2_X1    g01072(.A1(new_n248_), .A2(new_n1133_), .ZN(new_n1137_));
  AOI21_X1   g01073(.A1(new_n1132_), .A2(new_n1136_), .B(new_n1137_), .ZN(new_n1138_));
  NAND3_X1   g01074(.A1(new_n71_), .A2(new_n1108_), .A3(new_n863_), .ZN(new_n1139_));
  INV_X1     g01075(.I(new_n1139_), .ZN(new_n1140_));
  NAND3_X1   g01076(.A1(new_n117_), .A2(\a[26] ), .A3(\a[27] ), .ZN(new_n1141_));
  OAI21_X1   g01077(.A1(new_n1128_), .A2(new_n65_), .B(new_n863_), .ZN(new_n1142_));
  AOI22_X1   g01078(.A1(new_n1142_), .A2(new_n1141_), .B1(new_n71_), .B2(new_n1108_), .ZN(new_n1143_));
  NOR3_X1    g01079(.A1(new_n1143_), .A2(new_n1140_), .A3(new_n248_), .ZN(new_n1144_));
  OAI21_X1   g01080(.A1(new_n1143_), .A2(new_n1140_), .B(new_n248_), .ZN(new_n1145_));
  OAI21_X1   g01081(.A1(new_n1138_), .A2(new_n1144_), .B(new_n1145_), .ZN(new_n1146_));
  NAND3_X1   g01082(.A1(new_n925_), .A2(new_n71_), .A3(new_n924_), .ZN(new_n1147_));
  NAND2_X1   g01083(.A1(new_n926_), .A2(new_n118_), .ZN(new_n1148_));
  AOI21_X1   g01084(.A1(new_n1148_), .A2(new_n1147_), .B(new_n922_), .ZN(new_n1149_));
  AOI21_X1   g01085(.A1(new_n1110_), .A2(new_n1112_), .B(new_n1109_), .ZN(new_n1150_));
  OAI21_X1   g01086(.A1(new_n1149_), .A2(new_n1150_), .B(new_n248_), .ZN(new_n1151_));
  NOR3_X1    g01087(.A1(new_n928_), .A2(new_n118_), .A3(new_n923_), .ZN(new_n1152_));
  AOI21_X1   g01088(.A1(new_n925_), .A2(new_n924_), .B(new_n71_), .ZN(new_n1153_));
  OAI21_X1   g01089(.A1(new_n1152_), .A2(new_n1153_), .B(new_n1109_), .ZN(new_n1154_));
  AOI21_X1   g01090(.A1(new_n925_), .A2(new_n924_), .B(new_n118_), .ZN(new_n1155_));
  OAI21_X1   g01091(.A1(new_n1155_), .A2(new_n929_), .B(new_n922_), .ZN(new_n1156_));
  NAND3_X1   g01092(.A1(new_n1156_), .A2(new_n1154_), .A3(new_n189_), .ZN(new_n1157_));
  INV_X1     g01093(.I(new_n1157_), .ZN(new_n1158_));
  AOI21_X1   g01094(.A1(new_n1146_), .A2(new_n1151_), .B(new_n1158_), .ZN(new_n1159_));
  XOR2_X1    g01095(.A1(new_n933_), .A2(new_n71_), .Z(new_n1160_));
  OAI21_X1   g01096(.A1(new_n927_), .A2(new_n929_), .B(new_n1160_), .ZN(new_n1161_));
  NAND2_X1   g01097(.A1(new_n931_), .A2(new_n934_), .ZN(new_n1162_));
  NAND3_X1   g01098(.A1(new_n1111_), .A2(new_n1162_), .A3(new_n1112_), .ZN(new_n1163_));
  AOI21_X1   g01099(.A1(new_n1161_), .A2(new_n1163_), .B(new_n248_), .ZN(new_n1164_));
  NAND3_X1   g01100(.A1(new_n1161_), .A2(new_n248_), .A3(new_n1163_), .ZN(new_n1165_));
  OAI21_X1   g01101(.A1(new_n1159_), .A2(new_n1164_), .B(new_n1165_), .ZN(new_n1166_));
  NOR3_X1    g01102(.A1(new_n1117_), .A2(new_n1107_), .A3(new_n248_), .ZN(new_n1167_));
  INV_X1     g01103(.I(new_n1105_), .ZN(new_n1168_));
  AOI21_X1   g01104(.A1(new_n943_), .A2(new_n936_), .B(new_n71_), .ZN(new_n1169_));
  OAI22_X1   g01105(.A1(new_n1114_), .A2(new_n1115_), .B1(new_n1168_), .B2(new_n1169_), .ZN(new_n1170_));
  OAI21_X1   g01106(.A1(new_n949_), .A2(new_n946_), .B(new_n71_), .ZN(new_n1171_));
  NAND3_X1   g01107(.A1(new_n943_), .A2(new_n118_), .A3(new_n936_), .ZN(new_n1172_));
  NAND2_X1   g01108(.A1(new_n1171_), .A2(new_n1172_), .ZN(new_n1173_));
  NAND3_X1   g01109(.A1(new_n1173_), .A2(new_n932_), .A3(new_n934_), .ZN(new_n1174_));
  AOI21_X1   g01110(.A1(new_n1170_), .A2(new_n1174_), .B(new_n189_), .ZN(new_n1175_));
  NOR2_X1    g01111(.A1(new_n1167_), .A2(new_n1175_), .ZN(new_n1176_));
  OAI22_X1   g01112(.A1(new_n945_), .A2(new_n950_), .B1(new_n953_), .B2(new_n958_), .ZN(new_n1177_));
  OAI21_X1   g01113(.A1(new_n1114_), .A2(new_n1115_), .B(new_n1171_), .ZN(new_n1178_));
  AOI21_X1   g01114(.A1(new_n956_), .A2(new_n957_), .B(new_n71_), .ZN(new_n1179_));
  NOR3_X1    g01115(.A1(new_n951_), .A2(new_n118_), .A3(new_n952_), .ZN(new_n1180_));
  NOR2_X1    g01116(.A1(new_n1179_), .A2(new_n1180_), .ZN(new_n1181_));
  INV_X1     g01117(.I(new_n1181_), .ZN(new_n1182_));
  NAND3_X1   g01118(.A1(new_n1178_), .A2(new_n1182_), .A3(new_n1172_), .ZN(new_n1183_));
  AOI21_X1   g01119(.A1(new_n1177_), .A2(new_n1183_), .B(new_n189_), .ZN(new_n1184_));
  OAI21_X1   g01120(.A1(new_n1166_), .A2(new_n1176_), .B(new_n1184_), .ZN(new_n1185_));
  NAND2_X1   g01121(.A1(new_n919_), .A2(new_n920_), .ZN(new_n1186_));
  XOR2_X1    g01122(.A1(\a[20] ), .A2(\a[21] ), .Z(new_n1187_));
  NOR2_X1    g01123(.A1(new_n1187_), .A2(new_n68_), .ZN(new_n1188_));
  OAI21_X1   g01124(.A1(new_n248_), .A2(new_n1188_), .B(new_n1186_), .ZN(new_n1189_));
  AOI21_X1   g01125(.A1(new_n117_), .A2(\a[26] ), .B(new_n921_), .ZN(new_n1190_));
  OAI21_X1   g01126(.A1(new_n1190_), .A2(new_n1124_), .B(new_n189_), .ZN(new_n1191_));
  NOR3_X1    g01127(.A1(new_n1190_), .A2(new_n189_), .A3(new_n1124_), .ZN(new_n1192_));
  AOI21_X1   g01128(.A1(new_n1189_), .A2(new_n1191_), .B(new_n1192_), .ZN(new_n1193_));
  INV_X1     g01129(.I(new_n1137_), .ZN(new_n1194_));
  OAI21_X1   g01130(.A1(new_n1193_), .A2(new_n1135_), .B(new_n1194_), .ZN(new_n1195_));
  NOR3_X1    g01131(.A1(new_n1128_), .A2(new_n65_), .A3(new_n73_), .ZN(new_n1196_));
  AOI21_X1   g01132(.A1(new_n117_), .A2(\a[26] ), .B(new_n918_), .ZN(new_n1197_));
  OAI22_X1   g01133(.A1(new_n1196_), .A2(new_n1197_), .B1(new_n118_), .B2(new_n921_), .ZN(new_n1198_));
  NAND3_X1   g01134(.A1(new_n1198_), .A2(new_n189_), .A3(new_n1139_), .ZN(new_n1199_));
  INV_X1     g01135(.I(new_n1145_), .ZN(new_n1200_));
  AOI21_X1   g01136(.A1(new_n1195_), .A2(new_n1199_), .B(new_n1200_), .ZN(new_n1201_));
  AOI21_X1   g01137(.A1(new_n1156_), .A2(new_n1154_), .B(new_n189_), .ZN(new_n1202_));
  OAI21_X1   g01138(.A1(new_n1201_), .A2(new_n1202_), .B(new_n1157_), .ZN(new_n1203_));
  XOR2_X1    g01139(.A1(new_n933_), .A2(new_n118_), .Z(new_n1204_));
  AOI21_X1   g01140(.A1(new_n1111_), .A2(new_n1112_), .B(new_n1204_), .ZN(new_n1205_));
  INV_X1     g01141(.I(new_n1163_), .ZN(new_n1206_));
  OAI21_X1   g01142(.A1(new_n1206_), .A2(new_n1205_), .B(new_n189_), .ZN(new_n1207_));
  NOR3_X1    g01143(.A1(new_n1206_), .A2(new_n1205_), .A3(new_n189_), .ZN(new_n1208_));
  AOI21_X1   g01144(.A1(new_n1203_), .A2(new_n1207_), .B(new_n1208_), .ZN(new_n1209_));
  NAND3_X1   g01145(.A1(new_n1170_), .A2(new_n1174_), .A3(new_n189_), .ZN(new_n1210_));
  OAI21_X1   g01146(.A1(new_n1117_), .A2(new_n1107_), .B(new_n248_), .ZN(new_n1211_));
  NAND2_X1   g01147(.A1(new_n1211_), .A2(new_n1210_), .ZN(new_n1212_));
  AOI22_X1   g01148(.A1(new_n1178_), .A2(new_n1172_), .B1(new_n954_), .B2(new_n959_), .ZN(new_n1213_));
  NOR3_X1    g01149(.A1(new_n945_), .A2(new_n1181_), .A3(new_n950_), .ZN(new_n1214_));
  OAI21_X1   g01150(.A1(new_n1213_), .A2(new_n1214_), .B(new_n248_), .ZN(new_n1215_));
  NAND3_X1   g01151(.A1(new_n1209_), .A2(new_n1215_), .A3(new_n1212_), .ZN(new_n1216_));
  AOI21_X1   g01152(.A1(new_n1216_), .A2(new_n1185_), .B(new_n1119_), .ZN(new_n1217_));
  NOR2_X1    g01153(.A1(new_n1213_), .A2(new_n1214_), .ZN(new_n1218_));
  NOR2_X1    g01154(.A1(new_n1118_), .A2(new_n248_), .ZN(new_n1219_));
  NOR2_X1    g01155(.A1(new_n1217_), .A2(new_n1219_), .ZN(new_n1220_));
  NAND3_X1   g01156(.A1(new_n1156_), .A2(new_n1154_), .A3(new_n248_), .ZN(new_n1221_));
  OAI21_X1   g01157(.A1(new_n1149_), .A2(new_n1150_), .B(new_n189_), .ZN(new_n1222_));
  NAND2_X1   g01158(.A1(new_n1222_), .A2(new_n1221_), .ZN(new_n1223_));
  NAND2_X1   g01159(.A1(new_n1223_), .A2(new_n1146_), .ZN(new_n1224_));
  NAND2_X1   g01160(.A1(new_n1151_), .A2(new_n1157_), .ZN(new_n1225_));
  NAND2_X1   g01161(.A1(new_n1225_), .A2(new_n1201_), .ZN(new_n1226_));
  NAND2_X1   g01162(.A1(new_n1226_), .A2(new_n1224_), .ZN(new_n1227_));
  INV_X1     g01163(.I(new_n1227_), .ZN(new_n1228_));
  XOR2_X1    g01164(.A1(\a[17] ), .A2(\a[18] ), .Z(new_n1229_));
  NOR2_X1    g01165(.A1(new_n1229_), .A2(new_n90_), .ZN(new_n1230_));
  OAI21_X1   g01166(.A1(new_n273_), .A2(new_n1230_), .B(new_n1187_), .ZN(new_n1231_));
  NOR4_X1    g01167(.A1(new_n90_), .A2(new_n68_), .A3(\a[21] ), .A4(\a[22] ), .ZN(new_n1232_));
  NOR3_X1    g01168(.A1(new_n247_), .A2(new_n68_), .A3(new_n1187_), .ZN(new_n1233_));
  OAI21_X1   g01169(.A1(new_n1233_), .A2(new_n1232_), .B(new_n356_), .ZN(new_n1234_));
  NAND2_X1   g01170(.A1(new_n1234_), .A2(new_n1231_), .ZN(new_n1235_));
  INV_X1     g01171(.I(new_n1232_), .ZN(new_n1236_));
  NOR2_X1    g01172(.A1(new_n243_), .A2(\a[23] ), .ZN(new_n1237_));
  NOR2_X1    g01173(.A1(new_n68_), .A2(\a[21] ), .ZN(new_n1238_));
  OAI22_X1   g01174(.A1(new_n1237_), .A2(new_n1238_), .B1(new_n186_), .B2(new_n187_), .ZN(new_n1239_));
  NAND3_X1   g01175(.A1(new_n1239_), .A2(\a[23] ), .A3(new_n1121_), .ZN(new_n1240_));
  NAND3_X1   g01176(.A1(new_n1240_), .A2(new_n273_), .A3(new_n1236_), .ZN(new_n1241_));
  NOR4_X1    g01177(.A1(new_n90_), .A2(new_n68_), .A3(\a[21] ), .A4(\a[22] ), .ZN(new_n1242_));
  INV_X1     g01178(.I(new_n1242_), .ZN(new_n1243_));
  NOR2_X1    g01179(.A1(new_n356_), .A2(new_n1243_), .ZN(new_n1244_));
  AOI21_X1   g01180(.A1(new_n1235_), .A2(new_n1241_), .B(new_n1244_), .ZN(new_n1245_));
  NOR2_X1    g01181(.A1(new_n273_), .A2(new_n1242_), .ZN(new_n1246_));
  NAND3_X1   g01182(.A1(new_n189_), .A2(new_n1186_), .A3(new_n1188_), .ZN(new_n1247_));
  NOR3_X1    g01183(.A1(new_n1239_), .A2(new_n68_), .A3(new_n113_), .ZN(new_n1248_));
  NAND3_X1   g01184(.A1(new_n247_), .A2(\a[23] ), .A3(new_n1121_), .ZN(new_n1249_));
  NOR2_X1    g01185(.A1(new_n189_), .A2(new_n1120_), .ZN(new_n1250_));
  OAI21_X1   g01186(.A1(new_n1250_), .A2(new_n1248_), .B(new_n1249_), .ZN(new_n1251_));
  NAND3_X1   g01187(.A1(new_n1251_), .A2(new_n356_), .A3(new_n1247_), .ZN(new_n1252_));
  OAI21_X1   g01188(.A1(new_n1245_), .A2(new_n1246_), .B(new_n1252_), .ZN(new_n1253_));
  INV_X1     g01189(.I(new_n1247_), .ZN(new_n1254_));
  NAND2_X1   g01190(.A1(new_n189_), .A2(new_n1120_), .ZN(new_n1255_));
  OAI21_X1   g01191(.A1(new_n1239_), .A2(new_n68_), .B(new_n1186_), .ZN(new_n1256_));
  AOI22_X1   g01192(.A1(new_n1255_), .A2(new_n1256_), .B1(new_n189_), .B2(new_n1188_), .ZN(new_n1257_));
  OAI21_X1   g01193(.A1(new_n1257_), .A2(new_n1254_), .B(new_n273_), .ZN(new_n1258_));
  NAND3_X1   g01194(.A1(new_n1129_), .A2(new_n189_), .A3(new_n1125_), .ZN(new_n1259_));
  INV_X1     g01195(.I(new_n1259_), .ZN(new_n1260_));
  AOI21_X1   g01196(.A1(new_n1129_), .A2(new_n1125_), .B(new_n189_), .ZN(new_n1261_));
  OAI21_X1   g01197(.A1(new_n1260_), .A2(new_n1261_), .B(new_n1189_), .ZN(new_n1262_));
  OAI21_X1   g01198(.A1(new_n1130_), .A2(new_n1192_), .B(new_n1123_), .ZN(new_n1263_));
  AOI21_X1   g01199(.A1(new_n1262_), .A2(new_n1263_), .B(new_n356_), .ZN(new_n1264_));
  AOI21_X1   g01200(.A1(new_n1253_), .A2(new_n1258_), .B(new_n1264_), .ZN(new_n1265_));
  INV_X1     g01201(.I(new_n1261_), .ZN(new_n1266_));
  AOI21_X1   g01202(.A1(new_n1266_), .A2(new_n1259_), .B(new_n1123_), .ZN(new_n1267_));
  AOI21_X1   g01203(.A1(new_n1191_), .A2(new_n1131_), .B(new_n1189_), .ZN(new_n1268_));
  NOR3_X1    g01204(.A1(new_n1267_), .A2(new_n273_), .A3(new_n1268_), .ZN(new_n1269_));
  XOR2_X1    g01205(.A1(new_n189_), .A2(new_n1134_), .Z(new_n1270_));
  NAND2_X1   g01206(.A1(new_n1132_), .A2(new_n1270_), .ZN(new_n1271_));
  NAND2_X1   g01207(.A1(new_n1194_), .A2(new_n1136_), .ZN(new_n1272_));
  NAND2_X1   g01208(.A1(new_n1193_), .A2(new_n1272_), .ZN(new_n1273_));
  NAND2_X1   g01209(.A1(new_n1273_), .A2(new_n1271_), .ZN(new_n1274_));
  NAND2_X1   g01210(.A1(new_n1274_), .A2(new_n356_), .ZN(new_n1275_));
  OAI21_X1   g01211(.A1(new_n1265_), .A2(new_n1269_), .B(new_n1275_), .ZN(new_n1276_));
  NAND3_X1   g01212(.A1(new_n1273_), .A2(new_n1271_), .A3(new_n273_), .ZN(new_n1277_));
  NOR2_X1    g01213(.A1(new_n1143_), .A2(new_n1140_), .ZN(new_n1278_));
  NOR2_X1    g01214(.A1(new_n1278_), .A2(new_n248_), .ZN(new_n1279_));
  NAND2_X1   g01215(.A1(new_n1198_), .A2(new_n1139_), .ZN(new_n1280_));
  NOR2_X1    g01216(.A1(new_n1280_), .A2(new_n189_), .ZN(new_n1281_));
  OAI21_X1   g01217(.A1(new_n1279_), .A2(new_n1281_), .B(new_n1195_), .ZN(new_n1282_));
  NAND2_X1   g01218(.A1(new_n1145_), .A2(new_n1199_), .ZN(new_n1283_));
  NAND2_X1   g01219(.A1(new_n1283_), .A2(new_n1138_), .ZN(new_n1284_));
  NAND3_X1   g01220(.A1(new_n1282_), .A2(new_n1284_), .A3(new_n273_), .ZN(new_n1285_));
  NAND2_X1   g01221(.A1(new_n1280_), .A2(new_n189_), .ZN(new_n1286_));
  NAND2_X1   g01222(.A1(new_n1278_), .A2(new_n248_), .ZN(new_n1287_));
  AOI21_X1   g01223(.A1(new_n1286_), .A2(new_n1287_), .B(new_n1138_), .ZN(new_n1288_));
  AOI21_X1   g01224(.A1(new_n1199_), .A2(new_n1145_), .B(new_n1195_), .ZN(new_n1289_));
  OAI21_X1   g01225(.A1(new_n1289_), .A2(new_n1288_), .B(new_n356_), .ZN(new_n1290_));
  NAND4_X1   g01226(.A1(new_n1276_), .A2(new_n1277_), .A3(new_n1285_), .A4(new_n1290_), .ZN(new_n1291_));
  NOR2_X1    g01227(.A1(new_n1291_), .A2(new_n1228_), .ZN(new_n1292_));
  AOI21_X1   g01228(.A1(new_n1282_), .A2(new_n1284_), .B(new_n273_), .ZN(new_n1293_));
  NAND2_X1   g01229(.A1(new_n1293_), .A2(new_n273_), .ZN(new_n1294_));
  AOI21_X1   g01230(.A1(new_n1291_), .A2(new_n1228_), .B(new_n1294_), .ZN(new_n1295_));
  AOI21_X1   g01231(.A1(new_n1207_), .A2(new_n1165_), .B(new_n1159_), .ZN(new_n1296_));
  NOR3_X1    g01232(.A1(new_n1206_), .A2(new_n1205_), .A3(new_n248_), .ZN(new_n1297_));
  AOI21_X1   g01233(.A1(new_n1161_), .A2(new_n1163_), .B(new_n189_), .ZN(new_n1298_));
  NOR2_X1    g01234(.A1(new_n1297_), .A2(new_n1298_), .ZN(new_n1299_));
  NOR2_X1    g01235(.A1(new_n1299_), .A2(new_n1203_), .ZN(new_n1300_));
  NOR3_X1    g01236(.A1(new_n1296_), .A2(new_n1300_), .A3(new_n273_), .ZN(new_n1301_));
  NAND2_X1   g01237(.A1(new_n1191_), .A2(new_n1189_), .ZN(new_n1302_));
  AOI21_X1   g01238(.A1(new_n1302_), .A2(new_n1131_), .B(new_n1135_), .ZN(new_n1303_));
  OAI21_X1   g01239(.A1(new_n1303_), .A2(new_n1137_), .B(new_n1199_), .ZN(new_n1304_));
  AOI21_X1   g01240(.A1(new_n1304_), .A2(new_n1145_), .B(new_n1202_), .ZN(new_n1305_));
  OAI22_X1   g01241(.A1(new_n1305_), .A2(new_n1158_), .B1(new_n1208_), .B2(new_n1164_), .ZN(new_n1306_));
  NAND3_X1   g01242(.A1(new_n1161_), .A2(new_n189_), .A3(new_n1163_), .ZN(new_n1307_));
  OAI21_X1   g01243(.A1(new_n1206_), .A2(new_n1205_), .B(new_n248_), .ZN(new_n1308_));
  NAND2_X1   g01244(.A1(new_n1308_), .A2(new_n1307_), .ZN(new_n1309_));
  NAND2_X1   g01245(.A1(new_n1309_), .A2(new_n1159_), .ZN(new_n1310_));
  AOI21_X1   g01246(.A1(new_n1310_), .A2(new_n1306_), .B(new_n356_), .ZN(new_n1311_));
  NAND2_X1   g01247(.A1(new_n1129_), .A2(new_n1125_), .ZN(new_n1312_));
  AOI21_X1   g01248(.A1(new_n1312_), .A2(new_n189_), .B(new_n1123_), .ZN(new_n1313_));
  OAI21_X1   g01249(.A1(new_n1313_), .A2(new_n1192_), .B(new_n1136_), .ZN(new_n1314_));
  AOI21_X1   g01250(.A1(new_n1314_), .A2(new_n1194_), .B(new_n1144_), .ZN(new_n1315_));
  OAI21_X1   g01251(.A1(new_n1315_), .A2(new_n1200_), .B(new_n1151_), .ZN(new_n1316_));
  AOI21_X1   g01252(.A1(new_n1316_), .A2(new_n1157_), .B(new_n1164_), .ZN(new_n1317_));
  NOR3_X1    g01253(.A1(new_n1212_), .A2(new_n1317_), .A3(new_n1208_), .ZN(new_n1318_));
  NOR2_X1    g01254(.A1(new_n1209_), .A2(new_n1176_), .ZN(new_n1319_));
  NOR3_X1    g01255(.A1(new_n1319_), .A2(new_n1318_), .A3(new_n356_), .ZN(new_n1320_));
  OAI21_X1   g01256(.A1(new_n1305_), .A2(new_n1158_), .B(new_n1207_), .ZN(new_n1321_));
  NAND4_X1   g01257(.A1(new_n1321_), .A2(new_n1165_), .A3(new_n1210_), .A4(new_n1211_), .ZN(new_n1322_));
  NAND2_X1   g01258(.A1(new_n1166_), .A2(new_n1212_), .ZN(new_n1323_));
  AOI21_X1   g01259(.A1(new_n1323_), .A2(new_n1322_), .B(new_n273_), .ZN(new_n1324_));
  OAI22_X1   g01260(.A1(new_n1295_), .A2(new_n1292_), .B1(new_n1301_), .B2(new_n1311_), .ZN(new_n1326_));
  NOR2_X1    g01261(.A1(new_n1326_), .A2(new_n1220_), .ZN(new_n1327_));
  NAND2_X1   g01262(.A1(new_n1324_), .A2(new_n356_), .ZN(new_n1328_));
  AOI21_X1   g01263(.A1(new_n1326_), .A2(new_n1220_), .B(new_n1328_), .ZN(new_n1329_));
  NAND2_X1   g01264(.A1(new_n1177_), .A2(new_n1183_), .ZN(new_n1330_));
  NAND3_X1   g01265(.A1(new_n1209_), .A2(new_n1330_), .A3(new_n1212_), .ZN(new_n1331_));
  AOI21_X1   g01266(.A1(new_n1209_), .A2(new_n1212_), .B(new_n1330_), .ZN(new_n1332_));
  NAND2_X1   g01267(.A1(new_n1119_), .A2(new_n248_), .ZN(new_n1333_));
  OAI21_X1   g01268(.A1(new_n1332_), .A2(new_n1333_), .B(new_n1331_), .ZN(new_n1334_));
  INV_X1     g01269(.I(new_n969_), .ZN(new_n1335_));
  INV_X1     g01270(.I(new_n974_), .ZN(new_n1336_));
  AOI22_X1   g01271(.A1(new_n955_), .A2(new_n959_), .B1(new_n1335_), .B2(new_n1336_), .ZN(new_n1337_));
  AOI21_X1   g01272(.A1(new_n1178_), .A2(new_n1172_), .B(new_n953_), .ZN(new_n1338_));
  NOR3_X1    g01273(.A1(new_n973_), .A2(new_n118_), .A3(new_n963_), .ZN(new_n1339_));
  AOI21_X1   g01274(.A1(new_n968_), .A2(new_n964_), .B(new_n71_), .ZN(new_n1340_));
  NOR2_X1    g01275(.A1(new_n1339_), .A2(new_n1340_), .ZN(new_n1341_));
  NOR3_X1    g01276(.A1(new_n1338_), .A2(new_n1341_), .A3(new_n958_), .ZN(new_n1342_));
  NOR3_X1    g01277(.A1(new_n1337_), .A2(new_n1342_), .A3(new_n248_), .ZN(new_n1343_));
  OAI22_X1   g01278(.A1(new_n1338_), .A2(new_n958_), .B1(new_n969_), .B2(new_n974_), .ZN(new_n1344_));
  INV_X1     g01279(.I(new_n1341_), .ZN(new_n1345_));
  NAND3_X1   g01280(.A1(new_n1345_), .A2(new_n955_), .A3(new_n959_), .ZN(new_n1346_));
  AOI21_X1   g01281(.A1(new_n1344_), .A2(new_n1346_), .B(new_n189_), .ZN(new_n1347_));
  NOR2_X1    g01282(.A1(new_n1347_), .A2(new_n1343_), .ZN(new_n1348_));
  NOR2_X1    g01283(.A1(new_n1334_), .A2(new_n1348_), .ZN(new_n1349_));
  NOR3_X1    g01284(.A1(new_n1166_), .A2(new_n1176_), .A3(new_n1218_), .ZN(new_n1350_));
  OAI21_X1   g01285(.A1(new_n1166_), .A2(new_n1176_), .B(new_n1218_), .ZN(new_n1351_));
  INV_X1     g01286(.I(new_n1333_), .ZN(new_n1352_));
  AOI21_X1   g01287(.A1(new_n1352_), .A2(new_n1351_), .B(new_n1350_), .ZN(new_n1353_));
  NAND3_X1   g01288(.A1(new_n1344_), .A2(new_n1346_), .A3(new_n189_), .ZN(new_n1354_));
  OAI21_X1   g01289(.A1(new_n1337_), .A2(new_n1342_), .B(new_n248_), .ZN(new_n1355_));
  NAND2_X1   g01290(.A1(new_n1355_), .A2(new_n1354_), .ZN(new_n1356_));
  NOR2_X1    g01291(.A1(new_n1353_), .A2(new_n1356_), .ZN(new_n1357_));
  OAI21_X1   g01292(.A1(new_n1349_), .A2(new_n1357_), .B(new_n356_), .ZN(new_n1358_));
  OAI21_X1   g01293(.A1(new_n1327_), .A2(new_n1329_), .B(new_n1358_), .ZN(new_n1359_));
  NAND2_X1   g01294(.A1(new_n1353_), .A2(new_n1356_), .ZN(new_n1360_));
  NAND2_X1   g01295(.A1(new_n1334_), .A2(new_n1348_), .ZN(new_n1361_));
  NAND3_X1   g01296(.A1(new_n1361_), .A2(new_n1360_), .A3(new_n273_), .ZN(new_n1362_));
  OAI21_X1   g01297(.A1(new_n1338_), .A2(new_n958_), .B(new_n1335_), .ZN(new_n1363_));
  INV_X1     g01298(.I(new_n978_), .ZN(new_n1364_));
  AOI22_X1   g01299(.A1(new_n1363_), .A2(new_n1336_), .B1(new_n1364_), .B2(new_n980_), .ZN(new_n1365_));
  XOR2_X1    g01300(.A1(new_n976_), .A2(new_n118_), .Z(new_n1366_));
  NOR3_X1    g01301(.A1(new_n970_), .A2(new_n974_), .A3(new_n1366_), .ZN(new_n1367_));
  NOR3_X1    g01302(.A1(new_n1365_), .A2(new_n1367_), .A3(new_n248_), .ZN(new_n1368_));
  OAI22_X1   g01303(.A1(new_n970_), .A2(new_n974_), .B1(new_n978_), .B2(new_n979_), .ZN(new_n1369_));
  INV_X1     g01304(.I(new_n1366_), .ZN(new_n1370_));
  NAND3_X1   g01305(.A1(new_n1363_), .A2(new_n1336_), .A3(new_n1370_), .ZN(new_n1371_));
  AOI21_X1   g01306(.A1(new_n1369_), .A2(new_n1371_), .B(new_n189_), .ZN(new_n1372_));
  NOR3_X1    g01307(.A1(new_n1368_), .A2(new_n1372_), .A3(new_n1343_), .ZN(new_n1373_));
  NOR3_X1    g01308(.A1(new_n1373_), .A2(new_n1334_), .A3(new_n1348_), .ZN(new_n1374_));
  NAND3_X1   g01309(.A1(new_n1369_), .A2(new_n1371_), .A3(new_n189_), .ZN(new_n1375_));
  OAI21_X1   g01310(.A1(new_n1365_), .A2(new_n1367_), .B(new_n248_), .ZN(new_n1376_));
  NAND3_X1   g01311(.A1(new_n1376_), .A2(new_n1375_), .A3(new_n1354_), .ZN(new_n1377_));
  AOI21_X1   g01312(.A1(new_n1377_), .A2(new_n1356_), .B(new_n1353_), .ZN(new_n1378_));
  OAI21_X1   g01313(.A1(new_n1374_), .A2(new_n1378_), .B(new_n356_), .ZN(new_n1379_));
  NAND3_X1   g01314(.A1(new_n1377_), .A2(new_n1353_), .A3(new_n1356_), .ZN(new_n1380_));
  OAI21_X1   g01315(.A1(new_n1373_), .A2(new_n1348_), .B(new_n1334_), .ZN(new_n1381_));
  NAND3_X1   g01316(.A1(new_n1381_), .A2(new_n1380_), .A3(new_n273_), .ZN(new_n1382_));
  AOI22_X1   g01317(.A1(new_n1359_), .A2(new_n1362_), .B1(new_n1379_), .B2(new_n1382_), .ZN(new_n1383_));
  INV_X1     g01318(.I(new_n1118_), .ZN(new_n1384_));
  NAND2_X1   g01319(.A1(new_n1384_), .A2(new_n189_), .ZN(new_n1385_));
  AOI21_X1   g01320(.A1(new_n1209_), .A2(new_n1212_), .B(new_n1215_), .ZN(new_n1386_));
  NOR3_X1    g01321(.A1(new_n1166_), .A2(new_n1176_), .A3(new_n1184_), .ZN(new_n1387_));
  OAI21_X1   g01322(.A1(new_n1386_), .A2(new_n1387_), .B(new_n1385_), .ZN(new_n1388_));
  INV_X1     g01323(.I(new_n1219_), .ZN(new_n1389_));
  NAND2_X1   g01324(.A1(new_n1388_), .A2(new_n1389_), .ZN(new_n1390_));
  NOR3_X1    g01325(.A1(new_n1233_), .A2(new_n356_), .A3(new_n1232_), .ZN(new_n1391_));
  AOI21_X1   g01326(.A1(new_n1231_), .A2(new_n1234_), .B(new_n1391_), .ZN(new_n1392_));
  INV_X1     g01327(.I(new_n1246_), .ZN(new_n1393_));
  OAI21_X1   g01328(.A1(new_n1392_), .A2(new_n1244_), .B(new_n1393_), .ZN(new_n1394_));
  AOI21_X1   g01329(.A1(new_n1251_), .A2(new_n1247_), .B(new_n356_), .ZN(new_n1395_));
  AOI21_X1   g01330(.A1(new_n1394_), .A2(new_n1252_), .B(new_n1395_), .ZN(new_n1396_));
  NAND3_X1   g01331(.A1(new_n1262_), .A2(new_n356_), .A3(new_n1263_), .ZN(new_n1397_));
  OAI21_X1   g01332(.A1(new_n1396_), .A2(new_n1264_), .B(new_n1397_), .ZN(new_n1398_));
  INV_X1     g01333(.I(new_n1277_), .ZN(new_n1399_));
  AOI21_X1   g01334(.A1(new_n1398_), .A2(new_n1275_), .B(new_n1399_), .ZN(new_n1400_));
  NOR3_X1    g01335(.A1(new_n1289_), .A2(new_n1288_), .A3(new_n356_), .ZN(new_n1401_));
  NOR2_X1    g01336(.A1(new_n1401_), .A2(new_n1293_), .ZN(new_n1402_));
  NAND3_X1   g01337(.A1(new_n1402_), .A2(new_n1400_), .A3(new_n1227_), .ZN(new_n1403_));
  INV_X1     g01338(.I(new_n1231_), .ZN(new_n1404_));
  AOI21_X1   g01339(.A1(new_n1240_), .A2(new_n1236_), .B(new_n273_), .ZN(new_n1405_));
  NOR2_X1    g01340(.A1(new_n1404_), .A2(new_n1405_), .ZN(new_n1406_));
  INV_X1     g01341(.I(new_n1244_), .ZN(new_n1407_));
  OAI21_X1   g01342(.A1(new_n1406_), .A2(new_n1391_), .B(new_n1407_), .ZN(new_n1408_));
  NOR2_X1    g01343(.A1(new_n1257_), .A2(new_n1254_), .ZN(new_n1409_));
  AOI22_X1   g01344(.A1(new_n1408_), .A2(new_n1393_), .B1(new_n356_), .B2(new_n1409_), .ZN(new_n1410_));
  OAI21_X1   g01345(.A1(new_n1267_), .A2(new_n1268_), .B(new_n273_), .ZN(new_n1411_));
  OAI21_X1   g01346(.A1(new_n1410_), .A2(new_n1395_), .B(new_n1411_), .ZN(new_n1412_));
  AOI21_X1   g01347(.A1(new_n1273_), .A2(new_n1271_), .B(new_n273_), .ZN(new_n1413_));
  AOI21_X1   g01348(.A1(new_n1412_), .A2(new_n1397_), .B(new_n1413_), .ZN(new_n1414_));
  NAND2_X1   g01349(.A1(new_n1290_), .A2(new_n1285_), .ZN(new_n1415_));
  NOR3_X1    g01350(.A1(new_n1415_), .A2(new_n1414_), .A3(new_n1399_), .ZN(new_n1416_));
  INV_X1     g01351(.I(new_n1294_), .ZN(new_n1417_));
  OAI21_X1   g01352(.A1(new_n1416_), .A2(new_n1227_), .B(new_n1417_), .ZN(new_n1418_));
  NAND3_X1   g01353(.A1(new_n1310_), .A2(new_n1306_), .A3(new_n356_), .ZN(new_n1419_));
  OAI21_X1   g01354(.A1(new_n1296_), .A2(new_n1300_), .B(new_n273_), .ZN(new_n1420_));
  AOI22_X1   g01355(.A1(new_n1418_), .A2(new_n1403_), .B1(new_n1419_), .B2(new_n1420_), .ZN(new_n1421_));
  NAND2_X1   g01356(.A1(new_n1421_), .A2(new_n1390_), .ZN(new_n1422_));
  OAI21_X1   g01357(.A1(new_n1319_), .A2(new_n1318_), .B(new_n356_), .ZN(new_n1423_));
  NOR2_X1    g01358(.A1(new_n1423_), .A2(new_n273_), .ZN(new_n1424_));
  OAI21_X1   g01359(.A1(new_n1421_), .A2(new_n1390_), .B(new_n1424_), .ZN(new_n1425_));
  AOI21_X1   g01360(.A1(new_n1361_), .A2(new_n1360_), .B(new_n273_), .ZN(new_n1426_));
  AOI21_X1   g01361(.A1(new_n1425_), .A2(new_n1422_), .B(new_n1426_), .ZN(new_n1427_));
  NOR3_X1    g01362(.A1(new_n1349_), .A2(new_n1357_), .A3(new_n356_), .ZN(new_n1428_));
  NOR3_X1    g01363(.A1(new_n1374_), .A2(new_n1378_), .A3(new_n273_), .ZN(new_n1429_));
  AOI21_X1   g01364(.A1(new_n1381_), .A2(new_n1380_), .B(new_n356_), .ZN(new_n1430_));
  NOR2_X1    g01365(.A1(new_n1429_), .A2(new_n1430_), .ZN(new_n1431_));
  NOR3_X1    g01366(.A1(new_n1431_), .A2(new_n1427_), .A3(new_n1428_), .ZN(new_n1432_));
  NOR3_X1    g01367(.A1(new_n1432_), .A2(new_n568_), .A3(new_n1383_), .ZN(new_n1433_));
  NAND3_X1   g01368(.A1(new_n1326_), .A2(new_n1390_), .A3(new_n356_), .ZN(new_n1434_));
  OAI21_X1   g01369(.A1(new_n273_), .A2(new_n1220_), .B(new_n1421_), .ZN(new_n1435_));
  AOI21_X1   g01370(.A1(new_n1435_), .A2(new_n1434_), .B(new_n1324_), .ZN(new_n1436_));
  NOR3_X1    g01371(.A1(new_n1421_), .A2(new_n273_), .A3(new_n1220_), .ZN(new_n1437_));
  AOI21_X1   g01372(.A1(new_n356_), .A2(new_n1390_), .B(new_n1326_), .ZN(new_n1438_));
  NOR3_X1    g01373(.A1(new_n1437_), .A2(new_n1438_), .A3(new_n1423_), .ZN(new_n1439_));
  NOR2_X1    g01374(.A1(new_n1436_), .A2(new_n1439_), .ZN(new_n1440_));
  AOI21_X1   g01375(.A1(new_n1402_), .A2(new_n1400_), .B(new_n1227_), .ZN(new_n1441_));
  OAI21_X1   g01376(.A1(new_n1441_), .A2(new_n1294_), .B(new_n1403_), .ZN(new_n1442_));
  NOR2_X1    g01377(.A1(new_n1301_), .A2(new_n1311_), .ZN(new_n1443_));
  NOR2_X1    g01378(.A1(new_n1442_), .A2(new_n1443_), .ZN(new_n1444_));
  NAND2_X1   g01379(.A1(new_n1420_), .A2(new_n1419_), .ZN(new_n1445_));
  AOI21_X1   g01380(.A1(new_n1418_), .A2(new_n1403_), .B(new_n1445_), .ZN(new_n1446_));
  NOR2_X1    g01381(.A1(new_n1444_), .A2(new_n1446_), .ZN(new_n1447_));
  INV_X1     g01382(.I(new_n1447_), .ZN(new_n1448_));
  NOR3_X1    g01383(.A1(new_n1320_), .A2(new_n1324_), .A3(new_n1301_), .ZN(new_n1449_));
  NOR3_X1    g01384(.A1(new_n1449_), .A2(new_n1442_), .A3(new_n1443_), .ZN(new_n1450_));
  NOR2_X1    g01385(.A1(new_n1295_), .A2(new_n1292_), .ZN(new_n1451_));
  NAND3_X1   g01386(.A1(new_n1323_), .A2(new_n1322_), .A3(new_n273_), .ZN(new_n1452_));
  NAND3_X1   g01387(.A1(new_n1423_), .A2(new_n1452_), .A3(new_n1419_), .ZN(new_n1453_));
  AOI21_X1   g01388(.A1(new_n1453_), .A2(new_n1445_), .B(new_n1451_), .ZN(new_n1454_));
  NOR2_X1    g01389(.A1(new_n1450_), .A2(new_n1454_), .ZN(new_n1455_));
  AOI21_X1   g01390(.A1(new_n1455_), .A2(new_n1448_), .B(new_n568_), .ZN(new_n1456_));
  NAND3_X1   g01391(.A1(new_n1262_), .A2(new_n273_), .A3(new_n1263_), .ZN(new_n1457_));
  OAI21_X1   g01392(.A1(new_n1267_), .A2(new_n1268_), .B(new_n356_), .ZN(new_n1458_));
  AND2_X2    g01393(.A1(new_n1458_), .A2(new_n1457_), .Z(new_n1459_));
  OAI21_X1   g01394(.A1(new_n1264_), .A2(new_n1269_), .B(new_n1396_), .ZN(new_n1460_));
  OAI21_X1   g01395(.A1(new_n1459_), .A2(new_n1396_), .B(new_n1460_), .ZN(new_n1461_));
  NOR3_X1    g01396(.A1(new_n1233_), .A2(new_n273_), .A3(new_n1232_), .ZN(new_n1462_));
  AOI21_X1   g01397(.A1(new_n1240_), .A2(new_n1236_), .B(new_n356_), .ZN(new_n1463_));
  OAI21_X1   g01398(.A1(new_n1462_), .A2(new_n1463_), .B(new_n1231_), .ZN(new_n1464_));
  OAI21_X1   g01399(.A1(new_n1405_), .A2(new_n1391_), .B(new_n1404_), .ZN(new_n1465_));
  NAND2_X1   g01400(.A1(new_n1465_), .A2(new_n1464_), .ZN(new_n1466_));
  XNOR2_X1   g01401(.A1(\a[17] ), .A2(\a[18] ), .ZN(new_n1467_));
  XNOR2_X1   g01402(.A1(\a[14] ), .A2(\a[15] ), .ZN(new_n1468_));
  NAND2_X1   g01403(.A1(new_n1468_), .A2(\a[17] ), .ZN(new_n1469_));
  AOI21_X1   g01404(.A1(new_n443_), .A2(new_n1469_), .B(new_n1467_), .ZN(new_n1470_));
  INV_X1     g01405(.I(new_n1470_), .ZN(new_n1471_));
  NAND4_X1   g01406(.A1(new_n268_), .A2(new_n270_), .A3(\a[17] ), .A4(\a[20] ), .ZN(new_n1472_));
  INV_X1     g01407(.I(new_n1472_), .ZN(new_n1473_));
  NAND2_X1   g01408(.A1(new_n1467_), .A2(\a[20] ), .ZN(new_n1474_));
  NOR2_X1    g01409(.A1(new_n356_), .A2(new_n1474_), .ZN(new_n1475_));
  OAI21_X1   g01410(.A1(new_n1475_), .A2(new_n1473_), .B(new_n443_), .ZN(new_n1476_));
  NAND2_X1   g01411(.A1(new_n1476_), .A2(new_n1471_), .ZN(new_n1477_));
  NAND2_X1   g01412(.A1(new_n273_), .A2(new_n1230_), .ZN(new_n1478_));
  NAND3_X1   g01413(.A1(new_n1478_), .A2(new_n568_), .A3(new_n1472_), .ZN(new_n1479_));
  NAND4_X1   g01414(.A1(new_n268_), .A2(new_n270_), .A3(\a[17] ), .A4(\a[20] ), .ZN(new_n1480_));
  NOR2_X1    g01415(.A1(new_n443_), .A2(new_n1480_), .ZN(new_n1481_));
  INV_X1     g01416(.I(new_n1481_), .ZN(new_n1482_));
  NAND2_X1   g01417(.A1(new_n443_), .A2(new_n1480_), .ZN(new_n1483_));
  NAND3_X1   g01418(.A1(new_n356_), .A2(new_n1187_), .A3(new_n1230_), .ZN(new_n1484_));
  INV_X1     g01419(.I(new_n1484_), .ZN(new_n1485_));
  NOR4_X1    g01420(.A1(new_n355_), .A2(\a[18] ), .A3(new_n90_), .A4(new_n243_), .ZN(new_n1486_));
  INV_X1     g01421(.I(new_n1486_), .ZN(new_n1487_));
  NOR4_X1    g01422(.A1(new_n270_), .A2(new_n90_), .A3(\a[17] ), .A4(\a[18] ), .ZN(new_n1488_));
  NAND2_X1   g01423(.A1(new_n273_), .A2(new_n1187_), .ZN(new_n1489_));
  AOI21_X1   g01424(.A1(new_n1487_), .A2(new_n1489_), .B(new_n1488_), .ZN(new_n1490_));
  NOR3_X1    g01425(.A1(new_n1490_), .A2(new_n443_), .A3(new_n1485_), .ZN(new_n1491_));
  INV_X1     g01426(.I(new_n1488_), .ZN(new_n1492_));
  NOR2_X1    g01427(.A1(new_n356_), .A2(new_n1121_), .ZN(new_n1493_));
  OAI21_X1   g01428(.A1(new_n1493_), .A2(new_n1486_), .B(new_n1492_), .ZN(new_n1494_));
  AOI21_X1   g01429(.A1(new_n1494_), .A2(new_n1484_), .B(new_n568_), .ZN(new_n1495_));
  AOI22_X1   g01430(.A1(new_n1477_), .A2(new_n1479_), .B1(new_n1482_), .B2(new_n1483_), .ZN(new_n1497_));
  NAND2_X1   g01431(.A1(new_n1497_), .A2(new_n1466_), .ZN(new_n1498_));
  NAND3_X1   g01432(.A1(new_n1494_), .A2(new_n443_), .A3(new_n1484_), .ZN(new_n1499_));
  INV_X1     g01433(.I(new_n1499_), .ZN(new_n1500_));
  OAI21_X1   g01434(.A1(new_n1497_), .A2(new_n1466_), .B(new_n1500_), .ZN(new_n1501_));
  XOR2_X1    g01435(.A1(new_n273_), .A2(new_n1243_), .Z(new_n1502_));
  INV_X1     g01436(.I(new_n1502_), .ZN(new_n1503_));
  OAI21_X1   g01437(.A1(new_n1406_), .A2(new_n1391_), .B(new_n1503_), .ZN(new_n1504_));
  NOR2_X1    g01438(.A1(new_n1244_), .A2(new_n1246_), .ZN(new_n1505_));
  INV_X1     g01439(.I(new_n1505_), .ZN(new_n1506_));
  NAND2_X1   g01440(.A1(new_n1392_), .A2(new_n1506_), .ZN(new_n1507_));
  NAND2_X1   g01441(.A1(new_n1504_), .A2(new_n1507_), .ZN(new_n1508_));
  AOI22_X1   g01442(.A1(new_n1501_), .A2(new_n1498_), .B1(new_n1508_), .B2(new_n443_), .ZN(new_n1509_));
  NAND3_X1   g01443(.A1(new_n1504_), .A2(new_n1507_), .A3(new_n568_), .ZN(new_n1510_));
  INV_X1     g01444(.I(new_n1510_), .ZN(new_n1511_));
  OAI21_X1   g01445(.A1(new_n1257_), .A2(new_n1254_), .B(new_n356_), .ZN(new_n1512_));
  NAND3_X1   g01446(.A1(new_n1251_), .A2(new_n273_), .A3(new_n1247_), .ZN(new_n1513_));
  AOI22_X1   g01447(.A1(new_n1408_), .A2(new_n1393_), .B1(new_n1512_), .B2(new_n1513_), .ZN(new_n1514_));
  AOI21_X1   g01448(.A1(new_n1252_), .A2(new_n1258_), .B(new_n1394_), .ZN(new_n1515_));
  NOR3_X1    g01449(.A1(new_n1515_), .A2(new_n1514_), .A3(new_n443_), .ZN(new_n1516_));
  NAND2_X1   g01450(.A1(new_n1512_), .A2(new_n1513_), .ZN(new_n1517_));
  NAND2_X1   g01451(.A1(new_n1517_), .A2(new_n1394_), .ZN(new_n1518_));
  NAND2_X1   g01452(.A1(new_n1258_), .A2(new_n1252_), .ZN(new_n1519_));
  NAND3_X1   g01453(.A1(new_n1519_), .A2(new_n1408_), .A3(new_n1393_), .ZN(new_n1520_));
  AOI21_X1   g01454(.A1(new_n1520_), .A2(new_n1518_), .B(new_n568_), .ZN(new_n1521_));
  NOR4_X1    g01455(.A1(new_n1509_), .A2(new_n1516_), .A3(new_n1521_), .A4(new_n1511_), .ZN(new_n1522_));
  NAND2_X1   g01456(.A1(new_n1522_), .A2(new_n1461_), .ZN(new_n1523_));
  OAI21_X1   g01457(.A1(new_n1515_), .A2(new_n1514_), .B(new_n443_), .ZN(new_n1524_));
  NOR2_X1    g01458(.A1(new_n1524_), .A2(new_n443_), .ZN(new_n1525_));
  OAI21_X1   g01459(.A1(new_n1522_), .A2(new_n1461_), .B(new_n1525_), .ZN(new_n1526_));
  AOI22_X1   g01460(.A1(new_n1412_), .A2(new_n1397_), .B1(new_n1277_), .B2(new_n1275_), .ZN(new_n1527_));
  NAND3_X1   g01461(.A1(new_n1273_), .A2(new_n1271_), .A3(new_n356_), .ZN(new_n1528_));
  NAND2_X1   g01462(.A1(new_n1274_), .A2(new_n273_), .ZN(new_n1529_));
  AOI21_X1   g01463(.A1(new_n1528_), .A2(new_n1529_), .B(new_n1398_), .ZN(new_n1530_));
  NOR3_X1    g01464(.A1(new_n1530_), .A2(new_n1527_), .A3(new_n568_), .ZN(new_n1531_));
  AOI21_X1   g01465(.A1(new_n1526_), .A2(new_n1523_), .B(new_n1531_), .ZN(new_n1532_));
  NOR2_X1    g01466(.A1(new_n1530_), .A2(new_n1527_), .ZN(new_n1533_));
  NOR2_X1    g01467(.A1(new_n1533_), .A2(new_n443_), .ZN(new_n1534_));
  NOR2_X1    g01468(.A1(new_n1265_), .A2(new_n1269_), .ZN(new_n1535_));
  OAI21_X1   g01469(.A1(new_n1535_), .A2(new_n1413_), .B(new_n1277_), .ZN(new_n1536_));
  NAND2_X1   g01470(.A1(new_n1536_), .A2(new_n1415_), .ZN(new_n1537_));
  NAND3_X1   g01471(.A1(new_n1537_), .A2(new_n443_), .A3(new_n1291_), .ZN(new_n1538_));
  OAI21_X1   g01472(.A1(new_n1532_), .A2(new_n1534_), .B(new_n1538_), .ZN(new_n1539_));
  NAND2_X1   g01473(.A1(new_n1537_), .A2(new_n1291_), .ZN(new_n1540_));
  NAND2_X1   g01474(.A1(new_n1540_), .A2(new_n568_), .ZN(new_n1541_));
  AOI22_X1   g01475(.A1(new_n1304_), .A2(new_n1145_), .B1(new_n1222_), .B2(new_n1221_), .ZN(new_n1542_));
  AOI21_X1   g01476(.A1(new_n1151_), .A2(new_n1157_), .B(new_n1146_), .ZN(new_n1543_));
  OAI21_X1   g01477(.A1(new_n1543_), .A2(new_n1542_), .B(new_n273_), .ZN(new_n1544_));
  AOI21_X1   g01478(.A1(new_n1400_), .A2(new_n1402_), .B(new_n1544_), .ZN(new_n1545_));
  AOI21_X1   g01479(.A1(new_n1226_), .A2(new_n1224_), .B(new_n356_), .ZN(new_n1546_));
  NOR3_X1    g01480(.A1(new_n1536_), .A2(new_n1546_), .A3(new_n1415_), .ZN(new_n1547_));
  OAI21_X1   g01481(.A1(new_n1547_), .A2(new_n1545_), .B(new_n1290_), .ZN(new_n1548_));
  OAI21_X1   g01482(.A1(new_n1536_), .A2(new_n1415_), .B(new_n1546_), .ZN(new_n1549_));
  NAND3_X1   g01483(.A1(new_n1402_), .A2(new_n1544_), .A3(new_n1400_), .ZN(new_n1550_));
  NAND3_X1   g01484(.A1(new_n1549_), .A2(new_n1550_), .A3(new_n1293_), .ZN(new_n1551_));
  NAND2_X1   g01485(.A1(new_n1548_), .A2(new_n1551_), .ZN(new_n1552_));
  AOI22_X1   g01486(.A1(new_n1539_), .A2(new_n1541_), .B1(new_n1552_), .B2(new_n568_), .ZN(new_n1553_));
  NOR2_X1    g01487(.A1(new_n1552_), .A2(new_n568_), .ZN(new_n1554_));
  NOR2_X1    g01488(.A1(new_n1553_), .A2(new_n1554_), .ZN(new_n1555_));
  NOR3_X1    g01489(.A1(new_n1450_), .A2(new_n1454_), .A3(new_n568_), .ZN(new_n1556_));
  NAND3_X1   g01490(.A1(new_n1453_), .A2(new_n1451_), .A3(new_n1445_), .ZN(new_n1557_));
  OAI21_X1   g01491(.A1(new_n1449_), .A2(new_n1443_), .B(new_n1442_), .ZN(new_n1558_));
  AOI21_X1   g01492(.A1(new_n1558_), .A2(new_n1557_), .B(new_n443_), .ZN(new_n1559_));
  NOR3_X1    g01493(.A1(new_n1556_), .A2(new_n1559_), .A3(new_n1448_), .ZN(new_n1560_));
  NOR4_X1    g01494(.A1(new_n1440_), .A2(new_n1456_), .A3(new_n1560_), .A4(new_n1555_), .ZN(new_n1561_));
  NAND2_X1   g01495(.A1(new_n1558_), .A2(new_n1557_), .ZN(new_n1562_));
  OAI21_X1   g01496(.A1(new_n1562_), .A2(new_n1447_), .B(new_n443_), .ZN(new_n1563_));
  AOI21_X1   g01497(.A1(new_n1457_), .A2(new_n1458_), .B(new_n1396_), .ZN(new_n1564_));
  NOR2_X1    g01498(.A1(new_n1269_), .A2(new_n1264_), .ZN(new_n1565_));
  NOR3_X1    g01499(.A1(new_n1565_), .A2(new_n1410_), .A3(new_n1395_), .ZN(new_n1566_));
  NOR2_X1    g01500(.A1(new_n1566_), .A2(new_n1564_), .ZN(new_n1567_));
  NAND3_X1   g01501(.A1(new_n1240_), .A2(new_n356_), .A3(new_n1236_), .ZN(new_n1568_));
  OAI21_X1   g01502(.A1(new_n1233_), .A2(new_n1232_), .B(new_n273_), .ZN(new_n1569_));
  AOI21_X1   g01503(.A1(new_n1568_), .A2(new_n1569_), .B(new_n1404_), .ZN(new_n1570_));
  AOI21_X1   g01504(.A1(new_n1234_), .A2(new_n1241_), .B(new_n1231_), .ZN(new_n1571_));
  NOR2_X1    g01505(.A1(new_n1570_), .A2(new_n1571_), .ZN(new_n1572_));
  NAND2_X1   g01506(.A1(new_n1478_), .A2(new_n1472_), .ZN(new_n1573_));
  AOI21_X1   g01507(.A1(new_n1573_), .A2(new_n443_), .B(new_n1470_), .ZN(new_n1574_));
  NOR3_X1    g01508(.A1(new_n1475_), .A2(new_n1473_), .A3(new_n443_), .ZN(new_n1575_));
  INV_X1     g01509(.I(new_n1483_), .ZN(new_n1576_));
  OAI22_X1   g01510(.A1(new_n1574_), .A2(new_n1575_), .B1(new_n1481_), .B2(new_n1576_), .ZN(new_n1577_));
  NOR2_X1    g01511(.A1(new_n1577_), .A2(new_n1572_), .ZN(new_n1578_));
  AOI21_X1   g01512(.A1(new_n1577_), .A2(new_n1572_), .B(new_n1499_), .ZN(new_n1579_));
  NOR2_X1    g01513(.A1(new_n1392_), .A2(new_n1502_), .ZN(new_n1580_));
  NOR3_X1    g01514(.A1(new_n1406_), .A2(new_n1391_), .A3(new_n1505_), .ZN(new_n1581_));
  OAI21_X1   g01515(.A1(new_n1580_), .A2(new_n1581_), .B(new_n443_), .ZN(new_n1582_));
  OAI21_X1   g01516(.A1(new_n1579_), .A2(new_n1578_), .B(new_n1582_), .ZN(new_n1583_));
  NAND3_X1   g01517(.A1(new_n1520_), .A2(new_n1518_), .A3(new_n568_), .ZN(new_n1584_));
  NAND4_X1   g01518(.A1(new_n1524_), .A2(new_n1583_), .A3(new_n1584_), .A4(new_n1510_), .ZN(new_n1585_));
  NOR2_X1    g01519(.A1(new_n1585_), .A2(new_n1567_), .ZN(new_n1586_));
  NAND2_X1   g01520(.A1(new_n1521_), .A2(new_n568_), .ZN(new_n1587_));
  AOI21_X1   g01521(.A1(new_n1585_), .A2(new_n1567_), .B(new_n1587_), .ZN(new_n1588_));
  OAI21_X1   g01522(.A1(new_n1413_), .A2(new_n1399_), .B(new_n1398_), .ZN(new_n1589_));
  NAND2_X1   g01523(.A1(new_n1529_), .A2(new_n1528_), .ZN(new_n1590_));
  NAND2_X1   g01524(.A1(new_n1535_), .A2(new_n1590_), .ZN(new_n1591_));
  NAND3_X1   g01525(.A1(new_n1591_), .A2(new_n1589_), .A3(new_n443_), .ZN(new_n1592_));
  OAI21_X1   g01526(.A1(new_n1588_), .A2(new_n1586_), .B(new_n1592_), .ZN(new_n1593_));
  NAND2_X1   g01527(.A1(new_n1591_), .A2(new_n1589_), .ZN(new_n1594_));
  NAND2_X1   g01528(.A1(new_n1594_), .A2(new_n568_), .ZN(new_n1595_));
  NOR2_X1    g01529(.A1(new_n1402_), .A2(new_n1400_), .ZN(new_n1596_));
  NOR3_X1    g01530(.A1(new_n1416_), .A2(new_n1596_), .A3(new_n568_), .ZN(new_n1597_));
  AOI21_X1   g01531(.A1(new_n1593_), .A2(new_n1595_), .B(new_n1597_), .ZN(new_n1598_));
  NOR2_X1    g01532(.A1(new_n1416_), .A2(new_n1596_), .ZN(new_n1599_));
  NOR2_X1    g01533(.A1(new_n1599_), .A2(new_n443_), .ZN(new_n1600_));
  NOR2_X1    g01534(.A1(new_n1598_), .A2(new_n1600_), .ZN(new_n1601_));
  AOI21_X1   g01535(.A1(new_n1549_), .A2(new_n1550_), .B(new_n1293_), .ZN(new_n1602_));
  NOR3_X1    g01536(.A1(new_n1547_), .A2(new_n1545_), .A3(new_n1290_), .ZN(new_n1603_));
  NOR2_X1    g01537(.A1(new_n1603_), .A2(new_n1602_), .ZN(new_n1604_));
  NOR2_X1    g01538(.A1(new_n1604_), .A2(new_n443_), .ZN(new_n1605_));
  NAND2_X1   g01539(.A1(new_n1604_), .A2(new_n443_), .ZN(new_n1606_));
  OAI21_X1   g01540(.A1(new_n1601_), .A2(new_n1605_), .B(new_n1606_), .ZN(new_n1607_));
  NAND3_X1   g01541(.A1(new_n1558_), .A2(new_n1557_), .A3(new_n443_), .ZN(new_n1608_));
  OAI21_X1   g01542(.A1(new_n1450_), .A2(new_n1454_), .B(new_n568_), .ZN(new_n1609_));
  NAND3_X1   g01543(.A1(new_n1609_), .A2(new_n1608_), .A3(new_n1447_), .ZN(new_n1610_));
  NAND3_X1   g01544(.A1(new_n1610_), .A2(new_n1563_), .A3(new_n1607_), .ZN(new_n1611_));
  NAND2_X1   g01545(.A1(new_n1611_), .A2(new_n1440_), .ZN(new_n1612_));
  NAND2_X1   g01546(.A1(new_n1562_), .A2(new_n443_), .ZN(new_n1613_));
  NOR2_X1    g01547(.A1(new_n1613_), .A2(new_n443_), .ZN(new_n1614_));
  AOI21_X1   g01548(.A1(new_n1612_), .A2(new_n1614_), .B(new_n1561_), .ZN(new_n1615_));
  NAND2_X1   g01549(.A1(new_n1358_), .A2(new_n1362_), .ZN(new_n1616_));
  INV_X1     g01550(.I(\a[15] ), .ZN(new_n1617_));
  NOR2_X1    g01551(.A1(new_n1617_), .A2(\a[17] ), .ZN(new_n1618_));
  NOR2_X1    g01552(.A1(new_n126_), .A2(\a[15] ), .ZN(new_n1619_));
  OAI22_X1   g01553(.A1(new_n1618_), .A2(new_n1619_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n1620_));
  NOR3_X1    g01554(.A1(new_n439_), .A2(\a[14] ), .A3(\a[15] ), .ZN(new_n1621_));
  AOI21_X1   g01555(.A1(\a[15] ), .A2(new_n441_), .B(new_n1621_), .ZN(new_n1622_));
  NOR2_X1    g01556(.A1(new_n1620_), .A2(new_n1622_), .ZN(new_n1623_));
  NAND3_X1   g01557(.A1(new_n1425_), .A2(new_n1422_), .A3(new_n1623_), .ZN(new_n1624_));
  INV_X1     g01558(.I(new_n1623_), .ZN(new_n1625_));
  OAI21_X1   g01559(.A1(new_n1329_), .A2(new_n1327_), .B(new_n1625_), .ZN(new_n1626_));
  AOI21_X1   g01560(.A1(new_n1624_), .A2(new_n1626_), .B(new_n1616_), .ZN(new_n1627_));
  NOR2_X1    g01561(.A1(new_n1426_), .A2(new_n1428_), .ZN(new_n1628_));
  NOR3_X1    g01562(.A1(new_n1329_), .A2(new_n1327_), .A3(new_n1625_), .ZN(new_n1629_));
  AOI21_X1   g01563(.A1(new_n1425_), .A2(new_n1422_), .B(new_n1623_), .ZN(new_n1630_));
  NOR3_X1    g01564(.A1(new_n1630_), .A2(new_n1628_), .A3(new_n1629_), .ZN(new_n1631_));
  OAI21_X1   g01565(.A1(new_n1631_), .A2(new_n1627_), .B(new_n126_), .ZN(new_n1632_));
  OAI21_X1   g01566(.A1(new_n1630_), .A2(new_n1629_), .B(new_n1628_), .ZN(new_n1633_));
  NAND3_X1   g01567(.A1(new_n1624_), .A2(new_n1626_), .A3(new_n1616_), .ZN(new_n1634_));
  NAND3_X1   g01568(.A1(new_n1633_), .A2(new_n1634_), .A3(\a[17] ), .ZN(new_n1635_));
  NAND2_X1   g01569(.A1(new_n1632_), .A2(new_n1635_), .ZN(new_n1636_));
  NAND2_X1   g01570(.A1(new_n1616_), .A2(new_n126_), .ZN(new_n1637_));
  NAND2_X1   g01571(.A1(new_n1628_), .A2(\a[17] ), .ZN(new_n1638_));
  AOI22_X1   g01572(.A1(new_n1638_), .A2(new_n1637_), .B1(new_n1624_), .B2(new_n1626_), .ZN(new_n1639_));
  AOI21_X1   g01573(.A1(new_n1381_), .A2(new_n1380_), .B(new_n273_), .ZN(new_n1640_));
  NOR3_X1    g01574(.A1(new_n1374_), .A2(new_n1378_), .A3(new_n356_), .ZN(new_n1641_));
  OAI22_X1   g01575(.A1(new_n1427_), .A2(new_n1428_), .B1(new_n1640_), .B2(new_n1641_), .ZN(new_n1642_));
  NAND3_X1   g01576(.A1(new_n1381_), .A2(new_n1380_), .A3(new_n356_), .ZN(new_n1643_));
  OAI21_X1   g01577(.A1(new_n1374_), .A2(new_n1378_), .B(new_n273_), .ZN(new_n1644_));
  NAND2_X1   g01578(.A1(new_n1644_), .A2(new_n1643_), .ZN(new_n1645_));
  NAND3_X1   g01579(.A1(new_n1645_), .A2(new_n1359_), .A3(new_n1362_), .ZN(new_n1646_));
  NAND3_X1   g01580(.A1(new_n1646_), .A2(new_n1642_), .A3(new_n443_), .ZN(new_n1647_));
  OAI21_X1   g01581(.A1(new_n1432_), .A2(new_n1383_), .B(new_n568_), .ZN(new_n1648_));
  NAND2_X1   g01582(.A1(new_n1648_), .A2(new_n1647_), .ZN(new_n1649_));
  AOI21_X1   g01583(.A1(new_n1649_), .A2(new_n1639_), .B(new_n1636_), .ZN(new_n1650_));
  OAI21_X1   g01584(.A1(new_n1427_), .A2(new_n1428_), .B(new_n1379_), .ZN(new_n1651_));
  OAI21_X1   g01585(.A1(new_n1343_), .A2(new_n1347_), .B(new_n1334_), .ZN(new_n1652_));
  OR2_X2     g01586(.A1(new_n993_), .A2(new_n990_), .Z(new_n1653_));
  NAND2_X1   g01587(.A1(new_n981_), .A2(new_n1653_), .ZN(new_n1654_));
  XOR2_X1    g01588(.A1(new_n989_), .A2(new_n71_), .Z(new_n1655_));
  OAI21_X1   g01589(.A1(new_n981_), .A2(new_n1655_), .B(new_n1654_), .ZN(new_n1656_));
  NAND3_X1   g01590(.A1(new_n1656_), .A2(new_n1652_), .A3(new_n189_), .ZN(new_n1657_));
  AOI21_X1   g01591(.A1(new_n1354_), .A2(new_n1355_), .B(new_n1353_), .ZN(new_n1658_));
  NOR2_X1    g01592(.A1(new_n981_), .A2(new_n1655_), .ZN(new_n1659_));
  AOI21_X1   g01593(.A1(new_n981_), .A2(new_n1653_), .B(new_n1659_), .ZN(new_n1660_));
  OAI21_X1   g01594(.A1(new_n1660_), .A2(new_n248_), .B(new_n1658_), .ZN(new_n1661_));
  AOI21_X1   g01595(.A1(new_n1661_), .A2(new_n1657_), .B(new_n1368_), .ZN(new_n1662_));
  NOR3_X1    g01596(.A1(new_n1660_), .A2(new_n1658_), .A3(new_n248_), .ZN(new_n1663_));
  AOI21_X1   g01597(.A1(new_n1656_), .A2(new_n189_), .B(new_n1652_), .ZN(new_n1664_));
  NOR3_X1    g01598(.A1(new_n1664_), .A2(new_n1663_), .A3(new_n1375_), .ZN(new_n1665_));
  OAI21_X1   g01599(.A1(new_n1665_), .A2(new_n1662_), .B(new_n356_), .ZN(new_n1666_));
  OAI21_X1   g01600(.A1(new_n1664_), .A2(new_n1663_), .B(new_n1375_), .ZN(new_n1667_));
  NAND3_X1   g01601(.A1(new_n1661_), .A2(new_n1657_), .A3(new_n1368_), .ZN(new_n1668_));
  NAND3_X1   g01602(.A1(new_n1667_), .A2(new_n1668_), .A3(new_n273_), .ZN(new_n1669_));
  AOI22_X1   g01603(.A1(new_n1666_), .A2(new_n1669_), .B1(new_n1382_), .B2(new_n1651_), .ZN(new_n1670_));
  INV_X1     g01604(.I(new_n1670_), .ZN(new_n1671_));
  NAND3_X1   g01605(.A1(new_n1667_), .A2(new_n1668_), .A3(new_n356_), .ZN(new_n1672_));
  OAI21_X1   g01606(.A1(new_n1665_), .A2(new_n1662_), .B(new_n273_), .ZN(new_n1673_));
  NAND2_X1   g01607(.A1(new_n1673_), .A2(new_n1672_), .ZN(new_n1674_));
  NAND3_X1   g01608(.A1(new_n1674_), .A2(new_n1382_), .A3(new_n1651_), .ZN(new_n1675_));
  AOI21_X1   g01609(.A1(new_n1675_), .A2(new_n1671_), .B(new_n568_), .ZN(new_n1676_));
  OAI21_X1   g01610(.A1(new_n1615_), .A2(new_n1650_), .B(new_n1676_), .ZN(new_n1677_));
  NOR3_X1    g01611(.A1(new_n1676_), .A2(new_n1650_), .A3(new_n1615_), .ZN(new_n1678_));
  INV_X1     g01612(.I(new_n1678_), .ZN(new_n1679_));
  AOI21_X1   g01613(.A1(new_n1679_), .A2(new_n1677_), .B(new_n1433_), .ZN(new_n1680_));
  NOR2_X1    g01614(.A1(new_n1650_), .A2(new_n1615_), .ZN(new_n1681_));
  INV_X1     g01615(.I(new_n1676_), .ZN(new_n1682_));
  NOR2_X1    g01616(.A1(new_n1681_), .A2(new_n1682_), .ZN(new_n1683_));
  NOR3_X1    g01617(.A1(new_n1683_), .A2(new_n1647_), .A3(new_n1678_), .ZN(new_n1684_));
  NOR2_X1    g01618(.A1(new_n1680_), .A2(new_n1684_), .ZN(new_n1685_));
  INV_X1     g01619(.I(new_n1613_), .ZN(new_n1686_));
  NAND2_X1   g01620(.A1(new_n1686_), .A2(new_n568_), .ZN(new_n1687_));
  AOI21_X1   g01621(.A1(new_n1611_), .A2(new_n1440_), .B(new_n1687_), .ZN(new_n1688_));
  AOI21_X1   g01622(.A1(new_n1633_), .A2(new_n1634_), .B(\a[17] ), .ZN(new_n1689_));
  NOR3_X1    g01623(.A1(new_n1631_), .A2(new_n1627_), .A3(new_n126_), .ZN(new_n1690_));
  NOR2_X1    g01624(.A1(new_n1690_), .A2(new_n1689_), .ZN(new_n1691_));
  NOR3_X1    g01625(.A1(new_n1691_), .A2(new_n1688_), .A3(new_n1561_), .ZN(new_n1692_));
  NOR2_X1    g01626(.A1(new_n1615_), .A2(new_n1636_), .ZN(new_n1693_));
  NOR2_X1    g01627(.A1(new_n1693_), .A2(new_n1692_), .ZN(new_n1694_));
  NAND2_X1   g01628(.A1(new_n1624_), .A2(new_n1626_), .ZN(new_n1695_));
  NAND2_X1   g01629(.A1(new_n1638_), .A2(new_n1637_), .ZN(new_n1696_));
  NAND2_X1   g01630(.A1(new_n1696_), .A2(new_n1695_), .ZN(new_n1697_));
  NAND3_X1   g01631(.A1(new_n1648_), .A2(new_n1647_), .A3(new_n1697_), .ZN(new_n1698_));
  NAND3_X1   g01632(.A1(new_n1698_), .A2(new_n1615_), .A3(new_n1636_), .ZN(new_n1699_));
  AOI21_X1   g01633(.A1(new_n1646_), .A2(new_n1642_), .B(new_n443_), .ZN(new_n1700_));
  NOR3_X1    g01634(.A1(new_n1433_), .A2(new_n1700_), .A3(new_n1639_), .ZN(new_n1701_));
  OAI22_X1   g01635(.A1(new_n1701_), .A2(new_n1691_), .B1(new_n1561_), .B2(new_n1688_), .ZN(new_n1702_));
  NAND2_X1   g01636(.A1(new_n1702_), .A2(new_n1699_), .ZN(new_n1703_));
  INV_X1     g01637(.I(new_n1703_), .ZN(new_n1704_));
  OAI21_X1   g01638(.A1(new_n1704_), .A2(new_n1694_), .B(new_n644_), .ZN(new_n1705_));
  NOR2_X1    g01639(.A1(new_n1440_), .A2(new_n443_), .ZN(new_n1706_));
  NAND2_X1   g01640(.A1(new_n1706_), .A2(new_n1611_), .ZN(new_n1707_));
  NOR3_X1    g01641(.A1(new_n1560_), .A2(new_n1456_), .A3(new_n1555_), .ZN(new_n1708_));
  OAI21_X1   g01642(.A1(new_n1437_), .A2(new_n1438_), .B(new_n1423_), .ZN(new_n1709_));
  NAND3_X1   g01643(.A1(new_n1435_), .A2(new_n1324_), .A3(new_n1434_), .ZN(new_n1710_));
  NAND2_X1   g01644(.A1(new_n1710_), .A2(new_n1709_), .ZN(new_n1711_));
  NAND2_X1   g01645(.A1(new_n1711_), .A2(new_n568_), .ZN(new_n1712_));
  NAND2_X1   g01646(.A1(new_n1712_), .A2(new_n1708_), .ZN(new_n1713_));
  AOI21_X1   g01647(.A1(new_n1713_), .A2(new_n1707_), .B(new_n1686_), .ZN(new_n1714_));
  NOR2_X1    g01648(.A1(new_n1712_), .A2(new_n1708_), .ZN(new_n1715_));
  NOR2_X1    g01649(.A1(new_n1706_), .A2(new_n1611_), .ZN(new_n1716_));
  NOR3_X1    g01650(.A1(new_n1715_), .A2(new_n1716_), .A3(new_n1613_), .ZN(new_n1717_));
  NAND2_X1   g01651(.A1(new_n1494_), .A2(new_n1484_), .ZN(new_n1718_));
  NOR2_X1    g01652(.A1(new_n1718_), .A2(new_n568_), .ZN(new_n1719_));
  NAND3_X1   g01653(.A1(new_n1577_), .A2(new_n1466_), .A3(new_n443_), .ZN(new_n1720_));
  OAI21_X1   g01654(.A1(new_n568_), .A2(new_n1572_), .B(new_n1497_), .ZN(new_n1721_));
  AOI21_X1   g01655(.A1(new_n1721_), .A2(new_n1720_), .B(new_n1719_), .ZN(new_n1722_));
  INV_X1     g01656(.I(new_n1719_), .ZN(new_n1723_));
  NOR3_X1    g01657(.A1(new_n1497_), .A2(new_n1572_), .A3(new_n568_), .ZN(new_n1724_));
  AOI21_X1   g01658(.A1(new_n443_), .A2(new_n1466_), .B(new_n1577_), .ZN(new_n1725_));
  NOR3_X1    g01659(.A1(new_n1725_), .A2(new_n1724_), .A3(new_n1723_), .ZN(new_n1726_));
  NOR2_X1    g01660(.A1(new_n1722_), .A2(new_n1726_), .ZN(new_n1727_));
  NAND3_X1   g01661(.A1(new_n1478_), .A2(new_n443_), .A3(new_n1472_), .ZN(new_n1728_));
  OAI21_X1   g01662(.A1(new_n1475_), .A2(new_n1473_), .B(new_n568_), .ZN(new_n1729_));
  AOI21_X1   g01663(.A1(new_n1729_), .A2(new_n1728_), .B(new_n1470_), .ZN(new_n1730_));
  AOI21_X1   g01664(.A1(new_n1476_), .A2(new_n1479_), .B(new_n1471_), .ZN(new_n1731_));
  NOR2_X1    g01665(.A1(new_n1731_), .A2(new_n1730_), .ZN(new_n1732_));
  XNOR2_X1   g01666(.A1(\a[11] ), .A2(\a[12] ), .ZN(new_n1733_));
  NAND2_X1   g01667(.A1(new_n1733_), .A2(\a[14] ), .ZN(new_n1734_));
  AOI21_X1   g01668(.A1(new_n644_), .A2(new_n1734_), .B(new_n1468_), .ZN(new_n1735_));
  NAND2_X1   g01669(.A1(new_n443_), .A2(new_n1469_), .ZN(new_n1736_));
  NAND3_X1   g01670(.A1(new_n1620_), .A2(\a[17] ), .A3(new_n1468_), .ZN(new_n1737_));
  AOI21_X1   g01671(.A1(new_n1736_), .A2(new_n1737_), .B(new_n786_), .ZN(new_n1738_));
  NOR2_X1    g01672(.A1(new_n1738_), .A2(new_n1735_), .ZN(new_n1739_));
  NAND3_X1   g01673(.A1(new_n1736_), .A2(new_n786_), .A3(new_n1737_), .ZN(new_n1740_));
  INV_X1     g01674(.I(new_n1740_), .ZN(new_n1741_));
  NAND3_X1   g01675(.A1(new_n786_), .A2(new_n443_), .A3(new_n1469_), .ZN(new_n1742_));
  NAND2_X1   g01676(.A1(new_n443_), .A2(new_n1469_), .ZN(new_n1743_));
  NAND2_X1   g01677(.A1(new_n1743_), .A2(new_n644_), .ZN(new_n1744_));
  NOR3_X1    g01678(.A1(new_n568_), .A2(new_n1467_), .A3(new_n1469_), .ZN(new_n1745_));
  NAND2_X1   g01679(.A1(new_n443_), .A2(new_n1467_), .ZN(new_n1746_));
  XOR2_X1    g01680(.A1(\a[14] ), .A2(\a[15] ), .Z(new_n1747_));
  NOR2_X1    g01681(.A1(new_n1747_), .A2(new_n126_), .ZN(new_n1748_));
  NAND2_X1   g01682(.A1(new_n568_), .A2(new_n1229_), .ZN(new_n1749_));
  AOI22_X1   g01683(.A1(new_n1749_), .A2(new_n1746_), .B1(new_n443_), .B2(new_n1748_), .ZN(new_n1750_));
  NOR3_X1    g01684(.A1(new_n1750_), .A2(new_n644_), .A3(new_n1745_), .ZN(new_n1751_));
  INV_X1     g01685(.I(new_n1745_), .ZN(new_n1752_));
  INV_X1     g01686(.I(new_n1746_), .ZN(new_n1753_));
  NAND2_X1   g01687(.A1(new_n443_), .A2(new_n1748_), .ZN(new_n1754_));
  NOR2_X1    g01688(.A1(new_n443_), .A2(new_n1467_), .ZN(new_n1755_));
  OAI21_X1   g01689(.A1(new_n1753_), .A2(new_n1755_), .B(new_n1754_), .ZN(new_n1756_));
  AOI21_X1   g01690(.A1(new_n1756_), .A2(new_n1752_), .B(new_n786_), .ZN(new_n1757_));
  NAND2_X1   g01691(.A1(new_n1744_), .A2(new_n1742_), .ZN(new_n1759_));
  OAI21_X1   g01692(.A1(new_n1739_), .A2(new_n1741_), .B(new_n1759_), .ZN(new_n1760_));
  NOR2_X1    g01693(.A1(new_n1732_), .A2(new_n1760_), .ZN(new_n1761_));
  NAND3_X1   g01694(.A1(new_n1756_), .A2(new_n1752_), .A3(new_n644_), .ZN(new_n1762_));
  AOI21_X1   g01695(.A1(new_n1732_), .A2(new_n1760_), .B(new_n1762_), .ZN(new_n1763_));
  NOR2_X1    g01696(.A1(new_n1576_), .A2(new_n1481_), .ZN(new_n1764_));
  NOR3_X1    g01697(.A1(new_n1574_), .A2(new_n1764_), .A3(new_n1575_), .ZN(new_n1765_));
  NAND2_X1   g01698(.A1(new_n1482_), .A2(new_n1483_), .ZN(new_n1766_));
  AOI21_X1   g01699(.A1(new_n1477_), .A2(new_n1479_), .B(new_n1766_), .ZN(new_n1767_));
  OAI21_X1   g01700(.A1(new_n1767_), .A2(new_n1765_), .B(new_n644_), .ZN(new_n1768_));
  OAI21_X1   g01701(.A1(new_n1763_), .A2(new_n1761_), .B(new_n1768_), .ZN(new_n1769_));
  NAND3_X1   g01702(.A1(new_n1477_), .A2(new_n1479_), .A3(new_n1766_), .ZN(new_n1770_));
  OAI21_X1   g01703(.A1(new_n1574_), .A2(new_n1575_), .B(new_n1764_), .ZN(new_n1771_));
  NAND3_X1   g01704(.A1(new_n1770_), .A2(new_n1771_), .A3(new_n786_), .ZN(new_n1772_));
  NOR2_X1    g01705(.A1(new_n1574_), .A2(new_n1575_), .ZN(new_n1773_));
  NAND3_X1   g01706(.A1(new_n1494_), .A2(new_n568_), .A3(new_n1484_), .ZN(new_n1774_));
  OAI21_X1   g01707(.A1(new_n1490_), .A2(new_n1485_), .B(new_n443_), .ZN(new_n1775_));
  NAND3_X1   g01708(.A1(new_n1775_), .A2(new_n1774_), .A3(new_n1482_), .ZN(new_n1776_));
  NAND3_X1   g01709(.A1(new_n1776_), .A2(new_n1773_), .A3(new_n1766_), .ZN(new_n1777_));
  NAND2_X1   g01710(.A1(new_n1477_), .A2(new_n1479_), .ZN(new_n1778_));
  NOR3_X1    g01711(.A1(new_n1491_), .A2(new_n1495_), .A3(new_n1481_), .ZN(new_n1779_));
  OAI21_X1   g01712(.A1(new_n1779_), .A2(new_n1764_), .B(new_n1778_), .ZN(new_n1780_));
  NAND3_X1   g01713(.A1(new_n1780_), .A2(new_n1777_), .A3(new_n786_), .ZN(new_n1781_));
  NOR3_X1    g01714(.A1(new_n1779_), .A2(new_n1778_), .A3(new_n1764_), .ZN(new_n1782_));
  AOI21_X1   g01715(.A1(new_n1776_), .A2(new_n1766_), .B(new_n1773_), .ZN(new_n1783_));
  OAI21_X1   g01716(.A1(new_n1782_), .A2(new_n1783_), .B(new_n644_), .ZN(new_n1784_));
  NAND4_X1   g01717(.A1(new_n1769_), .A2(new_n1784_), .A3(new_n1781_), .A4(new_n1772_), .ZN(new_n1785_));
  NOR2_X1    g01718(.A1(new_n1785_), .A2(new_n1727_), .ZN(new_n1786_));
  AOI21_X1   g01719(.A1(new_n1780_), .A2(new_n1777_), .B(new_n786_), .ZN(new_n1787_));
  NAND2_X1   g01720(.A1(new_n1787_), .A2(new_n786_), .ZN(new_n1788_));
  AOI21_X1   g01721(.A1(new_n1785_), .A2(new_n1727_), .B(new_n1788_), .ZN(new_n1789_));
  NOR2_X1    g01722(.A1(new_n1789_), .A2(new_n1786_), .ZN(new_n1790_));
  NOR2_X1    g01723(.A1(new_n1579_), .A2(new_n1578_), .ZN(new_n1791_));
  AOI21_X1   g01724(.A1(new_n1582_), .A2(new_n1510_), .B(new_n1791_), .ZN(new_n1792_));
  XOR2_X1    g01725(.A1(new_n1508_), .A2(new_n443_), .Z(new_n1793_));
  AOI21_X1   g01726(.A1(new_n1791_), .A2(new_n1793_), .B(new_n1792_), .ZN(new_n1794_));
  NOR2_X1    g01727(.A1(new_n1790_), .A2(new_n1794_), .ZN(new_n1795_));
  AOI21_X1   g01728(.A1(new_n1790_), .A2(new_n1794_), .B(new_n279_), .ZN(new_n1796_));
  AOI22_X1   g01729(.A1(new_n1524_), .A2(new_n1584_), .B1(new_n1583_), .B2(new_n1510_), .ZN(new_n1797_));
  NOR2_X1    g01730(.A1(new_n1522_), .A2(new_n1797_), .ZN(new_n1798_));
  NAND2_X1   g01731(.A1(new_n1798_), .A2(new_n644_), .ZN(new_n1799_));
  OAI21_X1   g01732(.A1(new_n1796_), .A2(new_n1795_), .B(new_n1799_), .ZN(new_n1800_));
  NOR2_X1    g01733(.A1(new_n1798_), .A2(new_n644_), .ZN(new_n1801_));
  INV_X1     g01734(.I(new_n1801_), .ZN(new_n1802_));
  OAI21_X1   g01735(.A1(new_n1566_), .A2(new_n1564_), .B(new_n568_), .ZN(new_n1803_));
  NOR2_X1    g01736(.A1(new_n1522_), .A2(new_n1803_), .ZN(new_n1804_));
  AOI21_X1   g01737(.A1(new_n568_), .A2(new_n1461_), .B(new_n1585_), .ZN(new_n1805_));
  OAI21_X1   g01738(.A1(new_n1805_), .A2(new_n1804_), .B(new_n1524_), .ZN(new_n1806_));
  NAND3_X1   g01739(.A1(new_n1461_), .A2(new_n1585_), .A3(new_n568_), .ZN(new_n1807_));
  NAND2_X1   g01740(.A1(new_n1522_), .A2(new_n1803_), .ZN(new_n1808_));
  NAND3_X1   g01741(.A1(new_n1807_), .A2(new_n1808_), .A3(new_n1521_), .ZN(new_n1809_));
  AOI21_X1   g01742(.A1(new_n1806_), .A2(new_n1809_), .B(new_n644_), .ZN(new_n1810_));
  AOI21_X1   g01743(.A1(new_n1800_), .A2(new_n1802_), .B(new_n1810_), .ZN(new_n1811_));
  NAND2_X1   g01744(.A1(new_n1806_), .A2(new_n1809_), .ZN(new_n1812_));
  NOR2_X1    g01745(.A1(new_n1812_), .A2(new_n786_), .ZN(new_n1813_));
  NOR2_X1    g01746(.A1(new_n1588_), .A2(new_n1586_), .ZN(new_n1814_));
  NAND2_X1   g01747(.A1(new_n1594_), .A2(new_n443_), .ZN(new_n1815_));
  NAND2_X1   g01748(.A1(new_n1533_), .A2(new_n568_), .ZN(new_n1816_));
  AOI21_X1   g01749(.A1(new_n1815_), .A2(new_n1816_), .B(new_n1814_), .ZN(new_n1817_));
  OAI21_X1   g01750(.A1(new_n1531_), .A2(new_n1534_), .B(new_n1814_), .ZN(new_n1818_));
  INV_X1     g01751(.I(new_n1818_), .ZN(new_n1819_));
  OAI21_X1   g01752(.A1(new_n1819_), .A2(new_n1817_), .B(new_n644_), .ZN(new_n1820_));
  OAI21_X1   g01753(.A1(new_n1811_), .A2(new_n1813_), .B(new_n1820_), .ZN(new_n1821_));
  INV_X1     g01754(.I(new_n1814_), .ZN(new_n1822_));
  NAND2_X1   g01755(.A1(new_n1815_), .A2(new_n1816_), .ZN(new_n1823_));
  NAND2_X1   g01756(.A1(new_n1822_), .A2(new_n1823_), .ZN(new_n1824_));
  NAND2_X1   g01757(.A1(new_n1824_), .A2(new_n1818_), .ZN(new_n1825_));
  NOR2_X1    g01758(.A1(new_n1825_), .A2(new_n644_), .ZN(new_n1826_));
  INV_X1     g01759(.I(new_n1826_), .ZN(new_n1827_));
  NAND2_X1   g01760(.A1(new_n1593_), .A2(new_n1595_), .ZN(new_n1828_));
  NAND2_X1   g01761(.A1(new_n1540_), .A2(new_n443_), .ZN(new_n1829_));
  NAND2_X1   g01762(.A1(new_n1599_), .A2(new_n568_), .ZN(new_n1830_));
  NAND2_X1   g01763(.A1(new_n1829_), .A2(new_n1830_), .ZN(new_n1831_));
  NAND2_X1   g01764(.A1(new_n1831_), .A2(new_n1828_), .ZN(new_n1832_));
  NOR2_X1    g01765(.A1(new_n1532_), .A2(new_n1534_), .ZN(new_n1833_));
  OAI21_X1   g01766(.A1(new_n1597_), .A2(new_n1600_), .B(new_n1833_), .ZN(new_n1834_));
  AOI21_X1   g01767(.A1(new_n1832_), .A2(new_n1834_), .B(new_n786_), .ZN(new_n1835_));
  AOI21_X1   g01768(.A1(new_n1821_), .A2(new_n1827_), .B(new_n1835_), .ZN(new_n1836_));
  AOI21_X1   g01769(.A1(new_n1829_), .A2(new_n1830_), .B(new_n1833_), .ZN(new_n1837_));
  AOI21_X1   g01770(.A1(new_n1538_), .A2(new_n1541_), .B(new_n1828_), .ZN(new_n1838_));
  NOR3_X1    g01771(.A1(new_n1837_), .A2(new_n1838_), .A3(new_n644_), .ZN(new_n1839_));
  NAND2_X1   g01772(.A1(new_n1604_), .A2(new_n568_), .ZN(new_n1840_));
  NAND2_X1   g01773(.A1(new_n1552_), .A2(new_n443_), .ZN(new_n1841_));
  AOI21_X1   g01774(.A1(new_n1840_), .A2(new_n1841_), .B(new_n1601_), .ZN(new_n1842_));
  INV_X1     g01775(.I(new_n1601_), .ZN(new_n1843_));
  NOR2_X1    g01776(.A1(new_n1605_), .A2(new_n1554_), .ZN(new_n1844_));
  NOR2_X1    g01777(.A1(new_n1844_), .A2(new_n1843_), .ZN(new_n1845_));
  OAI21_X1   g01778(.A1(new_n1845_), .A2(new_n1842_), .B(new_n644_), .ZN(new_n1846_));
  OAI21_X1   g01779(.A1(new_n1836_), .A2(new_n1839_), .B(new_n1846_), .ZN(new_n1847_));
  NOR3_X1    g01780(.A1(new_n1845_), .A2(new_n644_), .A3(new_n1842_), .ZN(new_n1848_));
  INV_X1     g01781(.I(new_n1848_), .ZN(new_n1849_));
  NOR2_X1    g01782(.A1(new_n639_), .A2(\a[12] ), .ZN(new_n1850_));
  AOI21_X1   g01783(.A1(\a[12] ), .A2(new_n783_), .B(new_n1850_), .ZN(new_n1851_));
  NOR2_X1    g01784(.A1(new_n1851_), .A2(new_n643_), .ZN(new_n1852_));
  XOR2_X1    g01785(.A1(new_n1852_), .A2(new_n279_), .Z(new_n1853_));
  INV_X1     g01786(.I(new_n1853_), .ZN(new_n1854_));
  OAI22_X1   g01787(.A1(new_n1598_), .A2(new_n1600_), .B1(new_n1604_), .B2(new_n443_), .ZN(new_n1855_));
  OAI21_X1   g01788(.A1(new_n1444_), .A2(new_n1446_), .B(new_n443_), .ZN(new_n1856_));
  NAND3_X1   g01789(.A1(new_n1418_), .A2(new_n1445_), .A3(new_n1403_), .ZN(new_n1857_));
  NAND2_X1   g01790(.A1(new_n1442_), .A2(new_n1443_), .ZN(new_n1858_));
  NAND3_X1   g01791(.A1(new_n1858_), .A2(new_n1857_), .A3(new_n568_), .ZN(new_n1859_));
  AOI22_X1   g01792(.A1(new_n1855_), .A2(new_n1606_), .B1(new_n1856_), .B2(new_n1859_), .ZN(new_n1860_));
  NOR3_X1    g01793(.A1(new_n1444_), .A2(new_n1446_), .A3(new_n568_), .ZN(new_n1861_));
  AOI21_X1   g01794(.A1(new_n1858_), .A2(new_n1857_), .B(new_n443_), .ZN(new_n1862_));
  NOR2_X1    g01795(.A1(new_n1861_), .A2(new_n1862_), .ZN(new_n1863_));
  NOR2_X1    g01796(.A1(new_n1607_), .A2(new_n1863_), .ZN(new_n1864_));
  NOR3_X1    g01797(.A1(new_n1864_), .A2(new_n1854_), .A3(new_n1860_), .ZN(new_n1865_));
  AOI21_X1   g01798(.A1(new_n1858_), .A2(new_n1857_), .B(new_n568_), .ZN(new_n1866_));
  NOR3_X1    g01799(.A1(new_n1444_), .A2(new_n1446_), .A3(new_n443_), .ZN(new_n1867_));
  OAI22_X1   g01800(.A1(new_n1553_), .A2(new_n1554_), .B1(new_n1866_), .B2(new_n1867_), .ZN(new_n1868_));
  NAND3_X1   g01801(.A1(new_n1858_), .A2(new_n1857_), .A3(new_n443_), .ZN(new_n1869_));
  OAI21_X1   g01802(.A1(new_n1444_), .A2(new_n1446_), .B(new_n568_), .ZN(new_n1870_));
  NAND2_X1   g01803(.A1(new_n1870_), .A2(new_n1869_), .ZN(new_n1871_));
  NAND3_X1   g01804(.A1(new_n1871_), .A2(new_n1855_), .A3(new_n1606_), .ZN(new_n1872_));
  AOI21_X1   g01805(.A1(new_n1872_), .A2(new_n1868_), .B(new_n1853_), .ZN(new_n1873_));
  MUX2_X1    g01806(.I0(new_n1448_), .I1(new_n568_), .S(new_n1562_), .Z(new_n1874_));
  NAND2_X1   g01807(.A1(new_n1874_), .A2(new_n1555_), .ZN(new_n1875_));
  MUX2_X1    g01808(.I0(new_n1447_), .I1(new_n443_), .S(new_n1562_), .Z(new_n1876_));
  NAND2_X1   g01809(.A1(new_n1876_), .A2(new_n1607_), .ZN(new_n1877_));
  AOI21_X1   g01810(.A1(new_n1875_), .A2(new_n1877_), .B(new_n786_), .ZN(new_n1878_));
  NOR2_X1    g01811(.A1(new_n1876_), .A2(new_n1607_), .ZN(new_n1879_));
  NOR2_X1    g01812(.A1(new_n1874_), .A2(new_n1555_), .ZN(new_n1880_));
  NOR3_X1    g01813(.A1(new_n1879_), .A2(new_n1880_), .A3(new_n644_), .ZN(new_n1881_));
  NOR2_X1    g01814(.A1(new_n1865_), .A2(new_n1873_), .ZN(new_n1883_));
  AOI21_X1   g01815(.A1(new_n1847_), .A2(new_n1849_), .B(new_n1883_), .ZN(new_n1884_));
  OAI21_X1   g01816(.A1(new_n1714_), .A2(new_n1717_), .B(new_n1884_), .ZN(new_n1885_));
  NOR3_X1    g01817(.A1(new_n1884_), .A2(new_n1714_), .A3(new_n1717_), .ZN(new_n1886_));
  OAI21_X1   g01818(.A1(new_n1879_), .A2(new_n1880_), .B(new_n644_), .ZN(new_n1887_));
  NOR2_X1    g01819(.A1(new_n1887_), .A2(new_n786_), .ZN(new_n1888_));
  INV_X1     g01820(.I(new_n1888_), .ZN(new_n1889_));
  OAI21_X1   g01821(.A1(new_n1886_), .A2(new_n1889_), .B(new_n1885_), .ZN(new_n1890_));
  NAND3_X1   g01822(.A1(new_n1702_), .A2(new_n1699_), .A3(new_n786_), .ZN(new_n1891_));
  AOI21_X1   g01823(.A1(new_n1702_), .A2(new_n1699_), .B(new_n786_), .ZN(new_n1892_));
  INV_X1     g01824(.I(new_n1892_), .ZN(new_n1893_));
  NAND3_X1   g01825(.A1(new_n1893_), .A2(new_n1694_), .A3(new_n1891_), .ZN(new_n1894_));
  NAND3_X1   g01826(.A1(new_n1894_), .A2(new_n1705_), .A3(new_n1890_), .ZN(new_n1895_));
  NOR2_X1    g01827(.A1(new_n1895_), .A2(new_n1685_), .ZN(new_n1896_));
  NAND2_X1   g01828(.A1(new_n1892_), .A2(new_n786_), .ZN(new_n1897_));
  AOI21_X1   g01829(.A1(new_n1895_), .A2(new_n1685_), .B(new_n1897_), .ZN(new_n1898_));
  NAND2_X1   g01830(.A1(new_n1671_), .A2(new_n1675_), .ZN(new_n1899_));
  NAND2_X1   g01831(.A1(new_n1681_), .A2(new_n1899_), .ZN(new_n1900_));
  NOR2_X1    g01832(.A1(new_n1647_), .A2(new_n568_), .ZN(new_n1901_));
  OAI21_X1   g01833(.A1(new_n1681_), .A2(new_n1899_), .B(new_n1901_), .ZN(new_n1902_));
  NAND2_X1   g01834(.A1(new_n1651_), .A2(new_n1382_), .ZN(new_n1903_));
  NAND2_X1   g01835(.A1(new_n1903_), .A2(new_n1666_), .ZN(new_n1904_));
  NAND2_X1   g01836(.A1(new_n1904_), .A2(new_n1669_), .ZN(new_n1905_));
  NAND2_X1   g01837(.A1(new_n1656_), .A2(new_n1658_), .ZN(new_n1906_));
  NOR2_X1    g01838(.A1(new_n1375_), .A2(new_n248_), .ZN(new_n1907_));
  OAI21_X1   g01839(.A1(new_n1656_), .A2(new_n1658_), .B(new_n1907_), .ZN(new_n1908_));
  NAND2_X1   g01840(.A1(new_n1908_), .A2(new_n1906_), .ZN(new_n1909_));
  NOR2_X1    g01841(.A1(new_n1000_), .A2(new_n998_), .ZN(new_n1910_));
  NOR2_X1    g01842(.A1(new_n994_), .A2(new_n1910_), .ZN(new_n1911_));
  INV_X1     g01843(.I(new_n1911_), .ZN(new_n1912_));
  XOR2_X1    g01844(.A1(new_n997_), .A2(new_n71_), .Z(new_n1913_));
  INV_X1     g01845(.I(new_n1913_), .ZN(new_n1914_));
  NAND2_X1   g01846(.A1(new_n994_), .A2(new_n1914_), .ZN(new_n1915_));
  AOI21_X1   g01847(.A1(new_n1912_), .A2(new_n1915_), .B(new_n248_), .ZN(new_n1916_));
  NAND3_X1   g01848(.A1(new_n1912_), .A2(new_n248_), .A3(new_n1915_), .ZN(new_n1917_));
  INV_X1     g01849(.I(new_n1917_), .ZN(new_n1918_));
  OAI21_X1   g01850(.A1(new_n1918_), .A2(new_n1916_), .B(new_n1909_), .ZN(new_n1919_));
  INV_X1     g01851(.I(new_n1919_), .ZN(new_n1920_));
  NAND3_X1   g01852(.A1(new_n1912_), .A2(new_n189_), .A3(new_n1915_), .ZN(new_n1921_));
  AOI21_X1   g01853(.A1(new_n1912_), .A2(new_n1915_), .B(new_n189_), .ZN(new_n1922_));
  INV_X1     g01854(.I(new_n1922_), .ZN(new_n1923_));
  AOI21_X1   g01855(.A1(new_n1923_), .A2(new_n1921_), .B(new_n1909_), .ZN(new_n1924_));
  OAI21_X1   g01856(.A1(new_n1920_), .A2(new_n1924_), .B(new_n356_), .ZN(new_n1925_));
  NOR2_X1    g01857(.A1(new_n1660_), .A2(new_n1652_), .ZN(new_n1926_));
  NAND2_X1   g01858(.A1(new_n1660_), .A2(new_n1652_), .ZN(new_n1927_));
  AOI21_X1   g01859(.A1(new_n1927_), .A2(new_n1907_), .B(new_n1926_), .ZN(new_n1928_));
  INV_X1     g01860(.I(new_n1921_), .ZN(new_n1929_));
  OAI21_X1   g01861(.A1(new_n1929_), .A2(new_n1922_), .B(new_n1928_), .ZN(new_n1930_));
  NAND3_X1   g01862(.A1(new_n1930_), .A2(new_n1919_), .A3(new_n273_), .ZN(new_n1931_));
  NAND2_X1   g01863(.A1(new_n1925_), .A2(new_n1931_), .ZN(new_n1932_));
  NAND2_X1   g01864(.A1(new_n1932_), .A2(new_n1905_), .ZN(new_n1933_));
  INV_X1     g01865(.I(new_n1669_), .ZN(new_n1934_));
  AOI21_X1   g01866(.A1(new_n1903_), .A2(new_n1666_), .B(new_n1934_), .ZN(new_n1935_));
  NOR3_X1    g01867(.A1(new_n1920_), .A2(new_n1924_), .A3(new_n273_), .ZN(new_n1936_));
  AOI21_X1   g01868(.A1(new_n1930_), .A2(new_n1919_), .B(new_n356_), .ZN(new_n1937_));
  OAI21_X1   g01869(.A1(new_n1936_), .A2(new_n1937_), .B(new_n1935_), .ZN(new_n1938_));
  AOI21_X1   g01870(.A1(new_n1933_), .A2(new_n1938_), .B(new_n568_), .ZN(new_n1939_));
  AOI21_X1   g01871(.A1(new_n1925_), .A2(new_n1931_), .B(new_n1935_), .ZN(new_n1940_));
  NOR2_X1    g01872(.A1(new_n1936_), .A2(new_n1937_), .ZN(new_n1941_));
  NOR2_X1    g01873(.A1(new_n1941_), .A2(new_n1905_), .ZN(new_n1942_));
  NOR3_X1    g01874(.A1(new_n1942_), .A2(new_n1940_), .A3(new_n443_), .ZN(new_n1943_));
  NOR2_X1    g01875(.A1(new_n1939_), .A2(new_n1943_), .ZN(new_n1944_));
  AOI21_X1   g01876(.A1(new_n1900_), .A2(new_n1902_), .B(new_n1944_), .ZN(new_n1945_));
  NAND3_X1   g01877(.A1(new_n1933_), .A2(new_n1938_), .A3(new_n443_), .ZN(new_n1946_));
  OAI21_X1   g01878(.A1(new_n1942_), .A2(new_n1940_), .B(new_n568_), .ZN(new_n1947_));
  NAND2_X1   g01879(.A1(new_n1947_), .A2(new_n1946_), .ZN(new_n1948_));
  NAND3_X1   g01880(.A1(new_n1948_), .A2(new_n1900_), .A3(new_n1902_), .ZN(new_n1949_));
  INV_X1     g01881(.I(new_n1949_), .ZN(new_n1950_));
  OAI21_X1   g01882(.A1(new_n1950_), .A2(new_n1945_), .B(new_n644_), .ZN(new_n1951_));
  OAI21_X1   g01883(.A1(new_n1898_), .A2(new_n1896_), .B(new_n1951_), .ZN(new_n1952_));
  NAND2_X1   g01884(.A1(new_n1902_), .A2(new_n1900_), .ZN(new_n1953_));
  INV_X1     g01885(.I(new_n1944_), .ZN(new_n1954_));
  NAND2_X1   g01886(.A1(new_n1954_), .A2(new_n1953_), .ZN(new_n1955_));
  NAND3_X1   g01887(.A1(new_n1955_), .A2(new_n1949_), .A3(new_n786_), .ZN(new_n1956_));
  INV_X1     g01888(.I(new_n1953_), .ZN(new_n1957_));
  INV_X1     g01889(.I(new_n1947_), .ZN(new_n1958_));
  NAND2_X1   g01890(.A1(new_n1905_), .A2(new_n1925_), .ZN(new_n1959_));
  NOR4_X1    g01891(.A1(new_n981_), .A2(new_n71_), .A3(new_n989_), .A4(new_n997_), .ZN(new_n1960_));
  INV_X1     g01892(.I(new_n1960_), .ZN(new_n1961_));
  NAND4_X1   g01893(.A1(new_n981_), .A2(new_n71_), .A3(new_n989_), .A4(new_n997_), .ZN(new_n1962_));
  AOI21_X1   g01894(.A1(new_n1961_), .A2(new_n1962_), .B(new_n995_), .ZN(new_n1963_));
  INV_X1     g01895(.I(new_n995_), .ZN(new_n1964_));
  AOI21_X1   g01896(.A1(new_n994_), .A2(new_n118_), .B(new_n1964_), .ZN(new_n1965_));
  OAI21_X1   g01897(.A1(new_n1963_), .A2(new_n1965_), .B(new_n1004_), .ZN(new_n1966_));
  INV_X1     g01898(.I(new_n1004_), .ZN(new_n1967_));
  INV_X1     g01899(.I(new_n1962_), .ZN(new_n1968_));
  OAI21_X1   g01900(.A1(new_n1968_), .A2(new_n1960_), .B(new_n1964_), .ZN(new_n1969_));
  INV_X1     g01901(.I(new_n1965_), .ZN(new_n1970_));
  NAND3_X1   g01902(.A1(new_n1969_), .A2(new_n1970_), .A3(new_n1967_), .ZN(new_n1971_));
  NOR2_X1    g01903(.A1(new_n245_), .A2(\a[21] ), .ZN(new_n1972_));
  AOI21_X1   g01904(.A1(\a[21] ), .A2(new_n187_), .B(new_n1972_), .ZN(new_n1973_));
  NOR2_X1    g01905(.A1(new_n1973_), .A2(new_n1239_), .ZN(new_n1974_));
  XOR2_X1    g01906(.A1(new_n1974_), .A2(new_n68_), .Z(new_n1975_));
  AOI21_X1   g01907(.A1(new_n1966_), .A2(new_n1971_), .B(new_n1975_), .ZN(new_n1976_));
  AOI21_X1   g01908(.A1(new_n1969_), .A2(new_n1970_), .B(new_n1967_), .ZN(new_n1977_));
  NOR3_X1    g01909(.A1(new_n1963_), .A2(new_n1004_), .A3(new_n1965_), .ZN(new_n1978_));
  XOR2_X1    g01910(.A1(new_n1974_), .A2(\a[23] ), .Z(new_n1979_));
  NOR3_X1    g01911(.A1(new_n1978_), .A2(new_n1977_), .A3(new_n1979_), .ZN(new_n1980_));
  NOR2_X1    g01912(.A1(new_n1980_), .A2(new_n1976_), .ZN(new_n1981_));
  AOI21_X1   g01913(.A1(new_n1909_), .A2(new_n1921_), .B(new_n1922_), .ZN(new_n1982_));
  INV_X1     g01914(.I(new_n1982_), .ZN(new_n1983_));
  NAND2_X1   g01915(.A1(new_n1981_), .A2(new_n1983_), .ZN(new_n1984_));
  INV_X1     g01916(.I(new_n1975_), .ZN(new_n1985_));
  OAI21_X1   g01917(.A1(new_n1978_), .A2(new_n1977_), .B(new_n1985_), .ZN(new_n1986_));
  INV_X1     g01918(.I(new_n1979_), .ZN(new_n1987_));
  NAND3_X1   g01919(.A1(new_n1966_), .A2(new_n1971_), .A3(new_n1987_), .ZN(new_n1988_));
  NAND2_X1   g01920(.A1(new_n1986_), .A2(new_n1988_), .ZN(new_n1989_));
  NAND2_X1   g01921(.A1(new_n1989_), .A2(new_n1982_), .ZN(new_n1990_));
  NAND3_X1   g01922(.A1(new_n1984_), .A2(new_n1990_), .A3(new_n273_), .ZN(new_n1991_));
  NOR2_X1    g01923(.A1(new_n1989_), .A2(new_n1982_), .ZN(new_n1992_));
  NOR2_X1    g01924(.A1(new_n1981_), .A2(new_n1983_), .ZN(new_n1993_));
  OAI21_X1   g01925(.A1(new_n1993_), .A2(new_n1992_), .B(new_n356_), .ZN(new_n1994_));
  NAND4_X1   g01926(.A1(new_n1959_), .A2(new_n1991_), .A3(new_n1994_), .A4(new_n1931_), .ZN(new_n1995_));
  INV_X1     g01927(.I(new_n1931_), .ZN(new_n1996_));
  NAND2_X1   g01928(.A1(new_n1930_), .A2(new_n1919_), .ZN(new_n1997_));
  AOI22_X1   g01929(.A1(new_n1904_), .A2(new_n1669_), .B1(new_n1997_), .B2(new_n356_), .ZN(new_n1998_));
  NOR3_X1    g01930(.A1(new_n1993_), .A2(new_n1992_), .A3(new_n356_), .ZN(new_n1999_));
  AOI21_X1   g01931(.A1(new_n1984_), .A2(new_n1990_), .B(new_n273_), .ZN(new_n2000_));
  OAI22_X1   g01932(.A1(new_n1999_), .A2(new_n2000_), .B1(new_n1998_), .B2(new_n1996_), .ZN(new_n2001_));
  XOR2_X1    g01933(.A1(new_n1623_), .A2(new_n126_), .Z(new_n2002_));
  AOI21_X1   g01934(.A1(new_n1995_), .A2(new_n2001_), .B(new_n2002_), .ZN(new_n2003_));
  NOR4_X1    g01935(.A1(new_n1998_), .A2(new_n2000_), .A3(new_n1999_), .A4(new_n1996_), .ZN(new_n2004_));
  AOI22_X1   g01936(.A1(new_n1959_), .A2(new_n1931_), .B1(new_n1994_), .B2(new_n1991_), .ZN(new_n2005_));
  XOR2_X1    g01937(.A1(new_n1623_), .A2(\a[17] ), .Z(new_n2006_));
  NOR3_X1    g01938(.A1(new_n2005_), .A2(new_n2004_), .A3(new_n2006_), .ZN(new_n2007_));
  NOR2_X1    g01939(.A1(new_n2007_), .A2(new_n2003_), .ZN(new_n2008_));
  NOR3_X1    g01940(.A1(new_n2008_), .A2(new_n1944_), .A3(new_n1958_), .ZN(new_n2009_));
  NOR2_X1    g01941(.A1(new_n1942_), .A2(new_n1940_), .ZN(new_n2010_));
  NOR2_X1    g01942(.A1(new_n2010_), .A2(new_n443_), .ZN(new_n2011_));
  OAI21_X1   g01943(.A1(new_n2009_), .A2(new_n2011_), .B(new_n1957_), .ZN(new_n2012_));
  INV_X1     g01944(.I(new_n2002_), .ZN(new_n2013_));
  OAI21_X1   g01945(.A1(new_n2005_), .A2(new_n2004_), .B(new_n2013_), .ZN(new_n2014_));
  INV_X1     g01946(.I(new_n2006_), .ZN(new_n2015_));
  NAND3_X1   g01947(.A1(new_n1995_), .A2(new_n2001_), .A3(new_n2015_), .ZN(new_n2016_));
  NAND2_X1   g01948(.A1(new_n2014_), .A2(new_n2016_), .ZN(new_n2017_));
  NAND3_X1   g01949(.A1(new_n2017_), .A2(new_n1954_), .A3(new_n1947_), .ZN(new_n2018_));
  INV_X1     g01950(.I(new_n2011_), .ZN(new_n2019_));
  NAND3_X1   g01951(.A1(new_n2018_), .A2(new_n1953_), .A3(new_n2019_), .ZN(new_n2020_));
  NAND3_X1   g01952(.A1(new_n2012_), .A2(new_n2020_), .A3(new_n786_), .ZN(new_n2021_));
  AOI21_X1   g01953(.A1(new_n2018_), .A2(new_n2019_), .B(new_n1953_), .ZN(new_n2022_));
  NOR3_X1    g01954(.A1(new_n2009_), .A2(new_n1957_), .A3(new_n2011_), .ZN(new_n2023_));
  OAI21_X1   g01955(.A1(new_n2023_), .A2(new_n2022_), .B(new_n644_), .ZN(new_n2024_));
  NAND4_X1   g01956(.A1(new_n2024_), .A2(new_n2021_), .A3(new_n1952_), .A4(new_n1956_), .ZN(new_n2025_));
  NAND2_X1   g01957(.A1(new_n1952_), .A2(new_n1956_), .ZN(new_n2026_));
  NAND2_X1   g01958(.A1(new_n2024_), .A2(new_n2021_), .ZN(new_n2027_));
  NAND2_X1   g01959(.A1(new_n2027_), .A2(new_n2026_), .ZN(new_n2028_));
  NAND3_X1   g01960(.A1(new_n2028_), .A2(new_n294_), .A3(new_n2025_), .ZN(new_n2029_));
  INV_X1     g01961(.I(new_n1694_), .ZN(new_n2030_));
  AOI21_X1   g01962(.A1(new_n2030_), .A2(new_n1703_), .B(new_n786_), .ZN(new_n2031_));
  OAI21_X1   g01963(.A1(new_n1715_), .A2(new_n1716_), .B(new_n1613_), .ZN(new_n2032_));
  NAND3_X1   g01964(.A1(new_n1713_), .A2(new_n1707_), .A3(new_n1686_), .ZN(new_n2033_));
  INV_X1     g01965(.I(new_n1794_), .ZN(new_n2034_));
  OAI21_X1   g01966(.A1(new_n1786_), .A2(new_n1789_), .B(new_n2034_), .ZN(new_n2035_));
  OAI21_X1   g01967(.A1(new_n1725_), .A2(new_n1724_), .B(new_n1723_), .ZN(new_n2036_));
  NAND3_X1   g01968(.A1(new_n1721_), .A2(new_n1719_), .A3(new_n1720_), .ZN(new_n2037_));
  NAND2_X1   g01969(.A1(new_n2037_), .A2(new_n2036_), .ZN(new_n2038_));
  INV_X1     g01970(.I(new_n1728_), .ZN(new_n2039_));
  AOI21_X1   g01971(.A1(new_n1478_), .A2(new_n1472_), .B(new_n443_), .ZN(new_n2040_));
  OAI21_X1   g01972(.A1(new_n2039_), .A2(new_n2040_), .B(new_n1471_), .ZN(new_n2041_));
  AOI21_X1   g01973(.A1(new_n1478_), .A2(new_n1472_), .B(new_n568_), .ZN(new_n2042_));
  OAI21_X1   g01974(.A1(new_n2042_), .A2(new_n1575_), .B(new_n1470_), .ZN(new_n2043_));
  NAND2_X1   g01975(.A1(new_n2041_), .A2(new_n2043_), .ZN(new_n2044_));
  XOR2_X1    g01976(.A1(\a[11] ), .A2(\a[12] ), .Z(new_n2045_));
  NOR2_X1    g01977(.A1(new_n2045_), .A2(new_n279_), .ZN(new_n2046_));
  OAI21_X1   g01978(.A1(new_n786_), .A2(new_n2046_), .B(new_n1747_), .ZN(new_n2047_));
  NOR3_X1    g01979(.A1(new_n1620_), .A2(new_n126_), .A3(new_n1468_), .ZN(new_n2048_));
  NOR2_X1    g01980(.A1(new_n443_), .A2(new_n1469_), .ZN(new_n2049_));
  OAI21_X1   g01981(.A1(new_n2049_), .A2(new_n2048_), .B(new_n644_), .ZN(new_n2050_));
  NAND2_X1   g01982(.A1(new_n2050_), .A2(new_n2047_), .ZN(new_n2051_));
  AOI22_X1   g01983(.A1(new_n2051_), .A2(new_n1740_), .B1(new_n1742_), .B2(new_n1744_), .ZN(new_n2052_));
  NAND2_X1   g01984(.A1(new_n2044_), .A2(new_n2052_), .ZN(new_n2053_));
  NOR3_X1    g01985(.A1(new_n1750_), .A2(new_n786_), .A3(new_n1745_), .ZN(new_n2054_));
  OAI21_X1   g01986(.A1(new_n2044_), .A2(new_n2052_), .B(new_n2054_), .ZN(new_n2055_));
  AOI21_X1   g01987(.A1(new_n1770_), .A2(new_n1771_), .B(new_n786_), .ZN(new_n2056_));
  AOI21_X1   g01988(.A1(new_n2055_), .A2(new_n2053_), .B(new_n2056_), .ZN(new_n2057_));
  INV_X1     g01989(.I(new_n1772_), .ZN(new_n2058_));
  NOR3_X1    g01990(.A1(new_n1782_), .A2(new_n1783_), .A3(new_n644_), .ZN(new_n2059_));
  NOR4_X1    g01991(.A1(new_n2057_), .A2(new_n2059_), .A3(new_n1787_), .A4(new_n2058_), .ZN(new_n2060_));
  NAND2_X1   g01992(.A1(new_n2060_), .A2(new_n2038_), .ZN(new_n2061_));
  NOR2_X1    g01993(.A1(new_n1784_), .A2(new_n644_), .ZN(new_n2062_));
  OAI21_X1   g01994(.A1(new_n2060_), .A2(new_n2038_), .B(new_n2062_), .ZN(new_n2063_));
  NAND3_X1   g01995(.A1(new_n2063_), .A2(new_n2061_), .A3(new_n1794_), .ZN(new_n2064_));
  NAND2_X1   g01996(.A1(new_n2064_), .A2(\a[14] ), .ZN(new_n2065_));
  INV_X1     g01997(.I(new_n1799_), .ZN(new_n2066_));
  AOI21_X1   g01998(.A1(new_n2065_), .A2(new_n2035_), .B(new_n2066_), .ZN(new_n2067_));
  INV_X1     g01999(.I(new_n1810_), .ZN(new_n2068_));
  OAI21_X1   g02000(.A1(new_n2067_), .A2(new_n1801_), .B(new_n2068_), .ZN(new_n2069_));
  INV_X1     g02001(.I(new_n1813_), .ZN(new_n2070_));
  AOI21_X1   g02002(.A1(new_n1824_), .A2(new_n1818_), .B(new_n786_), .ZN(new_n2071_));
  AOI21_X1   g02003(.A1(new_n2069_), .A2(new_n2070_), .B(new_n2071_), .ZN(new_n2072_));
  OAI21_X1   g02004(.A1(new_n1837_), .A2(new_n1838_), .B(new_n644_), .ZN(new_n2073_));
  OAI21_X1   g02005(.A1(new_n2072_), .A2(new_n1826_), .B(new_n2073_), .ZN(new_n2074_));
  INV_X1     g02006(.I(new_n1839_), .ZN(new_n2075_));
  INV_X1     g02007(.I(new_n1842_), .ZN(new_n2076_));
  OAI21_X1   g02008(.A1(new_n1605_), .A2(new_n1554_), .B(new_n1601_), .ZN(new_n2077_));
  AOI21_X1   g02009(.A1(new_n2076_), .A2(new_n2077_), .B(new_n786_), .ZN(new_n2078_));
  AOI21_X1   g02010(.A1(new_n2074_), .A2(new_n2075_), .B(new_n2078_), .ZN(new_n2079_));
  NAND3_X1   g02011(.A1(new_n1872_), .A2(new_n1868_), .A3(new_n1853_), .ZN(new_n2080_));
  OAI21_X1   g02012(.A1(new_n1864_), .A2(new_n1860_), .B(new_n1854_), .ZN(new_n2081_));
  NAND2_X1   g02013(.A1(new_n2081_), .A2(new_n2080_), .ZN(new_n2082_));
  OAI21_X1   g02014(.A1(new_n2079_), .A2(new_n1848_), .B(new_n2082_), .ZN(new_n2083_));
  AOI21_X1   g02015(.A1(new_n2032_), .A2(new_n2033_), .B(new_n2083_), .ZN(new_n2084_));
  NAND3_X1   g02016(.A1(new_n2083_), .A2(new_n2032_), .A3(new_n2033_), .ZN(new_n2085_));
  AOI21_X1   g02017(.A1(new_n2085_), .A2(new_n1888_), .B(new_n2084_), .ZN(new_n2086_));
  INV_X1     g02018(.I(new_n1891_), .ZN(new_n2087_));
  NOR3_X1    g02019(.A1(new_n2087_), .A2(new_n2030_), .A3(new_n1892_), .ZN(new_n2088_));
  NOR3_X1    g02020(.A1(new_n2088_), .A2(new_n2031_), .A3(new_n2086_), .ZN(new_n2089_));
  OAI21_X1   g02021(.A1(new_n1680_), .A2(new_n1684_), .B(new_n786_), .ZN(new_n2090_));
  NOR2_X1    g02022(.A1(new_n2089_), .A2(new_n2090_), .ZN(new_n2091_));
  OAI21_X1   g02023(.A1(new_n1683_), .A2(new_n1678_), .B(new_n1647_), .ZN(new_n2092_));
  NAND3_X1   g02024(.A1(new_n1679_), .A2(new_n1677_), .A3(new_n1433_), .ZN(new_n2093_));
  AOI21_X1   g02025(.A1(new_n2092_), .A2(new_n2093_), .B(new_n644_), .ZN(new_n2094_));
  NOR2_X1    g02026(.A1(new_n1895_), .A2(new_n2094_), .ZN(new_n2095_));
  OAI21_X1   g02027(.A1(new_n2091_), .A2(new_n2095_), .B(new_n1893_), .ZN(new_n2096_));
  NAND2_X1   g02028(.A1(new_n1895_), .A2(new_n2094_), .ZN(new_n2097_));
  NAND2_X1   g02029(.A1(new_n2089_), .A2(new_n2090_), .ZN(new_n2098_));
  NAND3_X1   g02030(.A1(new_n2098_), .A2(new_n2097_), .A3(new_n1892_), .ZN(new_n2099_));
  AND2_X2    g02031(.A1(new_n2096_), .A2(new_n2099_), .Z(new_n2100_));
  NAND2_X1   g02032(.A1(new_n2032_), .A2(new_n2033_), .ZN(new_n2101_));
  NAND3_X1   g02033(.A1(new_n2101_), .A2(new_n644_), .A3(new_n2083_), .ZN(new_n2102_));
  OAI21_X1   g02034(.A1(new_n1714_), .A2(new_n1717_), .B(new_n644_), .ZN(new_n2103_));
  NAND2_X1   g02035(.A1(new_n2103_), .A2(new_n1884_), .ZN(new_n2104_));
  AOI21_X1   g02036(.A1(new_n2104_), .A2(new_n2102_), .B(new_n1878_), .ZN(new_n2105_));
  NOR2_X1    g02037(.A1(new_n2103_), .A2(new_n1884_), .ZN(new_n2106_));
  AOI21_X1   g02038(.A1(new_n2101_), .A2(new_n644_), .B(new_n2083_), .ZN(new_n2107_));
  NOR3_X1    g02039(.A1(new_n2106_), .A2(new_n2107_), .A3(new_n1887_), .ZN(new_n2108_));
  NOR2_X1    g02040(.A1(new_n2108_), .A2(new_n2105_), .ZN(new_n2109_));
  INV_X1     g02041(.I(new_n2109_), .ZN(new_n2110_));
  NOR2_X1    g02042(.A1(new_n2079_), .A2(new_n1848_), .ZN(new_n2111_));
  NOR2_X1    g02043(.A1(new_n1865_), .A2(new_n1873_), .ZN(new_n2112_));
  INV_X1     g02044(.I(new_n2112_), .ZN(new_n2113_));
  NAND2_X1   g02045(.A1(new_n2111_), .A2(new_n2113_), .ZN(new_n2114_));
  NAND2_X1   g02046(.A1(new_n1847_), .A2(new_n1849_), .ZN(new_n2115_));
  NAND2_X1   g02047(.A1(new_n2115_), .A2(new_n2112_), .ZN(new_n2116_));
  NAND2_X1   g02048(.A1(new_n2114_), .A2(new_n2116_), .ZN(new_n2117_));
  NOR3_X1    g02049(.A1(new_n1878_), .A2(new_n1881_), .A3(new_n1865_), .ZN(new_n2118_));
  NOR3_X1    g02050(.A1(new_n2118_), .A2(new_n2115_), .A3(new_n2112_), .ZN(new_n2119_));
  NAND3_X1   g02051(.A1(new_n1875_), .A2(new_n1877_), .A3(new_n786_), .ZN(new_n2120_));
  NAND3_X1   g02052(.A1(new_n1887_), .A2(new_n2120_), .A3(new_n2080_), .ZN(new_n2121_));
  AOI21_X1   g02053(.A1(new_n2121_), .A2(new_n2113_), .B(new_n2111_), .ZN(new_n2122_));
  NOR2_X1    g02054(.A1(new_n2119_), .A2(new_n2122_), .ZN(new_n2123_));
  AOI21_X1   g02055(.A1(new_n2123_), .A2(new_n2117_), .B(new_n806_), .ZN(new_n2124_));
  NOR3_X1    g02056(.A1(new_n1845_), .A2(new_n786_), .A3(new_n1842_), .ZN(new_n2125_));
  AOI21_X1   g02057(.A1(new_n2076_), .A2(new_n2077_), .B(new_n644_), .ZN(new_n2126_));
  OAI22_X1   g02058(.A1(new_n2126_), .A2(new_n2125_), .B1(new_n1836_), .B2(new_n1839_), .ZN(new_n2127_));
  NOR2_X1    g02059(.A1(new_n1836_), .A2(new_n1839_), .ZN(new_n2128_));
  OAI21_X1   g02060(.A1(new_n2078_), .A2(new_n1848_), .B(new_n2128_), .ZN(new_n2129_));
  AND2_X2    g02061(.A1(new_n2129_), .A2(new_n2127_), .Z(new_n2130_));
  NOR3_X1    g02062(.A1(new_n1750_), .A2(new_n786_), .A3(new_n1745_), .ZN(new_n2131_));
  NOR3_X1    g02063(.A1(new_n1732_), .A2(new_n2052_), .A3(new_n786_), .ZN(new_n2132_));
  INV_X1     g02064(.I(new_n2132_), .ZN(new_n2133_));
  OAI21_X1   g02065(.A1(new_n786_), .A2(new_n1732_), .B(new_n2052_), .ZN(new_n2134_));
  AOI21_X1   g02066(.A1(new_n2133_), .A2(new_n2134_), .B(new_n2131_), .ZN(new_n2135_));
  INV_X1     g02067(.I(new_n2131_), .ZN(new_n2136_));
  INV_X1     g02068(.I(new_n2134_), .ZN(new_n2137_));
  NOR3_X1    g02069(.A1(new_n2137_), .A2(new_n2136_), .A3(new_n2132_), .ZN(new_n2138_));
  NOR2_X1    g02070(.A1(new_n2138_), .A2(new_n2135_), .ZN(new_n2139_));
  NAND3_X1   g02071(.A1(new_n1736_), .A2(new_n644_), .A3(new_n1737_), .ZN(new_n2140_));
  INV_X1     g02072(.I(new_n2140_), .ZN(new_n2141_));
  AOI21_X1   g02073(.A1(new_n1736_), .A2(new_n1737_), .B(new_n644_), .ZN(new_n2142_));
  OAI21_X1   g02074(.A1(new_n2141_), .A2(new_n2142_), .B(new_n2047_), .ZN(new_n2143_));
  OAI21_X1   g02075(.A1(new_n1741_), .A2(new_n1738_), .B(new_n1735_), .ZN(new_n2144_));
  NAND3_X1   g02076(.A1(new_n785_), .A2(new_n1734_), .A3(\a[14] ), .ZN(new_n2145_));
  NAND2_X1   g02077(.A1(new_n786_), .A2(new_n2046_), .ZN(new_n2146_));
  NOR4_X1    g02078(.A1(new_n801_), .A2(new_n294_), .A3(\a[8] ), .A4(\a[9] ), .ZN(new_n2147_));
  NOR2_X1    g02079(.A1(new_n2045_), .A2(new_n2147_), .ZN(new_n2148_));
  NAND4_X1   g02080(.A1(new_n498_), .A2(new_n1075_), .A3(\a[10] ), .A4(\a[11] ), .ZN(new_n2149_));
  NOR2_X1    g02081(.A1(new_n1733_), .A2(new_n2149_), .ZN(new_n2150_));
  AOI21_X1   g02082(.A1(new_n2146_), .A2(new_n2145_), .B(new_n1079_), .ZN(new_n2151_));
  NAND4_X1   g02083(.A1(new_n642_), .A2(new_n638_), .A3(new_n2045_), .A4(\a[14] ), .ZN(new_n2152_));
  NOR2_X1    g02084(.A1(new_n1079_), .A2(new_n2152_), .ZN(new_n2153_));
  INV_X1     g02085(.I(new_n2152_), .ZN(new_n2154_));
  NOR2_X1    g02086(.A1(new_n2154_), .A2(new_n806_), .ZN(new_n2155_));
  NOR3_X1    g02087(.A1(new_n786_), .A2(new_n1468_), .A3(new_n1734_), .ZN(new_n2156_));
  NAND2_X1   g02088(.A1(new_n644_), .A2(new_n1468_), .ZN(new_n2157_));
  NAND2_X1   g02089(.A1(new_n786_), .A2(new_n1747_), .ZN(new_n2158_));
  AOI22_X1   g02090(.A1(new_n2158_), .A2(new_n2157_), .B1(new_n644_), .B2(new_n2046_), .ZN(new_n2159_));
  NOR3_X1    g02091(.A1(new_n2159_), .A2(new_n1079_), .A3(new_n2156_), .ZN(new_n2160_));
  INV_X1     g02092(.I(new_n2156_), .ZN(new_n2161_));
  NOR2_X1    g02093(.A1(new_n786_), .A2(new_n1747_), .ZN(new_n2162_));
  NAND2_X1   g02094(.A1(new_n644_), .A2(new_n2046_), .ZN(new_n2163_));
  NOR2_X1    g02095(.A1(new_n644_), .A2(new_n1468_), .ZN(new_n2164_));
  OAI21_X1   g02096(.A1(new_n2162_), .A2(new_n2164_), .B(new_n2163_), .ZN(new_n2165_));
  AOI21_X1   g02097(.A1(new_n2165_), .A2(new_n2161_), .B(new_n806_), .ZN(new_n2166_));
  OAI21_X1   g02098(.A1(new_n2153_), .A2(new_n2155_), .B(new_n2151_), .ZN(new_n2167_));
  AOI21_X1   g02099(.A1(new_n2143_), .A2(new_n2144_), .B(new_n2167_), .ZN(new_n2168_));
  INV_X1     g02100(.I(new_n2142_), .ZN(new_n2169_));
  NAND2_X1   g02101(.A1(new_n2169_), .A2(new_n2140_), .ZN(new_n2170_));
  AOI21_X1   g02102(.A1(new_n2050_), .A2(new_n1740_), .B(new_n2047_), .ZN(new_n2171_));
  AOI21_X1   g02103(.A1(new_n2170_), .A2(new_n2047_), .B(new_n2171_), .ZN(new_n2172_));
  NAND3_X1   g02104(.A1(new_n2165_), .A2(new_n1079_), .A3(new_n2161_), .ZN(new_n2173_));
  AOI21_X1   g02105(.A1(new_n2172_), .A2(new_n2167_), .B(new_n2173_), .ZN(new_n2174_));
  NAND2_X1   g02106(.A1(new_n2051_), .A2(new_n1740_), .ZN(new_n2175_));
  NAND2_X1   g02107(.A1(new_n1744_), .A2(new_n1742_), .ZN(new_n2176_));
  INV_X1     g02108(.I(new_n2176_), .ZN(new_n2177_));
  NOR2_X1    g02109(.A1(new_n2175_), .A2(new_n2177_), .ZN(new_n2178_));
  NOR2_X1    g02110(.A1(new_n1739_), .A2(new_n1741_), .ZN(new_n2179_));
  NOR2_X1    g02111(.A1(new_n2179_), .A2(new_n2176_), .ZN(new_n2180_));
  OAI21_X1   g02112(.A1(new_n2180_), .A2(new_n2178_), .B(new_n1079_), .ZN(new_n2181_));
  OAI21_X1   g02113(.A1(new_n2174_), .A2(new_n2168_), .B(new_n2181_), .ZN(new_n2182_));
  NAND2_X1   g02114(.A1(new_n2179_), .A2(new_n2176_), .ZN(new_n2183_));
  NAND2_X1   g02115(.A1(new_n2175_), .A2(new_n2177_), .ZN(new_n2184_));
  NAND3_X1   g02116(.A1(new_n2183_), .A2(new_n2184_), .A3(new_n806_), .ZN(new_n2185_));
  NAND3_X1   g02117(.A1(new_n1756_), .A2(new_n1752_), .A3(new_n786_), .ZN(new_n2186_));
  OAI21_X1   g02118(.A1(new_n1750_), .A2(new_n1745_), .B(new_n644_), .ZN(new_n2187_));
  NAND3_X1   g02119(.A1(new_n2187_), .A2(new_n2186_), .A3(new_n1742_), .ZN(new_n2188_));
  NAND3_X1   g02120(.A1(new_n2188_), .A2(new_n2179_), .A3(new_n2176_), .ZN(new_n2189_));
  INV_X1     g02121(.I(new_n1742_), .ZN(new_n2190_));
  NOR3_X1    g02122(.A1(new_n1751_), .A2(new_n1757_), .A3(new_n2190_), .ZN(new_n2191_));
  OAI21_X1   g02123(.A1(new_n2191_), .A2(new_n2177_), .B(new_n2175_), .ZN(new_n2192_));
  NAND3_X1   g02124(.A1(new_n2192_), .A2(new_n2189_), .A3(new_n806_), .ZN(new_n2193_));
  NOR3_X1    g02125(.A1(new_n2191_), .A2(new_n2175_), .A3(new_n2177_), .ZN(new_n2194_));
  AOI21_X1   g02126(.A1(new_n2188_), .A2(new_n2176_), .B(new_n2179_), .ZN(new_n2195_));
  OAI21_X1   g02127(.A1(new_n2194_), .A2(new_n2195_), .B(new_n1079_), .ZN(new_n2196_));
  NAND4_X1   g02128(.A1(new_n2193_), .A2(new_n2196_), .A3(new_n2182_), .A4(new_n2185_), .ZN(new_n2197_));
  NOR2_X1    g02129(.A1(new_n2197_), .A2(new_n2139_), .ZN(new_n2198_));
  AOI21_X1   g02130(.A1(new_n2192_), .A2(new_n2189_), .B(new_n806_), .ZN(new_n2199_));
  NAND2_X1   g02131(.A1(new_n2199_), .A2(new_n806_), .ZN(new_n2200_));
  AOI21_X1   g02132(.A1(new_n2197_), .A2(new_n2139_), .B(new_n2200_), .ZN(new_n2201_));
  NAND2_X1   g02133(.A1(new_n2055_), .A2(new_n2053_), .ZN(new_n2202_));
  NAND2_X1   g02134(.A1(new_n1768_), .A2(new_n1772_), .ZN(new_n2203_));
  NAND2_X1   g02135(.A1(new_n2202_), .A2(new_n2203_), .ZN(new_n2204_));
  NAND2_X1   g02136(.A1(new_n1770_), .A2(new_n1771_), .ZN(new_n2205_));
  XOR2_X1    g02137(.A1(new_n2205_), .A2(new_n786_), .Z(new_n2206_));
  OAI21_X1   g02138(.A1(new_n2202_), .A2(new_n2206_), .B(new_n2204_), .ZN(new_n2207_));
  OAI21_X1   g02139(.A1(new_n2201_), .A2(new_n2198_), .B(new_n2207_), .ZN(new_n2208_));
  NOR3_X1    g02140(.A1(new_n2201_), .A2(new_n2198_), .A3(new_n2207_), .ZN(new_n2209_));
  OAI21_X1   g02141(.A1(new_n294_), .A2(new_n2209_), .B(new_n2208_), .ZN(new_n2210_));
  AOI22_X1   g02142(.A1(new_n1784_), .A2(new_n1781_), .B1(new_n1769_), .B2(new_n1772_), .ZN(new_n2211_));
  NOR2_X1    g02143(.A1(new_n2060_), .A2(new_n2211_), .ZN(new_n2212_));
  NAND2_X1   g02144(.A1(new_n2212_), .A2(new_n1079_), .ZN(new_n2213_));
  NOR2_X1    g02145(.A1(new_n2212_), .A2(new_n1079_), .ZN(new_n2214_));
  AOI21_X1   g02146(.A1(new_n2210_), .A2(new_n2213_), .B(new_n2214_), .ZN(new_n2215_));
  NOR2_X1    g02147(.A1(new_n1727_), .A2(new_n644_), .ZN(new_n2216_));
  XOR2_X1    g02148(.A1(new_n2216_), .A2(new_n2060_), .Z(new_n2217_));
  NAND2_X1   g02149(.A1(new_n2217_), .A2(new_n1784_), .ZN(new_n2218_));
  XOR2_X1    g02150(.A1(new_n2216_), .A2(new_n1785_), .Z(new_n2219_));
  NAND2_X1   g02151(.A1(new_n2219_), .A2(new_n1787_), .ZN(new_n2220_));
  AOI21_X1   g02152(.A1(new_n2220_), .A2(new_n2218_), .B(new_n1079_), .ZN(new_n2221_));
  NAND3_X1   g02153(.A1(new_n2220_), .A2(new_n2218_), .A3(new_n1079_), .ZN(new_n2222_));
  OAI21_X1   g02154(.A1(new_n2215_), .A2(new_n2221_), .B(new_n2222_), .ZN(new_n2223_));
  NAND2_X1   g02155(.A1(new_n1790_), .A2(new_n2034_), .ZN(new_n2224_));
  NOR2_X1    g02156(.A1(new_n1790_), .A2(new_n2034_), .ZN(new_n2225_));
  INV_X1     g02157(.I(new_n2225_), .ZN(new_n2226_));
  AOI21_X1   g02158(.A1(new_n2226_), .A2(new_n2224_), .B(\a[14] ), .ZN(new_n2227_));
  INV_X1     g02159(.I(new_n2224_), .ZN(new_n2228_));
  NOR3_X1    g02160(.A1(new_n2228_), .A2(new_n279_), .A3(new_n2225_), .ZN(new_n2229_));
  OAI21_X1   g02161(.A1(new_n2227_), .A2(new_n2229_), .B(new_n1079_), .ZN(new_n2230_));
  NOR3_X1    g02162(.A1(new_n2227_), .A2(new_n2229_), .A3(new_n1079_), .ZN(new_n2231_));
  AOI21_X1   g02163(.A1(new_n2223_), .A2(new_n2230_), .B(new_n2231_), .ZN(new_n2232_));
  NAND2_X1   g02164(.A1(new_n2065_), .A2(new_n2035_), .ZN(new_n2233_));
  XOR2_X1    g02165(.A1(new_n1798_), .A2(new_n786_), .Z(new_n2234_));
  INV_X1     g02166(.I(new_n2234_), .ZN(new_n2235_));
  NAND2_X1   g02167(.A1(new_n2233_), .A2(new_n2235_), .ZN(new_n2236_));
  NOR2_X1    g02168(.A1(new_n1796_), .A2(new_n1795_), .ZN(new_n2237_));
  NAND2_X1   g02169(.A1(new_n1802_), .A2(new_n1799_), .ZN(new_n2238_));
  NAND2_X1   g02170(.A1(new_n2237_), .A2(new_n2238_), .ZN(new_n2239_));
  AOI21_X1   g02171(.A1(new_n2236_), .A2(new_n2239_), .B(new_n806_), .ZN(new_n2240_));
  NAND3_X1   g02172(.A1(new_n2236_), .A2(new_n2239_), .A3(new_n806_), .ZN(new_n2241_));
  OAI21_X1   g02173(.A1(new_n2232_), .A2(new_n2240_), .B(new_n2241_), .ZN(new_n2242_));
  NAND2_X1   g02174(.A1(new_n1800_), .A2(new_n1802_), .ZN(new_n2243_));
  NAND3_X1   g02175(.A1(new_n1806_), .A2(new_n1809_), .A3(new_n786_), .ZN(new_n2244_));
  NAND2_X1   g02176(.A1(new_n1812_), .A2(new_n644_), .ZN(new_n2245_));
  NAND2_X1   g02177(.A1(new_n2245_), .A2(new_n2244_), .ZN(new_n2246_));
  NAND2_X1   g02178(.A1(new_n2243_), .A2(new_n2246_), .ZN(new_n2247_));
  INV_X1     g02179(.I(new_n2247_), .ZN(new_n2248_));
  AOI21_X1   g02180(.A1(new_n2068_), .A2(new_n2070_), .B(new_n2243_), .ZN(new_n2249_));
  OAI21_X1   g02181(.A1(new_n2248_), .A2(new_n2249_), .B(new_n1079_), .ZN(new_n2250_));
  NOR2_X1    g02182(.A1(new_n2067_), .A2(new_n1801_), .ZN(new_n2251_));
  OAI21_X1   g02183(.A1(new_n1810_), .A2(new_n1813_), .B(new_n2251_), .ZN(new_n2252_));
  NAND3_X1   g02184(.A1(new_n2252_), .A2(new_n806_), .A3(new_n2247_), .ZN(new_n2253_));
  INV_X1     g02185(.I(new_n2253_), .ZN(new_n2254_));
  AOI21_X1   g02186(.A1(new_n2242_), .A2(new_n2250_), .B(new_n2254_), .ZN(new_n2255_));
  INV_X1     g02187(.I(new_n2255_), .ZN(new_n2256_));
  NOR3_X1    g02188(.A1(new_n801_), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n2257_));
  AOI21_X1   g02189(.A1(\a[9] ), .A2(new_n803_), .B(new_n2257_), .ZN(new_n2258_));
  NOR2_X1    g02190(.A1(new_n1078_), .A2(new_n2258_), .ZN(new_n2259_));
  XOR2_X1    g02191(.A1(new_n2259_), .A2(new_n294_), .Z(new_n2260_));
  NAND2_X1   g02192(.A1(new_n2069_), .A2(new_n2070_), .ZN(new_n2261_));
  OAI21_X1   g02193(.A1(new_n2071_), .A2(new_n1826_), .B(new_n2261_), .ZN(new_n2262_));
  NOR2_X1    g02194(.A1(new_n1811_), .A2(new_n1813_), .ZN(new_n2263_));
  NAND3_X1   g02195(.A1(new_n1824_), .A2(new_n1818_), .A3(new_n644_), .ZN(new_n2264_));
  NAND2_X1   g02196(.A1(new_n1825_), .A2(new_n786_), .ZN(new_n2265_));
  NAND2_X1   g02197(.A1(new_n2265_), .A2(new_n2264_), .ZN(new_n2266_));
  NAND2_X1   g02198(.A1(new_n2266_), .A2(new_n2263_), .ZN(new_n2267_));
  NAND3_X1   g02199(.A1(new_n2262_), .A2(new_n2260_), .A3(new_n2267_), .ZN(new_n2268_));
  INV_X1     g02200(.I(new_n2260_), .ZN(new_n2269_));
  AOI21_X1   g02201(.A1(new_n1820_), .A2(new_n1827_), .B(new_n2263_), .ZN(new_n2270_));
  AOI21_X1   g02202(.A1(new_n2264_), .A2(new_n2265_), .B(new_n2261_), .ZN(new_n2271_));
  OAI21_X1   g02203(.A1(new_n2271_), .A2(new_n2270_), .B(new_n2269_), .ZN(new_n2272_));
  AOI22_X1   g02204(.A1(new_n2073_), .A2(new_n2075_), .B1(new_n1821_), .B2(new_n1827_), .ZN(new_n2273_));
  NAND3_X1   g02205(.A1(new_n1832_), .A2(new_n1834_), .A3(new_n644_), .ZN(new_n2274_));
  OAI21_X1   g02206(.A1(new_n1837_), .A2(new_n1838_), .B(new_n786_), .ZN(new_n2275_));
  NAND2_X1   g02207(.A1(new_n2274_), .A2(new_n2275_), .ZN(new_n2276_));
  NAND3_X1   g02208(.A1(new_n2276_), .A2(new_n1821_), .A3(new_n1827_), .ZN(new_n2277_));
  INV_X1     g02209(.I(new_n2277_), .ZN(new_n2278_));
  NOR3_X1    g02210(.A1(new_n2278_), .A2(new_n806_), .A3(new_n2273_), .ZN(new_n2279_));
  INV_X1     g02211(.I(new_n2273_), .ZN(new_n2280_));
  AOI21_X1   g02212(.A1(new_n2280_), .A2(new_n2277_), .B(new_n1079_), .ZN(new_n2281_));
  NAND2_X1   g02213(.A1(new_n2272_), .A2(new_n2268_), .ZN(new_n2283_));
  NAND2_X1   g02214(.A1(new_n2256_), .A2(new_n2283_), .ZN(new_n2284_));
  NOR2_X1    g02215(.A1(new_n2284_), .A2(new_n2130_), .ZN(new_n2285_));
  NAND2_X1   g02216(.A1(new_n2279_), .A2(new_n1079_), .ZN(new_n2286_));
  AOI21_X1   g02217(.A1(new_n2284_), .A2(new_n2130_), .B(new_n2286_), .ZN(new_n2287_));
  NOR2_X1    g02218(.A1(new_n2287_), .A2(new_n2285_), .ZN(new_n2288_));
  NOR3_X1    g02219(.A1(new_n2119_), .A2(new_n2122_), .A3(new_n806_), .ZN(new_n2289_));
  NAND3_X1   g02220(.A1(new_n2121_), .A2(new_n2111_), .A3(new_n2113_), .ZN(new_n2290_));
  OAI21_X1   g02221(.A1(new_n2118_), .A2(new_n2112_), .B(new_n2115_), .ZN(new_n2291_));
  AOI21_X1   g02222(.A1(new_n2291_), .A2(new_n2290_), .B(new_n1079_), .ZN(new_n2292_));
  NOR3_X1    g02223(.A1(new_n2289_), .A2(new_n2292_), .A3(new_n2117_), .ZN(new_n2293_));
  NOR3_X1    g02224(.A1(new_n2293_), .A2(new_n2124_), .A3(new_n2288_), .ZN(new_n2294_));
  NAND2_X1   g02225(.A1(new_n2294_), .A2(new_n2110_), .ZN(new_n2295_));
  NAND2_X1   g02226(.A1(new_n2291_), .A2(new_n2290_), .ZN(new_n2296_));
  NAND2_X1   g02227(.A1(new_n2296_), .A2(new_n1079_), .ZN(new_n2297_));
  NOR2_X1    g02228(.A1(new_n2297_), .A2(new_n1079_), .ZN(new_n2298_));
  OAI21_X1   g02229(.A1(new_n2294_), .A2(new_n2110_), .B(new_n2298_), .ZN(new_n2299_));
  NAND2_X1   g02230(.A1(new_n2299_), .A2(new_n2295_), .ZN(new_n2300_));
  NAND2_X1   g02231(.A1(new_n2085_), .A2(new_n1888_), .ZN(new_n2301_));
  NAND2_X1   g02232(.A1(new_n1708_), .A2(new_n1711_), .ZN(new_n2302_));
  OAI21_X1   g02233(.A1(new_n1708_), .A2(new_n1711_), .B(new_n1614_), .ZN(new_n2303_));
  NAND3_X1   g02234(.A1(new_n1636_), .A2(new_n2303_), .A3(new_n2302_), .ZN(new_n2304_));
  OAI21_X1   g02235(.A1(new_n1561_), .A2(new_n1688_), .B(new_n1691_), .ZN(new_n2305_));
  NAND3_X1   g02236(.A1(new_n2305_), .A2(new_n786_), .A3(new_n2304_), .ZN(new_n2306_));
  OAI21_X1   g02237(.A1(new_n1693_), .A2(new_n1692_), .B(new_n644_), .ZN(new_n2307_));
  NAND2_X1   g02238(.A1(new_n2307_), .A2(new_n2306_), .ZN(new_n2308_));
  NAND3_X1   g02239(.A1(new_n2308_), .A2(new_n1885_), .A3(new_n2301_), .ZN(new_n2309_));
  NOR3_X1    g02240(.A1(new_n1693_), .A2(new_n1692_), .A3(new_n644_), .ZN(new_n2310_));
  AOI21_X1   g02241(.A1(new_n2305_), .A2(new_n2304_), .B(new_n786_), .ZN(new_n2311_));
  NOR2_X1    g02242(.A1(new_n2310_), .A2(new_n2311_), .ZN(new_n2312_));
  NAND2_X1   g02243(.A1(new_n1890_), .A2(new_n2312_), .ZN(new_n2313_));
  AOI21_X1   g02244(.A1(new_n2313_), .A2(new_n2309_), .B(new_n2259_), .ZN(new_n2314_));
  INV_X1     g02245(.I(new_n2259_), .ZN(new_n2315_));
  NOR2_X1    g02246(.A1(new_n1890_), .A2(new_n2312_), .ZN(new_n2316_));
  NOR2_X1    g02247(.A1(new_n2086_), .A2(new_n2308_), .ZN(new_n2317_));
  NOR3_X1    g02248(.A1(new_n2317_), .A2(new_n2316_), .A3(new_n2315_), .ZN(new_n2318_));
  OAI21_X1   g02249(.A1(new_n2318_), .A2(new_n2314_), .B(new_n294_), .ZN(new_n2319_));
  OAI21_X1   g02250(.A1(new_n2317_), .A2(new_n2316_), .B(new_n2315_), .ZN(new_n2320_));
  NAND3_X1   g02251(.A1(new_n2313_), .A2(new_n2309_), .A3(new_n2259_), .ZN(new_n2321_));
  NAND3_X1   g02252(.A1(new_n2320_), .A2(new_n2321_), .A3(\a[11] ), .ZN(new_n2322_));
  NAND2_X1   g02253(.A1(new_n2319_), .A2(new_n2322_), .ZN(new_n2323_));
  XOR2_X1    g02254(.A1(new_n2308_), .A2(\a[11] ), .Z(new_n2324_));
  XOR2_X1    g02255(.A1(new_n1890_), .A2(new_n2259_), .Z(new_n2325_));
  NAND2_X1   g02256(.A1(new_n2325_), .A2(new_n2324_), .ZN(new_n2326_));
  MUX2_X1    g02257(.I0(new_n786_), .I1(new_n2030_), .S(new_n1703_), .Z(new_n2327_));
  NAND2_X1   g02258(.A1(new_n2327_), .A2(new_n2086_), .ZN(new_n2328_));
  MUX2_X1    g02259(.I0(new_n644_), .I1(new_n1694_), .S(new_n1703_), .Z(new_n2329_));
  NAND2_X1   g02260(.A1(new_n2329_), .A2(new_n1890_), .ZN(new_n2330_));
  NAND3_X1   g02261(.A1(new_n2328_), .A2(new_n2330_), .A3(new_n1079_), .ZN(new_n2331_));
  NOR2_X1    g02262(.A1(new_n2329_), .A2(new_n1890_), .ZN(new_n2332_));
  NOR2_X1    g02263(.A1(new_n2327_), .A2(new_n2086_), .ZN(new_n2333_));
  OAI21_X1   g02264(.A1(new_n2332_), .A2(new_n2333_), .B(new_n806_), .ZN(new_n2334_));
  AOI21_X1   g02265(.A1(new_n2334_), .A2(new_n2331_), .B(new_n2326_), .ZN(new_n2335_));
  OAI21_X1   g02266(.A1(new_n2335_), .A2(new_n2323_), .B(new_n2300_), .ZN(new_n2336_));
  NOR2_X1    g02267(.A1(new_n2100_), .A2(new_n2336_), .ZN(new_n2337_));
  NOR2_X1    g02268(.A1(new_n2331_), .A2(new_n806_), .ZN(new_n2338_));
  INV_X1     g02269(.I(new_n2338_), .ZN(new_n2339_));
  AOI21_X1   g02270(.A1(new_n2100_), .A2(new_n2336_), .B(new_n2339_), .ZN(new_n2340_));
  NOR2_X1    g02271(.A1(new_n2340_), .A2(new_n2337_), .ZN(new_n2341_));
  NOR2_X1    g02272(.A1(new_n1898_), .A2(new_n1896_), .ZN(new_n2342_));
  AOI21_X1   g02273(.A1(new_n1955_), .A2(new_n1949_), .B(new_n786_), .ZN(new_n2343_));
  NOR3_X1    g02274(.A1(new_n1950_), .A2(new_n644_), .A3(new_n1945_), .ZN(new_n2344_));
  NOR3_X1    g02275(.A1(new_n2344_), .A2(new_n2343_), .A3(new_n806_), .ZN(new_n2345_));
  INV_X1     g02276(.I(new_n2345_), .ZN(new_n2346_));
  OAI21_X1   g02277(.A1(new_n2344_), .A2(new_n2343_), .B(new_n806_), .ZN(new_n2347_));
  AOI21_X1   g02278(.A1(new_n2346_), .A2(new_n2347_), .B(new_n2342_), .ZN(new_n2348_));
  AOI21_X1   g02279(.A1(new_n1951_), .A2(new_n1956_), .B(new_n806_), .ZN(new_n2349_));
  INV_X1     g02280(.I(new_n2349_), .ZN(new_n2350_));
  NOR2_X1    g02281(.A1(new_n2344_), .A2(new_n2343_), .ZN(new_n2351_));
  NAND2_X1   g02282(.A1(new_n2351_), .A2(new_n806_), .ZN(new_n2352_));
  NAND2_X1   g02283(.A1(new_n2352_), .A2(new_n2350_), .ZN(new_n2353_));
  AOI21_X1   g02284(.A1(new_n2342_), .A2(new_n2353_), .B(new_n2348_), .ZN(new_n2354_));
  NAND2_X1   g02285(.A1(new_n2028_), .A2(new_n2025_), .ZN(new_n2355_));
  XOR2_X1    g02286(.A1(new_n2342_), .A2(new_n2351_), .Z(new_n2356_));
  NAND4_X1   g02287(.A1(new_n2355_), .A2(\a[11] ), .A3(new_n805_), .A4(new_n2356_), .ZN(new_n2357_));
  AOI21_X1   g02288(.A1(new_n2357_), .A2(new_n2354_), .B(new_n2341_), .ZN(new_n2358_));
  AOI21_X1   g02289(.A1(new_n2012_), .A2(new_n2020_), .B(new_n786_), .ZN(new_n2359_));
  INV_X1     g02290(.I(new_n2010_), .ZN(new_n2360_));
  AOI21_X1   g02291(.A1(new_n2017_), .A2(new_n568_), .B(new_n2360_), .ZN(new_n2361_));
  OAI21_X1   g02292(.A1(new_n2017_), .A2(new_n568_), .B(new_n1953_), .ZN(new_n2362_));
  NOR2_X1    g02293(.A1(new_n2361_), .A2(new_n2362_), .ZN(new_n2363_));
  NOR2_X1    g02294(.A1(new_n1009_), .A2(new_n1011_), .ZN(new_n2364_));
  AOI21_X1   g02295(.A1(new_n1007_), .A2(new_n1003_), .B(new_n2364_), .ZN(new_n2365_));
  XOR2_X1    g02296(.A1(new_n1008_), .A2(new_n71_), .Z(new_n2366_));
  INV_X1     g02297(.I(new_n2366_), .ZN(new_n2367_));
  NAND3_X1   g02298(.A1(new_n1007_), .A2(new_n1003_), .A3(new_n2367_), .ZN(new_n2368_));
  INV_X1     g02299(.I(new_n2368_), .ZN(new_n2369_));
  OAI21_X1   g02300(.A1(new_n2369_), .A2(new_n2365_), .B(new_n248_), .ZN(new_n2370_));
  AOI21_X1   g02301(.A1(new_n1981_), .A2(new_n1982_), .B(new_n2370_), .ZN(new_n2371_));
  INV_X1     g02302(.I(new_n2365_), .ZN(new_n2372_));
  AOI21_X1   g02303(.A1(new_n2372_), .A2(new_n2368_), .B(new_n189_), .ZN(new_n2373_));
  NOR3_X1    g02304(.A1(new_n1989_), .A2(new_n2373_), .A3(new_n1983_), .ZN(new_n2374_));
  OAI21_X1   g02305(.A1(new_n2371_), .A2(new_n2374_), .B(new_n1988_), .ZN(new_n2375_));
  OAI21_X1   g02306(.A1(new_n1989_), .A2(new_n1983_), .B(new_n2373_), .ZN(new_n2376_));
  NAND3_X1   g02307(.A1(new_n1981_), .A2(new_n2370_), .A3(new_n1982_), .ZN(new_n2377_));
  NAND3_X1   g02308(.A1(new_n2376_), .A2(new_n2377_), .A3(new_n1980_), .ZN(new_n2378_));
  AOI21_X1   g02309(.A1(new_n2375_), .A2(new_n2378_), .B(new_n273_), .ZN(new_n2379_));
  NAND2_X1   g02310(.A1(new_n1995_), .A2(new_n2379_), .ZN(new_n2380_));
  AOI21_X1   g02311(.A1(new_n2376_), .A2(new_n2377_), .B(new_n1980_), .ZN(new_n2381_));
  NOR3_X1    g02312(.A1(new_n2371_), .A2(new_n2374_), .A3(new_n1988_), .ZN(new_n2382_));
  OAI21_X1   g02313(.A1(new_n2382_), .A2(new_n2381_), .B(new_n356_), .ZN(new_n2383_));
  NAND2_X1   g02314(.A1(new_n2004_), .A2(new_n2383_), .ZN(new_n2384_));
  AOI21_X1   g02315(.A1(new_n2380_), .A2(new_n2384_), .B(new_n2000_), .ZN(new_n2385_));
  NOR2_X1    g02316(.A1(new_n2004_), .A2(new_n2383_), .ZN(new_n2386_));
  NOR2_X1    g02317(.A1(new_n1995_), .A2(new_n2379_), .ZN(new_n2387_));
  NOR3_X1    g02318(.A1(new_n2387_), .A2(new_n2386_), .A3(new_n1994_), .ZN(new_n2388_));
  OAI21_X1   g02319(.A1(new_n2385_), .A2(new_n2388_), .B(new_n568_), .ZN(new_n2389_));
  NOR2_X1    g02320(.A1(new_n2363_), .A2(new_n2389_), .ZN(new_n2390_));
  OAI21_X1   g02321(.A1(new_n2387_), .A2(new_n2386_), .B(new_n1994_), .ZN(new_n2391_));
  NAND3_X1   g02322(.A1(new_n2380_), .A2(new_n2384_), .A3(new_n2000_), .ZN(new_n2392_));
  AOI21_X1   g02323(.A1(new_n2391_), .A2(new_n2392_), .B(new_n443_), .ZN(new_n2393_));
  NOR3_X1    g02324(.A1(new_n2393_), .A2(new_n2361_), .A3(new_n2362_), .ZN(new_n2394_));
  OAI21_X1   g02325(.A1(new_n2390_), .A2(new_n2394_), .B(new_n2016_), .ZN(new_n2395_));
  OAI21_X1   g02326(.A1(new_n2361_), .A2(new_n2362_), .B(new_n2393_), .ZN(new_n2396_));
  OR3_X2     g02327(.A1(new_n2393_), .A2(new_n2361_), .A3(new_n2362_), .Z(new_n2397_));
  NAND3_X1   g02328(.A1(new_n2397_), .A2(new_n2396_), .A3(new_n2007_), .ZN(new_n2398_));
  NAND2_X1   g02329(.A1(new_n2395_), .A2(new_n2398_), .ZN(new_n2399_));
  NAND3_X1   g02330(.A1(new_n2399_), .A2(new_n2025_), .A3(new_n644_), .ZN(new_n2400_));
  NOR2_X1    g02331(.A1(new_n2027_), .A2(new_n2026_), .ZN(new_n2401_));
  AOI21_X1   g02332(.A1(new_n2397_), .A2(new_n2396_), .B(new_n2007_), .ZN(new_n2402_));
  NOR3_X1    g02333(.A1(new_n2390_), .A2(new_n2394_), .A3(new_n2016_), .ZN(new_n2403_));
  OAI21_X1   g02334(.A1(new_n2403_), .A2(new_n2402_), .B(new_n644_), .ZN(new_n2404_));
  NAND2_X1   g02335(.A1(new_n2401_), .A2(new_n2404_), .ZN(new_n2405_));
  AOI21_X1   g02336(.A1(new_n2405_), .A2(new_n2400_), .B(new_n2359_), .ZN(new_n2406_));
  NOR2_X1    g02337(.A1(new_n2401_), .A2(new_n2404_), .ZN(new_n2407_));
  AOI21_X1   g02338(.A1(new_n2399_), .A2(new_n644_), .B(new_n2025_), .ZN(new_n2408_));
  NOR3_X1    g02339(.A1(new_n2407_), .A2(new_n2408_), .A3(new_n2024_), .ZN(new_n2409_));
  OAI21_X1   g02340(.A1(new_n2409_), .A2(new_n2406_), .B(new_n806_), .ZN(new_n2410_));
  NOR2_X1    g02341(.A1(new_n2410_), .A2(new_n2358_), .ZN(new_n2411_));
  NAND2_X1   g02342(.A1(new_n2096_), .A2(new_n2099_), .ZN(new_n2412_));
  NOR4_X1    g02343(.A1(new_n2109_), .A2(new_n2293_), .A3(new_n2124_), .A4(new_n2288_), .ZN(new_n2413_));
  INV_X1     g02344(.I(new_n2117_), .ZN(new_n2414_));
  OAI21_X1   g02345(.A1(new_n2296_), .A2(new_n2414_), .B(new_n1079_), .ZN(new_n2415_));
  NAND2_X1   g02346(.A1(new_n2129_), .A2(new_n2127_), .ZN(new_n2416_));
  AOI21_X1   g02347(.A1(new_n2268_), .A2(new_n2272_), .B(new_n2255_), .ZN(new_n2417_));
  NAND2_X1   g02348(.A1(new_n2417_), .A2(new_n2416_), .ZN(new_n2418_));
  NAND3_X1   g02349(.A1(new_n2280_), .A2(new_n1079_), .A3(new_n2277_), .ZN(new_n2419_));
  NOR2_X1    g02350(.A1(new_n2419_), .A2(new_n806_), .ZN(new_n2420_));
  OAI21_X1   g02351(.A1(new_n2417_), .A2(new_n2416_), .B(new_n2420_), .ZN(new_n2421_));
  NAND2_X1   g02352(.A1(new_n2421_), .A2(new_n2418_), .ZN(new_n2422_));
  NAND3_X1   g02353(.A1(new_n2291_), .A2(new_n2290_), .A3(new_n1079_), .ZN(new_n2423_));
  OAI21_X1   g02354(.A1(new_n2119_), .A2(new_n2122_), .B(new_n806_), .ZN(new_n2424_));
  NAND3_X1   g02355(.A1(new_n2424_), .A2(new_n2423_), .A3(new_n2414_), .ZN(new_n2425_));
  NAND3_X1   g02356(.A1(new_n2425_), .A2(new_n2415_), .A3(new_n2422_), .ZN(new_n2426_));
  NAND2_X1   g02357(.A1(new_n2426_), .A2(new_n2109_), .ZN(new_n2427_));
  AOI21_X1   g02358(.A1(new_n2427_), .A2(new_n2298_), .B(new_n2413_), .ZN(new_n2428_));
  AOI21_X1   g02359(.A1(new_n2320_), .A2(new_n2321_), .B(\a[11] ), .ZN(new_n2429_));
  NOR3_X1    g02360(.A1(new_n2318_), .A2(new_n2314_), .A3(new_n294_), .ZN(new_n2430_));
  NOR2_X1    g02361(.A1(new_n2430_), .A2(new_n2429_), .ZN(new_n2431_));
  XOR2_X1    g02362(.A1(new_n2308_), .A2(new_n294_), .Z(new_n2432_));
  XOR2_X1    g02363(.A1(new_n1890_), .A2(new_n2315_), .Z(new_n2433_));
  NOR2_X1    g02364(.A1(new_n2433_), .A2(new_n2432_), .ZN(new_n2434_));
  NOR3_X1    g02365(.A1(new_n2332_), .A2(new_n2333_), .A3(new_n806_), .ZN(new_n2435_));
  AOI21_X1   g02366(.A1(new_n2328_), .A2(new_n2330_), .B(new_n1079_), .ZN(new_n2436_));
  OAI21_X1   g02367(.A1(new_n2436_), .A2(new_n2435_), .B(new_n2434_), .ZN(new_n2437_));
  AOI21_X1   g02368(.A1(new_n2437_), .A2(new_n2431_), .B(new_n2428_), .ZN(new_n2438_));
  NAND2_X1   g02369(.A1(new_n2438_), .A2(new_n2412_), .ZN(new_n2439_));
  OAI21_X1   g02370(.A1(new_n2438_), .A2(new_n2412_), .B(new_n2338_), .ZN(new_n2440_));
  NAND2_X1   g02371(.A1(new_n2440_), .A2(new_n2439_), .ZN(new_n2441_));
  OR2_X2     g02372(.A1(new_n1898_), .A2(new_n1896_), .Z(new_n2442_));
  AOI21_X1   g02373(.A1(new_n1951_), .A2(new_n1956_), .B(new_n1079_), .ZN(new_n2443_));
  OAI22_X1   g02374(.A1(new_n2345_), .A2(new_n2443_), .B1(new_n1896_), .B2(new_n1898_), .ZN(new_n2444_));
  NAND2_X1   g02375(.A1(new_n1951_), .A2(new_n1956_), .ZN(new_n2445_));
  NOR2_X1    g02376(.A1(new_n2445_), .A2(new_n1079_), .ZN(new_n2446_));
  NOR2_X1    g02377(.A1(new_n2446_), .A2(new_n2349_), .ZN(new_n2447_));
  OAI21_X1   g02378(.A1(new_n2447_), .A2(new_n2442_), .B(new_n2444_), .ZN(new_n2448_));
  NAND2_X1   g02379(.A1(new_n2356_), .A2(new_n1079_), .ZN(new_n2449_));
  AOI22_X1   g02380(.A1(new_n2024_), .A2(new_n2021_), .B1(new_n1952_), .B2(new_n1956_), .ZN(new_n2450_));
  OAI21_X1   g02381(.A1(new_n2401_), .A2(new_n2450_), .B(\a[11] ), .ZN(new_n2451_));
  AOI21_X1   g02382(.A1(new_n2451_), .A2(new_n2029_), .B(new_n2449_), .ZN(new_n2452_));
  OAI21_X1   g02383(.A1(new_n2452_), .A2(new_n2448_), .B(new_n2441_), .ZN(new_n2453_));
  OAI21_X1   g02384(.A1(new_n2407_), .A2(new_n2408_), .B(new_n2024_), .ZN(new_n2454_));
  NAND3_X1   g02385(.A1(new_n2405_), .A2(new_n2400_), .A3(new_n2359_), .ZN(new_n2455_));
  AOI21_X1   g02386(.A1(new_n2454_), .A2(new_n2455_), .B(new_n1079_), .ZN(new_n2456_));
  NOR2_X1    g02387(.A1(new_n2453_), .A2(new_n2456_), .ZN(new_n2457_));
  OAI21_X1   g02388(.A1(new_n2457_), .A2(new_n2411_), .B(new_n2029_), .ZN(new_n2458_));
  NOR3_X1    g02389(.A1(new_n2401_), .A2(\a[11] ), .A3(new_n2450_), .ZN(new_n2459_));
  NAND2_X1   g02390(.A1(new_n2453_), .A2(new_n2456_), .ZN(new_n2460_));
  NAND2_X1   g02391(.A1(new_n2410_), .A2(new_n2358_), .ZN(new_n2461_));
  NAND3_X1   g02392(.A1(new_n2460_), .A2(new_n2461_), .A3(new_n2459_), .ZN(new_n2462_));
  NAND2_X1   g02393(.A1(new_n2458_), .A2(new_n2462_), .ZN(new_n2463_));
  XNOR2_X1   g02394(.A1(\a[6] ), .A2(\a[8] ), .ZN(new_n2464_));
  INV_X1     g02395(.I(\a[7] ), .ZN(new_n2465_));
  NOR2_X1    g02396(.A1(new_n2465_), .A2(\a[5] ), .ZN(new_n2466_));
  NOR2_X1    g02397(.A1(new_n452_), .A2(\a[7] ), .ZN(new_n2467_));
  NOR2_X1    g02398(.A1(new_n2466_), .A2(new_n2467_), .ZN(new_n2468_));
  NOR2_X1    g02399(.A1(new_n2468_), .A2(new_n2464_), .ZN(new_n2469_));
  NAND2_X1   g02400(.A1(new_n2469_), .A2(\a[8] ), .ZN(new_n2470_));
  NOR3_X1    g02401(.A1(new_n2354_), .A2(new_n2340_), .A3(new_n2337_), .ZN(new_n2471_));
  AOI21_X1   g02402(.A1(new_n2440_), .A2(new_n2439_), .B(new_n2448_), .ZN(new_n2472_));
  NOR2_X1    g02403(.A1(new_n2471_), .A2(new_n2472_), .ZN(new_n2473_));
  INV_X1     g02404(.I(new_n2473_), .ZN(new_n2474_));
  NAND3_X1   g02405(.A1(new_n2451_), .A2(new_n2029_), .A3(new_n2449_), .ZN(new_n2475_));
  NAND3_X1   g02406(.A1(new_n2475_), .A2(new_n2341_), .A3(new_n2448_), .ZN(new_n2476_));
  XOR2_X1    g02407(.A1(new_n2342_), .A2(new_n2445_), .Z(new_n2477_));
  NOR2_X1    g02408(.A1(new_n2477_), .A2(new_n806_), .ZN(new_n2478_));
  AOI21_X1   g02409(.A1(new_n2028_), .A2(new_n2025_), .B(new_n294_), .ZN(new_n2479_));
  NOR3_X1    g02410(.A1(new_n2459_), .A2(new_n2479_), .A3(new_n2478_), .ZN(new_n2480_));
  OAI21_X1   g02411(.A1(new_n2480_), .A2(new_n2354_), .B(new_n2441_), .ZN(new_n2481_));
  NAND2_X1   g02412(.A1(new_n2481_), .A2(new_n2476_), .ZN(new_n2482_));
  AOI21_X1   g02413(.A1(new_n2482_), .A2(new_n2474_), .B(new_n2470_), .ZN(new_n2483_));
  AOI21_X1   g02414(.A1(new_n2096_), .A2(new_n2099_), .B(new_n806_), .ZN(new_n2484_));
  NAND2_X1   g02415(.A1(new_n2336_), .A2(new_n2484_), .ZN(new_n2485_));
  NOR2_X1    g02416(.A1(new_n2336_), .A2(new_n2484_), .ZN(new_n2486_));
  INV_X1     g02417(.I(new_n2486_), .ZN(new_n2487_));
  AOI21_X1   g02418(.A1(new_n2487_), .A2(new_n2485_), .B(new_n2435_), .ZN(new_n2488_));
  NOR3_X1    g02419(.A1(new_n2100_), .A2(new_n2438_), .A3(new_n806_), .ZN(new_n2489_));
  NOR3_X1    g02420(.A1(new_n2489_), .A2(new_n2486_), .A3(new_n2331_), .ZN(new_n2490_));
  NOR2_X1    g02421(.A1(new_n2488_), .A2(new_n2490_), .ZN(new_n2491_));
  INV_X1     g02422(.I(\a[6] ), .ZN(new_n2492_));
  NOR2_X1    g02423(.A1(new_n2492_), .A2(\a[8] ), .ZN(new_n2493_));
  NOR2_X1    g02424(.A1(new_n498_), .A2(\a[6] ), .ZN(new_n2494_));
  OAI22_X1   g02425(.A1(new_n2493_), .A2(new_n2494_), .B1(new_n2466_), .B2(new_n2467_), .ZN(new_n2495_));
  NOR2_X1    g02426(.A1(new_n2495_), .A2(new_n498_), .ZN(new_n2496_));
  XOR2_X1    g02427(.A1(new_n2428_), .A2(new_n2323_), .Z(new_n2497_));
  NAND3_X1   g02428(.A1(new_n2334_), .A2(new_n2331_), .A3(new_n2326_), .ZN(new_n2498_));
  NAND3_X1   g02429(.A1(new_n2498_), .A2(new_n2428_), .A3(new_n2323_), .ZN(new_n2499_));
  NOR3_X1    g02430(.A1(new_n2436_), .A2(new_n2435_), .A3(new_n2434_), .ZN(new_n2500_));
  OAI21_X1   g02431(.A1(new_n2500_), .A2(new_n2431_), .B(new_n2300_), .ZN(new_n2501_));
  NAND2_X1   g02432(.A1(new_n2501_), .A2(new_n2499_), .ZN(new_n2502_));
  OAI21_X1   g02433(.A1(new_n2497_), .A2(new_n2502_), .B(new_n2496_), .ZN(new_n2503_));
  NOR2_X1    g02434(.A1(new_n2109_), .A2(new_n1079_), .ZN(new_n2504_));
  NAND2_X1   g02435(.A1(new_n2504_), .A2(new_n2426_), .ZN(new_n2505_));
  INV_X1     g02436(.I(new_n2505_), .ZN(new_n2506_));
  NOR2_X1    g02437(.A1(new_n2504_), .A2(new_n2426_), .ZN(new_n2507_));
  OAI21_X1   g02438(.A1(new_n2506_), .A2(new_n2507_), .B(new_n2297_), .ZN(new_n2508_));
  INV_X1     g02439(.I(new_n2297_), .ZN(new_n2509_));
  INV_X1     g02440(.I(new_n2507_), .ZN(new_n2510_));
  NAND3_X1   g02441(.A1(new_n2510_), .A2(new_n2509_), .A3(new_n2505_), .ZN(new_n2511_));
  NAND2_X1   g02442(.A1(new_n2508_), .A2(new_n2511_), .ZN(new_n2512_));
  NAND3_X1   g02443(.A1(new_n2284_), .A2(new_n2416_), .A3(new_n1079_), .ZN(new_n2513_));
  OAI21_X1   g02444(.A1(new_n2130_), .A2(new_n806_), .B(new_n2417_), .ZN(new_n2514_));
  AOI21_X1   g02445(.A1(new_n2514_), .A2(new_n2513_), .B(new_n2279_), .ZN(new_n2515_));
  NOR3_X1    g02446(.A1(new_n2130_), .A2(new_n2417_), .A3(new_n806_), .ZN(new_n2516_));
  AOI21_X1   g02447(.A1(new_n1079_), .A2(new_n2416_), .B(new_n2284_), .ZN(new_n2517_));
  NOR3_X1    g02448(.A1(new_n2517_), .A2(new_n2516_), .A3(new_n2419_), .ZN(new_n2518_));
  NOR2_X1    g02449(.A1(new_n2518_), .A2(new_n2515_), .ZN(new_n2519_));
  NAND2_X1   g02450(.A1(new_n2272_), .A2(new_n2268_), .ZN(new_n2520_));
  NAND2_X1   g02451(.A1(new_n2520_), .A2(new_n2255_), .ZN(new_n2521_));
  AND2_X2    g02452(.A1(new_n2272_), .A2(new_n2268_), .Z(new_n2522_));
  NAND2_X1   g02453(.A1(new_n2256_), .A2(new_n2522_), .ZN(new_n2523_));
  NAND2_X1   g02454(.A1(new_n2523_), .A2(new_n2521_), .ZN(new_n2524_));
  INV_X1     g02455(.I(new_n2524_), .ZN(new_n2525_));
  INV_X1     g02456(.I(new_n2268_), .ZN(new_n2526_));
  NOR3_X1    g02457(.A1(new_n2281_), .A2(new_n2279_), .A3(new_n2526_), .ZN(new_n2527_));
  NOR3_X1    g02458(.A1(new_n2527_), .A2(new_n2522_), .A3(new_n2256_), .ZN(new_n2528_));
  OAI21_X1   g02459(.A1(new_n2278_), .A2(new_n2273_), .B(new_n806_), .ZN(new_n2529_));
  NAND3_X1   g02460(.A1(new_n2419_), .A2(new_n2529_), .A3(new_n2268_), .ZN(new_n2530_));
  AOI21_X1   g02461(.A1(new_n2530_), .A2(new_n2520_), .B(new_n2255_), .ZN(new_n2531_));
  NOR2_X1    g02462(.A1(new_n2528_), .A2(new_n2531_), .ZN(new_n2532_));
  OAI21_X1   g02463(.A1(new_n2525_), .A2(new_n2532_), .B(new_n2496_), .ZN(new_n2533_));
  NAND3_X1   g02464(.A1(new_n2220_), .A2(new_n2218_), .A3(new_n806_), .ZN(new_n2534_));
  NOR2_X1    g02465(.A1(new_n2219_), .A2(new_n1787_), .ZN(new_n2535_));
  NOR2_X1    g02466(.A1(new_n2217_), .A2(new_n1784_), .ZN(new_n2536_));
  OAI21_X1   g02467(.A1(new_n2535_), .A2(new_n2536_), .B(new_n1079_), .ZN(new_n2537_));
  AOI21_X1   g02468(.A1(new_n2534_), .A2(new_n2537_), .B(new_n2215_), .ZN(new_n2538_));
  OAI21_X1   g02469(.A1(new_n2535_), .A2(new_n2536_), .B(new_n806_), .ZN(new_n2539_));
  NAND2_X1   g02470(.A1(new_n2539_), .A2(new_n2222_), .ZN(new_n2540_));
  AOI21_X1   g02471(.A1(new_n2215_), .A2(new_n2540_), .B(new_n2538_), .ZN(new_n2541_));
  OAI21_X1   g02472(.A1(new_n2137_), .A2(new_n2132_), .B(new_n2136_), .ZN(new_n2542_));
  NAND3_X1   g02473(.A1(new_n2133_), .A2(new_n2131_), .A3(new_n2134_), .ZN(new_n2543_));
  AOI21_X1   g02474(.A1(new_n2542_), .A2(new_n2543_), .B(new_n1079_), .ZN(new_n2544_));
  NAND2_X1   g02475(.A1(new_n2197_), .A2(new_n2544_), .ZN(new_n2545_));
  NOR2_X1    g02476(.A1(new_n2174_), .A2(new_n2168_), .ZN(new_n2546_));
  AOI21_X1   g02477(.A1(new_n2183_), .A2(new_n2184_), .B(new_n806_), .ZN(new_n2547_));
  OAI21_X1   g02478(.A1(new_n2546_), .A2(new_n2547_), .B(new_n2185_), .ZN(new_n2548_));
  NOR3_X1    g02479(.A1(new_n2194_), .A2(new_n2195_), .A3(new_n1079_), .ZN(new_n2549_));
  NOR3_X1    g02480(.A1(new_n2548_), .A2(new_n2549_), .A3(new_n2199_), .ZN(new_n2550_));
  OAI21_X1   g02481(.A1(new_n2138_), .A2(new_n2135_), .B(new_n806_), .ZN(new_n2551_));
  NAND2_X1   g02482(.A1(new_n2550_), .A2(new_n2551_), .ZN(new_n2552_));
  AOI21_X1   g02483(.A1(new_n2552_), .A2(new_n2545_), .B(new_n2199_), .ZN(new_n2553_));
  NOR2_X1    g02484(.A1(new_n2550_), .A2(new_n2551_), .ZN(new_n2554_));
  NOR2_X1    g02485(.A1(new_n2197_), .A2(new_n2544_), .ZN(new_n2555_));
  NOR3_X1    g02486(.A1(new_n2554_), .A2(new_n2555_), .A3(new_n2196_), .ZN(new_n2556_));
  NOR2_X1    g02487(.A1(new_n2556_), .A2(new_n2553_), .ZN(new_n2557_));
  NAND2_X1   g02488(.A1(new_n2165_), .A2(new_n2161_), .ZN(new_n2558_));
  NOR2_X1    g02489(.A1(new_n2558_), .A2(new_n806_), .ZN(new_n2559_));
  NAND2_X1   g02490(.A1(new_n2143_), .A2(new_n2144_), .ZN(new_n2560_));
  NAND3_X1   g02491(.A1(new_n2560_), .A2(new_n1079_), .A3(new_n2167_), .ZN(new_n2561_));
  NOR3_X1    g02492(.A1(new_n643_), .A2(new_n2046_), .A3(new_n279_), .ZN(new_n2562_));
  NOR2_X1    g02493(.A1(new_n644_), .A2(new_n1734_), .ZN(new_n2563_));
  OAI21_X1   g02494(.A1(new_n2563_), .A2(new_n2562_), .B(new_n806_), .ZN(new_n2564_));
  NOR2_X1    g02495(.A1(new_n2155_), .A2(new_n2153_), .ZN(new_n2565_));
  NOR2_X1    g02496(.A1(new_n2565_), .A2(new_n2564_), .ZN(new_n2566_));
  OAI21_X1   g02497(.A1(new_n2172_), .A2(new_n806_), .B(new_n2566_), .ZN(new_n2567_));
  AOI21_X1   g02498(.A1(new_n2561_), .A2(new_n2567_), .B(new_n2559_), .ZN(new_n2568_));
  NOR3_X1    g02499(.A1(new_n2172_), .A2(new_n806_), .A3(new_n2566_), .ZN(new_n2569_));
  AOI21_X1   g02500(.A1(new_n2560_), .A2(new_n1079_), .B(new_n2167_), .ZN(new_n2570_));
  NOR4_X1    g02501(.A1(new_n2570_), .A2(new_n2569_), .A3(new_n806_), .A4(new_n2558_), .ZN(new_n2571_));
  NOR2_X1    g02502(.A1(new_n2571_), .A2(new_n2568_), .ZN(new_n2572_));
  XNOR2_X1   g02503(.A1(\a[8] ), .A2(\a[9] ), .ZN(new_n2573_));
  NAND2_X1   g02504(.A1(new_n2573_), .A2(\a[11] ), .ZN(new_n2574_));
  NOR4_X1    g02505(.A1(new_n1079_), .A2(new_n279_), .A3(new_n785_), .A4(new_n2045_), .ZN(new_n2576_));
  INV_X1     g02506(.I(new_n2576_), .ZN(new_n2577_));
  NAND4_X1   g02507(.A1(new_n2146_), .A2(new_n806_), .A3(new_n2045_), .A4(new_n2145_), .ZN(new_n2578_));
  AOI21_X1   g02508(.A1(new_n2578_), .A2(new_n2577_), .B(new_n2150_), .ZN(new_n2579_));
  NOR4_X1    g02509(.A1(new_n2563_), .A2(new_n1079_), .A3(new_n1733_), .A4(new_n2562_), .ZN(new_n2580_));
  NOR4_X1    g02510(.A1(new_n2580_), .A2(new_n1733_), .A3(new_n2149_), .A4(new_n2576_), .ZN(new_n2581_));
  NOR2_X1    g02511(.A1(new_n2581_), .A2(new_n2579_), .ZN(new_n2582_));
  XNOR2_X1   g02512(.A1(\a[5] ), .A2(\a[6] ), .ZN(new_n2583_));
  NAND2_X1   g02513(.A1(new_n2583_), .A2(\a[8] ), .ZN(new_n2584_));
  NOR2_X1    g02514(.A1(new_n2470_), .A2(new_n2584_), .ZN(new_n2585_));
  NAND3_X1   g02515(.A1(new_n2469_), .A2(\a[8] ), .A3(new_n1075_), .ZN(new_n2586_));
  INV_X1     g02516(.I(new_n2586_), .ZN(new_n2587_));
  NOR3_X1    g02517(.A1(new_n1079_), .A2(new_n2496_), .A3(new_n2574_), .ZN(new_n2588_));
  NOR3_X1    g02518(.A1(new_n1078_), .A2(new_n294_), .A3(new_n2573_), .ZN(new_n2589_));
  NOR2_X1    g02519(.A1(new_n2470_), .A2(new_n2589_), .ZN(new_n2590_));
  NOR2_X1    g02520(.A1(new_n2590_), .A2(new_n2588_), .ZN(new_n2591_));
  NOR2_X1    g02521(.A1(new_n1079_), .A2(new_n1733_), .ZN(new_n2592_));
  NOR2_X1    g02522(.A1(new_n2150_), .A2(new_n2148_), .ZN(new_n2593_));
  NOR2_X1    g02523(.A1(new_n806_), .A2(new_n2593_), .ZN(new_n2594_));
  NOR3_X1    g02524(.A1(new_n2594_), .A2(new_n2592_), .A3(new_n2496_), .ZN(new_n2595_));
  OAI21_X1   g02525(.A1(new_n2594_), .A2(new_n2592_), .B(new_n2496_), .ZN(new_n2596_));
  INV_X1     g02526(.I(new_n2596_), .ZN(new_n2597_));
  OAI21_X1   g02527(.A1(new_n2597_), .A2(new_n2595_), .B(new_n2591_), .ZN(new_n2598_));
  NOR2_X1    g02528(.A1(new_n2582_), .A2(new_n2598_), .ZN(new_n2599_));
  NOR2_X1    g02529(.A1(new_n2594_), .A2(new_n2592_), .ZN(new_n2600_));
  NAND2_X1   g02530(.A1(new_n2600_), .A2(new_n2496_), .ZN(new_n2601_));
  AOI21_X1   g02531(.A1(new_n2582_), .A2(new_n2598_), .B(new_n2601_), .ZN(new_n2602_));
  NOR2_X1    g02532(.A1(new_n2155_), .A2(new_n2153_), .ZN(new_n2603_));
  XOR2_X1    g02533(.A1(new_n2603_), .A2(new_n2564_), .Z(new_n2604_));
  NAND2_X1   g02534(.A1(new_n2604_), .A2(new_n2496_), .ZN(new_n2605_));
  OAI21_X1   g02535(.A1(new_n2602_), .A2(new_n2599_), .B(new_n2605_), .ZN(new_n2606_));
  XOR2_X1    g02536(.A1(new_n2603_), .A2(new_n2151_), .Z(new_n2607_));
  NAND2_X1   g02537(.A1(new_n2607_), .A2(new_n2470_), .ZN(new_n2608_));
  INV_X1     g02538(.I(new_n2603_), .ZN(new_n2609_));
  INV_X1     g02539(.I(new_n2153_), .ZN(new_n2610_));
  NAND3_X1   g02540(.A1(new_n2165_), .A2(new_n806_), .A3(new_n2161_), .ZN(new_n2611_));
  OAI21_X1   g02541(.A1(new_n2159_), .A2(new_n2156_), .B(new_n1079_), .ZN(new_n2612_));
  NAND3_X1   g02542(.A1(new_n2612_), .A2(new_n2611_), .A3(new_n2610_), .ZN(new_n2613_));
  NAND3_X1   g02543(.A1(new_n2613_), .A2(new_n2564_), .A3(new_n2609_), .ZN(new_n2614_));
  NOR3_X1    g02544(.A1(new_n2160_), .A2(new_n2166_), .A3(new_n2153_), .ZN(new_n2615_));
  OAI21_X1   g02545(.A1(new_n2615_), .A2(new_n2603_), .B(new_n2151_), .ZN(new_n2616_));
  NAND3_X1   g02546(.A1(new_n2616_), .A2(new_n2614_), .A3(new_n2470_), .ZN(new_n2617_));
  NOR3_X1    g02547(.A1(new_n2615_), .A2(new_n2151_), .A3(new_n2603_), .ZN(new_n2618_));
  AOI21_X1   g02548(.A1(new_n2613_), .A2(new_n2609_), .B(new_n2564_), .ZN(new_n2619_));
  OAI21_X1   g02549(.A1(new_n2618_), .A2(new_n2619_), .B(new_n2496_), .ZN(new_n2620_));
  NAND4_X1   g02550(.A1(new_n2620_), .A2(new_n2617_), .A3(new_n2606_), .A4(new_n2608_), .ZN(new_n2621_));
  NOR2_X1    g02551(.A1(new_n2621_), .A2(new_n2572_), .ZN(new_n2622_));
  AOI21_X1   g02552(.A1(new_n2616_), .A2(new_n2614_), .B(new_n2470_), .ZN(new_n2623_));
  NAND2_X1   g02553(.A1(new_n2623_), .A2(new_n2470_), .ZN(new_n2624_));
  AOI21_X1   g02554(.A1(new_n2621_), .A2(new_n2572_), .B(new_n2624_), .ZN(new_n2625_));
  NAND2_X1   g02555(.A1(new_n2560_), .A2(new_n2566_), .ZN(new_n2626_));
  INV_X1     g02556(.I(new_n2173_), .ZN(new_n2627_));
  OAI21_X1   g02557(.A1(new_n2560_), .A2(new_n2566_), .B(new_n2627_), .ZN(new_n2628_));
  NAND2_X1   g02558(.A1(new_n2628_), .A2(new_n2626_), .ZN(new_n2629_));
  NAND2_X1   g02559(.A1(new_n2181_), .A2(new_n2185_), .ZN(new_n2630_));
  NAND2_X1   g02560(.A1(new_n2630_), .A2(new_n2629_), .ZN(new_n2631_));
  NAND3_X1   g02561(.A1(new_n2183_), .A2(new_n2184_), .A3(new_n1079_), .ZN(new_n2632_));
  OAI21_X1   g02562(.A1(new_n2180_), .A2(new_n2178_), .B(new_n806_), .ZN(new_n2633_));
  AND2_X2    g02563(.A1(new_n2633_), .A2(new_n2632_), .Z(new_n2634_));
  OAI21_X1   g02564(.A1(new_n2634_), .A2(new_n2629_), .B(new_n2631_), .ZN(new_n2635_));
  OAI21_X1   g02565(.A1(new_n2625_), .A2(new_n2622_), .B(new_n2635_), .ZN(new_n2636_));
  OR2_X2     g02566(.A1(new_n2571_), .A2(new_n2568_), .Z(new_n2637_));
  OAI22_X1   g02567(.A1(new_n2580_), .A2(new_n2576_), .B1(new_n1733_), .B2(new_n2149_), .ZN(new_n2638_));
  NAND3_X1   g02568(.A1(new_n2578_), .A2(new_n2150_), .A3(new_n2577_), .ZN(new_n2639_));
  NAND2_X1   g02569(.A1(new_n2638_), .A2(new_n2639_), .ZN(new_n2640_));
  INV_X1     g02570(.I(new_n2574_), .ZN(new_n2641_));
  NAND3_X1   g02571(.A1(new_n806_), .A2(new_n2470_), .A3(new_n2641_), .ZN(new_n2642_));
  OAI21_X1   g02572(.A1(new_n806_), .A2(new_n2641_), .B(new_n2496_), .ZN(new_n2643_));
  NAND2_X1   g02573(.A1(new_n2642_), .A2(new_n2643_), .ZN(new_n2644_));
  INV_X1     g02574(.I(new_n2595_), .ZN(new_n2645_));
  AOI21_X1   g02575(.A1(new_n2645_), .A2(new_n2596_), .B(new_n2644_), .ZN(new_n2646_));
  NAND2_X1   g02576(.A1(new_n2640_), .A2(new_n2646_), .ZN(new_n2647_));
  INV_X1     g02577(.I(new_n2601_), .ZN(new_n2648_));
  OAI21_X1   g02578(.A1(new_n2640_), .A2(new_n2646_), .B(new_n2648_), .ZN(new_n2649_));
  NOR2_X1    g02579(.A1(new_n2607_), .A2(new_n2470_), .ZN(new_n2650_));
  AOI21_X1   g02580(.A1(new_n2649_), .A2(new_n2647_), .B(new_n2650_), .ZN(new_n2651_));
  INV_X1     g02581(.I(new_n2608_), .ZN(new_n2652_));
  NOR3_X1    g02582(.A1(new_n2618_), .A2(new_n2619_), .A3(new_n2496_), .ZN(new_n2653_));
  NOR4_X1    g02583(.A1(new_n2653_), .A2(new_n2623_), .A3(new_n2651_), .A4(new_n2652_), .ZN(new_n2654_));
  NAND2_X1   g02584(.A1(new_n2654_), .A2(new_n2637_), .ZN(new_n2655_));
  NOR2_X1    g02585(.A1(new_n2620_), .A2(new_n2496_), .ZN(new_n2656_));
  OAI21_X1   g02586(.A1(new_n2654_), .A2(new_n2637_), .B(new_n2656_), .ZN(new_n2657_));
  NOR2_X1    g02587(.A1(new_n2634_), .A2(new_n2629_), .ZN(new_n2658_));
  AOI21_X1   g02588(.A1(new_n2630_), .A2(new_n2629_), .B(new_n2658_), .ZN(new_n2659_));
  NAND3_X1   g02589(.A1(new_n2657_), .A2(new_n2655_), .A3(new_n2659_), .ZN(new_n2660_));
  NAND2_X1   g02590(.A1(new_n2660_), .A2(\a[8] ), .ZN(new_n2661_));
  AOI22_X1   g02591(.A1(new_n2196_), .A2(new_n2193_), .B1(new_n2182_), .B2(new_n2185_), .ZN(new_n2662_));
  NOR3_X1    g02592(.A1(new_n2550_), .A2(new_n2662_), .A3(new_n2470_), .ZN(new_n2663_));
  OAI21_X1   g02593(.A1(new_n2549_), .A2(new_n2199_), .B(new_n2548_), .ZN(new_n2664_));
  AOI21_X1   g02594(.A1(new_n2664_), .A2(new_n2197_), .B(new_n2496_), .ZN(new_n2665_));
  NOR2_X1    g02595(.A1(new_n2665_), .A2(new_n2663_), .ZN(new_n2666_));
  NAND3_X1   g02596(.A1(new_n2661_), .A2(new_n2636_), .A3(new_n2666_), .ZN(new_n2667_));
  NOR2_X1    g02597(.A1(new_n2667_), .A2(new_n2557_), .ZN(new_n2668_));
  NAND3_X1   g02598(.A1(new_n2664_), .A2(new_n2197_), .A3(new_n2496_), .ZN(new_n2669_));
  NOR2_X1    g02599(.A1(new_n2669_), .A2(new_n2470_), .ZN(new_n2670_));
  INV_X1     g02600(.I(new_n2670_), .ZN(new_n2671_));
  AOI21_X1   g02601(.A1(new_n2667_), .A2(new_n2557_), .B(new_n2671_), .ZN(new_n2672_));
  INV_X1     g02602(.I(new_n2207_), .ZN(new_n2673_));
  NOR3_X1    g02603(.A1(new_n2201_), .A2(new_n2198_), .A3(new_n2673_), .ZN(new_n2674_));
  INV_X1     g02604(.I(new_n2674_), .ZN(new_n2675_));
  OAI21_X1   g02605(.A1(new_n2201_), .A2(new_n2198_), .B(new_n2673_), .ZN(new_n2676_));
  AOI21_X1   g02606(.A1(new_n2675_), .A2(new_n2676_), .B(\a[11] ), .ZN(new_n2677_));
  INV_X1     g02607(.I(new_n2676_), .ZN(new_n2678_));
  NOR3_X1    g02608(.A1(new_n2678_), .A2(new_n2674_), .A3(new_n294_), .ZN(new_n2679_));
  OAI21_X1   g02609(.A1(new_n2677_), .A2(new_n2679_), .B(new_n2496_), .ZN(new_n2680_));
  OAI21_X1   g02610(.A1(new_n2672_), .A2(new_n2668_), .B(new_n2680_), .ZN(new_n2681_));
  NOR3_X1    g02611(.A1(new_n2677_), .A2(new_n2679_), .A3(new_n2496_), .ZN(new_n2682_));
  INV_X1     g02612(.I(new_n2682_), .ZN(new_n2683_));
  XOR2_X1    g02613(.A1(new_n2212_), .A2(new_n1079_), .Z(new_n2684_));
  NAND2_X1   g02614(.A1(new_n2210_), .A2(new_n2684_), .ZN(new_n2685_));
  NAND2_X1   g02615(.A1(new_n2542_), .A2(new_n2543_), .ZN(new_n2686_));
  NAND2_X1   g02616(.A1(new_n2550_), .A2(new_n2686_), .ZN(new_n2687_));
  NOR2_X1    g02617(.A1(new_n2196_), .A2(new_n1079_), .ZN(new_n2688_));
  OAI21_X1   g02618(.A1(new_n2550_), .A2(new_n2686_), .B(new_n2688_), .ZN(new_n2689_));
  NAND3_X1   g02619(.A1(new_n2689_), .A2(new_n2687_), .A3(new_n2673_), .ZN(new_n2690_));
  NAND2_X1   g02620(.A1(new_n2690_), .A2(\a[11] ), .ZN(new_n2691_));
  INV_X1     g02621(.I(new_n2214_), .ZN(new_n2692_));
  NAND2_X1   g02622(.A1(new_n2692_), .A2(new_n2213_), .ZN(new_n2693_));
  NAND3_X1   g02623(.A1(new_n2691_), .A2(new_n2693_), .A3(new_n2208_), .ZN(new_n2694_));
  NAND3_X1   g02624(.A1(new_n2685_), .A2(new_n2694_), .A3(new_n2470_), .ZN(new_n2695_));
  XOR2_X1    g02625(.A1(new_n2212_), .A2(new_n806_), .Z(new_n2696_));
  AOI21_X1   g02626(.A1(new_n2691_), .A2(new_n2208_), .B(new_n2696_), .ZN(new_n2697_));
  INV_X1     g02627(.I(new_n2213_), .ZN(new_n2698_));
  NOR2_X1    g02628(.A1(new_n2698_), .A2(new_n2214_), .ZN(new_n2699_));
  NOR2_X1    g02629(.A1(new_n2210_), .A2(new_n2699_), .ZN(new_n2700_));
  OAI21_X1   g02630(.A1(new_n2700_), .A2(new_n2697_), .B(new_n2496_), .ZN(new_n2701_));
  NAND4_X1   g02631(.A1(new_n2681_), .A2(new_n2683_), .A3(new_n2695_), .A4(new_n2701_), .ZN(new_n2702_));
  NOR2_X1    g02632(.A1(new_n2702_), .A2(new_n2541_), .ZN(new_n2703_));
  NOR2_X1    g02633(.A1(new_n2701_), .A2(new_n2496_), .ZN(new_n2704_));
  INV_X1     g02634(.I(new_n2704_), .ZN(new_n2705_));
  AOI21_X1   g02635(.A1(new_n2702_), .A2(new_n2541_), .B(new_n2705_), .ZN(new_n2706_));
  OAI21_X1   g02636(.A1(new_n2228_), .A2(new_n2225_), .B(new_n279_), .ZN(new_n2707_));
  NAND3_X1   g02637(.A1(new_n2226_), .A2(\a[14] ), .A3(new_n2224_), .ZN(new_n2708_));
  AOI21_X1   g02638(.A1(new_n2707_), .A2(new_n2708_), .B(new_n806_), .ZN(new_n2709_));
  OAI21_X1   g02639(.A1(new_n2709_), .A2(new_n2231_), .B(new_n2223_), .ZN(new_n2710_));
  AOI21_X1   g02640(.A1(new_n2691_), .A2(new_n2208_), .B(new_n2698_), .ZN(new_n2711_));
  OAI21_X1   g02641(.A1(new_n2711_), .A2(new_n2214_), .B(new_n2539_), .ZN(new_n2712_));
  NAND3_X1   g02642(.A1(new_n2707_), .A2(new_n2708_), .A3(new_n1079_), .ZN(new_n2713_));
  OAI21_X1   g02643(.A1(new_n2227_), .A2(new_n2229_), .B(new_n806_), .ZN(new_n2714_));
  NAND2_X1   g02644(.A1(new_n2714_), .A2(new_n2713_), .ZN(new_n2715_));
  NAND3_X1   g02645(.A1(new_n2712_), .A2(new_n2715_), .A3(new_n2222_), .ZN(new_n2716_));
  NOR3_X1    g02646(.A1(new_n2465_), .A2(\a[5] ), .A3(\a[6] ), .ZN(new_n2717_));
  AOI21_X1   g02647(.A1(\a[6] ), .A2(new_n2467_), .B(new_n2717_), .ZN(new_n2718_));
  NOR2_X1    g02648(.A1(new_n2495_), .A2(new_n2718_), .ZN(new_n2719_));
  XOR2_X1    g02649(.A1(new_n2719_), .A2(new_n498_), .Z(new_n2720_));
  NAND3_X1   g02650(.A1(new_n2716_), .A2(new_n2710_), .A3(new_n2720_), .ZN(new_n2721_));
  OAI21_X1   g02651(.A1(new_n2706_), .A2(new_n2703_), .B(new_n2721_), .ZN(new_n2722_));
  AOI21_X1   g02652(.A1(new_n2716_), .A2(new_n2710_), .B(new_n2720_), .ZN(new_n2723_));
  INV_X1     g02653(.I(new_n2723_), .ZN(new_n2724_));
  INV_X1     g02654(.I(new_n2240_), .ZN(new_n2725_));
  AOI21_X1   g02655(.A1(new_n2725_), .A2(new_n2241_), .B(new_n2232_), .ZN(new_n2726_));
  AOI21_X1   g02656(.A1(new_n2712_), .A2(new_n2222_), .B(new_n2709_), .ZN(new_n2727_));
  NAND3_X1   g02657(.A1(new_n2236_), .A2(new_n2239_), .A3(new_n1079_), .ZN(new_n2728_));
  INV_X1     g02658(.I(new_n2728_), .ZN(new_n2729_));
  AOI21_X1   g02659(.A1(new_n2236_), .A2(new_n2239_), .B(new_n1079_), .ZN(new_n2730_));
  NOR2_X1    g02660(.A1(new_n2729_), .A2(new_n2730_), .ZN(new_n2731_));
  NOR3_X1    g02661(.A1(new_n2731_), .A2(new_n2727_), .A3(new_n2231_), .ZN(new_n2732_));
  NOR3_X1    g02662(.A1(new_n2726_), .A2(new_n2732_), .A3(new_n2470_), .ZN(new_n2733_));
  AOI21_X1   g02663(.A1(new_n2722_), .A2(new_n2724_), .B(new_n2733_), .ZN(new_n2734_));
  INV_X1     g02664(.I(new_n2241_), .ZN(new_n2735_));
  OAI22_X1   g02665(.A1(new_n2727_), .A2(new_n2231_), .B1(new_n2735_), .B2(new_n2240_), .ZN(new_n2736_));
  NOR2_X1    g02666(.A1(new_n2237_), .A2(new_n2234_), .ZN(new_n2737_));
  INV_X1     g02667(.I(new_n2239_), .ZN(new_n2738_));
  OAI21_X1   g02668(.A1(new_n2738_), .A2(new_n2737_), .B(new_n806_), .ZN(new_n2739_));
  NAND2_X1   g02669(.A1(new_n2739_), .A2(new_n2728_), .ZN(new_n2740_));
  NAND2_X1   g02670(.A1(new_n2740_), .A2(new_n2232_), .ZN(new_n2741_));
  AOI21_X1   g02671(.A1(new_n2736_), .A2(new_n2741_), .B(new_n2496_), .ZN(new_n2742_));
  NOR2_X1    g02672(.A1(new_n2734_), .A2(new_n2742_), .ZN(new_n2743_));
  NAND3_X1   g02673(.A1(new_n2252_), .A2(new_n1079_), .A3(new_n2247_), .ZN(new_n2744_));
  OAI21_X1   g02674(.A1(new_n2248_), .A2(new_n2249_), .B(new_n806_), .ZN(new_n2745_));
  NAND2_X1   g02675(.A1(new_n2745_), .A2(new_n2744_), .ZN(new_n2746_));
  NAND2_X1   g02676(.A1(new_n2746_), .A2(new_n2242_), .ZN(new_n2747_));
  OAI21_X1   g02677(.A1(new_n2727_), .A2(new_n2231_), .B(new_n2725_), .ZN(new_n2748_));
  NAND2_X1   g02678(.A1(new_n2250_), .A2(new_n2253_), .ZN(new_n2749_));
  NAND3_X1   g02679(.A1(new_n2749_), .A2(new_n2748_), .A3(new_n2241_), .ZN(new_n2750_));
  AOI21_X1   g02680(.A1(new_n2750_), .A2(new_n2747_), .B(new_n2496_), .ZN(new_n2751_));
  NAND3_X1   g02681(.A1(new_n2750_), .A2(new_n2747_), .A3(new_n2496_), .ZN(new_n2752_));
  OAI21_X1   g02682(.A1(new_n2743_), .A2(new_n2751_), .B(new_n2752_), .ZN(new_n2753_));
  NAND3_X1   g02683(.A1(new_n2530_), .A2(new_n2255_), .A3(new_n2520_), .ZN(new_n2754_));
  OAI21_X1   g02684(.A1(new_n2527_), .A2(new_n2522_), .B(new_n2256_), .ZN(new_n2755_));
  NAND3_X1   g02685(.A1(new_n2755_), .A2(new_n2754_), .A3(new_n2470_), .ZN(new_n2756_));
  OAI21_X1   g02686(.A1(new_n2528_), .A2(new_n2531_), .B(new_n2496_), .ZN(new_n2757_));
  NAND3_X1   g02687(.A1(new_n2525_), .A2(new_n2757_), .A3(new_n2756_), .ZN(new_n2758_));
  NAND3_X1   g02688(.A1(new_n2758_), .A2(new_n2533_), .A3(new_n2753_), .ZN(new_n2759_));
  NOR2_X1    g02689(.A1(new_n2759_), .A2(new_n2519_), .ZN(new_n2760_));
  NAND2_X1   g02690(.A1(new_n2759_), .A2(new_n2519_), .ZN(new_n2761_));
  NOR2_X1    g02691(.A1(new_n2757_), .A2(new_n2496_), .ZN(new_n2762_));
  AOI21_X1   g02692(.A1(new_n2761_), .A2(new_n2762_), .B(new_n2760_), .ZN(new_n2763_));
  XOR2_X1    g02693(.A1(new_n2117_), .A2(new_n1079_), .Z(new_n2764_));
  NAND3_X1   g02694(.A1(new_n2421_), .A2(new_n2418_), .A3(new_n2719_), .ZN(new_n2765_));
  INV_X1     g02695(.I(new_n2765_), .ZN(new_n2766_));
  AOI21_X1   g02696(.A1(new_n2421_), .A2(new_n2418_), .B(new_n2719_), .ZN(new_n2767_));
  OAI21_X1   g02697(.A1(new_n2766_), .A2(new_n2767_), .B(new_n2764_), .ZN(new_n2768_));
  XOR2_X1    g02698(.A1(new_n2117_), .A2(new_n806_), .Z(new_n2769_));
  INV_X1     g02699(.I(new_n2767_), .ZN(new_n2770_));
  NAND3_X1   g02700(.A1(new_n2770_), .A2(new_n2765_), .A3(new_n2769_), .ZN(new_n2771_));
  AOI21_X1   g02701(.A1(new_n2771_), .A2(new_n2768_), .B(\a[8] ), .ZN(new_n2772_));
  AOI21_X1   g02702(.A1(new_n2770_), .A2(new_n2765_), .B(new_n2769_), .ZN(new_n2773_));
  NOR3_X1    g02703(.A1(new_n2766_), .A2(new_n2764_), .A3(new_n2767_), .ZN(new_n2774_));
  NOR3_X1    g02704(.A1(new_n2773_), .A2(new_n2774_), .A3(new_n498_), .ZN(new_n2775_));
  NOR2_X1    g02705(.A1(new_n2772_), .A2(new_n2775_), .ZN(new_n2776_));
  NAND2_X1   g02706(.A1(new_n2769_), .A2(new_n498_), .ZN(new_n2777_));
  NAND2_X1   g02707(.A1(new_n2764_), .A2(\a[8] ), .ZN(new_n2778_));
  AOI22_X1   g02708(.A1(new_n2778_), .A2(new_n2777_), .B1(new_n2765_), .B2(new_n2770_), .ZN(new_n2779_));
  MUX2_X1    g02709(.I0(new_n2414_), .I1(new_n1079_), .S(new_n2296_), .Z(new_n2780_));
  NOR2_X1    g02710(.A1(new_n2780_), .A2(new_n2422_), .ZN(new_n2781_));
  MUX2_X1    g02711(.I0(new_n2117_), .I1(new_n806_), .S(new_n2296_), .Z(new_n2782_));
  NOR2_X1    g02712(.A1(new_n2782_), .A2(new_n2288_), .ZN(new_n2783_));
  NOR3_X1    g02713(.A1(new_n2781_), .A2(new_n2783_), .A3(new_n2496_), .ZN(new_n2784_));
  NAND2_X1   g02714(.A1(new_n2782_), .A2(new_n2288_), .ZN(new_n2785_));
  NAND2_X1   g02715(.A1(new_n2780_), .A2(new_n2422_), .ZN(new_n2786_));
  AOI21_X1   g02716(.A1(new_n2785_), .A2(new_n2786_), .B(new_n2470_), .ZN(new_n2787_));
  OAI21_X1   g02717(.A1(new_n2787_), .A2(new_n2784_), .B(new_n2779_), .ZN(new_n2788_));
  AOI21_X1   g02718(.A1(new_n2788_), .A2(new_n2776_), .B(new_n2763_), .ZN(new_n2789_));
  NAND2_X1   g02719(.A1(new_n2789_), .A2(new_n2512_), .ZN(new_n2790_));
  OAI21_X1   g02720(.A1(new_n2781_), .A2(new_n2783_), .B(new_n2496_), .ZN(new_n2791_));
  NOR2_X1    g02721(.A1(new_n2791_), .A2(new_n2470_), .ZN(new_n2792_));
  OAI21_X1   g02722(.A1(new_n2789_), .A2(new_n2512_), .B(new_n2792_), .ZN(new_n2793_));
  NAND2_X1   g02723(.A1(new_n2793_), .A2(new_n2790_), .ZN(new_n2794_));
  NAND3_X1   g02724(.A1(new_n2501_), .A2(new_n2499_), .A3(new_n2496_), .ZN(new_n2795_));
  AOI21_X1   g02725(.A1(new_n2501_), .A2(new_n2499_), .B(new_n2496_), .ZN(new_n2796_));
  INV_X1     g02726(.I(new_n2796_), .ZN(new_n2797_));
  NAND3_X1   g02727(.A1(new_n2797_), .A2(new_n2497_), .A3(new_n2795_), .ZN(new_n2798_));
  NAND3_X1   g02728(.A1(new_n2794_), .A2(new_n2798_), .A3(new_n2503_), .ZN(new_n2799_));
  NOR2_X1    g02729(.A1(new_n2799_), .A2(new_n2491_), .ZN(new_n2800_));
  NOR2_X1    g02730(.A1(new_n2797_), .A2(new_n2496_), .ZN(new_n2801_));
  INV_X1     g02731(.I(new_n2801_), .ZN(new_n2802_));
  AOI21_X1   g02732(.A1(new_n2799_), .A2(new_n2491_), .B(new_n2802_), .ZN(new_n2803_));
  NOR2_X1    g02733(.A1(new_n2803_), .A2(new_n2800_), .ZN(new_n2804_));
  NOR3_X1    g02734(.A1(new_n2480_), .A2(new_n2441_), .A3(new_n2354_), .ZN(new_n2805_));
  AOI21_X1   g02735(.A1(new_n2475_), .A2(new_n2448_), .B(new_n2341_), .ZN(new_n2806_));
  NOR3_X1    g02736(.A1(new_n2805_), .A2(new_n2806_), .A3(new_n2496_), .ZN(new_n2807_));
  AOI21_X1   g02737(.A1(new_n2481_), .A2(new_n2476_), .B(new_n2470_), .ZN(new_n2808_));
  NOR3_X1    g02738(.A1(new_n2807_), .A2(new_n2808_), .A3(new_n2474_), .ZN(new_n2809_));
  NOR3_X1    g02739(.A1(new_n2809_), .A2(new_n2804_), .A3(new_n2483_), .ZN(new_n2810_));
  NAND2_X1   g02740(.A1(new_n2810_), .A2(new_n2463_), .ZN(new_n2811_));
  OAI21_X1   g02741(.A1(new_n2805_), .A2(new_n2806_), .B(new_n2496_), .ZN(new_n2812_));
  NOR2_X1    g02742(.A1(new_n2812_), .A2(new_n2470_), .ZN(new_n2813_));
  OAI21_X1   g02743(.A1(new_n2810_), .A2(new_n2463_), .B(new_n2813_), .ZN(new_n2814_));
  NAND2_X1   g02744(.A1(new_n2814_), .A2(new_n2811_), .ZN(new_n2815_));
  NAND2_X1   g02745(.A1(new_n2454_), .A2(new_n2455_), .ZN(new_n2816_));
  NAND2_X1   g02746(.A1(new_n2358_), .A2(new_n2816_), .ZN(new_n2817_));
  NOR2_X1    g02747(.A1(new_n2029_), .A2(new_n1079_), .ZN(new_n2818_));
  OAI21_X1   g02748(.A1(new_n2358_), .A2(new_n2816_), .B(new_n2818_), .ZN(new_n2819_));
  NAND2_X1   g02749(.A1(new_n2819_), .A2(new_n2817_), .ZN(new_n2820_));
  INV_X1     g02750(.I(new_n2820_), .ZN(new_n2821_));
  NAND2_X1   g02751(.A1(new_n2391_), .A2(new_n2392_), .ZN(new_n2822_));
  NAND2_X1   g02752(.A1(new_n2363_), .A2(new_n2822_), .ZN(new_n2823_));
  NOR2_X1    g02753(.A1(new_n2016_), .A2(new_n443_), .ZN(new_n2824_));
  OAI21_X1   g02754(.A1(new_n2363_), .A2(new_n2822_), .B(new_n2824_), .ZN(new_n2825_));
  NAND2_X1   g02755(.A1(new_n2825_), .A2(new_n2823_), .ZN(new_n2826_));
  INV_X1     g02756(.I(new_n2826_), .ZN(new_n2827_));
  NAND2_X1   g02757(.A1(new_n2375_), .A2(new_n2378_), .ZN(new_n2828_));
  NAND2_X1   g02758(.A1(new_n2004_), .A2(new_n2828_), .ZN(new_n2829_));
  NOR2_X1    g02759(.A1(new_n1994_), .A2(new_n273_), .ZN(new_n2830_));
  OAI21_X1   g02760(.A1(new_n2004_), .A2(new_n2828_), .B(new_n2830_), .ZN(new_n2831_));
  NAND2_X1   g02761(.A1(new_n2831_), .A2(new_n2829_), .ZN(new_n2832_));
  INV_X1     g02762(.I(new_n2832_), .ZN(new_n2833_));
  NAND2_X1   g02763(.A1(new_n1981_), .A2(new_n1982_), .ZN(new_n2834_));
  NAND2_X1   g02764(.A1(new_n2372_), .A2(new_n2368_), .ZN(new_n2835_));
  INV_X1     g02765(.I(new_n2835_), .ZN(new_n2836_));
  NOR2_X1    g02766(.A1(new_n2834_), .A2(new_n2836_), .ZN(new_n2837_));
  NAND2_X1   g02767(.A1(new_n1980_), .A2(new_n248_), .ZN(new_n2838_));
  AOI21_X1   g02768(.A1(new_n2834_), .A2(new_n2836_), .B(new_n2838_), .ZN(new_n2839_));
  XOR2_X1    g02769(.A1(new_n1017_), .A2(new_n189_), .Z(new_n2840_));
  NOR2_X1    g02770(.A1(new_n1012_), .A2(new_n2840_), .ZN(new_n2841_));
  NOR2_X1    g02771(.A1(new_n1020_), .A2(new_n1018_), .ZN(new_n2842_));
  NOR3_X1    g02772(.A1(new_n1010_), .A2(new_n1011_), .A3(new_n2842_), .ZN(new_n2843_));
  NOR2_X1    g02773(.A1(new_n2841_), .A2(new_n2843_), .ZN(new_n2844_));
  XOR2_X1    g02774(.A1(new_n2844_), .A2(new_n273_), .Z(new_n2845_));
  OAI21_X1   g02775(.A1(new_n2837_), .A2(new_n2839_), .B(new_n2845_), .ZN(new_n2846_));
  NOR2_X1    g02776(.A1(new_n2839_), .A2(new_n2837_), .ZN(new_n2847_));
  OAI21_X1   g02777(.A1(new_n2841_), .A2(new_n2843_), .B(new_n356_), .ZN(new_n2848_));
  NAND2_X1   g02778(.A1(new_n2844_), .A2(new_n273_), .ZN(new_n2849_));
  NAND2_X1   g02779(.A1(new_n2849_), .A2(new_n2848_), .ZN(new_n2850_));
  NAND2_X1   g02780(.A1(new_n2847_), .A2(new_n2850_), .ZN(new_n2851_));
  NAND2_X1   g02781(.A1(new_n2846_), .A2(new_n2851_), .ZN(new_n2852_));
  INV_X1     g02782(.I(new_n2852_), .ZN(new_n2853_));
  NAND2_X1   g02783(.A1(new_n2853_), .A2(new_n2002_), .ZN(new_n2854_));
  NAND2_X1   g02784(.A1(new_n2852_), .A2(new_n2013_), .ZN(new_n2855_));
  AOI21_X1   g02785(.A1(new_n2854_), .A2(new_n2855_), .B(new_n2833_), .ZN(new_n2856_));
  NOR2_X1    g02786(.A1(new_n2852_), .A2(new_n2002_), .ZN(new_n2857_));
  INV_X1     g02787(.I(new_n2857_), .ZN(new_n2858_));
  NAND2_X1   g02788(.A1(new_n2852_), .A2(new_n2002_), .ZN(new_n2859_));
  AOI21_X1   g02789(.A1(new_n2858_), .A2(new_n2859_), .B(new_n2832_), .ZN(new_n2860_));
  NOR2_X1    g02790(.A1(new_n2860_), .A2(new_n2856_), .ZN(new_n2861_));
  XOR2_X1    g02791(.A1(new_n2861_), .A2(new_n644_), .Z(new_n2862_));
  OAI21_X1   g02792(.A1(new_n2860_), .A2(new_n2856_), .B(new_n644_), .ZN(new_n2863_));
  NAND2_X1   g02793(.A1(new_n2861_), .A2(new_n786_), .ZN(new_n2864_));
  NAND2_X1   g02794(.A1(new_n2864_), .A2(new_n2863_), .ZN(new_n2865_));
  NAND2_X1   g02795(.A1(new_n2827_), .A2(new_n2865_), .ZN(new_n2866_));
  OAI21_X1   g02796(.A1(new_n2827_), .A2(new_n2862_), .B(new_n2866_), .ZN(new_n2867_));
  NAND2_X1   g02797(.A1(new_n2401_), .A2(new_n2399_), .ZN(new_n2868_));
  NAND2_X1   g02798(.A1(new_n2359_), .A2(new_n644_), .ZN(new_n2869_));
  INV_X1     g02799(.I(new_n2869_), .ZN(new_n2870_));
  OAI21_X1   g02800(.A1(new_n2401_), .A2(new_n2399_), .B(new_n2870_), .ZN(new_n2871_));
  NAND3_X1   g02801(.A1(new_n2871_), .A2(new_n2868_), .A3(new_n2259_), .ZN(new_n2872_));
  NOR2_X1    g02802(.A1(new_n2403_), .A2(new_n2402_), .ZN(new_n2873_));
  NOR2_X1    g02803(.A1(new_n2873_), .A2(new_n2025_), .ZN(new_n2874_));
  AOI21_X1   g02804(.A1(new_n2873_), .A2(new_n2025_), .B(new_n2869_), .ZN(new_n2875_));
  OAI21_X1   g02805(.A1(new_n2875_), .A2(new_n2874_), .B(new_n2315_), .ZN(new_n2876_));
  AOI21_X1   g02806(.A1(new_n2872_), .A2(new_n2876_), .B(new_n2867_), .ZN(new_n2877_));
  NAND3_X1   g02807(.A1(new_n2872_), .A2(new_n2876_), .A3(new_n2867_), .ZN(new_n2878_));
  INV_X1     g02808(.I(new_n2878_), .ZN(new_n2879_));
  OAI21_X1   g02809(.A1(new_n2879_), .A2(new_n2877_), .B(new_n294_), .ZN(new_n2880_));
  INV_X1     g02810(.I(new_n2867_), .ZN(new_n2881_));
  NAND2_X1   g02811(.A1(new_n2872_), .A2(new_n2876_), .ZN(new_n2882_));
  NAND2_X1   g02812(.A1(new_n2882_), .A2(new_n2881_), .ZN(new_n2883_));
  NAND3_X1   g02813(.A1(new_n2883_), .A2(\a[11] ), .A3(new_n2878_), .ZN(new_n2884_));
  NAND3_X1   g02814(.A1(new_n2880_), .A2(new_n2884_), .A3(new_n2496_), .ZN(new_n2885_));
  AOI21_X1   g02815(.A1(new_n2883_), .A2(new_n2878_), .B(\a[11] ), .ZN(new_n2886_));
  NOR3_X1    g02816(.A1(new_n2879_), .A2(new_n2877_), .A3(new_n294_), .ZN(new_n2887_));
  OAI21_X1   g02817(.A1(new_n2887_), .A2(new_n2886_), .B(new_n2470_), .ZN(new_n2888_));
  AOI21_X1   g02818(.A1(new_n2888_), .A2(new_n2885_), .B(new_n2821_), .ZN(new_n2889_));
  OAI21_X1   g02819(.A1(new_n2887_), .A2(new_n2886_), .B(new_n2496_), .ZN(new_n2890_));
  NAND3_X1   g02820(.A1(new_n2880_), .A2(new_n2884_), .A3(new_n2470_), .ZN(new_n2891_));
  AOI21_X1   g02821(.A1(new_n2890_), .A2(new_n2891_), .B(new_n2820_), .ZN(new_n2892_));
  XNOR2_X1   g02822(.A1(\a[3] ), .A2(\a[5] ), .ZN(new_n2893_));
  INV_X1     g02823(.I(\a[4] ), .ZN(new_n2894_));
  NOR2_X1    g02824(.A1(new_n2894_), .A2(\a[2] ), .ZN(new_n2895_));
  NOR2_X1    g02825(.A1(new_n451_), .A2(\a[4] ), .ZN(new_n2896_));
  NOR2_X1    g02826(.A1(new_n2895_), .A2(new_n2896_), .ZN(new_n2897_));
  NOR2_X1    g02827(.A1(new_n2897_), .A2(new_n2893_), .ZN(new_n2898_));
  NAND2_X1   g02828(.A1(new_n2898_), .A2(\a[5] ), .ZN(new_n2899_));
  OAI21_X1   g02829(.A1(new_n2889_), .A2(new_n2892_), .B(new_n2899_), .ZN(new_n2900_));
  NOR3_X1    g02830(.A1(new_n2889_), .A2(new_n2892_), .A3(new_n2899_), .ZN(new_n2901_));
  AOI21_X1   g02831(.A1(new_n2815_), .A2(new_n2900_), .B(new_n2901_), .ZN(new_n2902_));
  NOR3_X1    g02832(.A1(new_n2887_), .A2(new_n2886_), .A3(new_n2496_), .ZN(new_n2903_));
  AOI21_X1   g02833(.A1(new_n2820_), .A2(new_n2890_), .B(new_n2903_), .ZN(new_n2904_));
  INV_X1     g02834(.I(new_n2899_), .ZN(new_n2905_));
  NAND2_X1   g02835(.A1(new_n2826_), .A2(new_n2863_), .ZN(new_n2906_));
  NAND2_X1   g02836(.A1(new_n2906_), .A2(new_n2864_), .ZN(new_n2907_));
  AOI21_X1   g02837(.A1(new_n1024_), .A2(new_n1025_), .B(new_n356_), .ZN(new_n2908_));
  XOR2_X1    g02838(.A1(new_n916_), .A2(new_n1022_), .Z(new_n2909_));
  NOR2_X1    g02839(.A1(new_n2909_), .A2(new_n273_), .ZN(new_n2910_));
  NOR2_X1    g02840(.A1(new_n2908_), .A2(new_n2910_), .ZN(new_n2911_));
  OAI21_X1   g02841(.A1(new_n2839_), .A2(new_n2837_), .B(new_n2848_), .ZN(new_n2912_));
  NAND2_X1   g02842(.A1(new_n2912_), .A2(new_n2849_), .ZN(new_n2913_));
  INV_X1     g02843(.I(new_n2913_), .ZN(new_n2914_));
  NAND2_X1   g02844(.A1(new_n2914_), .A2(new_n2911_), .ZN(new_n2915_));
  OAI21_X1   g02845(.A1(new_n2908_), .A2(new_n2910_), .B(new_n2913_), .ZN(new_n2916_));
  NAND2_X1   g02846(.A1(new_n2915_), .A2(new_n2916_), .ZN(new_n2917_));
  NAND2_X1   g02847(.A1(new_n2917_), .A2(new_n568_), .ZN(new_n2918_));
  XOR2_X1    g02848(.A1(new_n2911_), .A2(new_n2913_), .Z(new_n2919_));
  OAI21_X1   g02849(.A1(new_n2919_), .A2(new_n568_), .B(new_n2918_), .ZN(new_n2920_));
  AOI21_X1   g02850(.A1(new_n2832_), .A2(new_n2859_), .B(new_n2857_), .ZN(new_n2921_));
  NAND2_X1   g02851(.A1(new_n2921_), .A2(new_n786_), .ZN(new_n2922_));
  INV_X1     g02852(.I(new_n2922_), .ZN(new_n2923_));
  NOR2_X1    g02853(.A1(new_n2921_), .A2(new_n786_), .ZN(new_n2924_));
  OAI21_X1   g02854(.A1(new_n2923_), .A2(new_n2924_), .B(new_n2920_), .ZN(new_n2925_));
  XOR2_X1    g02855(.A1(new_n2921_), .A2(new_n644_), .Z(new_n2926_));
  OAI21_X1   g02856(.A1(new_n2920_), .A2(new_n2926_), .B(new_n2925_), .ZN(new_n2927_));
  NOR2_X1    g02857(.A1(new_n2907_), .A2(new_n2927_), .ZN(new_n2928_));
  AND2_X2    g02858(.A1(new_n2907_), .A2(new_n2927_), .Z(new_n2929_));
  OAI21_X1   g02859(.A1(new_n2929_), .A2(new_n2928_), .B(new_n806_), .ZN(new_n2930_));
  XNOR2_X1   g02860(.A1(new_n2907_), .A2(new_n2927_), .ZN(new_n2931_));
  OAI21_X1   g02861(.A1(new_n2931_), .A2(new_n806_), .B(new_n2930_), .ZN(new_n2932_));
  INV_X1     g02862(.I(new_n2932_), .ZN(new_n2933_));
  NAND2_X1   g02863(.A1(new_n2871_), .A2(new_n2868_), .ZN(new_n2934_));
  INV_X1     g02864(.I(new_n2934_), .ZN(new_n2935_));
  NOR2_X1    g02865(.A1(new_n2935_), .A2(new_n2881_), .ZN(new_n2936_));
  AOI21_X1   g02866(.A1(new_n2935_), .A2(new_n2881_), .B(new_n2260_), .ZN(new_n2937_));
  NOR2_X1    g02867(.A1(new_n2937_), .A2(new_n2936_), .ZN(new_n2938_));
  NAND2_X1   g02868(.A1(new_n2933_), .A2(new_n2938_), .ZN(new_n2939_));
  OAI21_X1   g02869(.A1(new_n2936_), .A2(new_n2937_), .B(new_n2932_), .ZN(new_n2940_));
  AOI21_X1   g02870(.A1(new_n2939_), .A2(new_n2940_), .B(new_n2496_), .ZN(new_n2941_));
  XOR2_X1    g02871(.A1(new_n2938_), .A2(new_n2932_), .Z(new_n2942_));
  NOR2_X1    g02872(.A1(new_n2942_), .A2(new_n2470_), .ZN(new_n2943_));
  NOR2_X1    g02873(.A1(new_n2943_), .A2(new_n2941_), .ZN(new_n2944_));
  XOR2_X1    g02874(.A1(new_n2944_), .A2(new_n2905_), .Z(new_n2945_));
  NOR3_X1    g02875(.A1(new_n2943_), .A2(new_n2905_), .A3(new_n2941_), .ZN(new_n2946_));
  NOR2_X1    g02876(.A1(new_n2944_), .A2(new_n2899_), .ZN(new_n2947_));
  NOR2_X1    g02877(.A1(new_n2947_), .A2(new_n2946_), .ZN(new_n2948_));
  MUX2_X1    g02878(.I0(new_n2945_), .I1(new_n2948_), .S(new_n2904_), .Z(new_n2949_));
  NOR2_X1    g02879(.A1(new_n2949_), .A2(new_n2902_), .ZN(new_n2950_));
  INV_X1     g02880(.I(new_n2950_), .ZN(new_n2951_));
  MUX2_X1    g02881(.I0(new_n2470_), .I1(new_n2474_), .S(new_n2482_), .Z(new_n2952_));
  XOR2_X1    g02882(.A1(new_n2952_), .A2(new_n2804_), .Z(new_n2953_));
  INV_X1     g02883(.I(new_n2953_), .ZN(new_n2954_));
  OAI21_X1   g02884(.A1(new_n2489_), .A2(new_n2486_), .B(new_n2331_), .ZN(new_n2955_));
  INV_X1     g02885(.I(new_n2490_), .ZN(new_n2956_));
  AOI21_X1   g02886(.A1(new_n2956_), .A2(new_n2955_), .B(new_n2496_), .ZN(new_n2957_));
  NAND2_X1   g02887(.A1(new_n2957_), .A2(new_n2799_), .ZN(new_n2958_));
  OAI21_X1   g02888(.A1(new_n2488_), .A2(new_n2490_), .B(new_n2470_), .ZN(new_n2959_));
  NAND4_X1   g02889(.A1(new_n2959_), .A2(new_n2503_), .A3(new_n2794_), .A4(new_n2798_), .ZN(new_n2960_));
  AOI21_X1   g02890(.A1(new_n2958_), .A2(new_n2960_), .B(new_n2796_), .ZN(new_n2961_));
  INV_X1     g02891(.I(new_n2503_), .ZN(new_n2962_));
  AOI21_X1   g02892(.A1(new_n2510_), .A2(new_n2505_), .B(new_n2509_), .ZN(new_n2963_));
  NOR3_X1    g02893(.A1(new_n2506_), .A2(new_n2297_), .A3(new_n2507_), .ZN(new_n2964_));
  NOR2_X1    g02894(.A1(new_n2963_), .A2(new_n2964_), .ZN(new_n2965_));
  OR2_X2     g02895(.A1(new_n2518_), .A2(new_n2515_), .Z(new_n2966_));
  NAND2_X1   g02896(.A1(new_n2755_), .A2(new_n2754_), .ZN(new_n2967_));
  AOI21_X1   g02897(.A1(new_n2967_), .A2(new_n2524_), .B(new_n2470_), .ZN(new_n2968_));
  INV_X1     g02898(.I(new_n2538_), .ZN(new_n2969_));
  NAND2_X1   g02899(.A1(new_n2540_), .A2(new_n2215_), .ZN(new_n2970_));
  NAND2_X1   g02900(.A1(new_n2969_), .A2(new_n2970_), .ZN(new_n2971_));
  INV_X1     g02901(.I(new_n2557_), .ZN(new_n2972_));
  NOR3_X1    g02902(.A1(new_n2625_), .A2(new_n2622_), .A3(new_n2635_), .ZN(new_n2973_));
  OAI21_X1   g02903(.A1(new_n498_), .A2(new_n2973_), .B(new_n2636_), .ZN(new_n2974_));
  INV_X1     g02904(.I(new_n2666_), .ZN(new_n2975_));
  NOR2_X1    g02905(.A1(new_n2974_), .A2(new_n2975_), .ZN(new_n2976_));
  NAND2_X1   g02906(.A1(new_n2976_), .A2(new_n2972_), .ZN(new_n2977_));
  OAI21_X1   g02907(.A1(new_n2976_), .A2(new_n2972_), .B(new_n2670_), .ZN(new_n2978_));
  OAI21_X1   g02908(.A1(new_n2678_), .A2(new_n2674_), .B(new_n294_), .ZN(new_n2979_));
  NAND3_X1   g02909(.A1(new_n2675_), .A2(\a[11] ), .A3(new_n2676_), .ZN(new_n2980_));
  AOI21_X1   g02910(.A1(new_n2979_), .A2(new_n2980_), .B(new_n2470_), .ZN(new_n2981_));
  AOI21_X1   g02911(.A1(new_n2978_), .A2(new_n2977_), .B(new_n2981_), .ZN(new_n2982_));
  NAND2_X1   g02912(.A1(new_n2701_), .A2(new_n2695_), .ZN(new_n2983_));
  NOR3_X1    g02913(.A1(new_n2982_), .A2(new_n2983_), .A3(new_n2682_), .ZN(new_n2984_));
  NAND2_X1   g02914(.A1(new_n2984_), .A2(new_n2971_), .ZN(new_n2985_));
  OAI21_X1   g02915(.A1(new_n2984_), .A2(new_n2971_), .B(new_n2704_), .ZN(new_n2986_));
  INV_X1     g02916(.I(new_n2710_), .ZN(new_n2987_));
  AOI21_X1   g02917(.A1(new_n2713_), .A2(new_n2714_), .B(new_n2223_), .ZN(new_n2988_));
  INV_X1     g02918(.I(new_n2720_), .ZN(new_n2989_));
  NOR3_X1    g02919(.A1(new_n2987_), .A2(new_n2988_), .A3(new_n2989_), .ZN(new_n2990_));
  AOI21_X1   g02920(.A1(new_n2986_), .A2(new_n2985_), .B(new_n2990_), .ZN(new_n2991_));
  NAND3_X1   g02921(.A1(new_n2736_), .A2(new_n2741_), .A3(new_n2496_), .ZN(new_n2992_));
  OAI21_X1   g02922(.A1(new_n2991_), .A2(new_n2723_), .B(new_n2992_), .ZN(new_n2993_));
  OAI21_X1   g02923(.A1(new_n2726_), .A2(new_n2732_), .B(new_n2470_), .ZN(new_n2994_));
  NAND2_X1   g02924(.A1(new_n2993_), .A2(new_n2994_), .ZN(new_n2995_));
  INV_X1     g02925(.I(new_n2751_), .ZN(new_n2996_));
  AOI22_X1   g02926(.A1(new_n2748_), .A2(new_n2241_), .B1(new_n2744_), .B2(new_n2745_), .ZN(new_n2997_));
  AOI21_X1   g02927(.A1(new_n2250_), .A2(new_n2253_), .B(new_n2242_), .ZN(new_n2998_));
  NOR3_X1    g02928(.A1(new_n2998_), .A2(new_n2997_), .A3(new_n2470_), .ZN(new_n2999_));
  AOI21_X1   g02929(.A1(new_n2995_), .A2(new_n2996_), .B(new_n2999_), .ZN(new_n3000_));
  NOR3_X1    g02930(.A1(new_n2528_), .A2(new_n2531_), .A3(new_n2496_), .ZN(new_n3001_));
  AOI21_X1   g02931(.A1(new_n2755_), .A2(new_n2754_), .B(new_n2470_), .ZN(new_n3002_));
  NOR3_X1    g02932(.A1(new_n3001_), .A2(new_n3002_), .A3(new_n2524_), .ZN(new_n3003_));
  NOR3_X1    g02933(.A1(new_n3003_), .A2(new_n3000_), .A3(new_n2968_), .ZN(new_n3004_));
  NAND2_X1   g02934(.A1(new_n2966_), .A2(new_n3004_), .ZN(new_n3005_));
  OAI21_X1   g02935(.A1(new_n2966_), .A2(new_n3004_), .B(new_n2762_), .ZN(new_n3006_));
  NAND2_X1   g02936(.A1(new_n3006_), .A2(new_n3005_), .ZN(new_n3007_));
  OAI21_X1   g02937(.A1(new_n2773_), .A2(new_n2774_), .B(new_n498_), .ZN(new_n3008_));
  NAND3_X1   g02938(.A1(new_n2771_), .A2(new_n2768_), .A3(\a[8] ), .ZN(new_n3009_));
  NAND2_X1   g02939(.A1(new_n3008_), .A2(new_n3009_), .ZN(new_n3010_));
  NAND2_X1   g02940(.A1(new_n2770_), .A2(new_n2765_), .ZN(new_n3011_));
  NAND2_X1   g02941(.A1(new_n2777_), .A2(new_n2778_), .ZN(new_n3012_));
  NAND2_X1   g02942(.A1(new_n3012_), .A2(new_n3011_), .ZN(new_n3013_));
  NAND3_X1   g02943(.A1(new_n2785_), .A2(new_n2786_), .A3(new_n2470_), .ZN(new_n3014_));
  AOI21_X1   g02944(.A1(new_n2791_), .A2(new_n3014_), .B(new_n3013_), .ZN(new_n3015_));
  OAI21_X1   g02945(.A1(new_n3015_), .A2(new_n3010_), .B(new_n3007_), .ZN(new_n3016_));
  NOR2_X1    g02946(.A1(new_n3016_), .A2(new_n2965_), .ZN(new_n3017_));
  INV_X1     g02947(.I(new_n2792_), .ZN(new_n3018_));
  AOI21_X1   g02948(.A1(new_n3016_), .A2(new_n2965_), .B(new_n3018_), .ZN(new_n3019_));
  NOR2_X1    g02949(.A1(new_n3019_), .A2(new_n3017_), .ZN(new_n3020_));
  NAND2_X1   g02950(.A1(new_n2428_), .A2(new_n2323_), .ZN(new_n3021_));
  NAND2_X1   g02951(.A1(new_n2300_), .A2(new_n2431_), .ZN(new_n3022_));
  NAND2_X1   g02952(.A1(new_n3022_), .A2(new_n3021_), .ZN(new_n3023_));
  INV_X1     g02953(.I(new_n2795_), .ZN(new_n3024_));
  NOR3_X1    g02954(.A1(new_n3024_), .A2(new_n3023_), .A3(new_n2796_), .ZN(new_n3025_));
  NOR3_X1    g02955(.A1(new_n3025_), .A2(new_n3020_), .A3(new_n2962_), .ZN(new_n3026_));
  NOR2_X1    g02956(.A1(new_n3026_), .A2(new_n2959_), .ZN(new_n3027_));
  NOR2_X1    g02957(.A1(new_n2957_), .A2(new_n2799_), .ZN(new_n3028_));
  NOR3_X1    g02958(.A1(new_n3027_), .A2(new_n3028_), .A3(new_n2797_), .ZN(new_n3029_));
  NOR2_X1    g02959(.A1(new_n3029_), .A2(new_n2961_), .ZN(new_n3030_));
  OAI21_X1   g02960(.A1(new_n2963_), .A2(new_n2964_), .B(new_n2496_), .ZN(new_n3031_));
  NOR2_X1    g02961(.A1(new_n2789_), .A2(new_n3031_), .ZN(new_n3032_));
  AOI21_X1   g02962(.A1(new_n2508_), .A2(new_n2511_), .B(new_n2470_), .ZN(new_n3033_));
  NOR2_X1    g02963(.A1(new_n3016_), .A2(new_n3033_), .ZN(new_n3034_));
  OAI21_X1   g02964(.A1(new_n3032_), .A2(new_n3034_), .B(new_n2791_), .ZN(new_n3035_));
  NAND2_X1   g02965(.A1(new_n3016_), .A2(new_n3033_), .ZN(new_n3036_));
  NAND2_X1   g02966(.A1(new_n2789_), .A2(new_n3031_), .ZN(new_n3037_));
  NAND3_X1   g02967(.A1(new_n3037_), .A2(new_n3036_), .A3(new_n2787_), .ZN(new_n3038_));
  NAND2_X1   g02968(.A1(new_n3035_), .A2(new_n3038_), .ZN(new_n3039_));
  INV_X1     g02969(.I(new_n2898_), .ZN(new_n3040_));
  NOR3_X1    g02970(.A1(new_n2894_), .A2(\a[2] ), .A3(\a[3] ), .ZN(new_n3041_));
  AOI21_X1   g02971(.A1(\a[3] ), .A2(new_n2896_), .B(new_n3041_), .ZN(new_n3042_));
  NOR2_X1    g02972(.A1(new_n3040_), .A2(new_n3042_), .ZN(new_n3043_));
  XOR2_X1    g02973(.A1(new_n3043_), .A2(new_n452_), .Z(new_n3044_));
  INV_X1     g02974(.I(new_n3044_), .ZN(new_n3045_));
  NAND3_X1   g02975(.A1(new_n2750_), .A2(new_n2747_), .A3(new_n2470_), .ZN(new_n3046_));
  OAI21_X1   g02976(.A1(new_n2998_), .A2(new_n2997_), .B(new_n2496_), .ZN(new_n3047_));
  NAND2_X1   g02977(.A1(new_n3047_), .A2(new_n3046_), .ZN(new_n3048_));
  NAND2_X1   g02978(.A1(new_n2995_), .A2(new_n3048_), .ZN(new_n3049_));
  NAND2_X1   g02979(.A1(new_n2996_), .A2(new_n2752_), .ZN(new_n3050_));
  NAND2_X1   g02980(.A1(new_n2743_), .A2(new_n3050_), .ZN(new_n3051_));
  NAND2_X1   g02981(.A1(new_n3049_), .A2(new_n3051_), .ZN(new_n3052_));
  NOR2_X1    g02982(.A1(new_n2982_), .A2(new_n2682_), .ZN(new_n3053_));
  XOR2_X1    g02983(.A1(new_n3053_), .A2(new_n2983_), .Z(new_n3054_));
  AOI22_X1   g02984(.A1(new_n2683_), .A2(new_n2680_), .B1(new_n2977_), .B2(new_n2978_), .ZN(new_n3055_));
  NAND2_X1   g02985(.A1(new_n2978_), .A2(new_n2977_), .ZN(new_n3056_));
  NAND3_X1   g02986(.A1(new_n2979_), .A2(new_n2980_), .A3(new_n2496_), .ZN(new_n3057_));
  OAI21_X1   g02987(.A1(new_n2677_), .A2(new_n2679_), .B(new_n2470_), .ZN(new_n3058_));
  AOI21_X1   g02988(.A1(new_n3057_), .A2(new_n3058_), .B(new_n3056_), .ZN(new_n3059_));
  NOR2_X1    g02989(.A1(new_n3059_), .A2(new_n3055_), .ZN(new_n3060_));
  INV_X1     g02990(.I(new_n3060_), .ZN(new_n3061_));
  AOI21_X1   g02991(.A1(new_n2657_), .A2(new_n2655_), .B(new_n2659_), .ZN(new_n3062_));
  AOI21_X1   g02992(.A1(\a[8] ), .A2(new_n2660_), .B(new_n3062_), .ZN(new_n3063_));
  OAI21_X1   g02993(.A1(new_n2556_), .A2(new_n2553_), .B(new_n2496_), .ZN(new_n3064_));
  AOI21_X1   g02994(.A1(new_n3063_), .A2(new_n2666_), .B(new_n3064_), .ZN(new_n3065_));
  OAI21_X1   g02995(.A1(new_n2554_), .A2(new_n2555_), .B(new_n2196_), .ZN(new_n3066_));
  NAND3_X1   g02996(.A1(new_n2552_), .A2(new_n2545_), .A3(new_n2199_), .ZN(new_n3067_));
  AOI21_X1   g02997(.A1(new_n3066_), .A2(new_n3067_), .B(new_n2470_), .ZN(new_n3068_));
  NOR3_X1    g02998(.A1(new_n2974_), .A2(new_n3068_), .A3(new_n2975_), .ZN(new_n3069_));
  OAI21_X1   g02999(.A1(new_n3065_), .A2(new_n3069_), .B(new_n2669_), .ZN(new_n3070_));
  OAI21_X1   g03000(.A1(new_n2974_), .A2(new_n2975_), .B(new_n3068_), .ZN(new_n3071_));
  NAND3_X1   g03001(.A1(new_n3063_), .A2(new_n3064_), .A3(new_n2666_), .ZN(new_n3072_));
  NAND3_X1   g03002(.A1(new_n3072_), .A2(new_n3071_), .A3(new_n2663_), .ZN(new_n3073_));
  NAND2_X1   g03003(.A1(new_n3070_), .A2(new_n3073_), .ZN(new_n3074_));
  NOR2_X1    g03004(.A1(new_n2651_), .A2(new_n2652_), .ZN(new_n3075_));
  NOR2_X1    g03005(.A1(new_n2653_), .A2(new_n2623_), .ZN(new_n3076_));
  NOR2_X1    g03006(.A1(new_n3076_), .A2(new_n3075_), .ZN(new_n3077_));
  NOR2_X1    g03007(.A1(new_n3077_), .A2(new_n2654_), .ZN(new_n3078_));
  INV_X1     g03008(.I(new_n3078_), .ZN(new_n3079_));
  NAND2_X1   g03009(.A1(new_n2649_), .A2(new_n2647_), .ZN(new_n3080_));
  NAND2_X1   g03010(.A1(new_n2608_), .A2(new_n2605_), .ZN(new_n3081_));
  NAND2_X1   g03011(.A1(new_n3081_), .A2(new_n3080_), .ZN(new_n3082_));
  XOR2_X1    g03012(.A1(new_n2604_), .A2(new_n2470_), .Z(new_n3083_));
  OAI21_X1   g03013(.A1(new_n3080_), .A2(new_n3083_), .B(new_n3082_), .ZN(new_n3084_));
  NAND2_X1   g03014(.A1(new_n2600_), .A2(new_n2496_), .ZN(new_n3085_));
  INV_X1     g03015(.I(new_n3085_), .ZN(new_n3086_));
  NAND3_X1   g03016(.A1(new_n2640_), .A2(new_n2598_), .A3(new_n2496_), .ZN(new_n3087_));
  OAI21_X1   g03017(.A1(new_n2582_), .A2(new_n2470_), .B(new_n2646_), .ZN(new_n3088_));
  AOI21_X1   g03018(.A1(new_n3088_), .A2(new_n3087_), .B(new_n3086_), .ZN(new_n3089_));
  NOR3_X1    g03019(.A1(new_n2582_), .A2(new_n2470_), .A3(new_n2646_), .ZN(new_n3090_));
  AOI21_X1   g03020(.A1(new_n2640_), .A2(new_n2496_), .B(new_n2598_), .ZN(new_n3091_));
  NOR3_X1    g03021(.A1(new_n3090_), .A2(new_n3091_), .A3(new_n3085_), .ZN(new_n3092_));
  NOR2_X1    g03022(.A1(new_n3092_), .A2(new_n3089_), .ZN(new_n3093_));
  NOR3_X1    g03023(.A1(new_n1079_), .A2(new_n2496_), .A3(new_n2574_), .ZN(new_n3094_));
  AOI21_X1   g03024(.A1(new_n1079_), .A2(new_n2574_), .B(new_n2470_), .ZN(new_n3095_));
  NOR2_X1    g03025(.A1(new_n3095_), .A2(new_n3094_), .ZN(new_n3096_));
  NAND2_X1   g03026(.A1(new_n2645_), .A2(new_n2596_), .ZN(new_n3097_));
  INV_X1     g03027(.I(new_n3097_), .ZN(new_n3098_));
  NAND2_X1   g03028(.A1(new_n2591_), .A2(new_n2899_), .ZN(new_n3099_));
  NAND2_X1   g03029(.A1(new_n2644_), .A2(new_n2905_), .ZN(new_n3100_));
  AOI22_X1   g03030(.A1(new_n3100_), .A2(new_n3099_), .B1(new_n2645_), .B2(new_n2596_), .ZN(new_n3101_));
  XOR2_X1    g03031(.A1(new_n2591_), .A2(new_n2899_), .Z(new_n3102_));
  AOI21_X1   g03032(.A1(new_n3098_), .A2(new_n3102_), .B(new_n3101_), .ZN(new_n3103_));
  OAI21_X1   g03033(.A1(new_n3103_), .A2(new_n3096_), .B(new_n2905_), .ZN(new_n3104_));
  INV_X1     g03034(.I(new_n2584_), .ZN(new_n3105_));
  NOR2_X1    g03035(.A1(new_n2470_), .A2(new_n3105_), .ZN(new_n3106_));
  NOR2_X1    g03036(.A1(new_n2496_), .A2(new_n2584_), .ZN(new_n3107_));
  NOR2_X1    g03037(.A1(new_n3106_), .A2(new_n3107_), .ZN(new_n3108_));
  NAND2_X1   g03038(.A1(new_n2496_), .A2(new_n2584_), .ZN(new_n3109_));
  OAI21_X1   g03039(.A1(new_n3108_), .A2(new_n2905_), .B(new_n3109_), .ZN(new_n3110_));
  INV_X1     g03040(.I(new_n3110_), .ZN(new_n3111_));
  NAND2_X1   g03041(.A1(new_n2496_), .A2(new_n3105_), .ZN(new_n3112_));
  NAND2_X1   g03042(.A1(new_n2496_), .A2(new_n2573_), .ZN(new_n3113_));
  XOR2_X1    g03043(.A1(new_n3112_), .A2(new_n3113_), .Z(new_n3114_));
  NAND2_X1   g03044(.A1(new_n3114_), .A2(new_n2905_), .ZN(new_n3115_));
  NOR2_X1    g03045(.A1(new_n3114_), .A2(new_n2905_), .ZN(new_n3116_));
  AOI21_X1   g03046(.A1(new_n3111_), .A2(new_n3115_), .B(new_n3116_), .ZN(new_n3117_));
  NOR2_X1    g03047(.A1(new_n2585_), .A2(new_n2586_), .ZN(new_n3118_));
  NOR2_X1    g03048(.A1(new_n2587_), .A2(new_n3112_), .ZN(new_n3119_));
  OAI21_X1   g03049(.A1(new_n3118_), .A2(new_n3119_), .B(new_n2470_), .ZN(new_n3120_));
  NOR2_X1    g03050(.A1(new_n806_), .A2(new_n2641_), .ZN(new_n3121_));
  NOR2_X1    g03051(.A1(new_n1079_), .A2(new_n2574_), .ZN(new_n3122_));
  OAI21_X1   g03052(.A1(new_n3121_), .A2(new_n3122_), .B(new_n2470_), .ZN(new_n3123_));
  NOR2_X1    g03053(.A1(new_n3112_), .A2(new_n2586_), .ZN(new_n3124_));
  NOR2_X1    g03054(.A1(new_n3123_), .A2(new_n3124_), .ZN(new_n3125_));
  XOR2_X1    g03055(.A1(new_n1079_), .A2(new_n2641_), .Z(new_n3126_));
  NAND2_X1   g03056(.A1(new_n2585_), .A2(new_n2587_), .ZN(new_n3127_));
  AOI21_X1   g03057(.A1(new_n3126_), .A2(new_n2470_), .B(new_n3127_), .ZN(new_n3128_));
  OAI21_X1   g03058(.A1(new_n3128_), .A2(new_n3125_), .B(new_n3120_), .ZN(new_n3129_));
  NAND2_X1   g03059(.A1(new_n2587_), .A2(new_n3112_), .ZN(new_n3130_));
  NAND2_X1   g03060(.A1(new_n2585_), .A2(new_n2586_), .ZN(new_n3131_));
  AOI21_X1   g03061(.A1(new_n3131_), .A2(new_n3130_), .B(new_n2496_), .ZN(new_n3132_));
  NAND2_X1   g03062(.A1(new_n3126_), .A2(new_n2470_), .ZN(new_n3133_));
  NAND2_X1   g03063(.A1(new_n3123_), .A2(new_n3124_), .ZN(new_n3134_));
  NAND3_X1   g03064(.A1(new_n3132_), .A2(new_n3133_), .A3(new_n3134_), .ZN(new_n3135_));
  AOI21_X1   g03065(.A1(new_n3129_), .A2(new_n3135_), .B(new_n2905_), .ZN(new_n3136_));
  NAND3_X1   g03066(.A1(new_n3129_), .A2(new_n3135_), .A3(new_n2905_), .ZN(new_n3137_));
  OAI21_X1   g03067(.A1(new_n3117_), .A2(new_n3136_), .B(new_n3137_), .ZN(new_n3138_));
  NAND2_X1   g03068(.A1(new_n3103_), .A2(new_n3096_), .ZN(new_n3139_));
  NAND3_X1   g03069(.A1(new_n3104_), .A2(new_n3138_), .A3(new_n3139_), .ZN(new_n3140_));
  NOR2_X1    g03070(.A1(new_n3140_), .A2(new_n3093_), .ZN(new_n3141_));
  XOR2_X1    g03071(.A1(new_n3097_), .A2(new_n2644_), .Z(new_n3142_));
  NOR2_X1    g03072(.A1(new_n3142_), .A2(new_n2899_), .ZN(new_n3143_));
  NAND2_X1   g03073(.A1(new_n3143_), .A2(new_n2899_), .ZN(new_n3144_));
  AOI21_X1   g03074(.A1(new_n3140_), .A2(new_n3093_), .B(new_n3144_), .ZN(new_n3145_));
  OAI21_X1   g03075(.A1(new_n3145_), .A2(new_n3141_), .B(new_n3084_), .ZN(new_n3146_));
  NOR3_X1    g03076(.A1(new_n3145_), .A2(new_n3141_), .A3(new_n3084_), .ZN(new_n3147_));
  OAI21_X1   g03077(.A1(new_n452_), .A2(new_n3147_), .B(new_n3146_), .ZN(new_n3148_));
  NAND3_X1   g03078(.A1(new_n3148_), .A2(new_n2905_), .A3(new_n3079_), .ZN(new_n3149_));
  NOR2_X1    g03079(.A1(new_n2572_), .A2(new_n2496_), .ZN(new_n3150_));
  XOR2_X1    g03080(.A1(new_n3150_), .A2(new_n2621_), .Z(new_n3151_));
  NOR2_X1    g03081(.A1(new_n3151_), .A2(new_n2623_), .ZN(new_n3152_));
  XOR2_X1    g03082(.A1(new_n3150_), .A2(new_n2654_), .Z(new_n3153_));
  NOR2_X1    g03083(.A1(new_n3153_), .A2(new_n2620_), .ZN(new_n3154_));
  NOR2_X1    g03084(.A1(new_n3154_), .A2(new_n3152_), .ZN(new_n3155_));
  INV_X1     g03085(.I(new_n3147_), .ZN(new_n3156_));
  NAND2_X1   g03086(.A1(new_n3156_), .A2(\a[5] ), .ZN(new_n3157_));
  NAND4_X1   g03087(.A1(new_n3157_), .A2(new_n2899_), .A3(new_n3078_), .A4(new_n3146_), .ZN(new_n3158_));
  NAND2_X1   g03088(.A1(new_n3158_), .A2(new_n3155_), .ZN(new_n3159_));
  NOR3_X1    g03089(.A1(new_n2665_), .A2(new_n2663_), .A3(new_n2899_), .ZN(new_n3160_));
  OAI21_X1   g03090(.A1(new_n2550_), .A2(new_n2662_), .B(new_n2470_), .ZN(new_n3161_));
  AOI21_X1   g03091(.A1(new_n2669_), .A2(new_n3161_), .B(new_n2905_), .ZN(new_n3162_));
  NOR2_X1    g03092(.A1(new_n3160_), .A2(new_n3162_), .ZN(new_n3163_));
  NOR2_X1    g03093(.A1(new_n3063_), .A2(new_n3163_), .ZN(new_n3164_));
  OAI21_X1   g03094(.A1(new_n2665_), .A2(new_n2663_), .B(new_n2905_), .ZN(new_n3165_));
  NAND3_X1   g03095(.A1(new_n2669_), .A2(new_n3161_), .A3(new_n2899_), .ZN(new_n3166_));
  AOI21_X1   g03096(.A1(new_n3165_), .A2(new_n3166_), .B(new_n2974_), .ZN(new_n3167_));
  OAI21_X1   g03097(.A1(new_n3167_), .A2(new_n3164_), .B(new_n2899_), .ZN(new_n3168_));
  NAND3_X1   g03098(.A1(new_n3168_), .A2(new_n3159_), .A3(new_n3149_), .ZN(new_n3169_));
  NOR2_X1    g03099(.A1(new_n3167_), .A2(new_n3164_), .ZN(new_n3170_));
  OAI21_X1   g03100(.A1(new_n2625_), .A2(new_n2622_), .B(new_n2659_), .ZN(new_n3171_));
  NOR2_X1    g03101(.A1(new_n2625_), .A2(new_n2622_), .ZN(new_n3172_));
  NAND2_X1   g03102(.A1(new_n3172_), .A2(new_n2635_), .ZN(new_n3173_));
  AOI21_X1   g03103(.A1(new_n3173_), .A2(new_n3171_), .B(\a[8] ), .ZN(new_n3174_));
  NOR2_X1    g03104(.A1(new_n3172_), .A2(new_n2635_), .ZN(new_n3175_));
  NOR3_X1    g03105(.A1(new_n2625_), .A2(new_n2659_), .A3(new_n2622_), .ZN(new_n3176_));
  NOR3_X1    g03106(.A1(new_n3175_), .A2(new_n498_), .A3(new_n3176_), .ZN(new_n3177_));
  NOR2_X1    g03107(.A1(new_n3177_), .A2(new_n3174_), .ZN(new_n3178_));
  AOI21_X1   g03108(.A1(new_n3170_), .A2(new_n2905_), .B(new_n3178_), .ZN(new_n3179_));
  NAND3_X1   g03109(.A1(new_n3169_), .A2(new_n3074_), .A3(new_n3179_), .ZN(new_n3180_));
  XOR2_X1    g03110(.A1(new_n3151_), .A2(new_n2620_), .Z(new_n3181_));
  NOR3_X1    g03111(.A1(new_n3148_), .A2(new_n2905_), .A3(new_n3079_), .ZN(new_n3182_));
  OAI21_X1   g03112(.A1(new_n3181_), .A2(new_n3182_), .B(new_n3149_), .ZN(new_n3183_));
  NOR2_X1    g03113(.A1(new_n2973_), .A2(new_n498_), .ZN(new_n3184_));
  OAI22_X1   g03114(.A1(new_n3184_), .A2(new_n3062_), .B1(new_n3160_), .B2(new_n3162_), .ZN(new_n3185_));
  NAND2_X1   g03115(.A1(new_n3165_), .A2(new_n3166_), .ZN(new_n3186_));
  NAND2_X1   g03116(.A1(new_n3063_), .A2(new_n3186_), .ZN(new_n3187_));
  AOI21_X1   g03117(.A1(new_n3187_), .A2(new_n3185_), .B(new_n2905_), .ZN(new_n3188_));
  NOR2_X1    g03118(.A1(new_n3183_), .A2(new_n3188_), .ZN(new_n3189_));
  OR2_X2     g03119(.A1(new_n3177_), .A2(new_n3174_), .Z(new_n3190_));
  NAND3_X1   g03120(.A1(new_n3187_), .A2(new_n3185_), .A3(new_n2905_), .ZN(new_n3191_));
  NAND2_X1   g03121(.A1(new_n3191_), .A2(new_n3190_), .ZN(new_n3192_));
  NOR2_X1    g03122(.A1(new_n3189_), .A2(new_n3192_), .ZN(new_n3193_));
  NOR2_X1    g03123(.A1(new_n3063_), .A2(new_n2975_), .ZN(new_n3194_));
  NOR2_X1    g03124(.A1(new_n2974_), .A2(new_n2666_), .ZN(new_n3195_));
  OAI21_X1   g03125(.A1(new_n3194_), .A2(new_n3195_), .B(new_n2905_), .ZN(new_n3196_));
  NOR2_X1    g03126(.A1(new_n3196_), .A2(new_n2905_), .ZN(new_n3197_));
  OAI21_X1   g03127(.A1(new_n3193_), .A2(new_n3074_), .B(new_n3197_), .ZN(new_n3198_));
  NAND2_X1   g03128(.A1(new_n3198_), .A2(new_n3180_), .ZN(new_n3199_));
  OAI21_X1   g03129(.A1(new_n3199_), .A2(new_n3045_), .B(new_n3061_), .ZN(new_n3200_));
  AOI21_X1   g03130(.A1(new_n3072_), .A2(new_n3071_), .B(new_n2663_), .ZN(new_n3201_));
  NOR3_X1    g03131(.A1(new_n3065_), .A2(new_n3069_), .A3(new_n2669_), .ZN(new_n3202_));
  NOR2_X1    g03132(.A1(new_n3202_), .A2(new_n3201_), .ZN(new_n3203_));
  NOR3_X1    g03133(.A1(new_n3203_), .A2(new_n3189_), .A3(new_n3192_), .ZN(new_n3204_));
  AOI21_X1   g03134(.A1(new_n3169_), .A2(new_n3179_), .B(new_n3074_), .ZN(new_n3205_));
  INV_X1     g03135(.I(new_n3197_), .ZN(new_n3206_));
  NOR2_X1    g03136(.A1(new_n3205_), .A2(new_n3206_), .ZN(new_n3207_));
  OAI21_X1   g03137(.A1(new_n3207_), .A2(new_n3204_), .B(new_n3045_), .ZN(new_n3208_));
  NAND2_X1   g03138(.A1(new_n3200_), .A2(new_n3208_), .ZN(new_n3209_));
  NAND3_X1   g03139(.A1(new_n3209_), .A2(new_n2905_), .A3(new_n3054_), .ZN(new_n3210_));
  NOR3_X1    g03140(.A1(new_n2984_), .A2(new_n2496_), .A3(new_n2541_), .ZN(new_n3211_));
  AOI21_X1   g03141(.A1(new_n2470_), .A2(new_n2971_), .B(new_n2702_), .ZN(new_n3212_));
  OAI21_X1   g03142(.A1(new_n3212_), .A2(new_n3211_), .B(new_n2701_), .ZN(new_n3213_));
  INV_X1     g03143(.I(new_n2701_), .ZN(new_n3214_));
  NAND3_X1   g03144(.A1(new_n2702_), .A2(new_n2971_), .A3(new_n2470_), .ZN(new_n3215_));
  OAI21_X1   g03145(.A1(new_n2496_), .A2(new_n2541_), .B(new_n2984_), .ZN(new_n3216_));
  NAND3_X1   g03146(.A1(new_n3216_), .A2(new_n3215_), .A3(new_n3214_), .ZN(new_n3217_));
  NAND2_X1   g03147(.A1(new_n3213_), .A2(new_n3217_), .ZN(new_n3218_));
  INV_X1     g03148(.I(new_n3218_), .ZN(new_n3219_));
  INV_X1     g03149(.I(new_n3054_), .ZN(new_n3220_));
  NAND4_X1   g03150(.A1(new_n3200_), .A2(new_n3220_), .A3(new_n2899_), .A4(new_n3208_), .ZN(new_n3221_));
  NAND2_X1   g03151(.A1(new_n3221_), .A2(new_n3219_), .ZN(new_n3222_));
  OAI21_X1   g03152(.A1(new_n2726_), .A2(new_n2732_), .B(new_n2496_), .ZN(new_n3223_));
  NAND3_X1   g03153(.A1(new_n2736_), .A2(new_n2741_), .A3(new_n2470_), .ZN(new_n3224_));
  NAND2_X1   g03154(.A1(new_n3223_), .A2(new_n3224_), .ZN(new_n3225_));
  OAI21_X1   g03155(.A1(new_n2991_), .A2(new_n2723_), .B(new_n3225_), .ZN(new_n3226_));
  NAND2_X1   g03156(.A1(new_n2994_), .A2(new_n2992_), .ZN(new_n3227_));
  NAND3_X1   g03157(.A1(new_n3227_), .A2(new_n2722_), .A3(new_n2724_), .ZN(new_n3228_));
  NAND3_X1   g03158(.A1(new_n3226_), .A2(new_n3228_), .A3(new_n2899_), .ZN(new_n3229_));
  NAND3_X1   g03159(.A1(new_n3222_), .A2(new_n3210_), .A3(new_n3229_), .ZN(new_n3230_));
  NAND2_X1   g03160(.A1(new_n2986_), .A2(new_n2985_), .ZN(new_n3231_));
  AOI21_X1   g03161(.A1(new_n2716_), .A2(new_n2710_), .B(new_n2989_), .ZN(new_n3232_));
  NOR3_X1    g03162(.A1(new_n2987_), .A2(new_n2988_), .A3(new_n2720_), .ZN(new_n3233_));
  NOR2_X1    g03163(.A1(new_n3233_), .A2(new_n3232_), .ZN(new_n3234_));
  NOR2_X1    g03164(.A1(new_n2990_), .A2(new_n2723_), .ZN(new_n3235_));
  MUX2_X1    g03165(.I0(new_n3235_), .I1(new_n3234_), .S(new_n3231_), .Z(new_n3236_));
  AOI22_X1   g03166(.A1(new_n2722_), .A2(new_n2724_), .B1(new_n3223_), .B2(new_n3224_), .ZN(new_n3237_));
  NOR2_X1    g03167(.A1(new_n2733_), .A2(new_n2742_), .ZN(new_n3238_));
  NOR3_X1    g03168(.A1(new_n3238_), .A2(new_n2991_), .A3(new_n2723_), .ZN(new_n3239_));
  NOR3_X1    g03169(.A1(new_n3239_), .A2(new_n3237_), .A3(new_n2899_), .ZN(new_n3240_));
  NOR2_X1    g03170(.A1(new_n3240_), .A2(new_n3236_), .ZN(new_n3241_));
  NAND3_X1   g03171(.A1(new_n3230_), .A2(new_n3052_), .A3(new_n3241_), .ZN(new_n3242_));
  AOI22_X1   g03172(.A1(new_n2993_), .A2(new_n2994_), .B1(new_n3046_), .B2(new_n3047_), .ZN(new_n3243_));
  NOR2_X1    g03173(.A1(new_n2999_), .A2(new_n2751_), .ZN(new_n3244_));
  NOR3_X1    g03174(.A1(new_n3244_), .A2(new_n2734_), .A3(new_n2742_), .ZN(new_n3245_));
  NOR2_X1    g03175(.A1(new_n3243_), .A2(new_n3245_), .ZN(new_n3246_));
  OAI21_X1   g03176(.A1(new_n3189_), .A2(new_n3192_), .B(new_n3203_), .ZN(new_n3247_));
  AOI21_X1   g03177(.A1(new_n3247_), .A2(new_n3197_), .B(new_n3204_), .ZN(new_n3248_));
  AOI21_X1   g03178(.A1(new_n3248_), .A2(new_n3044_), .B(new_n3060_), .ZN(new_n3249_));
  AOI21_X1   g03179(.A1(new_n3198_), .A2(new_n3180_), .B(new_n3044_), .ZN(new_n3250_));
  NOR2_X1    g03180(.A1(new_n3249_), .A2(new_n3250_), .ZN(new_n3251_));
  NOR3_X1    g03181(.A1(new_n3251_), .A2(new_n2899_), .A3(new_n3220_), .ZN(new_n3252_));
  NOR4_X1    g03182(.A1(new_n3249_), .A2(new_n2905_), .A3(new_n3054_), .A4(new_n3250_), .ZN(new_n3253_));
  NOR2_X1    g03183(.A1(new_n3253_), .A2(new_n3218_), .ZN(new_n3254_));
  NOR3_X1    g03184(.A1(new_n3239_), .A2(new_n3237_), .A3(new_n2905_), .ZN(new_n3255_));
  NOR3_X1    g03185(.A1(new_n3254_), .A2(new_n3252_), .A3(new_n3255_), .ZN(new_n3256_));
  NAND2_X1   g03186(.A1(new_n3226_), .A2(new_n3228_), .ZN(new_n3257_));
  OAI21_X1   g03187(.A1(new_n3233_), .A2(new_n3232_), .B(new_n3231_), .ZN(new_n3258_));
  OAI21_X1   g03188(.A1(new_n3231_), .A2(new_n3235_), .B(new_n3258_), .ZN(new_n3259_));
  OAI21_X1   g03189(.A1(new_n2899_), .A2(new_n3257_), .B(new_n3259_), .ZN(new_n3260_));
  OAI21_X1   g03190(.A1(new_n3256_), .A2(new_n3260_), .B(new_n3246_), .ZN(new_n3261_));
  AOI21_X1   g03191(.A1(new_n3226_), .A2(new_n3228_), .B(new_n2899_), .ZN(new_n3262_));
  NAND2_X1   g03192(.A1(new_n3262_), .A2(new_n2899_), .ZN(new_n3263_));
  INV_X1     g03193(.I(new_n3263_), .ZN(new_n3264_));
  NAND2_X1   g03194(.A1(new_n3261_), .A2(new_n3264_), .ZN(new_n3265_));
  NAND2_X1   g03195(.A1(new_n2524_), .A2(new_n2496_), .ZN(new_n3266_));
  NAND2_X1   g03196(.A1(new_n2525_), .A2(new_n2470_), .ZN(new_n3267_));
  AOI21_X1   g03197(.A1(new_n3266_), .A2(new_n3267_), .B(new_n3000_), .ZN(new_n3268_));
  NAND2_X1   g03198(.A1(new_n2525_), .A2(new_n2496_), .ZN(new_n3269_));
  NAND2_X1   g03199(.A1(new_n2524_), .A2(new_n2470_), .ZN(new_n3270_));
  AOI21_X1   g03200(.A1(new_n3269_), .A2(new_n3270_), .B(new_n2753_), .ZN(new_n3271_));
  NOR2_X1    g03201(.A1(new_n3268_), .A2(new_n3271_), .ZN(new_n3272_));
  AOI21_X1   g03202(.A1(new_n3265_), .A2(new_n3242_), .B(new_n3272_), .ZN(new_n3273_));
  NAND3_X1   g03203(.A1(new_n3265_), .A2(new_n3242_), .A3(new_n3272_), .ZN(new_n3274_));
  AOI21_X1   g03204(.A1(new_n3045_), .A2(new_n3274_), .B(new_n3273_), .ZN(new_n3275_));
  MUX2_X1    g03205(.I0(new_n2470_), .I1(new_n2524_), .S(new_n2967_), .Z(new_n3276_));
  XOR2_X1    g03206(.A1(new_n3276_), .A2(new_n2753_), .Z(new_n3277_));
  NOR2_X1    g03207(.A1(new_n3277_), .A2(new_n2899_), .ZN(new_n3278_));
  NAND2_X1   g03208(.A1(new_n3277_), .A2(new_n2899_), .ZN(new_n3279_));
  OAI21_X1   g03209(.A1(new_n3275_), .A2(new_n3278_), .B(new_n3279_), .ZN(new_n3280_));
  NOR2_X1    g03210(.A1(new_n2519_), .A2(new_n2496_), .ZN(new_n3281_));
  NAND2_X1   g03211(.A1(new_n3281_), .A2(new_n2759_), .ZN(new_n3282_));
  NOR2_X1    g03212(.A1(new_n3281_), .A2(new_n2759_), .ZN(new_n3283_));
  INV_X1     g03213(.I(new_n3283_), .ZN(new_n3284_));
  AOI21_X1   g03214(.A1(new_n3284_), .A2(new_n3282_), .B(new_n3002_), .ZN(new_n3285_));
  INV_X1     g03215(.I(new_n3282_), .ZN(new_n3286_));
  NOR3_X1    g03216(.A1(new_n3286_), .A2(new_n2757_), .A3(new_n3283_), .ZN(new_n3287_));
  OAI21_X1   g03217(.A1(new_n3285_), .A2(new_n3287_), .B(new_n2899_), .ZN(new_n3288_));
  NOR3_X1    g03218(.A1(new_n3285_), .A2(new_n3287_), .A3(new_n2899_), .ZN(new_n3289_));
  AOI21_X1   g03219(.A1(new_n3280_), .A2(new_n3288_), .B(new_n3289_), .ZN(new_n3290_));
  XOR2_X1    g03220(.A1(new_n3007_), .A2(new_n3010_), .Z(new_n3291_));
  NOR3_X1    g03221(.A1(new_n2787_), .A2(new_n2784_), .A3(new_n2779_), .ZN(new_n3292_));
  NOR3_X1    g03222(.A1(new_n3292_), .A2(new_n3007_), .A3(new_n2776_), .ZN(new_n3293_));
  NAND3_X1   g03223(.A1(new_n2791_), .A2(new_n3014_), .A3(new_n3013_), .ZN(new_n3294_));
  AOI21_X1   g03224(.A1(new_n3294_), .A2(new_n3010_), .B(new_n2763_), .ZN(new_n3295_));
  NOR3_X1    g03225(.A1(new_n3293_), .A2(new_n3295_), .A3(new_n2905_), .ZN(new_n3296_));
  NAND3_X1   g03226(.A1(new_n3294_), .A2(new_n2763_), .A3(new_n3010_), .ZN(new_n3297_));
  OAI21_X1   g03227(.A1(new_n3292_), .A2(new_n2776_), .B(new_n3007_), .ZN(new_n3298_));
  AOI21_X1   g03228(.A1(new_n3298_), .A2(new_n3297_), .B(new_n2899_), .ZN(new_n3299_));
  NOR3_X1    g03229(.A1(new_n3296_), .A2(new_n3299_), .A3(new_n3291_), .ZN(new_n3300_));
  NAND2_X1   g03230(.A1(new_n3298_), .A2(new_n3297_), .ZN(new_n3301_));
  AOI21_X1   g03231(.A1(new_n3301_), .A2(new_n3291_), .B(new_n2899_), .ZN(new_n3302_));
  NOR3_X1    g03232(.A1(new_n3300_), .A2(new_n3290_), .A3(new_n3302_), .ZN(new_n3303_));
  NAND2_X1   g03233(.A1(new_n3303_), .A2(new_n3039_), .ZN(new_n3304_));
  NOR2_X1    g03234(.A1(new_n3293_), .A2(new_n3295_), .ZN(new_n3305_));
  NOR2_X1    g03235(.A1(new_n3305_), .A2(new_n2905_), .ZN(new_n3306_));
  OAI21_X1   g03236(.A1(new_n3303_), .A2(new_n3039_), .B(new_n3306_), .ZN(new_n3307_));
  NAND2_X1   g03237(.A1(new_n3307_), .A2(new_n3304_), .ZN(new_n3308_));
  NAND2_X1   g03238(.A1(new_n2497_), .A2(new_n2470_), .ZN(new_n3309_));
  NAND2_X1   g03239(.A1(new_n3023_), .A2(new_n2496_), .ZN(new_n3310_));
  NAND2_X1   g03240(.A1(new_n3309_), .A2(new_n3310_), .ZN(new_n3311_));
  NAND3_X1   g03241(.A1(new_n2793_), .A2(new_n2790_), .A3(new_n3043_), .ZN(new_n3312_));
  INV_X1     g03242(.I(new_n3043_), .ZN(new_n3313_));
  OAI21_X1   g03243(.A1(new_n3019_), .A2(new_n3017_), .B(new_n3313_), .ZN(new_n3314_));
  AOI21_X1   g03244(.A1(new_n3312_), .A2(new_n3314_), .B(new_n3311_), .ZN(new_n3315_));
  XOR2_X1    g03245(.A1(new_n3023_), .A2(new_n2496_), .Z(new_n3316_));
  NOR3_X1    g03246(.A1(new_n3019_), .A2(new_n3017_), .A3(new_n3313_), .ZN(new_n3317_));
  AOI21_X1   g03247(.A1(new_n2793_), .A2(new_n2790_), .B(new_n3043_), .ZN(new_n3318_));
  NOR3_X1    g03248(.A1(new_n3318_), .A2(new_n3317_), .A3(new_n3316_), .ZN(new_n3319_));
  OAI21_X1   g03249(.A1(new_n3315_), .A2(new_n3319_), .B(new_n452_), .ZN(new_n3320_));
  OAI21_X1   g03250(.A1(new_n3318_), .A2(new_n3317_), .B(new_n3316_), .ZN(new_n3321_));
  NAND3_X1   g03251(.A1(new_n3312_), .A2(new_n3314_), .A3(new_n3311_), .ZN(new_n3322_));
  NAND3_X1   g03252(.A1(new_n3321_), .A2(new_n3322_), .A3(\a[5] ), .ZN(new_n3323_));
  NAND2_X1   g03253(.A1(new_n3320_), .A2(new_n3323_), .ZN(new_n3324_));
  NOR2_X1    g03254(.A1(new_n3316_), .A2(\a[5] ), .ZN(new_n3325_));
  NOR2_X1    g03255(.A1(new_n3311_), .A2(new_n452_), .ZN(new_n3326_));
  OAI22_X1   g03256(.A1(new_n3325_), .A2(new_n3326_), .B1(new_n3317_), .B2(new_n3318_), .ZN(new_n3327_));
  MUX2_X1    g03257(.I0(new_n3023_), .I1(new_n2470_), .S(new_n2502_), .Z(new_n3328_));
  NAND2_X1   g03258(.A1(new_n3328_), .A2(new_n3020_), .ZN(new_n3329_));
  MUX2_X1    g03259(.I0(new_n2497_), .I1(new_n2496_), .S(new_n2502_), .Z(new_n3330_));
  NAND2_X1   g03260(.A1(new_n3330_), .A2(new_n2794_), .ZN(new_n3331_));
  NAND3_X1   g03261(.A1(new_n3329_), .A2(new_n3331_), .A3(new_n2905_), .ZN(new_n3332_));
  NOR2_X1    g03262(.A1(new_n3330_), .A2(new_n2794_), .ZN(new_n3333_));
  NOR2_X1    g03263(.A1(new_n3328_), .A2(new_n3020_), .ZN(new_n3334_));
  OAI21_X1   g03264(.A1(new_n3333_), .A2(new_n3334_), .B(new_n2899_), .ZN(new_n3335_));
  AOI21_X1   g03265(.A1(new_n3335_), .A2(new_n3332_), .B(new_n3327_), .ZN(new_n3336_));
  OAI21_X1   g03266(.A1(new_n3336_), .A2(new_n3324_), .B(new_n3308_), .ZN(new_n3337_));
  NOR2_X1    g03267(.A1(new_n3337_), .A2(new_n3030_), .ZN(new_n3338_));
  NOR2_X1    g03268(.A1(new_n3332_), .A2(new_n2899_), .ZN(new_n3339_));
  INV_X1     g03269(.I(new_n3339_), .ZN(new_n3340_));
  AOI21_X1   g03270(.A1(new_n3337_), .A2(new_n3030_), .B(new_n3340_), .ZN(new_n3341_));
  OAI21_X1   g03271(.A1(new_n3341_), .A2(new_n3338_), .B(new_n2899_), .ZN(new_n3342_));
  OAI21_X1   g03272(.A1(new_n3027_), .A2(new_n3028_), .B(new_n2797_), .ZN(new_n3343_));
  NAND3_X1   g03273(.A1(new_n2958_), .A2(new_n2960_), .A3(new_n2796_), .ZN(new_n3344_));
  NAND2_X1   g03274(.A1(new_n3343_), .A2(new_n3344_), .ZN(new_n3345_));
  AOI21_X1   g03275(.A1(new_n3037_), .A2(new_n3036_), .B(new_n2787_), .ZN(new_n3346_));
  NOR3_X1    g03276(.A1(new_n3032_), .A2(new_n3034_), .A3(new_n2791_), .ZN(new_n3347_));
  NOR2_X1    g03277(.A1(new_n3346_), .A2(new_n3347_), .ZN(new_n3348_));
  AOI21_X1   g03278(.A1(new_n3230_), .A2(new_n3241_), .B(new_n3052_), .ZN(new_n3349_));
  OAI21_X1   g03279(.A1(new_n3349_), .A2(new_n3263_), .B(new_n3242_), .ZN(new_n3350_));
  INV_X1     g03280(.I(new_n3272_), .ZN(new_n3351_));
  NAND2_X1   g03281(.A1(new_n3350_), .A2(new_n3351_), .ZN(new_n3352_));
  OAI21_X1   g03282(.A1(new_n3350_), .A2(new_n3351_), .B(new_n3045_), .ZN(new_n3353_));
  NAND2_X1   g03283(.A1(new_n3353_), .A2(new_n3352_), .ZN(new_n3354_));
  INV_X1     g03284(.I(new_n3278_), .ZN(new_n3355_));
  INV_X1     g03285(.I(new_n3279_), .ZN(new_n3356_));
  AOI21_X1   g03286(.A1(new_n3354_), .A2(new_n3355_), .B(new_n3356_), .ZN(new_n3357_));
  OAI21_X1   g03287(.A1(new_n3286_), .A2(new_n3283_), .B(new_n2757_), .ZN(new_n3358_));
  INV_X1     g03288(.I(new_n3287_), .ZN(new_n3359_));
  AOI21_X1   g03289(.A1(new_n3359_), .A2(new_n3358_), .B(new_n2905_), .ZN(new_n3360_));
  NAND3_X1   g03290(.A1(new_n3359_), .A2(new_n3358_), .A3(new_n2905_), .ZN(new_n3361_));
  OAI21_X1   g03291(.A1(new_n3357_), .A2(new_n3360_), .B(new_n3361_), .ZN(new_n3362_));
  XOR2_X1    g03292(.A1(new_n3007_), .A2(new_n2776_), .Z(new_n3363_));
  NAND3_X1   g03293(.A1(new_n3298_), .A2(new_n3297_), .A3(new_n2899_), .ZN(new_n3364_));
  OAI21_X1   g03294(.A1(new_n3293_), .A2(new_n3295_), .B(new_n2905_), .ZN(new_n3365_));
  NAND3_X1   g03295(.A1(new_n3365_), .A2(new_n3364_), .A3(new_n3363_), .ZN(new_n3366_));
  OAI21_X1   g03296(.A1(new_n3305_), .A2(new_n3363_), .B(new_n2905_), .ZN(new_n3367_));
  NAND3_X1   g03297(.A1(new_n3362_), .A2(new_n3366_), .A3(new_n3367_), .ZN(new_n3368_));
  NOR2_X1    g03298(.A1(new_n3368_), .A2(new_n3348_), .ZN(new_n3369_));
  INV_X1     g03299(.I(new_n3306_), .ZN(new_n3370_));
  AOI21_X1   g03300(.A1(new_n3368_), .A2(new_n3348_), .B(new_n3370_), .ZN(new_n3371_));
  NOR2_X1    g03301(.A1(new_n3371_), .A2(new_n3369_), .ZN(new_n3372_));
  AOI21_X1   g03302(.A1(new_n3321_), .A2(new_n3322_), .B(\a[5] ), .ZN(new_n3373_));
  NOR3_X1    g03303(.A1(new_n3315_), .A2(new_n3319_), .A3(new_n452_), .ZN(new_n3374_));
  NOR2_X1    g03304(.A1(new_n3374_), .A2(new_n3373_), .ZN(new_n3375_));
  NAND2_X1   g03305(.A1(new_n3311_), .A2(new_n452_), .ZN(new_n3376_));
  NAND2_X1   g03306(.A1(new_n3316_), .A2(\a[5] ), .ZN(new_n3377_));
  AOI22_X1   g03307(.A1(new_n3377_), .A2(new_n3376_), .B1(new_n3312_), .B2(new_n3314_), .ZN(new_n3378_));
  NOR3_X1    g03308(.A1(new_n3333_), .A2(new_n3334_), .A3(new_n2899_), .ZN(new_n3379_));
  AOI21_X1   g03309(.A1(new_n3329_), .A2(new_n3331_), .B(new_n2905_), .ZN(new_n3380_));
  OAI21_X1   g03310(.A1(new_n3380_), .A2(new_n3379_), .B(new_n3378_), .ZN(new_n3381_));
  AOI21_X1   g03311(.A1(new_n3375_), .A2(new_n3381_), .B(new_n3372_), .ZN(new_n3382_));
  NAND2_X1   g03312(.A1(new_n3382_), .A2(new_n3345_), .ZN(new_n3383_));
  OAI21_X1   g03313(.A1(new_n3382_), .A2(new_n3345_), .B(new_n3339_), .ZN(new_n3384_));
  NAND3_X1   g03314(.A1(new_n3384_), .A2(new_n3383_), .A3(new_n2905_), .ZN(new_n3385_));
  NAND3_X1   g03315(.A1(new_n2440_), .A2(new_n2448_), .A3(new_n2439_), .ZN(new_n3386_));
  OAI21_X1   g03316(.A1(new_n2337_), .A2(new_n2340_), .B(new_n2354_), .ZN(new_n3387_));
  AOI21_X1   g03317(.A1(new_n3387_), .A2(new_n3386_), .B(new_n2470_), .ZN(new_n3388_));
  NOR3_X1    g03318(.A1(new_n2471_), .A2(new_n2472_), .A3(new_n2496_), .ZN(new_n3389_));
  NOR2_X1    g03319(.A1(new_n3388_), .A2(new_n3389_), .ZN(new_n3390_));
  XNOR2_X1   g03320(.A1(new_n2804_), .A2(new_n3390_), .ZN(new_n3391_));
  INV_X1     g03321(.I(new_n3391_), .ZN(new_n3392_));
  NAND2_X1   g03322(.A1(new_n3385_), .A2(new_n3392_), .ZN(new_n3393_));
  AOI21_X1   g03323(.A1(new_n3393_), .A2(new_n3342_), .B(new_n2954_), .ZN(new_n3394_));
  AOI21_X1   g03324(.A1(new_n3384_), .A2(new_n3383_), .B(new_n2905_), .ZN(new_n3395_));
  NOR2_X1    g03325(.A1(new_n3341_), .A2(new_n3338_), .ZN(new_n3396_));
  AOI21_X1   g03326(.A1(new_n3396_), .A2(new_n2905_), .B(new_n3391_), .ZN(new_n3397_));
  NOR3_X1    g03327(.A1(new_n3397_), .A2(new_n2953_), .A3(new_n3395_), .ZN(new_n3398_));
  OAI21_X1   g03328(.A1(new_n3394_), .A2(new_n3398_), .B(new_n452_), .ZN(new_n3399_));
  OAI21_X1   g03329(.A1(new_n3397_), .A2(new_n3395_), .B(new_n2953_), .ZN(new_n3400_));
  NAND3_X1   g03330(.A1(new_n3393_), .A2(new_n2954_), .A3(new_n3342_), .ZN(new_n3401_));
  NAND3_X1   g03331(.A1(new_n3400_), .A2(new_n3401_), .A3(\a[5] ), .ZN(new_n3402_));
  NAND2_X1   g03332(.A1(new_n3399_), .A2(new_n3402_), .ZN(new_n3403_));
  NOR3_X1    g03333(.A1(new_n3380_), .A2(new_n3379_), .A3(new_n3378_), .ZN(new_n3404_));
  OR3_X2     g03334(.A1(new_n3375_), .A2(new_n3404_), .A3(new_n3308_), .Z(new_n3405_));
  OAI21_X1   g03335(.A1(new_n3375_), .A2(new_n3404_), .B(new_n3308_), .ZN(new_n3406_));
  NAND2_X1   g03336(.A1(new_n3405_), .A2(new_n3406_), .ZN(new_n3407_));
  INV_X1     g03337(.I(new_n3407_), .ZN(new_n3408_));
  INV_X1     g03338(.I(\a[0] ), .ZN(new_n3409_));
  XNOR2_X1   g03339(.A1(\a[1] ), .A2(\a[2] ), .ZN(new_n3410_));
  NOR2_X1    g03340(.A1(new_n3410_), .A2(new_n3409_), .ZN(new_n3411_));
  NAND2_X1   g03341(.A1(new_n3411_), .A2(\a[2] ), .ZN(new_n3412_));
  INV_X1     g03342(.I(new_n3412_), .ZN(new_n3413_));
  INV_X1     g03343(.I(new_n3411_), .ZN(new_n3414_));
  NOR2_X1    g03344(.A1(\a[0] ), .A2(\a[1] ), .ZN(new_n3415_));
  INV_X1     g03345(.I(new_n3415_), .ZN(new_n3416_));
  OAI21_X1   g03346(.A1(new_n3414_), .A2(new_n3416_), .B(\a[2] ), .ZN(new_n3417_));
  NAND2_X1   g03347(.A1(new_n3108_), .A2(new_n2899_), .ZN(new_n3418_));
  XNOR2_X1   g03348(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n3419_));
  AND3_X2    g03349(.A1(new_n3411_), .A2(\a[2] ), .A3(new_n3419_), .Z(new_n3420_));
  NOR2_X1    g03350(.A1(new_n3420_), .A2(new_n2899_), .ZN(new_n3421_));
  AOI21_X1   g03351(.A1(new_n3420_), .A2(new_n2899_), .B(new_n451_), .ZN(new_n3422_));
  NOR3_X1    g03352(.A1(new_n3040_), .A2(new_n452_), .A3(new_n2492_), .ZN(new_n3423_));
  OAI22_X1   g03353(.A1(new_n3422_), .A2(new_n3421_), .B1(new_n3423_), .B2(new_n3412_), .ZN(new_n3424_));
  NAND2_X1   g03354(.A1(new_n3423_), .A2(new_n3412_), .ZN(new_n3425_));
  OAI21_X1   g03355(.A1(new_n3106_), .A2(new_n3107_), .B(new_n2905_), .ZN(new_n3426_));
  AOI22_X1   g03356(.A1(new_n3424_), .A2(new_n3425_), .B1(new_n3418_), .B2(new_n3426_), .ZN(new_n3427_));
  NAND4_X1   g03357(.A1(new_n3424_), .A2(new_n3418_), .A3(new_n3425_), .A4(new_n3426_), .ZN(new_n3428_));
  AOI21_X1   g03358(.A1(\a[2] ), .A2(new_n3428_), .B(new_n3427_), .ZN(new_n3429_));
  XOR2_X1    g03359(.A1(new_n3109_), .A2(new_n2899_), .Z(new_n3430_));
  XOR2_X1    g03360(.A1(new_n3430_), .A2(new_n3418_), .Z(new_n3431_));
  AOI21_X1   g03361(.A1(new_n3429_), .A2(new_n3431_), .B(new_n3413_), .ZN(new_n3432_));
  OAI21_X1   g03362(.A1(new_n3429_), .A2(new_n3431_), .B(new_n3413_), .ZN(new_n3433_));
  XOR2_X1    g03363(.A1(new_n3114_), .A2(new_n2905_), .Z(new_n3434_));
  XOR2_X1    g03364(.A1(new_n3434_), .A2(new_n3111_), .Z(new_n3435_));
  AOI21_X1   g03365(.A1(new_n3435_), .A2(new_n3433_), .B(new_n3432_), .ZN(new_n3436_));
  INV_X1     g03366(.I(new_n3117_), .ZN(new_n3437_));
  AOI21_X1   g03367(.A1(new_n3133_), .A2(new_n3134_), .B(new_n3132_), .ZN(new_n3438_));
  INV_X1     g03368(.I(new_n3135_), .ZN(new_n3439_));
  NOR3_X1    g03369(.A1(new_n3439_), .A2(new_n3438_), .A3(new_n2905_), .ZN(new_n3440_));
  AOI21_X1   g03370(.A1(new_n3129_), .A2(new_n3135_), .B(new_n2899_), .ZN(new_n3441_));
  OAI21_X1   g03371(.A1(new_n3440_), .A2(new_n3441_), .B(new_n3437_), .ZN(new_n3442_));
  NOR3_X1    g03372(.A1(new_n3439_), .A2(new_n3438_), .A3(new_n2899_), .ZN(new_n3443_));
  OAI21_X1   g03373(.A1(new_n3443_), .A2(new_n3136_), .B(new_n3117_), .ZN(new_n3444_));
  AOI21_X1   g03374(.A1(new_n3442_), .A2(new_n3444_), .B(new_n3412_), .ZN(new_n3445_));
  NAND3_X1   g03375(.A1(new_n3442_), .A2(new_n3444_), .A3(new_n3412_), .ZN(new_n3446_));
  OAI21_X1   g03376(.A1(new_n3436_), .A2(new_n3445_), .B(new_n3446_), .ZN(new_n3447_));
  NOR3_X1    g03377(.A1(new_n3095_), .A2(new_n3094_), .A3(new_n2899_), .ZN(new_n3448_));
  NOR2_X1    g03378(.A1(new_n3096_), .A2(new_n2905_), .ZN(new_n3449_));
  OAI21_X1   g03379(.A1(new_n3448_), .A2(new_n3449_), .B(new_n3138_), .ZN(new_n3450_));
  XOR2_X1    g03380(.A1(new_n3096_), .A2(new_n2899_), .Z(new_n3451_));
  OAI21_X1   g03381(.A1(new_n3138_), .A2(new_n3451_), .B(new_n3450_), .ZN(new_n3452_));
  NAND2_X1   g03382(.A1(new_n3447_), .A2(new_n3452_), .ZN(new_n3453_));
  XOR2_X1    g03383(.A1(\a[1] ), .A2(\a[2] ), .Z(new_n3454_));
  NOR2_X1    g03384(.A1(new_n3454_), .A2(new_n3409_), .ZN(new_n3455_));
  INV_X1     g03385(.I(new_n3455_), .ZN(new_n3456_));
  NOR2_X1    g03386(.A1(new_n3414_), .A2(new_n3456_), .ZN(new_n3457_));
  NOR2_X1    g03387(.A1(new_n3457_), .A2(new_n451_), .ZN(new_n3458_));
  NOR3_X1    g03388(.A1(new_n3414_), .A2(new_n3456_), .A3(\a[2] ), .ZN(new_n3459_));
  OAI22_X1   g03389(.A1(new_n3447_), .A2(new_n3452_), .B1(new_n3458_), .B2(new_n3459_), .ZN(new_n3460_));
  NOR3_X1    g03390(.A1(new_n3103_), .A2(new_n3449_), .A3(new_n3451_), .ZN(new_n3461_));
  INV_X1     g03391(.I(new_n3461_), .ZN(new_n3462_));
  NOR2_X1    g03392(.A1(new_n3096_), .A2(new_n2905_), .ZN(new_n3463_));
  INV_X1     g03393(.I(new_n3463_), .ZN(new_n3464_));
  AOI21_X1   g03394(.A1(new_n3462_), .A2(new_n3464_), .B(new_n3138_), .ZN(new_n3465_));
  INV_X1     g03395(.I(new_n3465_), .ZN(new_n3466_));
  NAND3_X1   g03396(.A1(new_n3462_), .A2(new_n3138_), .A3(new_n3464_), .ZN(new_n3467_));
  AOI21_X1   g03397(.A1(new_n3466_), .A2(new_n3467_), .B(new_n3412_), .ZN(new_n3468_));
  AOI21_X1   g03398(.A1(new_n3460_), .A2(new_n3453_), .B(new_n3468_), .ZN(new_n3469_));
  AND3_X2    g03399(.A1(new_n3466_), .A2(new_n3412_), .A3(new_n3467_), .Z(new_n3470_));
  INV_X1     g03400(.I(new_n3140_), .ZN(new_n3471_));
  OAI21_X1   g03401(.A1(new_n3092_), .A2(new_n3089_), .B(new_n2899_), .ZN(new_n3472_));
  NOR2_X1    g03402(.A1(new_n3471_), .A2(new_n3472_), .ZN(new_n3473_));
  INV_X1     g03403(.I(new_n3472_), .ZN(new_n3474_));
  NOR2_X1    g03404(.A1(new_n3474_), .A2(new_n3140_), .ZN(new_n3475_));
  OAI22_X1   g03405(.A1(new_n3473_), .A2(new_n3475_), .B1(new_n2899_), .B2(new_n3142_), .ZN(new_n3476_));
  NAND2_X1   g03406(.A1(new_n3474_), .A2(new_n3140_), .ZN(new_n3477_));
  NAND2_X1   g03407(.A1(new_n3471_), .A2(new_n3472_), .ZN(new_n3478_));
  NAND3_X1   g03408(.A1(new_n3478_), .A2(new_n3477_), .A3(new_n3143_), .ZN(new_n3479_));
  NAND2_X1   g03409(.A1(new_n3476_), .A2(new_n3479_), .ZN(new_n3480_));
  OAI21_X1   g03410(.A1(new_n3469_), .A2(new_n3470_), .B(new_n3480_), .ZN(new_n3481_));
  NOR3_X1    g03411(.A1(new_n3469_), .A2(new_n3480_), .A3(new_n3470_), .ZN(new_n3482_));
  OAI21_X1   g03412(.A1(new_n451_), .A2(new_n3482_), .B(new_n3481_), .ZN(new_n3483_));
  NOR2_X1    g03413(.A1(new_n3145_), .A2(new_n3141_), .ZN(new_n3484_));
  NAND2_X1   g03414(.A1(new_n3484_), .A2(new_n3084_), .ZN(new_n3485_));
  NOR2_X1    g03415(.A1(new_n3484_), .A2(new_n3084_), .ZN(new_n3486_));
  INV_X1     g03416(.I(new_n3486_), .ZN(new_n3487_));
  AOI21_X1   g03417(.A1(new_n3487_), .A2(new_n3485_), .B(\a[5] ), .ZN(new_n3488_));
  INV_X1     g03418(.I(new_n3485_), .ZN(new_n3489_));
  NOR3_X1    g03419(.A1(new_n3489_), .A2(new_n452_), .A3(new_n3486_), .ZN(new_n3490_));
  OAI21_X1   g03420(.A1(new_n3488_), .A2(new_n3490_), .B(new_n3413_), .ZN(new_n3491_));
  NOR3_X1    g03421(.A1(new_n3488_), .A2(new_n3490_), .A3(new_n3413_), .ZN(new_n3492_));
  AOI21_X1   g03422(.A1(new_n3483_), .A2(new_n3491_), .B(new_n3492_), .ZN(new_n3493_));
  XOR2_X1    g03423(.A1(new_n3078_), .A2(new_n2899_), .Z(new_n3494_));
  XNOR2_X1   g03424(.A1(new_n3494_), .A2(new_n3148_), .ZN(new_n3495_));
  AOI21_X1   g03425(.A1(new_n3493_), .A2(new_n3495_), .B(new_n3413_), .ZN(new_n3496_));
  OAI21_X1   g03426(.A1(new_n3493_), .A2(new_n3495_), .B(new_n3413_), .ZN(new_n3497_));
  OAI21_X1   g03427(.A1(new_n3148_), .A2(new_n2899_), .B(new_n3079_), .ZN(new_n3498_));
  NAND2_X1   g03428(.A1(new_n3148_), .A2(new_n2899_), .ZN(new_n3499_));
  NAND2_X1   g03429(.A1(new_n3498_), .A2(new_n3499_), .ZN(new_n3500_));
  NAND2_X1   g03430(.A1(new_n3155_), .A2(new_n2905_), .ZN(new_n3501_));
  OAI21_X1   g03431(.A1(new_n3154_), .A2(new_n3152_), .B(new_n2899_), .ZN(new_n3502_));
  NAND2_X1   g03432(.A1(new_n3501_), .A2(new_n3502_), .ZN(new_n3503_));
  XOR2_X1    g03433(.A1(new_n3503_), .A2(new_n3500_), .Z(new_n3504_));
  AOI21_X1   g03434(.A1(new_n3504_), .A2(new_n3497_), .B(new_n3496_), .ZN(new_n3505_));
  NOR2_X1    g03435(.A1(new_n3183_), .A2(new_n2899_), .ZN(new_n3506_));
  NAND2_X1   g03436(.A1(new_n3183_), .A2(new_n2899_), .ZN(new_n3507_));
  INV_X1     g03437(.I(new_n3507_), .ZN(new_n3508_));
  OAI21_X1   g03438(.A1(new_n3508_), .A2(new_n3506_), .B(new_n3190_), .ZN(new_n3509_));
  AOI21_X1   g03439(.A1(new_n3159_), .A2(new_n3149_), .B(new_n2899_), .ZN(new_n3510_));
  NOR2_X1    g03440(.A1(new_n3183_), .A2(new_n2905_), .ZN(new_n3511_));
  OAI21_X1   g03441(.A1(new_n3510_), .A2(new_n3511_), .B(new_n3178_), .ZN(new_n3512_));
  AOI21_X1   g03442(.A1(new_n3509_), .A2(new_n3512_), .B(new_n3412_), .ZN(new_n3513_));
  NAND3_X1   g03443(.A1(new_n3509_), .A2(new_n3512_), .A3(new_n3412_), .ZN(new_n3514_));
  OAI21_X1   g03444(.A1(new_n3505_), .A2(new_n3513_), .B(new_n3514_), .ZN(new_n3515_));
  INV_X1     g03445(.I(new_n3170_), .ZN(new_n3516_));
  OAI21_X1   g03446(.A1(new_n3510_), .A2(new_n3511_), .B(new_n3516_), .ZN(new_n3517_));
  NOR2_X1    g03447(.A1(new_n3517_), .A2(new_n3508_), .ZN(new_n3518_));
  NAND2_X1   g03448(.A1(new_n3183_), .A2(new_n2899_), .ZN(new_n3519_));
  INV_X1     g03449(.I(new_n3519_), .ZN(new_n3520_));
  OAI21_X1   g03450(.A1(new_n3518_), .A2(new_n3520_), .B(new_n3178_), .ZN(new_n3521_));
  NAND2_X1   g03451(.A1(new_n3183_), .A2(new_n2905_), .ZN(new_n3522_));
  NAND3_X1   g03452(.A1(new_n3159_), .A2(new_n2899_), .A3(new_n3149_), .ZN(new_n3523_));
  NAND2_X1   g03453(.A1(new_n3523_), .A2(new_n3522_), .ZN(new_n3524_));
  NAND3_X1   g03454(.A1(new_n3524_), .A2(new_n3516_), .A3(new_n3507_), .ZN(new_n3525_));
  NAND3_X1   g03455(.A1(new_n3525_), .A2(new_n3190_), .A3(new_n3519_), .ZN(new_n3526_));
  NAND2_X1   g03456(.A1(new_n3521_), .A2(new_n3526_), .ZN(new_n3527_));
  NAND2_X1   g03457(.A1(new_n3515_), .A2(new_n3527_), .ZN(new_n3528_));
  INV_X1     g03458(.I(new_n3417_), .ZN(new_n3529_));
  OAI21_X1   g03459(.A1(new_n3515_), .A2(new_n3527_), .B(new_n3529_), .ZN(new_n3530_));
  NAND2_X1   g03460(.A1(new_n3169_), .A2(new_n3179_), .ZN(new_n3531_));
  NAND3_X1   g03461(.A1(new_n3531_), .A2(new_n2899_), .A3(new_n3074_), .ZN(new_n3532_));
  NAND2_X1   g03462(.A1(new_n3074_), .A2(new_n2899_), .ZN(new_n3533_));
  NAND2_X1   g03463(.A1(new_n3533_), .A2(new_n3193_), .ZN(new_n3534_));
  NAND2_X1   g03464(.A1(new_n3532_), .A2(new_n3534_), .ZN(new_n3535_));
  NAND2_X1   g03465(.A1(new_n3535_), .A2(new_n3196_), .ZN(new_n3536_));
  INV_X1     g03466(.I(new_n3196_), .ZN(new_n3537_));
  NAND3_X1   g03467(.A1(new_n3532_), .A2(new_n3534_), .A3(new_n3537_), .ZN(new_n3538_));
  AOI21_X1   g03468(.A1(new_n3536_), .A2(new_n3538_), .B(new_n3413_), .ZN(new_n3539_));
  AOI21_X1   g03469(.A1(new_n3530_), .A2(new_n3528_), .B(new_n3539_), .ZN(new_n3540_));
  NAND3_X1   g03470(.A1(new_n3536_), .A2(new_n3413_), .A3(new_n3538_), .ZN(new_n3541_));
  INV_X1     g03471(.I(new_n3541_), .ZN(new_n3542_));
  XOR2_X1    g03472(.A1(new_n3248_), .A2(new_n3045_), .Z(new_n3543_));
  NOR2_X1    g03473(.A1(new_n3199_), .A2(new_n3045_), .ZN(new_n3544_));
  OAI21_X1   g03474(.A1(new_n3544_), .A2(new_n3250_), .B(new_n3060_), .ZN(new_n3545_));
  OAI21_X1   g03475(.A1(new_n3543_), .A2(new_n3060_), .B(new_n3545_), .ZN(new_n3546_));
  OAI21_X1   g03476(.A1(new_n3540_), .A2(new_n3542_), .B(new_n3546_), .ZN(new_n3547_));
  NOR3_X1    g03477(.A1(new_n3540_), .A2(new_n3546_), .A3(new_n3542_), .ZN(new_n3548_));
  OAI21_X1   g03478(.A1(new_n3417_), .A2(new_n3548_), .B(new_n3547_), .ZN(new_n3549_));
  XOR2_X1    g03479(.A1(new_n3054_), .A2(new_n2899_), .Z(new_n3550_));
  XOR2_X1    g03480(.A1(new_n3550_), .A2(new_n3209_), .Z(new_n3551_));
  INV_X1     g03481(.I(new_n3551_), .ZN(new_n3552_));
  OAI21_X1   g03482(.A1(new_n3549_), .A2(new_n3552_), .B(new_n3412_), .ZN(new_n3553_));
  INV_X1     g03483(.I(new_n3553_), .ZN(new_n3554_));
  AOI21_X1   g03484(.A1(new_n3549_), .A2(new_n3552_), .B(new_n3412_), .ZN(new_n3555_));
  OAI21_X1   g03485(.A1(new_n3209_), .A2(new_n2899_), .B(new_n3054_), .ZN(new_n3556_));
  OAI21_X1   g03486(.A1(new_n2905_), .A2(new_n3251_), .B(new_n3556_), .ZN(new_n3557_));
  XOR2_X1    g03487(.A1(new_n3218_), .A2(new_n2899_), .Z(new_n3558_));
  XOR2_X1    g03488(.A1(new_n3557_), .A2(new_n3558_), .Z(new_n3559_));
  NOR2_X1    g03489(.A1(new_n3555_), .A2(new_n3559_), .ZN(new_n3560_));
  NOR2_X1    g03490(.A1(new_n3254_), .A2(new_n3252_), .ZN(new_n3561_));
  NAND2_X1   g03491(.A1(new_n3561_), .A2(new_n2905_), .ZN(new_n3562_));
  NAND2_X1   g03492(.A1(new_n3222_), .A2(new_n3210_), .ZN(new_n3563_));
  NAND2_X1   g03493(.A1(new_n3563_), .A2(new_n2899_), .ZN(new_n3564_));
  AOI21_X1   g03494(.A1(new_n3564_), .A2(new_n3562_), .B(new_n3236_), .ZN(new_n3565_));
  NAND2_X1   g03495(.A1(new_n3563_), .A2(new_n2905_), .ZN(new_n3566_));
  NAND2_X1   g03496(.A1(new_n3561_), .A2(new_n2899_), .ZN(new_n3567_));
  AOI21_X1   g03497(.A1(new_n3566_), .A2(new_n3567_), .B(new_n3259_), .ZN(new_n3568_));
  OAI21_X1   g03498(.A1(new_n3565_), .A2(new_n3568_), .B(new_n3413_), .ZN(new_n3569_));
  OAI21_X1   g03499(.A1(new_n3560_), .A2(new_n3554_), .B(new_n3569_), .ZN(new_n3570_));
  NOR3_X1    g03500(.A1(new_n3565_), .A2(new_n3568_), .A3(new_n3413_), .ZN(new_n3571_));
  INV_X1     g03501(.I(new_n3571_), .ZN(new_n3572_));
  MUX2_X1    g03502(.I0(new_n2899_), .I1(new_n3563_), .S(new_n3257_), .Z(new_n3573_));
  NAND2_X1   g03503(.A1(new_n3573_), .A2(new_n3236_), .ZN(new_n3574_));
  NOR2_X1    g03504(.A1(new_n3573_), .A2(new_n3236_), .ZN(new_n3575_));
  INV_X1     g03505(.I(new_n3575_), .ZN(new_n3576_));
  AOI21_X1   g03506(.A1(new_n3576_), .A2(new_n3574_), .B(new_n3412_), .ZN(new_n3577_));
  AOI21_X1   g03507(.A1(new_n3570_), .A2(new_n3572_), .B(new_n3577_), .ZN(new_n3578_));
  NAND3_X1   g03508(.A1(new_n3576_), .A2(new_n3412_), .A3(new_n3574_), .ZN(new_n3579_));
  INV_X1     g03509(.I(new_n3579_), .ZN(new_n3580_));
  NOR2_X1    g03510(.A1(new_n3578_), .A2(new_n3580_), .ZN(new_n3581_));
  NOR2_X1    g03511(.A1(new_n3256_), .A2(new_n3260_), .ZN(new_n3582_));
  NOR2_X1    g03512(.A1(new_n3246_), .A2(new_n2905_), .ZN(new_n3583_));
  XNOR2_X1   g03513(.A1(new_n3582_), .A2(new_n3583_), .ZN(new_n3584_));
  XOR2_X1    g03514(.A1(new_n3584_), .A2(new_n3262_), .Z(new_n3585_));
  INV_X1     g03515(.I(new_n3585_), .ZN(new_n3586_));
  NOR3_X1    g03516(.A1(new_n3581_), .A2(new_n3413_), .A3(new_n3586_), .ZN(new_n3587_));
  NOR4_X1    g03517(.A1(new_n3578_), .A2(new_n3412_), .A3(new_n3580_), .A4(new_n3585_), .ZN(new_n3588_));
  NOR2_X1    g03518(.A1(new_n3272_), .A2(new_n3044_), .ZN(new_n3589_));
  XOR2_X1    g03519(.A1(new_n3043_), .A2(new_n452_), .Z(new_n3590_));
  AOI21_X1   g03520(.A1(new_n3272_), .A2(new_n3590_), .B(new_n3589_), .ZN(new_n3591_));
  XOR2_X1    g03521(.A1(new_n3591_), .A2(new_n3350_), .Z(new_n3592_));
  NOR2_X1    g03522(.A1(new_n3588_), .A2(new_n3592_), .ZN(new_n3593_));
  NOR2_X1    g03523(.A1(new_n3593_), .A2(new_n3587_), .ZN(new_n3594_));
  NOR2_X1    g03524(.A1(new_n3356_), .A2(new_n3278_), .ZN(new_n3595_));
  XOR2_X1    g03525(.A1(new_n3595_), .A2(new_n3275_), .Z(new_n3596_));
  INV_X1     g03526(.I(new_n3596_), .ZN(new_n3597_));
  NOR3_X1    g03527(.A1(new_n3594_), .A2(new_n3413_), .A3(new_n3597_), .ZN(new_n3598_));
  NOR4_X1    g03528(.A1(new_n3593_), .A2(new_n3587_), .A3(new_n3412_), .A4(new_n3596_), .ZN(new_n3599_));
  NAND2_X1   g03529(.A1(new_n3361_), .A2(new_n3288_), .ZN(new_n3600_));
  XOR2_X1    g03530(.A1(new_n3600_), .A2(new_n3357_), .Z(new_n3601_));
  NOR2_X1    g03531(.A1(new_n3599_), .A2(new_n3601_), .ZN(new_n3602_));
  XOR2_X1    g03532(.A1(new_n3291_), .A2(new_n2905_), .Z(new_n3603_));
  NAND2_X1   g03533(.A1(new_n3603_), .A2(new_n3362_), .ZN(new_n3604_));
  XOR2_X1    g03534(.A1(new_n3291_), .A2(new_n2899_), .Z(new_n3605_));
  NAND2_X1   g03535(.A1(new_n3605_), .A2(new_n3290_), .ZN(new_n3606_));
  NAND2_X1   g03536(.A1(new_n3604_), .A2(new_n3606_), .ZN(new_n3607_));
  NAND2_X1   g03537(.A1(new_n3607_), .A2(new_n3413_), .ZN(new_n3608_));
  OAI21_X1   g03538(.A1(new_n3602_), .A2(new_n3598_), .B(new_n3608_), .ZN(new_n3609_));
  NOR2_X1    g03539(.A1(new_n3607_), .A2(new_n3413_), .ZN(new_n3610_));
  INV_X1     g03540(.I(new_n3610_), .ZN(new_n3611_));
  NAND2_X1   g03541(.A1(new_n3609_), .A2(new_n3611_), .ZN(new_n3612_));
  MUX2_X1    g03542(.I0(new_n2899_), .I1(new_n3291_), .S(new_n3301_), .Z(new_n3613_));
  XOR2_X1    g03543(.A1(new_n3613_), .A2(new_n3290_), .Z(new_n3614_));
  NOR2_X1    g03544(.A1(new_n3614_), .A2(new_n3412_), .ZN(new_n3615_));
  INV_X1     g03545(.I(new_n3615_), .ZN(new_n3616_));
  NAND2_X1   g03546(.A1(new_n3614_), .A2(new_n3412_), .ZN(new_n3617_));
  INV_X1     g03547(.I(new_n3617_), .ZN(new_n3618_));
  AOI21_X1   g03548(.A1(new_n3612_), .A2(new_n3616_), .B(new_n3618_), .ZN(new_n3619_));
  NAND2_X1   g03549(.A1(new_n3301_), .A2(new_n2899_), .ZN(new_n3620_));
  NOR3_X1    g03550(.A1(new_n3303_), .A2(new_n2905_), .A3(new_n3348_), .ZN(new_n3621_));
  AOI21_X1   g03551(.A1(new_n2899_), .A2(new_n3039_), .B(new_n3368_), .ZN(new_n3622_));
  OAI21_X1   g03552(.A1(new_n3622_), .A2(new_n3621_), .B(new_n3620_), .ZN(new_n3623_));
  INV_X1     g03553(.I(new_n3620_), .ZN(new_n3624_));
  NAND3_X1   g03554(.A1(new_n3368_), .A2(new_n2899_), .A3(new_n3039_), .ZN(new_n3625_));
  OAI21_X1   g03555(.A1(new_n2905_), .A2(new_n3348_), .B(new_n3303_), .ZN(new_n3626_));
  NAND3_X1   g03556(.A1(new_n3626_), .A2(new_n3625_), .A3(new_n3624_), .ZN(new_n3627_));
  NAND2_X1   g03557(.A1(new_n3623_), .A2(new_n3627_), .ZN(new_n3628_));
  NAND3_X1   g03558(.A1(new_n3320_), .A2(new_n3323_), .A3(new_n3413_), .ZN(new_n3629_));
  OAI21_X1   g03559(.A1(new_n3374_), .A2(new_n3373_), .B(new_n3412_), .ZN(new_n3630_));
  AOI21_X1   g03560(.A1(new_n3630_), .A2(new_n3629_), .B(new_n3372_), .ZN(new_n3631_));
  OAI21_X1   g03561(.A1(new_n3374_), .A2(new_n3373_), .B(new_n3413_), .ZN(new_n3632_));
  NAND3_X1   g03562(.A1(new_n3320_), .A2(new_n3323_), .A3(new_n3412_), .ZN(new_n3633_));
  AOI21_X1   g03563(.A1(new_n3632_), .A2(new_n3633_), .B(new_n3308_), .ZN(new_n3634_));
  NOR3_X1    g03564(.A1(new_n3631_), .A2(new_n3634_), .A3(new_n3628_), .ZN(new_n3635_));
  AOI21_X1   g03565(.A1(new_n3626_), .A2(new_n3625_), .B(new_n3624_), .ZN(new_n3636_));
  NOR3_X1    g03566(.A1(new_n3622_), .A2(new_n3621_), .A3(new_n3620_), .ZN(new_n3637_));
  NOR2_X1    g03567(.A1(new_n3637_), .A2(new_n3636_), .ZN(new_n3638_));
  NOR3_X1    g03568(.A1(new_n3374_), .A2(new_n3373_), .A3(new_n3412_), .ZN(new_n3639_));
  AOI21_X1   g03569(.A1(new_n3320_), .A2(new_n3323_), .B(new_n3413_), .ZN(new_n3640_));
  OAI21_X1   g03570(.A1(new_n3639_), .A2(new_n3640_), .B(new_n3308_), .ZN(new_n3641_));
  AOI21_X1   g03571(.A1(new_n3320_), .A2(new_n3323_), .B(new_n3412_), .ZN(new_n3642_));
  NOR3_X1    g03572(.A1(new_n3374_), .A2(new_n3373_), .A3(new_n3413_), .ZN(new_n3643_));
  OAI21_X1   g03573(.A1(new_n3643_), .A2(new_n3642_), .B(new_n3372_), .ZN(new_n3644_));
  AOI21_X1   g03574(.A1(new_n3641_), .A2(new_n3644_), .B(new_n3638_), .ZN(new_n3645_));
  NOR2_X1    g03575(.A1(new_n3645_), .A2(new_n3413_), .ZN(new_n3646_));
  NOR4_X1    g03576(.A1(new_n3619_), .A2(new_n3646_), .A3(new_n3408_), .A4(new_n3635_), .ZN(new_n3647_));
  NAND3_X1   g03577(.A1(new_n3641_), .A2(new_n3644_), .A3(new_n3638_), .ZN(new_n3648_));
  OAI21_X1   g03578(.A1(new_n3413_), .A2(new_n3645_), .B(new_n3648_), .ZN(new_n3649_));
  OAI21_X1   g03579(.A1(new_n3649_), .A2(new_n3619_), .B(new_n3408_), .ZN(new_n3650_));
  XOR2_X1    g03580(.A1(new_n3324_), .A2(new_n3308_), .Z(new_n3651_));
  NAND2_X1   g03581(.A1(new_n3651_), .A2(new_n3413_), .ZN(new_n3652_));
  XOR2_X1    g03582(.A1(new_n3457_), .A2(\a[2] ), .Z(new_n3653_));
  NOR2_X1    g03583(.A1(new_n3652_), .A2(new_n3653_), .ZN(new_n3654_));
  AOI21_X1   g03584(.A1(new_n3650_), .A2(new_n3654_), .B(new_n3647_), .ZN(new_n3655_));
  AOI21_X1   g03585(.A1(new_n3343_), .A2(new_n3344_), .B(new_n2899_), .ZN(new_n3656_));
  NAND2_X1   g03586(.A1(new_n3337_), .A2(new_n3656_), .ZN(new_n3657_));
  OAI21_X1   g03587(.A1(new_n3029_), .A2(new_n2961_), .B(new_n2905_), .ZN(new_n3658_));
  NAND2_X1   g03588(.A1(new_n3382_), .A2(new_n3658_), .ZN(new_n3659_));
  AOI21_X1   g03589(.A1(new_n3659_), .A2(new_n3657_), .B(new_n3379_), .ZN(new_n3660_));
  NOR2_X1    g03590(.A1(new_n3382_), .A2(new_n3658_), .ZN(new_n3661_));
  NOR2_X1    g03591(.A1(new_n3337_), .A2(new_n3656_), .ZN(new_n3662_));
  NOR3_X1    g03592(.A1(new_n3661_), .A2(new_n3662_), .A3(new_n3332_), .ZN(new_n3663_));
  NOR2_X1    g03593(.A1(new_n3660_), .A2(new_n3663_), .ZN(new_n3664_));
  NOR3_X1    g03594(.A1(new_n3388_), .A2(new_n3389_), .A3(new_n2899_), .ZN(new_n3665_));
  OAI21_X1   g03595(.A1(new_n2471_), .A2(new_n2472_), .B(new_n2496_), .ZN(new_n3666_));
  NAND3_X1   g03596(.A1(new_n3387_), .A2(new_n3386_), .A3(new_n2470_), .ZN(new_n3667_));
  AOI21_X1   g03597(.A1(new_n3667_), .A2(new_n3666_), .B(new_n2905_), .ZN(new_n3668_));
  OAI22_X1   g03598(.A1(new_n2803_), .A2(new_n2800_), .B1(new_n3665_), .B2(new_n3668_), .ZN(new_n3669_));
  OAI21_X1   g03599(.A1(new_n3388_), .A2(new_n3389_), .B(new_n2905_), .ZN(new_n3670_));
  NAND3_X1   g03600(.A1(new_n3667_), .A2(new_n3666_), .A3(new_n2899_), .ZN(new_n3671_));
  NAND2_X1   g03601(.A1(new_n3670_), .A2(new_n3671_), .ZN(new_n3672_));
  NAND2_X1   g03602(.A1(new_n2804_), .A2(new_n3672_), .ZN(new_n3673_));
  NAND2_X1   g03603(.A1(new_n3673_), .A2(new_n3669_), .ZN(new_n3674_));
  NAND2_X1   g03604(.A1(new_n3674_), .A2(\a[2] ), .ZN(new_n3675_));
  NAND3_X1   g03605(.A1(new_n3673_), .A2(new_n451_), .A3(new_n3669_), .ZN(new_n3676_));
  AOI22_X1   g03606(.A1(new_n3384_), .A2(new_n3383_), .B1(new_n3675_), .B2(new_n3676_), .ZN(new_n3677_));
  NAND2_X1   g03607(.A1(new_n2956_), .A2(new_n2955_), .ZN(new_n3678_));
  NAND2_X1   g03608(.A1(new_n3026_), .A2(new_n3678_), .ZN(new_n3679_));
  OAI21_X1   g03609(.A1(new_n3026_), .A2(new_n3678_), .B(new_n2801_), .ZN(new_n3680_));
  NAND3_X1   g03610(.A1(new_n3667_), .A2(new_n3666_), .A3(new_n2905_), .ZN(new_n3681_));
  OAI21_X1   g03611(.A1(new_n3388_), .A2(new_n3389_), .B(new_n2899_), .ZN(new_n3682_));
  AOI22_X1   g03612(.A1(new_n3680_), .A2(new_n3679_), .B1(new_n3681_), .B2(new_n3682_), .ZN(new_n3683_));
  NAND2_X1   g03613(.A1(new_n3680_), .A2(new_n3679_), .ZN(new_n3684_));
  AOI21_X1   g03614(.A1(new_n3667_), .A2(new_n3666_), .B(new_n2899_), .ZN(new_n3685_));
  NOR3_X1    g03615(.A1(new_n3388_), .A2(new_n3389_), .A3(new_n2905_), .ZN(new_n3686_));
  NOR2_X1    g03616(.A1(new_n3686_), .A2(new_n3685_), .ZN(new_n3687_));
  NOR2_X1    g03617(.A1(new_n3684_), .A2(new_n3687_), .ZN(new_n3688_));
  NOR3_X1    g03618(.A1(new_n3688_), .A2(new_n451_), .A3(new_n3683_), .ZN(new_n3689_));
  AOI21_X1   g03619(.A1(new_n3673_), .A2(new_n3669_), .B(\a[2] ), .ZN(new_n3690_));
  NOR2_X1    g03620(.A1(new_n3689_), .A2(new_n3690_), .ZN(new_n3691_));
  NOR3_X1    g03621(.A1(new_n3691_), .A2(new_n3338_), .A3(new_n3341_), .ZN(new_n3692_));
  NOR2_X1    g03622(.A1(new_n3677_), .A2(new_n3692_), .ZN(new_n3693_));
  NAND2_X1   g03623(.A1(new_n3693_), .A2(new_n3664_), .ZN(new_n3694_));
  OAI21_X1   g03624(.A1(new_n3693_), .A2(new_n3664_), .B(new_n3413_), .ZN(new_n3695_));
  NAND2_X1   g03625(.A1(new_n3695_), .A2(new_n3694_), .ZN(new_n3696_));
  NOR2_X1    g03626(.A1(new_n3696_), .A2(new_n3655_), .ZN(new_n3697_));
  NAND2_X1   g03627(.A1(new_n3697_), .A2(new_n3403_), .ZN(new_n3698_));
  XNOR2_X1   g03628(.A1(new_n3396_), .A2(new_n3674_), .ZN(new_n3699_));
  NAND2_X1   g03629(.A1(new_n3699_), .A2(\a[2] ), .ZN(new_n3700_));
  NOR2_X1    g03630(.A1(new_n3700_), .A2(new_n3412_), .ZN(new_n3701_));
  OAI21_X1   g03631(.A1(new_n3697_), .A2(new_n3403_), .B(new_n3701_), .ZN(new_n3702_));
  NAND2_X1   g03632(.A1(new_n3702_), .A2(new_n3698_), .ZN(new_n3703_));
  AOI21_X1   g03633(.A1(new_n2460_), .A2(new_n2461_), .B(new_n2459_), .ZN(new_n3704_));
  NOR3_X1    g03634(.A1(new_n2457_), .A2(new_n2411_), .A3(new_n2029_), .ZN(new_n3705_));
  OAI21_X1   g03635(.A1(new_n3705_), .A2(new_n3704_), .B(new_n2496_), .ZN(new_n3706_));
  NOR2_X1    g03636(.A1(new_n2810_), .A2(new_n3706_), .ZN(new_n3707_));
  NAND3_X1   g03637(.A1(new_n2481_), .A2(new_n2476_), .A3(new_n2470_), .ZN(new_n3708_));
  NAND3_X1   g03638(.A1(new_n2812_), .A2(new_n3708_), .A3(new_n2473_), .ZN(new_n3709_));
  NAND2_X1   g03639(.A1(new_n3684_), .A2(new_n3709_), .ZN(new_n3710_));
  AOI21_X1   g03640(.A1(new_n2458_), .A2(new_n2462_), .B(new_n2470_), .ZN(new_n3711_));
  NOR3_X1    g03641(.A1(new_n3710_), .A2(new_n3711_), .A3(new_n2483_), .ZN(new_n3712_));
  OAI21_X1   g03642(.A1(new_n3712_), .A2(new_n3707_), .B(new_n2812_), .ZN(new_n3713_));
  OAI21_X1   g03643(.A1(new_n2483_), .A2(new_n3710_), .B(new_n3711_), .ZN(new_n3714_));
  NAND2_X1   g03644(.A1(new_n2810_), .A2(new_n3706_), .ZN(new_n3715_));
  NAND3_X1   g03645(.A1(new_n3714_), .A2(new_n3715_), .A3(new_n2808_), .ZN(new_n3716_));
  AOI21_X1   g03646(.A1(new_n3713_), .A2(new_n3716_), .B(new_n3045_), .ZN(new_n3717_));
  AOI21_X1   g03647(.A1(new_n3714_), .A2(new_n3715_), .B(new_n2808_), .ZN(new_n3718_));
  NOR3_X1    g03648(.A1(new_n3712_), .A2(new_n3707_), .A3(new_n2812_), .ZN(new_n3719_));
  NOR3_X1    g03649(.A1(new_n3718_), .A2(new_n3719_), .A3(new_n3044_), .ZN(new_n3720_));
  OAI21_X1   g03650(.A1(new_n3717_), .A2(new_n3720_), .B(new_n451_), .ZN(new_n3721_));
  OAI21_X1   g03651(.A1(new_n3718_), .A2(new_n3719_), .B(new_n3044_), .ZN(new_n3722_));
  NAND3_X1   g03652(.A1(new_n3713_), .A2(new_n3716_), .A3(new_n3045_), .ZN(new_n3723_));
  NAND3_X1   g03653(.A1(new_n3722_), .A2(new_n3723_), .A3(\a[2] ), .ZN(new_n3724_));
  NAND2_X1   g03654(.A1(new_n3721_), .A2(new_n3724_), .ZN(new_n3725_));
  AOI21_X1   g03655(.A1(new_n3713_), .A2(new_n3716_), .B(new_n3044_), .ZN(new_n3726_));
  NOR3_X1    g03656(.A1(new_n3718_), .A2(new_n3719_), .A3(new_n3045_), .ZN(new_n3727_));
  NOR2_X1    g03657(.A1(new_n3727_), .A2(new_n451_), .ZN(new_n3728_));
  NOR2_X1    g03658(.A1(new_n3728_), .A2(new_n3726_), .ZN(new_n3729_));
  AND2_X2    g03659(.A1(new_n2814_), .A2(new_n2811_), .Z(new_n3730_));
  NOR3_X1    g03660(.A1(new_n2889_), .A2(new_n2892_), .A3(new_n2905_), .ZN(new_n3731_));
  NOR3_X1    g03661(.A1(new_n2887_), .A2(new_n2886_), .A3(new_n2470_), .ZN(new_n3732_));
  AOI21_X1   g03662(.A1(new_n2880_), .A2(new_n2884_), .B(new_n2496_), .ZN(new_n3733_));
  OAI21_X1   g03663(.A1(new_n3732_), .A2(new_n3733_), .B(new_n2820_), .ZN(new_n3734_));
  AOI21_X1   g03664(.A1(new_n2880_), .A2(new_n2884_), .B(new_n2470_), .ZN(new_n3735_));
  OAI21_X1   g03665(.A1(new_n2903_), .A2(new_n3735_), .B(new_n2821_), .ZN(new_n3736_));
  AOI21_X1   g03666(.A1(new_n3736_), .A2(new_n3734_), .B(new_n2899_), .ZN(new_n3737_));
  NOR2_X1    g03667(.A1(new_n3737_), .A2(new_n3731_), .ZN(new_n3738_));
  NOR2_X1    g03668(.A1(new_n3738_), .A2(new_n3730_), .ZN(new_n3739_));
  INV_X1     g03669(.I(new_n2901_), .ZN(new_n3740_));
  NAND2_X1   g03670(.A1(new_n3740_), .A2(new_n2900_), .ZN(new_n3741_));
  AOI21_X1   g03671(.A1(new_n3730_), .A2(new_n3741_), .B(new_n3739_), .ZN(new_n3742_));
  NAND2_X1   g03672(.A1(new_n3729_), .A2(new_n3742_), .ZN(new_n3743_));
  OAI21_X1   g03673(.A1(new_n3731_), .A2(new_n3737_), .B(new_n2815_), .ZN(new_n3744_));
  INV_X1     g03674(.I(new_n2900_), .ZN(new_n3745_));
  NOR2_X1    g03675(.A1(new_n3745_), .A2(new_n2901_), .ZN(new_n3746_));
  OAI21_X1   g03676(.A1(new_n3746_), .A2(new_n2815_), .B(new_n3744_), .ZN(new_n3747_));
  OAI21_X1   g03677(.A1(new_n3726_), .A2(new_n3728_), .B(new_n3747_), .ZN(new_n3748_));
  NAND2_X1   g03678(.A1(new_n3743_), .A2(new_n3748_), .ZN(new_n3749_));
  NOR2_X1    g03679(.A1(new_n3749_), .A2(new_n3725_), .ZN(new_n3750_));
  NOR2_X1    g03680(.A1(new_n3397_), .A2(new_n3395_), .ZN(new_n3751_));
  NOR2_X1    g03681(.A1(new_n3751_), .A2(new_n2953_), .ZN(new_n3752_));
  AOI21_X1   g03682(.A1(new_n3751_), .A2(new_n2953_), .B(new_n452_), .ZN(new_n3753_));
  NOR2_X1    g03683(.A1(new_n3753_), .A2(new_n3752_), .ZN(new_n3754_));
  NAND2_X1   g03684(.A1(new_n3749_), .A2(new_n3725_), .ZN(new_n3755_));
  AOI21_X1   g03685(.A1(new_n3754_), .A2(new_n3755_), .B(new_n3750_), .ZN(new_n3756_));
  NAND2_X1   g03686(.A1(new_n3756_), .A2(new_n3703_), .ZN(new_n3757_));
  NAND2_X1   g03687(.A1(new_n3729_), .A2(new_n3747_), .ZN(new_n3758_));
  INV_X1     g03688(.I(new_n3758_), .ZN(new_n3759_));
  NAND2_X1   g03689(.A1(new_n2949_), .A2(new_n2902_), .ZN(new_n3760_));
  NAND2_X1   g03690(.A1(new_n3760_), .A2(new_n3759_), .ZN(new_n3761_));
  OAI21_X1   g03691(.A1(new_n3757_), .A2(new_n3761_), .B(new_n2951_), .ZN(new_n3762_));
  NOR2_X1    g03692(.A1(new_n2933_), .A2(new_n2938_), .ZN(new_n3763_));
  AOI21_X1   g03693(.A1(new_n2470_), .A2(new_n2939_), .B(new_n3763_), .ZN(new_n3764_));
  OAI21_X1   g03694(.A1(new_n1032_), .A2(new_n1029_), .B(new_n443_), .ZN(new_n3765_));
  XNOR2_X1   g03695(.A1(new_n914_), .A2(new_n1027_), .ZN(new_n3766_));
  NAND2_X1   g03696(.A1(new_n3766_), .A2(new_n568_), .ZN(new_n3767_));
  NAND2_X1   g03697(.A1(new_n3767_), .A2(new_n3765_), .ZN(new_n3768_));
  NAND2_X1   g03698(.A1(new_n2915_), .A2(new_n568_), .ZN(new_n3769_));
  NAND2_X1   g03699(.A1(new_n3769_), .A2(new_n2916_), .ZN(new_n3770_));
  XNOR2_X1   g03700(.A1(new_n3770_), .A2(new_n1852_), .ZN(new_n3771_));
  XOR2_X1    g03701(.A1(new_n3771_), .A2(new_n3768_), .Z(new_n3772_));
  NOR2_X1    g03702(.A1(new_n3772_), .A2(\a[14] ), .ZN(new_n3773_));
  AND2_X2    g03703(.A1(new_n3772_), .A2(\a[14] ), .Z(new_n3774_));
  NOR2_X1    g03704(.A1(new_n3774_), .A2(new_n3773_), .ZN(new_n3775_));
  AOI21_X1   g03705(.A1(new_n2920_), .A2(new_n2922_), .B(new_n2924_), .ZN(new_n3776_));
  NAND2_X1   g03706(.A1(new_n3775_), .A2(new_n3776_), .ZN(new_n3777_));
  INV_X1     g03707(.I(new_n3776_), .ZN(new_n3778_));
  OAI21_X1   g03708(.A1(new_n3774_), .A2(new_n3773_), .B(new_n3778_), .ZN(new_n3779_));
  AOI21_X1   g03709(.A1(new_n3777_), .A2(new_n3779_), .B(new_n806_), .ZN(new_n3780_));
  XOR2_X1    g03710(.A1(new_n3775_), .A2(new_n3778_), .Z(new_n3781_));
  NOR2_X1    g03711(.A1(new_n3781_), .A2(new_n1079_), .ZN(new_n3782_));
  NOR2_X1    g03712(.A1(new_n3782_), .A2(new_n3780_), .ZN(new_n3783_));
  NOR2_X1    g03713(.A1(new_n2928_), .A2(new_n1079_), .ZN(new_n3784_));
  NOR2_X1    g03714(.A1(new_n3784_), .A2(new_n2929_), .ZN(new_n3785_));
  NAND2_X1   g03715(.A1(new_n3783_), .A2(new_n3785_), .ZN(new_n3786_));
  OAI22_X1   g03716(.A1(new_n3782_), .A2(new_n3780_), .B1(new_n2929_), .B2(new_n3784_), .ZN(new_n3787_));
  AOI21_X1   g03717(.A1(new_n3786_), .A2(new_n3787_), .B(new_n2496_), .ZN(new_n3788_));
  XOR2_X1    g03718(.A1(new_n3783_), .A2(new_n3785_), .Z(new_n3789_));
  AOI21_X1   g03719(.A1(new_n3789_), .A2(new_n2496_), .B(new_n3788_), .ZN(new_n3790_));
  XOR2_X1    g03720(.A1(new_n3790_), .A2(new_n3764_), .Z(new_n3791_));
  XOR2_X1    g03721(.A1(new_n3791_), .A2(new_n452_), .Z(new_n3792_));
  NOR2_X1    g03722(.A1(new_n2946_), .A2(new_n2904_), .ZN(new_n3793_));
  NOR2_X1    g03723(.A1(new_n3793_), .A2(new_n2947_), .ZN(new_n3794_));
  NAND2_X1   g03724(.A1(new_n3792_), .A2(new_n3794_), .ZN(new_n3795_));
  NAND2_X1   g03725(.A1(new_n3762_), .A2(new_n3795_), .ZN(new_n3796_));
  OR2_X2     g03726(.A1(new_n3792_), .A2(new_n3794_), .Z(new_n3797_));
  NAND2_X1   g03727(.A1(new_n3796_), .A2(new_n3797_), .ZN(new_n3798_));
  NAND2_X1   g03728(.A1(new_n3786_), .A2(new_n2470_), .ZN(new_n3799_));
  NAND2_X1   g03729(.A1(new_n3799_), .A2(new_n3787_), .ZN(new_n3800_));
  NAND2_X1   g03730(.A1(new_n3777_), .A2(new_n1079_), .ZN(new_n3801_));
  NAND2_X1   g03731(.A1(new_n3801_), .A2(new_n3779_), .ZN(new_n3802_));
  INV_X1     g03732(.I(new_n3768_), .ZN(new_n3803_));
  INV_X1     g03733(.I(new_n3770_), .ZN(new_n3804_));
  AOI21_X1   g03734(.A1(new_n3803_), .A2(new_n3804_), .B(new_n1853_), .ZN(new_n3805_));
  AOI21_X1   g03735(.A1(new_n3768_), .A2(new_n3770_), .B(new_n3805_), .ZN(new_n3806_));
  XNOR2_X1   g03736(.A1(new_n910_), .A2(new_n1033_), .ZN(new_n3807_));
  OAI21_X1   g03737(.A1(new_n1035_), .A2(new_n1037_), .B(new_n443_), .ZN(new_n3808_));
  OAI21_X1   g03738(.A1(new_n443_), .A2(new_n3807_), .B(new_n3808_), .ZN(new_n3809_));
  XOR2_X1    g03739(.A1(new_n3809_), .A2(new_n3806_), .Z(new_n3810_));
  NAND2_X1   g03740(.A1(new_n3810_), .A2(new_n786_), .ZN(new_n3811_));
  NOR2_X1    g03741(.A1(new_n3809_), .A2(new_n3806_), .ZN(new_n3812_));
  NAND2_X1   g03742(.A1(new_n3809_), .A2(new_n3806_), .ZN(new_n3813_));
  INV_X1     g03743(.I(new_n3813_), .ZN(new_n3814_));
  OAI21_X1   g03744(.A1(new_n3814_), .A2(new_n3812_), .B(new_n644_), .ZN(new_n3815_));
  NAND2_X1   g03745(.A1(new_n3811_), .A2(new_n3815_), .ZN(new_n3816_));
  XOR2_X1    g03746(.A1(new_n3816_), .A2(new_n806_), .Z(new_n3817_));
  INV_X1     g03747(.I(new_n3817_), .ZN(new_n3818_));
  NAND3_X1   g03748(.A1(new_n3811_), .A2(new_n806_), .A3(new_n3815_), .ZN(new_n3819_));
  NAND2_X1   g03749(.A1(new_n3816_), .A2(new_n1079_), .ZN(new_n3820_));
  AOI21_X1   g03750(.A1(new_n3819_), .A2(new_n3820_), .B(new_n3802_), .ZN(new_n3821_));
  AOI21_X1   g03751(.A1(new_n3802_), .A2(new_n3818_), .B(new_n3821_), .ZN(new_n3822_));
  XOR2_X1    g03752(.A1(new_n3800_), .A2(new_n3822_), .Z(new_n3823_));
  XOR2_X1    g03753(.A1(new_n3823_), .A2(new_n498_), .Z(new_n3824_));
  INV_X1     g03754(.I(new_n3824_), .ZN(new_n3825_));
  NOR2_X1    g03755(.A1(new_n3790_), .A2(new_n3764_), .ZN(new_n3826_));
  AOI21_X1   g03756(.A1(new_n3790_), .A2(new_n3764_), .B(new_n452_), .ZN(new_n3827_));
  NOR2_X1    g03757(.A1(new_n3827_), .A2(new_n3826_), .ZN(new_n3828_));
  NAND2_X1   g03758(.A1(new_n3825_), .A2(new_n3828_), .ZN(new_n3829_));
  NAND2_X1   g03759(.A1(new_n3798_), .A2(new_n3829_), .ZN(new_n3830_));
  OAI21_X1   g03760(.A1(new_n3826_), .A2(new_n3827_), .B(new_n3824_), .ZN(new_n3831_));
  NAND2_X1   g03761(.A1(new_n3830_), .A2(new_n3831_), .ZN(new_n3832_));
  OAI21_X1   g03762(.A1(new_n1040_), .A2(new_n1042_), .B(new_n786_), .ZN(new_n3833_));
  XNOR2_X1   g03763(.A1(new_n906_), .A2(new_n1038_), .ZN(new_n3834_));
  OAI21_X1   g03764(.A1(new_n3834_), .A2(new_n786_), .B(new_n3833_), .ZN(new_n3835_));
  NOR2_X1    g03765(.A1(new_n3814_), .A2(new_n644_), .ZN(new_n3836_));
  NOR3_X1    g03766(.A1(new_n3835_), .A2(new_n3812_), .A3(new_n3836_), .ZN(new_n3837_));
  INV_X1     g03767(.I(new_n3835_), .ZN(new_n3838_));
  NOR2_X1    g03768(.A1(new_n3836_), .A2(new_n3812_), .ZN(new_n3839_));
  NOR2_X1    g03769(.A1(new_n3838_), .A2(new_n3839_), .ZN(new_n3840_));
  NOR2_X1    g03770(.A1(new_n3840_), .A2(new_n3837_), .ZN(new_n3841_));
  NOR2_X1    g03771(.A1(new_n3841_), .A2(new_n1079_), .ZN(new_n3842_));
  XOR2_X1    g03772(.A1(new_n3835_), .A2(new_n3839_), .Z(new_n3843_));
  NOR2_X1    g03773(.A1(new_n3843_), .A2(new_n806_), .ZN(new_n3844_));
  NOR2_X1    g03774(.A1(new_n3842_), .A2(new_n3844_), .ZN(new_n3845_));
  NAND2_X1   g03775(.A1(new_n3802_), .A2(new_n3820_), .ZN(new_n3846_));
  NAND2_X1   g03776(.A1(new_n3846_), .A2(new_n3819_), .ZN(new_n3847_));
  XOR2_X1    g03777(.A1(new_n3845_), .A2(new_n3847_), .Z(new_n3848_));
  NOR2_X1    g03778(.A1(new_n3848_), .A2(new_n2470_), .ZN(new_n3849_));
  INV_X1     g03779(.I(new_n3845_), .ZN(new_n3850_));
  NOR2_X1    g03780(.A1(new_n3850_), .A2(new_n3847_), .ZN(new_n3851_));
  INV_X1     g03781(.I(new_n3851_), .ZN(new_n3852_));
  NAND2_X1   g03782(.A1(new_n3850_), .A2(new_n3847_), .ZN(new_n3853_));
  AOI21_X1   g03783(.A1(new_n3852_), .A2(new_n3853_), .B(new_n2496_), .ZN(new_n3854_));
  NOR2_X1    g03784(.A1(new_n3854_), .A2(new_n3849_), .ZN(new_n3855_));
  INV_X1     g03785(.I(new_n3855_), .ZN(new_n3856_));
  INV_X1     g03786(.I(new_n3800_), .ZN(new_n3857_));
  NOR2_X1    g03787(.A1(new_n3857_), .A2(new_n3822_), .ZN(new_n3858_));
  AOI21_X1   g03788(.A1(new_n3857_), .A2(new_n3822_), .B(\a[8] ), .ZN(new_n3859_));
  NOR2_X1    g03789(.A1(new_n3859_), .A2(new_n3858_), .ZN(new_n3860_));
  NAND2_X1   g03790(.A1(new_n3856_), .A2(new_n3860_), .ZN(new_n3861_));
  NAND2_X1   g03791(.A1(new_n3832_), .A2(new_n3861_), .ZN(new_n3862_));
  NOR2_X1    g03792(.A1(new_n3856_), .A2(new_n3860_), .ZN(new_n3863_));
  INV_X1     g03793(.I(new_n3863_), .ZN(new_n3864_));
  NAND2_X1   g03794(.A1(new_n3862_), .A2(new_n3864_), .ZN(new_n3865_));
  OAI21_X1   g03795(.A1(new_n2470_), .A2(new_n3851_), .B(new_n3853_), .ZN(new_n3866_));
  XOR2_X1    g03796(.A1(new_n1049_), .A2(new_n1071_), .Z(new_n3867_));
  XOR2_X1    g03797(.A1(new_n3867_), .A2(\a[11] ), .Z(new_n3868_));
  AOI21_X1   g03798(.A1(new_n1046_), .A2(new_n1047_), .B(new_n1079_), .ZN(new_n3869_));
  XOR2_X1    g03799(.A1(new_n1043_), .A2(new_n901_), .Z(new_n3870_));
  NOR2_X1    g03800(.A1(new_n3870_), .A2(new_n806_), .ZN(new_n3871_));
  NOR2_X1    g03801(.A1(new_n3869_), .A2(new_n3871_), .ZN(new_n3872_));
  NOR2_X1    g03802(.A1(new_n3837_), .A2(new_n1079_), .ZN(new_n3873_));
  NOR2_X1    g03803(.A1(new_n3873_), .A2(new_n3840_), .ZN(new_n3874_));
  NOR2_X1    g03804(.A1(new_n3872_), .A2(new_n3874_), .ZN(new_n3875_));
  AOI21_X1   g03805(.A1(new_n3872_), .A2(new_n3874_), .B(new_n498_), .ZN(new_n3876_));
  NOR2_X1    g03806(.A1(new_n3876_), .A2(new_n3875_), .ZN(new_n3877_));
  XOR2_X1    g03807(.A1(new_n3868_), .A2(new_n3877_), .Z(new_n3878_));
  NOR2_X1    g03808(.A1(new_n3878_), .A2(new_n3866_), .ZN(new_n3879_));
  XOR2_X1    g03809(.A1(new_n3872_), .A2(new_n3874_), .Z(new_n3880_));
  XOR2_X1    g03810(.A1(new_n3880_), .A2(new_n498_), .Z(new_n3881_));
  INV_X1     g03811(.I(new_n3881_), .ZN(new_n3882_));
  AOI21_X1   g03812(.A1(new_n3878_), .A2(new_n3866_), .B(new_n3882_), .ZN(new_n3883_));
  NOR2_X1    g03813(.A1(new_n3883_), .A2(new_n3879_), .ZN(new_n3884_));
  NAND2_X1   g03814(.A1(new_n3868_), .A2(new_n3877_), .ZN(new_n3885_));
  INV_X1     g03815(.I(new_n3885_), .ZN(new_n3886_));
  NAND2_X1   g03816(.A1(new_n1104_), .A2(new_n1074_), .ZN(new_n3887_));
  NAND4_X1   g03817(.A1(new_n3865_), .A2(new_n3884_), .A3(new_n3886_), .A4(new_n3887_), .ZN(new_n3888_));
  OAI21_X1   g03818(.A1(new_n1074_), .A2(new_n1104_), .B(new_n3888_), .ZN(new_n3889_));
  INV_X1     g03819(.I(new_n1101_), .ZN(new_n3890_));
  OAI21_X1   g03820(.A1(new_n806_), .A2(new_n1100_), .B(new_n3890_), .ZN(new_n3891_));
  INV_X1     g03821(.I(new_n764_), .ZN(new_n3892_));
  OAI21_X1   g03822(.A1(new_n3892_), .A2(new_n763_), .B(new_n786_), .ZN(new_n3893_));
  XNOR2_X1   g03823(.A1(new_n708_), .A2(new_n762_), .ZN(new_n3894_));
  NAND2_X1   g03824(.A1(new_n3894_), .A2(new_n644_), .ZN(new_n3895_));
  NAND2_X1   g03825(.A1(new_n3893_), .A2(new_n3895_), .ZN(new_n3896_));
  INV_X1     g03826(.I(new_n3896_), .ZN(new_n3897_));
  NOR2_X1    g03827(.A1(new_n1086_), .A2(new_n644_), .ZN(new_n3898_));
  NOR2_X1    g03828(.A1(new_n3898_), .A2(new_n1089_), .ZN(new_n3899_));
  NOR2_X1    g03829(.A1(new_n3897_), .A2(new_n3899_), .ZN(new_n3900_));
  AOI21_X1   g03830(.A1(new_n3897_), .A2(new_n3899_), .B(new_n294_), .ZN(new_n3901_));
  NOR2_X1    g03831(.A1(new_n3901_), .A2(new_n3900_), .ZN(new_n3902_));
  XOR2_X1    g03832(.A1(new_n778_), .A2(new_n786_), .Z(new_n3903_));
  OAI21_X1   g03833(.A1(new_n779_), .A2(new_n787_), .B(new_n766_), .ZN(new_n3904_));
  OAI21_X1   g03834(.A1(new_n3903_), .A2(new_n766_), .B(new_n3904_), .ZN(new_n3905_));
  XOR2_X1    g03835(.A1(new_n3902_), .A2(new_n3905_), .Z(new_n3906_));
  NOR2_X1    g03836(.A1(new_n3906_), .A2(new_n3891_), .ZN(new_n3907_));
  XOR2_X1    g03837(.A1(new_n3896_), .A2(new_n3899_), .Z(new_n3908_));
  XOR2_X1    g03838(.A1(new_n3908_), .A2(\a[11] ), .Z(new_n3909_));
  NAND2_X1   g03839(.A1(new_n3906_), .A2(new_n3891_), .ZN(new_n3910_));
  AOI21_X1   g03840(.A1(new_n3909_), .A2(new_n3910_), .B(new_n3907_), .ZN(new_n3911_));
  NAND2_X1   g03841(.A1(new_n3902_), .A2(new_n3905_), .ZN(new_n3912_));
  INV_X1     g03842(.I(new_n3912_), .ZN(new_n3913_));
  OR4_X2     g03843(.A1(new_n780_), .A2(new_n794_), .A3(new_n787_), .A4(new_n798_), .Z(new_n3914_));
  NAND4_X1   g03844(.A1(new_n3889_), .A2(new_n3911_), .A3(new_n3913_), .A4(new_n3914_), .ZN(new_n3915_));
  NAND2_X1   g03845(.A1(new_n3915_), .A2(new_n799_), .ZN(new_n3916_));
  INV_X1     g03846(.I(new_n3916_), .ZN(new_n3917_));
  OAI21_X1   g03847(.A1(new_n786_), .A2(new_n795_), .B(new_n797_), .ZN(new_n3918_));
  XOR2_X1    g03848(.A1(new_n629_), .A2(new_n634_), .Z(new_n3919_));
  NOR2_X1    g03849(.A1(new_n3919_), .A2(new_n3918_), .ZN(new_n3920_));
  XOR2_X1    g03850(.A1(new_n626_), .A2(new_n576_), .Z(new_n3921_));
  XOR2_X1    g03851(.A1(new_n3921_), .A2(\a[14] ), .Z(new_n3922_));
  AOI21_X1   g03852(.A1(new_n3918_), .A2(new_n3919_), .B(new_n3922_), .ZN(new_n3923_));
  NOR3_X1    g03853(.A1(new_n3917_), .A2(new_n3920_), .A3(new_n3923_), .ZN(new_n3924_));
  OAI21_X1   g03854(.A1(new_n427_), .A2(new_n429_), .B(new_n273_), .ZN(new_n3925_));
  INV_X1     g03855(.I(new_n3925_), .ZN(new_n3926_));
  XOR2_X1    g03856(.A1(new_n391_), .A2(new_n425_), .Z(new_n3927_));
  AOI21_X1   g03857(.A1(new_n3927_), .A2(new_n356_), .B(new_n3926_), .ZN(new_n3928_));
  NOR2_X1    g03858(.A1(new_n562_), .A2(new_n356_), .ZN(new_n3929_));
  NOR2_X1    g03859(.A1(new_n3929_), .A2(new_n560_), .ZN(new_n3930_));
  INV_X1     g03860(.I(new_n3930_), .ZN(new_n3931_));
  NOR2_X1    g03861(.A1(new_n3931_), .A2(new_n443_), .ZN(new_n3932_));
  NOR2_X1    g03862(.A1(new_n3930_), .A2(new_n568_), .ZN(new_n3933_));
  NOR2_X1    g03863(.A1(new_n3932_), .A2(new_n3933_), .ZN(new_n3934_));
  NOR2_X1    g03864(.A1(new_n3934_), .A2(new_n3928_), .ZN(new_n3935_));
  XOR2_X1    g03865(.A1(new_n3930_), .A2(new_n568_), .Z(new_n3936_));
  AOI21_X1   g03866(.A1(new_n3928_), .A2(new_n3936_), .B(new_n3935_), .ZN(new_n3937_));
  NOR2_X1    g03867(.A1(new_n636_), .A2(new_n571_), .ZN(new_n3938_));
  NOR2_X1    g03868(.A1(new_n3938_), .A2(new_n3937_), .ZN(new_n3939_));
  NAND2_X1   g03869(.A1(new_n3924_), .A2(new_n3939_), .ZN(new_n3940_));
  NAND2_X1   g03870(.A1(new_n3940_), .A2(new_n637_), .ZN(new_n3941_));
  INV_X1     g03871(.I(new_n3933_), .ZN(new_n3942_));
  OAI21_X1   g03872(.A1(new_n3928_), .A2(new_n3932_), .B(new_n3942_), .ZN(new_n3943_));
  XOR2_X1    g03873(.A1(new_n433_), .A2(new_n437_), .Z(new_n3944_));
  NOR2_X1    g03874(.A1(new_n3944_), .A2(new_n3943_), .ZN(new_n3945_));
  XNOR2_X1   g03875(.A1(new_n387_), .A2(new_n430_), .ZN(new_n3946_));
  XOR2_X1    g03876(.A1(new_n3946_), .A2(\a[17] ), .Z(new_n3947_));
  NAND2_X1   g03877(.A1(new_n3944_), .A2(new_n3943_), .ZN(new_n3948_));
  AOI21_X1   g03878(.A1(new_n3947_), .A2(new_n3948_), .B(new_n3945_), .ZN(new_n3949_));
  OAI21_X1   g03879(.A1(new_n219_), .A2(new_n221_), .B(new_n118_), .ZN(new_n3950_));
  XNOR2_X1   g03880(.A1(new_n217_), .A2(new_n201_), .ZN(new_n3951_));
  OAI21_X1   g03881(.A1(new_n118_), .A2(new_n3951_), .B(new_n3950_), .ZN(new_n3952_));
  OAI21_X1   g03882(.A1(new_n71_), .A2(new_n366_), .B(new_n368_), .ZN(new_n3953_));
  NOR2_X1    g03883(.A1(new_n3953_), .A2(new_n3952_), .ZN(new_n3954_));
  INV_X1     g03884(.I(new_n3954_), .ZN(new_n3955_));
  NAND2_X1   g03885(.A1(new_n3953_), .A2(new_n3952_), .ZN(new_n3956_));
  AOI21_X1   g03886(.A1(new_n3955_), .A2(new_n3956_), .B(new_n189_), .ZN(new_n3957_));
  XNOR2_X1   g03887(.A1(new_n3953_), .A2(new_n3952_), .ZN(new_n3958_));
  NOR2_X1    g03888(.A1(new_n3958_), .A2(new_n248_), .ZN(new_n3959_));
  NOR2_X1    g03889(.A1(new_n3959_), .A2(new_n3957_), .ZN(new_n3960_));
  INV_X1     g03890(.I(new_n376_), .ZN(new_n3961_));
  AOI21_X1   g03891(.A1(new_n248_), .A2(new_n3961_), .B(new_n375_), .ZN(new_n3962_));
  AND2_X2    g03892(.A1(new_n3962_), .A2(new_n273_), .Z(new_n3963_));
  NOR2_X1    g03893(.A1(new_n3962_), .A2(new_n273_), .ZN(new_n3964_));
  NOR2_X1    g03894(.A1(new_n3963_), .A2(new_n3964_), .ZN(new_n3965_));
  NOR2_X1    g03895(.A1(new_n3965_), .A2(new_n3960_), .ZN(new_n3966_));
  INV_X1     g03896(.I(new_n3960_), .ZN(new_n3967_));
  XOR2_X1    g03897(.A1(new_n3962_), .A2(new_n356_), .Z(new_n3968_));
  NOR2_X1    g03898(.A1(new_n3968_), .A2(new_n3967_), .ZN(new_n3969_));
  NOR2_X1    g03899(.A1(new_n3966_), .A2(new_n3969_), .ZN(new_n3970_));
  AOI21_X1   g03900(.A1(new_n438_), .A2(new_n383_), .B(new_n3970_), .ZN(new_n3971_));
  NAND3_X1   g03901(.A1(new_n3941_), .A2(new_n3949_), .A3(new_n3971_), .ZN(new_n3972_));
  OAI21_X1   g03902(.A1(new_n383_), .A2(new_n438_), .B(new_n3972_), .ZN(new_n3973_));
  INV_X1     g03903(.I(new_n3963_), .ZN(new_n3974_));
  AOI21_X1   g03904(.A1(new_n3974_), .A2(new_n3967_), .B(new_n3964_), .ZN(new_n3975_));
  NOR2_X1    g03905(.A1(new_n250_), .A2(new_n240_), .ZN(new_n3976_));
  XOR2_X1    g03906(.A1(new_n249_), .A2(new_n248_), .Z(new_n3977_));
  NAND2_X1   g03907(.A1(new_n3977_), .A2(new_n228_), .ZN(new_n3978_));
  OAI21_X1   g03908(.A1(new_n228_), .A2(new_n3976_), .B(new_n3978_), .ZN(new_n3979_));
  OAI21_X1   g03909(.A1(new_n227_), .A2(new_n224_), .B(new_n248_), .ZN(new_n3980_));
  XOR2_X1    g03910(.A1(new_n226_), .A2(new_n223_), .Z(new_n3981_));
  OAI21_X1   g03911(.A1(new_n3981_), .A2(new_n248_), .B(new_n3980_), .ZN(new_n3982_));
  OAI21_X1   g03912(.A1(new_n189_), .A2(new_n3954_), .B(new_n3956_), .ZN(new_n3983_));
  NAND2_X1   g03913(.A1(new_n3982_), .A2(new_n3983_), .ZN(new_n3984_));
  OAI21_X1   g03914(.A1(new_n3982_), .A2(new_n3983_), .B(\a[20] ), .ZN(new_n3985_));
  NAND2_X1   g03915(.A1(new_n3985_), .A2(new_n3984_), .ZN(new_n3986_));
  XNOR2_X1   g03916(.A1(new_n3979_), .A2(new_n3986_), .ZN(new_n3987_));
  XNOR2_X1   g03917(.A1(new_n3982_), .A2(new_n3983_), .ZN(new_n3988_));
  NOR2_X1    g03918(.A1(new_n3988_), .A2(\a[20] ), .ZN(new_n3989_));
  NAND2_X1   g03919(.A1(new_n3988_), .A2(\a[20] ), .ZN(new_n3990_));
  INV_X1     g03920(.I(new_n3990_), .ZN(new_n3991_));
  NOR2_X1    g03921(.A1(new_n3991_), .A2(new_n3989_), .ZN(new_n3992_));
  INV_X1     g03922(.I(new_n3992_), .ZN(new_n3993_));
  NOR2_X1    g03923(.A1(new_n3987_), .A2(new_n3975_), .ZN(new_n3994_));
  NOR2_X1    g03924(.A1(new_n3994_), .A2(new_n3993_), .ZN(new_n3995_));
  AOI21_X1   g03925(.A1(new_n3975_), .A2(new_n3987_), .B(new_n3995_), .ZN(new_n3996_));
  NAND2_X1   g03926(.A1(new_n3973_), .A2(new_n3996_), .ZN(new_n3997_));
  INV_X1     g03927(.I(new_n3997_), .ZN(new_n3998_));
  NOR2_X1    g03928(.A1(new_n3979_), .A2(new_n3986_), .ZN(new_n3999_));
  INV_X1     g03929(.I(new_n3999_), .ZN(new_n4000_));
  AOI21_X1   g03930(.A1(new_n251_), .A2(new_n266_), .B(new_n4000_), .ZN(new_n4001_));
  AOI21_X1   g03931(.A1(new_n3998_), .A2(new_n4001_), .B(new_n267_), .ZN(new_n4002_));
  INV_X1     g03932(.I(new_n4002_), .ZN(new_n4003_));
  OAI21_X1   g03933(.A1(new_n263_), .A2(new_n259_), .B(new_n261_), .ZN(new_n4004_));
  NOR2_X1    g03934(.A1(new_n145_), .A2(new_n144_), .ZN(new_n4005_));
  XNOR2_X1   g03935(.A1(new_n4005_), .A2(new_n165_), .ZN(new_n4006_));
  NOR2_X1    g03936(.A1(new_n4006_), .A2(new_n4004_), .ZN(new_n4007_));
  XNOR2_X1   g03937(.A1(new_n143_), .A2(new_n121_), .ZN(new_n4008_));
  XOR2_X1    g03938(.A1(new_n4008_), .A2(\a[23] ), .Z(new_n4009_));
  NAND2_X1   g03939(.A1(new_n4006_), .A2(new_n4004_), .ZN(new_n4010_));
  AOI21_X1   g03940(.A1(new_n4009_), .A2(new_n4010_), .B(new_n4007_), .ZN(new_n4011_));
  NAND2_X1   g03941(.A1(new_n4003_), .A2(new_n4011_), .ZN(new_n4012_));
  XNOR2_X1   g03942(.A1(new_n4012_), .A2(new_n184_), .ZN(new_n4013_));
  NOR2_X1    g03943(.A1(new_n4013_), .A2(new_n166_), .ZN(new_n4014_));
  NAND2_X1   g03944(.A1(new_n4013_), .A2(new_n166_), .ZN(new_n4015_));
  INV_X1     g03945(.I(new_n4015_), .ZN(new_n4016_));
  NOR2_X1    g03946(.A1(new_n4016_), .A2(new_n4014_), .ZN(new_n4017_));
  INV_X1     g03947(.I(new_n4017_), .ZN(new_n4018_));
  INV_X1     g03948(.I(new_n4009_), .ZN(new_n4019_));
  NAND2_X1   g03949(.A1(new_n4019_), .A2(new_n4004_), .ZN(new_n4020_));
  XOR2_X1    g03950(.A1(new_n4009_), .A2(new_n4004_), .Z(new_n4021_));
  INV_X1     g03951(.I(new_n4021_), .ZN(new_n4022_));
  NAND2_X1   g03952(.A1(new_n4022_), .A2(new_n4006_), .ZN(new_n4023_));
  XNOR2_X1   g03953(.A1(new_n4023_), .A2(new_n4020_), .ZN(new_n4024_));
  NOR2_X1    g03954(.A1(new_n4003_), .A2(new_n4024_), .ZN(new_n4025_));
  NAND2_X1   g03955(.A1(new_n4003_), .A2(new_n4024_), .ZN(new_n4026_));
  INV_X1     g03956(.I(new_n4026_), .ZN(new_n4027_));
  NOR2_X1    g03957(.A1(new_n4027_), .A2(new_n4025_), .ZN(new_n4028_));
  INV_X1     g03958(.I(new_n4028_), .ZN(new_n4029_));
  NOR2_X1    g03959(.A1(new_n4018_), .A2(new_n4029_), .ZN(new_n4030_));
  INV_X1     g03960(.I(new_n4030_), .ZN(new_n4031_));
  NOR2_X1    g03961(.A1(new_n4002_), .A2(new_n4021_), .ZN(new_n4032_));
  XNOR2_X1   g03962(.A1(new_n4009_), .A2(new_n4004_), .ZN(new_n4033_));
  NOR2_X1    g03963(.A1(new_n4003_), .A2(new_n4033_), .ZN(new_n4034_));
  NOR2_X1    g03964(.A1(new_n4034_), .A2(new_n4032_), .ZN(new_n4035_));
  INV_X1     g03965(.I(new_n4035_), .ZN(new_n4036_));
  NOR2_X1    g03966(.A1(new_n4029_), .A2(new_n4036_), .ZN(new_n4037_));
  XOR2_X1    g03967(.A1(new_n3997_), .A2(new_n267_), .Z(new_n4038_));
  NOR2_X1    g03968(.A1(new_n4038_), .A2(new_n3999_), .ZN(new_n4039_));
  NAND2_X1   g03969(.A1(new_n4038_), .A2(new_n3999_), .ZN(new_n4040_));
  INV_X1     g03970(.I(new_n4040_), .ZN(new_n4041_));
  NOR2_X1    g03971(.A1(new_n4041_), .A2(new_n4039_), .ZN(new_n4042_));
  INV_X1     g03972(.I(new_n4042_), .ZN(new_n4043_));
  NOR2_X1    g03973(.A1(new_n4043_), .A2(new_n4036_), .ZN(new_n4044_));
  INV_X1     g03974(.I(new_n3975_), .ZN(new_n4045_));
  NAND2_X1   g03975(.A1(new_n3993_), .A2(new_n4045_), .ZN(new_n4046_));
  XOR2_X1    g03976(.A1(new_n3992_), .A2(new_n4045_), .Z(new_n4047_));
  NOR2_X1    g03977(.A1(new_n4047_), .A2(new_n3987_), .ZN(new_n4048_));
  XOR2_X1    g03978(.A1(new_n4048_), .A2(new_n4046_), .Z(new_n4049_));
  NOR2_X1    g03979(.A1(new_n3973_), .A2(new_n4049_), .ZN(new_n4050_));
  NAND2_X1   g03980(.A1(new_n3973_), .A2(new_n4049_), .ZN(new_n4051_));
  INV_X1     g03981(.I(new_n4051_), .ZN(new_n4052_));
  NOR2_X1    g03982(.A1(new_n4052_), .A2(new_n4050_), .ZN(new_n4053_));
  INV_X1     g03983(.I(new_n4053_), .ZN(new_n4054_));
  NOR2_X1    g03984(.A1(new_n4043_), .A2(new_n4054_), .ZN(new_n4055_));
  INV_X1     g03985(.I(new_n3973_), .ZN(new_n4056_));
  NOR2_X1    g03986(.A1(new_n4056_), .A2(new_n4047_), .ZN(new_n4057_));
  NAND2_X1   g03987(.A1(new_n3992_), .A2(new_n3975_), .ZN(new_n4058_));
  AOI21_X1   g03988(.A1(new_n4046_), .A2(new_n4058_), .B(new_n3973_), .ZN(new_n4059_));
  NOR2_X1    g03989(.A1(new_n4057_), .A2(new_n4059_), .ZN(new_n4060_));
  INV_X1     g03990(.I(new_n4060_), .ZN(new_n4061_));
  NOR2_X1    g03991(.A1(new_n4061_), .A2(new_n4054_), .ZN(new_n4062_));
  INV_X1     g03992(.I(new_n438_), .ZN(new_n4063_));
  NAND2_X1   g03993(.A1(new_n3941_), .A2(new_n3949_), .ZN(new_n4064_));
  NOR2_X1    g03994(.A1(new_n383_), .A2(new_n3970_), .ZN(new_n4065_));
  XOR2_X1    g03995(.A1(new_n4064_), .A2(new_n4065_), .Z(new_n4066_));
  NOR2_X1    g03996(.A1(new_n4066_), .A2(new_n4063_), .ZN(new_n4067_));
  NAND2_X1   g03997(.A1(new_n4066_), .A2(new_n4063_), .ZN(new_n4068_));
  INV_X1     g03998(.I(new_n4068_), .ZN(new_n4069_));
  NOR2_X1    g03999(.A1(new_n4069_), .A2(new_n4067_), .ZN(new_n4070_));
  INV_X1     g04000(.I(new_n4070_), .ZN(new_n4071_));
  NOR2_X1    g04001(.A1(new_n4071_), .A2(new_n4061_), .ZN(new_n4072_));
  INV_X1     g04002(.I(new_n3943_), .ZN(new_n4073_));
  NOR2_X1    g04003(.A1(new_n4073_), .A2(new_n3947_), .ZN(new_n4074_));
  XNOR2_X1   g04004(.A1(new_n3947_), .A2(new_n3943_), .ZN(new_n4075_));
  NAND2_X1   g04005(.A1(new_n4075_), .A2(new_n3944_), .ZN(new_n4076_));
  XOR2_X1    g04006(.A1(new_n4076_), .A2(new_n4074_), .Z(new_n4077_));
  NOR2_X1    g04007(.A1(new_n3941_), .A2(new_n4077_), .ZN(new_n4078_));
  NAND2_X1   g04008(.A1(new_n3941_), .A2(new_n4077_), .ZN(new_n4079_));
  INV_X1     g04009(.I(new_n4079_), .ZN(new_n4080_));
  NOR2_X1    g04010(.A1(new_n4080_), .A2(new_n4078_), .ZN(new_n4081_));
  INV_X1     g04011(.I(new_n4081_), .ZN(new_n4082_));
  NOR2_X1    g04012(.A1(new_n4071_), .A2(new_n4082_), .ZN(new_n4083_));
  INV_X1     g04013(.I(new_n4083_), .ZN(new_n4084_));
  NOR2_X1    g04014(.A1(new_n3937_), .A2(new_n570_), .ZN(new_n4085_));
  XNOR2_X1   g04015(.A1(new_n3924_), .A2(new_n4085_), .ZN(new_n4086_));
  NOR2_X1    g04016(.A1(new_n4086_), .A2(new_n636_), .ZN(new_n4087_));
  NAND2_X1   g04017(.A1(new_n4086_), .A2(new_n636_), .ZN(new_n4088_));
  INV_X1     g04018(.I(new_n4088_), .ZN(new_n4089_));
  NOR2_X1    g04019(.A1(new_n4089_), .A2(new_n4087_), .ZN(new_n4090_));
  INV_X1     g04020(.I(new_n4090_), .ZN(new_n4091_));
  NAND2_X1   g04021(.A1(new_n3922_), .A2(new_n3918_), .ZN(new_n4092_));
  XOR2_X1    g04022(.A1(new_n3922_), .A2(new_n3918_), .Z(new_n4093_));
  NAND2_X1   g04023(.A1(new_n4093_), .A2(new_n3919_), .ZN(new_n4094_));
  XNOR2_X1   g04024(.A1(new_n4094_), .A2(new_n4092_), .ZN(new_n4095_));
  NOR2_X1    g04025(.A1(new_n3916_), .A2(new_n4095_), .ZN(new_n4096_));
  NAND2_X1   g04026(.A1(new_n3916_), .A2(new_n4095_), .ZN(new_n4097_));
  INV_X1     g04027(.I(new_n4097_), .ZN(new_n4098_));
  NOR2_X1    g04028(.A1(new_n4098_), .A2(new_n4096_), .ZN(new_n4099_));
  INV_X1     g04029(.I(new_n4099_), .ZN(new_n4100_));
  NOR2_X1    g04030(.A1(new_n4091_), .A2(new_n4100_), .ZN(new_n4101_));
  INV_X1     g04031(.I(new_n4101_), .ZN(new_n4102_));
  NAND2_X1   g04032(.A1(new_n3916_), .A2(new_n4093_), .ZN(new_n4103_));
  XOR2_X1    g04033(.A1(new_n3922_), .A2(new_n3918_), .Z(new_n4104_));
  OAI21_X1   g04034(.A1(new_n3916_), .A2(new_n4104_), .B(new_n4103_), .ZN(new_n4105_));
  NOR2_X1    g04035(.A1(new_n4100_), .A2(new_n4105_), .ZN(new_n4106_));
  NAND2_X1   g04036(.A1(new_n3889_), .A2(new_n3911_), .ZN(new_n4107_));
  XNOR2_X1   g04037(.A1(new_n4107_), .A2(new_n799_), .ZN(new_n4108_));
  NOR2_X1    g04038(.A1(new_n4108_), .A2(new_n3913_), .ZN(new_n4109_));
  NAND2_X1   g04039(.A1(new_n4108_), .A2(new_n3913_), .ZN(new_n4110_));
  INV_X1     g04040(.I(new_n4110_), .ZN(new_n4111_));
  NOR2_X1    g04041(.A1(new_n4111_), .A2(new_n4109_), .ZN(new_n4112_));
  INV_X1     g04042(.I(new_n4112_), .ZN(new_n4113_));
  INV_X1     g04043(.I(new_n3909_), .ZN(new_n4114_));
  NAND2_X1   g04044(.A1(new_n4114_), .A2(new_n3891_), .ZN(new_n4115_));
  XOR2_X1    g04045(.A1(new_n3909_), .A2(new_n3891_), .Z(new_n4116_));
  INV_X1     g04046(.I(new_n4116_), .ZN(new_n4117_));
  NAND2_X1   g04047(.A1(new_n4117_), .A2(new_n3906_), .ZN(new_n4118_));
  XNOR2_X1   g04048(.A1(new_n4118_), .A2(new_n4115_), .ZN(new_n4119_));
  NOR2_X1    g04049(.A1(new_n3889_), .A2(new_n4119_), .ZN(new_n4120_));
  NAND2_X1   g04050(.A1(new_n3889_), .A2(new_n4119_), .ZN(new_n4121_));
  INV_X1     g04051(.I(new_n4121_), .ZN(new_n4122_));
  NOR2_X1    g04052(.A1(new_n4122_), .A2(new_n4120_), .ZN(new_n4123_));
  INV_X1     g04053(.I(new_n4123_), .ZN(new_n4124_));
  NOR2_X1    g04054(.A1(new_n1104_), .A2(new_n1074_), .ZN(new_n4125_));
  NAND2_X1   g04055(.A1(new_n3865_), .A2(new_n3884_), .ZN(new_n4126_));
  XOR2_X1    g04056(.A1(new_n4126_), .A2(new_n4125_), .Z(new_n4127_));
  NOR2_X1    g04057(.A1(new_n4127_), .A2(new_n3886_), .ZN(new_n4128_));
  XNOR2_X1   g04058(.A1(new_n4126_), .A2(new_n4125_), .ZN(new_n4129_));
  NOR2_X1    g04059(.A1(new_n4129_), .A2(new_n3885_), .ZN(new_n4130_));
  NOR2_X1    g04060(.A1(new_n4130_), .A2(new_n4128_), .ZN(new_n4131_));
  XOR2_X1    g04061(.A1(new_n3855_), .A2(new_n3860_), .Z(new_n4132_));
  AOI21_X1   g04062(.A1(new_n3830_), .A2(new_n3831_), .B(new_n4132_), .ZN(new_n4133_));
  AOI21_X1   g04063(.A1(new_n3861_), .A2(new_n3864_), .B(new_n3832_), .ZN(new_n4134_));
  NOR2_X1    g04064(.A1(new_n4134_), .A2(new_n4133_), .ZN(new_n4135_));
  INV_X1     g04065(.I(new_n4135_), .ZN(new_n4136_));
  XOR2_X1    g04066(.A1(new_n3824_), .A2(new_n3828_), .Z(new_n4137_));
  AOI21_X1   g04067(.A1(new_n3796_), .A2(new_n3797_), .B(new_n4137_), .ZN(new_n4138_));
  NAND2_X1   g04068(.A1(new_n3829_), .A2(new_n3831_), .ZN(new_n4139_));
  NAND3_X1   g04069(.A1(new_n3796_), .A2(new_n3797_), .A3(new_n4139_), .ZN(new_n4140_));
  INV_X1     g04070(.I(new_n4140_), .ZN(new_n4141_));
  NOR2_X1    g04071(.A1(new_n4141_), .A2(new_n4138_), .ZN(new_n4142_));
  INV_X1     g04072(.I(new_n4142_), .ZN(new_n4143_));
  AOI21_X1   g04073(.A1(new_n3756_), .A2(new_n3703_), .B(new_n2951_), .ZN(new_n4144_));
  INV_X1     g04074(.I(new_n4144_), .ZN(new_n4145_));
  NAND3_X1   g04075(.A1(new_n3756_), .A2(new_n2951_), .A3(new_n3703_), .ZN(new_n4146_));
  AOI21_X1   g04076(.A1(new_n4145_), .A2(new_n4146_), .B(new_n3759_), .ZN(new_n4147_));
  INV_X1     g04077(.I(new_n4146_), .ZN(new_n4148_));
  NOR3_X1    g04078(.A1(new_n4148_), .A2(new_n3758_), .A3(new_n4144_), .ZN(new_n4149_));
  NOR2_X1    g04079(.A1(new_n4147_), .A2(new_n4149_), .ZN(new_n4150_));
  INV_X1     g04080(.I(new_n3703_), .ZN(new_n4151_));
  OAI21_X1   g04081(.A1(new_n3753_), .A2(new_n3752_), .B(new_n3725_), .ZN(new_n4152_));
  NAND2_X1   g04082(.A1(new_n3393_), .A2(new_n3342_), .ZN(new_n4153_));
  NAND2_X1   g04083(.A1(new_n4153_), .A2(new_n2954_), .ZN(new_n4154_));
  OAI21_X1   g04084(.A1(new_n4153_), .A2(new_n2954_), .B(\a[5] ), .ZN(new_n4155_));
  NAND3_X1   g04085(.A1(new_n3725_), .A2(new_n4155_), .A3(new_n4154_), .ZN(new_n4156_));
  AOI21_X1   g04086(.A1(new_n3722_), .A2(new_n3723_), .B(\a[2] ), .ZN(new_n4157_));
  NOR3_X1    g04087(.A1(new_n3717_), .A2(new_n3720_), .A3(new_n451_), .ZN(new_n4158_));
  NOR2_X1    g04088(.A1(new_n4158_), .A2(new_n4157_), .ZN(new_n4159_));
  OAI21_X1   g04089(.A1(new_n3752_), .A2(new_n3753_), .B(new_n4159_), .ZN(new_n4160_));
  NAND2_X1   g04090(.A1(new_n4160_), .A2(new_n4156_), .ZN(new_n4161_));
  NAND3_X1   g04091(.A1(new_n4161_), .A2(new_n3749_), .A3(new_n4152_), .ZN(new_n4162_));
  INV_X1     g04092(.I(new_n4152_), .ZN(new_n4163_));
  NOR3_X1    g04093(.A1(new_n4159_), .A2(new_n3753_), .A3(new_n3752_), .ZN(new_n4164_));
  NOR2_X1    g04094(.A1(new_n3754_), .A2(new_n3725_), .ZN(new_n4165_));
  OAI21_X1   g04095(.A1(new_n4165_), .A2(new_n4164_), .B(new_n3749_), .ZN(new_n4166_));
  NAND2_X1   g04096(.A1(new_n4166_), .A2(new_n4163_), .ZN(new_n4167_));
  NAND2_X1   g04097(.A1(new_n4167_), .A2(new_n4162_), .ZN(new_n4168_));
  NAND2_X1   g04098(.A1(new_n4168_), .A2(new_n4151_), .ZN(new_n4169_));
  NAND3_X1   g04099(.A1(new_n4167_), .A2(new_n4162_), .A3(new_n3703_), .ZN(new_n4170_));
  NAND2_X1   g04100(.A1(new_n4169_), .A2(new_n4170_), .ZN(new_n4171_));
  AOI22_X1   g04101(.A1(new_n3702_), .A2(new_n3698_), .B1(new_n4156_), .B2(new_n4160_), .ZN(new_n4172_));
  XOR2_X1    g04102(.A1(new_n3754_), .A2(new_n4159_), .Z(new_n4173_));
  NOR2_X1    g04103(.A1(new_n3703_), .A2(new_n4173_), .ZN(new_n4174_));
  NOR2_X1    g04104(.A1(new_n4174_), .A2(new_n4172_), .ZN(new_n4175_));
  INV_X1     g04105(.I(new_n3700_), .ZN(new_n4176_));
  OAI21_X1   g04106(.A1(new_n3555_), .A2(new_n3559_), .B(new_n3553_), .ZN(new_n4177_));
  AOI21_X1   g04107(.A1(new_n4177_), .A2(new_n3569_), .B(new_n3571_), .ZN(new_n4178_));
  OAI21_X1   g04108(.A1(new_n4178_), .A2(new_n3577_), .B(new_n3579_), .ZN(new_n4179_));
  NAND3_X1   g04109(.A1(new_n4179_), .A2(new_n3412_), .A3(new_n3585_), .ZN(new_n4180_));
  OAI21_X1   g04110(.A1(new_n3588_), .A2(new_n3592_), .B(new_n4180_), .ZN(new_n4181_));
  NAND3_X1   g04111(.A1(new_n4181_), .A2(new_n3412_), .A3(new_n3596_), .ZN(new_n4182_));
  OAI21_X1   g04112(.A1(new_n3599_), .A2(new_n3601_), .B(new_n4182_), .ZN(new_n4183_));
  AOI21_X1   g04113(.A1(new_n4183_), .A2(new_n3608_), .B(new_n3610_), .ZN(new_n4184_));
  OAI21_X1   g04114(.A1(new_n4184_), .A2(new_n3615_), .B(new_n3617_), .ZN(new_n4185_));
  OAI21_X1   g04115(.A1(new_n3631_), .A2(new_n3634_), .B(new_n3628_), .ZN(new_n4186_));
  NAND2_X1   g04116(.A1(new_n4186_), .A2(new_n3412_), .ZN(new_n4187_));
  NAND4_X1   g04117(.A1(new_n4185_), .A2(new_n4187_), .A3(new_n3407_), .A4(new_n3648_), .ZN(new_n4188_));
  AOI21_X1   g04118(.A1(new_n3412_), .A2(new_n4186_), .B(new_n3635_), .ZN(new_n4189_));
  AOI21_X1   g04119(.A1(new_n4189_), .A2(new_n4185_), .B(new_n3407_), .ZN(new_n4190_));
  INV_X1     g04120(.I(new_n3654_), .ZN(new_n4191_));
  OAI21_X1   g04121(.A1(new_n4190_), .A2(new_n4191_), .B(new_n4188_), .ZN(new_n4192_));
  NAND3_X1   g04122(.A1(new_n4192_), .A2(new_n3694_), .A3(new_n3695_), .ZN(new_n4193_));
  NAND3_X1   g04123(.A1(new_n3403_), .A2(new_n3413_), .A3(new_n4193_), .ZN(new_n4194_));
  AOI21_X1   g04124(.A1(new_n3400_), .A2(new_n3401_), .B(\a[5] ), .ZN(new_n4195_));
  NOR3_X1    g04125(.A1(new_n3394_), .A2(new_n3398_), .A3(new_n452_), .ZN(new_n4196_));
  OAI21_X1   g04126(.A1(new_n4195_), .A2(new_n4196_), .B(new_n3413_), .ZN(new_n4197_));
  NAND2_X1   g04127(.A1(new_n4197_), .A2(new_n3697_), .ZN(new_n4198_));
  AOI21_X1   g04128(.A1(new_n4198_), .A2(new_n4194_), .B(new_n4176_), .ZN(new_n4199_));
  NOR2_X1    g04129(.A1(new_n4197_), .A2(new_n3697_), .ZN(new_n4200_));
  AOI21_X1   g04130(.A1(new_n3403_), .A2(new_n3413_), .B(new_n4193_), .ZN(new_n4201_));
  NOR3_X1    g04131(.A1(new_n4200_), .A2(new_n4201_), .A3(new_n3700_), .ZN(new_n4202_));
  NOR2_X1    g04132(.A1(new_n4202_), .A2(new_n4199_), .ZN(new_n4203_));
  OAI21_X1   g04133(.A1(new_n3660_), .A2(new_n3663_), .B(new_n3412_), .ZN(new_n4204_));
  INV_X1     g04134(.I(new_n4204_), .ZN(new_n4205_));
  OAI21_X1   g04135(.A1(new_n3661_), .A2(new_n3662_), .B(new_n3332_), .ZN(new_n4206_));
  NAND3_X1   g04136(.A1(new_n3659_), .A2(new_n3657_), .A3(new_n3379_), .ZN(new_n4207_));
  AOI21_X1   g04137(.A1(new_n4206_), .A2(new_n4207_), .B(new_n3412_), .ZN(new_n4208_));
  NOR3_X1    g04138(.A1(new_n3660_), .A2(new_n3663_), .A3(new_n3413_), .ZN(new_n4209_));
  NOR2_X1    g04139(.A1(new_n4209_), .A2(new_n4208_), .ZN(new_n4210_));
  NOR3_X1    g04140(.A1(new_n4210_), .A2(new_n3693_), .A3(new_n4205_), .ZN(new_n4211_));
  NOR2_X1    g04141(.A1(new_n3664_), .A2(new_n3413_), .ZN(new_n4212_));
  OAI21_X1   g04142(.A1(new_n4211_), .A2(new_n4212_), .B(new_n3655_), .ZN(new_n4213_));
  OR2_X2     g04143(.A1(new_n3677_), .A2(new_n3692_), .Z(new_n4214_));
  OAI21_X1   g04144(.A1(new_n3660_), .A2(new_n3663_), .B(new_n3413_), .ZN(new_n4215_));
  NAND3_X1   g04145(.A1(new_n4206_), .A2(new_n4207_), .A3(new_n3412_), .ZN(new_n4216_));
  NAND2_X1   g04146(.A1(new_n4215_), .A2(new_n4216_), .ZN(new_n4217_));
  NAND3_X1   g04147(.A1(new_n4217_), .A2(new_n4214_), .A3(new_n4204_), .ZN(new_n4218_));
  INV_X1     g04148(.I(new_n4212_), .ZN(new_n4219_));
  NAND3_X1   g04149(.A1(new_n4218_), .A2(new_n4192_), .A3(new_n4219_), .ZN(new_n4220_));
  NAND2_X1   g04150(.A1(new_n4213_), .A2(new_n4220_), .ZN(new_n4221_));
  NOR2_X1    g04151(.A1(new_n3631_), .A2(new_n3634_), .ZN(new_n4222_));
  NOR2_X1    g04152(.A1(new_n3638_), .A2(new_n3412_), .ZN(new_n4223_));
  XOR2_X1    g04153(.A1(new_n3628_), .A2(new_n3412_), .Z(new_n4224_));
  NOR3_X1    g04154(.A1(new_n4224_), .A2(new_n4222_), .A3(new_n4223_), .ZN(new_n4225_));
  NOR2_X1    g04155(.A1(new_n3638_), .A2(new_n3412_), .ZN(new_n4226_));
  OAI21_X1   g04156(.A1(new_n4225_), .A2(new_n4226_), .B(new_n3619_), .ZN(new_n4227_));
  INV_X1     g04157(.I(new_n4227_), .ZN(new_n4228_));
  NOR3_X1    g04158(.A1(new_n4225_), .A2(new_n3619_), .A3(new_n4226_), .ZN(new_n4229_));
  NOR2_X1    g04159(.A1(new_n4228_), .A2(new_n4229_), .ZN(new_n4230_));
  NAND2_X1   g04160(.A1(new_n3664_), .A2(new_n3413_), .ZN(new_n4231_));
  NAND2_X1   g04161(.A1(new_n4231_), .A2(new_n4204_), .ZN(new_n4232_));
  NOR2_X1    g04162(.A1(new_n4192_), .A2(new_n4210_), .ZN(new_n4233_));
  AOI21_X1   g04163(.A1(new_n4192_), .A2(new_n4232_), .B(new_n4233_), .ZN(new_n4234_));
  AOI21_X1   g04164(.A1(new_n3405_), .A2(new_n3406_), .B(new_n3653_), .ZN(new_n4235_));
  INV_X1     g04165(.I(new_n4235_), .ZN(new_n4236_));
  AOI21_X1   g04166(.A1(new_n4189_), .A2(new_n4185_), .B(new_n4236_), .ZN(new_n4237_));
  NOR3_X1    g04167(.A1(new_n3649_), .A2(new_n3619_), .A3(new_n4235_), .ZN(new_n4238_));
  OAI21_X1   g04168(.A1(new_n4238_), .A2(new_n4237_), .B(new_n3652_), .ZN(new_n4239_));
  INV_X1     g04169(.I(new_n3652_), .ZN(new_n4240_));
  OAI21_X1   g04170(.A1(new_n3649_), .A2(new_n3619_), .B(new_n4235_), .ZN(new_n4241_));
  NAND3_X1   g04171(.A1(new_n4189_), .A2(new_n4185_), .A3(new_n4236_), .ZN(new_n4242_));
  NAND3_X1   g04172(.A1(new_n4241_), .A2(new_n4242_), .A3(new_n4240_), .ZN(new_n4243_));
  AND2_X2    g04173(.A1(new_n4239_), .A2(new_n4243_), .Z(new_n4244_));
  NOR3_X1    g04174(.A1(new_n4221_), .A2(new_n4234_), .A3(new_n4230_), .ZN(new_n4245_));
  INV_X1     g04175(.I(new_n4245_), .ZN(new_n4246_));
  AOI21_X1   g04176(.A1(new_n4218_), .A2(new_n4219_), .B(new_n4192_), .ZN(new_n4247_));
  NOR3_X1    g04177(.A1(new_n4211_), .A2(new_n3655_), .A3(new_n4212_), .ZN(new_n4248_));
  NOR2_X1    g04178(.A1(new_n4248_), .A2(new_n4247_), .ZN(new_n4249_));
  INV_X1     g04179(.I(new_n4229_), .ZN(new_n4250_));
  NAND2_X1   g04180(.A1(new_n4250_), .A2(new_n4227_), .ZN(new_n4251_));
  NAND2_X1   g04181(.A1(new_n4239_), .A2(new_n4243_), .ZN(new_n4252_));
  NAND3_X1   g04182(.A1(new_n4221_), .A2(new_n4230_), .A3(new_n4252_), .ZN(new_n4253_));
  OAI21_X1   g04183(.A1(new_n4249_), .A2(new_n4244_), .B(new_n4251_), .ZN(new_n4254_));
  AOI21_X1   g04184(.A1(new_n4254_), .A2(new_n4253_), .B(new_n4234_), .ZN(new_n4255_));
  NOR3_X1    g04185(.A1(new_n4255_), .A2(new_n4249_), .A3(new_n4251_), .ZN(new_n4256_));
  NOR4_X1    g04186(.A1(new_n4171_), .A2(new_n4175_), .A3(new_n4203_), .A4(new_n4246_), .ZN(new_n4257_));
  OR2_X2     g04187(.A1(new_n4174_), .A2(new_n4172_), .Z(new_n4258_));
  NAND2_X1   g04188(.A1(new_n4192_), .A2(new_n4232_), .ZN(new_n4259_));
  OAI21_X1   g04189(.A1(new_n4192_), .A2(new_n4210_), .B(new_n4259_), .ZN(new_n4260_));
  NOR3_X1    g04190(.A1(new_n4249_), .A2(new_n4251_), .A3(new_n4244_), .ZN(new_n4261_));
  AOI21_X1   g04191(.A1(new_n4221_), .A2(new_n4252_), .B(new_n4230_), .ZN(new_n4262_));
  OAI21_X1   g04192(.A1(new_n4261_), .A2(new_n4262_), .B(new_n4260_), .ZN(new_n4263_));
  NAND4_X1   g04193(.A1(new_n4263_), .A2(new_n4203_), .A3(new_n4221_), .A4(new_n4230_), .ZN(new_n4264_));
  NOR2_X1    g04194(.A1(new_n4264_), .A2(new_n4258_), .ZN(new_n4265_));
  NOR3_X1    g04195(.A1(new_n4175_), .A2(new_n4203_), .A3(new_n4246_), .ZN(new_n4266_));
  INV_X1     g04196(.I(new_n4266_), .ZN(new_n4267_));
  NAND3_X1   g04197(.A1(new_n4267_), .A2(new_n4265_), .A3(new_n4171_), .ZN(new_n4268_));
  AOI21_X1   g04198(.A1(new_n4268_), .A2(new_n4150_), .B(new_n4257_), .ZN(new_n4269_));
  XOR2_X1    g04199(.A1(new_n3792_), .A2(new_n3794_), .Z(new_n4270_));
  AND2_X2    g04200(.A1(new_n3762_), .A2(new_n4270_), .Z(new_n4271_));
  AOI21_X1   g04201(.A1(new_n3795_), .A2(new_n3797_), .B(new_n3762_), .ZN(new_n4272_));
  NOR2_X1    g04202(.A1(new_n4271_), .A2(new_n4272_), .ZN(new_n4273_));
  INV_X1     g04203(.I(new_n4273_), .ZN(new_n4274_));
  NAND2_X1   g04204(.A1(new_n4269_), .A2(new_n4150_), .ZN(new_n4275_));
  NOR2_X1    g04205(.A1(new_n4275_), .A2(new_n4274_), .ZN(new_n4276_));
  NOR2_X1    g04206(.A1(new_n4273_), .A2(new_n4150_), .ZN(new_n4277_));
  INV_X1     g04207(.I(new_n4277_), .ZN(new_n4278_));
  OAI22_X1   g04208(.A1(new_n4276_), .A2(new_n4142_), .B1(new_n4269_), .B2(new_n4278_), .ZN(new_n4279_));
  INV_X1     g04209(.I(new_n4279_), .ZN(new_n4280_));
  AOI21_X1   g04210(.A1(new_n4280_), .A2(new_n4143_), .B(new_n4136_), .ZN(new_n4281_));
  XNOR2_X1   g04211(.A1(new_n3881_), .A2(new_n3866_), .ZN(new_n4282_));
  XNOR2_X1   g04212(.A1(new_n3881_), .A2(new_n3866_), .ZN(new_n4283_));
  NOR2_X1    g04213(.A1(new_n3865_), .A2(new_n4283_), .ZN(new_n4284_));
  AOI21_X1   g04214(.A1(new_n3865_), .A2(new_n4282_), .B(new_n4284_), .ZN(new_n4285_));
  NAND2_X1   g04215(.A1(new_n4279_), .A2(new_n4142_), .ZN(new_n4286_));
  NOR2_X1    g04216(.A1(new_n4279_), .A2(new_n4142_), .ZN(new_n4287_));
  NAND2_X1   g04217(.A1(new_n4286_), .A2(new_n4136_), .ZN(new_n4288_));
  AOI21_X1   g04218(.A1(new_n4285_), .A2(new_n4288_), .B(new_n4281_), .ZN(new_n4289_));
  INV_X1     g04219(.I(new_n4285_), .ZN(new_n4290_));
  NAND2_X1   g04220(.A1(new_n3882_), .A2(new_n3866_), .ZN(new_n4291_));
  NAND2_X1   g04221(.A1(new_n4282_), .A2(new_n3878_), .ZN(new_n4292_));
  XNOR2_X1   g04222(.A1(new_n4292_), .A2(new_n4291_), .ZN(new_n4293_));
  NOR2_X1    g04223(.A1(new_n3865_), .A2(new_n4293_), .ZN(new_n4294_));
  AND2_X2    g04224(.A1(new_n3865_), .A2(new_n4293_), .Z(new_n4295_));
  NOR2_X1    g04225(.A1(new_n4295_), .A2(new_n4294_), .ZN(new_n4296_));
  INV_X1     g04226(.I(new_n4296_), .ZN(new_n4297_));
  NOR2_X1    g04227(.A1(new_n4297_), .A2(new_n4290_), .ZN(new_n4298_));
  AOI21_X1   g04228(.A1(new_n4289_), .A2(new_n4298_), .B(new_n4131_), .ZN(new_n4299_));
  INV_X1     g04229(.I(new_n4289_), .ZN(new_n4300_));
  NOR2_X1    g04230(.A1(new_n4296_), .A2(new_n4285_), .ZN(new_n4301_));
  NAND2_X1   g04231(.A1(new_n4300_), .A2(new_n4301_), .ZN(new_n4302_));
  INV_X1     g04232(.I(new_n4302_), .ZN(new_n4303_));
  NOR2_X1    g04233(.A1(new_n4303_), .A2(new_n4299_), .ZN(new_n4304_));
  INV_X1     g04234(.I(new_n4304_), .ZN(new_n4305_));
  AND2_X2    g04235(.A1(new_n3889_), .A2(new_n4117_), .Z(new_n4306_));
  XNOR2_X1   g04236(.A1(new_n3909_), .A2(new_n3891_), .ZN(new_n4307_));
  NOR2_X1    g04237(.A1(new_n3889_), .A2(new_n4307_), .ZN(new_n4308_));
  NOR2_X1    g04238(.A1(new_n4306_), .A2(new_n4308_), .ZN(new_n4309_));
  NAND3_X1   g04239(.A1(new_n4304_), .A2(new_n4309_), .A3(new_n4131_), .ZN(new_n4310_));
  NOR2_X1    g04240(.A1(new_n4131_), .A2(new_n4309_), .ZN(new_n4311_));
  AOI22_X1   g04241(.A1(new_n4310_), .A2(new_n4124_), .B1(new_n4305_), .B2(new_n4311_), .ZN(new_n4312_));
  AOI21_X1   g04242(.A1(new_n4312_), .A2(new_n4124_), .B(new_n4113_), .ZN(new_n4313_));
  INV_X1     g04243(.I(new_n4313_), .ZN(new_n4314_));
  INV_X1     g04244(.I(new_n4105_), .ZN(new_n4315_));
  NOR2_X1    g04245(.A1(new_n4312_), .A2(new_n4124_), .ZN(new_n4316_));
  INV_X1     g04246(.I(new_n4312_), .ZN(new_n4317_));
  NOR2_X1    g04247(.A1(new_n4317_), .A2(new_n4123_), .ZN(new_n4318_));
  OAI21_X1   g04248(.A1(new_n4316_), .A2(new_n4112_), .B(new_n4315_), .ZN(new_n4319_));
  NOR2_X1    g04249(.A1(new_n4315_), .A2(new_n4099_), .ZN(new_n4320_));
  AOI21_X1   g04250(.A1(new_n4319_), .A2(new_n4314_), .B(new_n4320_), .ZN(new_n4321_));
  NOR2_X1    g04251(.A1(new_n4321_), .A2(new_n4106_), .ZN(new_n4322_));
  NOR2_X1    g04252(.A1(new_n4090_), .A2(new_n4099_), .ZN(new_n4323_));
  OAI21_X1   g04253(.A1(new_n4322_), .A2(new_n4323_), .B(new_n4102_), .ZN(new_n4324_));
  INV_X1     g04254(.I(new_n4324_), .ZN(new_n4325_));
  NAND2_X1   g04255(.A1(new_n3941_), .A2(new_n4075_), .ZN(new_n4326_));
  XNOR2_X1   g04256(.A1(new_n3947_), .A2(new_n3943_), .ZN(new_n4327_));
  OAI21_X1   g04257(.A1(new_n3941_), .A2(new_n4327_), .B(new_n4326_), .ZN(new_n4328_));
  NOR2_X1    g04258(.A1(new_n4091_), .A2(new_n4328_), .ZN(new_n4329_));
  AOI21_X1   g04259(.A1(new_n4325_), .A2(new_n4329_), .B(new_n4081_), .ZN(new_n4330_));
  INV_X1     g04260(.I(new_n4328_), .ZN(new_n4331_));
  NOR2_X1    g04261(.A1(new_n4090_), .A2(new_n4331_), .ZN(new_n4332_));
  INV_X1     g04262(.I(new_n4332_), .ZN(new_n4333_));
  NOR2_X1    g04263(.A1(new_n4325_), .A2(new_n4333_), .ZN(new_n4334_));
  NOR2_X1    g04264(.A1(new_n4330_), .A2(new_n4334_), .ZN(new_n4335_));
  NOR2_X1    g04265(.A1(new_n4070_), .A2(new_n4081_), .ZN(new_n4336_));
  OAI21_X1   g04266(.A1(new_n4335_), .A2(new_n4336_), .B(new_n4084_), .ZN(new_n4337_));
  INV_X1     g04267(.I(new_n4337_), .ZN(new_n4338_));
  NOR2_X1    g04268(.A1(new_n4070_), .A2(new_n4060_), .ZN(new_n4339_));
  NOR2_X1    g04269(.A1(new_n4338_), .A2(new_n4339_), .ZN(new_n4340_));
  NOR2_X1    g04270(.A1(new_n4340_), .A2(new_n4072_), .ZN(new_n4341_));
  NOR2_X1    g04271(.A1(new_n4060_), .A2(new_n4053_), .ZN(new_n4342_));
  NOR2_X1    g04272(.A1(new_n4341_), .A2(new_n4342_), .ZN(new_n4343_));
  NOR2_X1    g04273(.A1(new_n4343_), .A2(new_n4062_), .ZN(new_n4344_));
  INV_X1     g04274(.I(new_n4344_), .ZN(new_n4345_));
  NOR2_X1    g04275(.A1(new_n4042_), .A2(new_n4053_), .ZN(new_n4346_));
  INV_X1     g04276(.I(new_n4346_), .ZN(new_n4347_));
  AOI21_X1   g04277(.A1(new_n4345_), .A2(new_n4347_), .B(new_n4055_), .ZN(new_n4348_));
  NOR2_X1    g04278(.A1(new_n4042_), .A2(new_n4035_), .ZN(new_n4349_));
  NOR2_X1    g04279(.A1(new_n4348_), .A2(new_n4349_), .ZN(new_n4350_));
  NOR2_X1    g04280(.A1(new_n4350_), .A2(new_n4044_), .ZN(new_n4351_));
  NOR2_X1    g04281(.A1(new_n4028_), .A2(new_n4035_), .ZN(new_n4352_));
  NOR2_X1    g04282(.A1(new_n4351_), .A2(new_n4352_), .ZN(new_n4353_));
  NOR2_X1    g04283(.A1(new_n4353_), .A2(new_n4037_), .ZN(new_n4354_));
  NOR2_X1    g04284(.A1(new_n4017_), .A2(new_n4028_), .ZN(new_n4355_));
  OAI21_X1   g04285(.A1(new_n4354_), .A2(new_n4355_), .B(new_n4031_), .ZN(new_n4356_));
  OR4_X2     g04286(.A1(new_n162_), .A2(new_n179_), .A3(new_n167_), .A4(new_n183_), .Z(new_n4357_));
  NAND4_X1   g04287(.A1(new_n4003_), .A2(new_n166_), .A3(new_n4011_), .A4(new_n4357_), .ZN(new_n4358_));
  NOR2_X1    g04288(.A1(new_n174_), .A2(new_n80_), .ZN(new_n4359_));
  NOR2_X1    g04289(.A1(new_n4359_), .A2(new_n175_), .ZN(new_n4360_));
  XOR2_X1    g04290(.A1(new_n4360_), .A2(new_n93_), .Z(new_n4361_));
  XOR2_X1    g04291(.A1(new_n4361_), .A2(new_n102_), .Z(new_n4362_));
  XOR2_X1    g04292(.A1(new_n4362_), .A2(\a[26] ), .Z(new_n4363_));
  NAND2_X1   g04293(.A1(new_n182_), .A2(new_n71_), .ZN(new_n4364_));
  NAND2_X1   g04294(.A1(new_n4364_), .A2(new_n181_), .ZN(new_n4365_));
  INV_X1     g04295(.I(new_n4365_), .ZN(new_n4366_));
  NOR2_X1    g04296(.A1(new_n4363_), .A2(new_n4366_), .ZN(new_n4367_));
  INV_X1     g04297(.I(new_n4367_), .ZN(new_n4368_));
  NAND2_X1   g04298(.A1(new_n4363_), .A2(new_n4366_), .ZN(new_n4369_));
  AOI22_X1   g04299(.A1(new_n4358_), .A2(new_n184_), .B1(new_n4368_), .B2(new_n4369_), .ZN(new_n4370_));
  NAND2_X1   g04300(.A1(new_n4358_), .A2(new_n184_), .ZN(new_n4371_));
  XOR2_X1    g04301(.A1(new_n4363_), .A2(new_n4365_), .Z(new_n4372_));
  NOR2_X1    g04302(.A1(new_n4371_), .A2(new_n4372_), .ZN(new_n4373_));
  NOR2_X1    g04303(.A1(new_n4373_), .A2(new_n4370_), .ZN(new_n4374_));
  INV_X1     g04304(.I(new_n4374_), .ZN(new_n4375_));
  XOR2_X1    g04305(.A1(new_n4017_), .A2(new_n4375_), .Z(new_n4376_));
  INV_X1     g04306(.I(new_n4376_), .ZN(new_n4377_));
  XOR2_X1    g04307(.A1(new_n93_), .A2(new_n65_), .Z(new_n4378_));
  AND2_X2    g04308(.A1(new_n4378_), .A2(new_n102_), .Z(new_n4379_));
  INV_X1     g04309(.I(new_n4379_), .ZN(new_n4380_));
  NOR2_X1    g04310(.A1(new_n4378_), .A2(new_n102_), .ZN(new_n4381_));
  INV_X1     g04311(.I(new_n4381_), .ZN(new_n4382_));
  AOI22_X1   g04312(.A1(new_n4360_), .A2(new_n94_), .B1(new_n4380_), .B2(new_n4382_), .ZN(new_n4383_));
  NOR4_X1    g04313(.A1(new_n149_), .A2(\a[26] ), .A3(new_n102_), .A4(new_n93_), .ZN(new_n4384_));
  NOR2_X1    g04314(.A1(new_n4383_), .A2(new_n4384_), .ZN(new_n4385_));
  NOR2_X1    g04315(.A1(new_n4361_), .A2(new_n80_), .ZN(new_n4386_));
  NAND2_X1   g04316(.A1(new_n4361_), .A2(new_n80_), .ZN(new_n4387_));
  AOI21_X1   g04317(.A1(\a[26] ), .A2(new_n4387_), .B(new_n4386_), .ZN(new_n4388_));
  AND2_X2    g04318(.A1(new_n4388_), .A2(new_n4385_), .Z(new_n4389_));
  NOR2_X1    g04319(.A1(new_n4388_), .A2(new_n4385_), .ZN(new_n4390_));
  NOR2_X1    g04320(.A1(new_n4389_), .A2(new_n4390_), .ZN(new_n4391_));
  NOR2_X1    g04321(.A1(new_n4372_), .A2(new_n4391_), .ZN(new_n4392_));
  XOR2_X1    g04322(.A1(new_n4392_), .A2(new_n4368_), .Z(new_n4393_));
  NOR2_X1    g04323(.A1(new_n4371_), .A2(new_n4393_), .ZN(new_n4394_));
  NAND2_X1   g04324(.A1(new_n4371_), .A2(new_n4393_), .ZN(new_n4395_));
  INV_X1     g04325(.I(new_n4395_), .ZN(new_n4396_));
  NOR2_X1    g04326(.A1(new_n4396_), .A2(new_n4394_), .ZN(new_n4397_));
  NOR2_X1    g04327(.A1(new_n4375_), .A2(new_n4397_), .ZN(new_n4398_));
  INV_X1     g04328(.I(new_n4397_), .ZN(new_n4399_));
  NOR2_X1    g04329(.A1(new_n4399_), .A2(new_n4374_), .ZN(new_n4400_));
  OAI21_X1   g04330(.A1(new_n4398_), .A2(new_n4400_), .B(new_n4377_), .ZN(new_n4401_));
  INV_X1     g04331(.I(new_n4401_), .ZN(new_n4402_));
  XOR2_X1    g04332(.A1(new_n4356_), .A2(new_n4402_), .Z(new_n4403_));
  NOR2_X1    g04333(.A1(new_n4374_), .A2(new_n88_), .ZN(new_n4404_));
  INV_X1     g04334(.I(new_n4404_), .ZN(new_n4405_));
  INV_X1     g04335(.I(new_n92_), .ZN(new_n4406_));
  AOI22_X1   g04336(.A1(new_n4018_), .A2(new_n4406_), .B1(new_n962_), .B2(new_n4399_), .ZN(new_n4407_));
  AOI21_X1   g04337(.A1(new_n4407_), .A2(new_n4405_), .B(new_n82_), .ZN(new_n4408_));
  NAND2_X1   g04338(.A1(new_n4403_), .A2(new_n4408_), .ZN(new_n4409_));
  INV_X1     g04339(.I(new_n1973_), .ZN(new_n4410_));
  XNOR2_X1   g04340(.A1(\a[20] ), .A2(\a[23] ), .ZN(new_n4411_));
  NOR3_X1    g04341(.A1(new_n188_), .A2(new_n1121_), .A3(new_n4411_), .ZN(new_n4412_));
  NOR3_X1    g04342(.A1(new_n4410_), .A2(new_n247_), .A3(new_n4412_), .ZN(new_n4413_));
  NOR2_X1    g04343(.A1(new_n4413_), .A2(new_n68_), .ZN(new_n4414_));
  INV_X1     g04344(.I(new_n4414_), .ZN(new_n4415_));
  NAND2_X1   g04345(.A1(new_n4413_), .A2(new_n68_), .ZN(new_n4416_));
  AND2_X2    g04346(.A1(new_n4415_), .A2(new_n4416_), .Z(new_n4417_));
  NAND2_X1   g04347(.A1(new_n4391_), .A2(new_n4363_), .ZN(new_n4418_));
  OAI21_X1   g04348(.A1(new_n4391_), .A2(new_n4363_), .B(new_n4366_), .ZN(new_n4419_));
  AND3_X2    g04349(.A1(new_n4371_), .A2(new_n4418_), .A3(new_n4419_), .Z(new_n4420_));
  NAND2_X1   g04350(.A1(new_n4360_), .A2(new_n94_), .ZN(new_n4421_));
  AOI21_X1   g04351(.A1(new_n4421_), .A2(new_n4380_), .B(new_n4381_), .ZN(new_n4422_));
  NOR2_X1    g04352(.A1(new_n94_), .A2(new_n65_), .ZN(new_n4423_));
  NOR2_X1    g04353(.A1(new_n4423_), .A2(new_n80_), .ZN(new_n4424_));
  INV_X1     g04354(.I(new_n4423_), .ZN(new_n4425_));
  NOR2_X1    g04355(.A1(new_n4425_), .A2(new_n102_), .ZN(new_n4426_));
  OR2_X2     g04356(.A1(new_n4426_), .A2(new_n4424_), .Z(new_n4427_));
  NAND2_X1   g04357(.A1(new_n4425_), .A2(new_n80_), .ZN(new_n4428_));
  NAND2_X1   g04358(.A1(new_n4423_), .A2(new_n102_), .ZN(new_n4429_));
  AOI21_X1   g04359(.A1(new_n4428_), .A2(new_n4429_), .B(new_n965_), .ZN(new_n4430_));
  AOI21_X1   g04360(.A1(new_n4427_), .A2(new_n965_), .B(new_n4430_), .ZN(new_n4431_));
  NOR2_X1    g04361(.A1(new_n4422_), .A2(new_n4431_), .ZN(new_n4432_));
  XNOR2_X1   g04362(.A1(new_n4420_), .A2(new_n4432_), .ZN(new_n4433_));
  NOR2_X1    g04363(.A1(new_n4433_), .A2(new_n4389_), .ZN(new_n4434_));
  NAND2_X1   g04364(.A1(new_n4433_), .A2(new_n4389_), .ZN(new_n4435_));
  INV_X1     g04365(.I(new_n4435_), .ZN(new_n4436_));
  NOR2_X1    g04366(.A1(new_n4436_), .A2(new_n4434_), .ZN(new_n4437_));
  INV_X1     g04367(.I(new_n4437_), .ZN(new_n4438_));
  NOR2_X1    g04368(.A1(new_n4438_), .A2(new_n4399_), .ZN(new_n4439_));
  INV_X1     g04369(.I(new_n4439_), .ZN(new_n4440_));
  INV_X1     g04370(.I(new_n4356_), .ZN(new_n4441_));
  NOR2_X1    g04371(.A1(new_n4018_), .A2(new_n4375_), .ZN(new_n4442_));
  AOI21_X1   g04372(.A1(new_n4441_), .A2(new_n4442_), .B(new_n4397_), .ZN(new_n4443_));
  NOR2_X1    g04373(.A1(new_n4017_), .A2(new_n4374_), .ZN(new_n4444_));
  INV_X1     g04374(.I(new_n4444_), .ZN(new_n4445_));
  NOR2_X1    g04375(.A1(new_n4441_), .A2(new_n4445_), .ZN(new_n4446_));
  NOR2_X1    g04376(.A1(new_n4437_), .A2(new_n4397_), .ZN(new_n4447_));
  INV_X1     g04377(.I(new_n4447_), .ZN(new_n4448_));
  OAI21_X1   g04378(.A1(new_n4443_), .A2(new_n4446_), .B(new_n4448_), .ZN(new_n4449_));
  NAND2_X1   g04379(.A1(new_n4449_), .A2(new_n4440_), .ZN(new_n4450_));
  INV_X1     g04380(.I(new_n4450_), .ZN(new_n4451_));
  INV_X1     g04381(.I(new_n4422_), .ZN(new_n4452_));
  NAND2_X1   g04382(.A1(new_n4389_), .A2(new_n4452_), .ZN(new_n4453_));
  NOR2_X1    g04383(.A1(new_n4389_), .A2(new_n4452_), .ZN(new_n4454_));
  NOR2_X1    g04384(.A1(new_n4454_), .A2(new_n4431_), .ZN(new_n4455_));
  NAND2_X1   g04385(.A1(new_n4420_), .A2(new_n4455_), .ZN(new_n4456_));
  NAND2_X1   g04386(.A1(new_n4456_), .A2(new_n4453_), .ZN(new_n4457_));
  NAND3_X1   g04387(.A1(new_n4406_), .A2(\a[31] ), .A3(new_n81_), .ZN(new_n4458_));
  XOR2_X1    g04388(.A1(new_n4458_), .A2(new_n72_), .Z(new_n4459_));
  INV_X1     g04389(.I(new_n4459_), .ZN(new_n4460_));
  NOR2_X1    g04390(.A1(new_n4424_), .A2(new_n512_), .ZN(new_n4461_));
  NOR2_X1    g04391(.A1(new_n4461_), .A2(new_n4426_), .ZN(new_n4462_));
  XOR2_X1    g04392(.A1(new_n4462_), .A2(new_n4460_), .Z(new_n4463_));
  INV_X1     g04393(.I(new_n4463_), .ZN(new_n4464_));
  NOR2_X1    g04394(.A1(new_n4457_), .A2(new_n4464_), .ZN(new_n4465_));
  INV_X1     g04395(.I(new_n4457_), .ZN(new_n4466_));
  NOR2_X1    g04396(.A1(new_n4466_), .A2(new_n4463_), .ZN(new_n4467_));
  NOR2_X1    g04397(.A1(new_n4467_), .A2(new_n4465_), .ZN(new_n4468_));
  INV_X1     g04398(.I(new_n4468_), .ZN(new_n4469_));
  NOR2_X1    g04399(.A1(new_n4438_), .A2(new_n4469_), .ZN(new_n4470_));
  INV_X1     g04400(.I(new_n4470_), .ZN(new_n4471_));
  NOR2_X1    g04401(.A1(new_n4437_), .A2(new_n4468_), .ZN(new_n4472_));
  INV_X1     g04402(.I(new_n4472_), .ZN(new_n4473_));
  AOI21_X1   g04403(.A1(new_n4471_), .A2(new_n4473_), .B(new_n4451_), .ZN(new_n4474_));
  XNOR2_X1   g04404(.A1(new_n4437_), .A2(new_n4468_), .ZN(new_n4475_));
  NOR2_X1    g04405(.A1(new_n4450_), .A2(new_n4475_), .ZN(new_n4476_));
  NOR2_X1    g04406(.A1(new_n4474_), .A2(new_n4476_), .ZN(new_n4477_));
  INV_X1     g04407(.I(new_n4477_), .ZN(new_n4478_));
  NAND2_X1   g04408(.A1(new_n4438_), .A2(new_n87_), .ZN(new_n4479_));
  AOI22_X1   g04409(.A1(new_n4469_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n4399_), .ZN(new_n4480_));
  AOI21_X1   g04410(.A1(new_n4479_), .A2(new_n4480_), .B(new_n82_), .ZN(new_n4481_));
  AOI21_X1   g04411(.A1(new_n4478_), .A2(new_n4481_), .B(new_n4417_), .ZN(new_n4482_));
  INV_X1     g04412(.I(new_n4417_), .ZN(new_n4483_));
  NAND2_X1   g04413(.A1(new_n4478_), .A2(new_n4481_), .ZN(new_n4484_));
  NOR2_X1    g04414(.A1(new_n4484_), .A2(new_n4483_), .ZN(new_n4485_));
  NOR2_X1    g04415(.A1(new_n4485_), .A2(new_n4482_), .ZN(new_n4486_));
  NOR2_X1    g04416(.A1(new_n4486_), .A2(new_n4409_), .ZN(new_n4487_));
  INV_X1     g04417(.I(new_n4409_), .ZN(new_n4488_));
  XOR2_X1    g04418(.A1(new_n4484_), .A2(new_n4417_), .Z(new_n4489_));
  NOR2_X1    g04419(.A1(new_n4489_), .A2(new_n4488_), .ZN(new_n4490_));
  NOR2_X1    g04420(.A1(new_n4490_), .A2(new_n4487_), .ZN(new_n4491_));
  INV_X1     g04421(.I(new_n4491_), .ZN(new_n4492_));
  AOI21_X1   g04422(.A1(new_n4450_), .A2(new_n4473_), .B(new_n4470_), .ZN(new_n4493_));
  INV_X1     g04423(.I(new_n4493_), .ZN(new_n4494_));
  NAND2_X1   g04424(.A1(new_n4462_), .A2(new_n4459_), .ZN(new_n4495_));
  NAND4_X1   g04425(.A1(new_n4406_), .A2(new_n72_), .A3(\a[31] ), .A4(new_n81_), .ZN(new_n4496_));
  AOI21_X1   g04426(.A1(new_n4495_), .A2(new_n4496_), .B(new_n4463_), .ZN(new_n4497_));
  INV_X1     g04427(.I(new_n4497_), .ZN(new_n4498_));
  NOR2_X1    g04428(.A1(new_n4457_), .A2(new_n4498_), .ZN(new_n4499_));
  NOR2_X1    g04429(.A1(new_n4466_), .A2(new_n4497_), .ZN(new_n4500_));
  NOR2_X1    g04430(.A1(new_n4500_), .A2(new_n4499_), .ZN(new_n4501_));
  XNOR2_X1   g04431(.A1(new_n4468_), .A2(new_n4501_), .ZN(new_n4502_));
  INV_X1     g04432(.I(new_n4502_), .ZN(new_n4503_));
  AOI21_X1   g04433(.A1(new_n94_), .A2(new_n512_), .B(new_n72_), .ZN(new_n4504_));
  AOI21_X1   g04434(.A1(new_n93_), .A2(new_n965_), .B(new_n4504_), .ZN(new_n4505_));
  NOR2_X1    g04435(.A1(new_n965_), .A2(new_n72_), .ZN(new_n4506_));
  NOR2_X1    g04436(.A1(new_n512_), .A2(\a[29] ), .ZN(new_n4507_));
  OAI21_X1   g04437(.A1(new_n4506_), .A2(new_n4507_), .B(new_n4505_), .ZN(new_n4508_));
  INV_X1     g04438(.I(new_n4508_), .ZN(new_n4509_));
  OAI21_X1   g04439(.A1(new_n4495_), .A2(new_n4496_), .B(new_n4463_), .ZN(new_n4510_));
  NAND2_X1   g04440(.A1(new_n4457_), .A2(new_n4510_), .ZN(new_n4511_));
  XOR2_X1    g04441(.A1(new_n4511_), .A2(new_n4506_), .Z(new_n4512_));
  NOR2_X1    g04442(.A1(new_n4512_), .A2(new_n4509_), .ZN(new_n4513_));
  NAND2_X1   g04443(.A1(new_n4512_), .A2(new_n4509_), .ZN(new_n4514_));
  INV_X1     g04444(.I(new_n4514_), .ZN(new_n4515_));
  NOR2_X1    g04445(.A1(new_n4515_), .A2(new_n4513_), .ZN(new_n4516_));
  NOR2_X1    g04446(.A1(new_n4516_), .A2(new_n4469_), .ZN(new_n4517_));
  INV_X1     g04447(.I(new_n4516_), .ZN(new_n4518_));
  NOR2_X1    g04448(.A1(new_n4518_), .A2(new_n4468_), .ZN(new_n4519_));
  OAI21_X1   g04449(.A1(new_n4519_), .A2(new_n4517_), .B(new_n4503_), .ZN(new_n4520_));
  NOR2_X1    g04450(.A1(new_n4494_), .A2(new_n4520_), .ZN(new_n4521_));
  INV_X1     g04451(.I(new_n4520_), .ZN(new_n4522_));
  NOR2_X1    g04452(.A1(new_n4493_), .A2(new_n4522_), .ZN(new_n4523_));
  NOR2_X1    g04453(.A1(new_n4521_), .A2(new_n4523_), .ZN(new_n4524_));
  XNOR2_X1   g04454(.A1(\a[26] ), .A2(\a[29] ), .ZN(new_n4525_));
  NOR3_X1    g04455(.A1(new_n941_), .A2(new_n918_), .A3(new_n4525_), .ZN(new_n4526_));
  INV_X1     g04456(.I(new_n4526_), .ZN(new_n4527_));
  NOR2_X1    g04457(.A1(new_n99_), .A2(\a[27] ), .ZN(new_n4528_));
  AOI21_X1   g04458(.A1(\a[27] ), .A2(new_n78_), .B(new_n4528_), .ZN(new_n4529_));
  NOR2_X1    g04459(.A1(new_n4527_), .A2(new_n4529_), .ZN(new_n4530_));
  NOR2_X1    g04460(.A1(new_n4468_), .A2(new_n4501_), .ZN(new_n4531_));
  OAI22_X1   g04461(.A1(new_n4516_), .A2(new_n79_), .B1(new_n4530_), .B2(new_n4531_), .ZN(new_n4532_));
  AOI21_X1   g04462(.A1(new_n4532_), .A2(new_n72_), .B(new_n79_), .ZN(new_n4533_));
  XOR2_X1    g04463(.A1(new_n4524_), .A2(new_n4533_), .Z(new_n4534_));
  INV_X1     g04464(.I(new_n4534_), .ZN(new_n4535_));
  NOR2_X1    g04465(.A1(new_n4443_), .A2(new_n4446_), .ZN(new_n4536_));
  XOR2_X1    g04466(.A1(new_n4437_), .A2(new_n4399_), .Z(new_n4537_));
  NOR2_X1    g04467(.A1(new_n4536_), .A2(new_n4537_), .ZN(new_n4538_));
  NOR2_X1    g04468(.A1(new_n4439_), .A2(new_n4447_), .ZN(new_n4539_));
  NOR3_X1    g04469(.A1(new_n4443_), .A2(new_n4446_), .A3(new_n4539_), .ZN(new_n4540_));
  NOR2_X1    g04470(.A1(new_n4538_), .A2(new_n4540_), .ZN(new_n4541_));
  INV_X1     g04471(.I(new_n4541_), .ZN(new_n4542_));
  NOR2_X1    g04472(.A1(new_n4437_), .A2(new_n511_), .ZN(new_n4543_));
  INV_X1     g04473(.I(new_n4543_), .ZN(new_n4544_));
  NOR2_X1    g04474(.A1(new_n88_), .A2(new_n92_), .ZN(new_n4545_));
  NOR2_X1    g04475(.A1(new_n4397_), .A2(new_n4374_), .ZN(new_n4546_));
  NOR2_X1    g04476(.A1(new_n4546_), .A2(new_n4545_), .ZN(new_n4547_));
  AOI21_X1   g04477(.A1(new_n4544_), .A2(new_n4547_), .B(new_n82_), .ZN(new_n4548_));
  NAND2_X1   g04478(.A1(new_n4542_), .A2(new_n4548_), .ZN(new_n4549_));
  INV_X1     g04479(.I(new_n4549_), .ZN(new_n4550_));
  NOR2_X1    g04480(.A1(new_n4535_), .A2(new_n4550_), .ZN(new_n4551_));
  NOR2_X1    g04481(.A1(new_n4551_), .A2(new_n4488_), .ZN(new_n4552_));
  NOR2_X1    g04482(.A1(new_n4534_), .A2(new_n4549_), .ZN(new_n4553_));
  NOR2_X1    g04483(.A1(new_n4552_), .A2(new_n4553_), .ZN(new_n4554_));
  INV_X1     g04484(.I(new_n4501_), .ZN(new_n4555_));
  NOR2_X1    g04485(.A1(new_n4469_), .A2(new_n4555_), .ZN(new_n4556_));
  AOI21_X1   g04486(.A1(new_n4493_), .A2(new_n4556_), .B(new_n4516_), .ZN(new_n4557_));
  NOR3_X1    g04487(.A1(new_n4493_), .A2(new_n4468_), .A3(new_n4501_), .ZN(new_n4558_));
  NOR2_X1    g04488(.A1(new_n4558_), .A2(new_n4557_), .ZN(new_n4559_));
  INV_X1     g04489(.I(new_n4506_), .ZN(new_n4560_));
  NOR2_X1    g04490(.A1(new_n4508_), .A2(new_n4560_), .ZN(new_n4561_));
  AOI21_X1   g04491(.A1(new_n4560_), .A2(new_n4508_), .B(new_n4511_), .ZN(new_n4562_));
  NOR2_X1    g04492(.A1(new_n4562_), .A2(new_n4561_), .ZN(new_n4563_));
  INV_X1     g04493(.I(new_n4563_), .ZN(new_n4564_));
  XOR2_X1    g04494(.A1(new_n4516_), .A2(new_n4564_), .Z(new_n4565_));
  NOR2_X1    g04495(.A1(new_n4518_), .A2(new_n4564_), .ZN(new_n4566_));
  NOR2_X1    g04496(.A1(new_n4516_), .A2(new_n4563_), .ZN(new_n4567_));
  OAI21_X1   g04497(.A1(new_n4566_), .A2(new_n4567_), .B(new_n4559_), .ZN(new_n4568_));
  OAI21_X1   g04498(.A1(new_n4559_), .A2(new_n4565_), .B(new_n4568_), .ZN(new_n4569_));
  INV_X1     g04499(.I(new_n4529_), .ZN(new_n4570_));
  AOI22_X1   g04500(.A1(new_n4518_), .A2(new_n4526_), .B1(new_n4555_), .B2(new_n4570_), .ZN(new_n4571_));
  AOI21_X1   g04501(.A1(new_n101_), .A2(new_n4564_), .B(new_n4571_), .ZN(new_n4572_));
  OAI21_X1   g04502(.A1(new_n4572_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n4573_));
  XOR2_X1    g04503(.A1(new_n4569_), .A2(new_n4573_), .Z(new_n4574_));
  NAND2_X1   g04504(.A1(new_n4554_), .A2(new_n4574_), .ZN(new_n4575_));
  NOR2_X1    g04505(.A1(new_n4554_), .A2(new_n4574_), .ZN(new_n4576_));
  AOI21_X1   g04506(.A1(new_n4492_), .A2(new_n4575_), .B(new_n4576_), .ZN(new_n4577_));
  INV_X1     g04507(.I(new_n4482_), .ZN(new_n4578_));
  AOI21_X1   g04508(.A1(new_n4578_), .A2(new_n4488_), .B(new_n4485_), .ZN(new_n4579_));
  INV_X1     g04509(.I(new_n4579_), .ZN(new_n4580_));
  NOR2_X1    g04510(.A1(new_n4493_), .A2(new_n4502_), .ZN(new_n4581_));
  OAI21_X1   g04511(.A1(new_n4531_), .A2(new_n4556_), .B(new_n4493_), .ZN(new_n4582_));
  INV_X1     g04512(.I(new_n4582_), .ZN(new_n4583_));
  NOR2_X1    g04513(.A1(new_n4583_), .A2(new_n4581_), .ZN(new_n4584_));
  INV_X1     g04514(.I(new_n4584_), .ZN(new_n4585_));
  NAND2_X1   g04515(.A1(new_n4469_), .A2(new_n87_), .ZN(new_n4586_));
  AOI22_X1   g04516(.A1(new_n4438_), .A2(new_n4406_), .B1(new_n962_), .B2(new_n4555_), .ZN(new_n4587_));
  AOI21_X1   g04517(.A1(new_n4587_), .A2(new_n4586_), .B(new_n82_), .ZN(new_n4588_));
  NAND2_X1   g04518(.A1(new_n4585_), .A2(new_n4588_), .ZN(new_n4589_));
  INV_X1     g04519(.I(new_n4589_), .ZN(new_n4590_));
  NOR3_X1    g04520(.A1(new_n4558_), .A2(new_n4557_), .A3(new_n4565_), .ZN(new_n4591_));
  INV_X1     g04521(.I(new_n4565_), .ZN(new_n4592_));
  NOR2_X1    g04522(.A1(new_n4559_), .A2(new_n4592_), .ZN(new_n4593_));
  NOR2_X1    g04523(.A1(new_n4593_), .A2(new_n4591_), .ZN(new_n4594_));
  AOI22_X1   g04524(.A1(new_n4518_), .A2(new_n4570_), .B1(new_n4526_), .B2(new_n4564_), .ZN(new_n4595_));
  NOR2_X1    g04525(.A1(new_n4564_), .A2(new_n79_), .ZN(new_n4596_));
  OAI21_X1   g04526(.A1(new_n4595_), .A2(new_n4596_), .B(new_n72_), .ZN(new_n4597_));
  NAND2_X1   g04527(.A1(new_n4597_), .A2(new_n101_), .ZN(new_n4598_));
  XNOR2_X1   g04528(.A1(new_n4594_), .A2(new_n4598_), .ZN(new_n4599_));
  XOR2_X1    g04529(.A1(new_n4599_), .A2(new_n4590_), .Z(new_n4600_));
  NAND2_X1   g04530(.A1(new_n4600_), .A2(new_n4580_), .ZN(new_n4601_));
  AND2_X2    g04531(.A1(new_n4599_), .A2(new_n4590_), .Z(new_n4602_));
  NOR2_X1    g04532(.A1(new_n4599_), .A2(new_n4590_), .ZN(new_n4603_));
  OAI21_X1   g04533(.A1(new_n4602_), .A2(new_n4603_), .B(new_n4579_), .ZN(new_n4604_));
  NAND2_X1   g04534(.A1(new_n4601_), .A2(new_n4604_), .ZN(new_n4605_));
  INV_X1     g04535(.I(new_n4605_), .ZN(new_n4606_));
  INV_X1     g04536(.I(new_n4559_), .ZN(new_n4607_));
  NAND2_X1   g04537(.A1(new_n4559_), .A2(new_n4566_), .ZN(new_n4608_));
  AOI22_X1   g04538(.A1(new_n4608_), .A2(new_n4563_), .B1(new_n4607_), .B2(new_n4567_), .ZN(new_n4609_));
  NOR2_X1    g04539(.A1(new_n4609_), .A2(new_n4564_), .ZN(new_n4610_));
  NOR2_X1    g04540(.A1(new_n115_), .A2(\a[24] ), .ZN(new_n4611_));
  AOI21_X1   g04541(.A1(\a[24] ), .A2(new_n69_), .B(new_n4611_), .ZN(new_n4612_));
  INV_X1     g04542(.I(new_n4612_), .ZN(new_n4613_));
  NOR3_X1    g04543(.A1(new_n4564_), .A2(new_n1128_), .A3(new_n4613_), .ZN(new_n4614_));
  OAI21_X1   g04544(.A1(new_n4614_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n4615_));
  XOR2_X1    g04545(.A1(new_n4610_), .A2(new_n4615_), .Z(new_n4616_));
  INV_X1     g04546(.I(new_n4616_), .ZN(new_n4617_));
  NOR2_X1    g04547(.A1(new_n4606_), .A2(new_n4617_), .ZN(new_n4618_));
  NOR2_X1    g04548(.A1(new_n4618_), .A2(new_n4577_), .ZN(new_n4619_));
  NOR2_X1    g04549(.A1(new_n4605_), .A2(new_n4616_), .ZN(new_n4620_));
  NOR2_X1    g04550(.A1(new_n4619_), .A2(new_n4620_), .ZN(new_n4621_));
  NOR2_X1    g04551(.A1(new_n4602_), .A2(new_n4579_), .ZN(new_n4622_));
  NOR2_X1    g04552(.A1(new_n4622_), .A2(new_n4603_), .ZN(new_n4623_));
  INV_X1     g04553(.I(new_n4524_), .ZN(new_n4624_));
  NAND2_X1   g04554(.A1(new_n4518_), .A2(new_n962_), .ZN(new_n4625_));
  NOR2_X1    g04555(.A1(new_n4531_), .A2(new_n4545_), .ZN(new_n4626_));
  AOI21_X1   g04556(.A1(new_n4625_), .A2(new_n4626_), .B(new_n82_), .ZN(new_n4627_));
  NAND2_X1   g04557(.A1(new_n4624_), .A2(new_n4627_), .ZN(new_n4628_));
  XOR2_X1    g04558(.A1(new_n4589_), .A2(new_n4628_), .Z(new_n4629_));
  NOR2_X1    g04559(.A1(new_n4623_), .A2(new_n4629_), .ZN(new_n4630_));
  INV_X1     g04560(.I(new_n4623_), .ZN(new_n4631_));
  NOR2_X1    g04561(.A1(new_n4590_), .A2(new_n4628_), .ZN(new_n4632_));
  INV_X1     g04562(.I(new_n4628_), .ZN(new_n4633_));
  NOR2_X1    g04563(.A1(new_n4633_), .A2(new_n4589_), .ZN(new_n4634_));
  NOR2_X1    g04564(.A1(new_n4632_), .A2(new_n4634_), .ZN(new_n4635_));
  NOR2_X1    g04565(.A1(new_n4631_), .A2(new_n4635_), .ZN(new_n4636_));
  NOR2_X1    g04566(.A1(new_n4636_), .A2(new_n4630_), .ZN(new_n4637_));
  INV_X1     g04567(.I(new_n4637_), .ZN(new_n4638_));
  INV_X1     g04568(.I(new_n4530_), .ZN(new_n4639_));
  AOI21_X1   g04569(.A1(new_n4564_), .A2(new_n101_), .B(new_n4639_), .ZN(new_n4640_));
  OAI21_X1   g04570(.A1(new_n4640_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n4641_));
  XOR2_X1    g04571(.A1(new_n4609_), .A2(new_n4641_), .Z(new_n4642_));
  AND2_X2    g04572(.A1(new_n4642_), .A2(new_n118_), .Z(new_n4643_));
  NOR2_X1    g04573(.A1(new_n4642_), .A2(new_n118_), .ZN(new_n4644_));
  OAI21_X1   g04574(.A1(new_n4643_), .A2(new_n4644_), .B(new_n4638_), .ZN(new_n4645_));
  XOR2_X1    g04575(.A1(new_n4642_), .A2(new_n71_), .Z(new_n4646_));
  OAI21_X1   g04576(.A1(new_n4638_), .A2(new_n4646_), .B(new_n4645_), .ZN(new_n4647_));
  NAND2_X1   g04577(.A1(new_n4647_), .A2(new_n4621_), .ZN(new_n4648_));
  INV_X1     g04578(.I(new_n4648_), .ZN(new_n4649_));
  XNOR2_X1   g04579(.A1(new_n4060_), .A2(new_n4053_), .ZN(new_n4650_));
  OAI21_X1   g04580(.A1(new_n4062_), .A2(new_n4342_), .B(new_n4341_), .ZN(new_n4651_));
  OAI21_X1   g04581(.A1(new_n4341_), .A2(new_n4650_), .B(new_n4651_), .ZN(new_n4652_));
  NOR2_X1    g04582(.A1(new_n4060_), .A2(new_n88_), .ZN(new_n4653_));
  INV_X1     g04583(.I(new_n4653_), .ZN(new_n4654_));
  AOI22_X1   g04584(.A1(new_n4071_), .A2(new_n4406_), .B1(new_n962_), .B2(new_n4054_), .ZN(new_n4655_));
  AOI21_X1   g04585(.A1(new_n4655_), .A2(new_n4654_), .B(new_n82_), .ZN(new_n4656_));
  NAND2_X1   g04586(.A1(new_n4652_), .A2(new_n4656_), .ZN(new_n4657_));
  INV_X1     g04587(.I(new_n4657_), .ZN(new_n4658_));
  XNOR2_X1   g04588(.A1(\a[15] ), .A2(\a[17] ), .ZN(new_n4659_));
  NOR2_X1    g04589(.A1(new_n442_), .A2(new_n4659_), .ZN(new_n4660_));
  INV_X1     g04590(.I(new_n1622_), .ZN(new_n4661_));
  XNOR2_X1   g04591(.A1(\a[14] ), .A2(\a[17] ), .ZN(new_n4662_));
  NOR3_X1    g04592(.A1(new_n442_), .A2(new_n1468_), .A3(new_n4662_), .ZN(new_n4663_));
  NOR3_X1    g04593(.A1(new_n4661_), .A2(new_n4663_), .A3(new_n4660_), .ZN(new_n4664_));
  NOR2_X1    g04594(.A1(new_n4664_), .A2(new_n126_), .ZN(new_n4665_));
  INV_X1     g04595(.I(new_n4665_), .ZN(new_n4666_));
  NAND2_X1   g04596(.A1(new_n4664_), .A2(new_n126_), .ZN(new_n4667_));
  AND2_X2    g04597(.A1(new_n4666_), .A2(new_n4667_), .Z(new_n4668_));
  INV_X1     g04598(.I(new_n4348_), .ZN(new_n4669_));
  OAI21_X1   g04599(.A1(new_n4044_), .A2(new_n4349_), .B(new_n4669_), .ZN(new_n4670_));
  XNOR2_X1   g04600(.A1(new_n4042_), .A2(new_n4035_), .ZN(new_n4671_));
  OAI21_X1   g04601(.A1(new_n4669_), .A2(new_n4671_), .B(new_n4670_), .ZN(new_n4672_));
  NAND2_X1   g04602(.A1(new_n4043_), .A2(new_n87_), .ZN(new_n4673_));
  AOI22_X1   g04603(.A1(new_n4036_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n4054_), .ZN(new_n4674_));
  AOI21_X1   g04604(.A1(new_n4673_), .A2(new_n4674_), .B(new_n82_), .ZN(new_n4675_));
  NAND2_X1   g04605(.A1(new_n4672_), .A2(new_n4675_), .ZN(new_n4676_));
  INV_X1     g04606(.I(new_n4676_), .ZN(new_n4677_));
  NOR2_X1    g04607(.A1(new_n4677_), .A2(new_n4668_), .ZN(new_n4678_));
  INV_X1     g04608(.I(new_n4678_), .ZN(new_n4679_));
  INV_X1     g04609(.I(new_n4668_), .ZN(new_n4680_));
  NOR2_X1    g04610(.A1(new_n4676_), .A2(new_n4680_), .ZN(new_n4681_));
  AOI21_X1   g04611(.A1(new_n4679_), .A2(new_n4658_), .B(new_n4681_), .ZN(new_n4682_));
  OAI22_X1   g04612(.A1(new_n4350_), .A2(new_n4044_), .B1(new_n4037_), .B2(new_n4352_), .ZN(new_n4683_));
  NOR2_X1    g04613(.A1(new_n4029_), .A2(new_n4035_), .ZN(new_n4684_));
  NOR2_X1    g04614(.A1(new_n4036_), .A2(new_n4028_), .ZN(new_n4685_));
  OAI21_X1   g04615(.A1(new_n4684_), .A2(new_n4685_), .B(new_n4351_), .ZN(new_n4686_));
  NAND2_X1   g04616(.A1(new_n4686_), .A2(new_n4683_), .ZN(new_n4687_));
  NOR2_X1    g04617(.A1(new_n4035_), .A2(new_n88_), .ZN(new_n4688_));
  INV_X1     g04618(.I(new_n4688_), .ZN(new_n4689_));
  AOI22_X1   g04619(.A1(new_n4029_), .A2(new_n962_), .B1(new_n4043_), .B2(new_n4406_), .ZN(new_n4690_));
  AOI21_X1   g04620(.A1(new_n4690_), .A2(new_n4689_), .B(new_n82_), .ZN(new_n4691_));
  NAND2_X1   g04621(.A1(new_n4687_), .A2(new_n4691_), .ZN(new_n4692_));
  AOI22_X1   g04622(.A1(new_n4018_), .A2(new_n4570_), .B1(new_n4375_), .B2(new_n4526_), .ZN(new_n4693_));
  AOI21_X1   g04623(.A1(new_n101_), .A2(new_n4399_), .B(new_n4693_), .ZN(new_n4694_));
  OAI21_X1   g04624(.A1(new_n4694_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n4695_));
  XOR2_X1    g04625(.A1(new_n4403_), .A2(new_n4695_), .Z(new_n4696_));
  INV_X1     g04626(.I(new_n4696_), .ZN(new_n4697_));
  NOR2_X1    g04627(.A1(new_n4697_), .A2(new_n4692_), .ZN(new_n4698_));
  NOR2_X1    g04628(.A1(new_n4698_), .A2(new_n4682_), .ZN(new_n4699_));
  INV_X1     g04629(.I(new_n4692_), .ZN(new_n4700_));
  NOR2_X1    g04630(.A1(new_n4696_), .A2(new_n4700_), .ZN(new_n4701_));
  NOR2_X1    g04631(.A1(new_n4699_), .A2(new_n4701_), .ZN(new_n4702_));
  XOR2_X1    g04632(.A1(new_n4017_), .A2(new_n4029_), .Z(new_n4703_));
  OAI21_X1   g04633(.A1(new_n4030_), .A2(new_n4355_), .B(new_n4354_), .ZN(new_n4704_));
  OAI21_X1   g04634(.A1(new_n4354_), .A2(new_n4703_), .B(new_n4704_), .ZN(new_n4705_));
  NAND2_X1   g04635(.A1(new_n4018_), .A2(new_n962_), .ZN(new_n4706_));
  NOR2_X1    g04636(.A1(new_n4352_), .A2(new_n4545_), .ZN(new_n4707_));
  AOI21_X1   g04637(.A1(new_n4706_), .A2(new_n4707_), .B(new_n82_), .ZN(new_n4708_));
  NAND2_X1   g04638(.A1(new_n4705_), .A2(new_n4708_), .ZN(new_n4709_));
  NOR2_X1    g04639(.A1(new_n4709_), .A2(new_n4700_), .ZN(new_n4710_));
  INV_X1     g04640(.I(new_n4709_), .ZN(new_n4711_));
  NOR2_X1    g04641(.A1(new_n4711_), .A2(new_n4692_), .ZN(new_n4712_));
  INV_X1     g04642(.I(new_n4712_), .ZN(new_n4713_));
  OAI21_X1   g04643(.A1(new_n4702_), .A2(new_n4710_), .B(new_n4713_), .ZN(new_n4714_));
  INV_X1     g04644(.I(new_n4714_), .ZN(new_n4715_));
  XNOR2_X1   g04645(.A1(\a[18] ), .A2(\a[20] ), .ZN(new_n4716_));
  NOR2_X1    g04646(.A1(new_n355_), .A2(new_n4716_), .ZN(new_n4717_));
  NOR2_X1    g04647(.A1(new_n269_), .A2(\a[18] ), .ZN(new_n4718_));
  AOI21_X1   g04648(.A1(\a[18] ), .A2(new_n354_), .B(new_n4718_), .ZN(new_n4719_));
  INV_X1     g04649(.I(new_n4719_), .ZN(new_n4720_));
  XNOR2_X1   g04650(.A1(\a[17] ), .A2(\a[20] ), .ZN(new_n4721_));
  NOR3_X1    g04651(.A1(new_n355_), .A2(new_n1467_), .A3(new_n4721_), .ZN(new_n4722_));
  NOR3_X1    g04652(.A1(new_n4720_), .A2(new_n4717_), .A3(new_n4722_), .ZN(new_n4723_));
  NOR2_X1    g04653(.A1(new_n4723_), .A2(new_n90_), .ZN(new_n4724_));
  INV_X1     g04654(.I(new_n4724_), .ZN(new_n4725_));
  NAND2_X1   g04655(.A1(new_n4723_), .A2(new_n90_), .ZN(new_n4726_));
  AND2_X2    g04656(.A1(new_n4725_), .A2(new_n4726_), .Z(new_n4727_));
  NAND2_X1   g04657(.A1(new_n4356_), .A2(new_n4377_), .ZN(new_n4728_));
  OAI21_X1   g04658(.A1(new_n4442_), .A2(new_n4444_), .B(new_n4441_), .ZN(new_n4729_));
  NAND2_X1   g04659(.A1(new_n4729_), .A2(new_n4728_), .ZN(new_n4730_));
  NAND2_X1   g04660(.A1(new_n4018_), .A2(new_n87_), .ZN(new_n4731_));
  AOI22_X1   g04661(.A1(new_n4375_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n4029_), .ZN(new_n4732_));
  AOI21_X1   g04662(.A1(new_n4731_), .A2(new_n4732_), .B(new_n82_), .ZN(new_n4733_));
  NAND2_X1   g04663(.A1(new_n4730_), .A2(new_n4733_), .ZN(new_n4734_));
  XOR2_X1    g04664(.A1(new_n4734_), .A2(new_n4711_), .Z(new_n4735_));
  NOR2_X1    g04665(.A1(new_n4735_), .A2(new_n4727_), .ZN(new_n4736_));
  INV_X1     g04666(.I(new_n4727_), .ZN(new_n4737_));
  AOI21_X1   g04667(.A1(new_n4730_), .A2(new_n4733_), .B(new_n4711_), .ZN(new_n4738_));
  NOR2_X1    g04668(.A1(new_n4734_), .A2(new_n4709_), .ZN(new_n4739_));
  NOR2_X1    g04669(.A1(new_n4739_), .A2(new_n4738_), .ZN(new_n4740_));
  NOR2_X1    g04670(.A1(new_n4740_), .A2(new_n4737_), .ZN(new_n4741_));
  NOR2_X1    g04671(.A1(new_n4736_), .A2(new_n4741_), .ZN(new_n4742_));
  AOI22_X1   g04672(.A1(new_n4438_), .A2(new_n4526_), .B1(new_n4399_), .B2(new_n4570_), .ZN(new_n4743_));
  AOI21_X1   g04673(.A1(new_n101_), .A2(new_n4469_), .B(new_n4743_), .ZN(new_n4744_));
  OAI21_X1   g04674(.A1(new_n4744_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n4745_));
  XNOR2_X1   g04675(.A1(new_n4477_), .A2(new_n4745_), .ZN(new_n4746_));
  AND2_X2    g04676(.A1(new_n4746_), .A2(new_n4742_), .Z(new_n4747_));
  NOR2_X1    g04677(.A1(new_n4747_), .A2(new_n4715_), .ZN(new_n4748_));
  NOR2_X1    g04678(.A1(new_n4746_), .A2(new_n4742_), .ZN(new_n4749_));
  NOR2_X1    g04679(.A1(new_n4748_), .A2(new_n4749_), .ZN(new_n4750_));
  INV_X1     g04680(.I(new_n4738_), .ZN(new_n4751_));
  AOI21_X1   g04681(.A1(new_n4751_), .A2(new_n4727_), .B(new_n4739_), .ZN(new_n4752_));
  AOI22_X1   g04682(.A1(new_n4438_), .A2(new_n4570_), .B1(new_n4469_), .B2(new_n4526_), .ZN(new_n4753_));
  AOI21_X1   g04683(.A1(new_n101_), .A2(new_n4555_), .B(new_n4753_), .ZN(new_n4754_));
  OAI21_X1   g04684(.A1(new_n4754_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n4755_));
  XNOR2_X1   g04685(.A1(new_n4584_), .A2(new_n4755_), .ZN(new_n4756_));
  XOR2_X1    g04686(.A1(new_n4756_), .A2(new_n4409_), .Z(new_n4757_));
  NOR2_X1    g04687(.A1(new_n4757_), .A2(new_n4752_), .ZN(new_n4758_));
  INV_X1     g04688(.I(new_n4752_), .ZN(new_n4759_));
  AND2_X2    g04689(.A1(new_n4756_), .A2(new_n4488_), .Z(new_n4760_));
  NOR2_X1    g04690(.A1(new_n4756_), .A2(new_n4488_), .ZN(new_n4761_));
  NOR2_X1    g04691(.A1(new_n4760_), .A2(new_n4761_), .ZN(new_n4762_));
  NOR2_X1    g04692(.A1(new_n4762_), .A2(new_n4759_), .ZN(new_n4763_));
  NOR2_X1    g04693(.A1(new_n4763_), .A2(new_n4758_), .ZN(new_n4764_));
  NOR2_X1    g04694(.A1(new_n4564_), .A2(new_n1128_), .ZN(new_n4765_));
  XNOR2_X1   g04695(.A1(\a[23] ), .A2(\a[26] ), .ZN(new_n4766_));
  NOR3_X1    g04696(.A1(new_n70_), .A2(new_n1120_), .A3(new_n4766_), .ZN(new_n4767_));
  AOI22_X1   g04697(.A1(new_n4518_), .A2(new_n4613_), .B1(new_n4564_), .B2(new_n4767_), .ZN(new_n4768_));
  OAI21_X1   g04698(.A1(new_n4768_), .A2(new_n4765_), .B(new_n65_), .ZN(new_n4769_));
  NAND2_X1   g04699(.A1(new_n4769_), .A2(new_n117_), .ZN(new_n4770_));
  XNOR2_X1   g04700(.A1(new_n4594_), .A2(new_n4770_), .ZN(new_n4771_));
  INV_X1     g04701(.I(new_n4771_), .ZN(new_n4772_));
  NOR2_X1    g04702(.A1(new_n4764_), .A2(new_n4772_), .ZN(new_n4773_));
  NOR2_X1    g04703(.A1(new_n4773_), .A2(new_n4750_), .ZN(new_n4774_));
  NOR3_X1    g04704(.A1(new_n4763_), .A2(new_n4758_), .A3(new_n4771_), .ZN(new_n4775_));
  NOR2_X1    g04705(.A1(new_n4774_), .A2(new_n4775_), .ZN(new_n4776_));
  XOR2_X1    g04706(.A1(new_n4534_), .A2(new_n4550_), .Z(new_n4777_));
  OAI21_X1   g04707(.A1(new_n4551_), .A2(new_n4553_), .B(new_n4488_), .ZN(new_n4778_));
  OAI21_X1   g04708(.A1(new_n4777_), .A2(new_n4488_), .B(new_n4778_), .ZN(new_n4779_));
  INV_X1     g04709(.I(new_n4779_), .ZN(new_n4780_));
  INV_X1     g04710(.I(new_n4767_), .ZN(new_n4781_));
  NOR2_X1    g04711(.A1(new_n4781_), .A2(new_n4612_), .ZN(new_n4782_));
  INV_X1     g04712(.I(new_n4782_), .ZN(new_n4783_));
  AOI21_X1   g04713(.A1(new_n4564_), .A2(new_n117_), .B(new_n4783_), .ZN(new_n4784_));
  OAI21_X1   g04714(.A1(new_n4784_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n4785_));
  XOR2_X1    g04715(.A1(new_n4609_), .A2(new_n4785_), .Z(new_n4786_));
  INV_X1     g04716(.I(new_n4786_), .ZN(new_n4787_));
  INV_X1     g04717(.I(new_n4760_), .ZN(new_n4788_));
  AOI21_X1   g04718(.A1(new_n4788_), .A2(new_n4759_), .B(new_n4761_), .ZN(new_n4789_));
  XOR2_X1    g04719(.A1(new_n4789_), .A2(new_n4787_), .Z(new_n4790_));
  NOR2_X1    g04720(.A1(new_n4790_), .A2(new_n4780_), .ZN(new_n4791_));
  AND2_X2    g04721(.A1(new_n4789_), .A2(new_n4786_), .Z(new_n4792_));
  NOR2_X1    g04722(.A1(new_n4789_), .A2(new_n4786_), .ZN(new_n4793_));
  NOR2_X1    g04723(.A1(new_n4792_), .A2(new_n4793_), .ZN(new_n4794_));
  NOR2_X1    g04724(.A1(new_n4794_), .A2(new_n4779_), .ZN(new_n4795_));
  NOR2_X1    g04725(.A1(new_n4795_), .A2(new_n4791_), .ZN(new_n4796_));
  INV_X1     g04726(.I(new_n4796_), .ZN(new_n4797_));
  NOR2_X1    g04727(.A1(new_n4797_), .A2(new_n189_), .ZN(new_n4798_));
  NOR2_X1    g04728(.A1(new_n4798_), .A2(new_n4776_), .ZN(new_n4799_));
  NOR2_X1    g04729(.A1(new_n4796_), .A2(new_n248_), .ZN(new_n4800_));
  NOR2_X1    g04730(.A1(new_n4799_), .A2(new_n4800_), .ZN(new_n4801_));
  INV_X1     g04731(.I(new_n4776_), .ZN(new_n4802_));
  OAI21_X1   g04732(.A1(new_n4798_), .A2(new_n4800_), .B(new_n4802_), .ZN(new_n4803_));
  XOR2_X1    g04733(.A1(new_n4796_), .A2(new_n189_), .Z(new_n4804_));
  OAI21_X1   g04734(.A1(new_n4802_), .A2(new_n4804_), .B(new_n4803_), .ZN(new_n4805_));
  INV_X1     g04735(.I(new_n4805_), .ZN(new_n4806_));
  NOR2_X1    g04736(.A1(new_n4773_), .A2(new_n4775_), .ZN(new_n4807_));
  XOR2_X1    g04737(.A1(new_n4764_), .A2(new_n4772_), .Z(new_n4808_));
  NAND2_X1   g04738(.A1(new_n4808_), .A2(new_n4750_), .ZN(new_n4809_));
  OAI21_X1   g04739(.A1(new_n4750_), .A2(new_n4807_), .B(new_n4809_), .ZN(new_n4810_));
  OAI21_X1   g04740(.A1(new_n4747_), .A2(new_n4749_), .B(new_n4714_), .ZN(new_n4811_));
  XOR2_X1    g04741(.A1(new_n4746_), .A2(new_n4742_), .Z(new_n4812_));
  NAND2_X1   g04742(.A1(new_n4812_), .A2(new_n4715_), .ZN(new_n4813_));
  NAND2_X1   g04743(.A1(new_n4813_), .A2(new_n4811_), .ZN(new_n4814_));
  INV_X1     g04744(.I(new_n4814_), .ZN(new_n4815_));
  OAI22_X1   g04745(.A1(new_n4516_), .A2(new_n1128_), .B1(new_n4531_), .B2(new_n4782_), .ZN(new_n4816_));
  AOI21_X1   g04746(.A1(new_n4816_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n4817_));
  XOR2_X1    g04747(.A1(new_n4524_), .A2(new_n4817_), .Z(new_n4818_));
  OAI22_X1   g04748(.A1(new_n4437_), .A2(new_n79_), .B1(new_n4530_), .B2(new_n4546_), .ZN(new_n4819_));
  AOI21_X1   g04749(.A1(new_n4819_), .A2(new_n72_), .B(new_n79_), .ZN(new_n4820_));
  XOR2_X1    g04750(.A1(new_n4541_), .A2(new_n4820_), .Z(new_n4821_));
  NOR2_X1    g04751(.A1(new_n4818_), .A2(new_n4821_), .ZN(new_n4822_));
  INV_X1     g04752(.I(new_n4822_), .ZN(new_n4823_));
  XOR2_X1    g04753(.A1(new_n4709_), .A2(new_n4692_), .Z(new_n4824_));
  NOR2_X1    g04754(.A1(new_n4702_), .A2(new_n4824_), .ZN(new_n4825_));
  NOR2_X1    g04755(.A1(new_n4712_), .A2(new_n4710_), .ZN(new_n4826_));
  INV_X1     g04756(.I(new_n4826_), .ZN(new_n4827_));
  AOI21_X1   g04757(.A1(new_n4702_), .A2(new_n4827_), .B(new_n4825_), .ZN(new_n4828_));
  INV_X1     g04758(.I(new_n4828_), .ZN(new_n4829_));
  INV_X1     g04759(.I(new_n4818_), .ZN(new_n4830_));
  INV_X1     g04760(.I(new_n4821_), .ZN(new_n4831_));
  NOR2_X1    g04761(.A1(new_n4830_), .A2(new_n4831_), .ZN(new_n4832_));
  OAI21_X1   g04762(.A1(new_n4829_), .A2(new_n4832_), .B(new_n4823_), .ZN(new_n4833_));
  AOI22_X1   g04763(.A1(new_n4518_), .A2(new_n4767_), .B1(new_n4555_), .B2(new_n4613_), .ZN(new_n4834_));
  AOI21_X1   g04764(.A1(new_n117_), .A2(new_n4564_), .B(new_n4834_), .ZN(new_n4835_));
  OAI21_X1   g04765(.A1(new_n4835_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n4836_));
  XOR2_X1    g04766(.A1(new_n4569_), .A2(new_n4836_), .Z(new_n4837_));
  INV_X1     g04767(.I(new_n4837_), .ZN(new_n4838_));
  NOR2_X1    g04768(.A1(new_n4838_), .A2(new_n4833_), .ZN(new_n4839_));
  NAND2_X1   g04769(.A1(new_n4838_), .A2(new_n4833_), .ZN(new_n4840_));
  OAI21_X1   g04770(.A1(new_n4815_), .A2(new_n4839_), .B(new_n4840_), .ZN(new_n4841_));
  NAND3_X1   g04771(.A1(new_n4563_), .A2(new_n247_), .A3(new_n1973_), .ZN(new_n4842_));
  AOI21_X1   g04772(.A1(new_n4842_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n4843_));
  XNOR2_X1   g04773(.A1(new_n4610_), .A2(new_n4843_), .ZN(new_n4844_));
  INV_X1     g04774(.I(new_n4844_), .ZN(new_n4845_));
  NOR2_X1    g04775(.A1(new_n4841_), .A2(new_n4845_), .ZN(new_n4846_));
  INV_X1     g04776(.I(new_n4846_), .ZN(new_n4847_));
  NAND2_X1   g04777(.A1(new_n4841_), .A2(new_n4845_), .ZN(new_n4848_));
  INV_X1     g04778(.I(new_n4848_), .ZN(new_n4849_));
  AOI21_X1   g04779(.A1(new_n4810_), .A2(new_n4847_), .B(new_n4849_), .ZN(new_n4850_));
  NAND2_X1   g04780(.A1(new_n4806_), .A2(new_n4850_), .ZN(new_n4851_));
  NOR2_X1    g04781(.A1(new_n4851_), .A2(new_n4801_), .ZN(new_n4852_));
  INV_X1     g04782(.I(new_n4852_), .ZN(new_n4853_));
  XOR2_X1    g04783(.A1(new_n4818_), .A2(new_n4831_), .Z(new_n4854_));
  OAI21_X1   g04784(.A1(new_n4832_), .A2(new_n4822_), .B(new_n4828_), .ZN(new_n4855_));
  OAI21_X1   g04785(.A1(new_n4828_), .A2(new_n4854_), .B(new_n4855_), .ZN(new_n4856_));
  INV_X1     g04786(.I(new_n4856_), .ZN(new_n4857_));
  OAI22_X1   g04787(.A1(new_n4017_), .A2(new_n79_), .B1(new_n4352_), .B2(new_n4530_), .ZN(new_n4858_));
  AOI21_X1   g04788(.A1(new_n4858_), .A2(new_n72_), .B(new_n79_), .ZN(new_n4859_));
  XNOR2_X1   g04789(.A1(new_n4705_), .A2(new_n4859_), .ZN(new_n4860_));
  INV_X1     g04790(.I(new_n4860_), .ZN(new_n4861_));
  OAI21_X1   g04791(.A1(new_n4055_), .A2(new_n4346_), .B(new_n4345_), .ZN(new_n4862_));
  XOR2_X1    g04792(.A1(new_n4042_), .A2(new_n4054_), .Z(new_n4863_));
  OAI21_X1   g04793(.A1(new_n4345_), .A2(new_n4863_), .B(new_n4862_), .ZN(new_n4864_));
  NOR2_X1    g04794(.A1(new_n4042_), .A2(new_n511_), .ZN(new_n4865_));
  INV_X1     g04795(.I(new_n4865_), .ZN(new_n4866_));
  AOI22_X1   g04796(.A1(new_n4406_), .A2(new_n4061_), .B1(new_n4054_), .B2(new_n87_), .ZN(new_n4867_));
  AOI21_X1   g04797(.A1(new_n4866_), .A2(new_n4867_), .B(new_n82_), .ZN(new_n4868_));
  NAND2_X1   g04798(.A1(new_n4864_), .A2(new_n4868_), .ZN(new_n4869_));
  INV_X1     g04799(.I(new_n4869_), .ZN(new_n4870_));
  NOR2_X1    g04800(.A1(new_n4861_), .A2(new_n4870_), .ZN(new_n4871_));
  NOR2_X1    g04801(.A1(new_n4871_), .A2(new_n4658_), .ZN(new_n4872_));
  NOR2_X1    g04802(.A1(new_n4860_), .A2(new_n4869_), .ZN(new_n4873_));
  NOR2_X1    g04803(.A1(new_n4872_), .A2(new_n4873_), .ZN(new_n4874_));
  OAI21_X1   g04804(.A1(new_n4678_), .A2(new_n4681_), .B(new_n4658_), .ZN(new_n4875_));
  XOR2_X1    g04805(.A1(new_n4676_), .A2(new_n4668_), .Z(new_n4876_));
  OAI21_X1   g04806(.A1(new_n4658_), .A2(new_n4876_), .B(new_n4875_), .ZN(new_n4877_));
  AOI22_X1   g04807(.A1(new_n4018_), .A2(new_n4526_), .B1(new_n4029_), .B2(new_n4570_), .ZN(new_n4878_));
  AOI21_X1   g04808(.A1(new_n101_), .A2(new_n4375_), .B(new_n4878_), .ZN(new_n4879_));
  OAI21_X1   g04809(.A1(new_n4879_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n4880_));
  XOR2_X1    g04810(.A1(new_n4730_), .A2(new_n4880_), .Z(new_n4881_));
  INV_X1     g04811(.I(new_n4881_), .ZN(new_n4882_));
  NOR2_X1    g04812(.A1(new_n4882_), .A2(new_n4877_), .ZN(new_n4883_));
  NOR2_X1    g04813(.A1(new_n4874_), .A2(new_n4883_), .ZN(new_n4884_));
  INV_X1     g04814(.I(new_n4877_), .ZN(new_n4885_));
  NOR2_X1    g04815(.A1(new_n4881_), .A2(new_n4885_), .ZN(new_n4886_));
  NOR2_X1    g04816(.A1(new_n4884_), .A2(new_n4886_), .ZN(new_n4887_));
  INV_X1     g04817(.I(new_n4887_), .ZN(new_n4888_));
  XOR2_X1    g04818(.A1(new_n4696_), .A2(new_n4692_), .Z(new_n4889_));
  OAI21_X1   g04819(.A1(new_n4698_), .A2(new_n4701_), .B(new_n4682_), .ZN(new_n4890_));
  OAI21_X1   g04820(.A1(new_n4889_), .A2(new_n4682_), .B(new_n4890_), .ZN(new_n4891_));
  INV_X1     g04821(.I(new_n4891_), .ZN(new_n4892_));
  AOI22_X1   g04822(.A1(new_n4438_), .A2(new_n4613_), .B1(new_n4469_), .B2(new_n4767_), .ZN(new_n4893_));
  AOI21_X1   g04823(.A1(new_n117_), .A2(new_n4555_), .B(new_n4893_), .ZN(new_n4894_));
  OAI21_X1   g04824(.A1(new_n4894_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n4895_));
  XNOR2_X1   g04825(.A1(new_n4584_), .A2(new_n4895_), .ZN(new_n4896_));
  INV_X1     g04826(.I(new_n4896_), .ZN(new_n4897_));
  NOR2_X1    g04827(.A1(new_n4897_), .A2(new_n4892_), .ZN(new_n4898_));
  INV_X1     g04828(.I(new_n4898_), .ZN(new_n4899_));
  NOR2_X1    g04829(.A1(new_n4896_), .A2(new_n4891_), .ZN(new_n4900_));
  AOI21_X1   g04830(.A1(new_n4899_), .A2(new_n4888_), .B(new_n4900_), .ZN(new_n4901_));
  INV_X1     g04831(.I(new_n4412_), .ZN(new_n4902_));
  NOR2_X1    g04832(.A1(new_n4564_), .A2(new_n4902_), .ZN(new_n4903_));
  NOR2_X1    g04833(.A1(new_n4563_), .A2(new_n1973_), .ZN(new_n4904_));
  OAI22_X1   g04834(.A1(new_n4903_), .A2(new_n4904_), .B1(new_n1239_), .B2(new_n4563_), .ZN(new_n4905_));
  AOI21_X1   g04835(.A1(new_n4905_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n4906_));
  XNOR2_X1   g04836(.A1(new_n4609_), .A2(new_n4906_), .ZN(new_n4907_));
  AND2_X2    g04837(.A1(new_n4901_), .A2(new_n4907_), .Z(new_n4908_));
  NOR2_X1    g04838(.A1(new_n4901_), .A2(new_n4907_), .ZN(new_n4909_));
  NOR2_X1    g04839(.A1(new_n4908_), .A2(new_n4909_), .ZN(new_n4910_));
  NOR2_X1    g04840(.A1(new_n4910_), .A2(new_n4857_), .ZN(new_n4911_));
  XNOR2_X1   g04841(.A1(new_n4901_), .A2(new_n4907_), .ZN(new_n4912_));
  NOR2_X1    g04842(.A1(new_n4912_), .A2(new_n4856_), .ZN(new_n4913_));
  NOR2_X1    g04843(.A1(new_n4911_), .A2(new_n4913_), .ZN(new_n4914_));
  OAI21_X1   g04844(.A1(new_n4898_), .A2(new_n4900_), .B(new_n4888_), .ZN(new_n4915_));
  XOR2_X1    g04845(.A1(new_n4896_), .A2(new_n4892_), .Z(new_n4916_));
  OAI21_X1   g04846(.A1(new_n4888_), .A2(new_n4916_), .B(new_n4915_), .ZN(new_n4917_));
  INV_X1     g04847(.I(new_n4917_), .ZN(new_n4918_));
  INV_X1     g04848(.I(new_n4874_), .ZN(new_n4919_));
  OAI21_X1   g04849(.A1(new_n4883_), .A2(new_n4886_), .B(new_n4919_), .ZN(new_n4920_));
  XOR2_X1    g04850(.A1(new_n4881_), .A2(new_n4877_), .Z(new_n4921_));
  OAI21_X1   g04851(.A1(new_n4919_), .A2(new_n4921_), .B(new_n4920_), .ZN(new_n4922_));
  INV_X1     g04852(.I(new_n4336_), .ZN(new_n4923_));
  AOI21_X1   g04853(.A1(new_n4084_), .A2(new_n4923_), .B(new_n4335_), .ZN(new_n4924_));
  XOR2_X1    g04854(.A1(new_n4070_), .A2(new_n4082_), .Z(new_n4925_));
  INV_X1     g04855(.I(new_n4925_), .ZN(new_n4926_));
  AOI21_X1   g04856(.A1(new_n4335_), .A2(new_n4926_), .B(new_n4924_), .ZN(new_n4927_));
  INV_X1     g04857(.I(new_n4927_), .ZN(new_n4928_));
  NAND2_X1   g04858(.A1(new_n4071_), .A2(new_n962_), .ZN(new_n4929_));
  AOI22_X1   g04859(.A1(new_n4082_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n4328_), .ZN(new_n4930_));
  AOI21_X1   g04860(.A1(new_n4929_), .A2(new_n4930_), .B(new_n82_), .ZN(new_n4931_));
  NAND2_X1   g04861(.A1(new_n4928_), .A2(new_n4931_), .ZN(new_n4932_));
  XOR2_X1    g04862(.A1(new_n4070_), .A2(new_n4061_), .Z(new_n4933_));
  OAI21_X1   g04863(.A1(new_n4072_), .A2(new_n4339_), .B(new_n4338_), .ZN(new_n4934_));
  OAI21_X1   g04864(.A1(new_n4338_), .A2(new_n4933_), .B(new_n4934_), .ZN(new_n4935_));
  NAND2_X1   g04865(.A1(new_n4071_), .A2(new_n87_), .ZN(new_n4936_));
  AOI22_X1   g04866(.A1(new_n4061_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n4082_), .ZN(new_n4937_));
  AOI21_X1   g04867(.A1(new_n4936_), .A2(new_n4937_), .B(new_n82_), .ZN(new_n4938_));
  NAND2_X1   g04868(.A1(new_n4935_), .A2(new_n4938_), .ZN(new_n4939_));
  NOR2_X1    g04869(.A1(new_n4939_), .A2(new_n4932_), .ZN(new_n4940_));
  INV_X1     g04870(.I(new_n1851_), .ZN(new_n4941_));
  XNOR2_X1   g04871(.A1(\a[11] ), .A2(\a[14] ), .ZN(new_n4942_));
  NOR3_X1    g04872(.A1(new_n784_), .A2(new_n1733_), .A3(new_n4942_), .ZN(new_n4943_));
  NOR3_X1    g04873(.A1(new_n4941_), .A2(new_n785_), .A3(new_n4943_), .ZN(new_n4944_));
  NOR2_X1    g04874(.A1(new_n4944_), .A2(new_n279_), .ZN(new_n4945_));
  INV_X1     g04875(.I(new_n4945_), .ZN(new_n4946_));
  NAND2_X1   g04876(.A1(new_n4944_), .A2(new_n279_), .ZN(new_n4947_));
  AND2_X2    g04877(.A1(new_n4946_), .A2(new_n4947_), .Z(new_n4948_));
  NAND2_X1   g04878(.A1(new_n4939_), .A2(new_n4932_), .ZN(new_n4949_));
  AOI21_X1   g04879(.A1(new_n4948_), .A2(new_n4949_), .B(new_n4940_), .ZN(new_n4950_));
  INV_X1     g04880(.I(new_n4950_), .ZN(new_n4951_));
  AOI22_X1   g04881(.A1(new_n4043_), .A2(new_n4570_), .B1(new_n4036_), .B2(new_n4526_), .ZN(new_n4952_));
  AOI21_X1   g04882(.A1(new_n101_), .A2(new_n4029_), .B(new_n4952_), .ZN(new_n4953_));
  OAI21_X1   g04883(.A1(new_n4953_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n4954_));
  XOR2_X1    g04884(.A1(new_n4687_), .A2(new_n4954_), .Z(new_n4955_));
  INV_X1     g04885(.I(new_n4955_), .ZN(new_n4956_));
  NOR2_X1    g04886(.A1(new_n4956_), .A2(new_n4657_), .ZN(new_n4957_));
  INV_X1     g04887(.I(new_n4957_), .ZN(new_n4958_));
  NOR2_X1    g04888(.A1(new_n4955_), .A2(new_n4658_), .ZN(new_n4959_));
  AOI21_X1   g04889(.A1(new_n4958_), .A2(new_n4951_), .B(new_n4959_), .ZN(new_n4960_));
  OAI22_X1   g04890(.A1(new_n4437_), .A2(new_n1128_), .B1(new_n4546_), .B2(new_n4782_), .ZN(new_n4961_));
  AOI21_X1   g04891(.A1(new_n4961_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n4962_));
  XOR2_X1    g04892(.A1(new_n4541_), .A2(new_n4962_), .Z(new_n4963_));
  NOR2_X1    g04893(.A1(new_n4963_), .A2(new_n4960_), .ZN(new_n4964_));
  INV_X1     g04894(.I(new_n4964_), .ZN(new_n4965_));
  XOR2_X1    g04895(.A1(new_n4860_), .A2(new_n4870_), .Z(new_n4966_));
  OAI21_X1   g04896(.A1(new_n4871_), .A2(new_n4873_), .B(new_n4658_), .ZN(new_n4967_));
  OAI21_X1   g04897(.A1(new_n4966_), .A2(new_n4658_), .B(new_n4967_), .ZN(new_n4968_));
  AND2_X2    g04898(.A1(new_n4963_), .A2(new_n4960_), .Z(new_n4969_));
  OAI21_X1   g04899(.A1(new_n4968_), .A2(new_n4969_), .B(new_n4965_), .ZN(new_n4970_));
  AOI22_X1   g04900(.A1(new_n4438_), .A2(new_n4767_), .B1(new_n4399_), .B2(new_n4613_), .ZN(new_n4971_));
  AOI21_X1   g04901(.A1(new_n117_), .A2(new_n4469_), .B(new_n4971_), .ZN(new_n4972_));
  OAI21_X1   g04902(.A1(new_n4972_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n4973_));
  XNOR2_X1   g04903(.A1(new_n4477_), .A2(new_n4973_), .ZN(new_n4974_));
  INV_X1     g04904(.I(new_n4974_), .ZN(new_n4975_));
  NOR2_X1    g04905(.A1(new_n4975_), .A2(new_n4970_), .ZN(new_n4976_));
  INV_X1     g04906(.I(new_n4976_), .ZN(new_n4977_));
  NAND2_X1   g04907(.A1(new_n4975_), .A2(new_n4970_), .ZN(new_n4978_));
  INV_X1     g04908(.I(new_n4978_), .ZN(new_n4979_));
  AOI21_X1   g04909(.A1(new_n4922_), .A2(new_n4977_), .B(new_n4979_), .ZN(new_n4980_));
  NOR2_X1    g04910(.A1(new_n4902_), .A2(new_n1973_), .ZN(new_n4981_));
  OAI22_X1   g04911(.A1(new_n4567_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4564_), .ZN(new_n4982_));
  AOI21_X1   g04912(.A1(new_n4982_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n4983_));
  XOR2_X1    g04913(.A1(new_n4594_), .A2(new_n4983_), .Z(new_n4984_));
  AND2_X2    g04914(.A1(new_n4980_), .A2(new_n4984_), .Z(new_n4985_));
  NOR2_X1    g04915(.A1(new_n4918_), .A2(new_n4985_), .ZN(new_n4986_));
  NOR2_X1    g04916(.A1(new_n4980_), .A2(new_n4984_), .ZN(new_n4987_));
  NOR2_X1    g04917(.A1(new_n4986_), .A2(new_n4987_), .ZN(new_n4988_));
  INV_X1     g04918(.I(new_n4988_), .ZN(new_n4989_));
  NOR2_X1    g04919(.A1(new_n4989_), .A2(new_n356_), .ZN(new_n4990_));
  NOR2_X1    g04920(.A1(new_n4990_), .A2(new_n4914_), .ZN(new_n4991_));
  NOR2_X1    g04921(.A1(new_n4988_), .A2(new_n273_), .ZN(new_n4992_));
  NOR2_X1    g04922(.A1(new_n4991_), .A2(new_n4992_), .ZN(new_n4993_));
  INV_X1     g04923(.I(new_n4908_), .ZN(new_n4994_));
  AOI21_X1   g04924(.A1(new_n4994_), .A2(new_n4856_), .B(new_n4909_), .ZN(new_n4995_));
  XNOR2_X1   g04925(.A1(new_n4833_), .A2(new_n4837_), .ZN(new_n4996_));
  NAND2_X1   g04926(.A1(new_n4996_), .A2(new_n4814_), .ZN(new_n4997_));
  INV_X1     g04927(.I(new_n4840_), .ZN(new_n4998_));
  OAI21_X1   g04928(.A1(new_n4998_), .A2(new_n4839_), .B(new_n4815_), .ZN(new_n4999_));
  NAND2_X1   g04929(.A1(new_n4997_), .A2(new_n4999_), .ZN(new_n5000_));
  XOR2_X1    g04930(.A1(new_n4609_), .A2(new_n4563_), .Z(new_n5001_));
  NOR2_X1    g04931(.A1(new_n4902_), .A2(new_n1239_), .ZN(new_n5002_));
  AOI21_X1   g04932(.A1(new_n1973_), .A2(new_n5002_), .B(new_n4563_), .ZN(new_n5003_));
  AOI21_X1   g04933(.A1(new_n5003_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n5004_));
  XNOR2_X1   g04934(.A1(new_n5001_), .A2(new_n5004_), .ZN(new_n5005_));
  INV_X1     g04935(.I(new_n5005_), .ZN(new_n5006_));
  XOR2_X1    g04936(.A1(new_n5000_), .A2(new_n5006_), .Z(new_n5007_));
  NOR2_X1    g04937(.A1(new_n5007_), .A2(new_n4995_), .ZN(new_n5008_));
  INV_X1     g04938(.I(new_n4995_), .ZN(new_n5009_));
  AOI21_X1   g04939(.A1(new_n4997_), .A2(new_n4999_), .B(new_n5006_), .ZN(new_n5010_));
  NOR2_X1    g04940(.A1(new_n5000_), .A2(new_n5005_), .ZN(new_n5011_));
  NOR2_X1    g04941(.A1(new_n5011_), .A2(new_n5010_), .ZN(new_n5012_));
  NOR2_X1    g04942(.A1(new_n5012_), .A2(new_n5009_), .ZN(new_n5013_));
  NOR2_X1    g04943(.A1(new_n5008_), .A2(new_n5013_), .ZN(new_n5014_));
  NOR2_X1    g04944(.A1(new_n5014_), .A2(new_n4993_), .ZN(new_n5015_));
  NOR2_X1    g04945(.A1(new_n3415_), .A2(\a[2] ), .ZN(new_n5016_));
  NAND3_X1   g04946(.A1(new_n4280_), .A2(new_n4135_), .A3(new_n4143_), .ZN(new_n5017_));
  NOR2_X1    g04947(.A1(new_n4286_), .A2(new_n4135_), .ZN(new_n5018_));
  INV_X1     g04948(.I(new_n5018_), .ZN(new_n5019_));
  AOI21_X1   g04949(.A1(new_n5019_), .A2(new_n5017_), .B(new_n4285_), .ZN(new_n5020_));
  INV_X1     g04950(.I(new_n4281_), .ZN(new_n5021_));
  AOI21_X1   g04951(.A1(new_n5021_), .A2(new_n4288_), .B(new_n4290_), .ZN(new_n5022_));
  OR2_X2     g04952(.A1(new_n5022_), .A2(new_n5020_), .Z(new_n5023_));
  NAND2_X1   g04953(.A1(new_n4290_), .A2(new_n962_), .ZN(new_n5024_));
  AOI22_X1   g04954(.A1(new_n4136_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n4143_), .ZN(new_n5025_));
  AOI21_X1   g04955(.A1(new_n5024_), .A2(new_n5025_), .B(new_n82_), .ZN(new_n5026_));
  NAND2_X1   g04956(.A1(new_n5023_), .A2(new_n5026_), .ZN(new_n5027_));
  NOR2_X1    g04957(.A1(new_n5027_), .A2(new_n5016_), .ZN(new_n5028_));
  INV_X1     g04958(.I(new_n5028_), .ZN(new_n5029_));
  INV_X1     g04959(.I(new_n5016_), .ZN(new_n5030_));
  INV_X1     g04960(.I(new_n3042_), .ZN(new_n5031_));
  XNOR2_X1   g04961(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n5032_));
  NOR3_X1    g04962(.A1(new_n2897_), .A2(new_n3419_), .A3(new_n5032_), .ZN(new_n5033_));
  NOR3_X1    g04963(.A1(new_n5031_), .A2(new_n5033_), .A3(new_n2898_), .ZN(new_n5034_));
  NOR2_X1    g04964(.A1(new_n5034_), .A2(new_n452_), .ZN(new_n5035_));
  INV_X1     g04965(.I(new_n5034_), .ZN(new_n5036_));
  NOR2_X1    g04966(.A1(new_n5036_), .A2(\a[5] ), .ZN(new_n5037_));
  NOR2_X1    g04967(.A1(new_n5037_), .A2(new_n5035_), .ZN(new_n5038_));
  XOR2_X1    g04968(.A1(new_n5038_), .A2(new_n5030_), .Z(new_n5039_));
  INV_X1     g04969(.I(new_n5039_), .ZN(new_n5040_));
  INV_X1     g04970(.I(new_n4309_), .ZN(new_n5041_));
  INV_X1     g04971(.I(new_n4131_), .ZN(new_n5042_));
  XOR2_X1    g04972(.A1(new_n4304_), .A2(new_n5042_), .Z(new_n5043_));
  NAND2_X1   g04973(.A1(new_n5043_), .A2(new_n5041_), .ZN(new_n5044_));
  NOR2_X1    g04974(.A1(new_n4304_), .A2(new_n5042_), .ZN(new_n5045_));
  NAND2_X1   g04975(.A1(new_n4304_), .A2(new_n5042_), .ZN(new_n5046_));
  INV_X1     g04976(.I(new_n5046_), .ZN(new_n5047_));
  OAI21_X1   g04977(.A1(new_n5047_), .A2(new_n5045_), .B(new_n4309_), .ZN(new_n5048_));
  NAND2_X1   g04978(.A1(new_n5044_), .A2(new_n5048_), .ZN(new_n5049_));
  NOR2_X1    g04979(.A1(new_n4131_), .A2(new_n88_), .ZN(new_n5050_));
  INV_X1     g04980(.I(new_n5050_), .ZN(new_n5051_));
  AOI22_X1   g04981(.A1(new_n5041_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n4297_), .ZN(new_n5052_));
  AOI21_X1   g04982(.A1(new_n5052_), .A2(new_n5051_), .B(new_n82_), .ZN(new_n5053_));
  NAND2_X1   g04983(.A1(new_n5049_), .A2(new_n5053_), .ZN(new_n5054_));
  INV_X1     g04984(.I(new_n5054_), .ZN(new_n5055_));
  NOR2_X1    g04985(.A1(new_n5055_), .A2(new_n5040_), .ZN(new_n5056_));
  NOR2_X1    g04986(.A1(new_n5056_), .A2(new_n5029_), .ZN(new_n5057_));
  NOR2_X1    g04987(.A1(new_n5054_), .A2(new_n5039_), .ZN(new_n5058_));
  NOR2_X1    g04988(.A1(new_n5057_), .A2(new_n5058_), .ZN(new_n5059_));
  NAND2_X1   g04989(.A1(new_n5038_), .A2(new_n5016_), .ZN(new_n5060_));
  NOR2_X1    g04990(.A1(new_n5047_), .A2(new_n5045_), .ZN(new_n5061_));
  XOR2_X1    g04991(.A1(new_n4304_), .A2(new_n4124_), .Z(new_n5062_));
  NOR2_X1    g04992(.A1(new_n5061_), .A2(new_n5062_), .ZN(new_n5063_));
  NAND2_X1   g04993(.A1(new_n5063_), .A2(new_n4309_), .ZN(new_n5064_));
  NOR2_X1    g04994(.A1(new_n5063_), .A2(new_n4309_), .ZN(new_n5065_));
  INV_X1     g04995(.I(new_n5065_), .ZN(new_n5066_));
  NAND2_X1   g04996(.A1(new_n5066_), .A2(new_n5064_), .ZN(new_n5067_));
  NAND2_X1   g04997(.A1(new_n5041_), .A2(new_n87_), .ZN(new_n5068_));
  AOI22_X1   g04998(.A1(new_n5042_), .A2(new_n4406_), .B1(new_n4124_), .B2(new_n962_), .ZN(new_n5069_));
  AOI21_X1   g04999(.A1(new_n5069_), .A2(new_n5068_), .B(new_n82_), .ZN(new_n5070_));
  NAND2_X1   g05000(.A1(new_n5067_), .A2(new_n5070_), .ZN(new_n5071_));
  XNOR2_X1   g05001(.A1(new_n5071_), .A2(new_n5060_), .ZN(new_n5072_));
  INV_X1     g05002(.I(new_n5072_), .ZN(new_n5073_));
  NAND2_X1   g05003(.A1(new_n4319_), .A2(new_n4314_), .ZN(new_n5074_));
  NOR2_X1    g05004(.A1(new_n4099_), .A2(new_n4105_), .ZN(new_n5075_));
  NOR2_X1    g05005(.A1(new_n4100_), .A2(new_n4315_), .ZN(new_n5076_));
  OAI21_X1   g05006(.A1(new_n5075_), .A2(new_n5076_), .B(new_n5074_), .ZN(new_n5077_));
  NOR2_X1    g05007(.A1(new_n4106_), .A2(new_n4320_), .ZN(new_n5078_));
  OR2_X2     g05008(.A1(new_n5074_), .A2(new_n5078_), .Z(new_n5079_));
  NAND2_X1   g05009(.A1(new_n5079_), .A2(new_n5077_), .ZN(new_n5080_));
  AOI22_X1   g05010(.A1(new_n4113_), .A2(new_n4570_), .B1(new_n4105_), .B2(new_n4526_), .ZN(new_n5081_));
  AOI21_X1   g05011(.A1(new_n101_), .A2(new_n4100_), .B(new_n5081_), .ZN(new_n5082_));
  OAI21_X1   g05012(.A1(new_n5082_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n5083_));
  XOR2_X1    g05013(.A1(new_n5080_), .A2(new_n5083_), .Z(new_n5084_));
  AND2_X2    g05014(.A1(new_n5084_), .A2(new_n5073_), .Z(new_n5085_));
  NOR2_X1    g05015(.A1(new_n5084_), .A2(new_n5073_), .ZN(new_n5086_));
  INV_X1     g05016(.I(new_n5086_), .ZN(new_n5087_));
  OAI21_X1   g05017(.A1(new_n5059_), .A2(new_n5085_), .B(new_n5087_), .ZN(new_n5088_));
  NAND2_X1   g05018(.A1(new_n5071_), .A2(new_n5060_), .ZN(new_n5089_));
  INV_X1     g05019(.I(new_n5089_), .ZN(new_n5090_));
  OAI21_X1   g05020(.A1(new_n4318_), .A2(new_n4316_), .B(new_n4113_), .ZN(new_n5091_));
  INV_X1     g05021(.I(new_n5091_), .ZN(new_n5092_));
  NAND2_X1   g05022(.A1(new_n4312_), .A2(new_n4123_), .ZN(new_n5093_));
  NAND2_X1   g05023(.A1(new_n4317_), .A2(new_n4124_), .ZN(new_n5094_));
  AOI21_X1   g05024(.A1(new_n5094_), .A2(new_n5093_), .B(new_n4113_), .ZN(new_n5095_));
  NOR2_X1    g05025(.A1(new_n5092_), .A2(new_n5095_), .ZN(new_n5096_));
  INV_X1     g05026(.I(new_n5096_), .ZN(new_n5097_));
  NOR2_X1    g05027(.A1(new_n4112_), .A2(new_n511_), .ZN(new_n5098_));
  INV_X1     g05028(.I(new_n5098_), .ZN(new_n5099_));
  AOI22_X1   g05029(.A1(new_n87_), .A2(new_n4124_), .B1(new_n5041_), .B2(new_n4406_), .ZN(new_n5100_));
  AOI21_X1   g05030(.A1(new_n5099_), .A2(new_n5100_), .B(new_n82_), .ZN(new_n5101_));
  NAND2_X1   g05031(.A1(new_n5097_), .A2(new_n5101_), .ZN(new_n5102_));
  INV_X1     g05032(.I(new_n5102_), .ZN(new_n5103_));
  NOR2_X1    g05033(.A1(new_n5103_), .A2(new_n5090_), .ZN(new_n5104_));
  INV_X1     g05034(.I(new_n5104_), .ZN(new_n5105_));
  NOR2_X1    g05035(.A1(new_n5102_), .A2(new_n5089_), .ZN(new_n5106_));
  AOI21_X1   g05036(.A1(new_n5088_), .A2(new_n5105_), .B(new_n5106_), .ZN(new_n5107_));
  INV_X1     g05037(.I(new_n2718_), .ZN(new_n5108_));
  XNOR2_X1   g05038(.A1(\a[5] ), .A2(\a[8] ), .ZN(new_n5109_));
  NOR3_X1    g05039(.A1(new_n2468_), .A2(new_n2583_), .A3(new_n5109_), .ZN(new_n5110_));
  NOR3_X1    g05040(.A1(new_n5108_), .A2(new_n5110_), .A3(new_n2469_), .ZN(new_n5111_));
  NOR2_X1    g05041(.A1(new_n5111_), .A2(new_n498_), .ZN(new_n5112_));
  INV_X1     g05042(.I(new_n5112_), .ZN(new_n5113_));
  NAND2_X1   g05043(.A1(new_n5111_), .A2(new_n498_), .ZN(new_n5114_));
  AND2_X2    g05044(.A1(new_n5113_), .A2(new_n5114_), .Z(new_n5115_));
  NOR3_X1    g05045(.A1(new_n4317_), .A2(new_n4113_), .A3(new_n4123_), .ZN(new_n5116_));
  NOR3_X1    g05046(.A1(new_n4312_), .A2(new_n4112_), .A3(new_n4124_), .ZN(new_n5117_));
  OAI21_X1   g05047(.A1(new_n5116_), .A2(new_n5117_), .B(new_n4105_), .ZN(new_n5118_));
  NOR2_X1    g05048(.A1(new_n4316_), .A2(new_n4112_), .ZN(new_n5119_));
  OAI21_X1   g05049(.A1(new_n5119_), .A2(new_n4313_), .B(new_n4315_), .ZN(new_n5120_));
  NAND2_X1   g05050(.A1(new_n5120_), .A2(new_n5118_), .ZN(new_n5121_));
  NAND2_X1   g05051(.A1(new_n4113_), .A2(new_n87_), .ZN(new_n5122_));
  AOI22_X1   g05052(.A1(new_n4105_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n4124_), .ZN(new_n5123_));
  AOI21_X1   g05053(.A1(new_n5122_), .A2(new_n5123_), .B(new_n82_), .ZN(new_n5124_));
  AOI21_X1   g05054(.A1(new_n5121_), .A2(new_n5124_), .B(new_n5115_), .ZN(new_n5125_));
  INV_X1     g05055(.I(new_n5115_), .ZN(new_n5126_));
  NAND2_X1   g05056(.A1(new_n5121_), .A2(new_n5124_), .ZN(new_n5127_));
  NOR2_X1    g05057(.A1(new_n5127_), .A2(new_n5126_), .ZN(new_n5128_));
  NOR2_X1    g05058(.A1(new_n5128_), .A2(new_n5125_), .ZN(new_n5129_));
  NOR2_X1    g05059(.A1(new_n5129_), .A2(new_n5090_), .ZN(new_n5130_));
  XOR2_X1    g05060(.A1(new_n5127_), .A2(new_n5115_), .Z(new_n5131_));
  NOR2_X1    g05061(.A1(new_n5131_), .A2(new_n5089_), .ZN(new_n5132_));
  NOR2_X1    g05062(.A1(new_n5132_), .A2(new_n5130_), .ZN(new_n5133_));
  INV_X1     g05063(.I(new_n5133_), .ZN(new_n5134_));
  XOR2_X1    g05064(.A1(new_n4090_), .A2(new_n4328_), .Z(new_n5135_));
  NOR2_X1    g05065(.A1(new_n4325_), .A2(new_n5135_), .ZN(new_n5136_));
  NOR2_X1    g05066(.A1(new_n4329_), .A2(new_n4332_), .ZN(new_n5137_));
  NOR2_X1    g05067(.A1(new_n4324_), .A2(new_n5137_), .ZN(new_n5138_));
  NOR2_X1    g05068(.A1(new_n5136_), .A2(new_n5138_), .ZN(new_n5139_));
  AOI22_X1   g05069(.A1(new_n4091_), .A2(new_n4526_), .B1(new_n4100_), .B2(new_n4570_), .ZN(new_n5140_));
  AOI21_X1   g05070(.A1(new_n101_), .A2(new_n4328_), .B(new_n5140_), .ZN(new_n5141_));
  OAI21_X1   g05071(.A1(new_n5141_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n5142_));
  XNOR2_X1   g05072(.A1(new_n5139_), .A2(new_n5142_), .ZN(new_n5143_));
  INV_X1     g05073(.I(new_n5143_), .ZN(new_n5144_));
  NOR2_X1    g05074(.A1(new_n5144_), .A2(new_n5134_), .ZN(new_n5145_));
  NOR2_X1    g05075(.A1(new_n5107_), .A2(new_n5145_), .ZN(new_n5146_));
  NOR2_X1    g05076(.A1(new_n5143_), .A2(new_n5133_), .ZN(new_n5147_));
  NOR2_X1    g05077(.A1(new_n5146_), .A2(new_n5147_), .ZN(new_n5148_));
  INV_X1     g05078(.I(new_n5125_), .ZN(new_n5149_));
  AOI21_X1   g05079(.A1(new_n5149_), .A2(new_n5089_), .B(new_n5128_), .ZN(new_n5150_));
  NOR2_X1    g05080(.A1(new_n4315_), .A2(new_n88_), .ZN(new_n5151_));
  INV_X1     g05081(.I(new_n5151_), .ZN(new_n5152_));
  AOI22_X1   g05082(.A1(new_n4113_), .A2(new_n4406_), .B1(new_n962_), .B2(new_n4100_), .ZN(new_n5153_));
  AOI21_X1   g05083(.A1(new_n5153_), .A2(new_n5152_), .B(new_n82_), .ZN(new_n5154_));
  NAND2_X1   g05084(.A1(new_n5080_), .A2(new_n5154_), .ZN(new_n5155_));
  XOR2_X1    g05085(.A1(new_n4081_), .A2(new_n4328_), .Z(new_n5156_));
  NOR2_X1    g05086(.A1(new_n5135_), .A2(new_n5156_), .ZN(new_n5157_));
  INV_X1     g05087(.I(new_n5157_), .ZN(new_n5158_));
  NOR2_X1    g05088(.A1(new_n5158_), .A2(new_n4324_), .ZN(new_n5159_));
  NAND2_X1   g05089(.A1(new_n5158_), .A2(new_n4324_), .ZN(new_n5160_));
  INV_X1     g05090(.I(new_n5160_), .ZN(new_n5161_));
  NOR2_X1    g05091(.A1(new_n5161_), .A2(new_n5159_), .ZN(new_n5162_));
  AOI22_X1   g05092(.A1(new_n4091_), .A2(new_n4570_), .B1(new_n4328_), .B2(new_n4526_), .ZN(new_n5163_));
  AOI21_X1   g05093(.A1(new_n101_), .A2(new_n4082_), .B(new_n5163_), .ZN(new_n5164_));
  OAI21_X1   g05094(.A1(new_n5164_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n5165_));
  XNOR2_X1   g05095(.A1(new_n5162_), .A2(new_n5165_), .ZN(new_n5166_));
  XOR2_X1    g05096(.A1(new_n5166_), .A2(new_n5155_), .Z(new_n5167_));
  NOR2_X1    g05097(.A1(new_n5167_), .A2(new_n5150_), .ZN(new_n5168_));
  INV_X1     g05098(.I(new_n5150_), .ZN(new_n5169_));
  INV_X1     g05099(.I(new_n5155_), .ZN(new_n5170_));
  AND2_X2    g05100(.A1(new_n5166_), .A2(new_n5170_), .Z(new_n5171_));
  NOR2_X1    g05101(.A1(new_n5166_), .A2(new_n5170_), .ZN(new_n5172_));
  NOR2_X1    g05102(.A1(new_n5171_), .A2(new_n5172_), .ZN(new_n5173_));
  NOR2_X1    g05103(.A1(new_n5173_), .A2(new_n5169_), .ZN(new_n5174_));
  NOR2_X1    g05104(.A1(new_n5174_), .A2(new_n5168_), .ZN(new_n5175_));
  AOI22_X1   g05105(.A1(new_n4071_), .A2(new_n4613_), .B1(new_n4061_), .B2(new_n4767_), .ZN(new_n5176_));
  AOI21_X1   g05106(.A1(new_n117_), .A2(new_n4054_), .B(new_n5176_), .ZN(new_n5177_));
  OAI21_X1   g05107(.A1(new_n5177_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n5178_));
  XOR2_X1    g05108(.A1(new_n4652_), .A2(new_n5178_), .Z(new_n5179_));
  INV_X1     g05109(.I(new_n5179_), .ZN(new_n5180_));
  NOR2_X1    g05110(.A1(new_n5180_), .A2(new_n5175_), .ZN(new_n5181_));
  NOR2_X1    g05111(.A1(new_n5181_), .A2(new_n5148_), .ZN(new_n5182_));
  NOR3_X1    g05112(.A1(new_n5179_), .A2(new_n5168_), .A3(new_n5174_), .ZN(new_n5183_));
  NOR2_X1    g05113(.A1(new_n5182_), .A2(new_n5183_), .ZN(new_n5184_));
  INV_X1     g05114(.I(new_n5184_), .ZN(new_n5185_));
  INV_X1     g05115(.I(new_n5171_), .ZN(new_n5186_));
  AOI21_X1   g05116(.A1(new_n5186_), .A2(new_n5169_), .B(new_n5172_), .ZN(new_n5187_));
  OAI22_X1   g05117(.A1(new_n4331_), .A2(new_n4529_), .B1(new_n4081_), .B2(new_n4527_), .ZN(new_n5188_));
  OAI21_X1   g05118(.A1(new_n4070_), .A2(new_n79_), .B(new_n5188_), .ZN(new_n5189_));
  AOI21_X1   g05119(.A1(new_n5189_), .A2(new_n72_), .B(new_n79_), .ZN(new_n5190_));
  XOR2_X1    g05120(.A1(new_n4927_), .A2(new_n5190_), .Z(new_n5191_));
  XOR2_X1    g05121(.A1(new_n4090_), .A2(new_n4100_), .Z(new_n5192_));
  NOR2_X1    g05122(.A1(new_n4322_), .A2(new_n5192_), .ZN(new_n5193_));
  NOR2_X1    g05123(.A1(new_n4101_), .A2(new_n4323_), .ZN(new_n5194_));
  NOR3_X1    g05124(.A1(new_n5194_), .A2(new_n4106_), .A3(new_n4321_), .ZN(new_n5195_));
  NOR2_X1    g05125(.A1(new_n5195_), .A2(new_n5193_), .ZN(new_n5196_));
  INV_X1     g05126(.I(new_n5196_), .ZN(new_n5197_));
  NOR2_X1    g05127(.A1(new_n4090_), .A2(new_n511_), .ZN(new_n5198_));
  INV_X1     g05128(.I(new_n5198_), .ZN(new_n5199_));
  AOI22_X1   g05129(.A1(new_n4100_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n4105_), .ZN(new_n5200_));
  AOI21_X1   g05130(.A1(new_n5199_), .A2(new_n5200_), .B(new_n82_), .ZN(new_n5201_));
  NAND2_X1   g05131(.A1(new_n5197_), .A2(new_n5201_), .ZN(new_n5202_));
  INV_X1     g05132(.I(new_n5202_), .ZN(new_n5203_));
  XOR2_X1    g05133(.A1(new_n5191_), .A2(new_n5203_), .Z(new_n5204_));
  NOR2_X1    g05134(.A1(new_n5204_), .A2(new_n5170_), .ZN(new_n5205_));
  AND2_X2    g05135(.A1(new_n5191_), .A2(new_n5202_), .Z(new_n5206_));
  NOR2_X1    g05136(.A1(new_n5191_), .A2(new_n5202_), .ZN(new_n5207_));
  NOR2_X1    g05137(.A1(new_n5206_), .A2(new_n5207_), .ZN(new_n5208_));
  NOR2_X1    g05138(.A1(new_n5208_), .A2(new_n5155_), .ZN(new_n5209_));
  NOR2_X1    g05139(.A1(new_n5209_), .A2(new_n5205_), .ZN(new_n5210_));
  NOR2_X1    g05140(.A1(new_n4060_), .A2(new_n4612_), .ZN(new_n5211_));
  NOR2_X1    g05141(.A1(new_n4053_), .A2(new_n4781_), .ZN(new_n5212_));
  OAI22_X1   g05142(.A1(new_n4042_), .A2(new_n1128_), .B1(new_n5211_), .B2(new_n5212_), .ZN(new_n5213_));
  AOI21_X1   g05143(.A1(new_n5213_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n5214_));
  INV_X1     g05144(.I(new_n5214_), .ZN(new_n5215_));
  NOR2_X1    g05145(.A1(new_n4864_), .A2(new_n5215_), .ZN(new_n5216_));
  INV_X1     g05146(.I(new_n4864_), .ZN(new_n5217_));
  NOR2_X1    g05147(.A1(new_n5217_), .A2(new_n5214_), .ZN(new_n5218_));
  NOR2_X1    g05148(.A1(new_n5218_), .A2(new_n5216_), .ZN(new_n5219_));
  INV_X1     g05149(.I(new_n5219_), .ZN(new_n5220_));
  NOR2_X1    g05150(.A1(new_n5220_), .A2(new_n5210_), .ZN(new_n5221_));
  INV_X1     g05151(.I(new_n5221_), .ZN(new_n5222_));
  NAND2_X1   g05152(.A1(new_n5220_), .A2(new_n5210_), .ZN(new_n5223_));
  AOI21_X1   g05153(.A1(new_n5222_), .A2(new_n5223_), .B(new_n5187_), .ZN(new_n5224_));
  INV_X1     g05154(.I(new_n5187_), .ZN(new_n5225_));
  XOR2_X1    g05155(.A1(new_n5219_), .A2(new_n5210_), .Z(new_n5226_));
  NOR2_X1    g05156(.A1(new_n5226_), .A2(new_n5225_), .ZN(new_n5227_));
  NOR2_X1    g05157(.A1(new_n5224_), .A2(new_n5227_), .ZN(new_n5228_));
  INV_X1     g05158(.I(new_n5228_), .ZN(new_n5229_));
  OAI22_X1   g05159(.A1(new_n4028_), .A2(new_n4902_), .B1(new_n1973_), .B2(new_n4035_), .ZN(new_n5230_));
  OAI21_X1   g05160(.A1(new_n4017_), .A2(new_n1239_), .B(new_n5230_), .ZN(new_n5231_));
  AOI21_X1   g05161(.A1(new_n5231_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n5232_));
  XNOR2_X1   g05162(.A1(new_n4705_), .A2(new_n5232_), .ZN(new_n5233_));
  INV_X1     g05163(.I(new_n5233_), .ZN(new_n5234_));
  NOR2_X1    g05164(.A1(new_n5234_), .A2(new_n5229_), .ZN(new_n5235_));
  INV_X1     g05165(.I(new_n5235_), .ZN(new_n5236_));
  NOR2_X1    g05166(.A1(new_n5233_), .A2(new_n5228_), .ZN(new_n5237_));
  AOI21_X1   g05167(.A1(new_n5236_), .A2(new_n5185_), .B(new_n5237_), .ZN(new_n5238_));
  AOI22_X1   g05168(.A1(new_n4071_), .A2(new_n4526_), .B1(new_n4082_), .B2(new_n4570_), .ZN(new_n5239_));
  AOI21_X1   g05169(.A1(new_n101_), .A2(new_n4061_), .B(new_n5239_), .ZN(new_n5240_));
  OAI21_X1   g05170(.A1(new_n5240_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n5241_));
  XOR2_X1    g05171(.A1(new_n4935_), .A2(new_n5241_), .Z(new_n5242_));
  INV_X1     g05172(.I(new_n5242_), .ZN(new_n5243_));
  NOR2_X1    g05173(.A1(new_n5206_), .A2(new_n5170_), .ZN(new_n5244_));
  NOR2_X1    g05174(.A1(new_n5244_), .A2(new_n5207_), .ZN(new_n5245_));
  INV_X1     g05175(.I(new_n5139_), .ZN(new_n5246_));
  INV_X1     g05176(.I(new_n2258_), .ZN(new_n5247_));
  XNOR2_X1   g05177(.A1(\a[8] ), .A2(\a[11] ), .ZN(new_n5248_));
  NOR3_X1    g05178(.A1(new_n804_), .A2(new_n2573_), .A3(new_n5248_), .ZN(new_n5249_));
  NOR3_X1    g05179(.A1(new_n5247_), .A2(new_n5249_), .A3(new_n805_), .ZN(new_n5250_));
  NOR2_X1    g05180(.A1(new_n5250_), .A2(new_n294_), .ZN(new_n5251_));
  INV_X1     g05181(.I(new_n5251_), .ZN(new_n5252_));
  NAND2_X1   g05182(.A1(new_n5250_), .A2(new_n294_), .ZN(new_n5253_));
  AND2_X2    g05183(.A1(new_n5252_), .A2(new_n5253_), .Z(new_n5254_));
  NAND2_X1   g05184(.A1(new_n4091_), .A2(new_n87_), .ZN(new_n5255_));
  AOI22_X1   g05185(.A1(new_n4328_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n4100_), .ZN(new_n5256_));
  AOI21_X1   g05186(.A1(new_n5255_), .A2(new_n5256_), .B(new_n82_), .ZN(new_n5257_));
  AOI21_X1   g05187(.A1(new_n5246_), .A2(new_n5257_), .B(new_n5254_), .ZN(new_n5258_));
  INV_X1     g05188(.I(new_n5254_), .ZN(new_n5259_));
  NAND2_X1   g05189(.A1(new_n5246_), .A2(new_n5257_), .ZN(new_n5260_));
  NOR2_X1    g05190(.A1(new_n5260_), .A2(new_n5259_), .ZN(new_n5261_));
  NOR2_X1    g05191(.A1(new_n5261_), .A2(new_n5258_), .ZN(new_n5262_));
  NOR2_X1    g05192(.A1(new_n5262_), .A2(new_n5155_), .ZN(new_n5263_));
  XOR2_X1    g05193(.A1(new_n5260_), .A2(new_n5254_), .Z(new_n5264_));
  NOR2_X1    g05194(.A1(new_n5264_), .A2(new_n5170_), .ZN(new_n5265_));
  NOR2_X1    g05195(.A1(new_n5265_), .A2(new_n5263_), .ZN(new_n5266_));
  XOR2_X1    g05196(.A1(new_n5245_), .A2(new_n5266_), .Z(new_n5267_));
  OAI21_X1   g05197(.A1(new_n5187_), .A2(new_n5221_), .B(new_n5223_), .ZN(new_n5268_));
  AOI22_X1   g05198(.A1(new_n4043_), .A2(new_n4767_), .B1(new_n4054_), .B2(new_n4613_), .ZN(new_n5269_));
  AOI21_X1   g05199(.A1(new_n117_), .A2(new_n4036_), .B(new_n5269_), .ZN(new_n5270_));
  OAI21_X1   g05200(.A1(new_n5270_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n5271_));
  XOR2_X1    g05201(.A1(new_n4672_), .A2(new_n5271_), .Z(new_n5272_));
  INV_X1     g05202(.I(new_n5272_), .ZN(new_n5273_));
  XOR2_X1    g05203(.A1(new_n5268_), .A2(new_n5273_), .Z(new_n5274_));
  XOR2_X1    g05204(.A1(new_n5274_), .A2(new_n5267_), .Z(new_n5275_));
  XOR2_X1    g05205(.A1(new_n5275_), .A2(new_n5243_), .Z(new_n5276_));
  OAI22_X1   g05206(.A1(new_n4355_), .A2(new_n4981_), .B1(new_n4374_), .B2(new_n1239_), .ZN(new_n5277_));
  AOI21_X1   g05207(.A1(new_n5277_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n5278_));
  XNOR2_X1   g05208(.A1(new_n4730_), .A2(new_n5278_), .ZN(new_n5279_));
  INV_X1     g05209(.I(new_n5279_), .ZN(new_n5280_));
  NOR2_X1    g05210(.A1(new_n5276_), .A2(new_n5280_), .ZN(new_n5281_));
  NOR2_X1    g05211(.A1(new_n5281_), .A2(new_n5238_), .ZN(new_n5282_));
  AND2_X2    g05212(.A1(new_n5276_), .A2(new_n5280_), .Z(new_n5283_));
  AND2_X2    g05213(.A1(new_n5268_), .A2(new_n5273_), .Z(new_n5284_));
  NOR2_X1    g05214(.A1(new_n5268_), .A2(new_n5273_), .ZN(new_n5285_));
  XOR2_X1    g05215(.A1(new_n5267_), .A2(new_n5243_), .Z(new_n5286_));
  NOR2_X1    g05216(.A1(new_n5285_), .A2(new_n5286_), .ZN(new_n5287_));
  NOR2_X1    g05217(.A1(new_n5287_), .A2(new_n5284_), .ZN(new_n5288_));
  AOI21_X1   g05218(.A1(new_n5242_), .A2(new_n5266_), .B(new_n5245_), .ZN(new_n5289_));
  NOR2_X1    g05219(.A1(new_n5242_), .A2(new_n5266_), .ZN(new_n5290_));
  NOR2_X1    g05220(.A1(new_n5289_), .A2(new_n5290_), .ZN(new_n5291_));
  INV_X1     g05221(.I(new_n5258_), .ZN(new_n5292_));
  AOI21_X1   g05222(.A1(new_n5292_), .A2(new_n5170_), .B(new_n5261_), .ZN(new_n5293_));
  INV_X1     g05223(.I(new_n5162_), .ZN(new_n5294_));
  NOR2_X1    g05224(.A1(new_n4331_), .A2(new_n88_), .ZN(new_n5295_));
  INV_X1     g05225(.I(new_n5295_), .ZN(new_n5296_));
  AOI22_X1   g05226(.A1(new_n4091_), .A2(new_n4406_), .B1(new_n962_), .B2(new_n4082_), .ZN(new_n5297_));
  AOI21_X1   g05227(.A1(new_n5297_), .A2(new_n5296_), .B(new_n82_), .ZN(new_n5298_));
  NAND2_X1   g05228(.A1(new_n5294_), .A2(new_n5298_), .ZN(new_n5299_));
  AOI22_X1   g05229(.A1(new_n4071_), .A2(new_n4570_), .B1(new_n4061_), .B2(new_n4526_), .ZN(new_n5300_));
  AOI21_X1   g05230(.A1(new_n101_), .A2(new_n4054_), .B(new_n5300_), .ZN(new_n5301_));
  OAI21_X1   g05231(.A1(new_n5301_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n5302_));
  XOR2_X1    g05232(.A1(new_n4652_), .A2(new_n5302_), .Z(new_n5303_));
  XOR2_X1    g05233(.A1(new_n5303_), .A2(new_n5299_), .Z(new_n5304_));
  NOR2_X1    g05234(.A1(new_n5304_), .A2(new_n5293_), .ZN(new_n5305_));
  INV_X1     g05235(.I(new_n5293_), .ZN(new_n5306_));
  INV_X1     g05236(.I(new_n5299_), .ZN(new_n5307_));
  AND2_X2    g05237(.A1(new_n5303_), .A2(new_n5307_), .Z(new_n5308_));
  NOR2_X1    g05238(.A1(new_n5303_), .A2(new_n5307_), .ZN(new_n5309_));
  NOR2_X1    g05239(.A1(new_n5308_), .A2(new_n5309_), .ZN(new_n5310_));
  NOR2_X1    g05240(.A1(new_n5310_), .A2(new_n5306_), .ZN(new_n5311_));
  NOR2_X1    g05241(.A1(new_n5311_), .A2(new_n5305_), .ZN(new_n5312_));
  AOI22_X1   g05242(.A1(new_n4043_), .A2(new_n4613_), .B1(new_n4036_), .B2(new_n4767_), .ZN(new_n5313_));
  AOI21_X1   g05243(.A1(new_n117_), .A2(new_n4029_), .B(new_n5313_), .ZN(new_n5314_));
  OAI21_X1   g05244(.A1(new_n5314_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n5315_));
  XOR2_X1    g05245(.A1(new_n4687_), .A2(new_n5315_), .Z(new_n5316_));
  INV_X1     g05246(.I(new_n5316_), .ZN(new_n5317_));
  NOR2_X1    g05247(.A1(new_n5317_), .A2(new_n5312_), .ZN(new_n5318_));
  NOR3_X1    g05248(.A1(new_n5316_), .A2(new_n5305_), .A3(new_n5311_), .ZN(new_n5319_));
  NOR2_X1    g05249(.A1(new_n5318_), .A2(new_n5319_), .ZN(new_n5320_));
  XNOR2_X1   g05250(.A1(new_n5316_), .A2(new_n5312_), .ZN(new_n5321_));
  NAND2_X1   g05251(.A1(new_n5321_), .A2(new_n5291_), .ZN(new_n5322_));
  OAI21_X1   g05252(.A1(new_n5291_), .A2(new_n5320_), .B(new_n5322_), .ZN(new_n5323_));
  OAI22_X1   g05253(.A1(new_n4444_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4397_), .ZN(new_n5324_));
  AOI21_X1   g05254(.A1(new_n5324_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n5325_));
  XNOR2_X1   g05255(.A1(new_n4403_), .A2(new_n5325_), .ZN(new_n5326_));
  INV_X1     g05256(.I(new_n5326_), .ZN(new_n5327_));
  NOR2_X1    g05257(.A1(new_n5323_), .A2(new_n5327_), .ZN(new_n5328_));
  NAND2_X1   g05258(.A1(new_n5323_), .A2(new_n5327_), .ZN(new_n5329_));
  INV_X1     g05259(.I(new_n5329_), .ZN(new_n5330_));
  NOR2_X1    g05260(.A1(new_n5330_), .A2(new_n5328_), .ZN(new_n5331_));
  XOR2_X1    g05261(.A1(new_n5323_), .A2(new_n5327_), .Z(new_n5332_));
  NAND2_X1   g05262(.A1(new_n5332_), .A2(new_n5288_), .ZN(new_n5333_));
  OAI21_X1   g05263(.A1(new_n5288_), .A2(new_n5331_), .B(new_n5333_), .ZN(new_n5334_));
  INV_X1     g05264(.I(new_n4722_), .ZN(new_n5335_));
  NOR2_X1    g05265(.A1(new_n5335_), .A2(new_n4719_), .ZN(new_n5336_));
  INV_X1     g05266(.I(new_n5336_), .ZN(new_n5337_));
  AOI22_X1   g05267(.A1(new_n4473_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4555_), .ZN(new_n5338_));
  OAI21_X1   g05268(.A1(new_n5338_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n5339_));
  XNOR2_X1   g05269(.A1(new_n4584_), .A2(new_n5339_), .ZN(new_n5340_));
  INV_X1     g05270(.I(new_n5340_), .ZN(new_n5341_));
  NOR2_X1    g05271(.A1(new_n5341_), .A2(new_n5334_), .ZN(new_n5342_));
  NAND2_X1   g05272(.A1(new_n5341_), .A2(new_n5334_), .ZN(new_n5343_));
  INV_X1     g05273(.I(new_n5343_), .ZN(new_n5344_));
  OAI22_X1   g05274(.A1(new_n5344_), .A2(new_n5342_), .B1(new_n5282_), .B2(new_n5283_), .ZN(new_n5345_));
  NOR2_X1    g05275(.A1(new_n5282_), .A2(new_n5283_), .ZN(new_n5346_));
  XNOR2_X1   g05276(.A1(new_n5334_), .A2(new_n5340_), .ZN(new_n5347_));
  NAND2_X1   g05277(.A1(new_n5347_), .A2(new_n5346_), .ZN(new_n5348_));
  NAND2_X1   g05278(.A1(new_n5348_), .A2(new_n5345_), .ZN(new_n5349_));
  INV_X1     g05279(.I(new_n5349_), .ZN(new_n5350_));
  OAI21_X1   g05280(.A1(new_n5235_), .A2(new_n5237_), .B(new_n5185_), .ZN(new_n5351_));
  XNOR2_X1   g05281(.A1(new_n5233_), .A2(new_n5228_), .ZN(new_n5352_));
  OAI21_X1   g05282(.A1(new_n5352_), .A2(new_n5185_), .B(new_n5351_), .ZN(new_n5353_));
  INV_X1     g05283(.I(new_n5148_), .ZN(new_n5354_));
  OAI21_X1   g05284(.A1(new_n5181_), .A2(new_n5183_), .B(new_n5354_), .ZN(new_n5355_));
  XOR2_X1    g05285(.A1(new_n5179_), .A2(new_n5175_), .Z(new_n5356_));
  OAI21_X1   g05286(.A1(new_n5356_), .A2(new_n5354_), .B(new_n5355_), .ZN(new_n5357_));
  OAI22_X1   g05287(.A1(new_n4331_), .A2(new_n4612_), .B1(new_n4081_), .B2(new_n4781_), .ZN(new_n5358_));
  OAI21_X1   g05288(.A1(new_n4070_), .A2(new_n1128_), .B(new_n5358_), .ZN(new_n5359_));
  AOI21_X1   g05289(.A1(new_n5359_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n5360_));
  XOR2_X1    g05290(.A1(new_n4927_), .A2(new_n5360_), .Z(new_n5361_));
  OAI22_X1   g05291(.A1(new_n4315_), .A2(new_n4529_), .B1(new_n4099_), .B2(new_n4527_), .ZN(new_n5362_));
  OAI21_X1   g05292(.A1(new_n4090_), .A2(new_n79_), .B(new_n5362_), .ZN(new_n5363_));
  AOI21_X1   g05293(.A1(new_n5363_), .A2(new_n72_), .B(new_n79_), .ZN(new_n5364_));
  XOR2_X1    g05294(.A1(new_n5196_), .A2(new_n5364_), .Z(new_n5365_));
  NOR2_X1    g05295(.A1(new_n5361_), .A2(new_n5365_), .ZN(new_n5366_));
  INV_X1     g05296(.I(new_n5366_), .ZN(new_n5367_));
  INV_X1     g05297(.I(new_n5361_), .ZN(new_n5368_));
  INV_X1     g05298(.I(new_n5365_), .ZN(new_n5369_));
  XNOR2_X1   g05299(.A1(new_n5102_), .A2(new_n5089_), .ZN(new_n5370_));
  INV_X1     g05300(.I(new_n5370_), .ZN(new_n5371_));
  NOR2_X1    g05301(.A1(new_n5104_), .A2(new_n5106_), .ZN(new_n5372_));
  NOR2_X1    g05302(.A1(new_n5088_), .A2(new_n5372_), .ZN(new_n5373_));
  AOI21_X1   g05303(.A1(new_n5088_), .A2(new_n5371_), .B(new_n5373_), .ZN(new_n5374_));
  OAI21_X1   g05304(.A1(new_n5368_), .A2(new_n5369_), .B(new_n5374_), .ZN(new_n5375_));
  NAND2_X1   g05305(.A1(new_n5375_), .A2(new_n5367_), .ZN(new_n5376_));
  INV_X1     g05306(.I(new_n5376_), .ZN(new_n5377_));
  AOI22_X1   g05307(.A1(new_n4071_), .A2(new_n4767_), .B1(new_n4082_), .B2(new_n4613_), .ZN(new_n5378_));
  AOI21_X1   g05308(.A1(new_n117_), .A2(new_n4061_), .B(new_n5378_), .ZN(new_n5379_));
  OAI21_X1   g05309(.A1(new_n5379_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n5380_));
  XOR2_X1    g05310(.A1(new_n4935_), .A2(new_n5380_), .Z(new_n5381_));
  NOR2_X1    g05311(.A1(new_n5377_), .A2(new_n5381_), .ZN(new_n5382_));
  XOR2_X1    g05312(.A1(new_n5143_), .A2(new_n5134_), .Z(new_n5383_));
  NOR2_X1    g05313(.A1(new_n5145_), .A2(new_n5147_), .ZN(new_n5384_));
  MUX2_X1    g05314(.I0(new_n5383_), .I1(new_n5384_), .S(new_n5107_), .Z(new_n5385_));
  NAND2_X1   g05315(.A1(new_n5377_), .A2(new_n5381_), .ZN(new_n5386_));
  AOI21_X1   g05316(.A1(new_n5385_), .A2(new_n5386_), .B(new_n5382_), .ZN(new_n5387_));
  INV_X1     g05317(.I(new_n5387_), .ZN(new_n5388_));
  OAI22_X1   g05318(.A1(new_n4349_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4028_), .ZN(new_n5389_));
  AOI21_X1   g05319(.A1(new_n5389_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n5390_));
  XNOR2_X1   g05320(.A1(new_n4687_), .A2(new_n5390_), .ZN(new_n5391_));
  INV_X1     g05321(.I(new_n5391_), .ZN(new_n5392_));
  NOR2_X1    g05322(.A1(new_n5392_), .A2(new_n5388_), .ZN(new_n5393_));
  INV_X1     g05323(.I(new_n5393_), .ZN(new_n5394_));
  NOR2_X1    g05324(.A1(new_n5391_), .A2(new_n5387_), .ZN(new_n5395_));
  AOI21_X1   g05325(.A1(new_n5394_), .A2(new_n5357_), .B(new_n5395_), .ZN(new_n5396_));
  INV_X1     g05326(.I(new_n5396_), .ZN(new_n5397_));
  INV_X1     g05327(.I(new_n4717_), .ZN(new_n5398_));
  OAI22_X1   g05328(.A1(new_n4397_), .A2(new_n5335_), .B1(new_n4374_), .B2(new_n4719_), .ZN(new_n5399_));
  OAI21_X1   g05329(.A1(new_n4437_), .A2(new_n5398_), .B(new_n5399_), .ZN(new_n5400_));
  AOI21_X1   g05330(.A1(new_n5400_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n5401_));
  XOR2_X1    g05331(.A1(new_n4541_), .A2(new_n5401_), .Z(new_n5402_));
  INV_X1     g05332(.I(new_n5402_), .ZN(new_n5403_));
  NOR2_X1    g05333(.A1(new_n5403_), .A2(new_n5397_), .ZN(new_n5404_));
  INV_X1     g05334(.I(new_n5404_), .ZN(new_n5405_));
  NOR2_X1    g05335(.A1(new_n5402_), .A2(new_n5396_), .ZN(new_n5406_));
  AOI21_X1   g05336(.A1(new_n5405_), .A2(new_n5353_), .B(new_n5406_), .ZN(new_n5407_));
  AOI22_X1   g05337(.A1(new_n4448_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4469_), .ZN(new_n5408_));
  OAI21_X1   g05338(.A1(new_n5408_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n5409_));
  XNOR2_X1   g05339(.A1(new_n4477_), .A2(new_n5409_), .ZN(new_n5410_));
  INV_X1     g05340(.I(new_n5238_), .ZN(new_n5411_));
  XOR2_X1    g05341(.A1(new_n5276_), .A2(new_n5280_), .Z(new_n5412_));
  NAND2_X1   g05342(.A1(new_n5412_), .A2(new_n5411_), .ZN(new_n5413_));
  OAI21_X1   g05343(.A1(new_n5283_), .A2(new_n5281_), .B(new_n5238_), .ZN(new_n5414_));
  NAND2_X1   g05344(.A1(new_n5407_), .A2(new_n5410_), .ZN(new_n5415_));
  NAND3_X1   g05345(.A1(new_n5413_), .A2(new_n5414_), .A3(new_n5415_), .ZN(new_n5416_));
  OAI21_X1   g05346(.A1(new_n5407_), .A2(new_n5410_), .B(new_n5416_), .ZN(new_n5417_));
  INV_X1     g05347(.I(new_n4567_), .ZN(new_n5418_));
  INV_X1     g05348(.I(new_n4663_), .ZN(new_n5419_));
  NOR2_X1    g05349(.A1(new_n5419_), .A2(new_n1622_), .ZN(new_n5420_));
  INV_X1     g05350(.I(new_n5420_), .ZN(new_n5421_));
  AOI22_X1   g05351(.A1(new_n5418_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4563_), .ZN(new_n5422_));
  OAI21_X1   g05352(.A1(new_n5422_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n5423_));
  XNOR2_X1   g05353(.A1(new_n4594_), .A2(new_n5423_), .ZN(new_n5424_));
  INV_X1     g05354(.I(new_n5424_), .ZN(new_n5425_));
  NOR2_X1    g05355(.A1(new_n5417_), .A2(new_n5425_), .ZN(new_n5426_));
  NAND2_X1   g05356(.A1(new_n5417_), .A2(new_n5425_), .ZN(new_n5427_));
  OAI21_X1   g05357(.A1(new_n5350_), .A2(new_n5426_), .B(new_n5427_), .ZN(new_n5428_));
  OAI21_X1   g05358(.A1(new_n5346_), .A2(new_n5342_), .B(new_n5343_), .ZN(new_n5429_));
  INV_X1     g05359(.I(new_n5429_), .ZN(new_n5430_));
  NOR2_X1    g05360(.A1(new_n5308_), .A2(new_n5293_), .ZN(new_n5431_));
  NOR2_X1    g05361(.A1(new_n5431_), .A2(new_n5309_), .ZN(new_n5432_));
  XOR2_X1    g05362(.A1(new_n4932_), .A2(new_n5299_), .Z(new_n5433_));
  NOR2_X1    g05363(.A1(new_n5432_), .A2(new_n5433_), .ZN(new_n5434_));
  NOR2_X1    g05364(.A1(new_n4932_), .A2(new_n5307_), .ZN(new_n5435_));
  NAND2_X1   g05365(.A1(new_n4932_), .A2(new_n5307_), .ZN(new_n5436_));
  INV_X1     g05366(.I(new_n5436_), .ZN(new_n5437_));
  NOR2_X1    g05367(.A1(new_n5437_), .A2(new_n5435_), .ZN(new_n5438_));
  INV_X1     g05368(.I(new_n5438_), .ZN(new_n5439_));
  AOI21_X1   g05369(.A1(new_n5432_), .A2(new_n5439_), .B(new_n5434_), .ZN(new_n5440_));
  INV_X1     g05370(.I(new_n5440_), .ZN(new_n5441_));
  OAI22_X1   g05371(.A1(new_n4017_), .A2(new_n1128_), .B1(new_n4352_), .B2(new_n4782_), .ZN(new_n5442_));
  AOI21_X1   g05372(.A1(new_n5442_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n5443_));
  XNOR2_X1   g05373(.A1(new_n4705_), .A2(new_n5443_), .ZN(new_n5444_));
  OAI22_X1   g05374(.A1(new_n4060_), .A2(new_n4529_), .B1(new_n4053_), .B2(new_n4527_), .ZN(new_n5445_));
  OAI21_X1   g05375(.A1(new_n4042_), .A2(new_n79_), .B(new_n5445_), .ZN(new_n5446_));
  AOI21_X1   g05376(.A1(new_n5446_), .A2(new_n72_), .B(new_n79_), .ZN(new_n5447_));
  XNOR2_X1   g05377(.A1(new_n4864_), .A2(new_n5447_), .ZN(new_n5448_));
  INV_X1     g05378(.I(new_n5448_), .ZN(new_n5449_));
  XOR2_X1    g05379(.A1(new_n5444_), .A2(new_n5449_), .Z(new_n5450_));
  INV_X1     g05380(.I(new_n5450_), .ZN(new_n5451_));
  AND2_X2    g05381(.A1(new_n5444_), .A2(new_n5448_), .Z(new_n5452_));
  NOR2_X1    g05382(.A1(new_n5444_), .A2(new_n5448_), .ZN(new_n5453_));
  NOR2_X1    g05383(.A1(new_n5452_), .A2(new_n5453_), .ZN(new_n5454_));
  NOR2_X1    g05384(.A1(new_n5454_), .A2(new_n5441_), .ZN(new_n5455_));
  AOI21_X1   g05385(.A1(new_n5441_), .A2(new_n5451_), .B(new_n5455_), .ZN(new_n5456_));
  NOR2_X1    g05386(.A1(new_n5318_), .A2(new_n5291_), .ZN(new_n5457_));
  NOR2_X1    g05387(.A1(new_n5457_), .A2(new_n5319_), .ZN(new_n5458_));
  OAI22_X1   g05388(.A1(new_n4397_), .A2(new_n4902_), .B1(new_n1973_), .B2(new_n4374_), .ZN(new_n5459_));
  OAI21_X1   g05389(.A1(new_n4437_), .A2(new_n1239_), .B(new_n5459_), .ZN(new_n5460_));
  AOI21_X1   g05390(.A1(new_n5460_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n5461_));
  XOR2_X1    g05391(.A1(new_n4541_), .A2(new_n5461_), .Z(new_n5462_));
  AND2_X2    g05392(.A1(new_n5462_), .A2(new_n5458_), .Z(new_n5463_));
  INV_X1     g05393(.I(new_n5463_), .ZN(new_n5464_));
  NOR2_X1    g05394(.A1(new_n5462_), .A2(new_n5458_), .ZN(new_n5465_));
  INV_X1     g05395(.I(new_n5465_), .ZN(new_n5466_));
  AOI21_X1   g05396(.A1(new_n5464_), .A2(new_n5466_), .B(new_n5456_), .ZN(new_n5467_));
  INV_X1     g05397(.I(new_n5456_), .ZN(new_n5468_));
  XNOR2_X1   g05398(.A1(new_n5462_), .A2(new_n5458_), .ZN(new_n5469_));
  NOR2_X1    g05399(.A1(new_n5468_), .A2(new_n5469_), .ZN(new_n5470_));
  NOR2_X1    g05400(.A1(new_n5470_), .A2(new_n5467_), .ZN(new_n5471_));
  OAI21_X1   g05401(.A1(new_n5288_), .A2(new_n5328_), .B(new_n5329_), .ZN(new_n5472_));
  OAI22_X1   g05402(.A1(new_n4468_), .A2(new_n4719_), .B1(new_n4501_), .B2(new_n5335_), .ZN(new_n5473_));
  OAI21_X1   g05403(.A1(new_n4516_), .A2(new_n5398_), .B(new_n5473_), .ZN(new_n5474_));
  AOI21_X1   g05404(.A1(new_n5474_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n5475_));
  XOR2_X1    g05405(.A1(new_n4524_), .A2(new_n5475_), .Z(new_n5476_));
  INV_X1     g05406(.I(new_n5476_), .ZN(new_n5477_));
  NOR2_X1    g05407(.A1(new_n5477_), .A2(new_n5472_), .ZN(new_n5478_));
  INV_X1     g05408(.I(new_n5478_), .ZN(new_n5479_));
  NAND2_X1   g05409(.A1(new_n5477_), .A2(new_n5472_), .ZN(new_n5480_));
  AOI21_X1   g05410(.A1(new_n5479_), .A2(new_n5480_), .B(new_n5471_), .ZN(new_n5481_));
  INV_X1     g05411(.I(new_n5471_), .ZN(new_n5482_));
  XOR2_X1    g05412(.A1(new_n5476_), .A2(new_n5472_), .Z(new_n5483_));
  NOR2_X1    g05413(.A1(new_n5482_), .A2(new_n5483_), .ZN(new_n5484_));
  NAND2_X1   g05414(.A1(new_n4563_), .A2(new_n4663_), .ZN(new_n5485_));
  NAND2_X1   g05415(.A1(new_n4564_), .A2(new_n4661_), .ZN(new_n5486_));
  AOI22_X1   g05416(.A1(new_n5486_), .A2(new_n5485_), .B1(new_n4660_), .B2(new_n4564_), .ZN(new_n5487_));
  OAI21_X1   g05417(.A1(new_n5487_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n5488_));
  XOR2_X1    g05418(.A1(new_n4609_), .A2(new_n5488_), .Z(new_n5489_));
  INV_X1     g05419(.I(new_n5489_), .ZN(new_n5490_));
  NOR3_X1    g05420(.A1(new_n5481_), .A2(new_n5484_), .A3(new_n5490_), .ZN(new_n5491_));
  NOR2_X1    g05421(.A1(new_n5481_), .A2(new_n5484_), .ZN(new_n5492_));
  NOR2_X1    g05422(.A1(new_n5492_), .A2(new_n5489_), .ZN(new_n5493_));
  NOR2_X1    g05423(.A1(new_n5493_), .A2(new_n5491_), .ZN(new_n5494_));
  NOR2_X1    g05424(.A1(new_n5494_), .A2(new_n5430_), .ZN(new_n5495_));
  XOR2_X1    g05425(.A1(new_n5492_), .A2(new_n5490_), .Z(new_n5496_));
  NOR2_X1    g05426(.A1(new_n5496_), .A2(new_n5429_), .ZN(new_n5497_));
  NOR2_X1    g05427(.A1(new_n5497_), .A2(new_n5495_), .ZN(new_n5498_));
  INV_X1     g05428(.I(new_n5498_), .ZN(new_n5499_));
  NOR2_X1    g05429(.A1(new_n5499_), .A2(new_n644_), .ZN(new_n5500_));
  INV_X1     g05430(.I(new_n5500_), .ZN(new_n5501_));
  NOR2_X1    g05431(.A1(new_n5498_), .A2(new_n786_), .ZN(new_n5502_));
  AOI21_X1   g05432(.A1(new_n5501_), .A2(new_n5428_), .B(new_n5502_), .ZN(new_n5503_));
  INV_X1     g05433(.I(new_n5491_), .ZN(new_n5504_));
  AOI21_X1   g05434(.A1(new_n5504_), .A2(new_n5429_), .B(new_n5493_), .ZN(new_n5505_));
  OAI21_X1   g05435(.A1(new_n5432_), .A2(new_n5435_), .B(new_n5436_), .ZN(new_n5506_));
  INV_X1     g05436(.I(new_n5506_), .ZN(new_n5507_));
  XNOR2_X1   g05437(.A1(new_n4939_), .A2(new_n4932_), .ZN(new_n5508_));
  NOR2_X1    g05438(.A1(new_n5508_), .A2(new_n4948_), .ZN(new_n5509_));
  INV_X1     g05439(.I(new_n4940_), .ZN(new_n5510_));
  INV_X1     g05440(.I(new_n4948_), .ZN(new_n5511_));
  AOI21_X1   g05441(.A1(new_n5510_), .A2(new_n4949_), .B(new_n5511_), .ZN(new_n5512_));
  NOR2_X1    g05442(.A1(new_n5509_), .A2(new_n5512_), .ZN(new_n5513_));
  INV_X1     g05443(.I(new_n5513_), .ZN(new_n5514_));
  AOI22_X1   g05444(.A1(new_n4043_), .A2(new_n4526_), .B1(new_n4054_), .B2(new_n4570_), .ZN(new_n5515_));
  AOI21_X1   g05445(.A1(new_n101_), .A2(new_n4036_), .B(new_n5515_), .ZN(new_n5516_));
  OAI21_X1   g05446(.A1(new_n5516_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n5517_));
  XOR2_X1    g05447(.A1(new_n4672_), .A2(new_n5517_), .Z(new_n5518_));
  XOR2_X1    g05448(.A1(new_n5518_), .A2(new_n5514_), .Z(new_n5519_));
  NOR2_X1    g05449(.A1(new_n5519_), .A2(new_n5507_), .ZN(new_n5520_));
  AND2_X2    g05450(.A1(new_n5518_), .A2(new_n5513_), .Z(new_n5521_));
  NOR2_X1    g05451(.A1(new_n5518_), .A2(new_n5513_), .ZN(new_n5522_));
  NOR2_X1    g05452(.A1(new_n5521_), .A2(new_n5522_), .ZN(new_n5523_));
  NOR2_X1    g05453(.A1(new_n5523_), .A2(new_n5506_), .ZN(new_n5524_));
  NOR2_X1    g05454(.A1(new_n5524_), .A2(new_n5520_), .ZN(new_n5525_));
  NOR2_X1    g05455(.A1(new_n5452_), .A2(new_n5441_), .ZN(new_n5526_));
  AOI22_X1   g05456(.A1(new_n4018_), .A2(new_n4767_), .B1(new_n4029_), .B2(new_n4613_), .ZN(new_n5527_));
  AOI21_X1   g05457(.A1(new_n117_), .A2(new_n4375_), .B(new_n5527_), .ZN(new_n5528_));
  OAI21_X1   g05458(.A1(new_n5528_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n5529_));
  XOR2_X1    g05459(.A1(new_n4730_), .A2(new_n5529_), .Z(new_n5530_));
  INV_X1     g05460(.I(new_n5530_), .ZN(new_n5531_));
  NOR3_X1    g05461(.A1(new_n5526_), .A2(new_n5453_), .A3(new_n5531_), .ZN(new_n5532_));
  NOR2_X1    g05462(.A1(new_n5526_), .A2(new_n5453_), .ZN(new_n5533_));
  NOR2_X1    g05463(.A1(new_n5533_), .A2(new_n5530_), .ZN(new_n5534_));
  NOR2_X1    g05464(.A1(new_n5534_), .A2(new_n5532_), .ZN(new_n5535_));
  NOR2_X1    g05465(.A1(new_n5535_), .A2(new_n5525_), .ZN(new_n5536_));
  XOR2_X1    g05466(.A1(new_n5533_), .A2(new_n5531_), .Z(new_n5537_));
  NOR3_X1    g05467(.A1(new_n5537_), .A2(new_n5520_), .A3(new_n5524_), .ZN(new_n5538_));
  NOR2_X1    g05468(.A1(new_n5538_), .A2(new_n5536_), .ZN(new_n5539_));
  INV_X1     g05469(.I(new_n5539_), .ZN(new_n5540_));
  OAI21_X1   g05470(.A1(new_n5456_), .A2(new_n5463_), .B(new_n5466_), .ZN(new_n5541_));
  OAI22_X1   g05471(.A1(new_n4447_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4468_), .ZN(new_n5542_));
  AOI21_X1   g05472(.A1(new_n5542_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n5543_));
  XOR2_X1    g05473(.A1(new_n4477_), .A2(new_n5543_), .Z(new_n5544_));
  INV_X1     g05474(.I(new_n5544_), .ZN(new_n5545_));
  XOR2_X1    g05475(.A1(new_n5541_), .A2(new_n5545_), .Z(new_n5546_));
  INV_X1     g05476(.I(new_n5546_), .ZN(new_n5547_));
  XOR2_X1    g05477(.A1(new_n5541_), .A2(new_n5544_), .Z(new_n5548_));
  NOR2_X1    g05478(.A1(new_n5540_), .A2(new_n5548_), .ZN(new_n5549_));
  AOI21_X1   g05479(.A1(new_n5540_), .A2(new_n5547_), .B(new_n5549_), .ZN(new_n5550_));
  OAI21_X1   g05480(.A1(new_n5471_), .A2(new_n5478_), .B(new_n5480_), .ZN(new_n5551_));
  NOR2_X1    g05481(.A1(new_n4516_), .A2(new_n4501_), .ZN(new_n5552_));
  INV_X1     g05482(.I(new_n5552_), .ZN(new_n5553_));
  AOI22_X1   g05483(.A1(new_n5553_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4564_), .ZN(new_n5554_));
  OAI21_X1   g05484(.A1(new_n5554_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n5555_));
  XOR2_X1    g05485(.A1(new_n4569_), .A2(new_n5555_), .Z(new_n5556_));
  INV_X1     g05486(.I(new_n5556_), .ZN(new_n5557_));
  NOR2_X1    g05487(.A1(new_n5557_), .A2(new_n5551_), .ZN(new_n5558_));
  INV_X1     g05488(.I(new_n5558_), .ZN(new_n5559_));
  NAND2_X1   g05489(.A1(new_n5557_), .A2(new_n5551_), .ZN(new_n5560_));
  AOI21_X1   g05490(.A1(new_n5559_), .A2(new_n5560_), .B(new_n5550_), .ZN(new_n5561_));
  INV_X1     g05491(.I(new_n5550_), .ZN(new_n5562_));
  XOR2_X1    g05492(.A1(new_n5551_), .A2(new_n5556_), .Z(new_n5563_));
  NOR2_X1    g05493(.A1(new_n5562_), .A2(new_n5563_), .ZN(new_n5564_));
  NOR2_X1    g05494(.A1(new_n5564_), .A2(new_n5561_), .ZN(new_n5565_));
  NAND2_X1   g05495(.A1(new_n4663_), .A2(new_n4660_), .ZN(new_n5566_));
  OAI21_X1   g05496(.A1(new_n4661_), .A2(new_n5566_), .B(new_n4564_), .ZN(new_n5567_));
  OAI21_X1   g05497(.A1(new_n5567_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n5568_));
  XOR2_X1    g05498(.A1(new_n5001_), .A2(new_n5568_), .Z(new_n5569_));
  XOR2_X1    g05499(.A1(new_n5565_), .A2(new_n5569_), .Z(new_n5570_));
  NOR2_X1    g05500(.A1(new_n5570_), .A2(new_n5505_), .ZN(new_n5571_));
  INV_X1     g05501(.I(new_n5569_), .ZN(new_n5572_));
  NOR2_X1    g05502(.A1(new_n5565_), .A2(new_n5572_), .ZN(new_n5573_));
  INV_X1     g05503(.I(new_n5573_), .ZN(new_n5574_));
  NAND2_X1   g05504(.A1(new_n5565_), .A2(new_n5572_), .ZN(new_n5575_));
  NAND2_X1   g05505(.A1(new_n5574_), .A2(new_n5575_), .ZN(new_n5576_));
  AOI21_X1   g05506(.A1(new_n5505_), .A2(new_n5576_), .B(new_n5571_), .ZN(new_n5577_));
  NOR2_X1    g05507(.A1(new_n5577_), .A2(new_n5503_), .ZN(new_n5578_));
  INV_X1     g05508(.I(new_n5578_), .ZN(new_n5579_));
  NOR2_X1    g05509(.A1(new_n5393_), .A2(new_n5395_), .ZN(new_n5580_));
  XOR2_X1    g05510(.A1(new_n5391_), .A2(new_n5388_), .Z(new_n5581_));
  MUX2_X1    g05511(.I0(new_n5581_), .I1(new_n5580_), .S(new_n5357_), .Z(new_n5582_));
  XOR2_X1    g05512(.A1(new_n5361_), .A2(new_n5369_), .Z(new_n5583_));
  NOR2_X1    g05513(.A1(new_n5583_), .A2(new_n5374_), .ZN(new_n5584_));
  NOR2_X1    g05514(.A1(new_n5368_), .A2(new_n5369_), .ZN(new_n5585_));
  NOR2_X1    g05515(.A1(new_n5585_), .A2(new_n5366_), .ZN(new_n5586_));
  INV_X1     g05516(.I(new_n5586_), .ZN(new_n5587_));
  AOI21_X1   g05517(.A1(new_n5374_), .A2(new_n5587_), .B(new_n5584_), .ZN(new_n5588_));
  XOR2_X1    g05518(.A1(new_n5054_), .A2(new_n5040_), .Z(new_n5589_));
  OAI21_X1   g05519(.A1(new_n5056_), .A2(new_n5058_), .B(new_n5029_), .ZN(new_n5590_));
  OAI21_X1   g05520(.A1(new_n5029_), .A2(new_n5589_), .B(new_n5590_), .ZN(new_n5591_));
  NAND2_X1   g05521(.A1(new_n5027_), .A2(new_n5030_), .ZN(new_n5592_));
  XNOR2_X1   g05522(.A1(new_n4296_), .A2(new_n4285_), .ZN(new_n5593_));
  XOR2_X1    g05523(.A1(new_n4131_), .A2(new_n4297_), .Z(new_n5594_));
  NOR3_X1    g05524(.A1(new_n5594_), .A2(new_n4300_), .A3(new_n5593_), .ZN(new_n5595_));
  INV_X1     g05525(.I(new_n5593_), .ZN(new_n5596_));
  XOR2_X1    g05526(.A1(new_n4131_), .A2(new_n4296_), .Z(new_n5597_));
  AOI21_X1   g05527(.A1(new_n5597_), .A2(new_n5596_), .B(new_n4289_), .ZN(new_n5598_));
  OR2_X2     g05528(.A1(new_n5595_), .A2(new_n5598_), .Z(new_n5599_));
  NAND2_X1   g05529(.A1(new_n5042_), .A2(new_n962_), .ZN(new_n5600_));
  AOI22_X1   g05530(.A1(new_n4297_), .A2(new_n87_), .B1(new_n4290_), .B2(new_n4406_), .ZN(new_n5601_));
  AOI21_X1   g05531(.A1(new_n5600_), .A2(new_n5601_), .B(new_n82_), .ZN(new_n5602_));
  NAND2_X1   g05532(.A1(new_n5599_), .A2(new_n5602_), .ZN(new_n5603_));
  NAND2_X1   g05533(.A1(new_n5603_), .A2(new_n5592_), .ZN(new_n5604_));
  INV_X1     g05534(.I(new_n5604_), .ZN(new_n5605_));
  AOI22_X1   g05535(.A1(new_n4113_), .A2(new_n4526_), .B1(new_n4124_), .B2(new_n4570_), .ZN(new_n5606_));
  AOI21_X1   g05536(.A1(new_n101_), .A2(new_n4105_), .B(new_n5606_), .ZN(new_n5607_));
  OAI21_X1   g05537(.A1(new_n5607_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n5608_));
  XOR2_X1    g05538(.A1(new_n5121_), .A2(new_n5608_), .Z(new_n5609_));
  INV_X1     g05539(.I(new_n5609_), .ZN(new_n5610_));
  INV_X1     g05540(.I(new_n5591_), .ZN(new_n5611_));
  NOR2_X1    g05541(.A1(new_n5603_), .A2(new_n5592_), .ZN(new_n5612_));
  NOR2_X1    g05542(.A1(new_n5605_), .A2(new_n5612_), .ZN(new_n5613_));
  NAND2_X1   g05543(.A1(new_n5027_), .A2(new_n5030_), .ZN(new_n5614_));
  XOR2_X1    g05544(.A1(new_n5027_), .A2(new_n5030_), .Z(new_n5615_));
  INV_X1     g05545(.I(new_n5615_), .ZN(new_n5616_));
  INV_X1     g05546(.I(new_n4287_), .ZN(new_n5617_));
  AOI21_X1   g05547(.A1(new_n5617_), .A2(new_n4286_), .B(new_n4135_), .ZN(new_n5618_));
  INV_X1     g05548(.I(new_n5618_), .ZN(new_n5619_));
  NAND2_X1   g05549(.A1(new_n4280_), .A2(new_n4142_), .ZN(new_n5620_));
  NAND2_X1   g05550(.A1(new_n4279_), .A2(new_n4143_), .ZN(new_n5621_));
  AOI21_X1   g05551(.A1(new_n5620_), .A2(new_n5621_), .B(new_n4136_), .ZN(new_n5622_));
  INV_X1     g05552(.I(new_n5622_), .ZN(new_n5623_));
  NAND2_X1   g05553(.A1(new_n5619_), .A2(new_n5623_), .ZN(new_n5624_));
  AOI22_X1   g05554(.A1(new_n4143_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n4274_), .ZN(new_n5625_));
  OAI21_X1   g05555(.A1(new_n4135_), .A2(new_n511_), .B(new_n5625_), .ZN(new_n5626_));
  NOR2_X1    g05556(.A1(new_n4244_), .A2(new_n4230_), .ZN(new_n5627_));
  OAI22_X1   g05557(.A1(new_n4244_), .A2(new_n88_), .B1(new_n92_), .B2(new_n4230_), .ZN(new_n5628_));
  OAI21_X1   g05558(.A1(new_n511_), .A2(new_n4234_), .B(new_n5628_), .ZN(new_n5629_));
  OAI21_X1   g05559(.A1(new_n5629_), .A2(new_n5627_), .B(new_n4234_), .ZN(new_n5630_));
  AOI21_X1   g05560(.A1(new_n5627_), .A2(new_n5629_), .B(new_n5630_), .ZN(new_n5631_));
  NOR2_X1    g05561(.A1(new_n5631_), .A2(new_n82_), .ZN(new_n5632_));
  NAND2_X1   g05562(.A1(new_n4251_), .A2(new_n962_), .ZN(new_n5633_));
  NAND2_X1   g05563(.A1(new_n4252_), .A2(new_n4406_), .ZN(new_n5634_));
  NOR2_X1    g05564(.A1(new_n4230_), .A2(new_n4252_), .ZN(new_n5635_));
  NOR2_X1    g05565(.A1(new_n4244_), .A2(new_n4251_), .ZN(new_n5636_));
  NOR2_X1    g05566(.A1(new_n5636_), .A2(new_n5635_), .ZN(new_n5637_));
  AOI22_X1   g05567(.A1(new_n5637_), .A2(new_n961_), .B1(new_n5633_), .B2(new_n5634_), .ZN(new_n5638_));
  NAND2_X1   g05568(.A1(new_n5632_), .A2(new_n5638_), .ZN(new_n5639_));
  AOI21_X1   g05569(.A1(new_n4213_), .A2(new_n4220_), .B(new_n4251_), .ZN(new_n5640_));
  INV_X1     g05570(.I(new_n5640_), .ZN(new_n5641_));
  NAND3_X1   g05571(.A1(new_n4213_), .A2(new_n4220_), .A3(new_n4251_), .ZN(new_n5642_));
  NAND2_X1   g05572(.A1(new_n4249_), .A2(new_n4234_), .ZN(new_n5643_));
  NAND4_X1   g05573(.A1(new_n5643_), .A2(new_n5641_), .A3(new_n5642_), .A4(new_n4244_), .ZN(new_n5644_));
  INV_X1     g05574(.I(new_n5642_), .ZN(new_n5645_));
  NOR2_X1    g05575(.A1(new_n4221_), .A2(new_n4260_), .ZN(new_n5646_));
  OAI22_X1   g05576(.A1(new_n4252_), .A2(new_n5646_), .B1(new_n5645_), .B2(new_n5640_), .ZN(new_n5647_));
  NAND2_X1   g05577(.A1(new_n5647_), .A2(new_n5644_), .ZN(new_n5648_));
  AOI22_X1   g05578(.A1(new_n4221_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n4252_), .ZN(new_n5649_));
  OAI21_X1   g05579(.A1(new_n88_), .A2(new_n4234_), .B(new_n5649_), .ZN(new_n5650_));
  NAND3_X1   g05580(.A1(new_n5648_), .A2(new_n961_), .A3(new_n5650_), .ZN(new_n5651_));
  NOR2_X1    g05581(.A1(new_n5639_), .A2(new_n5651_), .ZN(new_n5652_));
  OAI21_X1   g05582(.A1(new_n4200_), .A2(new_n4201_), .B(new_n3700_), .ZN(new_n5653_));
  NAND3_X1   g05583(.A1(new_n4198_), .A2(new_n4194_), .A3(new_n4176_), .ZN(new_n5654_));
  NAND2_X1   g05584(.A1(new_n5653_), .A2(new_n5654_), .ZN(new_n5655_));
  OAI21_X1   g05585(.A1(new_n4256_), .A2(new_n4245_), .B(new_n5655_), .ZN(new_n5656_));
  AOI21_X1   g05586(.A1(new_n4251_), .A2(new_n4260_), .B(new_n4221_), .ZN(new_n5657_));
  AOI21_X1   g05587(.A1(new_n4263_), .A2(new_n4230_), .B(new_n4249_), .ZN(new_n5658_));
  OAI21_X1   g05588(.A1(new_n5658_), .A2(new_n5657_), .B(new_n4203_), .ZN(new_n5659_));
  NAND2_X1   g05589(.A1(new_n5659_), .A2(new_n5656_), .ZN(new_n5660_));
  NAND2_X1   g05590(.A1(new_n5655_), .A2(new_n962_), .ZN(new_n5661_));
  AOI22_X1   g05591(.A1(new_n4221_), .A2(new_n87_), .B1(new_n4260_), .B2(new_n4406_), .ZN(new_n5662_));
  AOI21_X1   g05592(.A1(new_n5661_), .A2(new_n5662_), .B(new_n82_), .ZN(new_n5663_));
  NAND3_X1   g05593(.A1(new_n5652_), .A2(new_n5660_), .A3(new_n5663_), .ZN(new_n5664_));
  NAND2_X1   g05594(.A1(new_n5655_), .A2(new_n4245_), .ZN(new_n5665_));
  AOI21_X1   g05595(.A1(new_n4264_), .A2(new_n5665_), .B(new_n4175_), .ZN(new_n5666_));
  INV_X1     g05596(.I(new_n5666_), .ZN(new_n5667_));
  AOI21_X1   g05597(.A1(new_n4256_), .A2(new_n4246_), .B(new_n5655_), .ZN(new_n5668_));
  NOR2_X1    g05598(.A1(new_n4203_), .A2(new_n4245_), .ZN(new_n5669_));
  OAI21_X1   g05599(.A1(new_n5668_), .A2(new_n5669_), .B(new_n4175_), .ZN(new_n5670_));
  NAND2_X1   g05600(.A1(new_n5670_), .A2(new_n5667_), .ZN(new_n5671_));
  NAND2_X1   g05601(.A1(new_n4258_), .A2(new_n962_), .ZN(new_n5672_));
  AOI22_X1   g05602(.A1(new_n5655_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n4221_), .ZN(new_n5673_));
  AOI21_X1   g05603(.A1(new_n5672_), .A2(new_n5673_), .B(new_n82_), .ZN(new_n5674_));
  NAND2_X1   g05604(.A1(new_n5671_), .A2(new_n5674_), .ZN(new_n5675_));
  NAND3_X1   g05605(.A1(new_n4263_), .A2(new_n4221_), .A3(new_n4230_), .ZN(new_n5676_));
  OAI21_X1   g05606(.A1(new_n5676_), .A2(new_n4245_), .B(new_n4203_), .ZN(new_n5677_));
  INV_X1     g05607(.I(new_n5669_), .ZN(new_n5678_));
  NAND2_X1   g05608(.A1(new_n5677_), .A2(new_n5678_), .ZN(new_n5679_));
  NAND2_X1   g05609(.A1(new_n5676_), .A2(new_n4203_), .ZN(new_n5680_));
  NAND3_X1   g05610(.A1(new_n5680_), .A2(new_n4171_), .A3(new_n4246_), .ZN(new_n5681_));
  AOI21_X1   g05611(.A1(new_n4167_), .A2(new_n4162_), .B(new_n3703_), .ZN(new_n5682_));
  INV_X1     g05612(.I(new_n4170_), .ZN(new_n5683_));
  NOR2_X1    g05613(.A1(new_n5683_), .A2(new_n5682_), .ZN(new_n5684_));
  NOR2_X1    g05614(.A1(new_n4256_), .A2(new_n5655_), .ZN(new_n5685_));
  OAI21_X1   g05615(.A1(new_n5685_), .A2(new_n4245_), .B(new_n5684_), .ZN(new_n5686_));
  NAND2_X1   g05616(.A1(new_n5686_), .A2(new_n5681_), .ZN(new_n5687_));
  NAND3_X1   g05617(.A1(new_n5687_), .A2(new_n4175_), .A3(new_n5679_), .ZN(new_n5688_));
  NOR3_X1    g05618(.A1(new_n5685_), .A2(new_n5684_), .A3(new_n4245_), .ZN(new_n5689_));
  AOI21_X1   g05619(.A1(new_n5680_), .A2(new_n4246_), .B(new_n4171_), .ZN(new_n5690_));
  OAI21_X1   g05620(.A1(new_n5690_), .A2(new_n5689_), .B(new_n5679_), .ZN(new_n5691_));
  NAND2_X1   g05621(.A1(new_n5691_), .A2(new_n4258_), .ZN(new_n5692_));
  NAND2_X1   g05622(.A1(new_n5692_), .A2(new_n5688_), .ZN(new_n5693_));
  NAND2_X1   g05623(.A1(new_n4258_), .A2(new_n87_), .ZN(new_n5694_));
  AOI22_X1   g05624(.A1(new_n4171_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n5655_), .ZN(new_n5695_));
  AOI21_X1   g05625(.A1(new_n5695_), .A2(new_n5694_), .B(new_n82_), .ZN(new_n5696_));
  NAND2_X1   g05626(.A1(new_n5693_), .A2(new_n5696_), .ZN(new_n5697_));
  NOR3_X1    g05627(.A1(new_n5697_), .A2(new_n5664_), .A3(new_n5675_), .ZN(new_n5698_));
  INV_X1     g05628(.I(new_n4257_), .ZN(new_n5699_));
  AOI21_X1   g05629(.A1(new_n5699_), .A2(new_n4268_), .B(new_n4150_), .ZN(new_n5700_));
  INV_X1     g05630(.I(new_n4150_), .ZN(new_n5701_));
  INV_X1     g05631(.I(new_n4265_), .ZN(new_n5702_));
  NAND2_X1   g05632(.A1(new_n5702_), .A2(new_n4171_), .ZN(new_n5703_));
  NAND3_X1   g05633(.A1(new_n5703_), .A2(new_n5684_), .A3(new_n4267_), .ZN(new_n5704_));
  OAI21_X1   g05634(.A1(new_n5702_), .A2(new_n4266_), .B(new_n4171_), .ZN(new_n5705_));
  AOI21_X1   g05635(.A1(new_n5704_), .A2(new_n5705_), .B(new_n5701_), .ZN(new_n5706_));
  NOR2_X1    g05636(.A1(new_n5706_), .A2(new_n5700_), .ZN(new_n5707_));
  NOR2_X1    g05637(.A1(new_n4150_), .A2(new_n511_), .ZN(new_n5708_));
  OAI22_X1   g05638(.A1(new_n5684_), .A2(new_n88_), .B1(new_n92_), .B2(new_n4175_), .ZN(new_n5709_));
  OAI21_X1   g05639(.A1(new_n5708_), .A2(new_n5709_), .B(new_n961_), .ZN(new_n5710_));
  NOR2_X1    g05640(.A1(new_n5707_), .A2(new_n5710_), .ZN(new_n5711_));
  NAND2_X1   g05641(.A1(new_n5698_), .A2(new_n5711_), .ZN(new_n5712_));
  NAND2_X1   g05642(.A1(new_n5701_), .A2(new_n4257_), .ZN(new_n5714_));
  AOI21_X1   g05643(.A1(new_n4275_), .A2(new_n5714_), .B(new_n4273_), .ZN(new_n5715_));
  INV_X1     g05644(.I(new_n5715_), .ZN(new_n5716_));
  NOR2_X1    g05645(.A1(new_n4269_), .A2(new_n5701_), .ZN(new_n5717_));
  NOR2_X1    g05646(.A1(new_n4150_), .A2(new_n4257_), .ZN(new_n5718_));
  NOR2_X1    g05647(.A1(new_n5717_), .A2(new_n5718_), .ZN(new_n5719_));
  NOR2_X1    g05648(.A1(new_n5719_), .A2(new_n4274_), .ZN(new_n5720_));
  INV_X1     g05649(.I(new_n5720_), .ZN(new_n5721_));
  NAND2_X1   g05650(.A1(new_n5721_), .A2(new_n5716_), .ZN(new_n5722_));
  NAND2_X1   g05651(.A1(new_n5701_), .A2(new_n87_), .ZN(new_n5723_));
  AOI22_X1   g05652(.A1(new_n4274_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n4171_), .ZN(new_n5724_));
  AOI21_X1   g05653(.A1(new_n5724_), .A2(new_n5723_), .B(new_n82_), .ZN(new_n5725_));
  NAND2_X1   g05654(.A1(new_n5722_), .A2(new_n5725_), .ZN(new_n5726_));
  NOR2_X1    g05655(.A1(new_n5726_), .A2(new_n5712_), .ZN(new_n5727_));
  INV_X1     g05656(.I(new_n5719_), .ZN(new_n5728_));
  XOR2_X1    g05657(.A1(new_n4142_), .A2(new_n4269_), .Z(new_n5729_));
  NAND3_X1   g05658(.A1(new_n5728_), .A2(new_n5729_), .A3(new_n4273_), .ZN(new_n5730_));
  XNOR2_X1   g05659(.A1(new_n4142_), .A2(new_n4269_), .ZN(new_n5731_));
  OAI21_X1   g05660(.A1(new_n5731_), .A2(new_n5719_), .B(new_n4274_), .ZN(new_n5732_));
  NAND2_X1   g05661(.A1(new_n5732_), .A2(new_n5730_), .ZN(new_n5733_));
  NOR2_X1    g05662(.A1(new_n4142_), .A2(new_n511_), .ZN(new_n5734_));
  INV_X1     g05663(.I(new_n5734_), .ZN(new_n5735_));
  AOI22_X1   g05664(.A1(new_n4274_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n5701_), .ZN(new_n5736_));
  AOI21_X1   g05665(.A1(new_n5735_), .A2(new_n5736_), .B(new_n82_), .ZN(new_n5737_));
  NAND2_X1   g05666(.A1(new_n5733_), .A2(new_n5737_), .ZN(new_n5738_));
  NOR2_X1    g05667(.A1(new_n5727_), .A2(new_n5738_), .ZN(new_n5739_));
  NAND4_X1   g05668(.A1(new_n5624_), .A2(new_n961_), .A3(new_n5626_), .A4(new_n5739_), .ZN(new_n5740_));
  OAI22_X1   g05669(.A1(new_n4131_), .A2(new_n4527_), .B1(new_n4296_), .B2(new_n4529_), .ZN(new_n5741_));
  OAI21_X1   g05670(.A1(new_n79_), .A2(new_n4309_), .B(new_n5741_), .ZN(new_n5742_));
  AOI21_X1   g05671(.A1(new_n5742_), .A2(new_n72_), .B(new_n79_), .ZN(new_n5743_));
  XNOR2_X1   g05672(.A1(new_n5049_), .A2(new_n5743_), .ZN(new_n5744_));
  NAND2_X1   g05673(.A1(new_n5744_), .A2(new_n5740_), .ZN(new_n5745_));
  NAND2_X1   g05674(.A1(new_n5745_), .A2(new_n5616_), .ZN(new_n5746_));
  OR2_X2     g05675(.A1(new_n5744_), .A2(new_n5740_), .Z(new_n5747_));
  NAND2_X1   g05676(.A1(new_n5746_), .A2(new_n5747_), .ZN(new_n5748_));
  INV_X1     g05677(.I(new_n5748_), .ZN(new_n5749_));
  NOR2_X1    g05678(.A1(new_n5593_), .A2(new_n4289_), .ZN(new_n5750_));
  INV_X1     g05679(.I(new_n5750_), .ZN(new_n5751_));
  NOR2_X1    g05680(.A1(new_n4298_), .A2(new_n4301_), .ZN(new_n5752_));
  OAI21_X1   g05681(.A1(new_n4300_), .A2(new_n5752_), .B(new_n5751_), .ZN(new_n5753_));
  NAND2_X1   g05682(.A1(new_n4290_), .A2(new_n87_), .ZN(new_n5754_));
  AOI22_X1   g05683(.A1(new_n4297_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n4136_), .ZN(new_n5755_));
  AOI21_X1   g05684(.A1(new_n5755_), .A2(new_n5754_), .B(new_n82_), .ZN(new_n5756_));
  NAND2_X1   g05685(.A1(new_n5753_), .A2(new_n5756_), .ZN(new_n5757_));
  AOI21_X1   g05686(.A1(new_n5749_), .A2(new_n5757_), .B(new_n5614_), .ZN(new_n5758_));
  NOR2_X1    g05687(.A1(new_n5749_), .A2(new_n5757_), .ZN(new_n5759_));
  NOR2_X1    g05688(.A1(new_n5758_), .A2(new_n5759_), .ZN(new_n5760_));
  NAND2_X1   g05689(.A1(new_n5760_), .A2(new_n5613_), .ZN(new_n5761_));
  AOI21_X1   g05690(.A1(new_n5611_), .A2(new_n5604_), .B(new_n5761_), .ZN(new_n5762_));
  AOI22_X1   g05691(.A1(new_n5762_), .A2(new_n5610_), .B1(new_n5591_), .B2(new_n5605_), .ZN(new_n5763_));
  XOR2_X1    g05692(.A1(new_n5084_), .A2(new_n5072_), .Z(new_n5764_));
  OAI21_X1   g05693(.A1(new_n5085_), .A2(new_n5086_), .B(new_n5059_), .ZN(new_n5765_));
  OAI21_X1   g05694(.A1(new_n5059_), .A2(new_n5764_), .B(new_n5765_), .ZN(new_n5766_));
  AOI22_X1   g05695(.A1(new_n4091_), .A2(new_n4613_), .B1(new_n4328_), .B2(new_n4767_), .ZN(new_n5767_));
  AOI21_X1   g05696(.A1(new_n117_), .A2(new_n4082_), .B(new_n5767_), .ZN(new_n5768_));
  OAI21_X1   g05697(.A1(new_n5768_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n5769_));
  XNOR2_X1   g05698(.A1(new_n5162_), .A2(new_n5769_), .ZN(new_n5770_));
  AND2_X2    g05699(.A1(new_n5766_), .A2(new_n5770_), .Z(new_n5771_));
  NOR2_X1    g05700(.A1(new_n5766_), .A2(new_n5770_), .ZN(new_n5772_));
  INV_X1     g05701(.I(new_n5772_), .ZN(new_n5773_));
  OAI21_X1   g05702(.A1(new_n5763_), .A2(new_n5771_), .B(new_n5773_), .ZN(new_n5774_));
  OAI22_X1   g05703(.A1(new_n4042_), .A2(new_n1239_), .B1(new_n4342_), .B2(new_n4981_), .ZN(new_n5775_));
  AOI21_X1   g05704(.A1(new_n5775_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n5776_));
  XNOR2_X1   g05705(.A1(new_n4864_), .A2(new_n5776_), .ZN(new_n5777_));
  INV_X1     g05706(.I(new_n5777_), .ZN(new_n5778_));
  NOR2_X1    g05707(.A1(new_n5778_), .A2(new_n5774_), .ZN(new_n5779_));
  NAND2_X1   g05708(.A1(new_n5778_), .A2(new_n5774_), .ZN(new_n5780_));
  OAI21_X1   g05709(.A1(new_n5588_), .A2(new_n5779_), .B(new_n5780_), .ZN(new_n5781_));
  INV_X1     g05710(.I(new_n5781_), .ZN(new_n5782_));
  INV_X1     g05711(.I(new_n4981_), .ZN(new_n5783_));
  AOI22_X1   g05712(.A1(new_n4347_), .A2(new_n5783_), .B1(new_n247_), .B2(new_n4036_), .ZN(new_n5784_));
  OAI21_X1   g05713(.A1(new_n5784_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n5785_));
  XOR2_X1    g05714(.A1(new_n4672_), .A2(new_n5785_), .Z(new_n5786_));
  NOR2_X1    g05715(.A1(new_n5782_), .A2(new_n5786_), .ZN(new_n5787_));
  XNOR2_X1   g05716(.A1(new_n5381_), .A2(new_n5385_), .ZN(new_n5788_));
  XOR2_X1    g05717(.A1(new_n5788_), .A2(new_n5376_), .Z(new_n5789_));
  AOI21_X1   g05718(.A1(new_n5782_), .A2(new_n5786_), .B(new_n5789_), .ZN(new_n5790_));
  NOR2_X1    g05719(.A1(new_n5790_), .A2(new_n5787_), .ZN(new_n5791_));
  AOI22_X1   g05720(.A1(new_n4445_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4399_), .ZN(new_n5792_));
  OAI21_X1   g05721(.A1(new_n5792_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n5793_));
  XOR2_X1    g05722(.A1(new_n4403_), .A2(new_n5793_), .Z(new_n5794_));
  AND2_X2    g05723(.A1(new_n5791_), .A2(new_n5794_), .Z(new_n5795_));
  NOR2_X1    g05724(.A1(new_n5791_), .A2(new_n5794_), .ZN(new_n5796_));
  NOR2_X1    g05725(.A1(new_n5795_), .A2(new_n5796_), .ZN(new_n5797_));
  NOR2_X1    g05726(.A1(new_n5797_), .A2(new_n5582_), .ZN(new_n5798_));
  XNOR2_X1   g05727(.A1(new_n5791_), .A2(new_n5794_), .ZN(new_n5799_));
  INV_X1     g05728(.I(new_n5799_), .ZN(new_n5800_));
  AOI21_X1   g05729(.A1(new_n5582_), .A2(new_n5800_), .B(new_n5798_), .ZN(new_n5801_));
  NOR2_X1    g05730(.A1(new_n5771_), .A2(new_n5772_), .ZN(new_n5802_));
  NOR2_X1    g05731(.A1(new_n5802_), .A2(new_n5763_), .ZN(new_n5803_));
  XNOR2_X1   g05732(.A1(new_n5766_), .A2(new_n5770_), .ZN(new_n5804_));
  INV_X1     g05733(.I(new_n5804_), .ZN(new_n5805_));
  AOI21_X1   g05734(.A1(new_n5763_), .A2(new_n5805_), .B(new_n5803_), .ZN(new_n5806_));
  INV_X1     g05735(.I(new_n5806_), .ZN(new_n5807_));
  NOR2_X1    g05736(.A1(new_n5611_), .A2(new_n5609_), .ZN(new_n5808_));
  XOR2_X1    g05737(.A1(new_n5761_), .A2(new_n5808_), .Z(new_n5809_));
  XOR2_X1    g05738(.A1(new_n5809_), .A2(new_n5605_), .Z(new_n5810_));
  INV_X1     g05739(.I(new_n5810_), .ZN(new_n5811_));
  OAI22_X1   g05740(.A1(new_n4315_), .A2(new_n4612_), .B1(new_n4099_), .B2(new_n4781_), .ZN(new_n5812_));
  OAI21_X1   g05741(.A1(new_n4090_), .A2(new_n1128_), .B(new_n5812_), .ZN(new_n5813_));
  AOI21_X1   g05742(.A1(new_n5813_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n5814_));
  XOR2_X1    g05743(.A1(new_n5196_), .A2(new_n5814_), .Z(new_n5815_));
  OAI22_X1   g05744(.A1(new_n4123_), .A2(new_n4527_), .B1(new_n4309_), .B2(new_n4529_), .ZN(new_n5816_));
  OAI21_X1   g05745(.A1(new_n4112_), .A2(new_n79_), .B(new_n5816_), .ZN(new_n5817_));
  AOI21_X1   g05746(.A1(new_n5817_), .A2(new_n72_), .B(new_n79_), .ZN(new_n5818_));
  XOR2_X1    g05747(.A1(new_n5096_), .A2(new_n5818_), .Z(new_n5819_));
  NOR2_X1    g05748(.A1(new_n5815_), .A2(new_n5819_), .ZN(new_n5820_));
  XNOR2_X1   g05749(.A1(new_n5760_), .A2(new_n5613_), .ZN(new_n5821_));
  INV_X1     g05750(.I(new_n5815_), .ZN(new_n5822_));
  INV_X1     g05751(.I(new_n5819_), .ZN(new_n5823_));
  NOR2_X1    g05752(.A1(new_n5822_), .A2(new_n5823_), .ZN(new_n5824_));
  INV_X1     g05753(.I(new_n5824_), .ZN(new_n5825_));
  AOI21_X1   g05754(.A1(new_n5821_), .A2(new_n5825_), .B(new_n5820_), .ZN(new_n5826_));
  INV_X1     g05755(.I(new_n5826_), .ZN(new_n5827_));
  AOI22_X1   g05756(.A1(new_n4091_), .A2(new_n4767_), .B1(new_n4100_), .B2(new_n4613_), .ZN(new_n5828_));
  AOI21_X1   g05757(.A1(new_n117_), .A2(new_n4328_), .B(new_n5828_), .ZN(new_n5829_));
  OAI21_X1   g05758(.A1(new_n5829_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n5830_));
  XNOR2_X1   g05759(.A1(new_n5139_), .A2(new_n5830_), .ZN(new_n5831_));
  INV_X1     g05760(.I(new_n5831_), .ZN(new_n5832_));
  NOR2_X1    g05761(.A1(new_n5827_), .A2(new_n5832_), .ZN(new_n5833_));
  INV_X1     g05762(.I(new_n5833_), .ZN(new_n5834_));
  NOR2_X1    g05763(.A1(new_n5826_), .A2(new_n5831_), .ZN(new_n5835_));
  AOI21_X1   g05764(.A1(new_n5811_), .A2(new_n5834_), .B(new_n5835_), .ZN(new_n5836_));
  INV_X1     g05765(.I(new_n5836_), .ZN(new_n5837_));
  OAI22_X1   g05766(.A1(new_n4339_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4053_), .ZN(new_n5838_));
  AOI21_X1   g05767(.A1(new_n5838_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n5839_));
  XNOR2_X1   g05768(.A1(new_n4652_), .A2(new_n5839_), .ZN(new_n5840_));
  INV_X1     g05769(.I(new_n5840_), .ZN(new_n5841_));
  NOR2_X1    g05770(.A1(new_n5837_), .A2(new_n5841_), .ZN(new_n5842_));
  INV_X1     g05771(.I(new_n5842_), .ZN(new_n5843_));
  NOR2_X1    g05772(.A1(new_n5836_), .A2(new_n5840_), .ZN(new_n5844_));
  AOI21_X1   g05773(.A1(new_n5843_), .A2(new_n5807_), .B(new_n5844_), .ZN(new_n5845_));
  OAI22_X1   g05774(.A1(new_n4028_), .A2(new_n5335_), .B1(new_n4035_), .B2(new_n4719_), .ZN(new_n5846_));
  OAI21_X1   g05775(.A1(new_n4017_), .A2(new_n5398_), .B(new_n5846_), .ZN(new_n5847_));
  AOI21_X1   g05776(.A1(new_n5847_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n5848_));
  XNOR2_X1   g05777(.A1(new_n4705_), .A2(new_n5848_), .ZN(new_n5849_));
  INV_X1     g05778(.I(new_n5780_), .ZN(new_n5850_));
  NOR2_X1    g05779(.A1(new_n5850_), .A2(new_n5779_), .ZN(new_n5851_));
  XNOR2_X1   g05780(.A1(new_n5777_), .A2(new_n5774_), .ZN(new_n5852_));
  NAND2_X1   g05781(.A1(new_n5852_), .A2(new_n5588_), .ZN(new_n5853_));
  OAI21_X1   g05782(.A1(new_n5588_), .A2(new_n5851_), .B(new_n5853_), .ZN(new_n5854_));
  INV_X1     g05783(.I(new_n5845_), .ZN(new_n5855_));
  INV_X1     g05784(.I(new_n5849_), .ZN(new_n5856_));
  OAI21_X1   g05785(.A1(new_n5856_), .A2(new_n5855_), .B(new_n5854_), .ZN(new_n5857_));
  OAI21_X1   g05786(.A1(new_n5845_), .A2(new_n5849_), .B(new_n5857_), .ZN(new_n5858_));
  INV_X1     g05787(.I(new_n4355_), .ZN(new_n5859_));
  AOI22_X1   g05788(.A1(new_n5859_), .A2(new_n5337_), .B1(new_n4375_), .B2(new_n4717_), .ZN(new_n5860_));
  OAI21_X1   g05789(.A1(new_n5860_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n5861_));
  XNOR2_X1   g05790(.A1(new_n4730_), .A2(new_n5861_), .ZN(new_n5862_));
  NAND2_X1   g05791(.A1(new_n5858_), .A2(new_n5862_), .ZN(new_n5863_));
  NOR2_X1    g05792(.A1(new_n5858_), .A2(new_n5862_), .ZN(new_n5864_));
  XOR2_X1    g05793(.A1(new_n5786_), .A2(new_n5377_), .Z(new_n5865_));
  NOR2_X1    g05794(.A1(new_n5865_), .A2(new_n5788_), .ZN(new_n5866_));
  INV_X1     g05795(.I(new_n5788_), .ZN(new_n5867_));
  XOR2_X1    g05796(.A1(new_n5786_), .A2(new_n5376_), .Z(new_n5868_));
  NOR2_X1    g05797(.A1(new_n5868_), .A2(new_n5867_), .ZN(new_n5869_));
  NOR2_X1    g05798(.A1(new_n5869_), .A2(new_n5866_), .ZN(new_n5870_));
  XOR2_X1    g05799(.A1(new_n5870_), .A2(new_n5781_), .Z(new_n5871_));
  OAI21_X1   g05800(.A1(new_n5864_), .A2(new_n5871_), .B(new_n5863_), .ZN(new_n5872_));
  AOI22_X1   g05801(.A1(new_n4473_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4555_), .ZN(new_n5873_));
  OAI21_X1   g05802(.A1(new_n5873_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n5874_));
  NOR2_X1    g05803(.A1(new_n4585_), .A2(new_n5874_), .ZN(new_n5875_));
  NAND2_X1   g05804(.A1(new_n4585_), .A2(new_n5874_), .ZN(new_n5876_));
  INV_X1     g05805(.I(new_n5876_), .ZN(new_n5877_));
  NOR2_X1    g05806(.A1(new_n5877_), .A2(new_n5875_), .ZN(new_n5878_));
  INV_X1     g05807(.I(new_n5878_), .ZN(new_n5879_));
  NOR2_X1    g05808(.A1(new_n5879_), .A2(new_n5872_), .ZN(new_n5880_));
  INV_X1     g05809(.I(new_n5880_), .ZN(new_n5881_));
  NAND2_X1   g05810(.A1(new_n5879_), .A2(new_n5872_), .ZN(new_n5882_));
  AOI21_X1   g05811(.A1(new_n5881_), .A2(new_n5882_), .B(new_n5801_), .ZN(new_n5883_));
  INV_X1     g05812(.I(new_n5801_), .ZN(new_n5884_));
  XOR2_X1    g05813(.A1(new_n5878_), .A2(new_n5872_), .Z(new_n5885_));
  NOR2_X1    g05814(.A1(new_n5885_), .A2(new_n5884_), .ZN(new_n5886_));
  NOR2_X1    g05815(.A1(new_n5883_), .A2(new_n5886_), .ZN(new_n5887_));
  XOR2_X1    g05816(.A1(new_n5849_), .A2(new_n5845_), .Z(new_n5888_));
  XOR2_X1    g05817(.A1(new_n5849_), .A2(new_n5855_), .Z(new_n5889_));
  MUX2_X1    g05818(.I0(new_n5889_), .I1(new_n5888_), .S(new_n5854_), .Z(new_n5890_));
  NOR2_X1    g05819(.A1(new_n5842_), .A2(new_n5844_), .ZN(new_n5891_));
  NOR2_X1    g05820(.A1(new_n5891_), .A2(new_n5806_), .ZN(new_n5892_));
  XNOR2_X1   g05821(.A1(new_n5836_), .A2(new_n5840_), .ZN(new_n5893_));
  NOR2_X1    g05822(.A1(new_n5893_), .A2(new_n5807_), .ZN(new_n5894_));
  NOR2_X1    g05823(.A1(new_n5892_), .A2(new_n5894_), .ZN(new_n5895_));
  INV_X1     g05824(.I(new_n5895_), .ZN(new_n5896_));
  XOR2_X1    g05825(.A1(new_n5815_), .A2(new_n5823_), .Z(new_n5897_));
  OR2_X2     g05826(.A1(new_n5821_), .A2(new_n5897_), .Z(new_n5898_));
  OAI21_X1   g05827(.A1(new_n5820_), .A2(new_n5824_), .B(new_n5821_), .ZN(new_n5899_));
  NAND2_X1   g05828(.A1(new_n5898_), .A2(new_n5899_), .ZN(new_n5900_));
  AOI22_X1   g05829(.A1(new_n4113_), .A2(new_n4613_), .B1(new_n4105_), .B2(new_n4767_), .ZN(new_n5901_));
  AOI21_X1   g05830(.A1(new_n117_), .A2(new_n4100_), .B(new_n5901_), .ZN(new_n5902_));
  OAI21_X1   g05831(.A1(new_n5902_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n5903_));
  XOR2_X1    g05832(.A1(new_n5080_), .A2(new_n5903_), .Z(new_n5904_));
  INV_X1     g05833(.I(new_n5064_), .ZN(new_n5905_));
  NOR2_X1    g05834(.A1(new_n5905_), .A2(new_n5065_), .ZN(new_n5906_));
  OAI22_X1   g05835(.A1(new_n4131_), .A2(new_n4529_), .B1(new_n4309_), .B2(new_n4527_), .ZN(new_n5907_));
  OAI21_X1   g05836(.A1(new_n79_), .A2(new_n4123_), .B(new_n5907_), .ZN(new_n5908_));
  AOI21_X1   g05837(.A1(new_n5908_), .A2(new_n72_), .B(new_n79_), .ZN(new_n5909_));
  XOR2_X1    g05838(.A1(new_n5906_), .A2(new_n5909_), .Z(new_n5910_));
  NOR2_X1    g05839(.A1(new_n5904_), .A2(new_n5910_), .ZN(new_n5911_));
  NAND2_X1   g05840(.A1(new_n5904_), .A2(new_n5910_), .ZN(new_n5912_));
  XOR2_X1    g05841(.A1(new_n5757_), .A2(new_n5614_), .Z(new_n5913_));
  XOR2_X1    g05842(.A1(new_n5748_), .A2(new_n5913_), .Z(new_n5914_));
  INV_X1     g05843(.I(new_n5914_), .ZN(new_n5915_));
  AOI21_X1   g05844(.A1(new_n5915_), .A2(new_n5912_), .B(new_n5911_), .ZN(new_n5916_));
  NOR2_X1    g05845(.A1(new_n4331_), .A2(new_n4081_), .ZN(new_n5917_));
  OAI22_X1   g05846(.A1(new_n4070_), .A2(new_n1239_), .B1(new_n4981_), .B2(new_n5917_), .ZN(new_n5918_));
  AOI21_X1   g05847(.A1(new_n5918_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n5919_));
  XOR2_X1    g05848(.A1(new_n4927_), .A2(new_n5919_), .Z(new_n5920_));
  NAND2_X1   g05849(.A1(new_n5920_), .A2(new_n5916_), .ZN(new_n5921_));
  NOR2_X1    g05850(.A1(new_n5920_), .A2(new_n5916_), .ZN(new_n5922_));
  AOI21_X1   g05851(.A1(new_n5900_), .A2(new_n5921_), .B(new_n5922_), .ZN(new_n5923_));
  OAI22_X1   g05852(.A1(new_n4336_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4060_), .ZN(new_n5924_));
  AOI21_X1   g05853(.A1(new_n5924_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n5925_));
  XNOR2_X1   g05854(.A1(new_n4935_), .A2(new_n5925_), .ZN(new_n5926_));
  NOR2_X1    g05855(.A1(new_n5923_), .A2(new_n5926_), .ZN(new_n5927_));
  XOR2_X1    g05856(.A1(new_n5826_), .A2(new_n5832_), .Z(new_n5928_));
  OAI21_X1   g05857(.A1(new_n5833_), .A2(new_n5835_), .B(new_n5810_), .ZN(new_n5929_));
  OAI21_X1   g05858(.A1(new_n5810_), .A2(new_n5928_), .B(new_n5929_), .ZN(new_n5930_));
  INV_X1     g05859(.I(new_n5930_), .ZN(new_n5931_));
  NAND2_X1   g05860(.A1(new_n5923_), .A2(new_n5926_), .ZN(new_n5932_));
  AOI21_X1   g05861(.A1(new_n5931_), .A2(new_n5932_), .B(new_n5927_), .ZN(new_n5933_));
  INV_X1     g05862(.I(new_n5933_), .ZN(new_n5934_));
  INV_X1     g05863(.I(new_n4349_), .ZN(new_n5935_));
  AOI22_X1   g05864(.A1(new_n5935_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4029_), .ZN(new_n5936_));
  OAI21_X1   g05865(.A1(new_n5936_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n5937_));
  XOR2_X1    g05866(.A1(new_n4687_), .A2(new_n5937_), .Z(new_n5938_));
  INV_X1     g05867(.I(new_n5938_), .ZN(new_n5939_));
  NOR2_X1    g05868(.A1(new_n5939_), .A2(new_n5934_), .ZN(new_n5940_));
  INV_X1     g05869(.I(new_n5940_), .ZN(new_n5941_));
  NOR2_X1    g05870(.A1(new_n5938_), .A2(new_n5933_), .ZN(new_n5942_));
  AOI21_X1   g05871(.A1(new_n5941_), .A2(new_n5896_), .B(new_n5942_), .ZN(new_n5943_));
  INV_X1     g05872(.I(new_n5943_), .ZN(new_n5944_));
  OAI22_X1   g05873(.A1(new_n4397_), .A2(new_n5419_), .B1(new_n1622_), .B2(new_n4374_), .ZN(new_n5945_));
  OAI21_X1   g05874(.A1(new_n4437_), .A2(new_n1620_), .B(new_n5945_), .ZN(new_n5946_));
  AOI21_X1   g05875(.A1(new_n5946_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n5947_));
  XOR2_X1    g05876(.A1(new_n4541_), .A2(new_n5947_), .Z(new_n5948_));
  INV_X1     g05877(.I(new_n5948_), .ZN(new_n5949_));
  NOR2_X1    g05878(.A1(new_n5949_), .A2(new_n5944_), .ZN(new_n5950_));
  NOR2_X1    g05879(.A1(new_n5950_), .A2(new_n5890_), .ZN(new_n5951_));
  NOR2_X1    g05880(.A1(new_n5948_), .A2(new_n5943_), .ZN(new_n5952_));
  NOR2_X1    g05881(.A1(new_n5951_), .A2(new_n5952_), .ZN(new_n5953_));
  AOI22_X1   g05882(.A1(new_n4448_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4469_), .ZN(new_n5954_));
  OAI21_X1   g05883(.A1(new_n5954_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n5955_));
  XNOR2_X1   g05884(.A1(new_n4477_), .A2(new_n5955_), .ZN(new_n5956_));
  NOR2_X1    g05885(.A1(new_n5953_), .A2(new_n5956_), .ZN(new_n5957_));
  XOR2_X1    g05886(.A1(new_n5862_), .A2(new_n5781_), .Z(new_n5958_));
  NOR2_X1    g05887(.A1(new_n5958_), .A2(new_n5870_), .ZN(new_n5959_));
  XOR2_X1    g05888(.A1(new_n5862_), .A2(new_n5782_), .Z(new_n5960_));
  NOR3_X1    g05889(.A1(new_n5960_), .A2(new_n5866_), .A3(new_n5869_), .ZN(new_n5961_));
  NOR2_X1    g05890(.A1(new_n5961_), .A2(new_n5959_), .ZN(new_n5962_));
  XOR2_X1    g05891(.A1(new_n5962_), .A2(new_n5858_), .Z(new_n5963_));
  AOI21_X1   g05892(.A1(new_n5953_), .A2(new_n5956_), .B(new_n5963_), .ZN(new_n5964_));
  NOR2_X1    g05893(.A1(new_n5964_), .A2(new_n5957_), .ZN(new_n5965_));
  INV_X1     g05894(.I(new_n4943_), .ZN(new_n5966_));
  NOR2_X1    g05895(.A1(new_n5966_), .A2(new_n1851_), .ZN(new_n5967_));
  INV_X1     g05896(.I(new_n5967_), .ZN(new_n5968_));
  AOI22_X1   g05897(.A1(new_n5418_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4563_), .ZN(new_n5969_));
  OAI21_X1   g05898(.A1(new_n5969_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n5970_));
  XNOR2_X1   g05899(.A1(new_n4594_), .A2(new_n5970_), .ZN(new_n5971_));
  AND2_X2    g05900(.A1(new_n5965_), .A2(new_n5971_), .Z(new_n5972_));
  NOR2_X1    g05901(.A1(new_n5972_), .A2(new_n5887_), .ZN(new_n5973_));
  NOR2_X1    g05902(.A1(new_n5965_), .A2(new_n5971_), .ZN(new_n5974_));
  NOR2_X1    g05903(.A1(new_n5973_), .A2(new_n5974_), .ZN(new_n5975_));
  OAI21_X1   g05904(.A1(new_n5404_), .A2(new_n5406_), .B(new_n5353_), .ZN(new_n5976_));
  XOR2_X1    g05905(.A1(new_n5402_), .A2(new_n5397_), .Z(new_n5977_));
  OAI21_X1   g05906(.A1(new_n5353_), .A2(new_n5977_), .B(new_n5976_), .ZN(new_n5978_));
  INV_X1     g05907(.I(new_n5978_), .ZN(new_n5979_));
  NOR2_X1    g05908(.A1(new_n5795_), .A2(new_n5582_), .ZN(new_n5980_));
  NOR2_X1    g05909(.A1(new_n5980_), .A2(new_n5796_), .ZN(new_n5981_));
  OAI22_X1   g05910(.A1(new_n1622_), .A2(new_n4468_), .B1(new_n4501_), .B2(new_n5419_), .ZN(new_n5982_));
  OAI21_X1   g05911(.A1(new_n4516_), .A2(new_n1620_), .B(new_n5982_), .ZN(new_n5983_));
  AOI21_X1   g05912(.A1(new_n5983_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n5984_));
  XOR2_X1    g05913(.A1(new_n4524_), .A2(new_n5984_), .Z(new_n5985_));
  AND2_X2    g05914(.A1(new_n5985_), .A2(new_n5981_), .Z(new_n5986_));
  NOR2_X1    g05915(.A1(new_n5985_), .A2(new_n5981_), .ZN(new_n5987_));
  NOR2_X1    g05916(.A1(new_n5986_), .A2(new_n5987_), .ZN(new_n5988_));
  NOR2_X1    g05917(.A1(new_n5988_), .A2(new_n5979_), .ZN(new_n5989_));
  XNOR2_X1   g05918(.A1(new_n5985_), .A2(new_n5981_), .ZN(new_n5990_));
  NOR2_X1    g05919(.A1(new_n5990_), .A2(new_n5978_), .ZN(new_n5991_));
  NOR2_X1    g05920(.A1(new_n5989_), .A2(new_n5991_), .ZN(new_n5992_));
  OAI21_X1   g05921(.A1(new_n5801_), .A2(new_n5880_), .B(new_n5882_), .ZN(new_n5993_));
  NAND2_X1   g05922(.A1(new_n4563_), .A2(new_n4943_), .ZN(new_n5994_));
  NAND2_X1   g05923(.A1(new_n4564_), .A2(new_n4941_), .ZN(new_n5995_));
  AOI22_X1   g05924(.A1(new_n5995_), .A2(new_n5994_), .B1(new_n785_), .B2(new_n4564_), .ZN(new_n5996_));
  OAI21_X1   g05925(.A1(new_n5996_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n5997_));
  XOR2_X1    g05926(.A1(new_n4609_), .A2(new_n5997_), .Z(new_n5998_));
  INV_X1     g05927(.I(new_n5998_), .ZN(new_n5999_));
  NOR2_X1    g05928(.A1(new_n5993_), .A2(new_n5999_), .ZN(new_n6000_));
  INV_X1     g05929(.I(new_n5993_), .ZN(new_n6001_));
  NOR2_X1    g05930(.A1(new_n6001_), .A2(new_n5998_), .ZN(new_n6002_));
  NOR2_X1    g05931(.A1(new_n6002_), .A2(new_n6000_), .ZN(new_n6003_));
  NOR2_X1    g05932(.A1(new_n6003_), .A2(new_n5992_), .ZN(new_n6004_));
  INV_X1     g05933(.I(new_n5992_), .ZN(new_n6005_));
  XOR2_X1    g05934(.A1(new_n5993_), .A2(new_n5998_), .Z(new_n6006_));
  NOR2_X1    g05935(.A1(new_n6006_), .A2(new_n6005_), .ZN(new_n6007_));
  NOR2_X1    g05936(.A1(new_n6004_), .A2(new_n6007_), .ZN(new_n6008_));
  INV_X1     g05937(.I(new_n6008_), .ZN(new_n6009_));
  NOR2_X1    g05938(.A1(new_n6009_), .A2(new_n1079_), .ZN(new_n6010_));
  NOR2_X1    g05939(.A1(new_n6010_), .A2(new_n5975_), .ZN(new_n6011_));
  NOR2_X1    g05940(.A1(new_n6008_), .A2(new_n806_), .ZN(new_n6012_));
  NOR2_X1    g05941(.A1(new_n6011_), .A2(new_n6012_), .ZN(new_n6013_));
  INV_X1     g05942(.I(new_n6000_), .ZN(new_n6014_));
  AOI21_X1   g05943(.A1(new_n6005_), .A2(new_n6014_), .B(new_n6002_), .ZN(new_n6015_));
  AOI22_X1   g05944(.A1(new_n5553_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4564_), .ZN(new_n6016_));
  OAI21_X1   g05945(.A1(new_n6016_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n6017_));
  XOR2_X1    g05946(.A1(new_n4569_), .A2(new_n6017_), .Z(new_n6018_));
  INV_X1     g05947(.I(new_n5986_), .ZN(new_n6019_));
  AOI21_X1   g05948(.A1(new_n6019_), .A2(new_n5978_), .B(new_n5987_), .ZN(new_n6020_));
  NAND2_X1   g05949(.A1(new_n5413_), .A2(new_n5414_), .ZN(new_n6021_));
  XOR2_X1    g05950(.A1(new_n6021_), .A2(new_n5410_), .Z(new_n6022_));
  XNOR2_X1   g05951(.A1(new_n6022_), .A2(new_n5407_), .ZN(new_n6023_));
  XNOR2_X1   g05952(.A1(new_n6023_), .A2(new_n6020_), .ZN(new_n6024_));
  XNOR2_X1   g05953(.A1(new_n6024_), .A2(new_n6018_), .ZN(new_n6025_));
  NAND2_X1   g05954(.A1(new_n4943_), .A2(new_n785_), .ZN(new_n6026_));
  OAI21_X1   g05955(.A1(new_n4941_), .A2(new_n6026_), .B(new_n4564_), .ZN(new_n6027_));
  OAI21_X1   g05956(.A1(new_n6027_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n6028_));
  XOR2_X1    g05957(.A1(new_n5001_), .A2(new_n6028_), .Z(new_n6029_));
  XOR2_X1    g05958(.A1(new_n6025_), .A2(new_n6029_), .Z(new_n6030_));
  NOR2_X1    g05959(.A1(new_n6030_), .A2(new_n6015_), .ZN(new_n6031_));
  INV_X1     g05960(.I(new_n6029_), .ZN(new_n6032_));
  NOR2_X1    g05961(.A1(new_n6025_), .A2(new_n6032_), .ZN(new_n6033_));
  INV_X1     g05962(.I(new_n6033_), .ZN(new_n6034_));
  NAND2_X1   g05963(.A1(new_n6025_), .A2(new_n6032_), .ZN(new_n6035_));
  NAND2_X1   g05964(.A1(new_n6034_), .A2(new_n6035_), .ZN(new_n6036_));
  AOI21_X1   g05965(.A1(new_n6015_), .A2(new_n6036_), .B(new_n6031_), .ZN(new_n6037_));
  NOR2_X1    g05966(.A1(new_n6037_), .A2(new_n6013_), .ZN(new_n6038_));
  AOI22_X1   g05967(.A1(new_n4445_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4399_), .ZN(new_n6039_));
  OAI21_X1   g05968(.A1(new_n6039_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n6040_));
  XOR2_X1    g05969(.A1(new_n4403_), .A2(new_n6040_), .Z(new_n6041_));
  INV_X1     g05970(.I(new_n6041_), .ZN(new_n6042_));
  INV_X1     g05971(.I(new_n5920_), .ZN(new_n6043_));
  XNOR2_X1   g05972(.A1(new_n5904_), .A2(new_n5913_), .ZN(new_n6044_));
  XOR2_X1    g05973(.A1(new_n6044_), .A2(new_n5748_), .Z(new_n6045_));
  XOR2_X1    g05974(.A1(new_n6045_), .A2(new_n5910_), .Z(new_n6046_));
  AOI22_X1   g05975(.A1(new_n5701_), .A2(new_n4526_), .B1(new_n4171_), .B2(new_n4570_), .ZN(new_n6047_));
  AOI21_X1   g05976(.A1(new_n101_), .A2(new_n4274_), .B(new_n6047_), .ZN(new_n6048_));
  OAI21_X1   g05977(.A1(new_n6048_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n6049_));
  XNOR2_X1   g05978(.A1(new_n5722_), .A2(new_n6049_), .ZN(new_n6050_));
  INV_X1     g05979(.I(new_n6050_), .ZN(new_n6051_));
  NOR2_X1    g05980(.A1(new_n4251_), .A2(new_n935_), .ZN(new_n6052_));
  INV_X1     g05981(.I(new_n6052_), .ZN(new_n6053_));
  NAND2_X1   g05982(.A1(new_n4252_), .A2(new_n4570_), .ZN(new_n6054_));
  OAI21_X1   g05983(.A1(new_n4234_), .A2(new_n4527_), .B(new_n6054_), .ZN(new_n6055_));
  OAI21_X1   g05984(.A1(new_n79_), .A2(new_n4249_), .B(new_n6055_), .ZN(new_n6056_));
  AOI21_X1   g05985(.A1(new_n6056_), .A2(new_n72_), .B(new_n79_), .ZN(new_n6057_));
  XOR2_X1    g05986(.A1(new_n5648_), .A2(new_n6057_), .Z(new_n6058_));
  NAND2_X1   g05987(.A1(new_n6058_), .A2(new_n6053_), .ZN(new_n6059_));
  NAND2_X1   g05988(.A1(new_n5627_), .A2(new_n79_), .ZN(new_n6060_));
  NAND2_X1   g05989(.A1(new_n4251_), .A2(new_n4252_), .ZN(new_n6061_));
  AOI21_X1   g05990(.A1(new_n101_), .A2(new_n6061_), .B(new_n4260_), .ZN(new_n6062_));
  OAI22_X1   g05991(.A1(new_n4244_), .A2(new_n4527_), .B1(new_n4230_), .B2(new_n4529_), .ZN(new_n6063_));
  OAI21_X1   g05992(.A1(new_n79_), .A2(new_n4234_), .B(new_n6063_), .ZN(new_n6064_));
  AOI21_X1   g05993(.A1(new_n6060_), .A2(new_n6062_), .B(new_n6064_), .ZN(new_n6065_));
  XOR2_X1    g05994(.A1(new_n6065_), .A2(new_n72_), .Z(new_n6066_));
  AOI21_X1   g05995(.A1(new_n4251_), .A2(new_n101_), .B(\a[29] ), .ZN(new_n6067_));
  NAND2_X1   g05996(.A1(new_n6067_), .A2(new_n6054_), .ZN(new_n6068_));
  NAND2_X1   g05997(.A1(new_n6068_), .A2(new_n101_), .ZN(new_n6069_));
  XNOR2_X1   g05998(.A1(new_n6069_), .A2(new_n5637_), .ZN(new_n6070_));
  INV_X1     g05999(.I(new_n6070_), .ZN(new_n6071_));
  NOR2_X1    g06000(.A1(new_n4251_), .A2(new_n918_), .ZN(new_n6072_));
  NOR2_X1    g06001(.A1(new_n6072_), .A2(new_n72_), .ZN(new_n6073_));
  INV_X1     g06002(.I(new_n6073_), .ZN(new_n6074_));
  NOR3_X1    g06003(.A1(new_n6066_), .A2(new_n6071_), .A3(new_n6074_), .ZN(new_n6075_));
  NOR2_X1    g06004(.A1(new_n6058_), .A2(new_n6053_), .ZN(new_n6076_));
  OAI21_X1   g06005(.A1(new_n6075_), .A2(new_n6076_), .B(new_n6059_), .ZN(new_n6077_));
  AOI21_X1   g06006(.A1(new_n5676_), .A2(new_n4246_), .B(new_n4203_), .ZN(new_n6078_));
  INV_X1     g06007(.I(new_n5657_), .ZN(new_n6079_));
  OAI21_X1   g06008(.A1(new_n4255_), .A2(new_n4251_), .B(new_n4221_), .ZN(new_n6080_));
  AOI21_X1   g06009(.A1(new_n6080_), .A2(new_n6079_), .B(new_n5655_), .ZN(new_n6081_));
  NOR2_X1    g06010(.A1(new_n6081_), .A2(new_n6078_), .ZN(new_n6082_));
  OAI22_X1   g06011(.A1(new_n4249_), .A2(new_n4527_), .B1(new_n4234_), .B2(new_n4529_), .ZN(new_n6083_));
  OAI21_X1   g06012(.A1(new_n4203_), .A2(new_n79_), .B(new_n6083_), .ZN(new_n6084_));
  AOI21_X1   g06013(.A1(new_n6084_), .A2(new_n72_), .B(new_n79_), .ZN(new_n6085_));
  XOR2_X1    g06014(.A1(new_n6082_), .A2(new_n6085_), .Z(new_n6086_));
  NAND2_X1   g06015(.A1(new_n6086_), .A2(new_n5638_), .ZN(new_n6087_));
  NOR2_X1    g06016(.A1(new_n6086_), .A2(new_n5638_), .ZN(new_n6088_));
  AOI21_X1   g06017(.A1(new_n6077_), .A2(new_n6087_), .B(new_n6088_), .ZN(new_n6089_));
  OAI22_X1   g06018(.A1(new_n4203_), .A2(new_n4527_), .B1(new_n4249_), .B2(new_n4529_), .ZN(new_n6090_));
  OAI21_X1   g06019(.A1(new_n79_), .A2(new_n4175_), .B(new_n6090_), .ZN(new_n6091_));
  AOI21_X1   g06020(.A1(new_n6091_), .A2(new_n72_), .B(new_n79_), .ZN(new_n6092_));
  XOR2_X1    g06021(.A1(new_n5671_), .A2(new_n6092_), .Z(new_n6093_));
  INV_X1     g06022(.I(new_n5638_), .ZN(new_n6094_));
  XOR2_X1    g06023(.A1(new_n5632_), .A2(new_n6094_), .Z(new_n6095_));
  INV_X1     g06024(.I(new_n6095_), .ZN(new_n6096_));
  NOR2_X1    g06025(.A1(new_n6093_), .A2(new_n6096_), .ZN(new_n6097_));
  NAND2_X1   g06026(.A1(new_n6093_), .A2(new_n6096_), .ZN(new_n6098_));
  OAI21_X1   g06027(.A1(new_n6089_), .A2(new_n6097_), .B(new_n6098_), .ZN(new_n6099_));
  NOR2_X1    g06028(.A1(new_n5691_), .A2(new_n4258_), .ZN(new_n6100_));
  AOI21_X1   g06029(.A1(new_n5687_), .A2(new_n5679_), .B(new_n4175_), .ZN(new_n6101_));
  NOR2_X1    g06030(.A1(new_n6100_), .A2(new_n6101_), .ZN(new_n6102_));
  OAI22_X1   g06031(.A1(new_n4175_), .A2(new_n4527_), .B1(new_n4203_), .B2(new_n4529_), .ZN(new_n6103_));
  OAI21_X1   g06032(.A1(new_n79_), .A2(new_n5684_), .B(new_n6103_), .ZN(new_n6104_));
  AOI21_X1   g06033(.A1(new_n6104_), .A2(new_n72_), .B(new_n79_), .ZN(new_n6105_));
  XOR2_X1    g06034(.A1(new_n6102_), .A2(new_n6105_), .Z(new_n6106_));
  XNOR2_X1   g06035(.A1(new_n5639_), .A2(new_n5651_), .ZN(new_n6107_));
  NAND2_X1   g06036(.A1(new_n6106_), .A2(new_n6107_), .ZN(new_n6108_));
  NAND2_X1   g06037(.A1(new_n6108_), .A2(new_n6099_), .ZN(new_n6109_));
  XOR2_X1    g06038(.A1(new_n5693_), .A2(new_n6105_), .Z(new_n6110_));
  INV_X1     g06039(.I(new_n6107_), .ZN(new_n6111_));
  NAND2_X1   g06040(.A1(new_n6110_), .A2(new_n6111_), .ZN(new_n6112_));
  OAI22_X1   g06041(.A1(new_n5684_), .A2(new_n4527_), .B1(new_n4175_), .B2(new_n4529_), .ZN(new_n6113_));
  OAI21_X1   g06042(.A1(new_n4150_), .A2(new_n79_), .B(new_n6113_), .ZN(new_n6114_));
  AOI21_X1   g06043(.A1(new_n6114_), .A2(new_n72_), .B(new_n79_), .ZN(new_n6115_));
  XOR2_X1    g06044(.A1(new_n5707_), .A2(new_n6115_), .Z(new_n6116_));
  NAND2_X1   g06045(.A1(new_n5660_), .A2(new_n5663_), .ZN(new_n6117_));
  XOR2_X1    g06046(.A1(new_n5652_), .A2(new_n6117_), .Z(new_n6118_));
  NAND2_X1   g06047(.A1(new_n6116_), .A2(new_n6118_), .ZN(new_n6119_));
  INV_X1     g06048(.I(new_n6119_), .ZN(new_n6120_));
  NOR2_X1    g06049(.A1(new_n6116_), .A2(new_n6118_), .ZN(new_n6121_));
  NOR2_X1    g06050(.A1(new_n6120_), .A2(new_n6121_), .ZN(new_n6122_));
  NAND3_X1   g06051(.A1(new_n6122_), .A2(new_n6109_), .A3(new_n6112_), .ZN(new_n6123_));
  NOR2_X1    g06052(.A1(new_n6123_), .A2(new_n6051_), .ZN(new_n6124_));
  XNOR2_X1   g06053(.A1(new_n5664_), .A2(new_n5675_), .ZN(new_n6125_));
  NOR2_X1    g06054(.A1(new_n6119_), .A2(new_n6125_), .ZN(new_n6126_));
  INV_X1     g06055(.I(new_n6126_), .ZN(new_n6127_));
  AOI21_X1   g06056(.A1(new_n6123_), .A2(new_n6051_), .B(new_n6127_), .ZN(new_n6128_));
  NOR2_X1    g06057(.A1(new_n6128_), .A2(new_n6124_), .ZN(new_n6129_));
  NOR2_X1    g06058(.A1(new_n5664_), .A2(new_n5675_), .ZN(new_n6130_));
  XOR2_X1    g06059(.A1(new_n5697_), .A2(new_n6130_), .Z(new_n6131_));
  NOR3_X1    g06060(.A1(new_n5731_), .A2(new_n5719_), .A3(new_n4274_), .ZN(new_n6132_));
  AOI21_X1   g06061(.A1(new_n5728_), .A2(new_n5729_), .B(new_n4273_), .ZN(new_n6133_));
  NOR2_X1    g06062(.A1(new_n6133_), .A2(new_n6132_), .ZN(new_n6134_));
  OAI22_X1   g06063(.A1(new_n4273_), .A2(new_n4527_), .B1(new_n4150_), .B2(new_n4529_), .ZN(new_n6135_));
  OAI21_X1   g06064(.A1(new_n79_), .A2(new_n4142_), .B(new_n6135_), .ZN(new_n6136_));
  AOI21_X1   g06065(.A1(new_n6136_), .A2(new_n72_), .B(new_n79_), .ZN(new_n6137_));
  XOR2_X1    g06066(.A1(new_n6134_), .A2(new_n6137_), .Z(new_n6138_));
  AND2_X2    g06067(.A1(new_n6138_), .A2(new_n6131_), .Z(new_n6139_));
  NOR2_X1    g06068(.A1(new_n6129_), .A2(new_n6139_), .ZN(new_n6140_));
  NOR2_X1    g06069(.A1(new_n6138_), .A2(new_n6131_), .ZN(new_n6141_));
  NOR2_X1    g06070(.A1(new_n6140_), .A2(new_n6141_), .ZN(new_n6142_));
  INV_X1     g06071(.I(new_n6142_), .ZN(new_n6143_));
  XNOR2_X1   g06072(.A1(new_n5698_), .A2(new_n5711_), .ZN(new_n6144_));
  INV_X1     g06073(.I(new_n6144_), .ZN(new_n6145_));
  AOI22_X1   g06074(.A1(new_n4143_), .A2(new_n4526_), .B1(new_n4274_), .B2(new_n4570_), .ZN(new_n6146_));
  NOR2_X1    g06075(.A1(new_n4135_), .A2(new_n79_), .ZN(new_n6147_));
  OAI21_X1   g06076(.A1(new_n6147_), .A2(new_n6146_), .B(new_n72_), .ZN(new_n6148_));
  NAND2_X1   g06077(.A1(new_n6148_), .A2(new_n101_), .ZN(new_n6149_));
  XOR2_X1    g06078(.A1(new_n5624_), .A2(new_n6149_), .Z(new_n6150_));
  INV_X1     g06079(.I(new_n6150_), .ZN(new_n6151_));
  NOR2_X1    g06080(.A1(new_n6151_), .A2(new_n6145_), .ZN(new_n6152_));
  INV_X1     g06081(.I(new_n6152_), .ZN(new_n6153_));
  NOR2_X1    g06082(.A1(new_n6150_), .A2(new_n6144_), .ZN(new_n6154_));
  AOI21_X1   g06083(.A1(new_n6143_), .A2(new_n6153_), .B(new_n6154_), .ZN(new_n6155_));
  INV_X1     g06084(.I(new_n6155_), .ZN(new_n6156_));
  XOR2_X1    g06085(.A1(new_n5726_), .A2(new_n5712_), .Z(new_n6157_));
  OAI22_X1   g06086(.A1(new_n4135_), .A2(new_n4527_), .B1(new_n4142_), .B2(new_n4529_), .ZN(new_n6158_));
  OAI21_X1   g06087(.A1(new_n4285_), .A2(new_n79_), .B(new_n6158_), .ZN(new_n6159_));
  AOI21_X1   g06088(.A1(new_n6159_), .A2(new_n72_), .B(new_n79_), .ZN(new_n6160_));
  XNOR2_X1   g06089(.A1(new_n5023_), .A2(new_n6160_), .ZN(new_n6161_));
  INV_X1     g06090(.I(new_n6161_), .ZN(new_n6162_));
  NOR2_X1    g06091(.A1(new_n6162_), .A2(new_n6157_), .ZN(new_n6163_));
  INV_X1     g06092(.I(new_n6163_), .ZN(new_n6164_));
  NAND2_X1   g06093(.A1(new_n6162_), .A2(new_n6157_), .ZN(new_n6165_));
  INV_X1     g06094(.I(new_n6165_), .ZN(new_n6166_));
  AOI21_X1   g06095(.A1(new_n6156_), .A2(new_n6164_), .B(new_n6166_), .ZN(new_n6167_));
  INV_X1     g06096(.I(new_n6167_), .ZN(new_n6168_));
  NAND2_X1   g06097(.A1(new_n5727_), .A2(new_n5738_), .ZN(new_n6169_));
  INV_X1     g06098(.I(new_n6169_), .ZN(new_n6170_));
  NOR2_X1    g06099(.A1(new_n6170_), .A2(new_n5739_), .ZN(new_n6171_));
  INV_X1     g06100(.I(new_n6171_), .ZN(new_n6172_));
  AOI22_X1   g06101(.A1(new_n4290_), .A2(new_n4526_), .B1(new_n4136_), .B2(new_n4570_), .ZN(new_n6173_));
  AOI21_X1   g06102(.A1(new_n101_), .A2(new_n4297_), .B(new_n6173_), .ZN(new_n6174_));
  OAI21_X1   g06103(.A1(new_n6174_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n6175_));
  XOR2_X1    g06104(.A1(new_n5753_), .A2(new_n6175_), .Z(new_n6176_));
  INV_X1     g06105(.I(new_n6176_), .ZN(new_n6177_));
  NOR2_X1    g06106(.A1(new_n6177_), .A2(new_n6172_), .ZN(new_n6178_));
  INV_X1     g06107(.I(new_n6178_), .ZN(new_n6179_));
  NOR2_X1    g06108(.A1(new_n6176_), .A2(new_n6171_), .ZN(new_n6180_));
  AOI21_X1   g06109(.A1(new_n6168_), .A2(new_n6179_), .B(new_n6180_), .ZN(new_n6181_));
  INV_X1     g06110(.I(new_n6181_), .ZN(new_n6182_));
  INV_X1     g06111(.I(new_n5738_), .ZN(new_n6183_));
  NAND2_X1   g06112(.A1(new_n6183_), .A2(new_n5727_), .ZN(new_n6184_));
  OAI22_X1   g06113(.A1(new_n4296_), .A2(new_n4527_), .B1(new_n4285_), .B2(new_n4529_), .ZN(new_n6185_));
  OAI21_X1   g06114(.A1(new_n4131_), .A2(new_n79_), .B(new_n6185_), .ZN(new_n6186_));
  AOI21_X1   g06115(.A1(new_n6186_), .A2(new_n72_), .B(new_n79_), .ZN(new_n6187_));
  XNOR2_X1   g06116(.A1(new_n5599_), .A2(new_n6187_), .ZN(new_n6188_));
  INV_X1     g06117(.I(new_n6188_), .ZN(new_n6189_));
  NOR2_X1    g06118(.A1(new_n6189_), .A2(new_n6184_), .ZN(new_n6190_));
  INV_X1     g06119(.I(new_n6190_), .ZN(new_n6191_));
  AOI21_X1   g06120(.A1(new_n5727_), .A2(new_n6183_), .B(new_n6188_), .ZN(new_n6192_));
  AOI21_X1   g06121(.A1(new_n6182_), .A2(new_n6191_), .B(new_n6192_), .ZN(new_n6193_));
  AOI22_X1   g06122(.A1(new_n4113_), .A2(new_n4767_), .B1(new_n4124_), .B2(new_n4613_), .ZN(new_n6194_));
  AOI21_X1   g06123(.A1(new_n117_), .A2(new_n4105_), .B(new_n6194_), .ZN(new_n6195_));
  OAI21_X1   g06124(.A1(new_n6195_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n6196_));
  XOR2_X1    g06125(.A1(new_n5121_), .A2(new_n6196_), .Z(new_n6197_));
  NOR2_X1    g06126(.A1(new_n6193_), .A2(new_n6197_), .ZN(new_n6198_));
  INV_X1     g06127(.I(new_n6198_), .ZN(new_n6199_));
  XNOR2_X1   g06128(.A1(new_n5744_), .A2(new_n5740_), .ZN(new_n6200_));
  NOR2_X1    g06129(.A1(new_n6200_), .A2(new_n5615_), .ZN(new_n6201_));
  AOI21_X1   g06130(.A1(new_n5747_), .A2(new_n5745_), .B(new_n5616_), .ZN(new_n6202_));
  NOR2_X1    g06131(.A1(new_n6201_), .A2(new_n6202_), .ZN(new_n6203_));
  INV_X1     g06132(.I(new_n6203_), .ZN(new_n6204_));
  INV_X1     g06133(.I(new_n6193_), .ZN(new_n6205_));
  INV_X1     g06134(.I(new_n6197_), .ZN(new_n6206_));
  NOR2_X1    g06135(.A1(new_n6205_), .A2(new_n6206_), .ZN(new_n6207_));
  OAI21_X1   g06136(.A1(new_n6204_), .A2(new_n6207_), .B(new_n6199_), .ZN(new_n6208_));
  OAI22_X1   g06137(.A1(new_n4332_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4081_), .ZN(new_n6209_));
  AOI21_X1   g06138(.A1(new_n6209_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6210_));
  XOR2_X1    g06139(.A1(new_n5162_), .A2(new_n6210_), .Z(new_n6211_));
  INV_X1     g06140(.I(new_n6211_), .ZN(new_n6212_));
  NOR2_X1    g06141(.A1(new_n6212_), .A2(new_n6208_), .ZN(new_n6213_));
  INV_X1     g06142(.I(new_n6213_), .ZN(new_n6214_));
  NAND2_X1   g06143(.A1(new_n6212_), .A2(new_n6208_), .ZN(new_n6215_));
  INV_X1     g06144(.I(new_n6215_), .ZN(new_n6216_));
  AOI21_X1   g06145(.A1(new_n6046_), .A2(new_n6214_), .B(new_n6216_), .ZN(new_n6217_));
  OAI22_X1   g06146(.A1(new_n4042_), .A2(new_n5398_), .B1(new_n4342_), .B2(new_n5336_), .ZN(new_n6218_));
  AOI21_X1   g06147(.A1(new_n6218_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n6219_));
  XNOR2_X1   g06148(.A1(new_n4864_), .A2(new_n6219_), .ZN(new_n6220_));
  XOR2_X1    g06149(.A1(new_n5900_), .A2(new_n5916_), .Z(new_n6221_));
  XOR2_X1    g06150(.A1(new_n6220_), .A2(new_n6221_), .Z(new_n6222_));
  XOR2_X1    g06151(.A1(new_n6222_), .A2(new_n6217_), .Z(new_n6223_));
  XOR2_X1    g06152(.A1(new_n6223_), .A2(new_n6043_), .Z(new_n6224_));
  INV_X1     g06153(.I(new_n6224_), .ZN(new_n6225_));
  OAI21_X1   g06154(.A1(new_n6213_), .A2(new_n6216_), .B(new_n6046_), .ZN(new_n6226_));
  XOR2_X1    g06155(.A1(new_n6208_), .A2(new_n6211_), .Z(new_n6227_));
  OAI21_X1   g06156(.A1(new_n6046_), .A2(new_n6227_), .B(new_n6226_), .ZN(new_n6228_));
  XOR2_X1    g06157(.A1(new_n6193_), .A2(new_n6206_), .Z(new_n6229_));
  NOR2_X1    g06158(.A1(new_n6229_), .A2(new_n6203_), .ZN(new_n6230_));
  NOR2_X1    g06159(.A1(new_n6207_), .A2(new_n6198_), .ZN(new_n6231_));
  INV_X1     g06160(.I(new_n6231_), .ZN(new_n6232_));
  AOI21_X1   g06161(.A1(new_n6203_), .A2(new_n6232_), .B(new_n6230_), .ZN(new_n6233_));
  INV_X1     g06162(.I(new_n6233_), .ZN(new_n6234_));
  XOR2_X1    g06163(.A1(new_n6150_), .A2(new_n6145_), .Z(new_n6235_));
  INV_X1     g06164(.I(new_n6235_), .ZN(new_n6236_));
  NOR2_X1    g06165(.A1(new_n6152_), .A2(new_n6154_), .ZN(new_n6237_));
  NOR2_X1    g06166(.A1(new_n6143_), .A2(new_n6237_), .ZN(new_n6238_));
  AOI21_X1   g06167(.A1(new_n6143_), .A2(new_n6236_), .B(new_n6238_), .ZN(new_n6239_));
  NAND2_X1   g06168(.A1(new_n6109_), .A2(new_n6112_), .ZN(new_n6240_));
  XNOR2_X1   g06169(.A1(new_n6122_), .A2(new_n6240_), .ZN(new_n6241_));
  INV_X1     g06170(.I(new_n6241_), .ZN(new_n6242_));
  NOR4_X1    g06171(.A1(new_n5646_), .A2(new_n5645_), .A3(new_n4252_), .A4(new_n5640_), .ZN(new_n6243_));
  AOI22_X1   g06172(.A1(new_n5643_), .A2(new_n4244_), .B1(new_n5641_), .B2(new_n5642_), .ZN(new_n6244_));
  NOR2_X1    g06173(.A1(new_n6244_), .A2(new_n6243_), .ZN(new_n6245_));
  NAND2_X1   g06174(.A1(new_n4252_), .A2(new_n4613_), .ZN(new_n6246_));
  OAI21_X1   g06175(.A1(new_n4234_), .A2(new_n4781_), .B(new_n6246_), .ZN(new_n6247_));
  OAI21_X1   g06176(.A1(new_n1128_), .A2(new_n4249_), .B(new_n6247_), .ZN(new_n6248_));
  AOI21_X1   g06177(.A1(new_n6248_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n6249_));
  XOR2_X1    g06178(.A1(new_n6245_), .A2(new_n6249_), .Z(new_n6250_));
  NOR2_X1    g06179(.A1(new_n6250_), .A2(new_n6072_), .ZN(new_n6251_));
  NAND2_X1   g06180(.A1(new_n5627_), .A2(new_n1128_), .ZN(new_n6252_));
  AOI21_X1   g06181(.A1(new_n117_), .A2(new_n6061_), .B(new_n4260_), .ZN(new_n6253_));
  OAI22_X1   g06182(.A1(new_n4244_), .A2(new_n4781_), .B1(new_n4230_), .B2(new_n4612_), .ZN(new_n6254_));
  OAI21_X1   g06183(.A1(new_n1128_), .A2(new_n4234_), .B(new_n6254_), .ZN(new_n6255_));
  AOI21_X1   g06184(.A1(new_n6252_), .A2(new_n6253_), .B(new_n6255_), .ZN(new_n6256_));
  XOR2_X1    g06185(.A1(new_n6256_), .A2(\a[26] ), .Z(new_n6257_));
  AOI21_X1   g06186(.A1(new_n4251_), .A2(new_n117_), .B(\a[26] ), .ZN(new_n6258_));
  AOI21_X1   g06187(.A1(new_n6258_), .A2(new_n6246_), .B(new_n1128_), .ZN(new_n6259_));
  XNOR2_X1   g06188(.A1(new_n5637_), .A2(new_n6259_), .ZN(new_n6260_));
  NOR2_X1    g06189(.A1(new_n4251_), .A2(new_n1120_), .ZN(new_n6261_));
  NOR2_X1    g06190(.A1(new_n6261_), .A2(new_n65_), .ZN(new_n6262_));
  INV_X1     g06191(.I(new_n6262_), .ZN(new_n6263_));
  NOR2_X1    g06192(.A1(new_n6260_), .A2(new_n6263_), .ZN(new_n6264_));
  NAND2_X1   g06193(.A1(new_n6257_), .A2(new_n6264_), .ZN(new_n6265_));
  NAND2_X1   g06194(.A1(new_n6250_), .A2(new_n6072_), .ZN(new_n6266_));
  AOI21_X1   g06195(.A1(new_n6265_), .A2(new_n6266_), .B(new_n6251_), .ZN(new_n6267_));
  XOR2_X1    g06196(.A1(new_n6070_), .A2(new_n6074_), .Z(new_n6268_));
  OAI22_X1   g06197(.A1(new_n4249_), .A2(new_n4781_), .B1(new_n4234_), .B2(new_n4612_), .ZN(new_n6269_));
  OAI21_X1   g06198(.A1(new_n4203_), .A2(new_n1128_), .B(new_n6269_), .ZN(new_n6270_));
  AOI21_X1   g06199(.A1(new_n6270_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n6271_));
  XOR2_X1    g06200(.A1(new_n5660_), .A2(new_n6271_), .Z(new_n6272_));
  NOR2_X1    g06201(.A1(new_n6272_), .A2(new_n6268_), .ZN(new_n6273_));
  NOR2_X1    g06202(.A1(new_n6273_), .A2(new_n6267_), .ZN(new_n6274_));
  INV_X1     g06203(.I(new_n6268_), .ZN(new_n6275_));
  XOR2_X1    g06204(.A1(new_n6082_), .A2(new_n6271_), .Z(new_n6276_));
  NOR2_X1    g06205(.A1(new_n6276_), .A2(new_n6275_), .ZN(new_n6277_));
  NOR2_X1    g06206(.A1(new_n6274_), .A2(new_n6277_), .ZN(new_n6278_));
  NOR2_X1    g06207(.A1(new_n6071_), .A2(new_n6074_), .ZN(new_n6279_));
  XOR2_X1    g06208(.A1(new_n6279_), .A2(new_n6066_), .Z(new_n6280_));
  OAI22_X1   g06209(.A1(new_n4203_), .A2(new_n4781_), .B1(new_n4249_), .B2(new_n4612_), .ZN(new_n6281_));
  OAI21_X1   g06210(.A1(new_n1128_), .A2(new_n4175_), .B(new_n6281_), .ZN(new_n6282_));
  AOI21_X1   g06211(.A1(new_n6282_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n6283_));
  XOR2_X1    g06212(.A1(new_n5671_), .A2(new_n6283_), .Z(new_n6284_));
  NOR2_X1    g06213(.A1(new_n6284_), .A2(new_n6280_), .ZN(new_n6285_));
  NAND2_X1   g06214(.A1(new_n6284_), .A2(new_n6280_), .ZN(new_n6286_));
  OAI21_X1   g06215(.A1(new_n6278_), .A2(new_n6285_), .B(new_n6286_), .ZN(new_n6287_));
  INV_X1     g06216(.I(new_n6075_), .ZN(new_n6288_));
  INV_X1     g06217(.I(new_n6076_), .ZN(new_n6289_));
  AOI21_X1   g06218(.A1(new_n6059_), .A2(new_n6289_), .B(new_n6288_), .ZN(new_n6290_));
  XOR2_X1    g06219(.A1(new_n6058_), .A2(new_n6052_), .Z(new_n6291_));
  NOR2_X1    g06220(.A1(new_n6291_), .A2(new_n6075_), .ZN(new_n6292_));
  OAI22_X1   g06221(.A1(new_n4175_), .A2(new_n4781_), .B1(new_n4203_), .B2(new_n4612_), .ZN(new_n6293_));
  OAI21_X1   g06222(.A1(new_n1128_), .A2(new_n5684_), .B(new_n6293_), .ZN(new_n6294_));
  AOI21_X1   g06223(.A1(new_n6294_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n6295_));
  XOR2_X1    g06224(.A1(new_n6102_), .A2(new_n6295_), .Z(new_n6296_));
  OAI21_X1   g06225(.A1(new_n6290_), .A2(new_n6292_), .B(new_n6296_), .ZN(new_n6297_));
  NAND2_X1   g06226(.A1(new_n6297_), .A2(new_n6287_), .ZN(new_n6298_));
  OR3_X2     g06227(.A1(new_n6296_), .A2(new_n6290_), .A3(new_n6292_), .Z(new_n6299_));
  NAND2_X1   g06228(.A1(new_n6298_), .A2(new_n6299_), .ZN(new_n6300_));
  INV_X1     g06229(.I(new_n6088_), .ZN(new_n6301_));
  NAND2_X1   g06230(.A1(new_n6301_), .A2(new_n6087_), .ZN(new_n6302_));
  NAND2_X1   g06231(.A1(new_n6302_), .A2(new_n6077_), .ZN(new_n6303_));
  XOR2_X1    g06232(.A1(new_n6086_), .A2(new_n6094_), .Z(new_n6304_));
  OAI21_X1   g06233(.A1(new_n6304_), .A2(new_n6077_), .B(new_n6303_), .ZN(new_n6305_));
  OAI22_X1   g06234(.A1(new_n5684_), .A2(new_n4781_), .B1(new_n4175_), .B2(new_n4612_), .ZN(new_n6306_));
  OAI21_X1   g06235(.A1(new_n4150_), .A2(new_n1128_), .B(new_n6306_), .ZN(new_n6307_));
  AOI21_X1   g06236(.A1(new_n6307_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n6308_));
  XNOR2_X1   g06237(.A1(new_n5707_), .A2(new_n6308_), .ZN(new_n6309_));
  OR2_X2     g06238(.A1(new_n6305_), .A2(new_n6309_), .Z(new_n6310_));
  NAND2_X1   g06239(.A1(new_n6310_), .A2(new_n6300_), .ZN(new_n6311_));
  NAND2_X1   g06240(.A1(new_n6305_), .A2(new_n6309_), .ZN(new_n6312_));
  NAND2_X1   g06241(.A1(new_n6311_), .A2(new_n6312_), .ZN(new_n6313_));
  XOR2_X1    g06242(.A1(new_n6093_), .A2(new_n6096_), .Z(new_n6314_));
  INV_X1     g06243(.I(new_n6314_), .ZN(new_n6315_));
  INV_X1     g06244(.I(new_n6098_), .ZN(new_n6316_));
  OAI21_X1   g06245(.A1(new_n6316_), .A2(new_n6097_), .B(new_n6089_), .ZN(new_n6317_));
  OAI21_X1   g06246(.A1(new_n6315_), .A2(new_n6089_), .B(new_n6317_), .ZN(new_n6318_));
  AOI22_X1   g06247(.A1(new_n5701_), .A2(new_n4767_), .B1(new_n4171_), .B2(new_n4613_), .ZN(new_n6319_));
  AOI21_X1   g06248(.A1(new_n117_), .A2(new_n4274_), .B(new_n6319_), .ZN(new_n6320_));
  OAI21_X1   g06249(.A1(new_n6320_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n6321_));
  XOR2_X1    g06250(.A1(new_n5722_), .A2(new_n6321_), .Z(new_n6322_));
  NOR2_X1    g06251(.A1(new_n6322_), .A2(new_n6318_), .ZN(new_n6323_));
  NAND2_X1   g06252(.A1(new_n6322_), .A2(new_n6318_), .ZN(new_n6324_));
  INV_X1     g06253(.I(new_n6324_), .ZN(new_n6325_));
  XOR2_X1    g06254(.A1(new_n6110_), .A2(new_n6111_), .Z(new_n6326_));
  AOI21_X1   g06255(.A1(new_n6108_), .A2(new_n6112_), .B(new_n6099_), .ZN(new_n6327_));
  AOI21_X1   g06256(.A1(new_n6326_), .A2(new_n6099_), .B(new_n6327_), .ZN(new_n6328_));
  OAI22_X1   g06257(.A1(new_n4273_), .A2(new_n4781_), .B1(new_n4150_), .B2(new_n4612_), .ZN(new_n6329_));
  OAI21_X1   g06258(.A1(new_n1128_), .A2(new_n4142_), .B(new_n6329_), .ZN(new_n6330_));
  AOI21_X1   g06259(.A1(new_n6330_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n6331_));
  XOR2_X1    g06260(.A1(new_n6134_), .A2(new_n6331_), .Z(new_n6332_));
  XNOR2_X1   g06261(.A1(new_n6328_), .A2(new_n6332_), .ZN(new_n6333_));
  OAI21_X1   g06262(.A1(new_n6323_), .A2(new_n6325_), .B(new_n6313_), .ZN(new_n6334_));
  NOR2_X1    g06263(.A1(new_n6334_), .A2(new_n6242_), .ZN(new_n6335_));
  INV_X1     g06264(.I(new_n6332_), .ZN(new_n6336_));
  NOR2_X1    g06265(.A1(new_n6336_), .A2(new_n6328_), .ZN(new_n6337_));
  AOI22_X1   g06266(.A1(new_n4143_), .A2(new_n4767_), .B1(new_n4274_), .B2(new_n4613_), .ZN(new_n6338_));
  NOR2_X1    g06267(.A1(new_n4135_), .A2(new_n1128_), .ZN(new_n6339_));
  OAI21_X1   g06268(.A1(new_n6339_), .A2(new_n6338_), .B(new_n65_), .ZN(new_n6340_));
  NAND2_X1   g06269(.A1(new_n6340_), .A2(new_n117_), .ZN(new_n6341_));
  XNOR2_X1   g06270(.A1(new_n5624_), .A2(new_n6341_), .ZN(new_n6342_));
  NAND2_X1   g06271(.A1(new_n6342_), .A2(new_n6337_), .ZN(new_n6343_));
  AOI21_X1   g06272(.A1(new_n6334_), .A2(new_n6242_), .B(new_n6343_), .ZN(new_n6344_));
  NOR2_X1    g06273(.A1(new_n6344_), .A2(new_n6335_), .ZN(new_n6345_));
  INV_X1     g06274(.I(new_n6345_), .ZN(new_n6346_));
  NOR2_X1    g06275(.A1(new_n6051_), .A2(new_n6125_), .ZN(new_n6347_));
  XOR2_X1    g06276(.A1(new_n6347_), .A2(new_n6123_), .Z(new_n6348_));
  XOR2_X1    g06277(.A1(new_n6348_), .A2(new_n6119_), .Z(new_n6349_));
  OAI22_X1   g06278(.A1(new_n4135_), .A2(new_n4781_), .B1(new_n4142_), .B2(new_n4612_), .ZN(new_n6350_));
  OAI21_X1   g06279(.A1(new_n4285_), .A2(new_n1128_), .B(new_n6350_), .ZN(new_n6351_));
  AOI21_X1   g06280(.A1(new_n6351_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n6352_));
  XNOR2_X1   g06281(.A1(new_n5023_), .A2(new_n6352_), .ZN(new_n6353_));
  NAND2_X1   g06282(.A1(new_n6349_), .A2(new_n6353_), .ZN(new_n6354_));
  NOR2_X1    g06283(.A1(new_n6349_), .A2(new_n6353_), .ZN(new_n6355_));
  AOI21_X1   g06284(.A1(new_n6346_), .A2(new_n6354_), .B(new_n6355_), .ZN(new_n6356_));
  XNOR2_X1   g06285(.A1(new_n6138_), .A2(new_n6131_), .ZN(new_n6357_));
  OAI21_X1   g06286(.A1(new_n6139_), .A2(new_n6141_), .B(new_n6129_), .ZN(new_n6358_));
  OAI21_X1   g06287(.A1(new_n6129_), .A2(new_n6357_), .B(new_n6358_), .ZN(new_n6359_));
  AOI22_X1   g06288(.A1(new_n4290_), .A2(new_n4767_), .B1(new_n4136_), .B2(new_n4613_), .ZN(new_n6360_));
  AOI21_X1   g06289(.A1(new_n117_), .A2(new_n4297_), .B(new_n6360_), .ZN(new_n6361_));
  OAI21_X1   g06290(.A1(new_n6361_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n6362_));
  XOR2_X1    g06291(.A1(new_n5753_), .A2(new_n6362_), .Z(new_n6363_));
  NOR2_X1    g06292(.A1(new_n6359_), .A2(new_n6363_), .ZN(new_n6364_));
  NAND2_X1   g06293(.A1(new_n6359_), .A2(new_n6363_), .ZN(new_n6365_));
  INV_X1     g06294(.I(new_n6365_), .ZN(new_n6366_));
  NOR2_X1    g06295(.A1(new_n6366_), .A2(new_n6364_), .ZN(new_n6367_));
  NAND2_X1   g06296(.A1(new_n6367_), .A2(new_n6356_), .ZN(new_n6368_));
  NAND2_X1   g06297(.A1(new_n6368_), .A2(new_n6239_), .ZN(new_n6369_));
  OAI22_X1   g06298(.A1(new_n4296_), .A2(new_n4781_), .B1(new_n4285_), .B2(new_n4612_), .ZN(new_n6370_));
  OAI21_X1   g06299(.A1(new_n4131_), .A2(new_n1128_), .B(new_n6370_), .ZN(new_n6371_));
  AOI21_X1   g06300(.A1(new_n6371_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n6372_));
  XNOR2_X1   g06301(.A1(new_n5599_), .A2(new_n6372_), .ZN(new_n6373_));
  NOR2_X1    g06302(.A1(new_n6373_), .A2(new_n6365_), .ZN(new_n6374_));
  NAND2_X1   g06303(.A1(new_n6369_), .A2(new_n6374_), .ZN(new_n6375_));
  OAI21_X1   g06304(.A1(new_n6239_), .A2(new_n6368_), .B(new_n6375_), .ZN(new_n6376_));
  XOR2_X1    g06305(.A1(new_n6161_), .A2(new_n6157_), .Z(new_n6377_));
  NOR2_X1    g06306(.A1(new_n6155_), .A2(new_n6377_), .ZN(new_n6378_));
  AOI21_X1   g06307(.A1(new_n6164_), .A2(new_n6165_), .B(new_n6156_), .ZN(new_n6379_));
  NOR2_X1    g06308(.A1(new_n6379_), .A2(new_n6378_), .ZN(new_n6380_));
  OAI22_X1   g06309(.A1(new_n4131_), .A2(new_n4781_), .B1(new_n4296_), .B2(new_n4612_), .ZN(new_n6381_));
  OAI21_X1   g06310(.A1(new_n1128_), .A2(new_n4309_), .B(new_n6381_), .ZN(new_n6382_));
  AOI21_X1   g06311(.A1(new_n6382_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n6383_));
  XNOR2_X1   g06312(.A1(new_n5049_), .A2(new_n6383_), .ZN(new_n6384_));
  INV_X1     g06313(.I(new_n6384_), .ZN(new_n6385_));
  NOR2_X1    g06314(.A1(new_n6380_), .A2(new_n6385_), .ZN(new_n6386_));
  INV_X1     g06315(.I(new_n6386_), .ZN(new_n6387_));
  NOR3_X1    g06316(.A1(new_n6384_), .A2(new_n6379_), .A3(new_n6378_), .ZN(new_n6388_));
  AOI21_X1   g06317(.A1(new_n6376_), .A2(new_n6387_), .B(new_n6388_), .ZN(new_n6389_));
  INV_X1     g06318(.I(new_n6389_), .ZN(new_n6390_));
  XOR2_X1    g06319(.A1(new_n6176_), .A2(new_n6172_), .Z(new_n6391_));
  OAI21_X1   g06320(.A1(new_n6178_), .A2(new_n6180_), .B(new_n6167_), .ZN(new_n6392_));
  OAI21_X1   g06321(.A1(new_n6167_), .A2(new_n6391_), .B(new_n6392_), .ZN(new_n6393_));
  INV_X1     g06322(.I(new_n6393_), .ZN(new_n6394_));
  OAI22_X1   g06323(.A1(new_n4131_), .A2(new_n4612_), .B1(new_n4309_), .B2(new_n4781_), .ZN(new_n6395_));
  OAI21_X1   g06324(.A1(new_n1128_), .A2(new_n4123_), .B(new_n6395_), .ZN(new_n6396_));
  AOI21_X1   g06325(.A1(new_n6396_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n6397_));
  XOR2_X1    g06326(.A1(new_n5906_), .A2(new_n6397_), .Z(new_n6398_));
  INV_X1     g06327(.I(new_n6398_), .ZN(new_n6399_));
  NOR2_X1    g06328(.A1(new_n6394_), .A2(new_n6399_), .ZN(new_n6400_));
  INV_X1     g06329(.I(new_n6400_), .ZN(new_n6401_));
  NOR2_X1    g06330(.A1(new_n6393_), .A2(new_n6398_), .ZN(new_n6402_));
  AOI21_X1   g06331(.A1(new_n6390_), .A2(new_n6401_), .B(new_n6402_), .ZN(new_n6403_));
  INV_X1     g06332(.I(new_n6403_), .ZN(new_n6404_));
  XOR2_X1    g06333(.A1(new_n6188_), .A2(new_n6184_), .Z(new_n6405_));
  OAI21_X1   g06334(.A1(new_n6190_), .A2(new_n6192_), .B(new_n6181_), .ZN(new_n6406_));
  OAI21_X1   g06335(.A1(new_n6181_), .A2(new_n6405_), .B(new_n6406_), .ZN(new_n6407_));
  INV_X1     g06336(.I(new_n6407_), .ZN(new_n6408_));
  OAI22_X1   g06337(.A1(new_n4123_), .A2(new_n4781_), .B1(new_n4309_), .B2(new_n4612_), .ZN(new_n6409_));
  OAI21_X1   g06338(.A1(new_n4112_), .A2(new_n1128_), .B(new_n6409_), .ZN(new_n6410_));
  AOI21_X1   g06339(.A1(new_n6410_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n6411_));
  XOR2_X1    g06340(.A1(new_n5096_), .A2(new_n6411_), .Z(new_n6412_));
  INV_X1     g06341(.I(new_n6412_), .ZN(new_n6413_));
  NOR2_X1    g06342(.A1(new_n6408_), .A2(new_n6413_), .ZN(new_n6414_));
  INV_X1     g06343(.I(new_n6414_), .ZN(new_n6415_));
  NOR2_X1    g06344(.A1(new_n6407_), .A2(new_n6412_), .ZN(new_n6416_));
  AOI21_X1   g06345(.A1(new_n6404_), .A2(new_n6415_), .B(new_n6416_), .ZN(new_n6417_));
  INV_X1     g06346(.I(new_n6417_), .ZN(new_n6418_));
  INV_X1     g06347(.I(new_n4323_), .ZN(new_n6419_));
  AOI22_X1   g06348(.A1(new_n6419_), .A2(new_n5783_), .B1(new_n247_), .B2(new_n4328_), .ZN(new_n6420_));
  OAI21_X1   g06349(.A1(new_n6420_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n6421_));
  XNOR2_X1   g06350(.A1(new_n5139_), .A2(new_n6421_), .ZN(new_n6422_));
  INV_X1     g06351(.I(new_n6422_), .ZN(new_n6423_));
  NOR2_X1    g06352(.A1(new_n6418_), .A2(new_n6423_), .ZN(new_n6424_));
  INV_X1     g06353(.I(new_n6424_), .ZN(new_n6425_));
  NOR2_X1    g06354(.A1(new_n6417_), .A2(new_n6422_), .ZN(new_n6426_));
  AOI21_X1   g06355(.A1(new_n6425_), .A2(new_n6234_), .B(new_n6426_), .ZN(new_n6427_));
  INV_X1     g06356(.I(new_n4339_), .ZN(new_n6428_));
  AOI22_X1   g06357(.A1(new_n6428_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4054_), .ZN(new_n6429_));
  OAI21_X1   g06358(.A1(new_n6429_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n6430_));
  XOR2_X1    g06359(.A1(new_n4652_), .A2(new_n6430_), .Z(new_n6431_));
  AND2_X2    g06360(.A1(new_n6431_), .A2(new_n6427_), .Z(new_n6432_));
  INV_X1     g06361(.I(new_n6432_), .ZN(new_n6433_));
  NOR2_X1    g06362(.A1(new_n6431_), .A2(new_n6427_), .ZN(new_n6434_));
  AOI21_X1   g06363(.A1(new_n6433_), .A2(new_n6228_), .B(new_n6434_), .ZN(new_n6435_));
  INV_X1     g06364(.I(new_n6435_), .ZN(new_n6436_));
  OAI22_X1   g06365(.A1(new_n4028_), .A2(new_n5419_), .B1(new_n1622_), .B2(new_n4035_), .ZN(new_n6437_));
  OAI21_X1   g06366(.A1(new_n4017_), .A2(new_n1620_), .B(new_n6437_), .ZN(new_n6438_));
  AOI21_X1   g06367(.A1(new_n6438_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n6439_));
  XNOR2_X1   g06368(.A1(new_n4705_), .A2(new_n6439_), .ZN(new_n6440_));
  INV_X1     g06369(.I(new_n6440_), .ZN(new_n6441_));
  NOR2_X1    g06370(.A1(new_n6441_), .A2(new_n6436_), .ZN(new_n6442_));
  INV_X1     g06371(.I(new_n6442_), .ZN(new_n6443_));
  NOR2_X1    g06372(.A1(new_n6440_), .A2(new_n6435_), .ZN(new_n6444_));
  AOI21_X1   g06373(.A1(new_n6225_), .A2(new_n6443_), .B(new_n6444_), .ZN(new_n6445_));
  AOI22_X1   g06374(.A1(new_n5859_), .A2(new_n5421_), .B1(new_n4375_), .B2(new_n4660_), .ZN(new_n6446_));
  OAI21_X1   g06375(.A1(new_n6446_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n6447_));
  XOR2_X1    g06376(.A1(new_n4730_), .A2(new_n6447_), .Z(new_n6448_));
  NOR2_X1    g06377(.A1(new_n6445_), .A2(new_n6448_), .ZN(new_n6449_));
  AOI22_X1   g06378(.A1(new_n4347_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4036_), .ZN(new_n6450_));
  OAI21_X1   g06379(.A1(new_n6450_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n6451_));
  XOR2_X1    g06380(.A1(new_n4672_), .A2(new_n6451_), .Z(new_n6452_));
  NOR2_X1    g06381(.A1(new_n6220_), .A2(new_n6217_), .ZN(new_n6453_));
  XOR2_X1    g06382(.A1(new_n6221_), .A2(new_n6043_), .Z(new_n6454_));
  AOI21_X1   g06383(.A1(new_n6220_), .A2(new_n6217_), .B(new_n6454_), .ZN(new_n6455_));
  NOR2_X1    g06384(.A1(new_n6455_), .A2(new_n6453_), .ZN(new_n6456_));
  XOR2_X1    g06385(.A1(new_n5930_), .A2(new_n5926_), .Z(new_n6457_));
  XNOR2_X1   g06386(.A1(new_n6457_), .A2(new_n5923_), .ZN(new_n6458_));
  XNOR2_X1   g06387(.A1(new_n6458_), .A2(new_n6456_), .ZN(new_n6459_));
  XNOR2_X1   g06388(.A1(new_n6459_), .A2(new_n6452_), .ZN(new_n6460_));
  INV_X1     g06389(.I(new_n6445_), .ZN(new_n6461_));
  INV_X1     g06390(.I(new_n6448_), .ZN(new_n6462_));
  NOR2_X1    g06391(.A1(new_n6461_), .A2(new_n6462_), .ZN(new_n6463_));
  INV_X1     g06392(.I(new_n6463_), .ZN(new_n6464_));
  AOI21_X1   g06393(.A1(new_n6464_), .A2(new_n6460_), .B(new_n6449_), .ZN(new_n6465_));
  OAI21_X1   g06394(.A1(new_n5940_), .A2(new_n5942_), .B(new_n5896_), .ZN(new_n6466_));
  XOR2_X1    g06395(.A1(new_n5938_), .A2(new_n5934_), .Z(new_n6467_));
  OAI21_X1   g06396(.A1(new_n5896_), .A2(new_n6467_), .B(new_n6466_), .ZN(new_n6468_));
  NOR2_X1    g06397(.A1(new_n6456_), .A2(new_n6452_), .ZN(new_n6469_));
  AOI21_X1   g06398(.A1(new_n6452_), .A2(new_n6456_), .B(new_n6458_), .ZN(new_n6470_));
  NOR2_X1    g06399(.A1(new_n6470_), .A2(new_n6469_), .ZN(new_n6471_));
  XOR2_X1    g06400(.A1(new_n6468_), .A2(new_n6471_), .Z(new_n6472_));
  AOI22_X1   g06401(.A1(new_n4473_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4555_), .ZN(new_n6473_));
  OAI21_X1   g06402(.A1(new_n6473_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n6474_));
  NOR2_X1    g06403(.A1(new_n4585_), .A2(new_n6474_), .ZN(new_n6475_));
  INV_X1     g06404(.I(new_n6475_), .ZN(new_n6476_));
  NAND2_X1   g06405(.A1(new_n4585_), .A2(new_n6474_), .ZN(new_n6477_));
  NAND2_X1   g06406(.A1(new_n6476_), .A2(new_n6477_), .ZN(new_n6478_));
  XOR2_X1    g06407(.A1(new_n6478_), .A2(new_n6472_), .Z(new_n6479_));
  XOR2_X1    g06408(.A1(new_n6479_), .A2(new_n6465_), .Z(new_n6480_));
  XOR2_X1    g06409(.A1(new_n6480_), .A2(new_n6042_), .Z(new_n6481_));
  OAI21_X1   g06410(.A1(new_n6442_), .A2(new_n6444_), .B(new_n6225_), .ZN(new_n6482_));
  XOR2_X1    g06411(.A1(new_n6440_), .A2(new_n6436_), .Z(new_n6483_));
  OAI21_X1   g06412(.A1(new_n6225_), .A2(new_n6483_), .B(new_n6482_), .ZN(new_n6484_));
  NOR2_X1    g06413(.A1(new_n6424_), .A2(new_n6426_), .ZN(new_n6485_));
  NOR2_X1    g06414(.A1(new_n6485_), .A2(new_n6233_), .ZN(new_n6486_));
  XOR2_X1    g06415(.A1(new_n6417_), .A2(new_n6423_), .Z(new_n6487_));
  NOR2_X1    g06416(.A1(new_n6487_), .A2(new_n6234_), .ZN(new_n6488_));
  NOR2_X1    g06417(.A1(new_n6486_), .A2(new_n6488_), .ZN(new_n6489_));
  XOR2_X1    g06418(.A1(new_n6407_), .A2(new_n6413_), .Z(new_n6490_));
  OAI21_X1   g06419(.A1(new_n6414_), .A2(new_n6416_), .B(new_n6403_), .ZN(new_n6491_));
  OAI21_X1   g06420(.A1(new_n6403_), .A2(new_n6490_), .B(new_n6491_), .ZN(new_n6492_));
  INV_X1     g06421(.I(new_n6492_), .ZN(new_n6493_));
  NOR2_X1    g06422(.A1(new_n6239_), .A2(new_n6373_), .ZN(new_n6494_));
  NAND2_X1   g06423(.A1(new_n6368_), .A2(new_n6494_), .ZN(new_n6495_));
  INV_X1     g06424(.I(new_n6495_), .ZN(new_n6496_));
  NOR2_X1    g06425(.A1(new_n6368_), .A2(new_n6494_), .ZN(new_n6497_));
  NOR2_X1    g06426(.A1(new_n6496_), .A2(new_n6497_), .ZN(new_n6498_));
  NOR2_X1    g06427(.A1(new_n6498_), .A2(new_n6366_), .ZN(new_n6499_));
  NOR3_X1    g06428(.A1(new_n6496_), .A2(new_n6365_), .A3(new_n6497_), .ZN(new_n6500_));
  NOR2_X1    g06429(.A1(new_n6499_), .A2(new_n6500_), .ZN(new_n6501_));
  NOR2_X1    g06430(.A1(new_n6325_), .A2(new_n6323_), .ZN(new_n6502_));
  XOR2_X1    g06431(.A1(new_n6502_), .A2(new_n6313_), .Z(new_n6503_));
  NOR2_X1    g06432(.A1(new_n4234_), .A2(new_n4244_), .ZN(new_n6504_));
  OAI22_X1   g06433(.A1(new_n6504_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4249_), .ZN(new_n6505_));
  NAND2_X1   g06434(.A1(new_n6505_), .A2(new_n68_), .ZN(new_n6506_));
  NAND2_X1   g06435(.A1(new_n6506_), .A2(new_n247_), .ZN(new_n6507_));
  XOR2_X1    g06436(.A1(new_n6507_), .A2(new_n5648_), .Z(new_n6508_));
  NOR2_X1    g06437(.A1(new_n6508_), .A2(new_n6261_), .ZN(new_n6509_));
  NAND2_X1   g06438(.A1(new_n5627_), .A2(new_n1239_), .ZN(new_n6510_));
  AOI21_X1   g06439(.A1(new_n247_), .A2(new_n6061_), .B(new_n4260_), .ZN(new_n6511_));
  OAI22_X1   g06440(.A1(new_n4244_), .A2(new_n4902_), .B1(new_n1973_), .B2(new_n4230_), .ZN(new_n6512_));
  OAI21_X1   g06441(.A1(new_n1239_), .A2(new_n4234_), .B(new_n6512_), .ZN(new_n6513_));
  AOI21_X1   g06442(.A1(new_n6510_), .A2(new_n6511_), .B(new_n6513_), .ZN(new_n6514_));
  XOR2_X1    g06443(.A1(new_n6514_), .A2(new_n68_), .Z(new_n6515_));
  NOR2_X1    g06444(.A1(new_n4244_), .A2(new_n1973_), .ZN(new_n6516_));
  OAI21_X1   g06445(.A1(new_n4230_), .A2(new_n1239_), .B(new_n68_), .ZN(new_n6517_));
  OAI21_X1   g06446(.A1(new_n6516_), .A2(new_n6517_), .B(new_n247_), .ZN(new_n6518_));
  XNOR2_X1   g06447(.A1(new_n6518_), .A2(new_n5637_), .ZN(new_n6519_));
  NOR2_X1    g06448(.A1(new_n4251_), .A2(new_n1121_), .ZN(new_n6520_));
  NOR2_X1    g06449(.A1(new_n6520_), .A2(new_n68_), .ZN(new_n6521_));
  NAND2_X1   g06450(.A1(new_n6519_), .A2(new_n6521_), .ZN(new_n6522_));
  NOR2_X1    g06451(.A1(new_n6515_), .A2(new_n6522_), .ZN(new_n6523_));
  INV_X1     g06452(.I(new_n6523_), .ZN(new_n6524_));
  NAND2_X1   g06453(.A1(new_n6508_), .A2(new_n6261_), .ZN(new_n6525_));
  AOI21_X1   g06454(.A1(new_n6524_), .A2(new_n6525_), .B(new_n6509_), .ZN(new_n6526_));
  XOR2_X1    g06455(.A1(new_n6260_), .A2(new_n6263_), .Z(new_n6527_));
  INV_X1     g06456(.I(new_n6527_), .ZN(new_n6528_));
  NOR2_X1    g06457(.A1(new_n4249_), .A2(new_n4234_), .ZN(new_n6529_));
  OAI22_X1   g06458(.A1(new_n4203_), .A2(new_n1239_), .B1(new_n4981_), .B2(new_n6529_), .ZN(new_n6530_));
  AOI21_X1   g06459(.A1(new_n6530_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6531_));
  XOR2_X1    g06460(.A1(new_n5660_), .A2(new_n6531_), .Z(new_n6532_));
  NOR2_X1    g06461(.A1(new_n6532_), .A2(new_n6528_), .ZN(new_n6533_));
  NOR2_X1    g06462(.A1(new_n6533_), .A2(new_n6526_), .ZN(new_n6534_));
  XOR2_X1    g06463(.A1(new_n6082_), .A2(new_n6531_), .Z(new_n6535_));
  NOR2_X1    g06464(.A1(new_n6535_), .A2(new_n6527_), .ZN(new_n6536_));
  NOR2_X1    g06465(.A1(new_n6534_), .A2(new_n6536_), .ZN(new_n6537_));
  XNOR2_X1   g06466(.A1(new_n6257_), .A2(new_n6264_), .ZN(new_n6538_));
  INV_X1     g06467(.I(new_n6538_), .ZN(new_n6539_));
  AOI21_X1   g06468(.A1(new_n5679_), .A2(new_n4175_), .B(new_n5666_), .ZN(new_n6540_));
  NAND2_X1   g06469(.A1(new_n5655_), .A2(new_n4221_), .ZN(new_n6541_));
  INV_X1     g06470(.I(new_n6541_), .ZN(new_n6542_));
  OAI22_X1   g06471(.A1(new_n6542_), .A2(new_n4981_), .B1(new_n4175_), .B2(new_n1239_), .ZN(new_n6543_));
  AOI21_X1   g06472(.A1(new_n6543_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6544_));
  XOR2_X1    g06473(.A1(new_n6540_), .A2(new_n6544_), .Z(new_n6545_));
  NAND2_X1   g06474(.A1(new_n6545_), .A2(new_n6539_), .ZN(new_n6546_));
  INV_X1     g06475(.I(new_n6546_), .ZN(new_n6547_));
  XOR2_X1    g06476(.A1(new_n5671_), .A2(new_n6544_), .Z(new_n6548_));
  NAND2_X1   g06477(.A1(new_n6548_), .A2(new_n6538_), .ZN(new_n6549_));
  OAI21_X1   g06478(.A1(new_n6537_), .A2(new_n6547_), .B(new_n6549_), .ZN(new_n6550_));
  INV_X1     g06479(.I(new_n6265_), .ZN(new_n6551_));
  XOR2_X1    g06480(.A1(new_n6250_), .A2(new_n6072_), .Z(new_n6552_));
  INV_X1     g06481(.I(new_n6251_), .ZN(new_n6553_));
  AOI21_X1   g06482(.A1(new_n6553_), .A2(new_n6266_), .B(new_n6551_), .ZN(new_n6554_));
  AOI21_X1   g06483(.A1(new_n6552_), .A2(new_n6551_), .B(new_n6554_), .ZN(new_n6555_));
  NOR2_X1    g06484(.A1(new_n4175_), .A2(new_n4203_), .ZN(new_n6556_));
  OAI22_X1   g06485(.A1(new_n5684_), .A2(new_n1239_), .B1(new_n6556_), .B2(new_n4981_), .ZN(new_n6557_));
  AOI21_X1   g06486(.A1(new_n6557_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6558_));
  XOR2_X1    g06487(.A1(new_n6102_), .A2(new_n6558_), .Z(new_n6559_));
  NAND2_X1   g06488(.A1(new_n6559_), .A2(new_n6555_), .ZN(new_n6560_));
  NAND2_X1   g06489(.A1(new_n6560_), .A2(new_n6550_), .ZN(new_n6561_));
  OR2_X2     g06490(.A1(new_n6559_), .A2(new_n6555_), .Z(new_n6562_));
  XOR2_X1    g06491(.A1(new_n6272_), .A2(new_n6275_), .Z(new_n6563_));
  OAI21_X1   g06492(.A1(new_n6277_), .A2(new_n6273_), .B(new_n6267_), .ZN(new_n6564_));
  OAI21_X1   g06493(.A1(new_n6563_), .A2(new_n6267_), .B(new_n6564_), .ZN(new_n6565_));
  INV_X1     g06494(.I(new_n6565_), .ZN(new_n6566_));
  NOR2_X1    g06495(.A1(new_n5684_), .A2(new_n4175_), .ZN(new_n6567_));
  OAI22_X1   g06496(.A1(new_n4150_), .A2(new_n1239_), .B1(new_n6567_), .B2(new_n4981_), .ZN(new_n6568_));
  AOI21_X1   g06497(.A1(new_n6568_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6569_));
  XNOR2_X1   g06498(.A1(new_n5707_), .A2(new_n6569_), .ZN(new_n6570_));
  NOR2_X1    g06499(.A1(new_n6566_), .A2(new_n6570_), .ZN(new_n6571_));
  AOI21_X1   g06500(.A1(new_n6561_), .A2(new_n6562_), .B(new_n6571_), .ZN(new_n6572_));
  INV_X1     g06501(.I(new_n6570_), .ZN(new_n6573_));
  NOR2_X1    g06502(.A1(new_n6573_), .A2(new_n6565_), .ZN(new_n6574_));
  NOR2_X1    g06503(.A1(new_n6572_), .A2(new_n6574_), .ZN(new_n6575_));
  XNOR2_X1   g06504(.A1(new_n6284_), .A2(new_n6280_), .ZN(new_n6576_));
  NOR2_X1    g06505(.A1(new_n6576_), .A2(new_n6278_), .ZN(new_n6577_));
  INV_X1     g06506(.I(new_n6285_), .ZN(new_n6578_));
  NAND2_X1   g06507(.A1(new_n6578_), .A2(new_n6286_), .ZN(new_n6579_));
  AND2_X2    g06508(.A1(new_n6579_), .A2(new_n6278_), .Z(new_n6580_));
  NOR2_X1    g06509(.A1(new_n6580_), .A2(new_n6577_), .ZN(new_n6581_));
  NAND2_X1   g06510(.A1(new_n5701_), .A2(new_n4171_), .ZN(new_n6582_));
  AOI22_X1   g06511(.A1(new_n6582_), .A2(new_n5783_), .B1(new_n247_), .B2(new_n4274_), .ZN(new_n6583_));
  OAI21_X1   g06512(.A1(new_n6583_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n6584_));
  XOR2_X1    g06513(.A1(new_n5722_), .A2(new_n6584_), .Z(new_n6585_));
  INV_X1     g06514(.I(new_n6585_), .ZN(new_n6586_));
  NOR2_X1    g06515(.A1(new_n6586_), .A2(new_n6581_), .ZN(new_n6587_));
  NAND2_X1   g06516(.A1(new_n6586_), .A2(new_n6581_), .ZN(new_n6588_));
  OAI21_X1   g06517(.A1(new_n6575_), .A2(new_n6587_), .B(new_n6588_), .ZN(new_n6589_));
  INV_X1     g06518(.I(new_n6287_), .ZN(new_n6590_));
  NOR2_X1    g06519(.A1(new_n6292_), .A2(new_n6290_), .ZN(new_n6591_));
  XOR2_X1    g06520(.A1(new_n6296_), .A2(new_n6591_), .Z(new_n6592_));
  NOR2_X1    g06521(.A1(new_n6592_), .A2(new_n6590_), .ZN(new_n6593_));
  AOI21_X1   g06522(.A1(new_n6299_), .A2(new_n6297_), .B(new_n6287_), .ZN(new_n6594_));
  OAI22_X1   g06523(.A1(new_n4142_), .A2(new_n1239_), .B1(new_n4277_), .B2(new_n4981_), .ZN(new_n6595_));
  AOI21_X1   g06524(.A1(new_n6595_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6596_));
  XOR2_X1    g06525(.A1(new_n6134_), .A2(new_n6596_), .Z(new_n6597_));
  OAI21_X1   g06526(.A1(new_n6593_), .A2(new_n6594_), .B(new_n6597_), .ZN(new_n6598_));
  NAND2_X1   g06527(.A1(new_n6589_), .A2(new_n6598_), .ZN(new_n6599_));
  NOR2_X1    g06528(.A1(new_n6593_), .A2(new_n6594_), .ZN(new_n6600_));
  INV_X1     g06529(.I(new_n6597_), .ZN(new_n6601_));
  NAND2_X1   g06530(.A1(new_n6600_), .A2(new_n6601_), .ZN(new_n6602_));
  NAND2_X1   g06531(.A1(new_n6599_), .A2(new_n6602_), .ZN(new_n6603_));
  AOI22_X1   g06532(.A1(new_n6310_), .A2(new_n6312_), .B1(new_n6298_), .B2(new_n6299_), .ZN(new_n6604_));
  XNOR2_X1   g06533(.A1(new_n6305_), .A2(new_n6309_), .ZN(new_n6605_));
  NOR2_X1    g06534(.A1(new_n6605_), .A2(new_n6300_), .ZN(new_n6606_));
  NOR2_X1    g06535(.A1(new_n6606_), .A2(new_n6604_), .ZN(new_n6607_));
  INV_X1     g06536(.I(new_n6607_), .ZN(new_n6608_));
  NAND2_X1   g06537(.A1(new_n4143_), .A2(new_n4274_), .ZN(new_n6609_));
  NAND2_X1   g06538(.A1(new_n6609_), .A2(new_n5783_), .ZN(new_n6610_));
  OAI21_X1   g06539(.A1(new_n4135_), .A2(new_n1239_), .B(new_n6610_), .ZN(new_n6611_));
  AOI21_X1   g06540(.A1(new_n6611_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6612_));
  XOR2_X1    g06541(.A1(new_n5624_), .A2(new_n6612_), .Z(new_n6613_));
  OR2_X2     g06542(.A1(new_n6608_), .A2(new_n6613_), .Z(new_n6614_));
  NAND2_X1   g06543(.A1(new_n6608_), .A2(new_n6613_), .ZN(new_n6615_));
  NAND2_X1   g06544(.A1(new_n6614_), .A2(new_n6615_), .ZN(new_n6616_));
  NOR2_X1    g06545(.A1(new_n6616_), .A2(new_n6603_), .ZN(new_n6617_));
  NAND2_X1   g06546(.A1(new_n6617_), .A2(new_n6503_), .ZN(new_n6618_));
  NOR2_X1    g06547(.A1(new_n6617_), .A2(new_n6503_), .ZN(new_n6619_));
  INV_X1     g06548(.I(new_n6614_), .ZN(new_n6620_));
  NOR2_X1    g06549(.A1(new_n4135_), .A2(new_n4142_), .ZN(new_n6621_));
  OAI22_X1   g06550(.A1(new_n4285_), .A2(new_n1239_), .B1(new_n4981_), .B2(new_n6621_), .ZN(new_n6622_));
  AOI21_X1   g06551(.A1(new_n6622_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6623_));
  XOR2_X1    g06552(.A1(new_n5023_), .A2(new_n6623_), .Z(new_n6624_));
  NAND2_X1   g06553(.A1(new_n6620_), .A2(new_n6624_), .ZN(new_n6625_));
  OAI21_X1   g06554(.A1(new_n6619_), .A2(new_n6625_), .B(new_n6618_), .ZN(new_n6626_));
  NOR2_X1    g06555(.A1(new_n4285_), .A2(new_n4135_), .ZN(new_n6627_));
  OAI22_X1   g06556(.A1(new_n6627_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4296_), .ZN(new_n6628_));
  AOI21_X1   g06557(.A1(new_n6628_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6629_));
  XOR2_X1    g06558(.A1(new_n5753_), .A2(new_n6629_), .Z(new_n6630_));
  INV_X1     g06559(.I(new_n6630_), .ZN(new_n6631_));
  NAND2_X1   g06560(.A1(new_n6333_), .A2(new_n6324_), .ZN(new_n6632_));
  OAI21_X1   g06561(.A1(new_n6323_), .A2(new_n6325_), .B(new_n6632_), .ZN(new_n6633_));
  XOR2_X1    g06562(.A1(new_n6633_), .A2(new_n6313_), .Z(new_n6634_));
  NAND2_X1   g06563(.A1(new_n6634_), .A2(new_n6631_), .ZN(new_n6635_));
  NAND2_X1   g06564(.A1(new_n6626_), .A2(new_n6635_), .ZN(new_n6636_));
  XNOR2_X1   g06565(.A1(new_n6633_), .A2(new_n6313_), .ZN(new_n6637_));
  NAND2_X1   g06566(.A1(new_n6637_), .A2(new_n6630_), .ZN(new_n6638_));
  NAND2_X1   g06567(.A1(new_n6636_), .A2(new_n6638_), .ZN(new_n6639_));
  NAND2_X1   g06568(.A1(new_n6342_), .A2(new_n6241_), .ZN(new_n6640_));
  XNOR2_X1   g06569(.A1(new_n6640_), .A2(new_n6334_), .ZN(new_n6641_));
  XOR2_X1    g06570(.A1(new_n6641_), .A2(new_n6337_), .Z(new_n6642_));
  INV_X1     g06571(.I(new_n6642_), .ZN(new_n6643_));
  OAI22_X1   g06572(.A1(new_n4131_), .A2(new_n1239_), .B1(new_n4301_), .B2(new_n4981_), .ZN(new_n6644_));
  AOI21_X1   g06573(.A1(new_n6644_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6645_));
  XNOR2_X1   g06574(.A1(new_n5599_), .A2(new_n6645_), .ZN(new_n6646_));
  INV_X1     g06575(.I(new_n6646_), .ZN(new_n6647_));
  NOR2_X1    g06576(.A1(new_n6643_), .A2(new_n6647_), .ZN(new_n6648_));
  INV_X1     g06577(.I(new_n6648_), .ZN(new_n6649_));
  NAND2_X1   g06578(.A1(new_n6643_), .A2(new_n6647_), .ZN(new_n6650_));
  INV_X1     g06579(.I(new_n6650_), .ZN(new_n6651_));
  AOI21_X1   g06580(.A1(new_n6639_), .A2(new_n6649_), .B(new_n6651_), .ZN(new_n6652_));
  INV_X1     g06581(.I(new_n6355_), .ZN(new_n6653_));
  AOI21_X1   g06582(.A1(new_n6653_), .A2(new_n6354_), .B(new_n6345_), .ZN(new_n6654_));
  XNOR2_X1   g06583(.A1(new_n6349_), .A2(new_n6353_), .ZN(new_n6655_));
  NOR2_X1    g06584(.A1(new_n6655_), .A2(new_n6346_), .ZN(new_n6656_));
  NOR2_X1    g06585(.A1(new_n6656_), .A2(new_n6654_), .ZN(new_n6657_));
  INV_X1     g06586(.I(new_n6657_), .ZN(new_n6658_));
  NOR2_X1    g06587(.A1(new_n4131_), .A2(new_n4296_), .ZN(new_n6659_));
  OAI22_X1   g06588(.A1(new_n6659_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4309_), .ZN(new_n6660_));
  AOI21_X1   g06589(.A1(new_n6660_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6661_));
  XNOR2_X1   g06590(.A1(new_n5049_), .A2(new_n6661_), .ZN(new_n6662_));
  INV_X1     g06591(.I(new_n6662_), .ZN(new_n6663_));
  NOR2_X1    g06592(.A1(new_n6658_), .A2(new_n6663_), .ZN(new_n6664_));
  NOR2_X1    g06593(.A1(new_n6657_), .A2(new_n6662_), .ZN(new_n6665_));
  INV_X1     g06594(.I(new_n6665_), .ZN(new_n6666_));
  OAI21_X1   g06595(.A1(new_n6652_), .A2(new_n6664_), .B(new_n6666_), .ZN(new_n6667_));
  AND2_X2    g06596(.A1(new_n6367_), .A2(new_n6356_), .Z(new_n6668_));
  NOR2_X1    g06597(.A1(new_n6367_), .A2(new_n6356_), .ZN(new_n6669_));
  NOR2_X1    g06598(.A1(new_n6668_), .A2(new_n6669_), .ZN(new_n6670_));
  OAI22_X1   g06599(.A1(new_n4311_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4123_), .ZN(new_n6671_));
  AOI21_X1   g06600(.A1(new_n6671_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6672_));
  XOR2_X1    g06601(.A1(new_n5906_), .A2(new_n6672_), .Z(new_n6673_));
  NAND2_X1   g06602(.A1(new_n6670_), .A2(new_n6673_), .ZN(new_n6674_));
  NOR2_X1    g06603(.A1(new_n6670_), .A2(new_n6673_), .ZN(new_n6675_));
  INV_X1     g06604(.I(new_n6675_), .ZN(new_n6676_));
  NAND2_X1   g06605(.A1(new_n6676_), .A2(new_n6674_), .ZN(new_n6677_));
  NOR2_X1    g06606(.A1(new_n6677_), .A2(new_n6667_), .ZN(new_n6678_));
  INV_X1     g06607(.I(new_n6678_), .ZN(new_n6679_));
  INV_X1     g06608(.I(new_n6674_), .ZN(new_n6680_));
  NAND2_X1   g06609(.A1(new_n6679_), .A2(new_n6501_), .ZN(new_n6681_));
  NOR2_X1    g06610(.A1(new_n4123_), .A2(new_n4309_), .ZN(new_n6682_));
  OAI22_X1   g06611(.A1(new_n4112_), .A2(new_n1239_), .B1(new_n4981_), .B2(new_n6682_), .ZN(new_n6683_));
  AOI21_X1   g06612(.A1(new_n6683_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6684_));
  XOR2_X1    g06613(.A1(new_n5096_), .A2(new_n6684_), .Z(new_n6685_));
  INV_X1     g06614(.I(new_n6685_), .ZN(new_n6686_));
  NAND3_X1   g06615(.A1(new_n6681_), .A2(new_n6680_), .A3(new_n6686_), .ZN(new_n6687_));
  OAI21_X1   g06616(.A1(new_n6501_), .A2(new_n6679_), .B(new_n6687_), .ZN(new_n6688_));
  OAI21_X1   g06617(.A1(new_n6386_), .A2(new_n6388_), .B(new_n6376_), .ZN(new_n6689_));
  XOR2_X1    g06618(.A1(new_n6380_), .A2(new_n6384_), .Z(new_n6690_));
  OAI21_X1   g06619(.A1(new_n6376_), .A2(new_n6690_), .B(new_n6689_), .ZN(new_n6691_));
  NOR2_X1    g06620(.A1(new_n4112_), .A2(new_n4123_), .ZN(new_n6692_));
  OAI22_X1   g06621(.A1(new_n6692_), .A2(new_n4981_), .B1(new_n4315_), .B2(new_n1239_), .ZN(new_n6693_));
  AOI21_X1   g06622(.A1(new_n6693_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6694_));
  XNOR2_X1   g06623(.A1(new_n5121_), .A2(new_n6694_), .ZN(new_n6695_));
  INV_X1     g06624(.I(new_n6695_), .ZN(new_n6696_));
  NOR2_X1    g06625(.A1(new_n6691_), .A2(new_n6696_), .ZN(new_n6697_));
  INV_X1     g06626(.I(new_n6697_), .ZN(new_n6698_));
  NAND2_X1   g06627(.A1(new_n6691_), .A2(new_n6696_), .ZN(new_n6699_));
  NOR2_X1    g06628(.A1(new_n6400_), .A2(new_n6402_), .ZN(new_n6700_));
  NOR2_X1    g06629(.A1(new_n6700_), .A2(new_n6389_), .ZN(new_n6701_));
  XOR2_X1    g06630(.A1(new_n6393_), .A2(new_n6398_), .Z(new_n6702_));
  AOI21_X1   g06631(.A1(new_n6389_), .A2(new_n6702_), .B(new_n6701_), .ZN(new_n6703_));
  NOR2_X1    g06632(.A1(new_n4112_), .A2(new_n4315_), .ZN(new_n6704_));
  OAI22_X1   g06633(.A1(new_n6704_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4099_), .ZN(new_n6705_));
  AOI21_X1   g06634(.A1(new_n6705_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6706_));
  XNOR2_X1   g06635(.A1(new_n5080_), .A2(new_n6706_), .ZN(new_n6707_));
  NAND2_X1   g06636(.A1(new_n6703_), .A2(new_n6707_), .ZN(new_n6708_));
  INV_X1     g06637(.I(new_n6708_), .ZN(new_n6709_));
  NOR2_X1    g06638(.A1(new_n6703_), .A2(new_n6707_), .ZN(new_n6710_));
  NOR2_X1    g06639(.A1(new_n6709_), .A2(new_n6710_), .ZN(new_n6711_));
  NAND2_X1   g06640(.A1(new_n6698_), .A2(new_n6699_), .ZN(new_n6712_));
  NAND2_X1   g06641(.A1(new_n6688_), .A2(new_n6712_), .ZN(new_n6713_));
  NAND2_X1   g06642(.A1(new_n6713_), .A2(new_n6493_), .ZN(new_n6714_));
  OAI22_X1   g06643(.A1(new_n4090_), .A2(new_n1239_), .B1(new_n4320_), .B2(new_n4981_), .ZN(new_n6715_));
  AOI21_X1   g06644(.A1(new_n6715_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n6716_));
  XOR2_X1    g06645(.A1(new_n5196_), .A2(new_n6716_), .Z(new_n6717_));
  NOR2_X1    g06646(.A1(new_n6708_), .A2(new_n6717_), .ZN(new_n6718_));
  NAND2_X1   g06647(.A1(new_n6714_), .A2(new_n6718_), .ZN(new_n6719_));
  OAI21_X1   g06648(.A1(new_n6493_), .A2(new_n6713_), .B(new_n6719_), .ZN(new_n6720_));
  AOI22_X1   g06649(.A1(new_n4923_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4061_), .ZN(new_n6721_));
  OAI21_X1   g06650(.A1(new_n6721_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n6722_));
  XOR2_X1    g06651(.A1(new_n4935_), .A2(new_n6722_), .Z(new_n6723_));
  INV_X1     g06652(.I(new_n6723_), .ZN(new_n6724_));
  NOR2_X1    g06653(.A1(new_n6720_), .A2(new_n6724_), .ZN(new_n6725_));
  NAND2_X1   g06654(.A1(new_n6720_), .A2(new_n6724_), .ZN(new_n6726_));
  OAI21_X1   g06655(.A1(new_n6489_), .A2(new_n6725_), .B(new_n6726_), .ZN(new_n6727_));
  AOI22_X1   g06656(.A1(new_n5935_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4029_), .ZN(new_n6728_));
  OAI21_X1   g06657(.A1(new_n6728_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n6729_));
  XNOR2_X1   g06658(.A1(new_n4687_), .A2(new_n6729_), .ZN(new_n6730_));
  NAND2_X1   g06659(.A1(new_n6730_), .A2(new_n6727_), .ZN(new_n6731_));
  NOR2_X1    g06660(.A1(new_n6730_), .A2(new_n6727_), .ZN(new_n6732_));
  INV_X1     g06661(.I(new_n6431_), .ZN(new_n6733_));
  XOR2_X1    g06662(.A1(new_n6228_), .A2(new_n6427_), .Z(new_n6734_));
  XOR2_X1    g06663(.A1(new_n6734_), .A2(new_n6733_), .Z(new_n6735_));
  OAI21_X1   g06664(.A1(new_n6735_), .A2(new_n6732_), .B(new_n6731_), .ZN(new_n6736_));
  OAI22_X1   g06665(.A1(new_n4397_), .A2(new_n5966_), .B1(new_n1851_), .B2(new_n4374_), .ZN(new_n6737_));
  OAI21_X1   g06666(.A1(new_n4437_), .A2(new_n643_), .B(new_n6737_), .ZN(new_n6738_));
  AOI21_X1   g06667(.A1(new_n6738_), .A2(new_n279_), .B(new_n643_), .ZN(new_n6739_));
  XOR2_X1    g06668(.A1(new_n4541_), .A2(new_n6739_), .Z(new_n6740_));
  INV_X1     g06669(.I(new_n6740_), .ZN(new_n6741_));
  OAI21_X1   g06670(.A1(new_n6736_), .A2(new_n6741_), .B(new_n6484_), .ZN(new_n6742_));
  NAND2_X1   g06671(.A1(new_n6741_), .A2(new_n6736_), .ZN(new_n6743_));
  NAND2_X1   g06672(.A1(new_n6742_), .A2(new_n6743_), .ZN(new_n6744_));
  AOI22_X1   g06673(.A1(new_n4448_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4469_), .ZN(new_n6745_));
  OAI21_X1   g06674(.A1(new_n6745_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n6746_));
  XNOR2_X1   g06675(.A1(new_n4477_), .A2(new_n6746_), .ZN(new_n6747_));
  INV_X1     g06676(.I(new_n6747_), .ZN(new_n6748_));
  NAND2_X1   g06677(.A1(new_n6744_), .A2(new_n6748_), .ZN(new_n6749_));
  NOR2_X1    g06678(.A1(new_n6463_), .A2(new_n6449_), .ZN(new_n6750_));
  NOR2_X1    g06679(.A1(new_n6750_), .A2(new_n6460_), .ZN(new_n6751_));
  XOR2_X1    g06680(.A1(new_n6445_), .A2(new_n6448_), .Z(new_n6752_));
  AOI21_X1   g06681(.A1(new_n6460_), .A2(new_n6752_), .B(new_n6751_), .ZN(new_n6753_));
  OAI21_X1   g06682(.A1(new_n6744_), .A2(new_n6748_), .B(new_n6753_), .ZN(new_n6754_));
  NAND2_X1   g06683(.A1(new_n6754_), .A2(new_n6749_), .ZN(new_n6755_));
  INV_X1     g06684(.I(new_n5249_), .ZN(new_n6756_));
  NOR2_X1    g06685(.A1(new_n6756_), .A2(new_n2258_), .ZN(new_n6757_));
  INV_X1     g06686(.I(new_n6757_), .ZN(new_n6758_));
  AOI22_X1   g06687(.A1(new_n5418_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4563_), .ZN(new_n6759_));
  OAI21_X1   g06688(.A1(new_n6759_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n6760_));
  XNOR2_X1   g06689(.A1(new_n4594_), .A2(new_n6760_), .ZN(new_n6761_));
  INV_X1     g06690(.I(new_n6761_), .ZN(new_n6762_));
  NOR2_X1    g06691(.A1(new_n6755_), .A2(new_n6762_), .ZN(new_n6763_));
  INV_X1     g06692(.I(new_n6763_), .ZN(new_n6764_));
  NAND2_X1   g06693(.A1(new_n6481_), .A2(new_n6764_), .ZN(new_n6765_));
  NAND2_X1   g06694(.A1(new_n6755_), .A2(new_n6762_), .ZN(new_n6766_));
  NAND2_X1   g06695(.A1(new_n6765_), .A2(new_n6766_), .ZN(new_n6767_));
  NOR2_X1    g06696(.A1(new_n6767_), .A2(new_n2496_), .ZN(new_n6768_));
  INV_X1     g06697(.I(new_n5890_), .ZN(new_n6769_));
  OAI21_X1   g06698(.A1(new_n5950_), .A2(new_n5952_), .B(new_n6769_), .ZN(new_n6770_));
  XOR2_X1    g06699(.A1(new_n5948_), .A2(new_n5944_), .Z(new_n6771_));
  OAI21_X1   g06700(.A1(new_n6769_), .A2(new_n6771_), .B(new_n6770_), .ZN(new_n6772_));
  NOR3_X1    g06701(.A1(new_n6042_), .A2(new_n6469_), .A3(new_n6470_), .ZN(new_n6773_));
  INV_X1     g06702(.I(new_n6773_), .ZN(new_n6774_));
  NOR2_X1    g06703(.A1(new_n6471_), .A2(new_n6041_), .ZN(new_n6775_));
  AOI21_X1   g06704(.A1(new_n6774_), .A2(new_n6468_), .B(new_n6775_), .ZN(new_n6776_));
  OAI22_X1   g06705(.A1(new_n1851_), .A2(new_n4468_), .B1(new_n4501_), .B2(new_n5966_), .ZN(new_n6777_));
  OAI21_X1   g06706(.A1(new_n4516_), .A2(new_n643_), .B(new_n6777_), .ZN(new_n6778_));
  AOI21_X1   g06707(.A1(new_n6778_), .A2(new_n279_), .B(new_n643_), .ZN(new_n6779_));
  XOR2_X1    g06708(.A1(new_n4524_), .A2(new_n6779_), .Z(new_n6780_));
  AND2_X2    g06709(.A1(new_n6780_), .A2(new_n6776_), .Z(new_n6781_));
  NOR2_X1    g06710(.A1(new_n6780_), .A2(new_n6776_), .ZN(new_n6782_));
  NOR2_X1    g06711(.A1(new_n6781_), .A2(new_n6782_), .ZN(new_n6783_));
  XNOR2_X1   g06712(.A1(new_n6780_), .A2(new_n6776_), .ZN(new_n6784_));
  MUX2_X1    g06713(.I0(new_n6784_), .I1(new_n6783_), .S(new_n6772_), .Z(new_n6785_));
  INV_X1     g06714(.I(new_n6478_), .ZN(new_n6786_));
  NOR2_X1    g06715(.A1(new_n6786_), .A2(new_n6465_), .ZN(new_n6787_));
  XOR2_X1    g06716(.A1(new_n6472_), .A2(new_n6042_), .Z(new_n6788_));
  AOI21_X1   g06717(.A1(new_n6786_), .A2(new_n6465_), .B(new_n6788_), .ZN(new_n6789_));
  NOR2_X1    g06718(.A1(new_n6789_), .A2(new_n6787_), .ZN(new_n6790_));
  XOR2_X1    g06719(.A1(new_n6785_), .A2(new_n6790_), .Z(new_n6791_));
  NAND2_X1   g06720(.A1(new_n4563_), .A2(new_n5249_), .ZN(new_n6792_));
  NAND2_X1   g06721(.A1(new_n4564_), .A2(new_n5247_), .ZN(new_n6793_));
  AOI22_X1   g06722(.A1(new_n6793_), .A2(new_n6792_), .B1(new_n805_), .B2(new_n4564_), .ZN(new_n6794_));
  OAI21_X1   g06723(.A1(new_n6794_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n6795_));
  XOR2_X1    g06724(.A1(new_n4609_), .A2(new_n6795_), .Z(new_n6796_));
  XOR2_X1    g06725(.A1(new_n6791_), .A2(new_n6796_), .Z(new_n6797_));
  NOR2_X1    g06726(.A1(new_n6768_), .A2(new_n6797_), .ZN(new_n6798_));
  AOI21_X1   g06727(.A1(new_n2496_), .A2(new_n6767_), .B(new_n6798_), .ZN(new_n6799_));
  AOI21_X1   g06728(.A1(new_n6790_), .A2(new_n6796_), .B(new_n6785_), .ZN(new_n6800_));
  NOR2_X1    g06729(.A1(new_n6790_), .A2(new_n6796_), .ZN(new_n6801_));
  NOR2_X1    g06730(.A1(new_n6800_), .A2(new_n6801_), .ZN(new_n6802_));
  AOI22_X1   g06731(.A1(new_n5553_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4564_), .ZN(new_n6803_));
  OAI21_X1   g06732(.A1(new_n6803_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n6804_));
  XOR2_X1    g06733(.A1(new_n4569_), .A2(new_n6804_), .Z(new_n6805_));
  INV_X1     g06734(.I(new_n6781_), .ZN(new_n6806_));
  AOI21_X1   g06735(.A1(new_n6806_), .A2(new_n6772_), .B(new_n6782_), .ZN(new_n6807_));
  XNOR2_X1   g06736(.A1(new_n5956_), .A2(new_n5858_), .ZN(new_n6808_));
  NOR2_X1    g06737(.A1(new_n6808_), .A2(new_n5962_), .ZN(new_n6809_));
  XOR2_X1    g06738(.A1(new_n5956_), .A2(new_n5858_), .Z(new_n6810_));
  INV_X1     g06739(.I(new_n6810_), .ZN(new_n6811_));
  AOI21_X1   g06740(.A1(new_n5962_), .A2(new_n6811_), .B(new_n6809_), .ZN(new_n6812_));
  XNOR2_X1   g06741(.A1(new_n6812_), .A2(new_n5953_), .ZN(new_n6813_));
  XNOR2_X1   g06742(.A1(new_n6813_), .A2(new_n6807_), .ZN(new_n6814_));
  XNOR2_X1   g06743(.A1(new_n6814_), .A2(new_n6805_), .ZN(new_n6815_));
  NAND2_X1   g06744(.A1(new_n5249_), .A2(new_n805_), .ZN(new_n6816_));
  OAI21_X1   g06745(.A1(new_n5247_), .A2(new_n6816_), .B(new_n4564_), .ZN(new_n6817_));
  OAI21_X1   g06746(.A1(new_n6817_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n6818_));
  XOR2_X1    g06747(.A1(new_n5001_), .A2(new_n6818_), .Z(new_n6819_));
  XOR2_X1    g06748(.A1(new_n6815_), .A2(new_n6819_), .Z(new_n6820_));
  NOR2_X1    g06749(.A1(new_n6820_), .A2(new_n6802_), .ZN(new_n6821_));
  INV_X1     g06750(.I(new_n6819_), .ZN(new_n6822_));
  NOR2_X1    g06751(.A1(new_n6815_), .A2(new_n6822_), .ZN(new_n6823_));
  INV_X1     g06752(.I(new_n6823_), .ZN(new_n6824_));
  NAND2_X1   g06753(.A1(new_n6815_), .A2(new_n6822_), .ZN(new_n6825_));
  NAND2_X1   g06754(.A1(new_n6824_), .A2(new_n6825_), .ZN(new_n6826_));
  AOI21_X1   g06755(.A1(new_n6802_), .A2(new_n6826_), .B(new_n6821_), .ZN(new_n6827_));
  NOR2_X1    g06756(.A1(new_n6827_), .A2(new_n6799_), .ZN(new_n6828_));
  XOR2_X1    g06757(.A1(new_n6730_), .A2(new_n6734_), .Z(new_n6829_));
  XOR2_X1    g06758(.A1(new_n6829_), .A2(new_n6727_), .Z(new_n6830_));
  XOR2_X1    g06759(.A1(new_n6830_), .A2(new_n6733_), .Z(new_n6831_));
  INV_X1     g06760(.I(new_n6831_), .ZN(new_n6832_));
  OAI21_X1   g06761(.A1(new_n6499_), .A2(new_n6500_), .B(new_n6686_), .ZN(new_n6833_));
  NOR2_X1    g06762(.A1(new_n6678_), .A2(new_n6833_), .ZN(new_n6834_));
  AND2_X2    g06763(.A1(new_n6678_), .A2(new_n6833_), .Z(new_n6835_));
  NOR2_X1    g06764(.A1(new_n6835_), .A2(new_n6834_), .ZN(new_n6836_));
  NOR2_X1    g06765(.A1(new_n6836_), .A2(new_n6680_), .ZN(new_n6837_));
  NOR3_X1    g06766(.A1(new_n6835_), .A2(new_n6674_), .A3(new_n6834_), .ZN(new_n6838_));
  NOR2_X1    g06767(.A1(new_n6837_), .A2(new_n6838_), .ZN(new_n6839_));
  XOR2_X1    g06768(.A1(new_n6642_), .A2(new_n6646_), .Z(new_n6840_));
  NAND2_X1   g06769(.A1(new_n6639_), .A2(new_n6840_), .ZN(new_n6841_));
  INV_X1     g06770(.I(new_n6639_), .ZN(new_n6842_));
  OAI21_X1   g06771(.A1(new_n6651_), .A2(new_n6648_), .B(new_n6842_), .ZN(new_n6843_));
  NAND2_X1   g06772(.A1(new_n6843_), .A2(new_n6841_), .ZN(new_n6844_));
  INV_X1     g06773(.I(new_n6844_), .ZN(new_n6845_));
  INV_X1     g06774(.I(new_n6589_), .ZN(new_n6846_));
  XOR2_X1    g06775(.A1(new_n6600_), .A2(new_n6597_), .Z(new_n6847_));
  NOR2_X1    g06776(.A1(new_n6847_), .A2(new_n6846_), .ZN(new_n6848_));
  AOI21_X1   g06777(.A1(new_n6598_), .A2(new_n6602_), .B(new_n6589_), .ZN(new_n6849_));
  NOR2_X1    g06778(.A1(new_n6848_), .A2(new_n6849_), .ZN(new_n6850_));
  NAND2_X1   g06779(.A1(new_n6609_), .A2(new_n5337_), .ZN(new_n6851_));
  OAI21_X1   g06780(.A1(new_n4135_), .A2(new_n5398_), .B(new_n6851_), .ZN(new_n6852_));
  AOI21_X1   g06781(.A1(new_n6852_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n6853_));
  XNOR2_X1   g06782(.A1(new_n5624_), .A2(new_n6853_), .ZN(new_n6854_));
  NAND2_X1   g06783(.A1(new_n6561_), .A2(new_n6562_), .ZN(new_n6855_));
  XNOR2_X1   g06784(.A1(new_n6570_), .A2(new_n6565_), .ZN(new_n6856_));
  NAND2_X1   g06785(.A1(new_n6856_), .A2(new_n6855_), .ZN(new_n6857_));
  NOR2_X1    g06786(.A1(new_n6574_), .A2(new_n6571_), .ZN(new_n6858_));
  OR2_X2     g06787(.A1(new_n6858_), .A2(new_n6855_), .Z(new_n6859_));
  NAND2_X1   g06788(.A1(new_n6859_), .A2(new_n6857_), .ZN(new_n6860_));
  INV_X1     g06789(.I(new_n6860_), .ZN(new_n6861_));
  INV_X1     g06790(.I(new_n6587_), .ZN(new_n6862_));
  AOI21_X1   g06791(.A1(new_n6862_), .A2(new_n6588_), .B(new_n6575_), .ZN(new_n6863_));
  XOR2_X1    g06792(.A1(new_n6581_), .A2(new_n6585_), .Z(new_n6864_));
  NOR3_X1    g06793(.A1(new_n6864_), .A2(new_n6572_), .A3(new_n6574_), .ZN(new_n6865_));
  NOR2_X1    g06794(.A1(new_n6865_), .A2(new_n6863_), .ZN(new_n6866_));
  OAI22_X1   g06795(.A1(new_n4285_), .A2(new_n5398_), .B1(new_n5336_), .B2(new_n6621_), .ZN(new_n6867_));
  AOI21_X1   g06796(.A1(new_n6867_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n6868_));
  XNOR2_X1   g06797(.A1(new_n5023_), .A2(new_n6868_), .ZN(new_n6869_));
  AND2_X2    g06798(.A1(new_n6866_), .A2(new_n6869_), .Z(new_n6870_));
  NOR2_X1    g06799(.A1(new_n6866_), .A2(new_n6869_), .ZN(new_n6871_));
  NOR2_X1    g06800(.A1(new_n6870_), .A2(new_n6871_), .ZN(new_n6872_));
  OAI21_X1   g06801(.A1(new_n6872_), .A2(new_n6861_), .B(new_n6854_), .ZN(new_n6873_));
  INV_X1     g06802(.I(new_n6520_), .ZN(new_n6874_));
  OAI22_X1   g06803(.A1(new_n6504_), .A2(new_n5336_), .B1(new_n5398_), .B2(new_n4249_), .ZN(new_n6875_));
  AOI21_X1   g06804(.A1(new_n6875_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n6876_));
  XOR2_X1    g06805(.A1(new_n5648_), .A2(new_n6876_), .Z(new_n6877_));
  NAND2_X1   g06806(.A1(new_n6877_), .A2(new_n6874_), .ZN(new_n6878_));
  NAND2_X1   g06807(.A1(new_n5627_), .A2(new_n5398_), .ZN(new_n6879_));
  AOI21_X1   g06808(.A1(new_n4717_), .A2(new_n6061_), .B(new_n4260_), .ZN(new_n6880_));
  OAI22_X1   g06809(.A1(new_n4244_), .A2(new_n5335_), .B1(new_n4230_), .B2(new_n4719_), .ZN(new_n6881_));
  OAI21_X1   g06810(.A1(new_n5398_), .A2(new_n4234_), .B(new_n6881_), .ZN(new_n6882_));
  AOI21_X1   g06811(.A1(new_n6879_), .A2(new_n6880_), .B(new_n6882_), .ZN(new_n6883_));
  XOR2_X1    g06812(.A1(new_n6883_), .A2(new_n90_), .Z(new_n6884_));
  NOR2_X1    g06813(.A1(new_n4244_), .A2(new_n4719_), .ZN(new_n6885_));
  OAI21_X1   g06814(.A1(new_n4230_), .A2(new_n5398_), .B(new_n90_), .ZN(new_n6886_));
  OAI21_X1   g06815(.A1(new_n6885_), .A2(new_n6886_), .B(new_n4717_), .ZN(new_n6887_));
  XNOR2_X1   g06816(.A1(new_n6887_), .A2(new_n5637_), .ZN(new_n6888_));
  NOR2_X1    g06817(.A1(new_n4251_), .A2(new_n1467_), .ZN(new_n6889_));
  NOR2_X1    g06818(.A1(new_n6889_), .A2(new_n90_), .ZN(new_n6890_));
  NAND2_X1   g06819(.A1(new_n6888_), .A2(new_n6890_), .ZN(new_n6891_));
  NOR2_X1    g06820(.A1(new_n6884_), .A2(new_n6891_), .ZN(new_n6892_));
  NOR2_X1    g06821(.A1(new_n6877_), .A2(new_n6874_), .ZN(new_n6893_));
  OAI21_X1   g06822(.A1(new_n6892_), .A2(new_n6893_), .B(new_n6878_), .ZN(new_n6894_));
  XOR2_X1    g06823(.A1(new_n6519_), .A2(new_n6521_), .Z(new_n6895_));
  OAI22_X1   g06824(.A1(new_n4203_), .A2(new_n5398_), .B1(new_n5336_), .B2(new_n6529_), .ZN(new_n6896_));
  AOI21_X1   g06825(.A1(new_n6896_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n6897_));
  XOR2_X1    g06826(.A1(new_n6082_), .A2(new_n6897_), .Z(new_n6898_));
  NAND2_X1   g06827(.A1(new_n6898_), .A2(new_n6895_), .ZN(new_n6899_));
  NOR2_X1    g06828(.A1(new_n6898_), .A2(new_n6895_), .ZN(new_n6900_));
  AOI21_X1   g06829(.A1(new_n6894_), .A2(new_n6899_), .B(new_n6900_), .ZN(new_n6901_));
  XNOR2_X1   g06830(.A1(new_n6515_), .A2(new_n6522_), .ZN(new_n6902_));
  AOI22_X1   g06831(.A1(new_n4258_), .A2(new_n4717_), .B1(new_n5337_), .B2(new_n6541_), .ZN(new_n6903_));
  OAI21_X1   g06832(.A1(new_n6903_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n6904_));
  XOR2_X1    g06833(.A1(new_n6540_), .A2(new_n6904_), .Z(new_n6905_));
  NOR2_X1    g06834(.A1(new_n6905_), .A2(new_n6902_), .ZN(new_n6906_));
  NAND2_X1   g06835(.A1(new_n6905_), .A2(new_n6902_), .ZN(new_n6907_));
  OAI21_X1   g06836(.A1(new_n6901_), .A2(new_n6906_), .B(new_n6907_), .ZN(new_n6908_));
  XOR2_X1    g06837(.A1(new_n6508_), .A2(new_n6261_), .Z(new_n6909_));
  NAND2_X1   g06838(.A1(new_n6909_), .A2(new_n6523_), .ZN(new_n6910_));
  INV_X1     g06839(.I(new_n6525_), .ZN(new_n6911_));
  OAI21_X1   g06840(.A1(new_n6911_), .A2(new_n6509_), .B(new_n6524_), .ZN(new_n6912_));
  OAI22_X1   g06841(.A1(new_n5684_), .A2(new_n5398_), .B1(new_n6556_), .B2(new_n5336_), .ZN(new_n6913_));
  AOI21_X1   g06842(.A1(new_n6913_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n6914_));
  XOR2_X1    g06843(.A1(new_n6102_), .A2(new_n6914_), .Z(new_n6915_));
  NAND3_X1   g06844(.A1(new_n6915_), .A2(new_n6910_), .A3(new_n6912_), .ZN(new_n6916_));
  NAND2_X1   g06845(.A1(new_n6916_), .A2(new_n6908_), .ZN(new_n6917_));
  NAND2_X1   g06846(.A1(new_n6910_), .A2(new_n6912_), .ZN(new_n6918_));
  INV_X1     g06847(.I(new_n6915_), .ZN(new_n6919_));
  NAND2_X1   g06848(.A1(new_n6919_), .A2(new_n6918_), .ZN(new_n6920_));
  XOR2_X1    g06849(.A1(new_n6532_), .A2(new_n6527_), .Z(new_n6921_));
  OAI21_X1   g06850(.A1(new_n6536_), .A2(new_n6533_), .B(new_n6526_), .ZN(new_n6922_));
  OAI21_X1   g06851(.A1(new_n6921_), .A2(new_n6526_), .B(new_n6922_), .ZN(new_n6923_));
  INV_X1     g06852(.I(new_n6923_), .ZN(new_n6924_));
  OAI22_X1   g06853(.A1(new_n4150_), .A2(new_n5398_), .B1(new_n6567_), .B2(new_n5336_), .ZN(new_n6925_));
  AOI21_X1   g06854(.A1(new_n6925_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n6926_));
  XNOR2_X1   g06855(.A1(new_n5707_), .A2(new_n6926_), .ZN(new_n6927_));
  NOR2_X1    g06856(.A1(new_n6924_), .A2(new_n6927_), .ZN(new_n6928_));
  AOI21_X1   g06857(.A1(new_n6917_), .A2(new_n6920_), .B(new_n6928_), .ZN(new_n6929_));
  INV_X1     g06858(.I(new_n6927_), .ZN(new_n6930_));
  NOR2_X1    g06859(.A1(new_n6930_), .A2(new_n6923_), .ZN(new_n6931_));
  NOR2_X1    g06860(.A1(new_n6929_), .A2(new_n6931_), .ZN(new_n6932_));
  XOR2_X1    g06861(.A1(new_n6545_), .A2(new_n6538_), .Z(new_n6933_));
  NOR2_X1    g06862(.A1(new_n6933_), .A2(new_n6537_), .ZN(new_n6934_));
  NAND2_X1   g06863(.A1(new_n6546_), .A2(new_n6549_), .ZN(new_n6935_));
  AND2_X2    g06864(.A1(new_n6935_), .A2(new_n6537_), .Z(new_n6936_));
  AOI22_X1   g06865(.A1(new_n6582_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4274_), .ZN(new_n6937_));
  OAI21_X1   g06866(.A1(new_n6937_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n6938_));
  XOR2_X1    g06867(.A1(new_n5722_), .A2(new_n6938_), .Z(new_n6939_));
  OAI21_X1   g06868(.A1(new_n6934_), .A2(new_n6936_), .B(new_n6939_), .ZN(new_n6940_));
  INV_X1     g06869(.I(new_n6940_), .ZN(new_n6941_));
  NOR2_X1    g06870(.A1(new_n6936_), .A2(new_n6934_), .ZN(new_n6942_));
  INV_X1     g06871(.I(new_n6939_), .ZN(new_n6943_));
  NAND2_X1   g06872(.A1(new_n6943_), .A2(new_n6942_), .ZN(new_n6944_));
  OAI21_X1   g06873(.A1(new_n6941_), .A2(new_n6932_), .B(new_n6944_), .ZN(new_n6945_));
  INV_X1     g06874(.I(new_n6550_), .ZN(new_n6946_));
  XNOR2_X1   g06875(.A1(new_n6559_), .A2(new_n6555_), .ZN(new_n6947_));
  NOR2_X1    g06876(.A1(new_n6947_), .A2(new_n6946_), .ZN(new_n6948_));
  AOI21_X1   g06877(.A1(new_n6562_), .A2(new_n6560_), .B(new_n6550_), .ZN(new_n6949_));
  OAI22_X1   g06878(.A1(new_n4142_), .A2(new_n5398_), .B1(new_n4277_), .B2(new_n5336_), .ZN(new_n6950_));
  AOI21_X1   g06879(.A1(new_n6950_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n6951_));
  XOR2_X1    g06880(.A1(new_n6134_), .A2(new_n6951_), .Z(new_n6952_));
  OAI21_X1   g06881(.A1(new_n6948_), .A2(new_n6949_), .B(new_n6952_), .ZN(new_n6953_));
  NAND2_X1   g06882(.A1(new_n6945_), .A2(new_n6953_), .ZN(new_n6954_));
  NOR2_X1    g06883(.A1(new_n6948_), .A2(new_n6949_), .ZN(new_n6955_));
  INV_X1     g06884(.I(new_n6952_), .ZN(new_n6956_));
  NAND2_X1   g06885(.A1(new_n6955_), .A2(new_n6956_), .ZN(new_n6957_));
  AOI22_X1   g06886(.A1(new_n6872_), .A2(new_n6861_), .B1(new_n6954_), .B2(new_n6957_), .ZN(new_n6958_));
  NAND2_X1   g06887(.A1(new_n6958_), .A2(new_n6873_), .ZN(new_n6959_));
  NOR2_X1    g06888(.A1(new_n6959_), .A2(new_n6850_), .ZN(new_n6960_));
  INV_X1     g06889(.I(new_n6627_), .ZN(new_n6961_));
  AOI22_X1   g06890(.A1(new_n6961_), .A2(new_n5337_), .B1(new_n4297_), .B2(new_n4717_), .ZN(new_n6962_));
  OAI21_X1   g06891(.A1(new_n6962_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n6963_));
  XOR2_X1    g06892(.A1(new_n5753_), .A2(new_n6963_), .Z(new_n6964_));
  INV_X1     g06893(.I(new_n6964_), .ZN(new_n6965_));
  NAND2_X1   g06894(.A1(new_n6965_), .A2(new_n6870_), .ZN(new_n6966_));
  AOI21_X1   g06895(.A1(new_n6959_), .A2(new_n6850_), .B(new_n6966_), .ZN(new_n6967_));
  NOR2_X1    g06896(.A1(new_n6967_), .A2(new_n6960_), .ZN(new_n6968_));
  OAI22_X1   g06897(.A1(new_n4131_), .A2(new_n5398_), .B1(new_n4301_), .B2(new_n5336_), .ZN(new_n6969_));
  AOI21_X1   g06898(.A1(new_n6969_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n6970_));
  XNOR2_X1   g06899(.A1(new_n5599_), .A2(new_n6970_), .ZN(new_n6971_));
  NOR2_X1    g06900(.A1(new_n6968_), .A2(new_n6971_), .ZN(new_n6972_));
  INV_X1     g06901(.I(new_n6603_), .ZN(new_n6973_));
  XOR2_X1    g06902(.A1(new_n6616_), .A2(new_n6973_), .Z(new_n6974_));
  AOI21_X1   g06903(.A1(new_n6968_), .A2(new_n6971_), .B(new_n6974_), .ZN(new_n6975_));
  NOR2_X1    g06904(.A1(new_n6975_), .A2(new_n6972_), .ZN(new_n6976_));
  NAND2_X1   g06905(.A1(new_n6503_), .A2(new_n6624_), .ZN(new_n6977_));
  XOR2_X1    g06906(.A1(new_n6617_), .A2(new_n6977_), .Z(new_n6978_));
  XOR2_X1    g06907(.A1(new_n6978_), .A2(new_n6620_), .Z(new_n6979_));
  INV_X1     g06908(.I(new_n6659_), .ZN(new_n6980_));
  AOI22_X1   g06909(.A1(new_n6980_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n5041_), .ZN(new_n6981_));
  OAI21_X1   g06910(.A1(new_n6981_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n6982_));
  XOR2_X1    g06911(.A1(new_n5049_), .A2(new_n6982_), .Z(new_n6983_));
  INV_X1     g06912(.I(new_n6983_), .ZN(new_n6984_));
  NOR2_X1    g06913(.A1(new_n6979_), .A2(new_n6984_), .ZN(new_n6985_));
  NOR2_X1    g06914(.A1(new_n6976_), .A2(new_n6985_), .ZN(new_n6986_));
  NAND2_X1   g06915(.A1(new_n6979_), .A2(new_n6984_), .ZN(new_n6987_));
  INV_X1     g06916(.I(new_n6987_), .ZN(new_n6988_));
  NOR2_X1    g06917(.A1(new_n6986_), .A2(new_n6988_), .ZN(new_n6989_));
  XOR2_X1    g06918(.A1(new_n6634_), .A2(new_n6631_), .Z(new_n6990_));
  NAND2_X1   g06919(.A1(new_n6638_), .A2(new_n6635_), .ZN(new_n6991_));
  MUX2_X1    g06920(.I0(new_n6991_), .I1(new_n6990_), .S(new_n6626_), .Z(new_n6992_));
  INV_X1     g06921(.I(new_n4311_), .ZN(new_n6993_));
  AOI22_X1   g06922(.A1(new_n6993_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4124_), .ZN(new_n6994_));
  OAI21_X1   g06923(.A1(new_n6994_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n6995_));
  XOR2_X1    g06924(.A1(new_n5067_), .A2(new_n6995_), .Z(new_n6996_));
  NOR2_X1    g06925(.A1(new_n6992_), .A2(new_n6996_), .ZN(new_n6997_));
  NAND2_X1   g06926(.A1(new_n6992_), .A2(new_n6996_), .ZN(new_n6998_));
  INV_X1     g06927(.I(new_n6998_), .ZN(new_n6999_));
  NOR2_X1    g06928(.A1(new_n6999_), .A2(new_n6997_), .ZN(new_n7000_));
  NAND2_X1   g06929(.A1(new_n6989_), .A2(new_n7000_), .ZN(new_n7001_));
  NOR2_X1    g06930(.A1(new_n7001_), .A2(new_n6845_), .ZN(new_n7002_));
  OAI22_X1   g06931(.A1(new_n4112_), .A2(new_n5398_), .B1(new_n5336_), .B2(new_n6682_), .ZN(new_n7003_));
  AOI21_X1   g06932(.A1(new_n7003_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n7004_));
  XNOR2_X1   g06933(.A1(new_n5096_), .A2(new_n7004_), .ZN(new_n7005_));
  NAND2_X1   g06934(.A1(new_n6999_), .A2(new_n7005_), .ZN(new_n7006_));
  AOI21_X1   g06935(.A1(new_n7001_), .A2(new_n6845_), .B(new_n7006_), .ZN(new_n7007_));
  NOR2_X1    g06936(.A1(new_n7007_), .A2(new_n7002_), .ZN(new_n7008_));
  INV_X1     g06937(.I(new_n7008_), .ZN(new_n7009_));
  XOR2_X1    g06938(.A1(new_n6657_), .A2(new_n6663_), .Z(new_n7010_));
  NOR2_X1    g06939(.A1(new_n7010_), .A2(new_n6652_), .ZN(new_n7011_));
  INV_X1     g06940(.I(new_n6652_), .ZN(new_n7012_));
  NOR2_X1    g06941(.A1(new_n6664_), .A2(new_n6665_), .ZN(new_n7013_));
  NOR2_X1    g06942(.A1(new_n7013_), .A2(new_n7012_), .ZN(new_n7014_));
  INV_X1     g06943(.I(new_n6692_), .ZN(new_n7015_));
  AOI22_X1   g06944(.A1(new_n7015_), .A2(new_n5337_), .B1(new_n4105_), .B2(new_n4717_), .ZN(new_n7016_));
  OAI21_X1   g06945(.A1(new_n7016_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n7017_));
  XOR2_X1    g06946(.A1(new_n5121_), .A2(new_n7017_), .Z(new_n7018_));
  OR3_X2     g06947(.A1(new_n7011_), .A2(new_n7014_), .A3(new_n7018_), .Z(new_n7019_));
  OAI21_X1   g06948(.A1(new_n7014_), .A2(new_n7011_), .B(new_n7018_), .ZN(new_n7020_));
  INV_X1     g06949(.I(new_n6704_), .ZN(new_n7021_));
  AOI22_X1   g06950(.A1(new_n7021_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4100_), .ZN(new_n7022_));
  OAI21_X1   g06951(.A1(new_n7022_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n7023_));
  NOR2_X1    g06952(.A1(new_n5080_), .A2(new_n7023_), .ZN(new_n7024_));
  AND2_X2    g06953(.A1(new_n5080_), .A2(new_n7023_), .Z(new_n7025_));
  NOR2_X1    g06954(.A1(new_n7025_), .A2(new_n7024_), .ZN(new_n7026_));
  INV_X1     g06955(.I(new_n7026_), .ZN(new_n7027_));
  NOR2_X1    g06956(.A1(new_n6677_), .A2(new_n7027_), .ZN(new_n7028_));
  INV_X1     g06957(.I(new_n6677_), .ZN(new_n7029_));
  NOR2_X1    g06958(.A1(new_n7029_), .A2(new_n7026_), .ZN(new_n7030_));
  OAI21_X1   g06959(.A1(new_n7030_), .A2(new_n7028_), .B(new_n6667_), .ZN(new_n7031_));
  INV_X1     g06960(.I(new_n6667_), .ZN(new_n7033_));
  NOR2_X1    g06961(.A1(new_n7029_), .A2(new_n7027_), .ZN(new_n7034_));
  NOR2_X1    g06962(.A1(new_n6677_), .A2(new_n7026_), .ZN(new_n7035_));
  OAI21_X1   g06963(.A1(new_n7034_), .A2(new_n7035_), .B(new_n7033_), .ZN(new_n7036_));
  NAND2_X1   g06964(.A1(new_n7019_), .A2(new_n7020_), .ZN(new_n7038_));
  NAND2_X1   g06965(.A1(new_n7009_), .A2(new_n7038_), .ZN(new_n7039_));
  NOR2_X1    g06966(.A1(new_n7039_), .A2(new_n6839_), .ZN(new_n7040_));
  XOR2_X1    g06967(.A1(new_n6677_), .A2(new_n6667_), .Z(new_n7041_));
  NAND2_X1   g06968(.A1(new_n7041_), .A2(new_n7026_), .ZN(new_n7042_));
  INV_X1     g06969(.I(new_n7042_), .ZN(new_n7043_));
  OAI22_X1   g06970(.A1(new_n4090_), .A2(new_n5398_), .B1(new_n4320_), .B2(new_n5336_), .ZN(new_n7044_));
  AOI21_X1   g06971(.A1(new_n7044_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n7045_));
  XOR2_X1    g06972(.A1(new_n5196_), .A2(new_n7045_), .Z(new_n7046_));
  INV_X1     g06973(.I(new_n7046_), .ZN(new_n7047_));
  NAND2_X1   g06974(.A1(new_n7043_), .A2(new_n7047_), .ZN(new_n7048_));
  AOI21_X1   g06975(.A1(new_n7039_), .A2(new_n6839_), .B(new_n7048_), .ZN(new_n7049_));
  NOR2_X1    g06976(.A1(new_n7049_), .A2(new_n7040_), .ZN(new_n7050_));
  AOI22_X1   g06977(.A1(new_n6419_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4328_), .ZN(new_n7051_));
  OAI21_X1   g06978(.A1(new_n7051_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n7052_));
  XNOR2_X1   g06979(.A1(new_n5139_), .A2(new_n7052_), .ZN(new_n7053_));
  NOR2_X1    g06980(.A1(new_n7050_), .A2(new_n7053_), .ZN(new_n7054_));
  NAND2_X1   g06981(.A1(new_n6698_), .A2(new_n6699_), .ZN(new_n7055_));
  XNOR2_X1   g06982(.A1(new_n6688_), .A2(new_n7055_), .ZN(new_n7056_));
  NAND2_X1   g06983(.A1(new_n7050_), .A2(new_n7053_), .ZN(new_n7057_));
  AOI21_X1   g06984(.A1(new_n7056_), .A2(new_n7057_), .B(new_n7054_), .ZN(new_n7058_));
  INV_X1     g06985(.I(new_n7058_), .ZN(new_n7059_));
  INV_X1     g06986(.I(new_n6688_), .ZN(new_n7060_));
  NAND2_X1   g06987(.A1(new_n6711_), .A2(new_n6698_), .ZN(new_n7061_));
  NAND3_X1   g06988(.A1(new_n7061_), .A2(new_n7060_), .A3(new_n7055_), .ZN(new_n7062_));
  INV_X1     g06989(.I(new_n7062_), .ZN(new_n7063_));
  AOI21_X1   g06990(.A1(new_n7061_), .A2(new_n7055_), .B(new_n7060_), .ZN(new_n7064_));
  NOR2_X1    g06991(.A1(new_n7063_), .A2(new_n7064_), .ZN(new_n7065_));
  AOI22_X1   g06992(.A1(new_n4333_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4082_), .ZN(new_n7066_));
  OAI21_X1   g06993(.A1(new_n7066_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n7067_));
  XNOR2_X1   g06994(.A1(new_n5162_), .A2(new_n7067_), .ZN(new_n7068_));
  INV_X1     g06995(.I(new_n7068_), .ZN(new_n7069_));
  NOR2_X1    g06996(.A1(new_n7065_), .A2(new_n7069_), .ZN(new_n7070_));
  INV_X1     g06997(.I(new_n7070_), .ZN(new_n7071_));
  NAND2_X1   g06998(.A1(new_n7059_), .A2(new_n7071_), .ZN(new_n7072_));
  NAND2_X1   g06999(.A1(new_n7065_), .A2(new_n7069_), .ZN(new_n7073_));
  NAND2_X1   g07000(.A1(new_n7072_), .A2(new_n7073_), .ZN(new_n7074_));
  NOR2_X1    g07001(.A1(new_n6493_), .A2(new_n6717_), .ZN(new_n7075_));
  XOR2_X1    g07002(.A1(new_n7075_), .A2(new_n6713_), .Z(new_n7076_));
  XOR2_X1    g07003(.A1(new_n7076_), .A2(new_n6709_), .Z(new_n7077_));
  OAI22_X1   g07004(.A1(new_n4070_), .A2(new_n5398_), .B1(new_n5336_), .B2(new_n5917_), .ZN(new_n7078_));
  AOI21_X1   g07005(.A1(new_n7078_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n7079_));
  XOR2_X1    g07006(.A1(new_n4927_), .A2(new_n7079_), .Z(new_n7080_));
  INV_X1     g07007(.I(new_n7080_), .ZN(new_n7081_));
  NOR2_X1    g07008(.A1(new_n7077_), .A2(new_n7081_), .ZN(new_n7082_));
  INV_X1     g07009(.I(new_n7082_), .ZN(new_n7083_));
  NAND2_X1   g07010(.A1(new_n7074_), .A2(new_n7083_), .ZN(new_n7084_));
  NAND2_X1   g07011(.A1(new_n7077_), .A2(new_n7081_), .ZN(new_n7085_));
  NAND2_X1   g07012(.A1(new_n7084_), .A2(new_n7085_), .ZN(new_n7086_));
  INV_X1     g07013(.I(new_n7086_), .ZN(new_n7087_));
  AOI22_X1   g07014(.A1(new_n4347_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4036_), .ZN(new_n7088_));
  OAI21_X1   g07015(.A1(new_n7088_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7089_));
  XOR2_X1    g07016(.A1(new_n4672_), .A2(new_n7089_), .Z(new_n7090_));
  NOR2_X1    g07017(.A1(new_n7087_), .A2(new_n7090_), .ZN(new_n7091_));
  NAND2_X1   g07018(.A1(new_n7087_), .A2(new_n7090_), .ZN(new_n7092_));
  XOR2_X1    g07019(.A1(new_n6720_), .A2(new_n6489_), .Z(new_n7093_));
  XOR2_X1    g07020(.A1(new_n7093_), .A2(new_n6723_), .Z(new_n7094_));
  AOI21_X1   g07021(.A1(new_n7092_), .A2(new_n7094_), .B(new_n7091_), .ZN(new_n7095_));
  AOI22_X1   g07022(.A1(new_n4445_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4399_), .ZN(new_n7096_));
  OAI21_X1   g07023(.A1(new_n7096_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7097_));
  XOR2_X1    g07024(.A1(new_n4403_), .A2(new_n7097_), .Z(new_n7098_));
  NAND2_X1   g07025(.A1(new_n7095_), .A2(new_n7098_), .ZN(new_n7099_));
  NAND2_X1   g07026(.A1(new_n6832_), .A2(new_n7099_), .ZN(new_n7100_));
  OR2_X2     g07027(.A1(new_n7095_), .A2(new_n7098_), .Z(new_n7101_));
  NAND2_X1   g07028(.A1(new_n7100_), .A2(new_n7101_), .ZN(new_n7102_));
  XOR2_X1    g07029(.A1(new_n6484_), .A2(new_n6736_), .Z(new_n7103_));
  OAI22_X1   g07030(.A1(new_n2258_), .A2(new_n4468_), .B1(new_n4501_), .B2(new_n6756_), .ZN(new_n7104_));
  OAI21_X1   g07031(.A1(new_n4516_), .A2(new_n1078_), .B(new_n7104_), .ZN(new_n7105_));
  AOI21_X1   g07032(.A1(new_n7105_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n7106_));
  XOR2_X1    g07033(.A1(new_n4524_), .A2(new_n7106_), .Z(new_n7107_));
  XOR2_X1    g07034(.A1(new_n7103_), .A2(new_n7107_), .Z(new_n7108_));
  XOR2_X1    g07035(.A1(new_n7108_), .A2(new_n7102_), .Z(new_n7109_));
  XOR2_X1    g07036(.A1(new_n7109_), .A2(new_n6741_), .Z(new_n7110_));
  NAND2_X1   g07037(.A1(new_n7101_), .A2(new_n7099_), .ZN(new_n7111_));
  NAND2_X1   g07038(.A1(new_n6832_), .A2(new_n7111_), .ZN(new_n7112_));
  XNOR2_X1   g07039(.A1(new_n7095_), .A2(new_n7098_), .ZN(new_n7113_));
  OAI21_X1   g07040(.A1(new_n6832_), .A2(new_n7113_), .B(new_n7112_), .ZN(new_n7114_));
  XNOR2_X1   g07041(.A1(new_n7090_), .A2(new_n7093_), .ZN(new_n7115_));
  XOR2_X1    g07042(.A1(new_n7115_), .A2(new_n7086_), .Z(new_n7116_));
  XOR2_X1    g07043(.A1(new_n7116_), .A2(new_n6724_), .Z(new_n7117_));
  INV_X1     g07044(.I(new_n7117_), .ZN(new_n7118_));
  XOR2_X1    g07045(.A1(new_n7077_), .A2(new_n7080_), .Z(new_n7119_));
  AOI21_X1   g07046(.A1(new_n7072_), .A2(new_n7073_), .B(new_n7119_), .ZN(new_n7120_));
  AOI21_X1   g07047(.A1(new_n7083_), .A2(new_n7085_), .B(new_n7074_), .ZN(new_n7121_));
  NOR2_X1    g07048(.A1(new_n7120_), .A2(new_n7121_), .ZN(new_n7122_));
  INV_X1     g07049(.I(new_n7122_), .ZN(new_n7123_));
  XNOR2_X1   g07050(.A1(new_n7050_), .A2(new_n7053_), .ZN(new_n7124_));
  NOR2_X1    g07051(.A1(new_n7124_), .A2(new_n7056_), .ZN(new_n7125_));
  INV_X1     g07052(.I(new_n7054_), .ZN(new_n7126_));
  INV_X1     g07053(.I(new_n7056_), .ZN(new_n7127_));
  AOI21_X1   g07054(.A1(new_n7126_), .A2(new_n7057_), .B(new_n7127_), .ZN(new_n7128_));
  NOR2_X1    g07055(.A1(new_n7125_), .A2(new_n7128_), .ZN(new_n7129_));
  AOI22_X1   g07056(.A1(new_n4923_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4061_), .ZN(new_n7130_));
  OAI21_X1   g07057(.A1(new_n7130_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7131_));
  XOR2_X1    g07058(.A1(new_n4935_), .A2(new_n7131_), .Z(new_n7132_));
  NAND2_X1   g07059(.A1(new_n7129_), .A2(new_n7132_), .ZN(new_n7133_));
  OR2_X2     g07060(.A1(new_n7129_), .A2(new_n7132_), .Z(new_n7134_));
  NAND2_X1   g07061(.A1(new_n7134_), .A2(new_n7133_), .ZN(new_n7135_));
  OAI21_X1   g07062(.A1(new_n6837_), .A2(new_n6838_), .B(new_n7047_), .ZN(new_n7136_));
  INV_X1     g07063(.I(new_n7136_), .ZN(new_n7137_));
  NAND2_X1   g07064(.A1(new_n7137_), .A2(new_n7039_), .ZN(new_n7138_));
  NAND3_X1   g07065(.A1(new_n7136_), .A2(new_n7009_), .A3(new_n7038_), .ZN(new_n7139_));
  AOI21_X1   g07066(.A1(new_n7138_), .A2(new_n7139_), .B(new_n7043_), .ZN(new_n7140_));
  INV_X1     g07067(.I(new_n7140_), .ZN(new_n7141_));
  NAND3_X1   g07068(.A1(new_n7138_), .A2(new_n7043_), .A3(new_n7139_), .ZN(new_n7142_));
  NAND2_X1   g07069(.A1(new_n7019_), .A2(new_n7020_), .ZN(new_n7143_));
  INV_X1     g07070(.I(new_n7143_), .ZN(new_n7144_));
  NAND2_X1   g07071(.A1(new_n7008_), .A2(new_n7144_), .ZN(new_n7145_));
  NOR2_X1    g07072(.A1(new_n7008_), .A2(new_n7144_), .ZN(new_n7146_));
  INV_X1     g07073(.I(new_n7146_), .ZN(new_n7147_));
  AOI22_X1   g07074(.A1(new_n6419_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4328_), .ZN(new_n7148_));
  OAI21_X1   g07075(.A1(new_n7148_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7149_));
  XNOR2_X1   g07076(.A1(new_n5139_), .A2(new_n7149_), .ZN(new_n7150_));
  NAND3_X1   g07077(.A1(new_n7147_), .A2(new_n7150_), .A3(new_n7145_), .ZN(new_n7151_));
  INV_X1     g07078(.I(new_n7145_), .ZN(new_n7152_));
  INV_X1     g07079(.I(new_n7150_), .ZN(new_n7153_));
  OAI21_X1   g07080(.A1(new_n7152_), .A2(new_n7146_), .B(new_n7153_), .ZN(new_n7154_));
  NAND2_X1   g07081(.A1(new_n7154_), .A2(new_n7151_), .ZN(new_n7155_));
  NAND2_X1   g07082(.A1(new_n6844_), .A2(new_n7005_), .ZN(new_n7156_));
  INV_X1     g07083(.I(new_n7156_), .ZN(new_n7157_));
  NAND2_X1   g07084(.A1(new_n7001_), .A2(new_n7157_), .ZN(new_n7158_));
  INV_X1     g07085(.I(new_n7000_), .ZN(new_n7159_));
  NOR3_X1    g07086(.A1(new_n7159_), .A2(new_n6986_), .A3(new_n6988_), .ZN(new_n7160_));
  NAND2_X1   g07087(.A1(new_n7160_), .A2(new_n7156_), .ZN(new_n7161_));
  AOI21_X1   g07088(.A1(new_n7161_), .A2(new_n7158_), .B(new_n6999_), .ZN(new_n7162_));
  AND3_X2    g07089(.A1(new_n7161_), .A2(new_n6999_), .A3(new_n7158_), .Z(new_n7163_));
  NOR2_X1    g07090(.A1(new_n7163_), .A2(new_n7162_), .ZN(new_n7164_));
  INV_X1     g07091(.I(new_n6971_), .ZN(new_n7165_));
  NAND2_X1   g07092(.A1(new_n6968_), .A2(new_n6616_), .ZN(new_n7166_));
  INV_X1     g07093(.I(new_n7166_), .ZN(new_n7167_));
  NOR2_X1    g07094(.A1(new_n6968_), .A2(new_n6616_), .ZN(new_n7168_));
  OAI21_X1   g07095(.A1(new_n7167_), .A2(new_n7168_), .B(new_n6973_), .ZN(new_n7169_));
  INV_X1     g07096(.I(new_n7168_), .ZN(new_n7170_));
  NAND3_X1   g07097(.A1(new_n7170_), .A2(new_n6603_), .A3(new_n7166_), .ZN(new_n7171_));
  AOI21_X1   g07098(.A1(new_n7169_), .A2(new_n7171_), .B(new_n7165_), .ZN(new_n7172_));
  AOI21_X1   g07099(.A1(new_n7170_), .A2(new_n7166_), .B(new_n6603_), .ZN(new_n7173_));
  NOR3_X1    g07100(.A1(new_n7167_), .A2(new_n6973_), .A3(new_n7168_), .ZN(new_n7174_));
  NOR3_X1    g07101(.A1(new_n7173_), .A2(new_n7174_), .A3(new_n6971_), .ZN(new_n7175_));
  NOR2_X1    g07102(.A1(new_n7172_), .A2(new_n7175_), .ZN(new_n7176_));
  NAND2_X1   g07103(.A1(new_n6957_), .A2(new_n6953_), .ZN(new_n7177_));
  XOR2_X1    g07104(.A1(new_n6955_), .A2(new_n6952_), .Z(new_n7178_));
  NOR2_X1    g07105(.A1(new_n7178_), .A2(new_n6945_), .ZN(new_n7179_));
  AOI21_X1   g07106(.A1(new_n6945_), .A2(new_n7177_), .B(new_n7179_), .ZN(new_n7180_));
  NAND2_X1   g07107(.A1(new_n6609_), .A2(new_n5421_), .ZN(new_n7181_));
  OAI21_X1   g07108(.A1(new_n4135_), .A2(new_n1620_), .B(new_n7181_), .ZN(new_n7182_));
  AOI21_X1   g07109(.A1(new_n7182_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n7183_));
  XNOR2_X1   g07110(.A1(new_n5624_), .A2(new_n7183_), .ZN(new_n7184_));
  NAND2_X1   g07111(.A1(new_n6917_), .A2(new_n6920_), .ZN(new_n7185_));
  XNOR2_X1   g07112(.A1(new_n6927_), .A2(new_n6923_), .ZN(new_n7186_));
  NAND2_X1   g07113(.A1(new_n7186_), .A2(new_n7185_), .ZN(new_n7187_));
  NOR2_X1    g07114(.A1(new_n6931_), .A2(new_n6928_), .ZN(new_n7188_));
  OR2_X2     g07115(.A1(new_n7188_), .A2(new_n7185_), .Z(new_n7189_));
  NAND2_X1   g07116(.A1(new_n7189_), .A2(new_n7187_), .ZN(new_n7190_));
  INV_X1     g07117(.I(new_n7190_), .ZN(new_n7191_));
  AOI21_X1   g07118(.A1(new_n6940_), .A2(new_n6944_), .B(new_n6932_), .ZN(new_n7192_));
  XNOR2_X1   g07119(.A1(new_n6939_), .A2(new_n6942_), .ZN(new_n7193_));
  AOI21_X1   g07120(.A1(new_n6932_), .A2(new_n7193_), .B(new_n7192_), .ZN(new_n7194_));
  OAI22_X1   g07121(.A1(new_n4285_), .A2(new_n1620_), .B1(new_n5420_), .B2(new_n6621_), .ZN(new_n7195_));
  AOI21_X1   g07122(.A1(new_n7195_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n7196_));
  XNOR2_X1   g07123(.A1(new_n5023_), .A2(new_n7196_), .ZN(new_n7197_));
  AND2_X2    g07124(.A1(new_n7194_), .A2(new_n7197_), .Z(new_n7198_));
  NOR2_X1    g07125(.A1(new_n7194_), .A2(new_n7197_), .ZN(new_n7199_));
  NOR2_X1    g07126(.A1(new_n7198_), .A2(new_n7199_), .ZN(new_n7200_));
  OAI21_X1   g07127(.A1(new_n7200_), .A2(new_n7191_), .B(new_n7184_), .ZN(new_n7201_));
  INV_X1     g07128(.I(new_n6889_), .ZN(new_n7202_));
  OAI22_X1   g07129(.A1(new_n6504_), .A2(new_n5420_), .B1(new_n1620_), .B2(new_n4249_), .ZN(new_n7203_));
  NAND2_X1   g07130(.A1(new_n7203_), .A2(new_n126_), .ZN(new_n7204_));
  NAND2_X1   g07131(.A1(new_n7204_), .A2(new_n4660_), .ZN(new_n7205_));
  XOR2_X1    g07132(.A1(new_n7205_), .A2(new_n5648_), .Z(new_n7206_));
  INV_X1     g07133(.I(new_n7206_), .ZN(new_n7207_));
  NAND2_X1   g07134(.A1(new_n7207_), .A2(new_n7202_), .ZN(new_n7208_));
  INV_X1     g07135(.I(new_n7208_), .ZN(new_n7209_));
  NAND2_X1   g07136(.A1(new_n5627_), .A2(new_n1620_), .ZN(new_n7210_));
  AOI21_X1   g07137(.A1(new_n4660_), .A2(new_n6061_), .B(new_n4260_), .ZN(new_n7211_));
  OAI22_X1   g07138(.A1(new_n4244_), .A2(new_n5419_), .B1(new_n1622_), .B2(new_n4230_), .ZN(new_n7212_));
  OAI21_X1   g07139(.A1(new_n1620_), .A2(new_n4234_), .B(new_n7212_), .ZN(new_n7213_));
  AOI21_X1   g07140(.A1(new_n7210_), .A2(new_n7211_), .B(new_n7213_), .ZN(new_n7214_));
  XOR2_X1    g07141(.A1(new_n7214_), .A2(\a[17] ), .Z(new_n7215_));
  NOR2_X1    g07142(.A1(new_n4244_), .A2(new_n1622_), .ZN(new_n7216_));
  OAI21_X1   g07143(.A1(new_n4230_), .A2(new_n1620_), .B(new_n126_), .ZN(new_n7217_));
  OAI21_X1   g07144(.A1(new_n7216_), .A2(new_n7217_), .B(new_n4660_), .ZN(new_n7218_));
  XOR2_X1    g07145(.A1(new_n7218_), .A2(new_n5637_), .Z(new_n7219_));
  NOR2_X1    g07146(.A1(new_n4251_), .A2(new_n1468_), .ZN(new_n7220_));
  NOR2_X1    g07147(.A1(new_n7220_), .A2(new_n126_), .ZN(new_n7221_));
  INV_X1     g07148(.I(new_n7221_), .ZN(new_n7222_));
  NOR2_X1    g07149(.A1(new_n7219_), .A2(new_n7222_), .ZN(new_n7223_));
  NAND2_X1   g07150(.A1(new_n7215_), .A2(new_n7223_), .ZN(new_n7224_));
  NAND2_X1   g07151(.A1(new_n7206_), .A2(new_n6889_), .ZN(new_n7225_));
  AOI21_X1   g07152(.A1(new_n7224_), .A2(new_n7225_), .B(new_n7209_), .ZN(new_n7226_));
  XNOR2_X1   g07153(.A1(new_n6888_), .A2(new_n6890_), .ZN(new_n7227_));
  OAI22_X1   g07154(.A1(new_n4203_), .A2(new_n1620_), .B1(new_n5420_), .B2(new_n6529_), .ZN(new_n7228_));
  AOI21_X1   g07155(.A1(new_n7228_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n7229_));
  XOR2_X1    g07156(.A1(new_n5660_), .A2(new_n7229_), .Z(new_n7230_));
  NOR2_X1    g07157(.A1(new_n7230_), .A2(new_n7227_), .ZN(new_n7231_));
  NOR2_X1    g07158(.A1(new_n7226_), .A2(new_n7231_), .ZN(new_n7232_));
  NAND2_X1   g07159(.A1(new_n7230_), .A2(new_n7227_), .ZN(new_n7233_));
  INV_X1     g07160(.I(new_n7233_), .ZN(new_n7234_));
  NOR2_X1    g07161(.A1(new_n7232_), .A2(new_n7234_), .ZN(new_n7235_));
  XNOR2_X1   g07162(.A1(new_n6884_), .A2(new_n6891_), .ZN(new_n7236_));
  INV_X1     g07163(.I(new_n7236_), .ZN(new_n7237_));
  AOI22_X1   g07164(.A1(new_n4258_), .A2(new_n4660_), .B1(new_n5421_), .B2(new_n6541_), .ZN(new_n7238_));
  OAI21_X1   g07165(.A1(new_n7238_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7239_));
  XOR2_X1    g07166(.A1(new_n5671_), .A2(new_n7239_), .Z(new_n7240_));
  AND2_X2    g07167(.A1(new_n7240_), .A2(new_n7237_), .Z(new_n7241_));
  NOR2_X1    g07168(.A1(new_n7240_), .A2(new_n7237_), .ZN(new_n7242_));
  INV_X1     g07169(.I(new_n7242_), .ZN(new_n7243_));
  OAI21_X1   g07170(.A1(new_n7235_), .A2(new_n7241_), .B(new_n7243_), .ZN(new_n7244_));
  INV_X1     g07171(.I(new_n6892_), .ZN(new_n7245_));
  XOR2_X1    g07172(.A1(new_n6877_), .A2(new_n6520_), .Z(new_n7246_));
  INV_X1     g07173(.I(new_n6878_), .ZN(new_n7247_));
  OAI22_X1   g07174(.A1(new_n7247_), .A2(new_n6893_), .B1(new_n6884_), .B2(new_n6891_), .ZN(new_n7248_));
  OAI21_X1   g07175(.A1(new_n7246_), .A2(new_n7245_), .B(new_n7248_), .ZN(new_n7249_));
  OAI22_X1   g07176(.A1(new_n5684_), .A2(new_n1620_), .B1(new_n6556_), .B2(new_n5420_), .ZN(new_n7250_));
  AOI21_X1   g07177(.A1(new_n7250_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n7251_));
  XOR2_X1    g07178(.A1(new_n6102_), .A2(new_n7251_), .Z(new_n7252_));
  INV_X1     g07179(.I(new_n7252_), .ZN(new_n7253_));
  OR2_X2     g07180(.A1(new_n7253_), .A2(new_n7249_), .Z(new_n7254_));
  NAND2_X1   g07181(.A1(new_n7254_), .A2(new_n7244_), .ZN(new_n7255_));
  NAND2_X1   g07182(.A1(new_n7253_), .A2(new_n7249_), .ZN(new_n7256_));
  INV_X1     g07183(.I(new_n6894_), .ZN(new_n7257_));
  XNOR2_X1   g07184(.A1(new_n6898_), .A2(new_n6895_), .ZN(new_n7258_));
  NOR2_X1    g07185(.A1(new_n7258_), .A2(new_n7257_), .ZN(new_n7259_));
  INV_X1     g07186(.I(new_n6900_), .ZN(new_n7260_));
  AOI21_X1   g07187(.A1(new_n7260_), .A2(new_n6899_), .B(new_n6894_), .ZN(new_n7261_));
  NOR2_X1    g07188(.A1(new_n7259_), .A2(new_n7261_), .ZN(new_n7262_));
  OAI22_X1   g07189(.A1(new_n4150_), .A2(new_n1620_), .B1(new_n6567_), .B2(new_n5420_), .ZN(new_n7263_));
  AOI21_X1   g07190(.A1(new_n7263_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n7264_));
  XOR2_X1    g07191(.A1(new_n5707_), .A2(new_n7264_), .Z(new_n7265_));
  INV_X1     g07192(.I(new_n7265_), .ZN(new_n7266_));
  NOR2_X1    g07193(.A1(new_n7266_), .A2(new_n7262_), .ZN(new_n7267_));
  AOI21_X1   g07194(.A1(new_n7255_), .A2(new_n7256_), .B(new_n7267_), .ZN(new_n7268_));
  INV_X1     g07195(.I(new_n7262_), .ZN(new_n7269_));
  NOR2_X1    g07196(.A1(new_n7269_), .A2(new_n7265_), .ZN(new_n7270_));
  NOR2_X1    g07197(.A1(new_n7268_), .A2(new_n7270_), .ZN(new_n7271_));
  XNOR2_X1   g07198(.A1(new_n6905_), .A2(new_n6902_), .ZN(new_n7272_));
  NOR2_X1    g07199(.A1(new_n7272_), .A2(new_n6901_), .ZN(new_n7273_));
  INV_X1     g07200(.I(new_n6901_), .ZN(new_n7274_));
  INV_X1     g07201(.I(new_n6906_), .ZN(new_n7275_));
  AOI21_X1   g07202(.A1(new_n7275_), .A2(new_n6907_), .B(new_n7274_), .ZN(new_n7276_));
  NOR2_X1    g07203(.A1(new_n7276_), .A2(new_n7273_), .ZN(new_n7277_));
  AOI22_X1   g07204(.A1(new_n6582_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4274_), .ZN(new_n7278_));
  OAI21_X1   g07205(.A1(new_n7278_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7279_));
  XOR2_X1    g07206(.A1(new_n5722_), .A2(new_n7279_), .Z(new_n7280_));
  INV_X1     g07207(.I(new_n7280_), .ZN(new_n7281_));
  NOR2_X1    g07208(.A1(new_n7281_), .A2(new_n7277_), .ZN(new_n7282_));
  INV_X1     g07209(.I(new_n7277_), .ZN(new_n7283_));
  NOR2_X1    g07210(.A1(new_n7283_), .A2(new_n7280_), .ZN(new_n7284_));
  INV_X1     g07211(.I(new_n7284_), .ZN(new_n7285_));
  OAI21_X1   g07212(.A1(new_n7271_), .A2(new_n7282_), .B(new_n7285_), .ZN(new_n7286_));
  INV_X1     g07213(.I(new_n6908_), .ZN(new_n7287_));
  XOR2_X1    g07214(.A1(new_n6915_), .A2(new_n6918_), .Z(new_n7288_));
  NOR2_X1    g07215(.A1(new_n7288_), .A2(new_n7287_), .ZN(new_n7289_));
  AOI21_X1   g07216(.A1(new_n6920_), .A2(new_n6916_), .B(new_n6908_), .ZN(new_n7290_));
  OAI22_X1   g07217(.A1(new_n4142_), .A2(new_n1620_), .B1(new_n4277_), .B2(new_n5420_), .ZN(new_n7291_));
  AOI21_X1   g07218(.A1(new_n7291_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n7292_));
  XOR2_X1    g07219(.A1(new_n6134_), .A2(new_n7292_), .Z(new_n7293_));
  OAI21_X1   g07220(.A1(new_n7289_), .A2(new_n7290_), .B(new_n7293_), .ZN(new_n7294_));
  NAND2_X1   g07221(.A1(new_n7286_), .A2(new_n7294_), .ZN(new_n7295_));
  NOR2_X1    g07222(.A1(new_n7289_), .A2(new_n7290_), .ZN(new_n7296_));
  INV_X1     g07223(.I(new_n7293_), .ZN(new_n7297_));
  NAND2_X1   g07224(.A1(new_n7296_), .A2(new_n7297_), .ZN(new_n7298_));
  AOI22_X1   g07225(.A1(new_n7200_), .A2(new_n7191_), .B1(new_n7295_), .B2(new_n7298_), .ZN(new_n7299_));
  NAND2_X1   g07226(.A1(new_n7299_), .A2(new_n7201_), .ZN(new_n7300_));
  OR2_X2     g07227(.A1(new_n7300_), .A2(new_n7180_), .Z(new_n7301_));
  NAND2_X1   g07228(.A1(new_n7300_), .A2(new_n7180_), .ZN(new_n7302_));
  INV_X1     g07229(.I(new_n7198_), .ZN(new_n7303_));
  AOI22_X1   g07230(.A1(new_n6961_), .A2(new_n5421_), .B1(new_n4297_), .B2(new_n4660_), .ZN(new_n7304_));
  OAI21_X1   g07231(.A1(new_n7304_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7305_));
  XOR2_X1    g07232(.A1(new_n5753_), .A2(new_n7305_), .Z(new_n7306_));
  NOR2_X1    g07233(.A1(new_n7303_), .A2(new_n7306_), .ZN(new_n7307_));
  NAND2_X1   g07234(.A1(new_n7302_), .A2(new_n7307_), .ZN(new_n7308_));
  NAND2_X1   g07235(.A1(new_n6861_), .A2(new_n6854_), .ZN(new_n7309_));
  NOR2_X1    g07236(.A1(new_n6861_), .A2(new_n6854_), .ZN(new_n7310_));
  INV_X1     g07237(.I(new_n7310_), .ZN(new_n7311_));
  AOI22_X1   g07238(.A1(new_n7311_), .A2(new_n7309_), .B1(new_n6954_), .B2(new_n6957_), .ZN(new_n7312_));
  NAND2_X1   g07239(.A1(new_n6954_), .A2(new_n6957_), .ZN(new_n7313_));
  XOR2_X1    g07240(.A1(new_n6854_), .A2(new_n6860_), .Z(new_n7314_));
  NOR2_X1    g07241(.A1(new_n7314_), .A2(new_n7313_), .ZN(new_n7315_));
  NOR2_X1    g07242(.A1(new_n7312_), .A2(new_n7315_), .ZN(new_n7316_));
  OAI22_X1   g07243(.A1(new_n4131_), .A2(new_n1620_), .B1(new_n4301_), .B2(new_n5420_), .ZN(new_n7317_));
  AOI21_X1   g07244(.A1(new_n7317_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n7318_));
  XNOR2_X1   g07245(.A1(new_n5599_), .A2(new_n7318_), .ZN(new_n7319_));
  INV_X1     g07246(.I(new_n7319_), .ZN(new_n7320_));
  NOR2_X1    g07247(.A1(new_n7320_), .A2(new_n7316_), .ZN(new_n7321_));
  AOI21_X1   g07248(.A1(new_n7308_), .A2(new_n7301_), .B(new_n7321_), .ZN(new_n7322_));
  NOR3_X1    g07249(.A1(new_n7312_), .A2(new_n7315_), .A3(new_n7319_), .ZN(new_n7323_));
  NOR2_X1    g07250(.A1(new_n6872_), .A2(new_n7314_), .ZN(new_n7324_));
  XOR2_X1    g07251(.A1(new_n7324_), .A2(new_n7311_), .Z(new_n7325_));
  NOR2_X1    g07252(.A1(new_n7325_), .A2(new_n7313_), .ZN(new_n7326_));
  XOR2_X1    g07253(.A1(new_n7324_), .A2(new_n7310_), .Z(new_n7327_));
  AOI21_X1   g07254(.A1(new_n6954_), .A2(new_n6957_), .B(new_n7327_), .ZN(new_n7328_));
  NOR2_X1    g07255(.A1(new_n7328_), .A2(new_n7326_), .ZN(new_n7329_));
  AOI22_X1   g07256(.A1(new_n6980_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n5041_), .ZN(new_n7330_));
  OAI21_X1   g07257(.A1(new_n7330_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7331_));
  XOR2_X1    g07258(.A1(new_n5049_), .A2(new_n7331_), .Z(new_n7332_));
  INV_X1     g07259(.I(new_n7332_), .ZN(new_n7333_));
  OAI22_X1   g07260(.A1(new_n7329_), .A2(new_n7333_), .B1(new_n7322_), .B2(new_n7323_), .ZN(new_n7334_));
  NOR3_X1    g07261(.A1(new_n7328_), .A2(new_n7326_), .A3(new_n7332_), .ZN(new_n7335_));
  INV_X1     g07262(.I(new_n7335_), .ZN(new_n7336_));
  NOR2_X1    g07263(.A1(new_n6850_), .A2(new_n6964_), .ZN(new_n7337_));
  INV_X1     g07264(.I(new_n7337_), .ZN(new_n7338_));
  AOI21_X1   g07265(.A1(new_n6958_), .A2(new_n6873_), .B(new_n7338_), .ZN(new_n7339_));
  INV_X1     g07266(.I(new_n7339_), .ZN(new_n7340_));
  NAND3_X1   g07267(.A1(new_n6958_), .A2(new_n6873_), .A3(new_n7338_), .ZN(new_n7341_));
  AOI21_X1   g07268(.A1(new_n7340_), .A2(new_n7341_), .B(new_n6870_), .ZN(new_n7342_));
  INV_X1     g07269(.I(new_n6870_), .ZN(new_n7343_));
  NAND2_X1   g07270(.A1(new_n7340_), .A2(new_n7341_), .ZN(new_n7344_));
  NOR2_X1    g07271(.A1(new_n7344_), .A2(new_n7343_), .ZN(new_n7345_));
  NOR2_X1    g07272(.A1(new_n7345_), .A2(new_n7342_), .ZN(new_n7346_));
  AOI22_X1   g07273(.A1(new_n6993_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4124_), .ZN(new_n7347_));
  OAI21_X1   g07274(.A1(new_n7347_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7348_));
  XOR2_X1    g07275(.A1(new_n5067_), .A2(new_n7348_), .Z(new_n7349_));
  NAND2_X1   g07276(.A1(new_n7346_), .A2(new_n7349_), .ZN(new_n7350_));
  INV_X1     g07277(.I(new_n7349_), .ZN(new_n7351_));
  OAI21_X1   g07278(.A1(new_n7345_), .A2(new_n7342_), .B(new_n7351_), .ZN(new_n7352_));
  NAND2_X1   g07279(.A1(new_n7350_), .A2(new_n7352_), .ZN(new_n7353_));
  NAND3_X1   g07280(.A1(new_n7353_), .A2(new_n7334_), .A3(new_n7336_), .ZN(new_n7354_));
  NOR2_X1    g07281(.A1(new_n7176_), .A2(new_n7354_), .ZN(new_n7355_));
  INV_X1     g07282(.I(new_n7355_), .ZN(new_n7356_));
  NOR2_X1    g07283(.A1(new_n7346_), .A2(new_n7351_), .ZN(new_n7357_));
  OAI22_X1   g07284(.A1(new_n4112_), .A2(new_n1620_), .B1(new_n5420_), .B2(new_n6682_), .ZN(new_n7358_));
  AOI21_X1   g07285(.A1(new_n7358_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n7359_));
  XOR2_X1    g07286(.A1(new_n5096_), .A2(new_n7359_), .Z(new_n7360_));
  INV_X1     g07287(.I(new_n7360_), .ZN(new_n7361_));
  NAND2_X1   g07288(.A1(new_n7357_), .A2(new_n7361_), .ZN(new_n7362_));
  AOI21_X1   g07289(.A1(new_n7176_), .A2(new_n7354_), .B(new_n7362_), .ZN(new_n7363_));
  INV_X1     g07290(.I(new_n7363_), .ZN(new_n7364_));
  NAND2_X1   g07291(.A1(new_n7364_), .A2(new_n7356_), .ZN(new_n7365_));
  INV_X1     g07292(.I(new_n6976_), .ZN(new_n7366_));
  OAI21_X1   g07293(.A1(new_n6985_), .A2(new_n6988_), .B(new_n7366_), .ZN(new_n7367_));
  XOR2_X1    g07294(.A1(new_n6979_), .A2(new_n6983_), .Z(new_n7368_));
  NOR2_X1    g07295(.A1(new_n7368_), .A2(new_n7366_), .ZN(new_n7369_));
  INV_X1     g07296(.I(new_n7369_), .ZN(new_n7370_));
  AOI22_X1   g07297(.A1(new_n7015_), .A2(new_n5421_), .B1(new_n4105_), .B2(new_n4660_), .ZN(new_n7371_));
  OAI21_X1   g07298(.A1(new_n7371_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7372_));
  XOR2_X1    g07299(.A1(new_n5121_), .A2(new_n7372_), .Z(new_n7373_));
  NAND3_X1   g07300(.A1(new_n7370_), .A2(new_n7367_), .A3(new_n7373_), .ZN(new_n7374_));
  NOR2_X1    g07301(.A1(new_n6988_), .A2(new_n6985_), .ZN(new_n7375_));
  NOR2_X1    g07302(.A1(new_n7375_), .A2(new_n6976_), .ZN(new_n7376_));
  INV_X1     g07303(.I(new_n7373_), .ZN(new_n7377_));
  OAI21_X1   g07304(.A1(new_n7376_), .A2(new_n7369_), .B(new_n7377_), .ZN(new_n7378_));
  NOR2_X1    g07305(.A1(new_n6989_), .A2(new_n7000_), .ZN(new_n7379_));
  AOI22_X1   g07306(.A1(new_n7021_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4100_), .ZN(new_n7380_));
  OAI21_X1   g07307(.A1(new_n7380_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7381_));
  XOR2_X1    g07308(.A1(new_n5080_), .A2(new_n7381_), .Z(new_n7382_));
  INV_X1     g07309(.I(new_n7382_), .ZN(new_n7383_));
  NOR3_X1    g07310(.A1(new_n7160_), .A2(new_n7379_), .A3(new_n7383_), .ZN(new_n7384_));
  OAI21_X1   g07311(.A1(new_n6986_), .A2(new_n6988_), .B(new_n7159_), .ZN(new_n7385_));
  AOI21_X1   g07312(.A1(new_n7385_), .A2(new_n7001_), .B(new_n7382_), .ZN(new_n7386_));
  NAND2_X1   g07313(.A1(new_n7374_), .A2(new_n7378_), .ZN(new_n7388_));
  NAND2_X1   g07314(.A1(new_n7365_), .A2(new_n7388_), .ZN(new_n7389_));
  NOR2_X1    g07315(.A1(new_n7389_), .A2(new_n7164_), .ZN(new_n7390_));
  OAI22_X1   g07316(.A1(new_n4090_), .A2(new_n1620_), .B1(new_n4320_), .B2(new_n5420_), .ZN(new_n7391_));
  AOI21_X1   g07317(.A1(new_n7391_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n7392_));
  XOR2_X1    g07318(.A1(new_n5196_), .A2(new_n7392_), .Z(new_n7393_));
  INV_X1     g07319(.I(new_n7393_), .ZN(new_n7394_));
  NAND2_X1   g07320(.A1(new_n7384_), .A2(new_n7394_), .ZN(new_n7395_));
  AOI21_X1   g07321(.A1(new_n7389_), .A2(new_n7164_), .B(new_n7395_), .ZN(new_n7396_));
  NOR2_X1    g07322(.A1(new_n7396_), .A2(new_n7390_), .ZN(new_n7397_));
  NAND3_X1   g07323(.A1(new_n7031_), .A2(new_n7036_), .A3(new_n7020_), .ZN(new_n7398_));
  NAND3_X1   g07324(.A1(new_n7008_), .A2(new_n7398_), .A3(new_n7143_), .ZN(new_n7399_));
  INV_X1     g07325(.I(new_n7399_), .ZN(new_n7400_));
  AOI21_X1   g07326(.A1(new_n7398_), .A2(new_n7143_), .B(new_n7008_), .ZN(new_n7401_));
  AOI22_X1   g07327(.A1(new_n4333_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4082_), .ZN(new_n7402_));
  OAI21_X1   g07328(.A1(new_n7402_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7403_));
  XNOR2_X1   g07329(.A1(new_n5162_), .A2(new_n7403_), .ZN(new_n7404_));
  INV_X1     g07330(.I(new_n7404_), .ZN(new_n7405_));
  NOR3_X1    g07331(.A1(new_n7400_), .A2(new_n7401_), .A3(new_n7405_), .ZN(new_n7406_));
  INV_X1     g07332(.I(new_n7401_), .ZN(new_n7407_));
  AOI21_X1   g07333(.A1(new_n7407_), .A2(new_n7399_), .B(new_n7404_), .ZN(new_n7408_));
  NOR2_X1    g07334(.A1(new_n7408_), .A2(new_n7406_), .ZN(new_n7409_));
  OAI21_X1   g07335(.A1(new_n7409_), .A2(new_n7151_), .B(new_n7397_), .ZN(new_n7410_));
  NAND2_X1   g07336(.A1(new_n7410_), .A2(new_n7155_), .ZN(new_n7411_));
  AOI21_X1   g07337(.A1(new_n7141_), .A2(new_n7142_), .B(new_n7411_), .ZN(new_n7412_));
  NAND3_X1   g07338(.A1(new_n7411_), .A2(new_n7141_), .A3(new_n7142_), .ZN(new_n7413_));
  OAI22_X1   g07339(.A1(new_n4070_), .A2(new_n1620_), .B1(new_n5420_), .B2(new_n5917_), .ZN(new_n7414_));
  AOI21_X1   g07340(.A1(new_n7414_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n7415_));
  XOR2_X1    g07341(.A1(new_n4927_), .A2(new_n7415_), .Z(new_n7416_));
  INV_X1     g07342(.I(new_n7416_), .ZN(new_n7417_));
  AND3_X2    g07343(.A1(new_n7413_), .A2(new_n7406_), .A3(new_n7417_), .Z(new_n7418_));
  NOR2_X1    g07344(.A1(new_n7418_), .A2(new_n7412_), .ZN(new_n7419_));
  AOI21_X1   g07345(.A1(new_n7071_), .A2(new_n7073_), .B(new_n7058_), .ZN(new_n7420_));
  NAND2_X1   g07346(.A1(new_n7065_), .A2(new_n7068_), .ZN(new_n7421_));
  OAI21_X1   g07347(.A1(new_n7063_), .A2(new_n7064_), .B(new_n7069_), .ZN(new_n7422_));
  AOI21_X1   g07348(.A1(new_n7421_), .A2(new_n7422_), .B(new_n7059_), .ZN(new_n7423_));
  AOI22_X1   g07349(.A1(new_n6428_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n4054_), .ZN(new_n7424_));
  OAI21_X1   g07350(.A1(new_n7424_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n7425_));
  XOR2_X1    g07351(.A1(new_n4652_), .A2(new_n7425_), .Z(new_n7426_));
  INV_X1     g07352(.I(new_n7426_), .ZN(new_n7427_));
  NOR3_X1    g07353(.A1(new_n7423_), .A2(new_n7420_), .A3(new_n7427_), .ZN(new_n7428_));
  NOR2_X1    g07354(.A1(new_n7423_), .A2(new_n7420_), .ZN(new_n7429_));
  NOR2_X1    g07355(.A1(new_n7429_), .A2(new_n7426_), .ZN(new_n7430_));
  NOR2_X1    g07356(.A1(new_n7430_), .A2(new_n7428_), .ZN(new_n7431_));
  OAI21_X1   g07357(.A1(new_n7431_), .A2(new_n7133_), .B(new_n7419_), .ZN(new_n7432_));
  NAND2_X1   g07358(.A1(new_n7432_), .A2(new_n7135_), .ZN(new_n7433_));
  INV_X1     g07359(.I(new_n7433_), .ZN(new_n7434_));
  OAI22_X1   g07360(.A1(new_n4042_), .A2(new_n1620_), .B1(new_n4342_), .B2(new_n5420_), .ZN(new_n7435_));
  AOI21_X1   g07361(.A1(new_n7435_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n7436_));
  XNOR2_X1   g07362(.A1(new_n4864_), .A2(new_n7436_), .ZN(new_n7437_));
  INV_X1     g07363(.I(new_n7437_), .ZN(new_n7438_));
  NAND2_X1   g07364(.A1(new_n7428_), .A2(new_n7438_), .ZN(new_n7439_));
  AOI21_X1   g07365(.A1(new_n7433_), .A2(new_n7122_), .B(new_n7439_), .ZN(new_n7440_));
  AOI21_X1   g07366(.A1(new_n7123_), .A2(new_n7434_), .B(new_n7440_), .ZN(new_n7441_));
  AOI22_X1   g07367(.A1(new_n5859_), .A2(new_n5968_), .B1(new_n4375_), .B2(new_n785_), .ZN(new_n7442_));
  OAI21_X1   g07368(.A1(new_n7442_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7443_));
  XOR2_X1    g07369(.A1(new_n4730_), .A2(new_n7443_), .Z(new_n7444_));
  NAND2_X1   g07370(.A1(new_n7441_), .A2(new_n7444_), .ZN(new_n7445_));
  NAND2_X1   g07371(.A1(new_n7445_), .A2(new_n7118_), .ZN(new_n7446_));
  OR2_X2     g07372(.A1(new_n7441_), .A2(new_n7444_), .Z(new_n7447_));
  NAND2_X1   g07373(.A1(new_n7446_), .A2(new_n7447_), .ZN(new_n7448_));
  AOI22_X1   g07374(.A1(new_n4473_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4555_), .ZN(new_n7449_));
  OAI21_X1   g07375(.A1(new_n7449_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n7450_));
  XNOR2_X1   g07376(.A1(new_n4584_), .A2(new_n7450_), .ZN(new_n7451_));
  INV_X1     g07377(.I(new_n7451_), .ZN(new_n7452_));
  OAI21_X1   g07378(.A1(new_n7448_), .A2(new_n7452_), .B(new_n7114_), .ZN(new_n7453_));
  NAND2_X1   g07379(.A1(new_n7452_), .A2(new_n7448_), .ZN(new_n7454_));
  NAND2_X1   g07380(.A1(new_n7453_), .A2(new_n7454_), .ZN(new_n7455_));
  NAND2_X1   g07381(.A1(new_n4563_), .A2(new_n5110_), .ZN(new_n7456_));
  NAND2_X1   g07382(.A1(new_n4564_), .A2(new_n5108_), .ZN(new_n7457_));
  AOI22_X1   g07383(.A1(new_n7457_), .A2(new_n7456_), .B1(new_n2469_), .B2(new_n4564_), .ZN(new_n7458_));
  OAI21_X1   g07384(.A1(new_n7458_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n7459_));
  XOR2_X1    g07385(.A1(new_n4609_), .A2(new_n7459_), .Z(new_n7460_));
  INV_X1     g07386(.I(new_n7460_), .ZN(new_n7461_));
  NOR2_X1    g07387(.A1(new_n7455_), .A2(new_n7461_), .ZN(new_n7462_));
  AOI21_X1   g07388(.A1(new_n7453_), .A2(new_n7454_), .B(new_n7460_), .ZN(new_n7463_));
  NOR2_X1    g07389(.A1(new_n7462_), .A2(new_n7463_), .ZN(new_n7464_));
  NOR2_X1    g07390(.A1(new_n7110_), .A2(new_n7464_), .ZN(new_n7465_));
  XOR2_X1    g07391(.A1(new_n7455_), .A2(new_n7460_), .Z(new_n7466_));
  INV_X1     g07392(.I(new_n7466_), .ZN(new_n7467_));
  AOI21_X1   g07393(.A1(new_n7110_), .A2(new_n7467_), .B(new_n7465_), .ZN(new_n7468_));
  NAND3_X1   g07394(.A1(new_n7407_), .A2(new_n7399_), .A3(new_n7404_), .ZN(new_n7469_));
  INV_X1     g07395(.I(new_n7142_), .ZN(new_n7470_));
  OAI21_X1   g07396(.A1(new_n7470_), .A2(new_n7140_), .B(new_n7417_), .ZN(new_n7471_));
  AOI21_X1   g07397(.A1(new_n7155_), .A2(new_n7410_), .B(new_n7471_), .ZN(new_n7472_));
  AOI21_X1   g07398(.A1(new_n7141_), .A2(new_n7142_), .B(new_n7416_), .ZN(new_n7473_));
  NOR2_X1    g07399(.A1(new_n7411_), .A2(new_n7473_), .ZN(new_n7474_));
  OAI21_X1   g07400(.A1(new_n7472_), .A2(new_n7474_), .B(new_n7469_), .ZN(new_n7475_));
  NAND2_X1   g07401(.A1(new_n7411_), .A2(new_n7473_), .ZN(new_n7476_));
  NAND3_X1   g07402(.A1(new_n7471_), .A2(new_n7155_), .A3(new_n7410_), .ZN(new_n7477_));
  NAND3_X1   g07403(.A1(new_n7476_), .A2(new_n7477_), .A3(new_n7406_), .ZN(new_n7478_));
  NAND2_X1   g07404(.A1(new_n7475_), .A2(new_n7478_), .ZN(new_n7479_));
  NAND3_X1   g07405(.A1(new_n7385_), .A2(new_n7001_), .A3(new_n7382_), .ZN(new_n7480_));
  AOI22_X1   g07406(.A1(new_n7364_), .A2(new_n7356_), .B1(new_n7374_), .B2(new_n7378_), .ZN(new_n7481_));
  NOR3_X1    g07407(.A1(new_n7164_), .A2(new_n7481_), .A3(new_n7393_), .ZN(new_n7482_));
  INV_X1     g07408(.I(new_n7162_), .ZN(new_n7483_));
  NAND3_X1   g07409(.A1(new_n7161_), .A2(new_n7158_), .A3(new_n6999_), .ZN(new_n7484_));
  AOI21_X1   g07410(.A1(new_n7483_), .A2(new_n7484_), .B(new_n7393_), .ZN(new_n7485_));
  NOR2_X1    g07411(.A1(new_n7485_), .A2(new_n7389_), .ZN(new_n7486_));
  OAI21_X1   g07412(.A1(new_n7486_), .A2(new_n7482_), .B(new_n7480_), .ZN(new_n7487_));
  NAND2_X1   g07413(.A1(new_n7485_), .A2(new_n7389_), .ZN(new_n7488_));
  OAI21_X1   g07414(.A1(new_n7164_), .A2(new_n7393_), .B(new_n7481_), .ZN(new_n7489_));
  NAND3_X1   g07415(.A1(new_n7488_), .A2(new_n7489_), .A3(new_n7384_), .ZN(new_n7490_));
  NAND2_X1   g07416(.A1(new_n7487_), .A2(new_n7490_), .ZN(new_n7491_));
  INV_X1     g07417(.I(new_n7354_), .ZN(new_n7492_));
  NOR3_X1    g07418(.A1(new_n7492_), .A2(new_n7176_), .A3(new_n7360_), .ZN(new_n7493_));
  OR2_X2     g07419(.A1(new_n7172_), .A2(new_n7175_), .Z(new_n7494_));
  AOI21_X1   g07420(.A1(new_n7494_), .A2(new_n7361_), .B(new_n7354_), .ZN(new_n7495_));
  OAI22_X1   g07421(.A1(new_n7495_), .A2(new_n7493_), .B1(new_n7346_), .B2(new_n7351_), .ZN(new_n7496_));
  NAND3_X1   g07422(.A1(new_n7494_), .A2(new_n7354_), .A3(new_n7361_), .ZN(new_n7497_));
  OAI21_X1   g07423(.A1(new_n7176_), .A2(new_n7360_), .B(new_n7492_), .ZN(new_n7498_));
  NAND3_X1   g07424(.A1(new_n7497_), .A2(new_n7498_), .A3(new_n7357_), .ZN(new_n7499_));
  NAND2_X1   g07425(.A1(new_n7496_), .A2(new_n7499_), .ZN(new_n7500_));
  NAND2_X1   g07426(.A1(new_n7308_), .A2(new_n7301_), .ZN(new_n7501_));
  XNOR2_X1   g07427(.A1(new_n7319_), .A2(new_n7316_), .ZN(new_n7502_));
  NOR2_X1    g07428(.A1(new_n7321_), .A2(new_n7323_), .ZN(new_n7503_));
  NOR2_X1    g07429(.A1(new_n7501_), .A2(new_n7503_), .ZN(new_n7504_));
  AOI21_X1   g07430(.A1(new_n7501_), .A2(new_n7502_), .B(new_n7504_), .ZN(new_n7505_));
  INV_X1     g07431(.I(new_n7286_), .ZN(new_n7506_));
  AOI21_X1   g07432(.A1(new_n7294_), .A2(new_n7298_), .B(new_n7506_), .ZN(new_n7507_));
  XOR2_X1    g07433(.A1(new_n7296_), .A2(new_n7293_), .Z(new_n7508_));
  NOR2_X1    g07434(.A1(new_n7508_), .A2(new_n7286_), .ZN(new_n7509_));
  NOR2_X1    g07435(.A1(new_n7507_), .A2(new_n7509_), .ZN(new_n7510_));
  INV_X1     g07436(.I(new_n7220_), .ZN(new_n7511_));
  OAI22_X1   g07437(.A1(new_n6504_), .A2(new_n5967_), .B1(new_n643_), .B2(new_n4249_), .ZN(new_n7512_));
  AOI21_X1   g07438(.A1(new_n7512_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7513_));
  XOR2_X1    g07439(.A1(new_n5648_), .A2(new_n7513_), .Z(new_n7514_));
  NAND2_X1   g07440(.A1(new_n7514_), .A2(new_n7511_), .ZN(new_n7515_));
  NAND2_X1   g07441(.A1(new_n5627_), .A2(new_n643_), .ZN(new_n7516_));
  AOI21_X1   g07442(.A1(new_n785_), .A2(new_n6061_), .B(new_n4260_), .ZN(new_n7517_));
  OAI22_X1   g07443(.A1(new_n4244_), .A2(new_n5966_), .B1(new_n1851_), .B2(new_n4230_), .ZN(new_n7518_));
  OAI21_X1   g07444(.A1(new_n643_), .A2(new_n4234_), .B(new_n7518_), .ZN(new_n7519_));
  AOI21_X1   g07445(.A1(new_n7516_), .A2(new_n7517_), .B(new_n7519_), .ZN(new_n7520_));
  XOR2_X1    g07446(.A1(new_n7520_), .A2(new_n279_), .Z(new_n7521_));
  NOR2_X1    g07447(.A1(new_n4244_), .A2(new_n1851_), .ZN(new_n7522_));
  OAI21_X1   g07448(.A1(new_n4230_), .A2(new_n643_), .B(new_n279_), .ZN(new_n7523_));
  OAI21_X1   g07449(.A1(new_n7522_), .A2(new_n7523_), .B(new_n785_), .ZN(new_n7524_));
  XNOR2_X1   g07450(.A1(new_n7524_), .A2(new_n5637_), .ZN(new_n7525_));
  NOR2_X1    g07451(.A1(new_n4251_), .A2(new_n1733_), .ZN(new_n7526_));
  NOR2_X1    g07452(.A1(new_n7526_), .A2(new_n279_), .ZN(new_n7527_));
  NAND2_X1   g07453(.A1(new_n7525_), .A2(new_n7527_), .ZN(new_n7528_));
  NOR2_X1    g07454(.A1(new_n7521_), .A2(new_n7528_), .ZN(new_n7529_));
  NOR2_X1    g07455(.A1(new_n7514_), .A2(new_n7511_), .ZN(new_n7530_));
  OAI21_X1   g07456(.A1(new_n7529_), .A2(new_n7530_), .B(new_n7515_), .ZN(new_n7531_));
  XOR2_X1    g07457(.A1(new_n7219_), .A2(new_n7222_), .Z(new_n7532_));
  OAI22_X1   g07458(.A1(new_n4203_), .A2(new_n643_), .B1(new_n5967_), .B2(new_n6529_), .ZN(new_n7533_));
  AOI21_X1   g07459(.A1(new_n7533_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7534_));
  XOR2_X1    g07460(.A1(new_n6082_), .A2(new_n7534_), .Z(new_n7535_));
  NAND2_X1   g07461(.A1(new_n7535_), .A2(new_n7532_), .ZN(new_n7536_));
  NAND2_X1   g07462(.A1(new_n7536_), .A2(new_n7531_), .ZN(new_n7537_));
  INV_X1     g07463(.I(new_n7532_), .ZN(new_n7538_));
  XOR2_X1    g07464(.A1(new_n5660_), .A2(new_n7534_), .Z(new_n7539_));
  NAND2_X1   g07465(.A1(new_n7539_), .A2(new_n7538_), .ZN(new_n7540_));
  NAND2_X1   g07466(.A1(new_n7537_), .A2(new_n7540_), .ZN(new_n7541_));
  AOI22_X1   g07467(.A1(new_n4258_), .A2(new_n785_), .B1(new_n5968_), .B2(new_n6541_), .ZN(new_n7542_));
  OAI21_X1   g07468(.A1(new_n7542_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7543_));
  XOR2_X1    g07469(.A1(new_n6540_), .A2(new_n7543_), .Z(new_n7544_));
  NAND2_X1   g07470(.A1(new_n7541_), .A2(new_n7544_), .ZN(new_n7545_));
  INV_X1     g07471(.I(new_n7224_), .ZN(new_n7546_));
  NOR2_X1    g07472(.A1(new_n7215_), .A2(new_n7223_), .ZN(new_n7547_));
  OAI22_X1   g07473(.A1(new_n7541_), .A2(new_n7544_), .B1(new_n7546_), .B2(new_n7547_), .ZN(new_n7548_));
  NAND2_X1   g07474(.A1(new_n7548_), .A2(new_n7545_), .ZN(new_n7549_));
  XOR2_X1    g07475(.A1(new_n7206_), .A2(new_n6889_), .Z(new_n7550_));
  AOI21_X1   g07476(.A1(new_n7208_), .A2(new_n7225_), .B(new_n7546_), .ZN(new_n7551_));
  AOI21_X1   g07477(.A1(new_n7550_), .A2(new_n7546_), .B(new_n7551_), .ZN(new_n7552_));
  OAI22_X1   g07478(.A1(new_n5684_), .A2(new_n643_), .B1(new_n6556_), .B2(new_n5967_), .ZN(new_n7553_));
  AOI21_X1   g07479(.A1(new_n7553_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7554_));
  XOR2_X1    g07480(.A1(new_n6102_), .A2(new_n7554_), .Z(new_n7555_));
  NAND2_X1   g07481(.A1(new_n7555_), .A2(new_n7552_), .ZN(new_n7556_));
  NAND2_X1   g07482(.A1(new_n7549_), .A2(new_n7556_), .ZN(new_n7557_));
  OR2_X2     g07483(.A1(new_n7555_), .A2(new_n7552_), .Z(new_n7558_));
  XOR2_X1    g07484(.A1(new_n7230_), .A2(new_n7227_), .Z(new_n7559_));
  INV_X1     g07485(.I(new_n7559_), .ZN(new_n7560_));
  OAI21_X1   g07486(.A1(new_n7234_), .A2(new_n7231_), .B(new_n7226_), .ZN(new_n7561_));
  OAI21_X1   g07487(.A1(new_n7560_), .A2(new_n7226_), .B(new_n7561_), .ZN(new_n7562_));
  OAI22_X1   g07488(.A1(new_n4150_), .A2(new_n643_), .B1(new_n6567_), .B2(new_n5967_), .ZN(new_n7563_));
  AOI21_X1   g07489(.A1(new_n7563_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7564_));
  XOR2_X1    g07490(.A1(new_n5707_), .A2(new_n7564_), .Z(new_n7565_));
  AOI22_X1   g07491(.A1(new_n7557_), .A2(new_n7558_), .B1(new_n7562_), .B2(new_n7565_), .ZN(new_n7566_));
  NOR2_X1    g07492(.A1(new_n7562_), .A2(new_n7565_), .ZN(new_n7567_));
  NOR2_X1    g07493(.A1(new_n7566_), .A2(new_n7567_), .ZN(new_n7568_));
  INV_X1     g07494(.I(new_n7568_), .ZN(new_n7569_));
  XOR2_X1    g07495(.A1(new_n7240_), .A2(new_n7236_), .Z(new_n7570_));
  OAI21_X1   g07496(.A1(new_n7241_), .A2(new_n7242_), .B(new_n7235_), .ZN(new_n7571_));
  OAI21_X1   g07497(.A1(new_n7235_), .A2(new_n7570_), .B(new_n7571_), .ZN(new_n7572_));
  AOI22_X1   g07498(.A1(new_n6582_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4274_), .ZN(new_n7573_));
  OAI21_X1   g07499(.A1(new_n7573_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7574_));
  XOR2_X1    g07500(.A1(new_n5722_), .A2(new_n7574_), .Z(new_n7575_));
  NAND2_X1   g07501(.A1(new_n7572_), .A2(new_n7575_), .ZN(new_n7576_));
  NAND2_X1   g07502(.A1(new_n7569_), .A2(new_n7576_), .ZN(new_n7577_));
  OR2_X2     g07503(.A1(new_n7572_), .A2(new_n7575_), .Z(new_n7578_));
  NAND2_X1   g07504(.A1(new_n7577_), .A2(new_n7578_), .ZN(new_n7579_));
  XNOR2_X1   g07505(.A1(new_n7252_), .A2(new_n7249_), .ZN(new_n7580_));
  NAND2_X1   g07506(.A1(new_n7254_), .A2(new_n7256_), .ZN(new_n7581_));
  MUX2_X1    g07507(.I0(new_n7581_), .I1(new_n7580_), .S(new_n7244_), .Z(new_n7582_));
  OAI22_X1   g07508(.A1(new_n4142_), .A2(new_n643_), .B1(new_n4277_), .B2(new_n5967_), .ZN(new_n7583_));
  AOI21_X1   g07509(.A1(new_n7583_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7584_));
  XOR2_X1    g07510(.A1(new_n6134_), .A2(new_n7584_), .Z(new_n7585_));
  NAND2_X1   g07511(.A1(new_n7582_), .A2(new_n7585_), .ZN(new_n7586_));
  NOR2_X1    g07512(.A1(new_n7582_), .A2(new_n7585_), .ZN(new_n7587_));
  AOI21_X1   g07513(.A1(new_n7579_), .A2(new_n7586_), .B(new_n7587_), .ZN(new_n7588_));
  NAND2_X1   g07514(.A1(new_n7255_), .A2(new_n7256_), .ZN(new_n7589_));
  XNOR2_X1   g07515(.A1(new_n7262_), .A2(new_n7265_), .ZN(new_n7590_));
  NOR2_X1    g07516(.A1(new_n7270_), .A2(new_n7267_), .ZN(new_n7591_));
  NOR2_X1    g07517(.A1(new_n7589_), .A2(new_n7591_), .ZN(new_n7592_));
  AOI21_X1   g07518(.A1(new_n7589_), .A2(new_n7590_), .B(new_n7592_), .ZN(new_n7593_));
  NAND2_X1   g07519(.A1(new_n6609_), .A2(new_n5968_), .ZN(new_n7594_));
  OAI21_X1   g07520(.A1(new_n4135_), .A2(new_n643_), .B(new_n7594_), .ZN(new_n7595_));
  AOI21_X1   g07521(.A1(new_n7595_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7596_));
  XNOR2_X1   g07522(.A1(new_n5624_), .A2(new_n7596_), .ZN(new_n7597_));
  INV_X1     g07523(.I(new_n7597_), .ZN(new_n7598_));
  NOR2_X1    g07524(.A1(new_n7598_), .A2(new_n7593_), .ZN(new_n7599_));
  NAND2_X1   g07525(.A1(new_n7598_), .A2(new_n7593_), .ZN(new_n7600_));
  OAI21_X1   g07526(.A1(new_n7588_), .A2(new_n7599_), .B(new_n7600_), .ZN(new_n7601_));
  NOR2_X1    g07527(.A1(new_n7282_), .A2(new_n7284_), .ZN(new_n7602_));
  XOR2_X1    g07528(.A1(new_n7280_), .A2(new_n7277_), .Z(new_n7603_));
  MUX2_X1    g07529(.I0(new_n7602_), .I1(new_n7603_), .S(new_n7271_), .Z(new_n7604_));
  OAI22_X1   g07530(.A1(new_n4285_), .A2(new_n643_), .B1(new_n5967_), .B2(new_n6621_), .ZN(new_n7605_));
  AOI21_X1   g07531(.A1(new_n7605_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7606_));
  XNOR2_X1   g07532(.A1(new_n5023_), .A2(new_n7606_), .ZN(new_n7607_));
  XNOR2_X1   g07533(.A1(new_n7604_), .A2(new_n7607_), .ZN(new_n7608_));
  NOR3_X1    g07534(.A1(new_n7608_), .A2(new_n7510_), .A3(new_n7601_), .ZN(new_n7609_));
  OAI21_X1   g07535(.A1(new_n7608_), .A2(new_n7601_), .B(new_n7510_), .ZN(new_n7610_));
  NAND2_X1   g07536(.A1(new_n7604_), .A2(new_n7607_), .ZN(new_n7611_));
  AOI22_X1   g07537(.A1(new_n6961_), .A2(new_n5968_), .B1(new_n4297_), .B2(new_n785_), .ZN(new_n7612_));
  OAI21_X1   g07538(.A1(new_n7612_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7613_));
  XOR2_X1    g07539(.A1(new_n5753_), .A2(new_n7613_), .Z(new_n7614_));
  NOR2_X1    g07540(.A1(new_n7611_), .A2(new_n7614_), .ZN(new_n7615_));
  AOI21_X1   g07541(.A1(new_n7610_), .A2(new_n7615_), .B(new_n7609_), .ZN(new_n7616_));
  NAND2_X1   g07542(.A1(new_n7191_), .A2(new_n7184_), .ZN(new_n7617_));
  NOR2_X1    g07543(.A1(new_n7191_), .A2(new_n7184_), .ZN(new_n7618_));
  INV_X1     g07544(.I(new_n7618_), .ZN(new_n7619_));
  AOI22_X1   g07545(.A1(new_n7619_), .A2(new_n7617_), .B1(new_n7295_), .B2(new_n7298_), .ZN(new_n7620_));
  NAND2_X1   g07546(.A1(new_n7295_), .A2(new_n7298_), .ZN(new_n7621_));
  XOR2_X1    g07547(.A1(new_n7184_), .A2(new_n7190_), .Z(new_n7622_));
  NOR2_X1    g07548(.A1(new_n7622_), .A2(new_n7621_), .ZN(new_n7623_));
  NOR2_X1    g07549(.A1(new_n7620_), .A2(new_n7623_), .ZN(new_n7624_));
  OAI22_X1   g07550(.A1(new_n4131_), .A2(new_n643_), .B1(new_n4301_), .B2(new_n5967_), .ZN(new_n7625_));
  AOI21_X1   g07551(.A1(new_n7625_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7626_));
  XNOR2_X1   g07552(.A1(new_n5599_), .A2(new_n7626_), .ZN(new_n7627_));
  INV_X1     g07553(.I(new_n7627_), .ZN(new_n7628_));
  NOR2_X1    g07554(.A1(new_n7628_), .A2(new_n7624_), .ZN(new_n7629_));
  NAND2_X1   g07555(.A1(new_n7628_), .A2(new_n7624_), .ZN(new_n7630_));
  OAI21_X1   g07556(.A1(new_n7616_), .A2(new_n7629_), .B(new_n7630_), .ZN(new_n7631_));
  INV_X1     g07557(.I(new_n7631_), .ZN(new_n7632_));
  NOR2_X1    g07558(.A1(new_n7200_), .A2(new_n7622_), .ZN(new_n7633_));
  XOR2_X1    g07559(.A1(new_n7633_), .A2(new_n7618_), .Z(new_n7634_));
  XNOR2_X1   g07560(.A1(new_n7634_), .A2(new_n7621_), .ZN(new_n7635_));
  AOI22_X1   g07561(.A1(new_n6980_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n5041_), .ZN(new_n7636_));
  OAI21_X1   g07562(.A1(new_n7636_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7637_));
  XOR2_X1    g07563(.A1(new_n5049_), .A2(new_n7637_), .Z(new_n7638_));
  INV_X1     g07564(.I(new_n7638_), .ZN(new_n7639_));
  NOR2_X1    g07565(.A1(new_n7635_), .A2(new_n7639_), .ZN(new_n7640_));
  NAND2_X1   g07566(.A1(new_n7635_), .A2(new_n7639_), .ZN(new_n7641_));
  OAI21_X1   g07567(.A1(new_n7632_), .A2(new_n7640_), .B(new_n7641_), .ZN(new_n7642_));
  NOR2_X1    g07568(.A1(new_n7180_), .A2(new_n7306_), .ZN(new_n7643_));
  INV_X1     g07569(.I(new_n7643_), .ZN(new_n7644_));
  AOI21_X1   g07570(.A1(new_n7299_), .A2(new_n7201_), .B(new_n7644_), .ZN(new_n7645_));
  NOR2_X1    g07571(.A1(new_n7300_), .A2(new_n7643_), .ZN(new_n7646_));
  NOR2_X1    g07572(.A1(new_n7646_), .A2(new_n7645_), .ZN(new_n7647_));
  NOR2_X1    g07573(.A1(new_n7647_), .A2(new_n7198_), .ZN(new_n7648_));
  NOR3_X1    g07574(.A1(new_n7646_), .A2(new_n7303_), .A3(new_n7645_), .ZN(new_n7649_));
  NOR2_X1    g07575(.A1(new_n7648_), .A2(new_n7649_), .ZN(new_n7650_));
  AOI22_X1   g07576(.A1(new_n6993_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4124_), .ZN(new_n7651_));
  OAI21_X1   g07577(.A1(new_n7651_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7652_));
  XOR2_X1    g07578(.A1(new_n5067_), .A2(new_n7652_), .Z(new_n7653_));
  INV_X1     g07579(.I(new_n7653_), .ZN(new_n7654_));
  NAND2_X1   g07580(.A1(new_n7650_), .A2(new_n7654_), .ZN(new_n7655_));
  OAI21_X1   g07581(.A1(new_n7648_), .A2(new_n7649_), .B(new_n7653_), .ZN(new_n7656_));
  NAND2_X1   g07582(.A1(new_n7655_), .A2(new_n7656_), .ZN(new_n7657_));
  NOR3_X1    g07583(.A1(new_n7642_), .A2(new_n7657_), .A3(new_n7505_), .ZN(new_n7658_));
  INV_X1     g07584(.I(new_n7505_), .ZN(new_n7659_));
  XOR2_X1    g07585(.A1(new_n7634_), .A2(new_n7621_), .Z(new_n7660_));
  NAND2_X1   g07586(.A1(new_n7660_), .A2(new_n7638_), .ZN(new_n7661_));
  NOR2_X1    g07587(.A1(new_n7660_), .A2(new_n7638_), .ZN(new_n7662_));
  AOI21_X1   g07588(.A1(new_n7631_), .A2(new_n7661_), .B(new_n7662_), .ZN(new_n7663_));
  AND2_X2    g07589(.A1(new_n7655_), .A2(new_n7656_), .Z(new_n7664_));
  AOI21_X1   g07590(.A1(new_n7664_), .A2(new_n7663_), .B(new_n7659_), .ZN(new_n7665_));
  OAI22_X1   g07591(.A1(new_n4112_), .A2(new_n643_), .B1(new_n5967_), .B2(new_n6682_), .ZN(new_n7666_));
  AOI21_X1   g07592(.A1(new_n7666_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7667_));
  XOR2_X1    g07593(.A1(new_n5096_), .A2(new_n7667_), .Z(new_n7668_));
  NOR2_X1    g07594(.A1(new_n7656_), .A2(new_n7668_), .ZN(new_n7669_));
  INV_X1     g07595(.I(new_n7669_), .ZN(new_n7670_));
  NOR2_X1    g07596(.A1(new_n7665_), .A2(new_n7670_), .ZN(new_n7671_));
  NOR2_X1    g07597(.A1(new_n7329_), .A2(new_n7333_), .ZN(new_n7672_));
  OAI22_X1   g07598(.A1(new_n7672_), .A2(new_n7335_), .B1(new_n7322_), .B2(new_n7323_), .ZN(new_n7673_));
  NOR2_X1    g07599(.A1(new_n7322_), .A2(new_n7323_), .ZN(new_n7674_));
  XOR2_X1    g07600(.A1(new_n7329_), .A2(new_n7333_), .Z(new_n7675_));
  NAND2_X1   g07601(.A1(new_n7675_), .A2(new_n7674_), .ZN(new_n7676_));
  AOI22_X1   g07602(.A1(new_n7015_), .A2(new_n5968_), .B1(new_n4105_), .B2(new_n785_), .ZN(new_n7677_));
  OAI21_X1   g07603(.A1(new_n7677_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7678_));
  XOR2_X1    g07604(.A1(new_n5121_), .A2(new_n7678_), .Z(new_n7679_));
  NAND3_X1   g07605(.A1(new_n7676_), .A2(new_n7673_), .A3(new_n7679_), .ZN(new_n7680_));
  OAI21_X1   g07606(.A1(new_n7671_), .A2(new_n7658_), .B(new_n7680_), .ZN(new_n7681_));
  INV_X1     g07607(.I(new_n7673_), .ZN(new_n7682_));
  XOR2_X1    g07608(.A1(new_n7329_), .A2(new_n7332_), .Z(new_n7683_));
  NOR3_X1    g07609(.A1(new_n7683_), .A2(new_n7322_), .A3(new_n7323_), .ZN(new_n7684_));
  INV_X1     g07610(.I(new_n7679_), .ZN(new_n7685_));
  OAI21_X1   g07611(.A1(new_n7684_), .A2(new_n7682_), .B(new_n7685_), .ZN(new_n7686_));
  NAND4_X1   g07612(.A1(new_n7334_), .A2(new_n7350_), .A3(new_n7336_), .A4(new_n7352_), .ZN(new_n7687_));
  INV_X1     g07613(.I(new_n7687_), .ZN(new_n7688_));
  AOI22_X1   g07614(.A1(new_n7334_), .A2(new_n7336_), .B1(new_n7350_), .B2(new_n7352_), .ZN(new_n7689_));
  AOI22_X1   g07615(.A1(new_n7021_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4100_), .ZN(new_n7690_));
  OAI21_X1   g07616(.A1(new_n7690_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7691_));
  XOR2_X1    g07617(.A1(new_n5080_), .A2(new_n7691_), .Z(new_n7692_));
  NOR3_X1    g07618(.A1(new_n7688_), .A2(new_n7689_), .A3(new_n7692_), .ZN(new_n7693_));
  NAND2_X1   g07619(.A1(new_n7334_), .A2(new_n7336_), .ZN(new_n7694_));
  NAND2_X1   g07620(.A1(new_n7694_), .A2(new_n7353_), .ZN(new_n7695_));
  INV_X1     g07621(.I(new_n7692_), .ZN(new_n7696_));
  AOI21_X1   g07622(.A1(new_n7695_), .A2(new_n7687_), .B(new_n7696_), .ZN(new_n7697_));
  NOR2_X1    g07623(.A1(new_n7693_), .A2(new_n7697_), .ZN(new_n7698_));
  NAND3_X1   g07624(.A1(new_n7681_), .A2(new_n7686_), .A3(new_n7698_), .ZN(new_n7699_));
  INV_X1     g07625(.I(new_n7699_), .ZN(new_n7700_));
  NAND2_X1   g07626(.A1(new_n7500_), .A2(new_n7700_), .ZN(new_n7701_));
  NAND3_X1   g07627(.A1(new_n7699_), .A2(new_n7496_), .A3(new_n7499_), .ZN(new_n7702_));
  OAI22_X1   g07628(.A1(new_n4090_), .A2(new_n643_), .B1(new_n4320_), .B2(new_n5967_), .ZN(new_n7703_));
  AOI21_X1   g07629(.A1(new_n7703_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7704_));
  XNOR2_X1   g07630(.A1(new_n5196_), .A2(new_n7704_), .ZN(new_n7705_));
  AND2_X2    g07631(.A1(new_n7697_), .A2(new_n7705_), .Z(new_n7706_));
  NAND2_X1   g07632(.A1(new_n7702_), .A2(new_n7706_), .ZN(new_n7707_));
  NAND2_X1   g07633(.A1(new_n7374_), .A2(new_n7378_), .ZN(new_n7708_));
  NAND3_X1   g07634(.A1(new_n7364_), .A2(new_n7356_), .A3(new_n7708_), .ZN(new_n7709_));
  AOI21_X1   g07635(.A1(new_n7364_), .A2(new_n7356_), .B(new_n7708_), .ZN(new_n7710_));
  INV_X1     g07636(.I(new_n7710_), .ZN(new_n7711_));
  AOI22_X1   g07637(.A1(new_n6419_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4328_), .ZN(new_n7712_));
  OAI21_X1   g07638(.A1(new_n7712_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7713_));
  XNOR2_X1   g07639(.A1(new_n5139_), .A2(new_n7713_), .ZN(new_n7714_));
  INV_X1     g07640(.I(new_n7714_), .ZN(new_n7715_));
  NAND3_X1   g07641(.A1(new_n7711_), .A2(new_n7709_), .A3(new_n7715_), .ZN(new_n7716_));
  INV_X1     g07642(.I(new_n7709_), .ZN(new_n7717_));
  OAI21_X1   g07643(.A1(new_n7717_), .A2(new_n7710_), .B(new_n7714_), .ZN(new_n7718_));
  INV_X1     g07644(.I(new_n7708_), .ZN(new_n7719_));
  NOR3_X1    g07645(.A1(new_n7376_), .A2(new_n7369_), .A3(new_n7377_), .ZN(new_n7720_));
  NOR3_X1    g07646(.A1(new_n7386_), .A2(new_n7384_), .A3(new_n7720_), .ZN(new_n7721_));
  NOR3_X1    g07647(.A1(new_n7365_), .A2(new_n7721_), .A3(new_n7719_), .ZN(new_n7722_));
  OAI21_X1   g07648(.A1(new_n7160_), .A2(new_n7379_), .B(new_n7383_), .ZN(new_n7723_));
  NAND3_X1   g07649(.A1(new_n7480_), .A2(new_n7723_), .A3(new_n7374_), .ZN(new_n7724_));
  AOI22_X1   g07650(.A1(new_n7724_), .A2(new_n7708_), .B1(new_n7356_), .B2(new_n7364_), .ZN(new_n7725_));
  AOI22_X1   g07651(.A1(new_n4333_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4082_), .ZN(new_n7726_));
  OAI21_X1   g07652(.A1(new_n7726_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7727_));
  XNOR2_X1   g07653(.A1(new_n5162_), .A2(new_n7727_), .ZN(new_n7728_));
  NOR3_X1    g07654(.A1(new_n7722_), .A2(new_n7725_), .A3(new_n7728_), .ZN(new_n7729_));
  NAND4_X1   g07655(.A1(new_n7724_), .A2(new_n7356_), .A3(new_n7364_), .A4(new_n7708_), .ZN(new_n7730_));
  OAI22_X1   g07656(.A1(new_n7721_), .A2(new_n7719_), .B1(new_n7355_), .B2(new_n7363_), .ZN(new_n7731_));
  INV_X1     g07657(.I(new_n7728_), .ZN(new_n7732_));
  AOI21_X1   g07658(.A1(new_n7731_), .A2(new_n7730_), .B(new_n7732_), .ZN(new_n7733_));
  AOI22_X1   g07659(.A1(new_n7707_), .A2(new_n7701_), .B1(new_n7718_), .B2(new_n7716_), .ZN(new_n7735_));
  NAND2_X1   g07660(.A1(new_n7491_), .A2(new_n7735_), .ZN(new_n7736_));
  OAI21_X1   g07661(.A1(new_n7722_), .A2(new_n7725_), .B(new_n7728_), .ZN(new_n7737_));
  OAI22_X1   g07662(.A1(new_n4070_), .A2(new_n643_), .B1(new_n5917_), .B2(new_n5967_), .ZN(new_n7738_));
  AOI21_X1   g07663(.A1(new_n7738_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7739_));
  XOR2_X1    g07664(.A1(new_n4927_), .A2(new_n7739_), .Z(new_n7740_));
  NOR2_X1    g07665(.A1(new_n7737_), .A2(new_n7740_), .ZN(new_n7741_));
  OAI21_X1   g07666(.A1(new_n7491_), .A2(new_n7735_), .B(new_n7741_), .ZN(new_n7742_));
  NAND2_X1   g07667(.A1(new_n7742_), .A2(new_n7736_), .ZN(new_n7743_));
  NOR2_X1    g07668(.A1(new_n7397_), .A2(new_n7155_), .ZN(new_n7744_));
  NAND2_X1   g07669(.A1(new_n7397_), .A2(new_n7155_), .ZN(new_n7745_));
  INV_X1     g07670(.I(new_n7745_), .ZN(new_n7746_));
  AOI22_X1   g07671(.A1(new_n4923_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4061_), .ZN(new_n7747_));
  OAI21_X1   g07672(.A1(new_n7747_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7748_));
  XOR2_X1    g07673(.A1(new_n4935_), .A2(new_n7748_), .Z(new_n7749_));
  NOR3_X1    g07674(.A1(new_n7746_), .A2(new_n7744_), .A3(new_n7749_), .ZN(new_n7750_));
  INV_X1     g07675(.I(new_n7744_), .ZN(new_n7751_));
  INV_X1     g07676(.I(new_n7749_), .ZN(new_n7752_));
  AOI21_X1   g07677(.A1(new_n7751_), .A2(new_n7745_), .B(new_n7752_), .ZN(new_n7753_));
  NOR3_X1    g07678(.A1(new_n7152_), .A2(new_n7146_), .A3(new_n7153_), .ZN(new_n7754_));
  NOR3_X1    g07679(.A1(new_n7408_), .A2(new_n7406_), .A3(new_n7754_), .ZN(new_n7755_));
  NOR3_X1    g07680(.A1(new_n7755_), .A2(new_n7155_), .A3(new_n7397_), .ZN(new_n7756_));
  INV_X1     g07681(.I(new_n7155_), .ZN(new_n7757_));
  INV_X1     g07682(.I(new_n7397_), .ZN(new_n7758_));
  OAI21_X1   g07683(.A1(new_n7400_), .A2(new_n7401_), .B(new_n7405_), .ZN(new_n7759_));
  NAND3_X1   g07684(.A1(new_n7469_), .A2(new_n7759_), .A3(new_n7151_), .ZN(new_n7760_));
  AOI21_X1   g07685(.A1(new_n7758_), .A2(new_n7760_), .B(new_n7757_), .ZN(new_n7761_));
  AOI22_X1   g07686(.A1(new_n6428_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4054_), .ZN(new_n7762_));
  OAI21_X1   g07687(.A1(new_n7762_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7763_));
  XOR2_X1    g07688(.A1(new_n4652_), .A2(new_n7763_), .Z(new_n7764_));
  NOR3_X1    g07689(.A1(new_n7761_), .A2(new_n7764_), .A3(new_n7756_), .ZN(new_n7765_));
  NAND3_X1   g07690(.A1(new_n7758_), .A2(new_n7757_), .A3(new_n7760_), .ZN(new_n7766_));
  OAI21_X1   g07691(.A1(new_n7755_), .A2(new_n7397_), .B(new_n7155_), .ZN(new_n7767_));
  INV_X1     g07692(.I(new_n7764_), .ZN(new_n7768_));
  AOI21_X1   g07693(.A1(new_n7766_), .A2(new_n7767_), .B(new_n7768_), .ZN(new_n7769_));
  OAI21_X1   g07694(.A1(new_n7750_), .A2(new_n7753_), .B(new_n7743_), .ZN(new_n7771_));
  INV_X1     g07695(.I(new_n7771_), .ZN(new_n7772_));
  NAND2_X1   g07696(.A1(new_n7479_), .A2(new_n7772_), .ZN(new_n7773_));
  NAND3_X1   g07697(.A1(new_n7771_), .A2(new_n7475_), .A3(new_n7478_), .ZN(new_n7774_));
  OAI22_X1   g07698(.A1(new_n4042_), .A2(new_n643_), .B1(new_n4342_), .B2(new_n5967_), .ZN(new_n7775_));
  AOI21_X1   g07699(.A1(new_n7775_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7776_));
  XOR2_X1    g07700(.A1(new_n4864_), .A2(new_n7776_), .Z(new_n7777_));
  NAND3_X1   g07701(.A1(new_n7774_), .A2(new_n7769_), .A3(new_n7777_), .ZN(new_n7778_));
  NAND2_X1   g07702(.A1(new_n7778_), .A2(new_n7773_), .ZN(new_n7779_));
  INV_X1     g07703(.I(new_n7779_), .ZN(new_n7780_));
  OR2_X2     g07704(.A1(new_n7135_), .A2(new_n7419_), .Z(new_n7781_));
  NAND2_X1   g07705(.A1(new_n7135_), .A2(new_n7419_), .ZN(new_n7782_));
  AOI22_X1   g07706(.A1(new_n4347_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4036_), .ZN(new_n7783_));
  OAI21_X1   g07707(.A1(new_n7783_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7784_));
  XOR2_X1    g07708(.A1(new_n4672_), .A2(new_n7784_), .Z(new_n7785_));
  INV_X1     g07709(.I(new_n7785_), .ZN(new_n7786_));
  AOI21_X1   g07710(.A1(new_n7781_), .A2(new_n7782_), .B(new_n7786_), .ZN(new_n7787_));
  NOR2_X1    g07711(.A1(new_n7787_), .A2(new_n7780_), .ZN(new_n7788_));
  NAND3_X1   g07712(.A1(new_n7781_), .A2(new_n7782_), .A3(new_n7786_), .ZN(new_n7789_));
  INV_X1     g07713(.I(new_n7789_), .ZN(new_n7790_));
  NOR2_X1    g07714(.A1(new_n7788_), .A2(new_n7790_), .ZN(new_n7791_));
  INV_X1     g07715(.I(new_n7133_), .ZN(new_n7792_));
  NOR3_X1    g07716(.A1(new_n7430_), .A2(new_n7792_), .A3(new_n7428_), .ZN(new_n7793_));
  NOR3_X1    g07717(.A1(new_n7793_), .A2(new_n7135_), .A3(new_n7419_), .ZN(new_n7794_));
  INV_X1     g07718(.I(new_n7794_), .ZN(new_n7795_));
  OAI21_X1   g07719(.A1(new_n7793_), .A2(new_n7419_), .B(new_n7135_), .ZN(new_n7796_));
  AOI22_X1   g07720(.A1(new_n5935_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n4029_), .ZN(new_n7797_));
  OAI21_X1   g07721(.A1(new_n7797_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n7798_));
  XOR2_X1    g07722(.A1(new_n4687_), .A2(new_n7798_), .Z(new_n7799_));
  INV_X1     g07723(.I(new_n7799_), .ZN(new_n7800_));
  AOI21_X1   g07724(.A1(new_n7795_), .A2(new_n7796_), .B(new_n7800_), .ZN(new_n7801_));
  INV_X1     g07725(.I(new_n7796_), .ZN(new_n7802_));
  NOR3_X1    g07726(.A1(new_n7802_), .A2(new_n7794_), .A3(new_n7799_), .ZN(new_n7803_));
  INV_X1     g07727(.I(new_n7803_), .ZN(new_n7804_));
  OAI21_X1   g07728(.A1(new_n7791_), .A2(new_n7801_), .B(new_n7804_), .ZN(new_n7805_));
  INV_X1     g07729(.I(new_n7805_), .ZN(new_n7806_));
  NAND3_X1   g07730(.A1(new_n7433_), .A2(new_n7123_), .A3(new_n7438_), .ZN(new_n7807_));
  NAND2_X1   g07731(.A1(new_n7123_), .A2(new_n7438_), .ZN(new_n7808_));
  NAND2_X1   g07732(.A1(new_n7434_), .A2(new_n7808_), .ZN(new_n7809_));
  AOI21_X1   g07733(.A1(new_n7809_), .A2(new_n7807_), .B(new_n7428_), .ZN(new_n7810_));
  INV_X1     g07734(.I(new_n7428_), .ZN(new_n7811_));
  NOR2_X1    g07735(.A1(new_n7434_), .A2(new_n7808_), .ZN(new_n7812_));
  AOI21_X1   g07736(.A1(new_n7123_), .A2(new_n7438_), .B(new_n7433_), .ZN(new_n7813_));
  NOR3_X1    g07737(.A1(new_n7812_), .A2(new_n7813_), .A3(new_n7811_), .ZN(new_n7814_));
  OAI22_X1   g07738(.A1(new_n4028_), .A2(new_n5966_), .B1(new_n1851_), .B2(new_n4035_), .ZN(new_n7815_));
  OAI21_X1   g07739(.A1(new_n4017_), .A2(new_n643_), .B(new_n7815_), .ZN(new_n7816_));
  AOI21_X1   g07740(.A1(new_n7816_), .A2(new_n279_), .B(new_n643_), .ZN(new_n7817_));
  XNOR2_X1   g07741(.A1(new_n4705_), .A2(new_n7817_), .ZN(new_n7818_));
  OAI21_X1   g07742(.A1(new_n7814_), .A2(new_n7810_), .B(new_n7818_), .ZN(new_n7819_));
  INV_X1     g07743(.I(new_n7819_), .ZN(new_n7820_));
  OAI21_X1   g07744(.A1(new_n7812_), .A2(new_n7813_), .B(new_n7811_), .ZN(new_n7821_));
  NAND3_X1   g07745(.A1(new_n7809_), .A2(new_n7428_), .A3(new_n7807_), .ZN(new_n7822_));
  INV_X1     g07746(.I(new_n7818_), .ZN(new_n7823_));
  NAND3_X1   g07747(.A1(new_n7821_), .A2(new_n7822_), .A3(new_n7823_), .ZN(new_n7824_));
  OAI21_X1   g07748(.A1(new_n7820_), .A2(new_n7806_), .B(new_n7824_), .ZN(new_n7825_));
  AOI22_X1   g07749(.A1(new_n4448_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4469_), .ZN(new_n7826_));
  OAI21_X1   g07750(.A1(new_n7826_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n7827_));
  XNOR2_X1   g07751(.A1(new_n4477_), .A2(new_n7827_), .ZN(new_n7828_));
  INV_X1     g07752(.I(new_n7828_), .ZN(new_n7829_));
  AOI21_X1   g07753(.A1(new_n7447_), .A2(new_n7445_), .B(new_n7117_), .ZN(new_n7830_));
  XOR2_X1    g07754(.A1(new_n7441_), .A2(new_n7444_), .Z(new_n7831_));
  AOI21_X1   g07755(.A1(new_n7117_), .A2(new_n7831_), .B(new_n7830_), .ZN(new_n7832_));
  NOR2_X1    g07756(.A1(new_n7825_), .A2(new_n7829_), .ZN(new_n7833_));
  NOR2_X1    g07757(.A1(new_n7833_), .A2(new_n7832_), .ZN(new_n7834_));
  AOI21_X1   g07758(.A1(new_n7825_), .A2(new_n7829_), .B(new_n7834_), .ZN(new_n7835_));
  INV_X1     g07759(.I(new_n5110_), .ZN(new_n7836_));
  NOR2_X1    g07760(.A1(new_n7836_), .A2(new_n2718_), .ZN(new_n7837_));
  INV_X1     g07761(.I(new_n7837_), .ZN(new_n7838_));
  AOI22_X1   g07762(.A1(new_n5418_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4563_), .ZN(new_n7839_));
  OAI21_X1   g07763(.A1(new_n7839_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n7840_));
  XNOR2_X1   g07764(.A1(new_n4594_), .A2(new_n7840_), .ZN(new_n7841_));
  NAND2_X1   g07765(.A1(new_n7835_), .A2(new_n7841_), .ZN(new_n7842_));
  XOR2_X1    g07766(.A1(new_n7114_), .A2(new_n7448_), .Z(new_n7843_));
  XOR2_X1    g07767(.A1(new_n7843_), .A2(new_n7452_), .Z(new_n7844_));
  NAND2_X1   g07768(.A1(new_n7844_), .A2(new_n7842_), .ZN(new_n7845_));
  OAI21_X1   g07769(.A1(new_n7835_), .A2(new_n7841_), .B(new_n7845_), .ZN(new_n7846_));
  NOR2_X1    g07770(.A1(new_n7846_), .A2(new_n2905_), .ZN(new_n7847_));
  NAND2_X1   g07771(.A1(new_n7846_), .A2(new_n2905_), .ZN(new_n7848_));
  OAI21_X1   g07772(.A1(new_n7468_), .A2(new_n7847_), .B(new_n7848_), .ZN(new_n7849_));
  INV_X1     g07773(.I(new_n7463_), .ZN(new_n7850_));
  OAI21_X1   g07774(.A1(new_n7110_), .A2(new_n7462_), .B(new_n7850_), .ZN(new_n7851_));
  AOI22_X1   g07775(.A1(new_n5553_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4564_), .ZN(new_n7852_));
  OAI21_X1   g07776(.A1(new_n7852_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n7853_));
  XOR2_X1    g07777(.A1(new_n4569_), .A2(new_n7853_), .Z(new_n7854_));
  INV_X1     g07778(.I(new_n7102_), .ZN(new_n7855_));
  NOR2_X1    g07779(.A1(new_n7855_), .A2(new_n7107_), .ZN(new_n7856_));
  XOR2_X1    g07780(.A1(new_n7103_), .A2(new_n6740_), .Z(new_n7857_));
  AOI21_X1   g07781(.A1(new_n7855_), .A2(new_n7107_), .B(new_n7857_), .ZN(new_n7858_));
  NOR2_X1    g07782(.A1(new_n7858_), .A2(new_n7856_), .ZN(new_n7859_));
  XOR2_X1    g07783(.A1(new_n6753_), .A2(new_n6748_), .Z(new_n7860_));
  XOR2_X1    g07784(.A1(new_n7860_), .A2(new_n6744_), .Z(new_n7861_));
  XNOR2_X1   g07785(.A1(new_n7861_), .A2(new_n7859_), .ZN(new_n7862_));
  XOR2_X1    g07786(.A1(new_n7862_), .A2(new_n7854_), .Z(new_n7863_));
  NAND2_X1   g07787(.A1(new_n5110_), .A2(new_n2469_), .ZN(new_n7864_));
  OAI21_X1   g07788(.A1(new_n5108_), .A2(new_n7864_), .B(new_n4564_), .ZN(new_n7865_));
  OAI21_X1   g07789(.A1(new_n7865_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n7866_));
  XOR2_X1    g07790(.A1(new_n5001_), .A2(new_n7866_), .Z(new_n7867_));
  XOR2_X1    g07791(.A1(new_n7863_), .A2(new_n7867_), .Z(new_n7868_));
  NAND2_X1   g07792(.A1(new_n7863_), .A2(new_n7867_), .ZN(new_n7869_));
  OR2_X2     g07793(.A1(new_n7863_), .A2(new_n7867_), .Z(new_n7870_));
  NAND2_X1   g07794(.A1(new_n7870_), .A2(new_n7869_), .ZN(new_n7871_));
  MUX2_X1    g07795(.I0(new_n7871_), .I1(new_n7868_), .S(new_n7851_), .Z(new_n7872_));
  NAND2_X1   g07796(.A1(new_n7872_), .A2(new_n7849_), .ZN(new_n7873_));
  NAND3_X1   g07797(.A1(new_n7821_), .A2(new_n7822_), .A3(new_n7818_), .ZN(new_n7874_));
  OAI21_X1   g07798(.A1(new_n7814_), .A2(new_n7810_), .B(new_n7823_), .ZN(new_n7875_));
  AOI21_X1   g07799(.A1(new_n7874_), .A2(new_n7875_), .B(new_n7806_), .ZN(new_n7876_));
  AOI21_X1   g07800(.A1(new_n7819_), .A2(new_n7824_), .B(new_n7805_), .ZN(new_n7877_));
  NOR2_X1    g07801(.A1(new_n7876_), .A2(new_n7877_), .ZN(new_n7878_));
  INV_X1     g07802(.I(new_n7787_), .ZN(new_n7879_));
  AOI21_X1   g07803(.A1(new_n7879_), .A2(new_n7789_), .B(new_n7780_), .ZN(new_n7880_));
  NAND3_X1   g07804(.A1(new_n7781_), .A2(new_n7782_), .A3(new_n7785_), .ZN(new_n7881_));
  NAND2_X1   g07805(.A1(new_n7781_), .A2(new_n7782_), .ZN(new_n7882_));
  NAND2_X1   g07806(.A1(new_n7882_), .A2(new_n7786_), .ZN(new_n7883_));
  AOI21_X1   g07807(.A1(new_n7883_), .A2(new_n7881_), .B(new_n7779_), .ZN(new_n7884_));
  AOI22_X1   g07808(.A1(new_n5859_), .A2(new_n6758_), .B1(new_n4375_), .B2(new_n805_), .ZN(new_n7885_));
  OAI21_X1   g07809(.A1(new_n7885_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n7886_));
  XOR2_X1    g07810(.A1(new_n4730_), .A2(new_n7886_), .Z(new_n7887_));
  INV_X1     g07811(.I(new_n7887_), .ZN(new_n7888_));
  NOR3_X1    g07812(.A1(new_n7880_), .A2(new_n7884_), .A3(new_n7888_), .ZN(new_n7889_));
  OAI21_X1   g07813(.A1(new_n7790_), .A2(new_n7787_), .B(new_n7779_), .ZN(new_n7890_));
  INV_X1     g07814(.I(new_n7884_), .ZN(new_n7891_));
  AOI21_X1   g07815(.A1(new_n7891_), .A2(new_n7890_), .B(new_n7887_), .ZN(new_n7892_));
  NOR2_X1    g07816(.A1(new_n7892_), .A2(new_n7889_), .ZN(new_n7893_));
  NAND3_X1   g07817(.A1(new_n7479_), .A2(new_n7771_), .A3(new_n7777_), .ZN(new_n7894_));
  AOI21_X1   g07818(.A1(new_n7476_), .A2(new_n7477_), .B(new_n7406_), .ZN(new_n7895_));
  NOR3_X1    g07819(.A1(new_n7472_), .A2(new_n7474_), .A3(new_n7469_), .ZN(new_n7896_));
  OAI21_X1   g07820(.A1(new_n7896_), .A2(new_n7895_), .B(new_n7777_), .ZN(new_n7897_));
  NAND2_X1   g07821(.A1(new_n7897_), .A2(new_n7772_), .ZN(new_n7898_));
  AOI21_X1   g07822(.A1(new_n7898_), .A2(new_n7894_), .B(new_n7769_), .ZN(new_n7899_));
  OAI21_X1   g07823(.A1(new_n7761_), .A2(new_n7756_), .B(new_n7764_), .ZN(new_n7900_));
  NOR2_X1    g07824(.A1(new_n7897_), .A2(new_n7772_), .ZN(new_n7901_));
  AOI21_X1   g07825(.A1(new_n7479_), .A2(new_n7777_), .B(new_n7771_), .ZN(new_n7902_));
  NOR3_X1    g07826(.A1(new_n7901_), .A2(new_n7902_), .A3(new_n7900_), .ZN(new_n7903_));
  NOR2_X1    g07827(.A1(new_n7903_), .A2(new_n7899_), .ZN(new_n7904_));
  NAND3_X1   g07828(.A1(new_n7751_), .A2(new_n7752_), .A3(new_n7745_), .ZN(new_n7905_));
  OAI21_X1   g07829(.A1(new_n7746_), .A2(new_n7744_), .B(new_n7749_), .ZN(new_n7906_));
  NAND2_X1   g07830(.A1(new_n7906_), .A2(new_n7905_), .ZN(new_n7907_));
  NOR2_X1    g07831(.A1(new_n7907_), .A2(new_n7743_), .ZN(new_n7908_));
  INV_X1     g07832(.I(new_n7743_), .ZN(new_n7909_));
  NOR2_X1    g07833(.A1(new_n7753_), .A2(new_n7750_), .ZN(new_n7910_));
  NOR2_X1    g07834(.A1(new_n7909_), .A2(new_n7910_), .ZN(new_n7911_));
  AOI22_X1   g07835(.A1(new_n4347_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4036_), .ZN(new_n7912_));
  OAI21_X1   g07836(.A1(new_n7912_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n7913_));
  XNOR2_X1   g07837(.A1(new_n4672_), .A2(new_n7913_), .ZN(new_n7914_));
  NOR3_X1    g07838(.A1(new_n7911_), .A2(new_n7908_), .A3(new_n7914_), .ZN(new_n7915_));
  NAND2_X1   g07839(.A1(new_n7909_), .A2(new_n7910_), .ZN(new_n7916_));
  NAND2_X1   g07840(.A1(new_n7907_), .A2(new_n7743_), .ZN(new_n7917_));
  XOR2_X1    g07841(.A1(new_n4672_), .A2(new_n7913_), .Z(new_n7918_));
  AOI21_X1   g07842(.A1(new_n7916_), .A2(new_n7917_), .B(new_n7918_), .ZN(new_n7919_));
  OR2_X2     g07843(.A1(new_n7915_), .A2(new_n7919_), .Z(new_n7920_));
  INV_X1     g07844(.I(new_n7735_), .ZN(new_n7921_));
  INV_X1     g07845(.I(new_n7740_), .ZN(new_n7922_));
  NAND3_X1   g07846(.A1(new_n7921_), .A2(new_n7491_), .A3(new_n7922_), .ZN(new_n7923_));
  AOI21_X1   g07847(.A1(new_n7488_), .A2(new_n7489_), .B(new_n7384_), .ZN(new_n7924_));
  NOR3_X1    g07848(.A1(new_n7486_), .A2(new_n7482_), .A3(new_n7480_), .ZN(new_n7925_));
  OAI21_X1   g07849(.A1(new_n7924_), .A2(new_n7925_), .B(new_n7922_), .ZN(new_n7926_));
  NAND2_X1   g07850(.A1(new_n7926_), .A2(new_n7735_), .ZN(new_n7927_));
  AOI21_X1   g07851(.A1(new_n7923_), .A2(new_n7927_), .B(new_n7733_), .ZN(new_n7928_));
  NOR2_X1    g07852(.A1(new_n7926_), .A2(new_n7735_), .ZN(new_n7929_));
  AOI21_X1   g07853(.A1(new_n7491_), .A2(new_n7922_), .B(new_n7921_), .ZN(new_n7930_));
  NOR3_X1    g07854(.A1(new_n7930_), .A2(new_n7737_), .A3(new_n7929_), .ZN(new_n7931_));
  NOR2_X1    g07855(.A1(new_n7931_), .A2(new_n7928_), .ZN(new_n7932_));
  AOI21_X1   g07856(.A1(new_n7496_), .A2(new_n7499_), .B(new_n7699_), .ZN(new_n7933_));
  AOI21_X1   g07857(.A1(new_n7702_), .A2(new_n7706_), .B(new_n7933_), .ZN(new_n7934_));
  NOR3_X1    g07858(.A1(new_n7717_), .A2(new_n7710_), .A3(new_n7714_), .ZN(new_n7935_));
  AOI21_X1   g07859(.A1(new_n7711_), .A2(new_n7709_), .B(new_n7715_), .ZN(new_n7936_));
  NOR2_X1    g07860(.A1(new_n7936_), .A2(new_n7935_), .ZN(new_n7937_));
  NAND2_X1   g07861(.A1(new_n7937_), .A2(new_n7934_), .ZN(new_n7938_));
  NAND2_X1   g07862(.A1(new_n7707_), .A2(new_n7701_), .ZN(new_n7939_));
  NAND2_X1   g07863(.A1(new_n7718_), .A2(new_n7716_), .ZN(new_n7940_));
  NAND2_X1   g07864(.A1(new_n7939_), .A2(new_n7940_), .ZN(new_n7941_));
  AOI22_X1   g07865(.A1(new_n4923_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4061_), .ZN(new_n7942_));
  OAI21_X1   g07866(.A1(new_n7942_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n7943_));
  NOR2_X1    g07867(.A1(new_n4935_), .A2(new_n7943_), .ZN(new_n7944_));
  AND2_X2    g07868(.A1(new_n4935_), .A2(new_n7943_), .Z(new_n7945_));
  NOR2_X1    g07869(.A1(new_n7945_), .A2(new_n7944_), .ZN(new_n7946_));
  NAND3_X1   g07870(.A1(new_n7941_), .A2(new_n7938_), .A3(new_n7946_), .ZN(new_n7947_));
  NOR2_X1    g07871(.A1(new_n7939_), .A2(new_n7940_), .ZN(new_n7948_));
  NOR2_X1    g07872(.A1(new_n7937_), .A2(new_n7934_), .ZN(new_n7949_));
  INV_X1     g07873(.I(new_n7946_), .ZN(new_n7950_));
  OAI21_X1   g07874(.A1(new_n7948_), .A2(new_n7949_), .B(new_n7950_), .ZN(new_n7951_));
  NAND2_X1   g07875(.A1(new_n7951_), .A2(new_n7947_), .ZN(new_n7952_));
  INV_X1     g07876(.I(new_n7697_), .ZN(new_n7953_));
  AOI21_X1   g07877(.A1(new_n7497_), .A2(new_n7498_), .B(new_n7357_), .ZN(new_n7954_));
  NOR4_X1    g07878(.A1(new_n7495_), .A2(new_n7346_), .A3(new_n7493_), .A4(new_n7351_), .ZN(new_n7955_));
  OAI21_X1   g07879(.A1(new_n7955_), .A2(new_n7954_), .B(new_n7705_), .ZN(new_n7956_));
  NOR2_X1    g07880(.A1(new_n7956_), .A2(new_n7700_), .ZN(new_n7957_));
  AOI21_X1   g07881(.A1(new_n7500_), .A2(new_n7705_), .B(new_n7699_), .ZN(new_n7958_));
  OAI21_X1   g07882(.A1(new_n7957_), .A2(new_n7958_), .B(new_n7953_), .ZN(new_n7959_));
  NAND3_X1   g07883(.A1(new_n7500_), .A2(new_n7699_), .A3(new_n7705_), .ZN(new_n7960_));
  NAND2_X1   g07884(.A1(new_n7956_), .A2(new_n7700_), .ZN(new_n7961_));
  NAND3_X1   g07885(.A1(new_n7961_), .A2(new_n7960_), .A3(new_n7697_), .ZN(new_n7962_));
  NAND2_X1   g07886(.A1(new_n7959_), .A2(new_n7962_), .ZN(new_n7963_));
  NOR2_X1    g07887(.A1(new_n7642_), .A2(new_n7657_), .ZN(new_n7964_));
  NOR2_X1    g07888(.A1(new_n7505_), .A2(new_n7668_), .ZN(new_n7965_));
  INV_X1     g07889(.I(new_n7965_), .ZN(new_n7966_));
  NOR2_X1    g07890(.A1(new_n7966_), .A2(new_n7964_), .ZN(new_n7967_));
  NAND2_X1   g07891(.A1(new_n7664_), .A2(new_n7663_), .ZN(new_n7968_));
  NOR2_X1    g07892(.A1(new_n7968_), .A2(new_n7965_), .ZN(new_n7969_));
  OAI21_X1   g07893(.A1(new_n7969_), .A2(new_n7967_), .B(new_n7656_), .ZN(new_n7970_));
  INV_X1     g07894(.I(new_n7656_), .ZN(new_n7971_));
  NAND2_X1   g07895(.A1(new_n7968_), .A2(new_n7965_), .ZN(new_n7972_));
  NAND2_X1   g07896(.A1(new_n7966_), .A2(new_n7964_), .ZN(new_n7973_));
  NAND3_X1   g07897(.A1(new_n7972_), .A2(new_n7973_), .A3(new_n7971_), .ZN(new_n7974_));
  NAND2_X1   g07898(.A1(new_n7970_), .A2(new_n7974_), .ZN(new_n7975_));
  XOR2_X1    g07899(.A1(new_n7627_), .A2(new_n7624_), .Z(new_n7976_));
  INV_X1     g07900(.I(new_n7630_), .ZN(new_n7977_));
  NOR2_X1    g07901(.A1(new_n7977_), .A2(new_n7629_), .ZN(new_n7978_));
  MUX2_X1    g07902(.I0(new_n7976_), .I1(new_n7978_), .S(new_n7616_), .Z(new_n7979_));
  INV_X1     g07903(.I(new_n7586_), .ZN(new_n7980_));
  OAI21_X1   g07904(.A1(new_n7980_), .A2(new_n7587_), .B(new_n7579_), .ZN(new_n7981_));
  XOR2_X1    g07905(.A1(new_n7582_), .A2(new_n7585_), .Z(new_n7982_));
  NAND3_X1   g07906(.A1(new_n7982_), .A2(new_n7577_), .A3(new_n7578_), .ZN(new_n7983_));
  NAND2_X1   g07907(.A1(new_n7981_), .A2(new_n7983_), .ZN(new_n7984_));
  INV_X1     g07908(.I(new_n7984_), .ZN(new_n7985_));
  OAI22_X1   g07909(.A1(new_n6504_), .A2(new_n6757_), .B1(new_n1078_), .B2(new_n4249_), .ZN(new_n7986_));
  NAND2_X1   g07910(.A1(new_n7986_), .A2(new_n294_), .ZN(new_n7987_));
  NAND2_X1   g07911(.A1(new_n7987_), .A2(new_n805_), .ZN(new_n7988_));
  XOR2_X1    g07912(.A1(new_n7988_), .A2(new_n5648_), .Z(new_n7989_));
  NOR2_X1    g07913(.A1(new_n7989_), .A2(new_n7526_), .ZN(new_n7990_));
  NAND2_X1   g07914(.A1(new_n5627_), .A2(new_n1078_), .ZN(new_n7991_));
  AOI21_X1   g07915(.A1(new_n805_), .A2(new_n6061_), .B(new_n4260_), .ZN(new_n7992_));
  OAI22_X1   g07916(.A1(new_n4244_), .A2(new_n6756_), .B1(new_n2258_), .B2(new_n4230_), .ZN(new_n7993_));
  OAI21_X1   g07917(.A1(new_n1078_), .A2(new_n4234_), .B(new_n7993_), .ZN(new_n7994_));
  AOI21_X1   g07918(.A1(new_n7991_), .A2(new_n7992_), .B(new_n7994_), .ZN(new_n7995_));
  XOR2_X1    g07919(.A1(new_n7995_), .A2(\a[11] ), .Z(new_n7996_));
  NOR2_X1    g07920(.A1(new_n4244_), .A2(new_n2258_), .ZN(new_n7997_));
  OAI21_X1   g07921(.A1(new_n4230_), .A2(new_n1078_), .B(new_n294_), .ZN(new_n7998_));
  OAI21_X1   g07922(.A1(new_n7997_), .A2(new_n7998_), .B(new_n805_), .ZN(new_n7999_));
  XOR2_X1    g07923(.A1(new_n7999_), .A2(new_n5637_), .Z(new_n8000_));
  NOR2_X1    g07924(.A1(new_n4251_), .A2(new_n2573_), .ZN(new_n8001_));
  NOR2_X1    g07925(.A1(new_n8001_), .A2(new_n294_), .ZN(new_n8002_));
  INV_X1     g07926(.I(new_n8002_), .ZN(new_n8003_));
  NOR2_X1    g07927(.A1(new_n8000_), .A2(new_n8003_), .ZN(new_n8004_));
  NAND2_X1   g07928(.A1(new_n7996_), .A2(new_n8004_), .ZN(new_n8005_));
  NAND2_X1   g07929(.A1(new_n7989_), .A2(new_n7526_), .ZN(new_n8006_));
  AOI21_X1   g07930(.A1(new_n8005_), .A2(new_n8006_), .B(new_n7990_), .ZN(new_n8007_));
  INV_X1     g07931(.I(new_n8007_), .ZN(new_n8008_));
  XNOR2_X1   g07932(.A1(new_n7525_), .A2(new_n7527_), .ZN(new_n8009_));
  INV_X1     g07933(.I(new_n8009_), .ZN(new_n8010_));
  OAI22_X1   g07934(.A1(new_n4203_), .A2(new_n1078_), .B1(new_n6529_), .B2(new_n6757_), .ZN(new_n8011_));
  AOI21_X1   g07935(.A1(new_n8011_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8012_));
  XOR2_X1    g07936(.A1(new_n6082_), .A2(new_n8012_), .Z(new_n8013_));
  NAND2_X1   g07937(.A1(new_n8013_), .A2(new_n8010_), .ZN(new_n8014_));
  NAND2_X1   g07938(.A1(new_n8008_), .A2(new_n8014_), .ZN(new_n8015_));
  XOR2_X1    g07939(.A1(new_n5660_), .A2(new_n8012_), .Z(new_n8016_));
  NAND2_X1   g07940(.A1(new_n8016_), .A2(new_n8009_), .ZN(new_n8017_));
  NAND2_X1   g07941(.A1(new_n8015_), .A2(new_n8017_), .ZN(new_n8018_));
  AOI22_X1   g07942(.A1(new_n4258_), .A2(new_n805_), .B1(new_n6541_), .B2(new_n6758_), .ZN(new_n8019_));
  OAI21_X1   g07943(.A1(new_n8019_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8020_));
  XOR2_X1    g07944(.A1(new_n5671_), .A2(new_n8020_), .Z(new_n8021_));
  INV_X1     g07945(.I(new_n8021_), .ZN(new_n8022_));
  NAND2_X1   g07946(.A1(new_n8018_), .A2(new_n8022_), .ZN(new_n8023_));
  AND2_X2    g07947(.A1(new_n7521_), .A2(new_n7528_), .Z(new_n8024_));
  OAI22_X1   g07948(.A1(new_n8018_), .A2(new_n8022_), .B1(new_n7529_), .B2(new_n8024_), .ZN(new_n8025_));
  NAND2_X1   g07949(.A1(new_n8025_), .A2(new_n8023_), .ZN(new_n8026_));
  XOR2_X1    g07950(.A1(new_n7514_), .A2(new_n7220_), .Z(new_n8027_));
  INV_X1     g07951(.I(new_n8027_), .ZN(new_n8028_));
  INV_X1     g07952(.I(new_n7530_), .ZN(new_n8029_));
  AOI21_X1   g07953(.A1(new_n8029_), .A2(new_n7515_), .B(new_n7529_), .ZN(new_n8030_));
  AOI21_X1   g07954(.A1(new_n8028_), .A2(new_n7529_), .B(new_n8030_), .ZN(new_n8031_));
  OAI22_X1   g07955(.A1(new_n5684_), .A2(new_n1078_), .B1(new_n6556_), .B2(new_n6757_), .ZN(new_n8032_));
  AOI21_X1   g07956(.A1(new_n8032_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8033_));
  XOR2_X1    g07957(.A1(new_n6102_), .A2(new_n8033_), .Z(new_n8034_));
  NAND2_X1   g07958(.A1(new_n8034_), .A2(new_n8031_), .ZN(new_n8035_));
  NAND2_X1   g07959(.A1(new_n8026_), .A2(new_n8035_), .ZN(new_n8036_));
  OR2_X2     g07960(.A1(new_n8034_), .A2(new_n8031_), .Z(new_n8037_));
  NAND2_X1   g07961(.A1(new_n8036_), .A2(new_n8037_), .ZN(new_n8038_));
  XOR2_X1    g07962(.A1(new_n7539_), .A2(new_n7538_), .Z(new_n8039_));
  AOI21_X1   g07963(.A1(new_n7536_), .A2(new_n7540_), .B(new_n7531_), .ZN(new_n8040_));
  AOI21_X1   g07964(.A1(new_n8039_), .A2(new_n7531_), .B(new_n8040_), .ZN(new_n8041_));
  OAI22_X1   g07965(.A1(new_n4150_), .A2(new_n1078_), .B1(new_n6567_), .B2(new_n6757_), .ZN(new_n8042_));
  AOI21_X1   g07966(.A1(new_n8042_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8043_));
  XNOR2_X1   g07967(.A1(new_n5707_), .A2(new_n8043_), .ZN(new_n8044_));
  NOR2_X1    g07968(.A1(new_n8044_), .A2(new_n8041_), .ZN(new_n8045_));
  INV_X1     g07969(.I(new_n8045_), .ZN(new_n8046_));
  AND2_X2    g07970(.A1(new_n8044_), .A2(new_n8041_), .Z(new_n8047_));
  AOI21_X1   g07971(.A1(new_n8038_), .A2(new_n8046_), .B(new_n8047_), .ZN(new_n8048_));
  INV_X1     g07972(.I(new_n8048_), .ZN(new_n8049_));
  XOR2_X1    g07973(.A1(new_n7541_), .A2(new_n7215_), .Z(new_n8050_));
  XOR2_X1    g07974(.A1(new_n8050_), .A2(new_n7544_), .Z(new_n8051_));
  XNOR2_X1   g07975(.A1(new_n8051_), .A2(new_n7223_), .ZN(new_n8052_));
  AOI22_X1   g07976(.A1(new_n6582_), .A2(new_n6758_), .B1(new_n4274_), .B2(new_n805_), .ZN(new_n8053_));
  OAI21_X1   g07977(.A1(new_n8053_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8054_));
  XOR2_X1    g07978(.A1(new_n5722_), .A2(new_n8054_), .Z(new_n8055_));
  NAND2_X1   g07979(.A1(new_n8052_), .A2(new_n8055_), .ZN(new_n8056_));
  NOR2_X1    g07980(.A1(new_n8052_), .A2(new_n8055_), .ZN(new_n8057_));
  AOI21_X1   g07981(.A1(new_n8049_), .A2(new_n8056_), .B(new_n8057_), .ZN(new_n8058_));
  XNOR2_X1   g07982(.A1(new_n7555_), .A2(new_n7552_), .ZN(new_n8059_));
  AOI21_X1   g07983(.A1(new_n7545_), .A2(new_n7548_), .B(new_n8059_), .ZN(new_n8060_));
  AOI21_X1   g07984(.A1(new_n7556_), .A2(new_n7558_), .B(new_n7549_), .ZN(new_n8061_));
  NOR2_X1    g07985(.A1(new_n8060_), .A2(new_n8061_), .ZN(new_n8062_));
  OAI22_X1   g07986(.A1(new_n4142_), .A2(new_n1078_), .B1(new_n4277_), .B2(new_n6757_), .ZN(new_n8063_));
  AOI21_X1   g07987(.A1(new_n8063_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8064_));
  XOR2_X1    g07988(.A1(new_n6134_), .A2(new_n8064_), .Z(new_n8065_));
  INV_X1     g07989(.I(new_n8065_), .ZN(new_n8066_));
  NOR2_X1    g07990(.A1(new_n8062_), .A2(new_n8066_), .ZN(new_n8067_));
  NOR2_X1    g07991(.A1(new_n8058_), .A2(new_n8067_), .ZN(new_n8068_));
  NOR3_X1    g07992(.A1(new_n8060_), .A2(new_n8061_), .A3(new_n8065_), .ZN(new_n8069_));
  NAND2_X1   g07993(.A1(new_n7557_), .A2(new_n7558_), .ZN(new_n8070_));
  XOR2_X1    g07994(.A1(new_n7562_), .A2(new_n7565_), .Z(new_n8071_));
  NAND2_X1   g07995(.A1(new_n7562_), .A2(new_n7565_), .ZN(new_n8072_));
  INV_X1     g07996(.I(new_n7567_), .ZN(new_n8073_));
  AOI21_X1   g07997(.A1(new_n8072_), .A2(new_n8073_), .B(new_n8070_), .ZN(new_n8074_));
  AOI21_X1   g07998(.A1(new_n8070_), .A2(new_n8071_), .B(new_n8074_), .ZN(new_n8075_));
  NAND2_X1   g07999(.A1(new_n6609_), .A2(new_n6758_), .ZN(new_n8076_));
  OAI21_X1   g08000(.A1(new_n4135_), .A2(new_n1078_), .B(new_n8076_), .ZN(new_n8077_));
  AOI21_X1   g08001(.A1(new_n8077_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8078_));
  XNOR2_X1   g08002(.A1(new_n5624_), .A2(new_n8078_), .ZN(new_n8079_));
  INV_X1     g08003(.I(new_n8079_), .ZN(new_n8080_));
  OAI22_X1   g08004(.A1(new_n8068_), .A2(new_n8069_), .B1(new_n8075_), .B2(new_n8080_), .ZN(new_n8081_));
  INV_X1     g08005(.I(new_n8075_), .ZN(new_n8082_));
  NOR2_X1    g08006(.A1(new_n8082_), .A2(new_n8079_), .ZN(new_n8083_));
  INV_X1     g08007(.I(new_n8083_), .ZN(new_n8084_));
  AOI21_X1   g08008(.A1(new_n7576_), .A2(new_n7578_), .B(new_n7568_), .ZN(new_n8085_));
  XNOR2_X1   g08009(.A1(new_n7572_), .A2(new_n7575_), .ZN(new_n8086_));
  NOR2_X1    g08010(.A1(new_n8086_), .A2(new_n7569_), .ZN(new_n8087_));
  NOR2_X1    g08011(.A1(new_n8087_), .A2(new_n8085_), .ZN(new_n8088_));
  OAI22_X1   g08012(.A1(new_n4285_), .A2(new_n1078_), .B1(new_n6621_), .B2(new_n6757_), .ZN(new_n8089_));
  AOI21_X1   g08013(.A1(new_n8089_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8090_));
  XNOR2_X1   g08014(.A1(new_n5023_), .A2(new_n8090_), .ZN(new_n8091_));
  NAND2_X1   g08015(.A1(new_n8088_), .A2(new_n8091_), .ZN(new_n8092_));
  INV_X1     g08016(.I(new_n8092_), .ZN(new_n8093_));
  NOR2_X1    g08017(.A1(new_n8088_), .A2(new_n8091_), .ZN(new_n8094_));
  NOR2_X1    g08018(.A1(new_n8093_), .A2(new_n8094_), .ZN(new_n8095_));
  NAND3_X1   g08019(.A1(new_n8081_), .A2(new_n8084_), .A3(new_n8095_), .ZN(new_n8096_));
  NOR2_X1    g08020(.A1(new_n8096_), .A2(new_n7985_), .ZN(new_n8097_));
  AOI22_X1   g08021(.A1(new_n6961_), .A2(new_n6758_), .B1(new_n4297_), .B2(new_n805_), .ZN(new_n8098_));
  OAI21_X1   g08022(.A1(new_n8098_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8099_));
  XOR2_X1    g08023(.A1(new_n5753_), .A2(new_n8099_), .Z(new_n8100_));
  NOR2_X1    g08024(.A1(new_n8092_), .A2(new_n8100_), .ZN(new_n8101_));
  INV_X1     g08025(.I(new_n8101_), .ZN(new_n8102_));
  AOI21_X1   g08026(.A1(new_n8096_), .A2(new_n7985_), .B(new_n8102_), .ZN(new_n8103_));
  NOR2_X1    g08027(.A1(new_n8103_), .A2(new_n8097_), .ZN(new_n8104_));
  XOR2_X1    g08028(.A1(new_n7593_), .A2(new_n7597_), .Z(new_n8105_));
  NOR2_X1    g08029(.A1(new_n8105_), .A2(new_n7588_), .ZN(new_n8106_));
  INV_X1     g08030(.I(new_n7599_), .ZN(new_n8107_));
  NAND2_X1   g08031(.A1(new_n8107_), .A2(new_n7600_), .ZN(new_n8108_));
  AOI21_X1   g08032(.A1(new_n7588_), .A2(new_n8108_), .B(new_n8106_), .ZN(new_n8109_));
  OAI22_X1   g08033(.A1(new_n4131_), .A2(new_n1078_), .B1(new_n4301_), .B2(new_n6757_), .ZN(new_n8110_));
  AOI21_X1   g08034(.A1(new_n8110_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8111_));
  XNOR2_X1   g08035(.A1(new_n5599_), .A2(new_n8111_), .ZN(new_n8112_));
  INV_X1     g08036(.I(new_n8112_), .ZN(new_n8113_));
  NOR2_X1    g08037(.A1(new_n8113_), .A2(new_n8109_), .ZN(new_n8114_));
  NAND2_X1   g08038(.A1(new_n8113_), .A2(new_n8109_), .ZN(new_n8115_));
  OAI21_X1   g08039(.A1(new_n8104_), .A2(new_n8114_), .B(new_n8115_), .ZN(new_n8116_));
  XNOR2_X1   g08040(.A1(new_n7608_), .A2(new_n7601_), .ZN(new_n8117_));
  INV_X1     g08041(.I(new_n8117_), .ZN(new_n8118_));
  AOI22_X1   g08042(.A1(new_n6980_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n5041_), .ZN(new_n8119_));
  OAI21_X1   g08043(.A1(new_n8119_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8120_));
  XOR2_X1    g08044(.A1(new_n5049_), .A2(new_n8120_), .Z(new_n8121_));
  NAND2_X1   g08045(.A1(new_n8118_), .A2(new_n8121_), .ZN(new_n8122_));
  NOR2_X1    g08046(.A1(new_n8118_), .A2(new_n8121_), .ZN(new_n8123_));
  AOI21_X1   g08047(.A1(new_n8116_), .A2(new_n8122_), .B(new_n8123_), .ZN(new_n8124_));
  INV_X1     g08048(.I(new_n7611_), .ZN(new_n8125_));
  NOR2_X1    g08049(.A1(new_n7510_), .A2(new_n7614_), .ZN(new_n8126_));
  OAI21_X1   g08050(.A1(new_n7601_), .A2(new_n7608_), .B(new_n8126_), .ZN(new_n8127_));
  NOR3_X1    g08051(.A1(new_n8126_), .A2(new_n7608_), .A3(new_n7601_), .ZN(new_n8128_));
  INV_X1     g08052(.I(new_n8128_), .ZN(new_n8129_));
  AOI21_X1   g08053(.A1(new_n8129_), .A2(new_n8127_), .B(new_n8125_), .ZN(new_n8130_));
  INV_X1     g08054(.I(new_n8130_), .ZN(new_n8131_));
  NAND3_X1   g08055(.A1(new_n8129_), .A2(new_n8125_), .A3(new_n8127_), .ZN(new_n8132_));
  AOI22_X1   g08056(.A1(new_n6993_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4124_), .ZN(new_n8133_));
  OAI21_X1   g08057(.A1(new_n8133_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8134_));
  XOR2_X1    g08058(.A1(new_n5906_), .A2(new_n8134_), .Z(new_n8135_));
  NAND3_X1   g08059(.A1(new_n8135_), .A2(new_n8131_), .A3(new_n8132_), .ZN(new_n8136_));
  INV_X1     g08060(.I(new_n8132_), .ZN(new_n8137_));
  XOR2_X1    g08061(.A1(new_n5067_), .A2(new_n8134_), .Z(new_n8138_));
  OAI21_X1   g08062(.A1(new_n8137_), .A2(new_n8130_), .B(new_n8138_), .ZN(new_n8139_));
  NAND2_X1   g08063(.A1(new_n8139_), .A2(new_n8136_), .ZN(new_n8140_));
  INV_X1     g08064(.I(new_n8140_), .ZN(new_n8141_));
  NAND2_X1   g08065(.A1(new_n8141_), .A2(new_n8124_), .ZN(new_n8142_));
  NOR2_X1    g08066(.A1(new_n8142_), .A2(new_n7979_), .ZN(new_n8143_));
  OAI22_X1   g08067(.A1(new_n4112_), .A2(new_n1078_), .B1(new_n6682_), .B2(new_n6757_), .ZN(new_n8144_));
  AOI21_X1   g08068(.A1(new_n8144_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8145_));
  XOR2_X1    g08069(.A1(new_n5096_), .A2(new_n8145_), .Z(new_n8146_));
  OR2_X2     g08070(.A1(new_n8139_), .A2(new_n8146_), .Z(new_n8147_));
  AOI21_X1   g08071(.A1(new_n8142_), .A2(new_n7979_), .B(new_n8147_), .ZN(new_n8148_));
  AOI21_X1   g08072(.A1(new_n7641_), .A2(new_n7661_), .B(new_n7632_), .ZN(new_n8149_));
  INV_X1     g08073(.I(new_n8149_), .ZN(new_n8150_));
  XOR2_X1    g08074(.A1(new_n7660_), .A2(new_n7638_), .Z(new_n8151_));
  NAND2_X1   g08075(.A1(new_n8151_), .A2(new_n7632_), .ZN(new_n8152_));
  AOI22_X1   g08076(.A1(new_n7015_), .A2(new_n6758_), .B1(new_n4105_), .B2(new_n805_), .ZN(new_n8153_));
  OAI21_X1   g08077(.A1(new_n8153_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8154_));
  XOR2_X1    g08078(.A1(new_n5121_), .A2(new_n8154_), .Z(new_n8155_));
  NAND3_X1   g08079(.A1(new_n8152_), .A2(new_n8150_), .A3(new_n8155_), .ZN(new_n8156_));
  OAI21_X1   g08080(.A1(new_n8148_), .A2(new_n8143_), .B(new_n8156_), .ZN(new_n8157_));
  AOI21_X1   g08081(.A1(new_n8152_), .A2(new_n8150_), .B(new_n8155_), .ZN(new_n8158_));
  INV_X1     g08082(.I(new_n8158_), .ZN(new_n8159_));
  NAND2_X1   g08083(.A1(new_n8157_), .A2(new_n8159_), .ZN(new_n8160_));
  NAND2_X1   g08084(.A1(new_n7642_), .A2(new_n7657_), .ZN(new_n8161_));
  AOI22_X1   g08085(.A1(new_n7021_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4100_), .ZN(new_n8162_));
  OAI21_X1   g08086(.A1(new_n8162_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8163_));
  XOR2_X1    g08087(.A1(new_n5080_), .A2(new_n8163_), .Z(new_n8164_));
  NAND3_X1   g08088(.A1(new_n7968_), .A2(new_n8161_), .A3(new_n8164_), .ZN(new_n8165_));
  NAND2_X1   g08089(.A1(new_n7968_), .A2(new_n8161_), .ZN(new_n8166_));
  INV_X1     g08090(.I(new_n8164_), .ZN(new_n8167_));
  NAND2_X1   g08091(.A1(new_n8166_), .A2(new_n8167_), .ZN(new_n8168_));
  NAND2_X1   g08092(.A1(new_n8168_), .A2(new_n8165_), .ZN(new_n8169_));
  NOR2_X1    g08093(.A1(new_n8160_), .A2(new_n8169_), .ZN(new_n8170_));
  AOI21_X1   g08094(.A1(new_n7972_), .A2(new_n7973_), .B(new_n7971_), .ZN(new_n8171_));
  NOR3_X1    g08095(.A1(new_n7969_), .A2(new_n7656_), .A3(new_n7967_), .ZN(new_n8172_));
  NOR2_X1    g08096(.A1(new_n8172_), .A2(new_n8171_), .ZN(new_n8173_));
  NAND4_X1   g08097(.A1(new_n8157_), .A2(new_n8168_), .A3(new_n8159_), .A4(new_n8165_), .ZN(new_n8174_));
  INV_X1     g08098(.I(new_n8165_), .ZN(new_n8175_));
  OAI22_X1   g08099(.A1(new_n4090_), .A2(new_n1078_), .B1(new_n4320_), .B2(new_n6757_), .ZN(new_n8176_));
  AOI21_X1   g08100(.A1(new_n8176_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8177_));
  XNOR2_X1   g08101(.A1(new_n5196_), .A2(new_n8177_), .ZN(new_n8178_));
  NAND2_X1   g08102(.A1(new_n8175_), .A2(new_n8178_), .ZN(new_n8179_));
  AOI21_X1   g08103(.A1(new_n8174_), .A2(new_n8173_), .B(new_n8179_), .ZN(new_n8180_));
  AOI21_X1   g08104(.A1(new_n7975_), .A2(new_n8170_), .B(new_n8180_), .ZN(new_n8181_));
  NAND3_X1   g08105(.A1(new_n7664_), .A2(new_n7659_), .A3(new_n7663_), .ZN(new_n8182_));
  OAI21_X1   g08106(.A1(new_n7665_), .A2(new_n7670_), .B(new_n8182_), .ZN(new_n8183_));
  OAI21_X1   g08107(.A1(new_n7684_), .A2(new_n7682_), .B(new_n7679_), .ZN(new_n8184_));
  NOR3_X1    g08108(.A1(new_n7684_), .A2(new_n7682_), .A3(new_n7679_), .ZN(new_n8185_));
  INV_X1     g08109(.I(new_n8185_), .ZN(new_n8186_));
  NAND2_X1   g08110(.A1(new_n8186_), .A2(new_n8184_), .ZN(new_n8187_));
  NAND2_X1   g08111(.A1(new_n8187_), .A2(new_n8183_), .ZN(new_n8188_));
  OAI21_X1   g08112(.A1(new_n7642_), .A2(new_n7657_), .B(new_n7505_), .ZN(new_n8189_));
  AOI21_X1   g08113(.A1(new_n8189_), .A2(new_n7669_), .B(new_n7658_), .ZN(new_n8190_));
  NOR3_X1    g08114(.A1(new_n7684_), .A2(new_n7682_), .A3(new_n7685_), .ZN(new_n8191_));
  AOI21_X1   g08115(.A1(new_n7676_), .A2(new_n7673_), .B(new_n7679_), .ZN(new_n8192_));
  OAI21_X1   g08116(.A1(new_n8191_), .A2(new_n8192_), .B(new_n8190_), .ZN(new_n8193_));
  AOI22_X1   g08117(.A1(new_n6419_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4328_), .ZN(new_n8194_));
  OAI21_X1   g08118(.A1(new_n8194_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8195_));
  NOR2_X1    g08119(.A1(new_n5246_), .A2(new_n8195_), .ZN(new_n8196_));
  INV_X1     g08120(.I(new_n8195_), .ZN(new_n8197_));
  NOR2_X1    g08121(.A1(new_n5139_), .A2(new_n8197_), .ZN(new_n8198_));
  NOR2_X1    g08122(.A1(new_n8196_), .A2(new_n8198_), .ZN(new_n8199_));
  INV_X1     g08123(.I(new_n8199_), .ZN(new_n8200_));
  NAND3_X1   g08124(.A1(new_n8188_), .A2(new_n8193_), .A3(new_n8200_), .ZN(new_n8201_));
  AOI21_X1   g08125(.A1(new_n8186_), .A2(new_n8184_), .B(new_n8190_), .ZN(new_n8202_));
  INV_X1     g08126(.I(new_n8193_), .ZN(new_n8203_));
  OAI21_X1   g08127(.A1(new_n8203_), .A2(new_n8202_), .B(new_n8199_), .ZN(new_n8204_));
  OAI21_X1   g08128(.A1(new_n8190_), .A2(new_n8191_), .B(new_n7686_), .ZN(new_n8205_));
  NOR2_X1    g08129(.A1(new_n8205_), .A2(new_n7698_), .ZN(new_n8206_));
  AOI21_X1   g08130(.A1(new_n8183_), .A2(new_n7680_), .B(new_n8192_), .ZN(new_n8207_));
  OR2_X2     g08131(.A1(new_n7693_), .A2(new_n7697_), .Z(new_n8208_));
  NOR2_X1    g08132(.A1(new_n8207_), .A2(new_n8208_), .ZN(new_n8209_));
  AOI22_X1   g08133(.A1(new_n4333_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4082_), .ZN(new_n8210_));
  OAI21_X1   g08134(.A1(new_n8210_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8211_));
  XNOR2_X1   g08135(.A1(new_n5162_), .A2(new_n8211_), .ZN(new_n8212_));
  INV_X1     g08136(.I(new_n8212_), .ZN(new_n8213_));
  NOR3_X1    g08137(.A1(new_n8209_), .A2(new_n8206_), .A3(new_n8213_), .ZN(new_n8214_));
  NAND2_X1   g08138(.A1(new_n8207_), .A2(new_n8208_), .ZN(new_n8215_));
  NAND2_X1   g08139(.A1(new_n8205_), .A2(new_n7698_), .ZN(new_n8216_));
  AOI21_X1   g08140(.A1(new_n8215_), .A2(new_n8216_), .B(new_n8212_), .ZN(new_n8217_));
  AOI21_X1   g08141(.A1(new_n8201_), .A2(new_n8204_), .B(new_n8181_), .ZN(new_n8219_));
  NAND2_X1   g08142(.A1(new_n7963_), .A2(new_n8219_), .ZN(new_n8220_));
  NOR2_X1    g08143(.A1(new_n8148_), .A2(new_n8143_), .ZN(new_n8221_));
  INV_X1     g08144(.I(new_n8221_), .ZN(new_n8222_));
  AOI21_X1   g08145(.A1(new_n8222_), .A2(new_n8156_), .B(new_n8158_), .ZN(new_n8223_));
  AOI21_X1   g08146(.A1(new_n7968_), .A2(new_n8161_), .B(new_n8164_), .ZN(new_n8224_));
  NOR2_X1    g08147(.A1(new_n8175_), .A2(new_n8224_), .ZN(new_n8225_));
  NAND3_X1   g08148(.A1(new_n7975_), .A2(new_n8223_), .A3(new_n8225_), .ZN(new_n8226_));
  AOI21_X1   g08149(.A1(new_n8223_), .A2(new_n8225_), .B(new_n7975_), .ZN(new_n8227_));
  OAI21_X1   g08150(.A1(new_n8227_), .A2(new_n8179_), .B(new_n8226_), .ZN(new_n8228_));
  NOR3_X1    g08151(.A1(new_n8203_), .A2(new_n8202_), .A3(new_n8199_), .ZN(new_n8229_));
  AOI21_X1   g08152(.A1(new_n8188_), .A2(new_n8193_), .B(new_n8200_), .ZN(new_n8230_));
  OAI21_X1   g08153(.A1(new_n8229_), .A2(new_n8230_), .B(new_n8228_), .ZN(new_n8231_));
  NAND3_X1   g08154(.A1(new_n8231_), .A2(new_n7959_), .A3(new_n7962_), .ZN(new_n8232_));
  NAND2_X1   g08155(.A1(new_n8215_), .A2(new_n8216_), .ZN(new_n8233_));
  NAND2_X1   g08156(.A1(new_n8233_), .A2(new_n8212_), .ZN(new_n8234_));
  OAI22_X1   g08157(.A1(new_n4070_), .A2(new_n1078_), .B1(new_n5917_), .B2(new_n6757_), .ZN(new_n8235_));
  AOI21_X1   g08158(.A1(new_n8235_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8236_));
  XOR2_X1    g08159(.A1(new_n4927_), .A2(new_n8236_), .Z(new_n8237_));
  NOR2_X1    g08160(.A1(new_n8234_), .A2(new_n8237_), .ZN(new_n8238_));
  NAND2_X1   g08161(.A1(new_n8232_), .A2(new_n8238_), .ZN(new_n8239_));
  NAND2_X1   g08162(.A1(new_n8239_), .A2(new_n8220_), .ZN(new_n8240_));
  NAND3_X1   g08163(.A1(new_n7731_), .A2(new_n7730_), .A3(new_n7732_), .ZN(new_n8241_));
  NAND3_X1   g08164(.A1(new_n7737_), .A2(new_n8241_), .A3(new_n7718_), .ZN(new_n8242_));
  NAND3_X1   g08165(.A1(new_n8242_), .A2(new_n7934_), .A3(new_n7940_), .ZN(new_n8243_));
  NOR3_X1    g08166(.A1(new_n7729_), .A2(new_n7733_), .A3(new_n7936_), .ZN(new_n8244_));
  OAI21_X1   g08167(.A1(new_n8244_), .A2(new_n7937_), .B(new_n7939_), .ZN(new_n8245_));
  AOI22_X1   g08168(.A1(new_n6428_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4054_), .ZN(new_n8246_));
  OAI21_X1   g08169(.A1(new_n8246_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8247_));
  XOR2_X1    g08170(.A1(new_n4652_), .A2(new_n8247_), .Z(new_n8248_));
  NAND3_X1   g08171(.A1(new_n8245_), .A2(new_n8243_), .A3(new_n8248_), .ZN(new_n8249_));
  NOR3_X1    g08172(.A1(new_n8244_), .A2(new_n7939_), .A3(new_n7937_), .ZN(new_n8250_));
  AOI21_X1   g08173(.A1(new_n8242_), .A2(new_n7940_), .B(new_n7934_), .ZN(new_n8251_));
  INV_X1     g08174(.I(new_n8248_), .ZN(new_n8252_));
  OAI21_X1   g08175(.A1(new_n8250_), .A2(new_n8251_), .B(new_n8252_), .ZN(new_n8253_));
  AOI21_X1   g08176(.A1(new_n8253_), .A2(new_n8249_), .B(new_n7947_), .ZN(new_n8254_));
  OAI21_X1   g08177(.A1(new_n8254_), .A2(new_n8240_), .B(new_n7952_), .ZN(new_n8255_));
  NOR2_X1    g08178(.A1(new_n8255_), .A2(new_n7932_), .ZN(new_n8256_));
  NOR3_X1    g08179(.A1(new_n8250_), .A2(new_n8251_), .A3(new_n8252_), .ZN(new_n8257_));
  OAI22_X1   g08180(.A1(new_n4042_), .A2(new_n1078_), .B1(new_n4342_), .B2(new_n6757_), .ZN(new_n8258_));
  AOI21_X1   g08181(.A1(new_n8258_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8259_));
  INV_X1     g08182(.I(new_n8259_), .ZN(new_n8260_));
  NOR2_X1    g08183(.A1(new_n4864_), .A2(new_n8260_), .ZN(new_n8261_));
  NOR2_X1    g08184(.A1(new_n5217_), .A2(new_n8259_), .ZN(new_n8262_));
  NOR2_X1    g08185(.A1(new_n8262_), .A2(new_n8261_), .ZN(new_n8263_));
  INV_X1     g08186(.I(new_n8263_), .ZN(new_n8264_));
  NAND2_X1   g08187(.A1(new_n8264_), .A2(new_n8257_), .ZN(new_n8265_));
  AOI21_X1   g08188(.A1(new_n8255_), .A2(new_n7932_), .B(new_n8265_), .ZN(new_n8266_));
  NOR2_X1    g08189(.A1(new_n8266_), .A2(new_n8256_), .ZN(new_n8267_));
  NOR3_X1    g08190(.A1(new_n7765_), .A2(new_n7769_), .A3(new_n7753_), .ZN(new_n8268_));
  NOR3_X1    g08191(.A1(new_n8268_), .A2(new_n7743_), .A3(new_n7910_), .ZN(new_n8269_));
  NAND3_X1   g08192(.A1(new_n7766_), .A2(new_n7767_), .A3(new_n7768_), .ZN(new_n8270_));
  NAND3_X1   g08193(.A1(new_n7900_), .A2(new_n8270_), .A3(new_n7906_), .ZN(new_n8271_));
  AOI21_X1   g08194(.A1(new_n8271_), .A2(new_n7907_), .B(new_n7909_), .ZN(new_n8272_));
  AOI22_X1   g08195(.A1(new_n5935_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4029_), .ZN(new_n8273_));
  OAI21_X1   g08196(.A1(new_n8273_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8274_));
  NOR2_X1    g08197(.A1(new_n4687_), .A2(new_n8274_), .ZN(new_n8275_));
  INV_X1     g08198(.I(new_n8274_), .ZN(new_n8276_));
  AOI21_X1   g08199(.A1(new_n4686_), .A2(new_n4683_), .B(new_n8276_), .ZN(new_n8277_));
  NOR2_X1    g08200(.A1(new_n8275_), .A2(new_n8277_), .ZN(new_n8278_));
  INV_X1     g08201(.I(new_n8278_), .ZN(new_n8279_));
  NOR3_X1    g08202(.A1(new_n8269_), .A2(new_n8272_), .A3(new_n8279_), .ZN(new_n8280_));
  NAND3_X1   g08203(.A1(new_n8271_), .A2(new_n7909_), .A3(new_n7907_), .ZN(new_n8281_));
  OAI21_X1   g08204(.A1(new_n8268_), .A2(new_n7910_), .B(new_n7743_), .ZN(new_n8282_));
  AOI21_X1   g08205(.A1(new_n8282_), .A2(new_n8281_), .B(new_n8278_), .ZN(new_n8283_));
  OAI21_X1   g08206(.A1(new_n8280_), .A2(new_n8283_), .B(new_n7915_), .ZN(new_n8284_));
  NAND2_X1   g08207(.A1(new_n8284_), .A2(new_n8267_), .ZN(new_n8285_));
  NAND2_X1   g08208(.A1(new_n8285_), .A2(new_n7920_), .ZN(new_n8286_));
  NOR2_X1    g08209(.A1(new_n8286_), .A2(new_n7904_), .ZN(new_n8287_));
  NAND3_X1   g08210(.A1(new_n8282_), .A2(new_n8281_), .A3(new_n8278_), .ZN(new_n8288_));
  NOR2_X1    g08211(.A1(new_n4028_), .A2(new_n6756_), .ZN(new_n8289_));
  NOR2_X1    g08212(.A1(new_n4035_), .A2(new_n2258_), .ZN(new_n8290_));
  OAI22_X1   g08213(.A1(new_n4017_), .A2(new_n1078_), .B1(new_n8289_), .B2(new_n8290_), .ZN(new_n8291_));
  AOI21_X1   g08214(.A1(new_n8291_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8292_));
  XNOR2_X1   g08215(.A1(new_n4705_), .A2(new_n8292_), .ZN(new_n8293_));
  NOR2_X1    g08216(.A1(new_n8293_), .A2(new_n8288_), .ZN(new_n8294_));
  INV_X1     g08217(.I(new_n8294_), .ZN(new_n8295_));
  AOI21_X1   g08218(.A1(new_n8286_), .A2(new_n7904_), .B(new_n8295_), .ZN(new_n8296_));
  NOR2_X1    g08219(.A1(new_n8296_), .A2(new_n8287_), .ZN(new_n8297_));
  INV_X1     g08220(.I(new_n8297_), .ZN(new_n8298_));
  OAI22_X1   g08221(.A1(new_n7788_), .A2(new_n7790_), .B1(new_n7801_), .B2(new_n7803_), .ZN(new_n8299_));
  NAND3_X1   g08222(.A1(new_n7795_), .A2(new_n7796_), .A3(new_n7799_), .ZN(new_n8300_));
  OAI21_X1   g08223(.A1(new_n7802_), .A2(new_n7794_), .B(new_n7800_), .ZN(new_n8301_));
  NAND2_X1   g08224(.A1(new_n8301_), .A2(new_n8300_), .ZN(new_n8302_));
  NAND2_X1   g08225(.A1(new_n7791_), .A2(new_n8302_), .ZN(new_n8303_));
  AOI22_X1   g08226(.A1(new_n4445_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n4399_), .ZN(new_n8304_));
  OAI21_X1   g08227(.A1(new_n8304_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n8305_));
  XOR2_X1    g08228(.A1(new_n4403_), .A2(new_n8305_), .Z(new_n8306_));
  NAND3_X1   g08229(.A1(new_n8303_), .A2(new_n8299_), .A3(new_n8306_), .ZN(new_n8307_));
  NOR2_X1    g08230(.A1(new_n7801_), .A2(new_n7803_), .ZN(new_n8308_));
  NOR2_X1    g08231(.A1(new_n7791_), .A2(new_n8308_), .ZN(new_n8309_));
  NOR3_X1    g08232(.A1(new_n7802_), .A2(new_n7794_), .A3(new_n7800_), .ZN(new_n8310_));
  AOI21_X1   g08233(.A1(new_n7795_), .A2(new_n7796_), .B(new_n7799_), .ZN(new_n8311_));
  NOR2_X1    g08234(.A1(new_n8311_), .A2(new_n8310_), .ZN(new_n8312_));
  NOR3_X1    g08235(.A1(new_n8312_), .A2(new_n7788_), .A3(new_n7790_), .ZN(new_n8313_));
  INV_X1     g08236(.I(new_n8306_), .ZN(new_n8314_));
  OAI21_X1   g08237(.A1(new_n8313_), .A2(new_n8309_), .B(new_n8314_), .ZN(new_n8315_));
  NAND2_X1   g08238(.A1(new_n8315_), .A2(new_n8307_), .ZN(new_n8316_));
  AOI21_X1   g08239(.A1(new_n8316_), .A2(new_n7889_), .B(new_n8298_), .ZN(new_n8317_));
  NOR2_X1    g08240(.A1(new_n8317_), .A2(new_n7893_), .ZN(new_n8318_));
  INV_X1     g08241(.I(new_n8318_), .ZN(new_n8319_));
  NOR2_X1    g08242(.A1(new_n8319_), .A2(new_n7878_), .ZN(new_n8320_));
  NOR3_X1    g08243(.A1(new_n8313_), .A2(new_n8309_), .A3(new_n8314_), .ZN(new_n8321_));
  OAI22_X1   g08244(.A1(new_n4397_), .A2(new_n6756_), .B1(new_n2258_), .B2(new_n4374_), .ZN(new_n8322_));
  OAI21_X1   g08245(.A1(new_n4437_), .A2(new_n1078_), .B(new_n8322_), .ZN(new_n8323_));
  AOI21_X1   g08246(.A1(new_n8323_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n8324_));
  XOR2_X1    g08247(.A1(new_n4541_), .A2(new_n8324_), .Z(new_n8325_));
  INV_X1     g08248(.I(new_n8325_), .ZN(new_n8326_));
  NAND2_X1   g08249(.A1(new_n8321_), .A2(new_n8326_), .ZN(new_n8327_));
  AOI21_X1   g08250(.A1(new_n8319_), .A2(new_n7878_), .B(new_n8327_), .ZN(new_n8328_));
  NOR2_X1    g08251(.A1(new_n8328_), .A2(new_n8320_), .ZN(new_n8329_));
  XOR2_X1    g08252(.A1(new_n7832_), .A2(new_n7825_), .Z(new_n8330_));
  AOI22_X1   g08253(.A1(new_n5553_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4564_), .ZN(new_n8331_));
  OAI21_X1   g08254(.A1(new_n8331_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8332_));
  XOR2_X1    g08255(.A1(new_n4569_), .A2(new_n8332_), .Z(new_n8333_));
  XOR2_X1    g08256(.A1(new_n8330_), .A2(new_n8333_), .Z(new_n8334_));
  NAND2_X1   g08257(.A1(new_n8334_), .A2(new_n8329_), .ZN(new_n8335_));
  INV_X1     g08258(.I(new_n8335_), .ZN(new_n8336_));
  NOR2_X1    g08259(.A1(new_n8334_), .A2(new_n8329_), .ZN(new_n8337_));
  NOR2_X1    g08260(.A1(new_n8336_), .A2(new_n8337_), .ZN(new_n8338_));
  NOR2_X1    g08261(.A1(new_n8338_), .A2(new_n7829_), .ZN(new_n8339_));
  NOR3_X1    g08262(.A1(new_n8336_), .A2(new_n7828_), .A3(new_n8337_), .ZN(new_n8340_));
  XOR2_X1    g08263(.A1(new_n4705_), .A2(new_n8292_), .Z(new_n8341_));
  OAI21_X1   g08264(.A1(new_n7903_), .A2(new_n7899_), .B(new_n8341_), .ZN(new_n8342_));
  AOI21_X1   g08265(.A1(new_n8285_), .A2(new_n7920_), .B(new_n8342_), .ZN(new_n8343_));
  OAI21_X1   g08266(.A1(new_n7901_), .A2(new_n7902_), .B(new_n7900_), .ZN(new_n8344_));
  NAND3_X1   g08267(.A1(new_n7898_), .A2(new_n7894_), .A3(new_n7769_), .ZN(new_n8345_));
  AOI21_X1   g08268(.A1(new_n8344_), .A2(new_n8345_), .B(new_n8293_), .ZN(new_n8346_));
  NOR2_X1    g08269(.A1(new_n8286_), .A2(new_n8346_), .ZN(new_n8347_));
  OAI21_X1   g08270(.A1(new_n8347_), .A2(new_n8343_), .B(new_n8288_), .ZN(new_n8348_));
  NOR2_X1    g08271(.A1(new_n7915_), .A2(new_n7919_), .ZN(new_n8349_));
  INV_X1     g08272(.I(new_n8267_), .ZN(new_n8350_));
  NAND3_X1   g08273(.A1(new_n7916_), .A2(new_n7917_), .A3(new_n7918_), .ZN(new_n8351_));
  OAI21_X1   g08274(.A1(new_n8269_), .A2(new_n8272_), .B(new_n8279_), .ZN(new_n8352_));
  AOI21_X1   g08275(.A1(new_n8352_), .A2(new_n8288_), .B(new_n8351_), .ZN(new_n8353_));
  NOR2_X1    g08276(.A1(new_n8350_), .A2(new_n8353_), .ZN(new_n8354_));
  OAI21_X1   g08277(.A1(new_n8354_), .A2(new_n8349_), .B(new_n8346_), .ZN(new_n8355_));
  NAND3_X1   g08278(.A1(new_n8342_), .A2(new_n8285_), .A3(new_n7920_), .ZN(new_n8356_));
  NAND3_X1   g08279(.A1(new_n8355_), .A2(new_n8356_), .A3(new_n8280_), .ZN(new_n8357_));
  NAND2_X1   g08280(.A1(new_n8348_), .A2(new_n8357_), .ZN(new_n8358_));
  INV_X1     g08281(.I(new_n8358_), .ZN(new_n8359_));
  OAI21_X1   g08282(.A1(new_n7930_), .A2(new_n7929_), .B(new_n7737_), .ZN(new_n8360_));
  NAND3_X1   g08283(.A1(new_n7923_), .A2(new_n7927_), .A3(new_n7733_), .ZN(new_n8361_));
  AOI21_X1   g08284(.A1(new_n8360_), .A2(new_n8361_), .B(new_n8263_), .ZN(new_n8362_));
  NAND2_X1   g08285(.A1(new_n8255_), .A2(new_n8362_), .ZN(new_n8363_));
  AOI21_X1   g08286(.A1(new_n7959_), .A2(new_n7962_), .B(new_n8231_), .ZN(new_n8364_));
  AOI21_X1   g08287(.A1(new_n8232_), .A2(new_n8238_), .B(new_n8364_), .ZN(new_n8365_));
  NOR3_X1    g08288(.A1(new_n7948_), .A2(new_n7949_), .A3(new_n7950_), .ZN(new_n8366_));
  AOI21_X1   g08289(.A1(new_n8245_), .A2(new_n8243_), .B(new_n8248_), .ZN(new_n8367_));
  OAI21_X1   g08290(.A1(new_n8257_), .A2(new_n8367_), .B(new_n8366_), .ZN(new_n8368_));
  NAND2_X1   g08291(.A1(new_n8368_), .A2(new_n8365_), .ZN(new_n8369_));
  OAI21_X1   g08292(.A1(new_n7931_), .A2(new_n7928_), .B(new_n8264_), .ZN(new_n8370_));
  NAND3_X1   g08293(.A1(new_n8370_), .A2(new_n8369_), .A3(new_n7952_), .ZN(new_n8371_));
  AOI21_X1   g08294(.A1(new_n8371_), .A2(new_n8363_), .B(new_n8257_), .ZN(new_n8372_));
  AOI21_X1   g08295(.A1(new_n8369_), .A2(new_n7952_), .B(new_n8370_), .ZN(new_n8373_));
  NOR2_X1    g08296(.A1(new_n8255_), .A2(new_n8362_), .ZN(new_n8374_));
  NOR3_X1    g08297(.A1(new_n8373_), .A2(new_n8374_), .A3(new_n8249_), .ZN(new_n8375_));
  NOR2_X1    g08298(.A1(new_n8375_), .A2(new_n8372_), .ZN(new_n8376_));
  AOI21_X1   g08299(.A1(new_n7961_), .A2(new_n7960_), .B(new_n7697_), .ZN(new_n8377_));
  NOR3_X1    g08300(.A1(new_n7957_), .A2(new_n7958_), .A3(new_n7953_), .ZN(new_n8378_));
  INV_X1     g08301(.I(new_n8237_), .ZN(new_n8379_));
  OAI21_X1   g08302(.A1(new_n8378_), .A2(new_n8377_), .B(new_n8379_), .ZN(new_n8380_));
  NOR2_X1    g08303(.A1(new_n8380_), .A2(new_n8219_), .ZN(new_n8381_));
  AOI21_X1   g08304(.A1(new_n7963_), .A2(new_n8379_), .B(new_n8231_), .ZN(new_n8382_));
  OAI21_X1   g08305(.A1(new_n8381_), .A2(new_n8382_), .B(new_n8234_), .ZN(new_n8383_));
  INV_X1     g08306(.I(new_n8234_), .ZN(new_n8384_));
  NAND3_X1   g08307(.A1(new_n7963_), .A2(new_n8231_), .A3(new_n8379_), .ZN(new_n8385_));
  NAND2_X1   g08308(.A1(new_n8380_), .A2(new_n8219_), .ZN(new_n8386_));
  NAND3_X1   g08309(.A1(new_n8386_), .A2(new_n8385_), .A3(new_n8384_), .ZN(new_n8387_));
  NAND2_X1   g08310(.A1(new_n8383_), .A2(new_n8387_), .ZN(new_n8388_));
  NAND2_X1   g08311(.A1(new_n8201_), .A2(new_n8204_), .ZN(new_n8389_));
  NOR2_X1    g08312(.A1(new_n8228_), .A2(new_n8389_), .ZN(new_n8390_));
  NOR2_X1    g08313(.A1(new_n8230_), .A2(new_n8229_), .ZN(new_n8391_));
  NOR2_X1    g08314(.A1(new_n8181_), .A2(new_n8391_), .ZN(new_n8392_));
  AOI22_X1   g08315(.A1(new_n4923_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4061_), .ZN(new_n8393_));
  OAI21_X1   g08316(.A1(new_n8393_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8394_));
  NOR2_X1    g08317(.A1(new_n4935_), .A2(new_n8394_), .ZN(new_n8395_));
  AND2_X2    g08318(.A1(new_n4935_), .A2(new_n8394_), .Z(new_n8396_));
  NOR2_X1    g08319(.A1(new_n8396_), .A2(new_n8395_), .ZN(new_n8397_));
  INV_X1     g08320(.I(new_n8397_), .ZN(new_n8398_));
  NOR3_X1    g08321(.A1(new_n8392_), .A2(new_n8390_), .A3(new_n8398_), .ZN(new_n8399_));
  NAND2_X1   g08322(.A1(new_n8181_), .A2(new_n8391_), .ZN(new_n8400_));
  NAND2_X1   g08323(.A1(new_n8228_), .A2(new_n8389_), .ZN(new_n8401_));
  AOI21_X1   g08324(.A1(new_n8400_), .A2(new_n8401_), .B(new_n8397_), .ZN(new_n8402_));
  NOR2_X1    g08325(.A1(new_n8402_), .A2(new_n8399_), .ZN(new_n8403_));
  OAI21_X1   g08326(.A1(new_n8172_), .A2(new_n8171_), .B(new_n8178_), .ZN(new_n8404_));
  NOR2_X1    g08327(.A1(new_n8170_), .A2(new_n8404_), .ZN(new_n8405_));
  AOI21_X1   g08328(.A1(new_n7975_), .A2(new_n8178_), .B(new_n8174_), .ZN(new_n8406_));
  OAI21_X1   g08329(.A1(new_n8405_), .A2(new_n8406_), .B(new_n8165_), .ZN(new_n8407_));
  NAND3_X1   g08330(.A1(new_n8174_), .A2(new_n7975_), .A3(new_n8178_), .ZN(new_n8408_));
  NAND2_X1   g08331(.A1(new_n8170_), .A2(new_n8404_), .ZN(new_n8409_));
  NAND3_X1   g08332(.A1(new_n8409_), .A2(new_n8175_), .A3(new_n8408_), .ZN(new_n8410_));
  NAND2_X1   g08333(.A1(new_n8407_), .A2(new_n8410_), .ZN(new_n8411_));
  NOR2_X1    g08334(.A1(new_n7979_), .A2(new_n8146_), .ZN(new_n8412_));
  NAND2_X1   g08335(.A1(new_n8142_), .A2(new_n8412_), .ZN(new_n8413_));
  OR2_X2     g08336(.A1(new_n8142_), .A2(new_n8412_), .Z(new_n8414_));
  NAND2_X1   g08337(.A1(new_n8414_), .A2(new_n8413_), .ZN(new_n8415_));
  NAND2_X1   g08338(.A1(new_n8415_), .A2(new_n8139_), .ZN(new_n8416_));
  INV_X1     g08339(.I(new_n8139_), .ZN(new_n8417_));
  NAND3_X1   g08340(.A1(new_n8414_), .A2(new_n8417_), .A3(new_n8413_), .ZN(new_n8418_));
  NAND2_X1   g08341(.A1(new_n8416_), .A2(new_n8418_), .ZN(new_n8419_));
  XOR2_X1    g08342(.A1(new_n8109_), .A2(new_n8112_), .Z(new_n8420_));
  OR2_X2     g08343(.A1(new_n8104_), .A2(new_n8420_), .Z(new_n8421_));
  INV_X1     g08344(.I(new_n8115_), .ZN(new_n8422_));
  OAI21_X1   g08345(.A1(new_n8114_), .A2(new_n8422_), .B(new_n8104_), .ZN(new_n8423_));
  NAND2_X1   g08346(.A1(new_n8421_), .A2(new_n8423_), .ZN(new_n8424_));
  XOR2_X1    g08347(.A1(new_n8051_), .A2(new_n7223_), .Z(new_n8425_));
  INV_X1     g08348(.I(new_n8055_), .ZN(new_n8426_));
  NOR2_X1    g08349(.A1(new_n8425_), .A2(new_n8426_), .ZN(new_n8427_));
  NOR2_X1    g08350(.A1(new_n8427_), .A2(new_n8048_), .ZN(new_n8428_));
  OAI22_X1   g08351(.A1(new_n8428_), .A2(new_n8057_), .B1(new_n8067_), .B2(new_n8069_), .ZN(new_n8429_));
  XOR2_X1    g08352(.A1(new_n8062_), .A2(new_n8065_), .Z(new_n8430_));
  INV_X1     g08353(.I(new_n8430_), .ZN(new_n8431_));
  NAND2_X1   g08354(.A1(new_n8058_), .A2(new_n8431_), .ZN(new_n8432_));
  NAND2_X1   g08355(.A1(new_n8432_), .A2(new_n8429_), .ZN(new_n8433_));
  OAI21_X1   g08356(.A1(new_n8057_), .A2(new_n8427_), .B(new_n8049_), .ZN(new_n8434_));
  NOR2_X1    g08357(.A1(new_n8052_), .A2(new_n8426_), .ZN(new_n8435_));
  NOR2_X1    g08358(.A1(new_n8425_), .A2(new_n8055_), .ZN(new_n8436_));
  OAI21_X1   g08359(.A1(new_n8435_), .A2(new_n8436_), .B(new_n8048_), .ZN(new_n8437_));
  OAI22_X1   g08360(.A1(new_n4285_), .A2(new_n2495_), .B1(new_n6621_), .B2(new_n7837_), .ZN(new_n8438_));
  NAND2_X1   g08361(.A1(new_n8438_), .A2(new_n498_), .ZN(new_n8439_));
  NAND2_X1   g08362(.A1(new_n8439_), .A2(new_n2469_), .ZN(new_n8440_));
  XOR2_X1    g08363(.A1(new_n5023_), .A2(new_n8440_), .Z(new_n8441_));
  NAND3_X1   g08364(.A1(new_n8434_), .A2(new_n8437_), .A3(new_n8441_), .ZN(new_n8442_));
  INV_X1     g08365(.I(new_n8442_), .ZN(new_n8443_));
  AOI21_X1   g08366(.A1(new_n8434_), .A2(new_n8437_), .B(new_n8441_), .ZN(new_n8444_));
  NOR2_X1    g08367(.A1(new_n8443_), .A2(new_n8444_), .ZN(new_n8445_));
  INV_X1     g08368(.I(new_n8445_), .ZN(new_n8446_));
  INV_X1     g08369(.I(new_n7528_), .ZN(new_n8447_));
  XOR2_X1    g08370(.A1(new_n8018_), .A2(new_n7521_), .Z(new_n8448_));
  XOR2_X1    g08371(.A1(new_n8448_), .A2(new_n8021_), .Z(new_n8449_));
  XOR2_X1    g08372(.A1(new_n8449_), .A2(new_n8447_), .Z(new_n8450_));
  XNOR2_X1   g08373(.A1(new_n7989_), .A2(new_n7526_), .ZN(new_n8451_));
  INV_X1     g08374(.I(new_n8006_), .ZN(new_n8452_));
  OAI21_X1   g08375(.A1(new_n8452_), .A2(new_n7990_), .B(new_n8005_), .ZN(new_n8453_));
  OAI21_X1   g08376(.A1(new_n8451_), .A2(new_n8005_), .B(new_n8453_), .ZN(new_n8454_));
  OAI22_X1   g08377(.A1(new_n5684_), .A2(new_n2495_), .B1(new_n6556_), .B2(new_n7837_), .ZN(new_n8455_));
  AOI21_X1   g08378(.A1(new_n8455_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8456_));
  NAND2_X1   g08379(.A1(new_n6102_), .A2(new_n8456_), .ZN(new_n8457_));
  INV_X1     g08380(.I(new_n8456_), .ZN(new_n8458_));
  NAND2_X1   g08381(.A1(new_n5693_), .A2(new_n8458_), .ZN(new_n8459_));
  NAND2_X1   g08382(.A1(new_n8457_), .A2(new_n8459_), .ZN(new_n8460_));
  INV_X1     g08383(.I(new_n8460_), .ZN(new_n8461_));
  XOR2_X1    g08384(.A1(new_n8016_), .A2(new_n8010_), .Z(new_n8462_));
  NAND2_X1   g08385(.A1(new_n8014_), .A2(new_n8017_), .ZN(new_n8463_));
  NAND2_X1   g08386(.A1(new_n8463_), .A2(new_n8007_), .ZN(new_n8464_));
  OAI21_X1   g08387(.A1(new_n8007_), .A2(new_n8462_), .B(new_n8464_), .ZN(new_n8465_));
  OAI22_X1   g08388(.A1(new_n4150_), .A2(new_n2495_), .B1(new_n6567_), .B2(new_n7837_), .ZN(new_n8466_));
  AOI21_X1   g08389(.A1(new_n8466_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8467_));
  XOR2_X1    g08390(.A1(new_n5707_), .A2(new_n8467_), .Z(new_n8468_));
  NOR2_X1    g08391(.A1(new_n8465_), .A2(new_n8468_), .ZN(new_n8469_));
  AND2_X2    g08392(.A1(new_n8465_), .A2(new_n8468_), .Z(new_n8470_));
  NOR2_X1    g08393(.A1(new_n8470_), .A2(new_n8469_), .ZN(new_n8471_));
  NOR2_X1    g08394(.A1(new_n8471_), .A2(new_n8461_), .ZN(new_n8472_));
  NOR2_X1    g08395(.A1(new_n8472_), .A2(new_n8454_), .ZN(new_n8473_));
  OAI22_X1   g08396(.A1(new_n6504_), .A2(new_n7837_), .B1(new_n2495_), .B2(new_n4249_), .ZN(new_n8474_));
  NAND2_X1   g08397(.A1(new_n8474_), .A2(new_n498_), .ZN(new_n8475_));
  NAND2_X1   g08398(.A1(new_n8475_), .A2(new_n2469_), .ZN(new_n8476_));
  XOR2_X1    g08399(.A1(new_n8476_), .A2(new_n6245_), .Z(new_n8477_));
  INV_X1     g08400(.I(new_n8477_), .ZN(new_n8478_));
  NOR2_X1    g08401(.A1(new_n8478_), .A2(new_n8001_), .ZN(new_n8479_));
  NAND2_X1   g08402(.A1(new_n5627_), .A2(new_n2495_), .ZN(new_n8480_));
  AOI21_X1   g08403(.A1(new_n2469_), .A2(new_n6061_), .B(new_n4260_), .ZN(new_n8481_));
  OAI22_X1   g08404(.A1(new_n4244_), .A2(new_n7836_), .B1(new_n2718_), .B2(new_n4230_), .ZN(new_n8482_));
  OAI21_X1   g08405(.A1(new_n2495_), .A2(new_n4234_), .B(new_n8482_), .ZN(new_n8483_));
  AOI21_X1   g08406(.A1(new_n8480_), .A2(new_n8481_), .B(new_n8483_), .ZN(new_n8484_));
  XOR2_X1    g08407(.A1(new_n8484_), .A2(\a[8] ), .Z(new_n8485_));
  NOR2_X1    g08408(.A1(new_n4244_), .A2(new_n2718_), .ZN(new_n8486_));
  OAI21_X1   g08409(.A1(new_n4230_), .A2(new_n2495_), .B(new_n498_), .ZN(new_n8487_));
  OAI21_X1   g08410(.A1(new_n8486_), .A2(new_n8487_), .B(new_n2469_), .ZN(new_n8488_));
  XOR2_X1    g08411(.A1(new_n8488_), .A2(new_n5637_), .Z(new_n8489_));
  NOR2_X1    g08412(.A1(new_n4251_), .A2(new_n2583_), .ZN(new_n8490_));
  NOR2_X1    g08413(.A1(new_n8490_), .A2(new_n498_), .ZN(new_n8491_));
  INV_X1     g08414(.I(new_n8491_), .ZN(new_n8492_));
  NOR2_X1    g08415(.A1(new_n8489_), .A2(new_n8492_), .ZN(new_n8493_));
  NAND2_X1   g08416(.A1(new_n8485_), .A2(new_n8493_), .ZN(new_n8494_));
  INV_X1     g08417(.I(new_n8494_), .ZN(new_n8495_));
  INV_X1     g08418(.I(new_n8001_), .ZN(new_n8496_));
  NOR2_X1    g08419(.A1(new_n8477_), .A2(new_n8496_), .ZN(new_n8497_));
  NOR2_X1    g08420(.A1(new_n8495_), .A2(new_n8497_), .ZN(new_n8498_));
  NOR2_X1    g08421(.A1(new_n8498_), .A2(new_n8479_), .ZN(new_n8499_));
  XOR2_X1    g08422(.A1(new_n8000_), .A2(new_n8002_), .Z(new_n8500_));
  OAI22_X1   g08423(.A1(new_n4203_), .A2(new_n2495_), .B1(new_n6529_), .B2(new_n7837_), .ZN(new_n8501_));
  AOI21_X1   g08424(.A1(new_n8501_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8502_));
  XOR2_X1    g08425(.A1(new_n5660_), .A2(new_n8502_), .Z(new_n8503_));
  NOR2_X1    g08426(.A1(new_n8503_), .A2(new_n8500_), .ZN(new_n8504_));
  NAND2_X1   g08427(.A1(new_n8503_), .A2(new_n8500_), .ZN(new_n8505_));
  OAI21_X1   g08428(.A1(new_n8499_), .A2(new_n8504_), .B(new_n8505_), .ZN(new_n8506_));
  INV_X1     g08429(.I(new_n8506_), .ZN(new_n8507_));
  XNOR2_X1   g08430(.A1(new_n7996_), .A2(new_n8004_), .ZN(new_n8508_));
  AOI22_X1   g08431(.A1(new_n4258_), .A2(new_n2469_), .B1(new_n6541_), .B2(new_n7838_), .ZN(new_n8509_));
  OAI21_X1   g08432(.A1(new_n8509_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8510_));
  XOR2_X1    g08433(.A1(new_n6540_), .A2(new_n8510_), .Z(new_n8511_));
  NOR2_X1    g08434(.A1(new_n8511_), .A2(new_n8508_), .ZN(new_n8512_));
  NAND2_X1   g08435(.A1(new_n8511_), .A2(new_n8508_), .ZN(new_n8513_));
  OAI21_X1   g08436(.A1(new_n8507_), .A2(new_n8512_), .B(new_n8513_), .ZN(new_n8514_));
  NAND2_X1   g08437(.A1(new_n8471_), .A2(new_n8461_), .ZN(new_n8515_));
  NAND2_X1   g08438(.A1(new_n8515_), .A2(new_n8514_), .ZN(new_n8516_));
  OR2_X2     g08439(.A1(new_n8473_), .A2(new_n8516_), .Z(new_n8517_));
  NOR2_X1    g08440(.A1(new_n8517_), .A2(new_n8450_), .ZN(new_n8518_));
  AOI22_X1   g08441(.A1(new_n6582_), .A2(new_n7838_), .B1(new_n4274_), .B2(new_n2469_), .ZN(new_n8519_));
  OAI21_X1   g08442(.A1(new_n8519_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8520_));
  XNOR2_X1   g08443(.A1(new_n5722_), .A2(new_n8520_), .ZN(new_n8521_));
  NAND2_X1   g08444(.A1(new_n8521_), .A2(new_n8470_), .ZN(new_n8522_));
  AOI21_X1   g08445(.A1(new_n8517_), .A2(new_n8450_), .B(new_n8522_), .ZN(new_n8523_));
  NOR2_X1    g08446(.A1(new_n8523_), .A2(new_n8518_), .ZN(new_n8524_));
  XOR2_X1    g08447(.A1(new_n8034_), .A2(new_n8031_), .Z(new_n8525_));
  AOI21_X1   g08448(.A1(new_n8037_), .A2(new_n8035_), .B(new_n8026_), .ZN(new_n8526_));
  AOI21_X1   g08449(.A1(new_n8026_), .A2(new_n8525_), .B(new_n8526_), .ZN(new_n8527_));
  OAI22_X1   g08450(.A1(new_n4142_), .A2(new_n2495_), .B1(new_n4277_), .B2(new_n7837_), .ZN(new_n8528_));
  AOI21_X1   g08451(.A1(new_n8528_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8529_));
  XOR2_X1    g08452(.A1(new_n6134_), .A2(new_n8529_), .Z(new_n8530_));
  INV_X1     g08453(.I(new_n8530_), .ZN(new_n8531_));
  NOR2_X1    g08454(.A1(new_n8527_), .A2(new_n8531_), .ZN(new_n8532_));
  NAND2_X1   g08455(.A1(new_n8527_), .A2(new_n8531_), .ZN(new_n8533_));
  OAI21_X1   g08456(.A1(new_n8524_), .A2(new_n8532_), .B(new_n8533_), .ZN(new_n8534_));
  XOR2_X1    g08457(.A1(new_n8044_), .A2(new_n8041_), .Z(new_n8535_));
  NAND2_X1   g08458(.A1(new_n8038_), .A2(new_n8535_), .ZN(new_n8536_));
  NOR2_X1    g08459(.A1(new_n8047_), .A2(new_n8045_), .ZN(new_n8537_));
  OAI21_X1   g08460(.A1(new_n8038_), .A2(new_n8537_), .B(new_n8536_), .ZN(new_n8538_));
  NAND2_X1   g08461(.A1(new_n6609_), .A2(new_n7838_), .ZN(new_n8539_));
  OAI21_X1   g08462(.A1(new_n4135_), .A2(new_n2495_), .B(new_n8539_), .ZN(new_n8540_));
  AOI21_X1   g08463(.A1(new_n8540_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8541_));
  XNOR2_X1   g08464(.A1(new_n5624_), .A2(new_n8541_), .ZN(new_n8542_));
  NAND2_X1   g08465(.A1(new_n8538_), .A2(new_n8542_), .ZN(new_n8543_));
  NOR2_X1    g08466(.A1(new_n8538_), .A2(new_n8542_), .ZN(new_n8544_));
  AOI21_X1   g08467(.A1(new_n8534_), .A2(new_n8543_), .B(new_n8544_), .ZN(new_n8545_));
  INV_X1     g08468(.I(new_n8545_), .ZN(new_n8546_));
  NOR2_X1    g08469(.A1(new_n8446_), .A2(new_n8546_), .ZN(new_n8547_));
  NAND2_X1   g08470(.A1(new_n8547_), .A2(new_n8433_), .ZN(new_n8548_));
  AOI22_X1   g08471(.A1(new_n6961_), .A2(new_n7838_), .B1(new_n4297_), .B2(new_n2469_), .ZN(new_n8549_));
  OAI21_X1   g08472(.A1(new_n8549_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8550_));
  XOR2_X1    g08473(.A1(new_n5753_), .A2(new_n8550_), .Z(new_n8551_));
  NOR2_X1    g08474(.A1(new_n8442_), .A2(new_n8551_), .ZN(new_n8552_));
  OAI21_X1   g08475(.A1(new_n8547_), .A2(new_n8433_), .B(new_n8552_), .ZN(new_n8553_));
  NOR2_X1    g08476(.A1(new_n8068_), .A2(new_n8069_), .ZN(new_n8554_));
  XOR2_X1    g08477(.A1(new_n8075_), .A2(new_n8079_), .Z(new_n8555_));
  NOR2_X1    g08478(.A1(new_n8554_), .A2(new_n8555_), .ZN(new_n8556_));
  INV_X1     g08479(.I(new_n8556_), .ZN(new_n8557_));
  NOR2_X1    g08480(.A1(new_n8080_), .A2(new_n8075_), .ZN(new_n8558_));
  OAI21_X1   g08481(.A1(new_n8558_), .A2(new_n8083_), .B(new_n8554_), .ZN(new_n8559_));
  OAI22_X1   g08482(.A1(new_n4131_), .A2(new_n2495_), .B1(new_n4301_), .B2(new_n7837_), .ZN(new_n8560_));
  AOI21_X1   g08483(.A1(new_n8560_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8561_));
  XNOR2_X1   g08484(.A1(new_n5599_), .A2(new_n8561_), .ZN(new_n8562_));
  INV_X1     g08485(.I(new_n8562_), .ZN(new_n8563_));
  AOI21_X1   g08486(.A1(new_n8557_), .A2(new_n8559_), .B(new_n8563_), .ZN(new_n8564_));
  AOI21_X1   g08487(.A1(new_n8553_), .A2(new_n8548_), .B(new_n8564_), .ZN(new_n8565_));
  INV_X1     g08488(.I(new_n8559_), .ZN(new_n8566_));
  NOR3_X1    g08489(.A1(new_n8566_), .A2(new_n8556_), .A3(new_n8562_), .ZN(new_n8567_));
  NOR2_X1    g08490(.A1(new_n8565_), .A2(new_n8567_), .ZN(new_n8568_));
  AOI22_X1   g08491(.A1(new_n6980_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n5041_), .ZN(new_n8569_));
  OAI21_X1   g08492(.A1(new_n8569_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8570_));
  XOR2_X1    g08493(.A1(new_n5049_), .A2(new_n8570_), .Z(new_n8571_));
  NOR2_X1    g08494(.A1(new_n8568_), .A2(new_n8571_), .ZN(new_n8572_));
  NAND2_X1   g08495(.A1(new_n8081_), .A2(new_n8084_), .ZN(new_n8573_));
  XOR2_X1    g08496(.A1(new_n8573_), .A2(new_n8095_), .Z(new_n8574_));
  AOI21_X1   g08497(.A1(new_n8568_), .A2(new_n8571_), .B(new_n8574_), .ZN(new_n8575_));
  INV_X1     g08498(.I(new_n8573_), .ZN(new_n8576_));
  INV_X1     g08499(.I(new_n8100_), .ZN(new_n8577_));
  NAND2_X1   g08500(.A1(new_n7984_), .A2(new_n8577_), .ZN(new_n8578_));
  AOI21_X1   g08501(.A1(new_n8576_), .A2(new_n8095_), .B(new_n8578_), .ZN(new_n8579_));
  AOI21_X1   g08502(.A1(new_n7984_), .A2(new_n8577_), .B(new_n8096_), .ZN(new_n8580_));
  OAI21_X1   g08503(.A1(new_n8579_), .A2(new_n8580_), .B(new_n8092_), .ZN(new_n8581_));
  OR3_X2     g08504(.A1(new_n8579_), .A2(new_n8092_), .A3(new_n8580_), .Z(new_n8582_));
  AOI22_X1   g08505(.A1(new_n6993_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4124_), .ZN(new_n8583_));
  OAI21_X1   g08506(.A1(new_n8583_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8584_));
  XOR2_X1    g08507(.A1(new_n5067_), .A2(new_n8584_), .Z(new_n8585_));
  INV_X1     g08508(.I(new_n8585_), .ZN(new_n8586_));
  NAND3_X1   g08509(.A1(new_n8582_), .A2(new_n8581_), .A3(new_n8586_), .ZN(new_n8587_));
  INV_X1     g08510(.I(new_n8587_), .ZN(new_n8588_));
  AOI21_X1   g08511(.A1(new_n8582_), .A2(new_n8581_), .B(new_n8586_), .ZN(new_n8589_));
  NOR4_X1    g08512(.A1(new_n8588_), .A2(new_n8575_), .A3(new_n8572_), .A4(new_n8589_), .ZN(new_n8590_));
  NAND2_X1   g08513(.A1(new_n8590_), .A2(new_n8424_), .ZN(new_n8591_));
  INV_X1     g08514(.I(new_n8589_), .ZN(new_n8592_));
  OAI22_X1   g08515(.A1(new_n4112_), .A2(new_n2495_), .B1(new_n6682_), .B2(new_n7837_), .ZN(new_n8593_));
  AOI21_X1   g08516(.A1(new_n8593_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8594_));
  XOR2_X1    g08517(.A1(new_n5096_), .A2(new_n8594_), .Z(new_n8595_));
  NOR2_X1    g08518(.A1(new_n8592_), .A2(new_n8595_), .ZN(new_n8596_));
  OAI21_X1   g08519(.A1(new_n8590_), .A2(new_n8424_), .B(new_n8596_), .ZN(new_n8597_));
  INV_X1     g08520(.I(new_n8116_), .ZN(new_n8598_));
  INV_X1     g08521(.I(new_n8123_), .ZN(new_n8599_));
  AOI21_X1   g08522(.A1(new_n8122_), .A2(new_n8599_), .B(new_n8598_), .ZN(new_n8600_));
  XOR2_X1    g08523(.A1(new_n8117_), .A2(new_n8121_), .Z(new_n8601_));
  NOR2_X1    g08524(.A1(new_n8116_), .A2(new_n8601_), .ZN(new_n8602_));
  NOR2_X1    g08525(.A1(new_n8600_), .A2(new_n8602_), .ZN(new_n8603_));
  AOI22_X1   g08526(.A1(new_n7015_), .A2(new_n7838_), .B1(new_n4105_), .B2(new_n2469_), .ZN(new_n8604_));
  OAI21_X1   g08527(.A1(new_n8604_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8605_));
  XOR2_X1    g08528(.A1(new_n5121_), .A2(new_n8605_), .Z(new_n8606_));
  AOI22_X1   g08529(.A1(new_n8597_), .A2(new_n8591_), .B1(new_n8603_), .B2(new_n8606_), .ZN(new_n8607_));
  NOR2_X1    g08530(.A1(new_n8603_), .A2(new_n8606_), .ZN(new_n8608_));
  AOI22_X1   g08531(.A1(new_n7021_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4100_), .ZN(new_n8609_));
  OAI21_X1   g08532(.A1(new_n8609_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8610_));
  XOR2_X1    g08533(.A1(new_n5080_), .A2(new_n8610_), .Z(new_n8611_));
  XNOR2_X1   g08534(.A1(new_n8140_), .A2(new_n8611_), .ZN(new_n8612_));
  NOR2_X1    g08535(.A1(new_n8612_), .A2(new_n8124_), .ZN(new_n8613_));
  INV_X1     g08536(.I(new_n8124_), .ZN(new_n8614_));
  XOR2_X1    g08537(.A1(new_n8140_), .A2(new_n8611_), .Z(new_n8615_));
  NOR2_X1    g08538(.A1(new_n8615_), .A2(new_n8614_), .ZN(new_n8616_));
  NOR4_X1    g08539(.A1(new_n8607_), .A2(new_n8608_), .A3(new_n8613_), .A4(new_n8616_), .ZN(new_n8617_));
  NAND2_X1   g08540(.A1(new_n8617_), .A2(new_n8419_), .ZN(new_n8618_));
  XNOR2_X1   g08541(.A1(new_n8124_), .A2(new_n8140_), .ZN(new_n8619_));
  NAND2_X1   g08542(.A1(new_n8619_), .A2(new_n8611_), .ZN(new_n8620_));
  OAI22_X1   g08543(.A1(new_n4090_), .A2(new_n2495_), .B1(new_n4320_), .B2(new_n7837_), .ZN(new_n8621_));
  AOI21_X1   g08544(.A1(new_n8621_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8622_));
  XOR2_X1    g08545(.A1(new_n5196_), .A2(new_n8622_), .Z(new_n8623_));
  NOR2_X1    g08546(.A1(new_n8620_), .A2(new_n8623_), .ZN(new_n8624_));
  OAI21_X1   g08547(.A1(new_n8617_), .A2(new_n8419_), .B(new_n8624_), .ZN(new_n8625_));
  NAND2_X1   g08548(.A1(new_n8152_), .A2(new_n8150_), .ZN(new_n8626_));
  NAND2_X1   g08549(.A1(new_n8626_), .A2(new_n8155_), .ZN(new_n8627_));
  OR2_X2     g08550(.A1(new_n8626_), .A2(new_n8155_), .Z(new_n8628_));
  AOI21_X1   g08551(.A1(new_n8628_), .A2(new_n8627_), .B(new_n8221_), .ZN(new_n8629_));
  INV_X1     g08552(.I(new_n8629_), .ZN(new_n8630_));
  AOI21_X1   g08553(.A1(new_n8156_), .A2(new_n8159_), .B(new_n8222_), .ZN(new_n8631_));
  INV_X1     g08554(.I(new_n8631_), .ZN(new_n8632_));
  AOI22_X1   g08555(.A1(new_n6419_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4328_), .ZN(new_n8633_));
  OAI21_X1   g08556(.A1(new_n8633_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8634_));
  XOR2_X1    g08557(.A1(new_n5139_), .A2(new_n8634_), .Z(new_n8635_));
  NAND3_X1   g08558(.A1(new_n8630_), .A2(new_n8632_), .A3(new_n8635_), .ZN(new_n8636_));
  INV_X1     g08559(.I(new_n8635_), .ZN(new_n8637_));
  OAI21_X1   g08560(.A1(new_n8629_), .A2(new_n8631_), .B(new_n8637_), .ZN(new_n8638_));
  NOR2_X1    g08561(.A1(new_n8160_), .A2(new_n8225_), .ZN(new_n8639_));
  NOR2_X1    g08562(.A1(new_n8223_), .A2(new_n8169_), .ZN(new_n8640_));
  AOI22_X1   g08563(.A1(new_n4333_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4082_), .ZN(new_n8641_));
  OAI21_X1   g08564(.A1(new_n8641_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8642_));
  XNOR2_X1   g08565(.A1(new_n5162_), .A2(new_n8642_), .ZN(new_n8643_));
  NOR3_X1    g08566(.A1(new_n8639_), .A2(new_n8640_), .A3(new_n8643_), .ZN(new_n8644_));
  OAI21_X1   g08567(.A1(new_n8639_), .A2(new_n8640_), .B(new_n8643_), .ZN(new_n8645_));
  INV_X1     g08568(.I(new_n8645_), .ZN(new_n8646_));
  AOI22_X1   g08569(.A1(new_n8636_), .A2(new_n8638_), .B1(new_n8625_), .B2(new_n8618_), .ZN(new_n8648_));
  NAND2_X1   g08570(.A1(new_n8411_), .A2(new_n8648_), .ZN(new_n8649_));
  OAI22_X1   g08571(.A1(new_n4070_), .A2(new_n2495_), .B1(new_n5917_), .B2(new_n7837_), .ZN(new_n8650_));
  AOI21_X1   g08572(.A1(new_n8650_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8651_));
  AND2_X2    g08573(.A1(new_n4927_), .A2(new_n8651_), .Z(new_n8652_));
  NOR2_X1    g08574(.A1(new_n4927_), .A2(new_n8651_), .ZN(new_n8653_));
  NOR2_X1    g08575(.A1(new_n8652_), .A2(new_n8653_), .ZN(new_n8654_));
  NOR2_X1    g08576(.A1(new_n8645_), .A2(new_n8654_), .ZN(new_n8655_));
  OAI21_X1   g08577(.A1(new_n8411_), .A2(new_n8648_), .B(new_n8655_), .ZN(new_n8656_));
  NAND2_X1   g08578(.A1(new_n8656_), .A2(new_n8649_), .ZN(new_n8657_));
  INV_X1     g08579(.I(new_n8657_), .ZN(new_n8658_));
  NOR3_X1    g08580(.A1(new_n8214_), .A2(new_n8217_), .A3(new_n8230_), .ZN(new_n8659_));
  NOR3_X1    g08581(.A1(new_n8659_), .A2(new_n8228_), .A3(new_n8391_), .ZN(new_n8660_));
  NAND3_X1   g08582(.A1(new_n8215_), .A2(new_n8216_), .A3(new_n8212_), .ZN(new_n8661_));
  OAI21_X1   g08583(.A1(new_n8209_), .A2(new_n8206_), .B(new_n8213_), .ZN(new_n8662_));
  NAND3_X1   g08584(.A1(new_n8662_), .A2(new_n8661_), .A3(new_n8204_), .ZN(new_n8663_));
  AOI21_X1   g08585(.A1(new_n8663_), .A2(new_n8389_), .B(new_n8181_), .ZN(new_n8664_));
  AOI22_X1   g08586(.A1(new_n6428_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4054_), .ZN(new_n8665_));
  OAI21_X1   g08587(.A1(new_n8665_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8666_));
  XOR2_X1    g08588(.A1(new_n4652_), .A2(new_n8666_), .Z(new_n8667_));
  NOR3_X1    g08589(.A1(new_n8664_), .A2(new_n8660_), .A3(new_n8667_), .ZN(new_n8668_));
  NAND3_X1   g08590(.A1(new_n8663_), .A2(new_n8181_), .A3(new_n8389_), .ZN(new_n8669_));
  OAI21_X1   g08591(.A1(new_n8659_), .A2(new_n8391_), .B(new_n8228_), .ZN(new_n8670_));
  INV_X1     g08592(.I(new_n8667_), .ZN(new_n8671_));
  AOI21_X1   g08593(.A1(new_n8670_), .A2(new_n8669_), .B(new_n8671_), .ZN(new_n8672_));
  OAI21_X1   g08594(.A1(new_n8668_), .A2(new_n8672_), .B(new_n8399_), .ZN(new_n8673_));
  AOI21_X1   g08595(.A1(new_n8658_), .A2(new_n8673_), .B(new_n8403_), .ZN(new_n8674_));
  NAND2_X1   g08596(.A1(new_n8388_), .A2(new_n8674_), .ZN(new_n8675_));
  OAI22_X1   g08597(.A1(new_n4042_), .A2(new_n2495_), .B1(new_n4342_), .B2(new_n7837_), .ZN(new_n8676_));
  AOI21_X1   g08598(.A1(new_n8676_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8677_));
  XOR2_X1    g08599(.A1(new_n4864_), .A2(new_n8677_), .Z(new_n8678_));
  AND2_X2    g08600(.A1(new_n8678_), .A2(new_n8672_), .Z(new_n8679_));
  OAI21_X1   g08601(.A1(new_n8388_), .A2(new_n8674_), .B(new_n8679_), .ZN(new_n8680_));
  AOI21_X1   g08602(.A1(new_n7941_), .A2(new_n7938_), .B(new_n7946_), .ZN(new_n8681_));
  NOR2_X1    g08603(.A1(new_n8681_), .A2(new_n8366_), .ZN(new_n8682_));
  NAND2_X1   g08604(.A1(new_n8240_), .A2(new_n8682_), .ZN(new_n8683_));
  NAND2_X1   g08605(.A1(new_n8365_), .A2(new_n7952_), .ZN(new_n8684_));
  AOI22_X1   g08606(.A1(new_n4347_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4036_), .ZN(new_n8685_));
  OAI21_X1   g08607(.A1(new_n8685_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8686_));
  XNOR2_X1   g08608(.A1(new_n4672_), .A2(new_n8686_), .ZN(new_n8687_));
  NAND3_X1   g08609(.A1(new_n8683_), .A2(new_n8684_), .A3(new_n8687_), .ZN(new_n8688_));
  NOR2_X1    g08610(.A1(new_n8365_), .A2(new_n7952_), .ZN(new_n8689_));
  NOR2_X1    g08611(.A1(new_n8240_), .A2(new_n8682_), .ZN(new_n8690_));
  XOR2_X1    g08612(.A1(new_n4672_), .A2(new_n8686_), .Z(new_n8691_));
  OAI21_X1   g08613(.A1(new_n8690_), .A2(new_n8689_), .B(new_n8691_), .ZN(new_n8692_));
  NOR3_X1    g08614(.A1(new_n8257_), .A2(new_n8367_), .A3(new_n8366_), .ZN(new_n8693_));
  NOR3_X1    g08615(.A1(new_n8693_), .A2(new_n7952_), .A3(new_n8365_), .ZN(new_n8694_));
  NAND3_X1   g08616(.A1(new_n8253_), .A2(new_n8249_), .A3(new_n7947_), .ZN(new_n8695_));
  AOI21_X1   g08617(.A1(new_n8695_), .A2(new_n8240_), .B(new_n8682_), .ZN(new_n8696_));
  AOI22_X1   g08618(.A1(new_n5935_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4029_), .ZN(new_n8697_));
  OAI21_X1   g08619(.A1(new_n8697_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8698_));
  XOR2_X1    g08620(.A1(new_n4687_), .A2(new_n8698_), .Z(new_n8699_));
  NOR3_X1    g08621(.A1(new_n8694_), .A2(new_n8696_), .A3(new_n8699_), .ZN(new_n8700_));
  NAND3_X1   g08622(.A1(new_n8695_), .A2(new_n8240_), .A3(new_n8682_), .ZN(new_n8701_));
  OAI21_X1   g08623(.A1(new_n8693_), .A2(new_n8365_), .B(new_n7952_), .ZN(new_n8702_));
  INV_X1     g08624(.I(new_n8698_), .ZN(new_n8703_));
  XOR2_X1    g08625(.A1(new_n4687_), .A2(new_n8703_), .Z(new_n8704_));
  AOI21_X1   g08626(.A1(new_n8702_), .A2(new_n8701_), .B(new_n8704_), .ZN(new_n8705_));
  AOI22_X1   g08627(.A1(new_n8680_), .A2(new_n8675_), .B1(new_n8692_), .B2(new_n8688_), .ZN(new_n8707_));
  INV_X1     g08628(.I(new_n8707_), .ZN(new_n8708_));
  NOR2_X1    g08629(.A1(new_n8376_), .A2(new_n8708_), .ZN(new_n8709_));
  NOR2_X1    g08630(.A1(new_n4028_), .A2(new_n7836_), .ZN(new_n8710_));
  NOR2_X1    g08631(.A1(new_n4035_), .A2(new_n2718_), .ZN(new_n8711_));
  OAI22_X1   g08632(.A1(new_n4017_), .A2(new_n2495_), .B1(new_n8710_), .B2(new_n8711_), .ZN(new_n8712_));
  AOI21_X1   g08633(.A1(new_n8712_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8713_));
  XOR2_X1    g08634(.A1(new_n4705_), .A2(new_n8713_), .Z(new_n8714_));
  NAND2_X1   g08635(.A1(new_n8714_), .A2(new_n8705_), .ZN(new_n8715_));
  AOI21_X1   g08636(.A1(new_n8376_), .A2(new_n8708_), .B(new_n8715_), .ZN(new_n8716_));
  NOR2_X1    g08637(.A1(new_n7920_), .A2(new_n8267_), .ZN(new_n8717_));
  NOR2_X1    g08638(.A1(new_n8350_), .A2(new_n8349_), .ZN(new_n8718_));
  AOI22_X1   g08639(.A1(new_n5859_), .A2(new_n7838_), .B1(new_n4375_), .B2(new_n2469_), .ZN(new_n8719_));
  OAI21_X1   g08640(.A1(new_n8719_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8720_));
  XOR2_X1    g08641(.A1(new_n4730_), .A2(new_n8720_), .Z(new_n8721_));
  NOR3_X1    g08642(.A1(new_n8718_), .A2(new_n8717_), .A3(new_n8721_), .ZN(new_n8722_));
  NAND2_X1   g08643(.A1(new_n8350_), .A2(new_n8349_), .ZN(new_n8723_));
  NAND2_X1   g08644(.A1(new_n7920_), .A2(new_n8267_), .ZN(new_n8724_));
  XNOR2_X1   g08645(.A1(new_n4730_), .A2(new_n8720_), .ZN(new_n8725_));
  AOI21_X1   g08646(.A1(new_n8723_), .A2(new_n8724_), .B(new_n8725_), .ZN(new_n8726_));
  NOR3_X1    g08647(.A1(new_n8280_), .A2(new_n8283_), .A3(new_n7915_), .ZN(new_n8727_));
  NOR3_X1    g08648(.A1(new_n7920_), .A2(new_n8727_), .A3(new_n8267_), .ZN(new_n8728_));
  NAND3_X1   g08649(.A1(new_n8352_), .A2(new_n8288_), .A3(new_n8351_), .ZN(new_n8729_));
  AOI21_X1   g08650(.A1(new_n8350_), .A2(new_n8729_), .B(new_n8349_), .ZN(new_n8730_));
  AOI22_X1   g08651(.A1(new_n4445_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4399_), .ZN(new_n8731_));
  OAI21_X1   g08652(.A1(new_n8731_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8732_));
  XOR2_X1    g08653(.A1(new_n4403_), .A2(new_n8732_), .Z(new_n8733_));
  NOR3_X1    g08654(.A1(new_n8728_), .A2(new_n8730_), .A3(new_n8733_), .ZN(new_n8734_));
  NAND3_X1   g08655(.A1(new_n8350_), .A2(new_n8729_), .A3(new_n8349_), .ZN(new_n8735_));
  OAI21_X1   g08656(.A1(new_n8727_), .A2(new_n8267_), .B(new_n7920_), .ZN(new_n8736_));
  INV_X1     g08657(.I(new_n8733_), .ZN(new_n8737_));
  AOI21_X1   g08658(.A1(new_n8736_), .A2(new_n8735_), .B(new_n8737_), .ZN(new_n8738_));
  OAI22_X1   g08659(.A1(new_n8726_), .A2(new_n8722_), .B1(new_n8709_), .B2(new_n8716_), .ZN(new_n8740_));
  NOR2_X1    g08660(.A1(new_n8359_), .A2(new_n8740_), .ZN(new_n8741_));
  INV_X1     g08661(.I(new_n8741_), .ZN(new_n8742_));
  NAND2_X1   g08662(.A1(new_n8359_), .A2(new_n8740_), .ZN(new_n8743_));
  NOR2_X1    g08663(.A1(new_n4397_), .A2(new_n7836_), .ZN(new_n8744_));
  NOR2_X1    g08664(.A1(new_n4374_), .A2(new_n2718_), .ZN(new_n8745_));
  OAI22_X1   g08665(.A1(new_n4437_), .A2(new_n2495_), .B1(new_n8744_), .B2(new_n8745_), .ZN(new_n8746_));
  AOI21_X1   g08666(.A1(new_n8746_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8747_));
  XNOR2_X1   g08667(.A1(new_n4541_), .A2(new_n8747_), .ZN(new_n8748_));
  NAND3_X1   g08668(.A1(new_n8743_), .A2(new_n8738_), .A3(new_n8748_), .ZN(new_n8749_));
  NAND2_X1   g08669(.A1(new_n8749_), .A2(new_n8742_), .ZN(new_n8750_));
  NAND2_X1   g08670(.A1(new_n7893_), .A2(new_n8298_), .ZN(new_n8751_));
  INV_X1     g08671(.I(new_n8751_), .ZN(new_n8752_));
  NOR2_X1    g08672(.A1(new_n7893_), .A2(new_n8298_), .ZN(new_n8753_));
  AOI22_X1   g08673(.A1(new_n4448_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4469_), .ZN(new_n8754_));
  OAI21_X1   g08674(.A1(new_n8754_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8755_));
  XNOR2_X1   g08675(.A1(new_n4477_), .A2(new_n8755_), .ZN(new_n8756_));
  OAI21_X1   g08676(.A1(new_n8752_), .A2(new_n8753_), .B(new_n8756_), .ZN(new_n8757_));
  NAND2_X1   g08677(.A1(new_n8757_), .A2(new_n8750_), .ZN(new_n8758_));
  NOR3_X1    g08678(.A1(new_n8752_), .A2(new_n8753_), .A3(new_n8756_), .ZN(new_n8759_));
  INV_X1     g08679(.I(new_n8759_), .ZN(new_n8760_));
  NAND2_X1   g08680(.A1(new_n8758_), .A2(new_n8760_), .ZN(new_n8761_));
  INV_X1     g08681(.I(new_n7889_), .ZN(new_n8762_));
  NAND3_X1   g08682(.A1(new_n8315_), .A2(new_n8307_), .A3(new_n8762_), .ZN(new_n8763_));
  NAND3_X1   g08683(.A1(new_n8763_), .A2(new_n7893_), .A3(new_n8298_), .ZN(new_n8764_));
  INV_X1     g08684(.I(new_n8764_), .ZN(new_n8765_));
  AOI21_X1   g08685(.A1(new_n8763_), .A2(new_n8298_), .B(new_n7893_), .ZN(new_n8766_));
  AOI22_X1   g08686(.A1(new_n4473_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n4555_), .ZN(new_n8767_));
  OAI21_X1   g08687(.A1(new_n8767_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n8768_));
  XNOR2_X1   g08688(.A1(new_n4584_), .A2(new_n8768_), .ZN(new_n8769_));
  OAI21_X1   g08689(.A1(new_n8765_), .A2(new_n8766_), .B(new_n8769_), .ZN(new_n8770_));
  NOR3_X1    g08690(.A1(new_n8765_), .A2(new_n8766_), .A3(new_n8769_), .ZN(new_n8771_));
  AOI21_X1   g08691(.A1(new_n8761_), .A2(new_n8770_), .B(new_n8771_), .ZN(new_n8772_));
  INV_X1     g08692(.I(new_n7893_), .ZN(new_n8773_));
  AOI21_X1   g08693(.A1(new_n8303_), .A2(new_n8299_), .B(new_n8306_), .ZN(new_n8774_));
  NOR2_X1    g08694(.A1(new_n8321_), .A2(new_n8774_), .ZN(new_n8775_));
  OAI21_X1   g08695(.A1(new_n8775_), .A2(new_n8762_), .B(new_n8297_), .ZN(new_n8776_));
  OAI21_X1   g08696(.A1(new_n7876_), .A2(new_n7877_), .B(new_n8326_), .ZN(new_n8777_));
  AOI21_X1   g08697(.A1(new_n8776_), .A2(new_n8773_), .B(new_n8777_), .ZN(new_n8778_));
  INV_X1     g08698(.I(new_n7874_), .ZN(new_n8779_));
  AOI21_X1   g08699(.A1(new_n7821_), .A2(new_n7822_), .B(new_n7818_), .ZN(new_n8780_));
  OAI21_X1   g08700(.A1(new_n8779_), .A2(new_n8780_), .B(new_n7805_), .ZN(new_n8781_));
  INV_X1     g08701(.I(new_n7877_), .ZN(new_n8782_));
  AOI21_X1   g08702(.A1(new_n8782_), .A2(new_n8781_), .B(new_n8325_), .ZN(new_n8783_));
  NOR3_X1    g08703(.A1(new_n8783_), .A2(new_n8317_), .A3(new_n7893_), .ZN(new_n8784_));
  OAI21_X1   g08704(.A1(new_n8784_), .A2(new_n8778_), .B(new_n8307_), .ZN(new_n8785_));
  OAI21_X1   g08705(.A1(new_n7893_), .A2(new_n8317_), .B(new_n8783_), .ZN(new_n8786_));
  NAND3_X1   g08706(.A1(new_n8776_), .A2(new_n8777_), .A3(new_n8773_), .ZN(new_n8787_));
  NAND3_X1   g08707(.A1(new_n8786_), .A2(new_n8321_), .A3(new_n8787_), .ZN(new_n8788_));
  OAI22_X1   g08708(.A1(new_n2718_), .A2(new_n4468_), .B1(new_n4501_), .B2(new_n7836_), .ZN(new_n8789_));
  OAI21_X1   g08709(.A1(new_n4516_), .A2(new_n2495_), .B(new_n8789_), .ZN(new_n8790_));
  AOI21_X1   g08710(.A1(new_n8790_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n8791_));
  XOR2_X1    g08711(.A1(new_n4524_), .A2(new_n8791_), .Z(new_n8792_));
  INV_X1     g08712(.I(new_n8792_), .ZN(new_n8793_));
  AOI21_X1   g08713(.A1(new_n8788_), .A2(new_n8785_), .B(new_n8793_), .ZN(new_n8794_));
  AOI21_X1   g08714(.A1(new_n8786_), .A2(new_n8787_), .B(new_n8321_), .ZN(new_n8795_));
  NOR3_X1    g08715(.A1(new_n8784_), .A2(new_n8778_), .A3(new_n8307_), .ZN(new_n8796_));
  NOR3_X1    g08716(.A1(new_n8795_), .A2(new_n8796_), .A3(new_n8792_), .ZN(new_n8797_));
  INV_X1     g08717(.I(new_n8797_), .ZN(new_n8798_));
  OAI21_X1   g08718(.A1(new_n8772_), .A2(new_n8794_), .B(new_n8798_), .ZN(new_n8799_));
  NAND2_X1   g08719(.A1(new_n5033_), .A2(new_n2898_), .ZN(new_n8800_));
  OAI21_X1   g08720(.A1(new_n5031_), .A2(new_n8800_), .B(new_n4564_), .ZN(new_n8801_));
  OAI21_X1   g08721(.A1(new_n8801_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n8802_));
  XOR2_X1    g08722(.A1(new_n5001_), .A2(new_n8802_), .Z(new_n8803_));
  INV_X1     g08723(.I(new_n8803_), .ZN(new_n8804_));
  NOR2_X1    g08724(.A1(new_n8799_), .A2(new_n8804_), .ZN(new_n8805_));
  NAND2_X1   g08725(.A1(new_n8799_), .A2(new_n8804_), .ZN(new_n8806_));
  INV_X1     g08726(.I(new_n8806_), .ZN(new_n8807_));
  OAI22_X1   g08727(.A1(new_n8339_), .A2(new_n8340_), .B1(new_n8805_), .B2(new_n8807_), .ZN(new_n8808_));
  NOR2_X1    g08728(.A1(new_n8339_), .A2(new_n8340_), .ZN(new_n8809_));
  XOR2_X1    g08729(.A1(new_n8799_), .A2(new_n8804_), .Z(new_n8810_));
  NAND2_X1   g08730(.A1(new_n8809_), .A2(new_n8810_), .ZN(new_n8811_));
  AND2_X2    g08731(.A1(new_n8811_), .A2(new_n8808_), .Z(new_n8812_));
  OAI21_X1   g08732(.A1(new_n8728_), .A2(new_n8730_), .B(new_n8733_), .ZN(new_n8813_));
  INV_X1     g08733(.I(new_n8740_), .ZN(new_n8814_));
  AOI21_X1   g08734(.A1(new_n8355_), .A2(new_n8356_), .B(new_n8280_), .ZN(new_n8815_));
  NOR3_X1    g08735(.A1(new_n8347_), .A2(new_n8343_), .A3(new_n8288_), .ZN(new_n8816_));
  OAI21_X1   g08736(.A1(new_n8816_), .A2(new_n8815_), .B(new_n8748_), .ZN(new_n8817_));
  NOR2_X1    g08737(.A1(new_n8817_), .A2(new_n8814_), .ZN(new_n8818_));
  AOI21_X1   g08738(.A1(new_n8358_), .A2(new_n8748_), .B(new_n8740_), .ZN(new_n8819_));
  OAI21_X1   g08739(.A1(new_n8818_), .A2(new_n8819_), .B(new_n8813_), .ZN(new_n8820_));
  NAND3_X1   g08740(.A1(new_n8358_), .A2(new_n8740_), .A3(new_n8748_), .ZN(new_n8821_));
  NAND2_X1   g08741(.A1(new_n8817_), .A2(new_n8814_), .ZN(new_n8822_));
  NAND3_X1   g08742(.A1(new_n8822_), .A2(new_n8821_), .A3(new_n8738_), .ZN(new_n8823_));
  NAND2_X1   g08743(.A1(new_n8820_), .A2(new_n8823_), .ZN(new_n8824_));
  NOR2_X1    g08744(.A1(new_n8716_), .A2(new_n8709_), .ZN(new_n8825_));
  NOR2_X1    g08745(.A1(new_n8726_), .A2(new_n8722_), .ZN(new_n8826_));
  NAND2_X1   g08746(.A1(new_n8826_), .A2(new_n8825_), .ZN(new_n8827_));
  NOR2_X1    g08747(.A1(new_n8826_), .A2(new_n8825_), .ZN(new_n8828_));
  INV_X1     g08748(.I(new_n8828_), .ZN(new_n8829_));
  INV_X1     g08749(.I(new_n5033_), .ZN(new_n8830_));
  NOR2_X1    g08750(.A1(new_n8830_), .A2(new_n3042_), .ZN(new_n8831_));
  INV_X1     g08751(.I(new_n8831_), .ZN(new_n8832_));
  AOI22_X1   g08752(.A1(new_n4448_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4469_), .ZN(new_n8833_));
  OAI21_X1   g08753(.A1(new_n8833_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n8834_));
  XNOR2_X1   g08754(.A1(new_n4477_), .A2(new_n8834_), .ZN(new_n8835_));
  NAND3_X1   g08755(.A1(new_n8829_), .A2(new_n8835_), .A3(new_n8827_), .ZN(new_n8836_));
  INV_X1     g08756(.I(new_n8827_), .ZN(new_n8837_));
  XOR2_X1    g08757(.A1(new_n4477_), .A2(new_n8834_), .Z(new_n8838_));
  OAI21_X1   g08758(.A1(new_n8837_), .A2(new_n8828_), .B(new_n8838_), .ZN(new_n8839_));
  NAND2_X1   g08759(.A1(new_n8839_), .A2(new_n8836_), .ZN(new_n8840_));
  OAI21_X1   g08760(.A1(new_n8373_), .A2(new_n8374_), .B(new_n8249_), .ZN(new_n8841_));
  NAND3_X1   g08761(.A1(new_n8371_), .A2(new_n8363_), .A3(new_n8257_), .ZN(new_n8842_));
  NAND2_X1   g08762(.A1(new_n8841_), .A2(new_n8842_), .ZN(new_n8843_));
  NAND3_X1   g08763(.A1(new_n8843_), .A2(new_n8708_), .A3(new_n8714_), .ZN(new_n8844_));
  INV_X1     g08764(.I(new_n8714_), .ZN(new_n8845_));
  OAI21_X1   g08765(.A1(new_n8376_), .A2(new_n8845_), .B(new_n8707_), .ZN(new_n8846_));
  AOI21_X1   g08766(.A1(new_n8846_), .A2(new_n8844_), .B(new_n8705_), .ZN(new_n8847_));
  OAI21_X1   g08767(.A1(new_n8694_), .A2(new_n8696_), .B(new_n8699_), .ZN(new_n8848_));
  NOR3_X1    g08768(.A1(new_n8376_), .A2(new_n8845_), .A3(new_n8707_), .ZN(new_n8849_));
  AOI21_X1   g08769(.A1(new_n8843_), .A2(new_n8714_), .B(new_n8708_), .ZN(new_n8850_));
  NOR3_X1    g08770(.A1(new_n8849_), .A2(new_n8850_), .A3(new_n8848_), .ZN(new_n8851_));
  NOR2_X1    g08771(.A1(new_n8851_), .A2(new_n8847_), .ZN(new_n8852_));
  NAND3_X1   g08772(.A1(new_n8400_), .A2(new_n8401_), .A3(new_n8397_), .ZN(new_n8853_));
  OAI21_X1   g08773(.A1(new_n8392_), .A2(new_n8390_), .B(new_n8398_), .ZN(new_n8854_));
  NAND2_X1   g08774(.A1(new_n8854_), .A2(new_n8853_), .ZN(new_n8855_));
  NAND3_X1   g08775(.A1(new_n8670_), .A2(new_n8669_), .A3(new_n8671_), .ZN(new_n8856_));
  OAI21_X1   g08776(.A1(new_n8664_), .A2(new_n8660_), .B(new_n8667_), .ZN(new_n8857_));
  AOI21_X1   g08777(.A1(new_n8857_), .A2(new_n8856_), .B(new_n8853_), .ZN(new_n8858_));
  OAI21_X1   g08778(.A1(new_n8858_), .A2(new_n8657_), .B(new_n8855_), .ZN(new_n8859_));
  AOI21_X1   g08779(.A1(new_n8383_), .A2(new_n8387_), .B(new_n8859_), .ZN(new_n8860_));
  NAND3_X1   g08780(.A1(new_n8859_), .A2(new_n8383_), .A3(new_n8387_), .ZN(new_n8861_));
  AOI21_X1   g08781(.A1(new_n8861_), .A2(new_n8679_), .B(new_n8860_), .ZN(new_n8862_));
  NOR3_X1    g08782(.A1(new_n8690_), .A2(new_n8689_), .A3(new_n8691_), .ZN(new_n8863_));
  AOI21_X1   g08783(.A1(new_n8683_), .A2(new_n8684_), .B(new_n8687_), .ZN(new_n8864_));
  NOR2_X1    g08784(.A1(new_n8864_), .A2(new_n8863_), .ZN(new_n8865_));
  NAND2_X1   g08785(.A1(new_n8862_), .A2(new_n8865_), .ZN(new_n8866_));
  NAND2_X1   g08786(.A1(new_n8680_), .A2(new_n8675_), .ZN(new_n8867_));
  NAND2_X1   g08787(.A1(new_n8692_), .A2(new_n8688_), .ZN(new_n8868_));
  NAND2_X1   g08788(.A1(new_n8867_), .A2(new_n8868_), .ZN(new_n8869_));
  AOI22_X1   g08789(.A1(new_n5859_), .A2(new_n8832_), .B1(new_n4375_), .B2(new_n2898_), .ZN(new_n8870_));
  OAI21_X1   g08790(.A1(new_n8870_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n8871_));
  INV_X1     g08791(.I(new_n8871_), .ZN(new_n8872_));
  NAND3_X1   g08792(.A1(new_n4729_), .A2(new_n4728_), .A3(new_n8872_), .ZN(new_n8873_));
  INV_X1     g08793(.I(new_n8873_), .ZN(new_n8874_));
  AOI21_X1   g08794(.A1(new_n4729_), .A2(new_n4728_), .B(new_n8872_), .ZN(new_n8875_));
  NOR2_X1    g08795(.A1(new_n8874_), .A2(new_n8875_), .ZN(new_n8876_));
  NAND3_X1   g08796(.A1(new_n8866_), .A2(new_n8876_), .A3(new_n8869_), .ZN(new_n8877_));
  NOR2_X1    g08797(.A1(new_n8867_), .A2(new_n8868_), .ZN(new_n8878_));
  INV_X1     g08798(.I(new_n8869_), .ZN(new_n8879_));
  INV_X1     g08799(.I(new_n8875_), .ZN(new_n8880_));
  NAND2_X1   g08800(.A1(new_n8880_), .A2(new_n8873_), .ZN(new_n8881_));
  OAI21_X1   g08801(.A1(new_n8879_), .A2(new_n8878_), .B(new_n8881_), .ZN(new_n8882_));
  NAND2_X1   g08802(.A1(new_n8882_), .A2(new_n8877_), .ZN(new_n8883_));
  NAND3_X1   g08803(.A1(new_n8388_), .A2(new_n8859_), .A3(new_n8678_), .ZN(new_n8884_));
  AOI21_X1   g08804(.A1(new_n8388_), .A2(new_n8678_), .B(new_n8859_), .ZN(new_n8885_));
  INV_X1     g08805(.I(new_n8885_), .ZN(new_n8886_));
  AOI21_X1   g08806(.A1(new_n8886_), .A2(new_n8884_), .B(new_n8672_), .ZN(new_n8887_));
  INV_X1     g08807(.I(new_n8884_), .ZN(new_n8888_));
  NOR3_X1    g08808(.A1(new_n8888_), .A2(new_n8857_), .A3(new_n8885_), .ZN(new_n8889_));
  INV_X1     g08809(.I(new_n8620_), .ZN(new_n8890_));
  AOI21_X1   g08810(.A1(new_n8416_), .A2(new_n8418_), .B(new_n8623_), .ZN(new_n8891_));
  INV_X1     g08811(.I(new_n8891_), .ZN(new_n8892_));
  NOR2_X1    g08812(.A1(new_n8892_), .A2(new_n8617_), .ZN(new_n8893_));
  INV_X1     g08813(.I(new_n8893_), .ZN(new_n8894_));
  NAND2_X1   g08814(.A1(new_n8892_), .A2(new_n8617_), .ZN(new_n8895_));
  AOI21_X1   g08815(.A1(new_n8894_), .A2(new_n8895_), .B(new_n8890_), .ZN(new_n8896_));
  INV_X1     g08816(.I(new_n8895_), .ZN(new_n8897_));
  NOR3_X1    g08817(.A1(new_n8897_), .A2(new_n8893_), .A3(new_n8620_), .ZN(new_n8898_));
  NOR2_X1    g08818(.A1(new_n8896_), .A2(new_n8898_), .ZN(new_n8899_));
  NAND3_X1   g08819(.A1(new_n8557_), .A2(new_n8559_), .A3(new_n8562_), .ZN(new_n8900_));
  OAI21_X1   g08820(.A1(new_n8566_), .A2(new_n8556_), .B(new_n8563_), .ZN(new_n8901_));
  AOI22_X1   g08821(.A1(new_n8553_), .A2(new_n8548_), .B1(new_n8901_), .B2(new_n8900_), .ZN(new_n8902_));
  NAND2_X1   g08822(.A1(new_n8553_), .A2(new_n8548_), .ZN(new_n8903_));
  NOR2_X1    g08823(.A1(new_n8567_), .A2(new_n8564_), .ZN(new_n8904_));
  NOR2_X1    g08824(.A1(new_n8903_), .A2(new_n8904_), .ZN(new_n8905_));
  NOR2_X1    g08825(.A1(new_n8905_), .A2(new_n8902_), .ZN(new_n8906_));
  AOI22_X1   g08826(.A1(new_n6961_), .A2(new_n8832_), .B1(new_n4297_), .B2(new_n2898_), .ZN(new_n8907_));
  OAI21_X1   g08827(.A1(new_n8907_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n8908_));
  XOR2_X1    g08828(.A1(new_n5753_), .A2(new_n8908_), .Z(new_n8909_));
  XNOR2_X1   g08829(.A1(new_n8511_), .A2(new_n8508_), .ZN(new_n8910_));
  NOR2_X1    g08830(.A1(new_n8910_), .A2(new_n8507_), .ZN(new_n8911_));
  INV_X1     g08831(.I(new_n8512_), .ZN(new_n8912_));
  AOI21_X1   g08832(.A1(new_n8912_), .A2(new_n8513_), .B(new_n8506_), .ZN(new_n8913_));
  NOR2_X1    g08833(.A1(new_n8911_), .A2(new_n8913_), .ZN(new_n8914_));
  INV_X1     g08834(.I(new_n8914_), .ZN(new_n8915_));
  OAI21_X1   g08835(.A1(new_n4234_), .A2(new_n4244_), .B(new_n8832_), .ZN(new_n8916_));
  NAND2_X1   g08836(.A1(new_n4221_), .A2(new_n2898_), .ZN(new_n8917_));
  AOI21_X1   g08837(.A1(new_n8917_), .A2(new_n8916_), .B(\a[5] ), .ZN(new_n8918_));
  NOR2_X1    g08838(.A1(new_n8918_), .A2(new_n3040_), .ZN(new_n8919_));
  INV_X1     g08839(.I(new_n8919_), .ZN(new_n8920_));
  NOR2_X1    g08840(.A1(new_n8920_), .A2(new_n5648_), .ZN(new_n8921_));
  NOR2_X1    g08841(.A1(new_n6245_), .A2(new_n8919_), .ZN(new_n8922_));
  NOR2_X1    g08842(.A1(new_n8921_), .A2(new_n8922_), .ZN(new_n8923_));
  NOR2_X1    g08843(.A1(new_n8923_), .A2(new_n8490_), .ZN(new_n8924_));
  INV_X1     g08844(.I(new_n8924_), .ZN(new_n8925_));
  NOR2_X1    g08845(.A1(new_n6061_), .A2(new_n2898_), .ZN(new_n8926_));
  OAI21_X1   g08846(.A1(new_n5627_), .A2(new_n3040_), .B(new_n4234_), .ZN(new_n8927_));
  NOR2_X1    g08847(.A1(new_n8927_), .A2(new_n8926_), .ZN(new_n8928_));
  OAI22_X1   g08848(.A1(new_n4244_), .A2(new_n8830_), .B1(new_n3042_), .B2(new_n4230_), .ZN(new_n8929_));
  OAI21_X1   g08849(.A1(new_n3040_), .A2(new_n4234_), .B(new_n8929_), .ZN(new_n8930_));
  NOR2_X1    g08850(.A1(new_n8928_), .A2(new_n8930_), .ZN(new_n8931_));
  NOR2_X1    g08851(.A1(new_n8931_), .A2(\a[5] ), .ZN(new_n8932_));
  NAND2_X1   g08852(.A1(new_n8931_), .A2(\a[5] ), .ZN(new_n8933_));
  INV_X1     g08853(.I(new_n8933_), .ZN(new_n8934_));
  NOR2_X1    g08854(.A1(new_n8934_), .A2(new_n8932_), .ZN(new_n8935_));
  INV_X1     g08855(.I(new_n5637_), .ZN(new_n8936_));
  AOI21_X1   g08856(.A1(new_n4251_), .A2(new_n2898_), .B(\a[5] ), .ZN(new_n8937_));
  OAI21_X1   g08857(.A1(new_n3042_), .A2(new_n4244_), .B(new_n8937_), .ZN(new_n8938_));
  NAND2_X1   g08858(.A1(new_n8938_), .A2(new_n2898_), .ZN(new_n8939_));
  NOR2_X1    g08859(.A1(new_n8939_), .A2(new_n8936_), .ZN(new_n8940_));
  AOI21_X1   g08860(.A1(new_n2898_), .A2(new_n8938_), .B(new_n5637_), .ZN(new_n8941_));
  NOR2_X1    g08861(.A1(new_n4251_), .A2(new_n3419_), .ZN(new_n8942_));
  NOR4_X1    g08862(.A1(new_n8941_), .A2(new_n8940_), .A3(new_n452_), .A4(new_n8942_), .ZN(new_n8943_));
  NAND2_X1   g08863(.A1(new_n8935_), .A2(new_n8943_), .ZN(new_n8944_));
  NAND2_X1   g08864(.A1(new_n8923_), .A2(new_n8490_), .ZN(new_n8945_));
  NAND2_X1   g08865(.A1(new_n8944_), .A2(new_n8945_), .ZN(new_n8946_));
  NAND2_X1   g08866(.A1(new_n8946_), .A2(new_n8925_), .ZN(new_n8947_));
  XOR2_X1    g08867(.A1(new_n8489_), .A2(new_n8491_), .Z(new_n8948_));
  OAI22_X1   g08868(.A1(new_n4203_), .A2(new_n3040_), .B1(new_n6529_), .B2(new_n8831_), .ZN(new_n8949_));
  AOI21_X1   g08869(.A1(new_n8949_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n8950_));
  NAND2_X1   g08870(.A1(new_n6082_), .A2(new_n8950_), .ZN(new_n8951_));
  INV_X1     g08871(.I(new_n8950_), .ZN(new_n8952_));
  NAND2_X1   g08872(.A1(new_n5660_), .A2(new_n8952_), .ZN(new_n8953_));
  NAND2_X1   g08873(.A1(new_n8953_), .A2(new_n8951_), .ZN(new_n8954_));
  OAI21_X1   g08874(.A1(new_n8948_), .A2(new_n8954_), .B(new_n8947_), .ZN(new_n8955_));
  INV_X1     g08875(.I(new_n8948_), .ZN(new_n8956_));
  NOR2_X1    g08876(.A1(new_n5660_), .A2(new_n8952_), .ZN(new_n8957_));
  NOR2_X1    g08877(.A1(new_n6082_), .A2(new_n8950_), .ZN(new_n8958_));
  NOR2_X1    g08878(.A1(new_n8957_), .A2(new_n8958_), .ZN(new_n8959_));
  NOR2_X1    g08879(.A1(new_n8959_), .A2(new_n8956_), .ZN(new_n8960_));
  INV_X1     g08880(.I(new_n8960_), .ZN(new_n8961_));
  NAND2_X1   g08881(.A1(new_n8955_), .A2(new_n8961_), .ZN(new_n8962_));
  XNOR2_X1   g08882(.A1(new_n8485_), .A2(new_n8493_), .ZN(new_n8963_));
  INV_X1     g08883(.I(new_n8963_), .ZN(new_n8964_));
  AOI22_X1   g08884(.A1(new_n4258_), .A2(new_n2898_), .B1(new_n6541_), .B2(new_n8832_), .ZN(new_n8965_));
  OAI21_X1   g08885(.A1(new_n8965_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n8966_));
  XOR2_X1    g08886(.A1(new_n5671_), .A2(new_n8966_), .Z(new_n8967_));
  NAND2_X1   g08887(.A1(new_n8967_), .A2(new_n8964_), .ZN(new_n8968_));
  NOR2_X1    g08888(.A1(new_n8967_), .A2(new_n8964_), .ZN(new_n8969_));
  AOI21_X1   g08889(.A1(new_n8962_), .A2(new_n8968_), .B(new_n8969_), .ZN(new_n8970_));
  INV_X1     g08890(.I(new_n8970_), .ZN(new_n8971_));
  XOR2_X1    g08891(.A1(new_n8477_), .A2(new_n8496_), .Z(new_n8972_));
  NAND2_X1   g08892(.A1(new_n8972_), .A2(new_n8495_), .ZN(new_n8973_));
  OAI21_X1   g08893(.A1(new_n8479_), .A2(new_n8497_), .B(new_n8494_), .ZN(new_n8974_));
  NAND2_X1   g08894(.A1(new_n8973_), .A2(new_n8974_), .ZN(new_n8975_));
  INV_X1     g08895(.I(new_n8975_), .ZN(new_n8976_));
  OAI22_X1   g08896(.A1(new_n5684_), .A2(new_n3040_), .B1(new_n6556_), .B2(new_n8831_), .ZN(new_n8977_));
  AOI21_X1   g08897(.A1(new_n8977_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n8978_));
  XOR2_X1    g08898(.A1(new_n6102_), .A2(new_n8978_), .Z(new_n8979_));
  NAND2_X1   g08899(.A1(new_n8979_), .A2(new_n8976_), .ZN(new_n8980_));
  NAND2_X1   g08900(.A1(new_n8971_), .A2(new_n8980_), .ZN(new_n8981_));
  XOR2_X1    g08901(.A1(new_n5693_), .A2(new_n8978_), .Z(new_n8982_));
  NAND2_X1   g08902(.A1(new_n8982_), .A2(new_n8975_), .ZN(new_n8983_));
  NAND2_X1   g08903(.A1(new_n8981_), .A2(new_n8983_), .ZN(new_n8984_));
  INV_X1     g08904(.I(new_n8500_), .ZN(new_n8985_));
  XOR2_X1    g08905(.A1(new_n8503_), .A2(new_n8985_), .Z(new_n8986_));
  NOR2_X1    g08906(.A1(new_n8986_), .A2(new_n8499_), .ZN(new_n8987_));
  INV_X1     g08907(.I(new_n8499_), .ZN(new_n8988_));
  INV_X1     g08908(.I(new_n8504_), .ZN(new_n8989_));
  AOI21_X1   g08909(.A1(new_n8989_), .A2(new_n8505_), .B(new_n8988_), .ZN(new_n8990_));
  NOR2_X1    g08910(.A1(new_n8987_), .A2(new_n8990_), .ZN(new_n8991_));
  OAI22_X1   g08911(.A1(new_n4150_), .A2(new_n3040_), .B1(new_n6567_), .B2(new_n8831_), .ZN(new_n8992_));
  AOI21_X1   g08912(.A1(new_n8992_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n8993_));
  XOR2_X1    g08913(.A1(new_n5707_), .A2(new_n8993_), .Z(new_n8994_));
  INV_X1     g08914(.I(new_n8994_), .ZN(new_n8995_));
  NAND2_X1   g08915(.A1(new_n8995_), .A2(new_n8991_), .ZN(new_n8996_));
  OAI21_X1   g08916(.A1(new_n8987_), .A2(new_n8990_), .B(new_n8994_), .ZN(new_n8997_));
  NAND2_X1   g08917(.A1(new_n8996_), .A2(new_n8997_), .ZN(new_n8998_));
  NOR2_X1    g08918(.A1(new_n8984_), .A2(new_n8998_), .ZN(new_n8999_));
  NAND2_X1   g08919(.A1(new_n8999_), .A2(new_n8915_), .ZN(new_n9000_));
  AOI22_X1   g08920(.A1(new_n6582_), .A2(new_n8832_), .B1(new_n4274_), .B2(new_n2898_), .ZN(new_n9001_));
  OAI21_X1   g08921(.A1(new_n9001_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9002_));
  XOR2_X1    g08922(.A1(new_n5722_), .A2(new_n9002_), .Z(new_n9003_));
  NOR2_X1    g08923(.A1(new_n9003_), .A2(new_n8997_), .ZN(new_n9004_));
  OAI21_X1   g08924(.A1(new_n8999_), .A2(new_n8915_), .B(new_n9004_), .ZN(new_n9005_));
  NAND2_X1   g08925(.A1(new_n9005_), .A2(new_n9000_), .ZN(new_n9006_));
  INV_X1     g08926(.I(new_n8514_), .ZN(new_n9007_));
  XNOR2_X1   g08927(.A1(new_n8460_), .A2(new_n8454_), .ZN(new_n9008_));
  NOR2_X1    g08928(.A1(new_n9008_), .A2(new_n9007_), .ZN(new_n9009_));
  OR2_X2     g08929(.A1(new_n8460_), .A2(new_n8454_), .Z(new_n9010_));
  NAND2_X1   g08930(.A1(new_n8460_), .A2(new_n8454_), .ZN(new_n9011_));
  AOI21_X1   g08931(.A1(new_n9010_), .A2(new_n9011_), .B(new_n8514_), .ZN(new_n9012_));
  NOR2_X1    g08932(.A1(new_n9009_), .A2(new_n9012_), .ZN(new_n9013_));
  INV_X1     g08933(.I(new_n9013_), .ZN(new_n9014_));
  OAI22_X1   g08934(.A1(new_n4142_), .A2(new_n3040_), .B1(new_n4277_), .B2(new_n8831_), .ZN(new_n9015_));
  AOI21_X1   g08935(.A1(new_n9015_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n9016_));
  XOR2_X1    g08936(.A1(new_n6134_), .A2(new_n9016_), .Z(new_n9017_));
  NAND2_X1   g08937(.A1(new_n9014_), .A2(new_n9017_), .ZN(new_n9018_));
  NAND2_X1   g08938(.A1(new_n9006_), .A2(new_n9018_), .ZN(new_n9019_));
  INV_X1     g08939(.I(new_n9017_), .ZN(new_n9020_));
  NAND2_X1   g08940(.A1(new_n9013_), .A2(new_n9020_), .ZN(new_n9021_));
  NAND2_X1   g08941(.A1(new_n9019_), .A2(new_n9021_), .ZN(new_n9022_));
  INV_X1     g08942(.I(new_n9022_), .ZN(new_n9023_));
  NOR2_X1    g08943(.A1(new_n8471_), .A2(new_n9008_), .ZN(new_n9024_));
  NAND2_X1   g08944(.A1(new_n9024_), .A2(new_n9011_), .ZN(new_n9025_));
  NAND2_X1   g08945(.A1(new_n8460_), .A2(new_n8454_), .ZN(new_n9026_));
  AOI21_X1   g08946(.A1(new_n9025_), .A2(new_n9026_), .B(new_n8514_), .ZN(new_n9027_));
  INV_X1     g08947(.I(new_n9027_), .ZN(new_n9028_));
  NAND3_X1   g08948(.A1(new_n9025_), .A2(new_n8514_), .A3(new_n9026_), .ZN(new_n9029_));
  NAND2_X1   g08949(.A1(new_n6609_), .A2(new_n8832_), .ZN(new_n9030_));
  OAI21_X1   g08950(.A1(new_n4135_), .A2(new_n3040_), .B(new_n9030_), .ZN(new_n9031_));
  AOI21_X1   g08951(.A1(new_n9031_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n9032_));
  XNOR2_X1   g08952(.A1(new_n5624_), .A2(new_n9032_), .ZN(new_n9033_));
  INV_X1     g08953(.I(new_n9033_), .ZN(new_n9034_));
  AOI21_X1   g08954(.A1(new_n9028_), .A2(new_n9029_), .B(new_n9034_), .ZN(new_n9035_));
  NAND3_X1   g08955(.A1(new_n9028_), .A2(new_n9029_), .A3(new_n9034_), .ZN(new_n9036_));
  OAI21_X1   g08956(.A1(new_n9023_), .A2(new_n9035_), .B(new_n9036_), .ZN(new_n9037_));
  INV_X1     g08957(.I(new_n9037_), .ZN(new_n9038_));
  OAI22_X1   g08958(.A1(new_n4285_), .A2(new_n3040_), .B1(new_n6621_), .B2(new_n8831_), .ZN(new_n9039_));
  NAND2_X1   g08959(.A1(new_n9039_), .A2(new_n452_), .ZN(new_n9040_));
  NAND2_X1   g08960(.A1(new_n9040_), .A2(new_n2898_), .ZN(new_n9041_));
  XOR2_X1    g08961(.A1(new_n5023_), .A2(new_n9041_), .Z(new_n9042_));
  XOR2_X1    g08962(.A1(new_n8449_), .A2(new_n7528_), .Z(new_n9043_));
  NAND3_X1   g08963(.A1(new_n8517_), .A2(new_n9043_), .A3(new_n8521_), .ZN(new_n9044_));
  NOR2_X1    g08964(.A1(new_n8473_), .A2(new_n8516_), .ZN(new_n9045_));
  INV_X1     g08965(.I(new_n8521_), .ZN(new_n9046_));
  OAI21_X1   g08966(.A1(new_n8450_), .A2(new_n9046_), .B(new_n9045_), .ZN(new_n9047_));
  AOI21_X1   g08967(.A1(new_n9044_), .A2(new_n9047_), .B(new_n8470_), .ZN(new_n9048_));
  INV_X1     g08968(.I(new_n9048_), .ZN(new_n9049_));
  NAND3_X1   g08969(.A1(new_n9044_), .A2(new_n9047_), .A3(new_n8470_), .ZN(new_n9050_));
  NAND3_X1   g08970(.A1(new_n9049_), .A2(new_n9050_), .A3(new_n9042_), .ZN(new_n9051_));
  INV_X1     g08971(.I(new_n9042_), .ZN(new_n9052_));
  INV_X1     g08972(.I(new_n9050_), .ZN(new_n9053_));
  OAI21_X1   g08973(.A1(new_n9053_), .A2(new_n9048_), .B(new_n9052_), .ZN(new_n9054_));
  NAND3_X1   g08974(.A1(new_n9051_), .A2(new_n9054_), .A3(new_n9038_), .ZN(new_n9055_));
  NOR2_X1    g08975(.A1(new_n9055_), .A2(new_n8909_), .ZN(new_n9056_));
  NOR3_X1    g08976(.A1(new_n9053_), .A2(new_n9052_), .A3(new_n9048_), .ZN(new_n9057_));
  INV_X1     g08977(.I(new_n8533_), .ZN(new_n9058_));
  OAI22_X1   g08978(.A1(new_n8523_), .A2(new_n8518_), .B1(new_n8532_), .B2(new_n9058_), .ZN(new_n9059_));
  XOR2_X1    g08979(.A1(new_n8527_), .A2(new_n8531_), .Z(new_n9060_));
  NAND2_X1   g08980(.A1(new_n8524_), .A2(new_n9060_), .ZN(new_n9061_));
  NAND2_X1   g08981(.A1(new_n9061_), .A2(new_n9059_), .ZN(new_n9062_));
  NAND2_X1   g08982(.A1(new_n9057_), .A2(new_n9062_), .ZN(new_n9063_));
  AOI21_X1   g08983(.A1(new_n9055_), .A2(new_n8909_), .B(new_n9063_), .ZN(new_n9064_));
  XOR2_X1    g08984(.A1(new_n8538_), .A2(new_n8542_), .Z(new_n9065_));
  AND2_X2    g08985(.A1(new_n8534_), .A2(new_n9065_), .Z(new_n9066_));
  INV_X1     g08986(.I(new_n8543_), .ZN(new_n9067_));
  NOR2_X1    g08987(.A1(new_n9067_), .A2(new_n8544_), .ZN(new_n9068_));
  NOR2_X1    g08988(.A1(new_n8534_), .A2(new_n9068_), .ZN(new_n9069_));
  OAI22_X1   g08989(.A1(new_n4131_), .A2(new_n3040_), .B1(new_n4301_), .B2(new_n8831_), .ZN(new_n9070_));
  AOI21_X1   g08990(.A1(new_n9070_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n9071_));
  XNOR2_X1   g08991(.A1(new_n5599_), .A2(new_n9071_), .ZN(new_n9072_));
  OAI21_X1   g08992(.A1(new_n9066_), .A2(new_n9069_), .B(new_n9072_), .ZN(new_n9073_));
  OAI21_X1   g08993(.A1(new_n9064_), .A2(new_n9056_), .B(new_n9073_), .ZN(new_n9074_));
  NAND2_X1   g08994(.A1(new_n8534_), .A2(new_n9065_), .ZN(new_n9075_));
  INV_X1     g08995(.I(new_n9069_), .ZN(new_n9076_));
  INV_X1     g08996(.I(new_n9072_), .ZN(new_n9077_));
  NAND3_X1   g08997(.A1(new_n9076_), .A2(new_n9075_), .A3(new_n9077_), .ZN(new_n9078_));
  NAND2_X1   g08998(.A1(new_n9074_), .A2(new_n9078_), .ZN(new_n9079_));
  NAND2_X1   g08999(.A1(new_n8546_), .A2(new_n8445_), .ZN(new_n9080_));
  NAND2_X1   g09000(.A1(new_n8446_), .A2(new_n8545_), .ZN(new_n9081_));
  NAND2_X1   g09001(.A1(new_n9081_), .A2(new_n9080_), .ZN(new_n9082_));
  AOI22_X1   g09002(.A1(new_n6980_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n5041_), .ZN(new_n9083_));
  OAI21_X1   g09003(.A1(new_n9083_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9084_));
  XOR2_X1    g09004(.A1(new_n5049_), .A2(new_n9084_), .Z(new_n9085_));
  NOR2_X1    g09005(.A1(new_n9082_), .A2(new_n9085_), .ZN(new_n9086_));
  INV_X1     g09006(.I(new_n9085_), .ZN(new_n9087_));
  AOI21_X1   g09007(.A1(new_n9081_), .A2(new_n9080_), .B(new_n9087_), .ZN(new_n9088_));
  AOI21_X1   g09008(.A1(new_n8432_), .A2(new_n8429_), .B(new_n8551_), .ZN(new_n9089_));
  INV_X1     g09009(.I(new_n9089_), .ZN(new_n9090_));
  AOI21_X1   g09010(.A1(new_n8545_), .A2(new_n8445_), .B(new_n9090_), .ZN(new_n9091_));
  NAND3_X1   g09011(.A1(new_n9090_), .A2(new_n8445_), .A3(new_n8545_), .ZN(new_n9092_));
  INV_X1     g09012(.I(new_n9092_), .ZN(new_n9093_));
  OAI21_X1   g09013(.A1(new_n9093_), .A2(new_n9091_), .B(new_n8442_), .ZN(new_n9094_));
  INV_X1     g09014(.I(new_n9094_), .ZN(new_n9095_));
  NOR3_X1    g09015(.A1(new_n9093_), .A2(new_n9091_), .A3(new_n8442_), .ZN(new_n9096_));
  AOI22_X1   g09016(.A1(new_n6993_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4124_), .ZN(new_n9097_));
  OAI21_X1   g09017(.A1(new_n9097_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9098_));
  XOR2_X1    g09018(.A1(new_n5067_), .A2(new_n9098_), .Z(new_n9099_));
  NOR3_X1    g09019(.A1(new_n9095_), .A2(new_n9099_), .A3(new_n9096_), .ZN(new_n9100_));
  INV_X1     g09020(.I(new_n9096_), .ZN(new_n9101_));
  INV_X1     g09021(.I(new_n9099_), .ZN(new_n9102_));
  AOI21_X1   g09022(.A1(new_n9101_), .A2(new_n9094_), .B(new_n9102_), .ZN(new_n9103_));
  OR2_X2     g09023(.A1(new_n9086_), .A2(new_n9088_), .Z(new_n9104_));
  NAND2_X1   g09024(.A1(new_n9104_), .A2(new_n9079_), .ZN(new_n9105_));
  NOR2_X1    g09025(.A1(new_n9105_), .A2(new_n8906_), .ZN(new_n9106_));
  NAND2_X1   g09026(.A1(new_n9105_), .A2(new_n8906_), .ZN(new_n9107_));
  OAI22_X1   g09027(.A1(new_n4112_), .A2(new_n3040_), .B1(new_n6682_), .B2(new_n8831_), .ZN(new_n9108_));
  AOI21_X1   g09028(.A1(new_n9108_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n9109_));
  XOR2_X1    g09029(.A1(new_n5096_), .A2(new_n9109_), .Z(new_n9110_));
  INV_X1     g09030(.I(new_n9110_), .ZN(new_n9111_));
  NAND2_X1   g09031(.A1(new_n9103_), .A2(new_n9111_), .ZN(new_n9112_));
  INV_X1     g09032(.I(new_n9112_), .ZN(new_n9113_));
  AOI21_X1   g09033(.A1(new_n9107_), .A2(new_n9113_), .B(new_n9106_), .ZN(new_n9114_));
  INV_X1     g09034(.I(new_n8571_), .ZN(new_n9115_));
  NOR3_X1    g09035(.A1(new_n8565_), .A2(new_n8095_), .A3(new_n8567_), .ZN(new_n9116_));
  OAI21_X1   g09036(.A1(new_n8565_), .A2(new_n8567_), .B(new_n8095_), .ZN(new_n9117_));
  INV_X1     g09037(.I(new_n9117_), .ZN(new_n9118_));
  OAI21_X1   g09038(.A1(new_n9118_), .A2(new_n9116_), .B(new_n8576_), .ZN(new_n9119_));
  INV_X1     g09039(.I(new_n9116_), .ZN(new_n9120_));
  NAND3_X1   g09040(.A1(new_n9120_), .A2(new_n8573_), .A3(new_n9117_), .ZN(new_n9121_));
  AOI21_X1   g09041(.A1(new_n9119_), .A2(new_n9121_), .B(new_n9115_), .ZN(new_n9122_));
  AOI21_X1   g09042(.A1(new_n9120_), .A2(new_n9117_), .B(new_n8573_), .ZN(new_n9123_));
  INV_X1     g09043(.I(new_n9121_), .ZN(new_n9124_));
  NOR3_X1    g09044(.A1(new_n9124_), .A2(new_n9123_), .A3(new_n8571_), .ZN(new_n9125_));
  AOI22_X1   g09045(.A1(new_n7015_), .A2(new_n8832_), .B1(new_n4105_), .B2(new_n2898_), .ZN(new_n9126_));
  OAI21_X1   g09046(.A1(new_n9126_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9127_));
  XOR2_X1    g09047(.A1(new_n5121_), .A2(new_n9127_), .Z(new_n9128_));
  INV_X1     g09048(.I(new_n9128_), .ZN(new_n9129_));
  NOR3_X1    g09049(.A1(new_n9125_), .A2(new_n9122_), .A3(new_n9129_), .ZN(new_n9130_));
  NOR2_X1    g09050(.A1(new_n9130_), .A2(new_n9114_), .ZN(new_n9131_));
  OAI21_X1   g09051(.A1(new_n9124_), .A2(new_n9123_), .B(new_n8571_), .ZN(new_n9132_));
  NAND3_X1   g09052(.A1(new_n9119_), .A2(new_n9121_), .A3(new_n9115_), .ZN(new_n9133_));
  AOI21_X1   g09053(.A1(new_n9132_), .A2(new_n9133_), .B(new_n9128_), .ZN(new_n9134_));
  NOR2_X1    g09054(.A1(new_n8575_), .A2(new_n8572_), .ZN(new_n9135_));
  AOI21_X1   g09055(.A1(new_n8587_), .A2(new_n8592_), .B(new_n9135_), .ZN(new_n9136_));
  AOI22_X1   g09056(.A1(new_n7021_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4100_), .ZN(new_n9137_));
  OAI21_X1   g09057(.A1(new_n9137_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9138_));
  XOR2_X1    g09058(.A1(new_n5080_), .A2(new_n9138_), .Z(new_n9139_));
  INV_X1     g09059(.I(new_n9139_), .ZN(new_n9140_));
  NOR3_X1    g09060(.A1(new_n9136_), .A2(new_n8590_), .A3(new_n9140_), .ZN(new_n9141_));
  INV_X1     g09061(.I(new_n9141_), .ZN(new_n9142_));
  OAI21_X1   g09062(.A1(new_n9131_), .A2(new_n9134_), .B(new_n9142_), .ZN(new_n9143_));
  OAI21_X1   g09063(.A1(new_n9136_), .A2(new_n8590_), .B(new_n9140_), .ZN(new_n9144_));
  NAND2_X1   g09064(.A1(new_n9143_), .A2(new_n9144_), .ZN(new_n9145_));
  INV_X1     g09065(.I(new_n8590_), .ZN(new_n9146_));
  INV_X1     g09066(.I(new_n8424_), .ZN(new_n9147_));
  NOR2_X1    g09067(.A1(new_n9147_), .A2(new_n8595_), .ZN(new_n9148_));
  NAND2_X1   g09068(.A1(new_n9146_), .A2(new_n9148_), .ZN(new_n9149_));
  OAI21_X1   g09069(.A1(new_n9147_), .A2(new_n8595_), .B(new_n8590_), .ZN(new_n9150_));
  AOI21_X1   g09070(.A1(new_n9149_), .A2(new_n9150_), .B(new_n8589_), .ZN(new_n9151_));
  NAND3_X1   g09071(.A1(new_n9149_), .A2(new_n8589_), .A3(new_n9150_), .ZN(new_n9152_));
  INV_X1     g09072(.I(new_n9152_), .ZN(new_n9153_));
  OAI22_X1   g09073(.A1(new_n4090_), .A2(new_n3040_), .B1(new_n4320_), .B2(new_n8831_), .ZN(new_n9154_));
  AOI21_X1   g09074(.A1(new_n9154_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n9155_));
  XOR2_X1    g09075(.A1(new_n5196_), .A2(new_n9155_), .Z(new_n9156_));
  OAI21_X1   g09076(.A1(new_n9153_), .A2(new_n9151_), .B(new_n9156_), .ZN(new_n9157_));
  INV_X1     g09077(.I(new_n9151_), .ZN(new_n9158_));
  INV_X1     g09078(.I(new_n9156_), .ZN(new_n9159_));
  NAND3_X1   g09079(.A1(new_n9158_), .A2(new_n9152_), .A3(new_n9159_), .ZN(new_n9160_));
  INV_X1     g09080(.I(new_n9160_), .ZN(new_n9161_));
  AOI21_X1   g09081(.A1(new_n9145_), .A2(new_n9157_), .B(new_n9161_), .ZN(new_n9162_));
  NAND2_X1   g09082(.A1(new_n8597_), .A2(new_n8591_), .ZN(new_n9163_));
  XOR2_X1    g09083(.A1(new_n8603_), .A2(new_n8606_), .Z(new_n9164_));
  NAND2_X1   g09084(.A1(new_n9163_), .A2(new_n9164_), .ZN(new_n9165_));
  XNOR2_X1   g09085(.A1(new_n8603_), .A2(new_n8606_), .ZN(new_n9166_));
  NAND3_X1   g09086(.A1(new_n9166_), .A2(new_n8591_), .A3(new_n8597_), .ZN(new_n9167_));
  NAND2_X1   g09087(.A1(new_n9167_), .A2(new_n9165_), .ZN(new_n9168_));
  AOI22_X1   g09088(.A1(new_n6419_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4328_), .ZN(new_n9169_));
  OAI21_X1   g09089(.A1(new_n9169_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9170_));
  XNOR2_X1   g09090(.A1(new_n5139_), .A2(new_n9170_), .ZN(new_n9171_));
  NOR2_X1    g09091(.A1(new_n9168_), .A2(new_n9171_), .ZN(new_n9172_));
  NAND2_X1   g09092(.A1(new_n9168_), .A2(new_n9171_), .ZN(new_n9173_));
  INV_X1     g09093(.I(new_n9173_), .ZN(new_n9174_));
  NOR2_X1    g09094(.A1(new_n8613_), .A2(new_n8616_), .ZN(new_n9175_));
  AOI22_X1   g09095(.A1(new_n4333_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4082_), .ZN(new_n9176_));
  OAI21_X1   g09096(.A1(new_n9176_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9177_));
  XNOR2_X1   g09097(.A1(new_n5162_), .A2(new_n9177_), .ZN(new_n9178_));
  XNOR2_X1   g09098(.A1(new_n9175_), .A2(new_n9178_), .ZN(new_n9179_));
  OAI21_X1   g09099(.A1(new_n8607_), .A2(new_n8608_), .B(new_n9179_), .ZN(new_n9180_));
  NOR2_X1    g09100(.A1(new_n8607_), .A2(new_n8608_), .ZN(new_n9181_));
  XOR2_X1    g09101(.A1(new_n9175_), .A2(new_n9178_), .Z(new_n9182_));
  NAND2_X1   g09102(.A1(new_n9182_), .A2(new_n9181_), .ZN(new_n9183_));
  NAND2_X1   g09103(.A1(new_n9180_), .A2(new_n9183_), .ZN(new_n9184_));
  NOR2_X1    g09104(.A1(new_n9174_), .A2(new_n9172_), .ZN(new_n9186_));
  NOR2_X1    g09105(.A1(new_n9162_), .A2(new_n9186_), .ZN(new_n9187_));
  INV_X1     g09106(.I(new_n9187_), .ZN(new_n9188_));
  NOR2_X1    g09107(.A1(new_n9188_), .A2(new_n8899_), .ZN(new_n9189_));
  XOR2_X1    g09108(.A1(new_n9181_), .A2(new_n9175_), .Z(new_n9190_));
  NAND2_X1   g09109(.A1(new_n9190_), .A2(new_n9178_), .ZN(new_n9191_));
  OAI22_X1   g09110(.A1(new_n4070_), .A2(new_n3040_), .B1(new_n5917_), .B2(new_n8831_), .ZN(new_n9192_));
  AOI21_X1   g09111(.A1(new_n9192_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n9193_));
  XOR2_X1    g09112(.A1(new_n4927_), .A2(new_n9193_), .Z(new_n9194_));
  NOR2_X1    g09113(.A1(new_n9191_), .A2(new_n9194_), .ZN(new_n9195_));
  INV_X1     g09114(.I(new_n9195_), .ZN(new_n9196_));
  AOI21_X1   g09115(.A1(new_n9188_), .A2(new_n8899_), .B(new_n9196_), .ZN(new_n9197_));
  NAND2_X1   g09116(.A1(new_n8625_), .A2(new_n8618_), .ZN(new_n9198_));
  NAND2_X1   g09117(.A1(new_n8636_), .A2(new_n8638_), .ZN(new_n9199_));
  NOR2_X1    g09118(.A1(new_n9199_), .A2(new_n9198_), .ZN(new_n9200_));
  INV_X1     g09119(.I(new_n9198_), .ZN(new_n9201_));
  INV_X1     g09120(.I(new_n9199_), .ZN(new_n9202_));
  NOR2_X1    g09121(.A1(new_n9202_), .A2(new_n9201_), .ZN(new_n9203_));
  AOI22_X1   g09122(.A1(new_n4923_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4061_), .ZN(new_n9204_));
  OAI21_X1   g09123(.A1(new_n9204_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9205_));
  XOR2_X1    g09124(.A1(new_n4935_), .A2(new_n9205_), .Z(new_n9206_));
  INV_X1     g09125(.I(new_n9206_), .ZN(new_n9207_));
  NOR3_X1    g09126(.A1(new_n9203_), .A2(new_n9200_), .A3(new_n9207_), .ZN(new_n9208_));
  INV_X1     g09127(.I(new_n9208_), .ZN(new_n9209_));
  OAI21_X1   g09128(.A1(new_n9197_), .A2(new_n9189_), .B(new_n9209_), .ZN(new_n9210_));
  OAI21_X1   g09129(.A1(new_n9203_), .A2(new_n9200_), .B(new_n9207_), .ZN(new_n9211_));
  INV_X1     g09130(.I(new_n8638_), .ZN(new_n9212_));
  NOR3_X1    g09131(.A1(new_n8646_), .A2(new_n9212_), .A3(new_n8644_), .ZN(new_n9213_));
  NOR3_X1    g09132(.A1(new_n9213_), .A2(new_n9198_), .A3(new_n9202_), .ZN(new_n9214_));
  INV_X1     g09133(.I(new_n9214_), .ZN(new_n9215_));
  OAI21_X1   g09134(.A1(new_n9213_), .A2(new_n9202_), .B(new_n9198_), .ZN(new_n9216_));
  AOI22_X1   g09135(.A1(new_n6428_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4054_), .ZN(new_n9217_));
  OAI21_X1   g09136(.A1(new_n9217_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9218_));
  XOR2_X1    g09137(.A1(new_n4652_), .A2(new_n9218_), .Z(new_n9219_));
  NAND3_X1   g09138(.A1(new_n9215_), .A2(new_n9216_), .A3(new_n9219_), .ZN(new_n9220_));
  INV_X1     g09139(.I(new_n9220_), .ZN(new_n9221_));
  AOI21_X1   g09140(.A1(new_n9210_), .A2(new_n9211_), .B(new_n9221_), .ZN(new_n9222_));
  AOI21_X1   g09141(.A1(new_n9215_), .A2(new_n9216_), .B(new_n9219_), .ZN(new_n9223_));
  INV_X1     g09142(.I(new_n8648_), .ZN(new_n9224_));
  AOI21_X1   g09143(.A1(new_n8407_), .A2(new_n8410_), .B(new_n8654_), .ZN(new_n9225_));
  NAND2_X1   g09144(.A1(new_n9225_), .A2(new_n9224_), .ZN(new_n9226_));
  NOR2_X1    g09145(.A1(new_n9225_), .A2(new_n9224_), .ZN(new_n9227_));
  INV_X1     g09146(.I(new_n9227_), .ZN(new_n9228_));
  AOI21_X1   g09147(.A1(new_n9228_), .A2(new_n9226_), .B(new_n8646_), .ZN(new_n9229_));
  INV_X1     g09148(.I(new_n9226_), .ZN(new_n9230_));
  NOR3_X1    g09149(.A1(new_n9230_), .A2(new_n8645_), .A3(new_n9227_), .ZN(new_n9231_));
  OAI22_X1   g09150(.A1(new_n4042_), .A2(new_n3040_), .B1(new_n4342_), .B2(new_n8831_), .ZN(new_n9232_));
  AOI21_X1   g09151(.A1(new_n9232_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n9233_));
  XNOR2_X1   g09152(.A1(new_n4864_), .A2(new_n9233_), .ZN(new_n9234_));
  OAI21_X1   g09153(.A1(new_n9229_), .A2(new_n9231_), .B(new_n9234_), .ZN(new_n9235_));
  OAI21_X1   g09154(.A1(new_n9222_), .A2(new_n9223_), .B(new_n9235_), .ZN(new_n9236_));
  NOR3_X1    g09155(.A1(new_n9229_), .A2(new_n9231_), .A3(new_n9234_), .ZN(new_n9237_));
  INV_X1     g09156(.I(new_n9237_), .ZN(new_n9238_));
  NAND2_X1   g09157(.A1(new_n8403_), .A2(new_n8657_), .ZN(new_n9239_));
  INV_X1     g09158(.I(new_n9239_), .ZN(new_n9240_));
  NOR2_X1    g09159(.A1(new_n8403_), .A2(new_n8657_), .ZN(new_n9241_));
  AOI22_X1   g09160(.A1(new_n4347_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4036_), .ZN(new_n9242_));
  OAI21_X1   g09161(.A1(new_n9242_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9243_));
  XOR2_X1    g09162(.A1(new_n4672_), .A2(new_n9243_), .Z(new_n9244_));
  NOR3_X1    g09163(.A1(new_n9240_), .A2(new_n9241_), .A3(new_n9244_), .ZN(new_n9245_));
  NAND2_X1   g09164(.A1(new_n8658_), .A2(new_n8855_), .ZN(new_n9246_));
  XNOR2_X1   g09165(.A1(new_n4672_), .A2(new_n9243_), .ZN(new_n9247_));
  AOI21_X1   g09166(.A1(new_n9246_), .A2(new_n9239_), .B(new_n9247_), .ZN(new_n9248_));
  NOR3_X1    g09167(.A1(new_n8668_), .A2(new_n8672_), .A3(new_n8399_), .ZN(new_n9249_));
  OR3_X2     g09168(.A1(new_n8658_), .A2(new_n8855_), .A3(new_n9249_), .Z(new_n9250_));
  OAI21_X1   g09169(.A1(new_n8658_), .A2(new_n9249_), .B(new_n8855_), .ZN(new_n9251_));
  NAND2_X1   g09170(.A1(new_n9250_), .A2(new_n9251_), .ZN(new_n9252_));
  INV_X1     g09171(.I(new_n9252_), .ZN(new_n9253_));
  AOI22_X1   g09172(.A1(new_n5935_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4029_), .ZN(new_n9254_));
  OAI21_X1   g09173(.A1(new_n9254_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9255_));
  XOR2_X1    g09174(.A1(new_n4687_), .A2(new_n9255_), .Z(new_n9256_));
  NAND2_X1   g09175(.A1(new_n9253_), .A2(new_n9256_), .ZN(new_n9257_));
  INV_X1     g09176(.I(new_n9256_), .ZN(new_n9258_));
  NAND2_X1   g09177(.A1(new_n9252_), .A2(new_n9258_), .ZN(new_n9259_));
  NOR2_X1    g09178(.A1(new_n9245_), .A2(new_n9248_), .ZN(new_n9261_));
  AOI21_X1   g09179(.A1(new_n9236_), .A2(new_n9238_), .B(new_n9261_), .ZN(new_n9262_));
  OAI21_X1   g09180(.A1(new_n8889_), .A2(new_n8887_), .B(new_n9262_), .ZN(new_n9263_));
  OAI21_X1   g09181(.A1(new_n8888_), .A2(new_n8885_), .B(new_n8857_), .ZN(new_n9264_));
  NAND3_X1   g09182(.A1(new_n8886_), .A2(new_n8672_), .A3(new_n8884_), .ZN(new_n9265_));
  NAND2_X1   g09183(.A1(new_n9265_), .A2(new_n9264_), .ZN(new_n9266_));
  NOR2_X1    g09184(.A1(new_n9266_), .A2(new_n9262_), .ZN(new_n9267_));
  NAND2_X1   g09185(.A1(new_n9252_), .A2(new_n9256_), .ZN(new_n9268_));
  OAI22_X1   g09186(.A1(new_n4028_), .A2(new_n8830_), .B1(new_n3042_), .B2(new_n4035_), .ZN(new_n9269_));
  OAI21_X1   g09187(.A1(new_n4017_), .A2(new_n3040_), .B(new_n9269_), .ZN(new_n9270_));
  AOI21_X1   g09188(.A1(new_n9270_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n9271_));
  XNOR2_X1   g09189(.A1(new_n4705_), .A2(new_n9271_), .ZN(new_n9272_));
  NOR2_X1    g09190(.A1(new_n9272_), .A2(new_n9268_), .ZN(new_n9273_));
  INV_X1     g09191(.I(new_n9273_), .ZN(new_n9274_));
  OAI21_X1   g09192(.A1(new_n9267_), .A2(new_n9274_), .B(new_n9263_), .ZN(new_n9275_));
  NAND3_X1   g09193(.A1(new_n8702_), .A2(new_n8701_), .A3(new_n8704_), .ZN(new_n9276_));
  NAND3_X1   g09194(.A1(new_n8848_), .A2(new_n9276_), .A3(new_n8692_), .ZN(new_n9277_));
  NAND3_X1   g09195(.A1(new_n9277_), .A2(new_n8862_), .A3(new_n8868_), .ZN(new_n9278_));
  NOR3_X1    g09196(.A1(new_n8700_), .A2(new_n8705_), .A3(new_n8864_), .ZN(new_n9279_));
  OAI21_X1   g09197(.A1(new_n9279_), .A2(new_n8865_), .B(new_n8867_), .ZN(new_n9280_));
  AOI22_X1   g09198(.A1(new_n4445_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4399_), .ZN(new_n9281_));
  OAI21_X1   g09199(.A1(new_n9281_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9282_));
  XOR2_X1    g09200(.A1(new_n4403_), .A2(new_n9282_), .Z(new_n9283_));
  NAND3_X1   g09201(.A1(new_n9280_), .A2(new_n9278_), .A3(new_n9283_), .ZN(new_n9284_));
  NOR3_X1    g09202(.A1(new_n9279_), .A2(new_n8867_), .A3(new_n8865_), .ZN(new_n9285_));
  AOI21_X1   g09203(.A1(new_n8868_), .A2(new_n9277_), .B(new_n8862_), .ZN(new_n9286_));
  XNOR2_X1   g09204(.A1(new_n4403_), .A2(new_n9282_), .ZN(new_n9287_));
  OAI21_X1   g09205(.A1(new_n9286_), .A2(new_n9285_), .B(new_n9287_), .ZN(new_n9288_));
  AOI21_X1   g09206(.A1(new_n9288_), .A2(new_n9284_), .B(new_n8877_), .ZN(new_n9289_));
  OAI21_X1   g09207(.A1(new_n9289_), .A2(new_n9275_), .B(new_n8883_), .ZN(new_n9290_));
  NOR2_X1    g09208(.A1(new_n9290_), .A2(new_n8852_), .ZN(new_n9291_));
  NOR3_X1    g09209(.A1(new_n9286_), .A2(new_n9285_), .A3(new_n9287_), .ZN(new_n9292_));
  NOR2_X1    g09210(.A1(new_n4397_), .A2(new_n8830_), .ZN(new_n9293_));
  NOR2_X1    g09211(.A1(new_n4374_), .A2(new_n3042_), .ZN(new_n9294_));
  OAI22_X1   g09212(.A1(new_n4437_), .A2(new_n3040_), .B1(new_n9293_), .B2(new_n9294_), .ZN(new_n9295_));
  AOI21_X1   g09213(.A1(new_n9295_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n9296_));
  INV_X1     g09214(.I(new_n9296_), .ZN(new_n9297_));
  NOR3_X1    g09215(.A1(new_n4538_), .A2(new_n4540_), .A3(new_n9297_), .ZN(new_n9298_));
  NOR2_X1    g09216(.A1(new_n4541_), .A2(new_n9296_), .ZN(new_n9299_));
  NOR2_X1    g09217(.A1(new_n9299_), .A2(new_n9298_), .ZN(new_n9300_));
  INV_X1     g09218(.I(new_n9300_), .ZN(new_n9301_));
  NAND2_X1   g09219(.A1(new_n9301_), .A2(new_n9292_), .ZN(new_n9302_));
  AOI21_X1   g09220(.A1(new_n9290_), .A2(new_n8852_), .B(new_n9302_), .ZN(new_n9303_));
  NOR2_X1    g09221(.A1(new_n9303_), .A2(new_n9291_), .ZN(new_n9304_));
  INV_X1     g09222(.I(new_n9304_), .ZN(new_n9305_));
  NAND3_X1   g09223(.A1(new_n8723_), .A2(new_n8725_), .A3(new_n8724_), .ZN(new_n9306_));
  OAI21_X1   g09224(.A1(new_n8718_), .A2(new_n8717_), .B(new_n8721_), .ZN(new_n9307_));
  NAND2_X1   g09225(.A1(new_n9306_), .A2(new_n9307_), .ZN(new_n9308_));
  NAND3_X1   g09226(.A1(new_n8736_), .A2(new_n8735_), .A3(new_n8737_), .ZN(new_n9309_));
  NAND3_X1   g09227(.A1(new_n8813_), .A2(new_n9309_), .A3(new_n9307_), .ZN(new_n9310_));
  NAND3_X1   g09228(.A1(new_n9310_), .A2(new_n8825_), .A3(new_n9308_), .ZN(new_n9311_));
  INV_X1     g09229(.I(new_n8825_), .ZN(new_n9312_));
  NOR3_X1    g09230(.A1(new_n8738_), .A2(new_n8734_), .A3(new_n8726_), .ZN(new_n9313_));
  OAI21_X1   g09231(.A1(new_n9313_), .A2(new_n8826_), .B(new_n9312_), .ZN(new_n9314_));
  INV_X1     g09232(.I(new_n4581_), .ZN(new_n9315_));
  AOI22_X1   g09233(.A1(new_n4473_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4555_), .ZN(new_n9316_));
  OAI21_X1   g09234(.A1(new_n9316_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9317_));
  INV_X1     g09235(.I(new_n9317_), .ZN(new_n9318_));
  NAND3_X1   g09236(.A1(new_n9315_), .A2(new_n4582_), .A3(new_n9318_), .ZN(new_n9319_));
  INV_X1     g09237(.I(new_n9319_), .ZN(new_n9320_));
  AOI21_X1   g09238(.A1(new_n9315_), .A2(new_n4582_), .B(new_n9318_), .ZN(new_n9321_));
  NOR2_X1    g09239(.A1(new_n9320_), .A2(new_n9321_), .ZN(new_n9322_));
  NAND3_X1   g09240(.A1(new_n9314_), .A2(new_n9322_), .A3(new_n9311_), .ZN(new_n9323_));
  NOR3_X1    g09241(.A1(new_n9313_), .A2(new_n9312_), .A3(new_n8826_), .ZN(new_n9324_));
  AOI21_X1   g09242(.A1(new_n9310_), .A2(new_n9308_), .B(new_n8825_), .ZN(new_n9325_));
  OAI21_X1   g09243(.A1(new_n4583_), .A2(new_n4581_), .B(new_n9317_), .ZN(new_n9326_));
  NAND2_X1   g09244(.A1(new_n9326_), .A2(new_n9319_), .ZN(new_n9327_));
  OAI21_X1   g09245(.A1(new_n9324_), .A2(new_n9325_), .B(new_n9327_), .ZN(new_n9328_));
  AOI21_X1   g09246(.A1(new_n9323_), .A2(new_n9328_), .B(new_n8836_), .ZN(new_n9329_));
  OAI21_X1   g09247(.A1(new_n9329_), .A2(new_n9305_), .B(new_n8840_), .ZN(new_n9330_));
  INV_X1     g09248(.I(new_n9330_), .ZN(new_n9331_));
  NAND2_X1   g09249(.A1(new_n9331_), .A2(new_n8824_), .ZN(new_n9332_));
  OAI22_X1   g09250(.A1(new_n3042_), .A2(new_n4468_), .B1(new_n4501_), .B2(new_n8830_), .ZN(new_n9333_));
  OAI21_X1   g09251(.A1(new_n4516_), .A2(new_n3040_), .B(new_n9333_), .ZN(new_n9334_));
  AOI21_X1   g09252(.A1(new_n9334_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n9335_));
  XOR2_X1    g09253(.A1(new_n4524_), .A2(new_n9335_), .Z(new_n9336_));
  NOR2_X1    g09254(.A1(new_n9323_), .A2(new_n9336_), .ZN(new_n9337_));
  OAI21_X1   g09255(.A1(new_n9331_), .A2(new_n8824_), .B(new_n9337_), .ZN(new_n9338_));
  NAND2_X1   g09256(.A1(new_n9338_), .A2(new_n9332_), .ZN(new_n9339_));
  INV_X1     g09257(.I(new_n9339_), .ZN(new_n9340_));
  AOI22_X1   g09258(.A1(new_n8760_), .A2(new_n8757_), .B1(new_n8742_), .B2(new_n8749_), .ZN(new_n9341_));
  INV_X1     g09259(.I(new_n8753_), .ZN(new_n9342_));
  NAND3_X1   g09260(.A1(new_n9342_), .A2(new_n8751_), .A3(new_n8756_), .ZN(new_n9343_));
  INV_X1     g09261(.I(new_n8756_), .ZN(new_n9344_));
  OAI21_X1   g09262(.A1(new_n8752_), .A2(new_n8753_), .B(new_n9344_), .ZN(new_n9345_));
  AOI21_X1   g09263(.A1(new_n9345_), .A2(new_n9343_), .B(new_n8750_), .ZN(new_n9346_));
  AOI22_X1   g09264(.A1(new_n5553_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4564_), .ZN(new_n9347_));
  OAI21_X1   g09265(.A1(new_n9347_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n9348_));
  XOR2_X1    g09266(.A1(new_n4569_), .A2(new_n9348_), .Z(new_n9349_));
  OAI21_X1   g09267(.A1(new_n9341_), .A2(new_n9346_), .B(new_n9349_), .ZN(new_n9350_));
  NAND2_X1   g09268(.A1(new_n8760_), .A2(new_n8757_), .ZN(new_n9351_));
  NAND2_X1   g09269(.A1(new_n9351_), .A2(new_n8750_), .ZN(new_n9352_));
  INV_X1     g09270(.I(new_n9346_), .ZN(new_n9353_));
  INV_X1     g09271(.I(new_n9349_), .ZN(new_n9354_));
  NAND3_X1   g09272(.A1(new_n9352_), .A2(new_n9353_), .A3(new_n9354_), .ZN(new_n9355_));
  AOI21_X1   g09273(.A1(new_n9355_), .A2(new_n9350_), .B(new_n9340_), .ZN(new_n9356_));
  NAND3_X1   g09274(.A1(new_n9352_), .A2(new_n9353_), .A3(new_n9349_), .ZN(new_n9357_));
  OAI21_X1   g09275(.A1(new_n9341_), .A2(new_n9346_), .B(new_n9354_), .ZN(new_n9358_));
  AOI21_X1   g09276(.A1(new_n9357_), .A2(new_n9358_), .B(new_n9339_), .ZN(new_n9359_));
  NOR2_X1    g09277(.A1(new_n9356_), .A2(new_n9359_), .ZN(new_n9360_));
  INV_X1     g09278(.I(new_n9360_), .ZN(new_n9361_));
  XNOR2_X1   g09279(.A1(new_n8840_), .A2(new_n9304_), .ZN(new_n9362_));
  OAI21_X1   g09280(.A1(new_n8897_), .A2(new_n8893_), .B(new_n8620_), .ZN(new_n9363_));
  NAND3_X1   g09281(.A1(new_n8894_), .A2(new_n8890_), .A3(new_n8895_), .ZN(new_n9364_));
  NAND2_X1   g09282(.A1(new_n9363_), .A2(new_n9364_), .ZN(new_n9365_));
  NAND2_X1   g09283(.A1(new_n9365_), .A2(new_n9187_), .ZN(new_n9366_));
  OAI21_X1   g09284(.A1(new_n9365_), .A2(new_n9187_), .B(new_n9195_), .ZN(new_n9367_));
  AOI21_X1   g09285(.A1(new_n9367_), .A2(new_n9366_), .B(new_n9208_), .ZN(new_n9368_));
  INV_X1     g09286(.I(new_n9211_), .ZN(new_n9369_));
  OAI21_X1   g09287(.A1(new_n9368_), .A2(new_n9369_), .B(new_n9220_), .ZN(new_n9370_));
  INV_X1     g09288(.I(new_n9223_), .ZN(new_n9371_));
  OAI21_X1   g09289(.A1(new_n9230_), .A2(new_n9227_), .B(new_n8645_), .ZN(new_n9372_));
  NAND3_X1   g09290(.A1(new_n9228_), .A2(new_n8646_), .A3(new_n9226_), .ZN(new_n9373_));
  INV_X1     g09291(.I(new_n9234_), .ZN(new_n9374_));
  AOI21_X1   g09292(.A1(new_n9372_), .A2(new_n9373_), .B(new_n9374_), .ZN(new_n9375_));
  AOI21_X1   g09293(.A1(new_n9370_), .A2(new_n9371_), .B(new_n9375_), .ZN(new_n9376_));
  OAI22_X1   g09294(.A1(new_n9376_), .A2(new_n9237_), .B1(new_n9245_), .B2(new_n9248_), .ZN(new_n9377_));
  AOI21_X1   g09295(.A1(new_n9264_), .A2(new_n9265_), .B(new_n9377_), .ZN(new_n9378_));
  NOR2_X1    g09296(.A1(new_n8887_), .A2(new_n8889_), .ZN(new_n9379_));
  NAND2_X1   g09297(.A1(new_n9379_), .A2(new_n9377_), .ZN(new_n9380_));
  AOI21_X1   g09298(.A1(new_n9380_), .A2(new_n9273_), .B(new_n9378_), .ZN(new_n9381_));
  XOR2_X1    g09299(.A1(new_n9381_), .A2(new_n8883_), .Z(new_n9382_));
  NAND3_X1   g09300(.A1(new_n9028_), .A2(new_n9029_), .A3(new_n9033_), .ZN(new_n9383_));
  INV_X1     g09301(.I(new_n9029_), .ZN(new_n9384_));
  OAI21_X1   g09302(.A1(new_n9384_), .A2(new_n9027_), .B(new_n9034_), .ZN(new_n9385_));
  NAND2_X1   g09303(.A1(new_n9383_), .A2(new_n9385_), .ZN(new_n9386_));
  OAI21_X1   g09304(.A1(new_n9384_), .A2(new_n9027_), .B(new_n9033_), .ZN(new_n9387_));
  AOI21_X1   g09305(.A1(new_n9036_), .A2(new_n9387_), .B(new_n9022_), .ZN(new_n9388_));
  AOI21_X1   g09306(.A1(new_n9022_), .A2(new_n9386_), .B(new_n9388_), .ZN(new_n9389_));
  NOR2_X1    g09307(.A1(new_n8954_), .A2(new_n8956_), .ZN(new_n9390_));
  NOR2_X1    g09308(.A1(new_n8959_), .A2(new_n8948_), .ZN(new_n9391_));
  OAI21_X1   g09309(.A1(new_n9391_), .A2(new_n9390_), .B(new_n8947_), .ZN(new_n9392_));
  AOI21_X1   g09310(.A1(new_n8944_), .A2(new_n8945_), .B(new_n8924_), .ZN(new_n9393_));
  NOR2_X1    g09311(.A1(new_n8954_), .A2(new_n8948_), .ZN(new_n9394_));
  OAI21_X1   g09312(.A1(new_n8960_), .A2(new_n9394_), .B(new_n9393_), .ZN(new_n9395_));
  NAND2_X1   g09313(.A1(new_n9392_), .A2(new_n9395_), .ZN(new_n9396_));
  INV_X1     g09314(.I(new_n8932_), .ZN(new_n9397_));
  NAND2_X1   g09315(.A1(new_n9397_), .A2(new_n8933_), .ZN(new_n9398_));
  NOR2_X1    g09316(.A1(new_n9398_), .A2(new_n8943_), .ZN(new_n9399_));
  INV_X1     g09317(.I(new_n8943_), .ZN(new_n9400_));
  NOR2_X1    g09318(.A1(new_n8935_), .A2(new_n9400_), .ZN(new_n9401_));
  NOR2_X1    g09319(.A1(new_n9401_), .A2(new_n9399_), .ZN(new_n9402_));
  INV_X1     g09320(.I(new_n8942_), .ZN(new_n9403_));
  NOR2_X1    g09321(.A1(new_n3416_), .A2(new_n451_), .ZN(new_n9404_));
  INV_X1     g09322(.I(new_n9404_), .ZN(new_n9405_));
  INV_X1     g09323(.I(\a[1] ), .ZN(new_n9406_));
  NOR2_X1    g09324(.A1(new_n9406_), .A2(\a[0] ), .ZN(new_n9407_));
  INV_X1     g09325(.I(new_n9407_), .ZN(new_n9408_));
  OAI22_X1   g09326(.A1(new_n4244_), .A2(new_n9405_), .B1(new_n4230_), .B2(new_n9408_), .ZN(new_n9409_));
  NAND2_X1   g09327(.A1(new_n9409_), .A2(\a[2] ), .ZN(new_n9410_));
  AOI21_X1   g09328(.A1(new_n9410_), .A2(new_n3456_), .B(new_n4234_), .ZN(new_n9411_));
  NOR2_X1    g09329(.A1(new_n4260_), .A2(new_n6061_), .ZN(new_n9412_));
  NOR2_X1    g09330(.A1(new_n5627_), .A2(new_n4234_), .ZN(new_n9413_));
  OAI21_X1   g09331(.A1(new_n9413_), .A2(new_n9412_), .B(new_n3413_), .ZN(new_n9414_));
  NAND2_X1   g09332(.A1(new_n5637_), .A2(new_n3413_), .ZN(new_n9415_));
  NOR2_X1    g09333(.A1(new_n3456_), .A2(new_n451_), .ZN(new_n9416_));
  NAND2_X1   g09334(.A1(new_n4252_), .A2(new_n9416_), .ZN(new_n9417_));
  OAI21_X1   g09335(.A1(new_n4230_), .A2(new_n451_), .B(new_n9406_), .ZN(new_n9418_));
  AND3_X2    g09336(.A1(new_n9418_), .A2(\a[0] ), .A3(new_n9417_), .Z(new_n9419_));
  NAND3_X1   g09337(.A1(new_n9414_), .A2(new_n9415_), .A3(new_n9419_), .ZN(new_n9420_));
  NOR3_X1    g09338(.A1(new_n9420_), .A2(new_n9403_), .A3(new_n9411_), .ZN(new_n9421_));
  INV_X1     g09339(.I(new_n9421_), .ZN(new_n9422_));
  OAI21_X1   g09340(.A1(new_n9420_), .A2(new_n9411_), .B(new_n9403_), .ZN(new_n9423_));
  NAND2_X1   g09341(.A1(new_n4221_), .A2(new_n3455_), .ZN(new_n9424_));
  NOR2_X1    g09342(.A1(new_n9405_), .A2(new_n9408_), .ZN(new_n9425_));
  AOI21_X1   g09343(.A1(new_n4260_), .A2(new_n4252_), .B(new_n9425_), .ZN(new_n9426_));
  AOI21_X1   g09344(.A1(new_n9426_), .A2(new_n9424_), .B(new_n3414_), .ZN(new_n9427_));
  AOI21_X1   g09345(.A1(new_n5648_), .A2(new_n9427_), .B(new_n451_), .ZN(new_n9428_));
  OAI21_X1   g09346(.A1(new_n6244_), .A2(new_n6243_), .B(new_n9427_), .ZN(new_n9429_));
  NOR2_X1    g09347(.A1(new_n9429_), .A2(\a[2] ), .ZN(new_n9430_));
  OAI21_X1   g09348(.A1(new_n9430_), .A2(new_n9428_), .B(new_n9423_), .ZN(new_n9431_));
  NAND2_X1   g09349(.A1(new_n9431_), .A2(new_n9422_), .ZN(new_n9432_));
  INV_X1     g09350(.I(new_n9425_), .ZN(new_n9433_));
  OAI21_X1   g09351(.A1(new_n4249_), .A2(new_n4234_), .B(new_n9433_), .ZN(new_n9434_));
  OAI21_X1   g09352(.A1(new_n4203_), .A2(new_n3456_), .B(new_n9434_), .ZN(new_n9435_));
  AOI21_X1   g09353(.A1(new_n9435_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n9436_));
  NAND3_X1   g09354(.A1(new_n5659_), .A2(new_n9436_), .A3(new_n5656_), .ZN(new_n9437_));
  INV_X1     g09355(.I(new_n9434_), .ZN(new_n9438_));
  AOI21_X1   g09356(.A1(new_n5653_), .A2(new_n5654_), .B(new_n3456_), .ZN(new_n9439_));
  OAI21_X1   g09357(.A1(new_n9439_), .A2(new_n9438_), .B(new_n451_), .ZN(new_n9440_));
  NAND2_X1   g09358(.A1(new_n9440_), .A2(new_n3411_), .ZN(new_n9441_));
  OAI21_X1   g09359(.A1(new_n6078_), .A2(new_n6081_), .B(new_n9441_), .ZN(new_n9442_));
  NAND2_X1   g09360(.A1(new_n9437_), .A2(new_n9442_), .ZN(new_n9443_));
  NAND2_X1   g09361(.A1(new_n9443_), .A2(new_n9432_), .ZN(new_n9444_));
  NOR2_X1    g09362(.A1(new_n8940_), .A2(new_n8941_), .ZN(new_n9445_));
  NOR2_X1    g09363(.A1(new_n8942_), .A2(new_n452_), .ZN(new_n9446_));
  NOR2_X1    g09364(.A1(new_n9445_), .A2(new_n9446_), .ZN(new_n9447_));
  NOR2_X1    g09365(.A1(new_n9447_), .A2(new_n8943_), .ZN(new_n9448_));
  INV_X1     g09366(.I(new_n9448_), .ZN(new_n9449_));
  OAI21_X1   g09367(.A1(new_n9443_), .A2(new_n9432_), .B(new_n9449_), .ZN(new_n9450_));
  AOI21_X1   g09368(.A1(new_n9450_), .A2(new_n9444_), .B(new_n9402_), .ZN(new_n9451_));
  NAND3_X1   g09369(.A1(new_n9450_), .A2(new_n9444_), .A3(new_n9402_), .ZN(new_n9452_));
  NAND2_X1   g09370(.A1(new_n4258_), .A2(new_n3455_), .ZN(new_n9453_));
  NOR2_X1    g09371(.A1(new_n6542_), .A2(new_n9425_), .ZN(new_n9454_));
  AOI21_X1   g09372(.A1(new_n9454_), .A2(new_n9453_), .B(new_n3414_), .ZN(new_n9455_));
  INV_X1     g09373(.I(new_n9455_), .ZN(new_n9456_));
  OAI21_X1   g09374(.A1(new_n9456_), .A2(new_n6540_), .B(\a[2] ), .ZN(new_n9457_));
  NAND3_X1   g09375(.A1(new_n5671_), .A2(new_n451_), .A3(new_n9455_), .ZN(new_n9458_));
  NAND2_X1   g09376(.A1(new_n9457_), .A2(new_n9458_), .ZN(new_n9459_));
  AOI21_X1   g09377(.A1(new_n9452_), .A2(new_n9459_), .B(new_n9451_), .ZN(new_n9460_));
  OAI22_X1   g09378(.A1(new_n5684_), .A2(new_n3456_), .B1(new_n6556_), .B2(new_n9425_), .ZN(new_n9461_));
  AOI21_X1   g09379(.A1(new_n9461_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n9462_));
  INV_X1     g09380(.I(new_n9462_), .ZN(new_n9463_));
  NOR3_X1    g09381(.A1(new_n6100_), .A2(new_n6101_), .A3(new_n9463_), .ZN(new_n9464_));
  AOI21_X1   g09382(.A1(new_n5692_), .A2(new_n5688_), .B(new_n9462_), .ZN(new_n9465_));
  NOR2_X1    g09383(.A1(new_n9464_), .A2(new_n9465_), .ZN(new_n9466_));
  NOR2_X1    g09384(.A1(new_n9460_), .A2(new_n9466_), .ZN(new_n9467_));
  AOI21_X1   g09385(.A1(new_n8935_), .A2(new_n8943_), .B(new_n8490_), .ZN(new_n9468_));
  NAND3_X1   g09386(.A1(new_n8935_), .A2(new_n8490_), .A3(new_n8943_), .ZN(new_n9469_));
  INV_X1     g09387(.I(new_n9469_), .ZN(new_n9470_));
  NOR3_X1    g09388(.A1(new_n9470_), .A2(new_n9468_), .A3(new_n8923_), .ZN(new_n9471_));
  INV_X1     g09389(.I(new_n8923_), .ZN(new_n9472_));
  INV_X1     g09390(.I(new_n9468_), .ZN(new_n9473_));
  AOI21_X1   g09391(.A1(new_n9473_), .A2(new_n9469_), .B(new_n9472_), .ZN(new_n9474_));
  NOR2_X1    g09392(.A1(new_n9474_), .A2(new_n9471_), .ZN(new_n9475_));
  AOI21_X1   g09393(.A1(new_n9460_), .A2(new_n9466_), .B(new_n9475_), .ZN(new_n9476_));
  OAI21_X1   g09394(.A1(new_n9476_), .A2(new_n9467_), .B(new_n9396_), .ZN(new_n9477_));
  NOR3_X1    g09395(.A1(new_n9476_), .A2(new_n9467_), .A3(new_n9396_), .ZN(new_n9478_));
  NAND2_X1   g09396(.A1(new_n5701_), .A2(new_n3455_), .ZN(new_n9479_));
  NOR2_X1    g09397(.A1(new_n6567_), .A2(new_n9425_), .ZN(new_n9480_));
  AOI21_X1   g09398(.A1(new_n9479_), .A2(new_n9480_), .B(new_n3414_), .ZN(new_n9481_));
  INV_X1     g09399(.I(new_n9481_), .ZN(new_n9482_));
  NOR2_X1    g09400(.A1(new_n5707_), .A2(new_n9482_), .ZN(new_n9483_));
  XOR2_X1    g09401(.A1(new_n9483_), .A2(new_n451_), .Z(new_n9484_));
  OAI21_X1   g09402(.A1(new_n9478_), .A2(new_n9484_), .B(new_n9477_), .ZN(new_n9485_));
  NAND2_X1   g09403(.A1(new_n8967_), .A2(new_n8963_), .ZN(new_n9486_));
  OR2_X2     g09404(.A1(new_n8967_), .A2(new_n8963_), .Z(new_n9487_));
  AOI22_X1   g09405(.A1(new_n9487_), .A2(new_n9486_), .B1(new_n8955_), .B2(new_n8961_), .ZN(new_n9488_));
  INV_X1     g09406(.I(new_n8969_), .ZN(new_n9489_));
  AOI21_X1   g09407(.A1(new_n8968_), .A2(new_n9489_), .B(new_n8962_), .ZN(new_n9490_));
  NOR2_X1    g09408(.A1(new_n9490_), .A2(new_n9488_), .ZN(new_n9491_));
  INV_X1     g09409(.I(new_n9491_), .ZN(new_n9492_));
  NAND2_X1   g09410(.A1(new_n9485_), .A2(new_n9492_), .ZN(new_n9493_));
  NOR3_X1    g09411(.A1(new_n5720_), .A2(new_n3414_), .A3(new_n5715_), .ZN(new_n9494_));
  AOI22_X1   g09412(.A1(new_n6582_), .A2(new_n9433_), .B1(new_n4274_), .B2(new_n3455_), .ZN(new_n9495_));
  INV_X1     g09413(.I(new_n9495_), .ZN(new_n9496_));
  NOR3_X1    g09414(.A1(new_n9494_), .A2(new_n451_), .A3(new_n9496_), .ZN(new_n9497_));
  INV_X1     g09415(.I(new_n9497_), .ZN(new_n9498_));
  OAI21_X1   g09416(.A1(new_n9494_), .A2(new_n9496_), .B(new_n451_), .ZN(new_n9499_));
  NAND2_X1   g09417(.A1(new_n9498_), .A2(new_n9499_), .ZN(new_n9500_));
  OAI21_X1   g09418(.A1(new_n9485_), .A2(new_n9492_), .B(new_n9500_), .ZN(new_n9501_));
  NAND2_X1   g09419(.A1(new_n8979_), .A2(new_n8975_), .ZN(new_n9502_));
  NAND2_X1   g09420(.A1(new_n8976_), .A2(new_n8982_), .ZN(new_n9503_));
  AOI21_X1   g09421(.A1(new_n9503_), .A2(new_n9502_), .B(new_n8970_), .ZN(new_n9504_));
  NAND2_X1   g09422(.A1(new_n8980_), .A2(new_n8983_), .ZN(new_n9505_));
  AOI21_X1   g09423(.A1(new_n8970_), .A2(new_n9505_), .B(new_n9504_), .ZN(new_n9506_));
  AOI21_X1   g09424(.A1(new_n9501_), .A2(new_n9493_), .B(new_n9506_), .ZN(new_n9507_));
  AND2_X2    g09425(.A1(new_n9392_), .A2(new_n9395_), .Z(new_n9508_));
  NAND2_X1   g09426(.A1(new_n8935_), .A2(new_n9400_), .ZN(new_n9509_));
  NAND2_X1   g09427(.A1(new_n9398_), .A2(new_n8943_), .ZN(new_n9510_));
  NAND2_X1   g09428(.A1(new_n9509_), .A2(new_n9510_), .ZN(new_n9511_));
  NAND2_X1   g09429(.A1(new_n9429_), .A2(\a[2] ), .ZN(new_n9512_));
  NAND3_X1   g09430(.A1(new_n5648_), .A2(new_n451_), .A3(new_n9427_), .ZN(new_n9513_));
  NAND2_X1   g09431(.A1(new_n9512_), .A2(new_n9513_), .ZN(new_n9514_));
  AOI21_X1   g09432(.A1(new_n9514_), .A2(new_n9423_), .B(new_n9421_), .ZN(new_n9515_));
  NOR3_X1    g09433(.A1(new_n6078_), .A2(new_n6081_), .A3(new_n9441_), .ZN(new_n9516_));
  AOI21_X1   g09434(.A1(new_n5656_), .A2(new_n5659_), .B(new_n9436_), .ZN(new_n9517_));
  NOR2_X1    g09435(.A1(new_n9517_), .A2(new_n9516_), .ZN(new_n9518_));
  NOR2_X1    g09436(.A1(new_n9518_), .A2(new_n9515_), .ZN(new_n9519_));
  AOI21_X1   g09437(.A1(new_n9518_), .A2(new_n9515_), .B(new_n9448_), .ZN(new_n9520_));
  OAI21_X1   g09438(.A1(new_n9520_), .A2(new_n9519_), .B(new_n9511_), .ZN(new_n9521_));
  NOR3_X1    g09439(.A1(new_n9520_), .A2(new_n9519_), .A3(new_n9511_), .ZN(new_n9522_));
  AOI21_X1   g09440(.A1(new_n5671_), .A2(new_n9455_), .B(new_n451_), .ZN(new_n9523_));
  NOR3_X1    g09441(.A1(new_n9456_), .A2(new_n6540_), .A3(\a[2] ), .ZN(new_n9524_));
  NOR2_X1    g09442(.A1(new_n9524_), .A2(new_n9523_), .ZN(new_n9525_));
  OAI21_X1   g09443(.A1(new_n9522_), .A2(new_n9525_), .B(new_n9521_), .ZN(new_n9526_));
  NAND3_X1   g09444(.A1(new_n5692_), .A2(new_n5688_), .A3(new_n9462_), .ZN(new_n9527_));
  OAI21_X1   g09445(.A1(new_n6100_), .A2(new_n6101_), .B(new_n9463_), .ZN(new_n9528_));
  NAND2_X1   g09446(.A1(new_n9528_), .A2(new_n9527_), .ZN(new_n9529_));
  NAND2_X1   g09447(.A1(new_n9526_), .A2(new_n9529_), .ZN(new_n9530_));
  OR2_X2     g09448(.A1(new_n9474_), .A2(new_n9471_), .Z(new_n9531_));
  OAI21_X1   g09449(.A1(new_n9526_), .A2(new_n9529_), .B(new_n9531_), .ZN(new_n9532_));
  NAND3_X1   g09450(.A1(new_n9532_), .A2(new_n9508_), .A3(new_n9530_), .ZN(new_n9533_));
  OAI21_X1   g09451(.A1(new_n5707_), .A2(new_n9482_), .B(\a[2] ), .ZN(new_n9534_));
  NAND2_X1   g09452(.A1(new_n9483_), .A2(new_n451_), .ZN(new_n9535_));
  NAND2_X1   g09453(.A1(new_n9535_), .A2(new_n9534_), .ZN(new_n9536_));
  NAND2_X1   g09454(.A1(new_n9533_), .A2(new_n9536_), .ZN(new_n9537_));
  AOI21_X1   g09455(.A1(new_n9537_), .A2(new_n9477_), .B(new_n9491_), .ZN(new_n9538_));
  NAND3_X1   g09456(.A1(new_n9537_), .A2(new_n9477_), .A3(new_n9491_), .ZN(new_n9539_));
  AOI21_X1   g09457(.A1(new_n9539_), .A2(new_n9500_), .B(new_n9538_), .ZN(new_n9540_));
  NOR2_X1    g09458(.A1(new_n5733_), .A2(new_n3414_), .ZN(new_n9541_));
  AOI22_X1   g09459(.A1(new_n4143_), .A2(new_n3455_), .B1(new_n4278_), .B2(new_n9433_), .ZN(new_n9542_));
  INV_X1     g09460(.I(new_n9542_), .ZN(new_n9543_));
  NOR3_X1    g09461(.A1(new_n9541_), .A2(new_n451_), .A3(new_n9543_), .ZN(new_n9544_));
  NAND2_X1   g09462(.A1(new_n6134_), .A2(new_n3411_), .ZN(new_n9545_));
  AOI21_X1   g09463(.A1(new_n9545_), .A2(new_n9542_), .B(\a[2] ), .ZN(new_n9546_));
  NOR2_X1    g09464(.A1(new_n9546_), .A2(new_n9544_), .ZN(new_n9547_));
  AOI21_X1   g09465(.A1(new_n9540_), .A2(new_n9506_), .B(new_n9547_), .ZN(new_n9548_));
  NAND2_X1   g09466(.A1(new_n6609_), .A2(new_n9433_), .ZN(new_n9549_));
  OAI21_X1   g09467(.A1(new_n4135_), .A2(new_n3456_), .B(new_n9549_), .ZN(new_n9550_));
  AOI21_X1   g09468(.A1(new_n9550_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n9551_));
  INV_X1     g09469(.I(new_n9551_), .ZN(new_n9552_));
  NOR3_X1    g09470(.A1(new_n5618_), .A2(new_n5622_), .A3(new_n9552_), .ZN(new_n9553_));
  AOI21_X1   g09471(.A1(new_n5619_), .A2(new_n5623_), .B(new_n9551_), .ZN(new_n9554_));
  NOR2_X1    g09472(.A1(new_n9554_), .A2(new_n9553_), .ZN(new_n9555_));
  INV_X1     g09473(.I(new_n9555_), .ZN(new_n9556_));
  OAI21_X1   g09474(.A1(new_n9548_), .A2(new_n9507_), .B(new_n9556_), .ZN(new_n9557_));
  AOI21_X1   g09475(.A1(new_n9532_), .A2(new_n9530_), .B(new_n9508_), .ZN(new_n9558_));
  AOI21_X1   g09476(.A1(new_n9533_), .A2(new_n9536_), .B(new_n9558_), .ZN(new_n9559_));
  INV_X1     g09477(.I(new_n9499_), .ZN(new_n9560_));
  NOR2_X1    g09478(.A1(new_n9560_), .A2(new_n9497_), .ZN(new_n9561_));
  AOI21_X1   g09479(.A1(new_n9559_), .A2(new_n9491_), .B(new_n9561_), .ZN(new_n9562_));
  INV_X1     g09480(.I(new_n9504_), .ZN(new_n9563_));
  NAND2_X1   g09481(.A1(new_n9505_), .A2(new_n8970_), .ZN(new_n9564_));
  NAND2_X1   g09482(.A1(new_n9563_), .A2(new_n9564_), .ZN(new_n9565_));
  OAI21_X1   g09483(.A1(new_n9562_), .A2(new_n9538_), .B(new_n9565_), .ZN(new_n9566_));
  NAND3_X1   g09484(.A1(new_n9501_), .A2(new_n9493_), .A3(new_n9506_), .ZN(new_n9567_));
  INV_X1     g09485(.I(new_n9547_), .ZN(new_n9568_));
  NAND2_X1   g09486(.A1(new_n9567_), .A2(new_n9568_), .ZN(new_n9569_));
  NAND3_X1   g09487(.A1(new_n9569_), .A2(new_n9566_), .A3(new_n9555_), .ZN(new_n9570_));
  XNOR2_X1   g09488(.A1(new_n8984_), .A2(new_n8998_), .ZN(new_n9571_));
  INV_X1     g09489(.I(new_n9571_), .ZN(new_n9572_));
  NAND2_X1   g09490(.A1(new_n9570_), .A2(new_n9572_), .ZN(new_n9573_));
  INV_X1     g09491(.I(new_n8997_), .ZN(new_n9574_));
  NOR2_X1    g09492(.A1(new_n9003_), .A2(new_n8914_), .ZN(new_n9575_));
  OAI21_X1   g09493(.A1(new_n8998_), .A2(new_n8984_), .B(new_n9575_), .ZN(new_n9576_));
  XNOR2_X1   g09494(.A1(new_n5722_), .A2(new_n9002_), .ZN(new_n9577_));
  NAND2_X1   g09495(.A1(new_n9577_), .A2(new_n8915_), .ZN(new_n9578_));
  NAND2_X1   g09496(.A1(new_n8999_), .A2(new_n9578_), .ZN(new_n9579_));
  AOI21_X1   g09497(.A1(new_n9579_), .A2(new_n9576_), .B(new_n9574_), .ZN(new_n9580_));
  NOR2_X1    g09498(.A1(new_n8999_), .A2(new_n9578_), .ZN(new_n9581_));
  NOR3_X1    g09499(.A1(new_n9575_), .A2(new_n8984_), .A3(new_n8998_), .ZN(new_n9582_));
  NOR3_X1    g09500(.A1(new_n9581_), .A2(new_n8997_), .A3(new_n9582_), .ZN(new_n9583_));
  NOR2_X1    g09501(.A1(new_n9583_), .A2(new_n9580_), .ZN(new_n9584_));
  AOI21_X1   g09502(.A1(new_n9573_), .A2(new_n9557_), .B(new_n9584_), .ZN(new_n9585_));
  AOI21_X1   g09503(.A1(new_n9569_), .A2(new_n9566_), .B(new_n9555_), .ZN(new_n9586_));
  AOI21_X1   g09504(.A1(new_n9570_), .A2(new_n9572_), .B(new_n9586_), .ZN(new_n9587_));
  NAND2_X1   g09505(.A1(new_n4290_), .A2(new_n3455_), .ZN(new_n9588_));
  NOR2_X1    g09506(.A1(new_n6621_), .A2(new_n9425_), .ZN(new_n9589_));
  AOI21_X1   g09507(.A1(new_n9588_), .A2(new_n9589_), .B(new_n3414_), .ZN(new_n9590_));
  NAND2_X1   g09508(.A1(new_n5023_), .A2(new_n9590_), .ZN(new_n9591_));
  XOR2_X1    g09509(.A1(new_n9591_), .A2(\a[2] ), .Z(new_n9592_));
  AOI21_X1   g09510(.A1(new_n9587_), .A2(new_n9584_), .B(new_n9592_), .ZN(new_n9593_));
  XOR2_X1    g09511(.A1(new_n9013_), .A2(new_n9020_), .Z(new_n9594_));
  NAND2_X1   g09512(.A1(new_n9006_), .A2(new_n9594_), .ZN(new_n9595_));
  AND2_X2    g09513(.A1(new_n9018_), .A2(new_n9021_), .Z(new_n9596_));
  OAI21_X1   g09514(.A1(new_n9006_), .A2(new_n9596_), .B(new_n9595_), .ZN(new_n9597_));
  OAI21_X1   g09515(.A1(new_n9593_), .A2(new_n9585_), .B(new_n9597_), .ZN(new_n9598_));
  AOI21_X1   g09516(.A1(new_n9567_), .A2(new_n9568_), .B(new_n9507_), .ZN(new_n9599_));
  AOI21_X1   g09517(.A1(new_n9599_), .A2(new_n9555_), .B(new_n9571_), .ZN(new_n9600_));
  OAI21_X1   g09518(.A1(new_n9581_), .A2(new_n9582_), .B(new_n8997_), .ZN(new_n9601_));
  NAND3_X1   g09519(.A1(new_n9579_), .A2(new_n9576_), .A3(new_n9574_), .ZN(new_n9602_));
  NAND2_X1   g09520(.A1(new_n9601_), .A2(new_n9602_), .ZN(new_n9603_));
  OAI21_X1   g09521(.A1(new_n9600_), .A2(new_n9586_), .B(new_n9603_), .ZN(new_n9604_));
  NOR3_X1    g09522(.A1(new_n9600_), .A2(new_n9603_), .A3(new_n9586_), .ZN(new_n9605_));
  OAI21_X1   g09523(.A1(new_n9605_), .A2(new_n9592_), .B(new_n9604_), .ZN(new_n9606_));
  NAND2_X1   g09524(.A1(new_n4297_), .A2(new_n3455_), .ZN(new_n9607_));
  NOR2_X1    g09525(.A1(new_n6627_), .A2(new_n9425_), .ZN(new_n9608_));
  AOI21_X1   g09526(.A1(new_n9607_), .A2(new_n9608_), .B(new_n3414_), .ZN(new_n9609_));
  NAND2_X1   g09527(.A1(new_n5753_), .A2(new_n9609_), .ZN(new_n9610_));
  XOR2_X1    g09528(.A1(new_n9610_), .A2(\a[2] ), .Z(new_n9611_));
  INV_X1     g09529(.I(new_n9611_), .ZN(new_n9612_));
  OAI21_X1   g09530(.A1(new_n9606_), .A2(new_n9597_), .B(new_n9612_), .ZN(new_n9613_));
  AOI21_X1   g09531(.A1(new_n9613_), .A2(new_n9598_), .B(new_n9389_), .ZN(new_n9614_));
  NOR3_X1    g09532(.A1(new_n9548_), .A2(new_n9507_), .A3(new_n9556_), .ZN(new_n9615_));
  OAI21_X1   g09533(.A1(new_n9615_), .A2(new_n9571_), .B(new_n9557_), .ZN(new_n9616_));
  XOR2_X1    g09534(.A1(new_n9591_), .A2(new_n451_), .Z(new_n9617_));
  OAI21_X1   g09535(.A1(new_n9616_), .A2(new_n9603_), .B(new_n9617_), .ZN(new_n9618_));
  NOR2_X1    g09536(.A1(new_n9596_), .A2(new_n9006_), .ZN(new_n9619_));
  AOI21_X1   g09537(.A1(new_n9006_), .A2(new_n9594_), .B(new_n9619_), .ZN(new_n9620_));
  AOI21_X1   g09538(.A1(new_n9618_), .A2(new_n9604_), .B(new_n9620_), .ZN(new_n9621_));
  NAND3_X1   g09539(.A1(new_n9618_), .A2(new_n9604_), .A3(new_n9620_), .ZN(new_n9622_));
  AOI21_X1   g09540(.A1(new_n9622_), .A2(new_n9612_), .B(new_n9621_), .ZN(new_n9623_));
  NAND2_X1   g09541(.A1(new_n5042_), .A2(new_n3455_), .ZN(new_n9624_));
  NOR2_X1    g09542(.A1(new_n4301_), .A2(new_n9425_), .ZN(new_n9625_));
  AOI21_X1   g09543(.A1(new_n9624_), .A2(new_n9625_), .B(new_n3414_), .ZN(new_n9626_));
  AOI21_X1   g09544(.A1(new_n5599_), .A2(new_n9626_), .B(new_n451_), .ZN(new_n9627_));
  AND3_X2    g09545(.A1(new_n5599_), .A2(new_n451_), .A3(new_n9626_), .Z(new_n9628_));
  NOR2_X1    g09546(.A1(new_n9628_), .A2(new_n9627_), .ZN(new_n9629_));
  AOI21_X1   g09547(.A1(new_n9623_), .A2(new_n9389_), .B(new_n9629_), .ZN(new_n9630_));
  AOI22_X1   g09548(.A1(new_n6980_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n5041_), .ZN(new_n9631_));
  OAI21_X1   g09549(.A1(new_n9631_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n9632_));
  NOR2_X1    g09550(.A1(new_n5049_), .A2(new_n9632_), .ZN(new_n9633_));
  AND2_X2    g09551(.A1(new_n5049_), .A2(new_n9632_), .Z(new_n9634_));
  NOR2_X1    g09552(.A1(new_n9634_), .A2(new_n9633_), .ZN(new_n9635_));
  INV_X1     g09553(.I(new_n9635_), .ZN(new_n9636_));
  OAI21_X1   g09554(.A1(new_n9630_), .A2(new_n9614_), .B(new_n9636_), .ZN(new_n9637_));
  NAND2_X1   g09555(.A1(new_n9036_), .A2(new_n9387_), .ZN(new_n9638_));
  MUX2_X1    g09556(.I0(new_n9638_), .I1(new_n9386_), .S(new_n9022_), .Z(new_n9639_));
  NAND3_X1   g09557(.A1(new_n9573_), .A2(new_n9557_), .A3(new_n9584_), .ZN(new_n9640_));
  AOI21_X1   g09558(.A1(new_n9640_), .A2(new_n9617_), .B(new_n9585_), .ZN(new_n9641_));
  AOI21_X1   g09559(.A1(new_n9641_), .A2(new_n9620_), .B(new_n9611_), .ZN(new_n9642_));
  OAI21_X1   g09560(.A1(new_n9642_), .A2(new_n9621_), .B(new_n9639_), .ZN(new_n9643_));
  NOR3_X1    g09561(.A1(new_n9593_), .A2(new_n9585_), .A3(new_n9597_), .ZN(new_n9644_));
  OAI21_X1   g09562(.A1(new_n9644_), .A2(new_n9611_), .B(new_n9598_), .ZN(new_n9645_));
  INV_X1     g09563(.I(new_n9629_), .ZN(new_n9646_));
  OAI21_X1   g09564(.A1(new_n9645_), .A2(new_n9639_), .B(new_n9646_), .ZN(new_n9647_));
  NAND3_X1   g09565(.A1(new_n9647_), .A2(new_n9643_), .A3(new_n9635_), .ZN(new_n9648_));
  AOI21_X1   g09566(.A1(new_n9049_), .A2(new_n9050_), .B(new_n9042_), .ZN(new_n9649_));
  OAI21_X1   g09567(.A1(new_n9649_), .A2(new_n9057_), .B(new_n9038_), .ZN(new_n9650_));
  NAND3_X1   g09568(.A1(new_n9051_), .A2(new_n9054_), .A3(new_n9037_), .ZN(new_n9651_));
  NAND2_X1   g09569(.A1(new_n9650_), .A2(new_n9651_), .ZN(new_n9652_));
  NAND2_X1   g09570(.A1(new_n9648_), .A2(new_n9652_), .ZN(new_n9653_));
  AOI22_X1   g09571(.A1(new_n6993_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n4124_), .ZN(new_n9654_));
  OAI21_X1   g09572(.A1(new_n9654_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n9655_));
  NOR2_X1    g09573(.A1(new_n5067_), .A2(new_n9655_), .ZN(new_n9656_));
  INV_X1     g09574(.I(new_n9655_), .ZN(new_n9657_));
  NOR2_X1    g09575(.A1(new_n5906_), .A2(new_n9657_), .ZN(new_n9658_));
  NOR2_X1    g09576(.A1(new_n9658_), .A2(new_n9656_), .ZN(new_n9659_));
  AOI21_X1   g09577(.A1(new_n9653_), .A2(new_n9637_), .B(new_n9659_), .ZN(new_n9660_));
  AOI21_X1   g09578(.A1(new_n9647_), .A2(new_n9643_), .B(new_n9635_), .ZN(new_n9661_));
  AOI21_X1   g09579(.A1(new_n9648_), .A2(new_n9652_), .B(new_n9661_), .ZN(new_n9662_));
  NAND3_X1   g09580(.A1(new_n9061_), .A2(new_n8909_), .A3(new_n9059_), .ZN(new_n9663_));
  AOI21_X1   g09581(.A1(new_n9061_), .A2(new_n9059_), .B(new_n8909_), .ZN(new_n9664_));
  INV_X1     g09582(.I(new_n9664_), .ZN(new_n9665_));
  AOI22_X1   g09583(.A1(new_n9055_), .A2(new_n9051_), .B1(new_n9663_), .B2(new_n9665_), .ZN(new_n9666_));
  OAI21_X1   g09584(.A1(new_n9037_), .A2(new_n9649_), .B(new_n9051_), .ZN(new_n9667_));
  NAND2_X1   g09585(.A1(new_n9665_), .A2(new_n9663_), .ZN(new_n9668_));
  NOR2_X1    g09586(.A1(new_n9668_), .A2(new_n9667_), .ZN(new_n9669_));
  NOR2_X1    g09587(.A1(new_n9669_), .A2(new_n9666_), .ZN(new_n9670_));
  AOI21_X1   g09588(.A1(new_n9662_), .A2(new_n9659_), .B(new_n9670_), .ZN(new_n9671_));
  NAND3_X1   g09589(.A1(new_n9076_), .A2(new_n9075_), .A3(new_n9072_), .ZN(new_n9672_));
  OAI21_X1   g09590(.A1(new_n9066_), .A2(new_n9069_), .B(new_n9077_), .ZN(new_n9673_));
  NAND2_X1   g09591(.A1(new_n9672_), .A2(new_n9673_), .ZN(new_n9674_));
  OAI21_X1   g09592(.A1(new_n9056_), .A2(new_n9064_), .B(new_n9674_), .ZN(new_n9675_));
  INV_X1     g09593(.I(new_n9056_), .ZN(new_n9676_));
  INV_X1     g09594(.I(new_n9064_), .ZN(new_n9677_));
  NAND2_X1   g09595(.A1(new_n9078_), .A2(new_n9073_), .ZN(new_n9678_));
  NAND3_X1   g09596(.A1(new_n9677_), .A2(new_n9678_), .A3(new_n9676_), .ZN(new_n9679_));
  NAND2_X1   g09597(.A1(new_n9675_), .A2(new_n9679_), .ZN(new_n9680_));
  OAI21_X1   g09598(.A1(new_n9671_), .A2(new_n9660_), .B(new_n9680_), .ZN(new_n9681_));
  NAND3_X1   g09599(.A1(new_n9613_), .A2(new_n9389_), .A3(new_n9598_), .ZN(new_n9682_));
  AOI21_X1   g09600(.A1(new_n9682_), .A2(new_n9646_), .B(new_n9614_), .ZN(new_n9683_));
  AOI21_X1   g09601(.A1(new_n9051_), .A2(new_n9054_), .B(new_n9037_), .ZN(new_n9684_));
  NOR3_X1    g09602(.A1(new_n9649_), .A2(new_n9057_), .A3(new_n9038_), .ZN(new_n9685_));
  NOR2_X1    g09603(.A1(new_n9684_), .A2(new_n9685_), .ZN(new_n9686_));
  AOI21_X1   g09604(.A1(new_n9683_), .A2(new_n9635_), .B(new_n9686_), .ZN(new_n9687_));
  INV_X1     g09605(.I(new_n9659_), .ZN(new_n9688_));
  OAI21_X1   g09606(.A1(new_n9687_), .A2(new_n9661_), .B(new_n9688_), .ZN(new_n9689_));
  NOR3_X1    g09607(.A1(new_n9687_), .A2(new_n9661_), .A3(new_n9688_), .ZN(new_n9690_));
  OAI21_X1   g09608(.A1(new_n9690_), .A2(new_n9670_), .B(new_n9689_), .ZN(new_n9691_));
  NOR2_X1    g09609(.A1(new_n5096_), .A2(new_n3414_), .ZN(new_n9692_));
  OAI22_X1   g09610(.A1(new_n4112_), .A2(new_n3456_), .B1(new_n6682_), .B2(new_n9425_), .ZN(new_n9693_));
  OR3_X2     g09611(.A1(new_n9692_), .A2(new_n451_), .A3(new_n9693_), .Z(new_n9694_));
  OAI21_X1   g09612(.A1(new_n9692_), .A2(new_n9693_), .B(new_n451_), .ZN(new_n9695_));
  NAND2_X1   g09613(.A1(new_n9694_), .A2(new_n9695_), .ZN(new_n9696_));
  OAI21_X1   g09614(.A1(new_n9691_), .A2(new_n9680_), .B(new_n9696_), .ZN(new_n9697_));
  NAND2_X1   g09615(.A1(new_n4105_), .A2(new_n3455_), .ZN(new_n9698_));
  NOR2_X1    g09616(.A1(new_n6692_), .A2(new_n9425_), .ZN(new_n9699_));
  AOI21_X1   g09617(.A1(new_n9699_), .A2(new_n9698_), .B(new_n3414_), .ZN(new_n9700_));
  AOI21_X1   g09618(.A1(new_n5121_), .A2(new_n9700_), .B(new_n451_), .ZN(new_n9701_));
  AND3_X2    g09619(.A1(new_n5121_), .A2(new_n451_), .A3(new_n9700_), .Z(new_n9702_));
  NOR2_X1    g09620(.A1(new_n9702_), .A2(new_n9701_), .ZN(new_n9703_));
  AOI21_X1   g09621(.A1(new_n9697_), .A2(new_n9681_), .B(new_n9703_), .ZN(new_n9704_));
  NOR3_X1    g09622(.A1(new_n9630_), .A2(new_n9614_), .A3(new_n9636_), .ZN(new_n9705_));
  OAI21_X1   g09623(.A1(new_n9705_), .A2(new_n9686_), .B(new_n9637_), .ZN(new_n9706_));
  INV_X1     g09624(.I(new_n9670_), .ZN(new_n9707_));
  OAI21_X1   g09625(.A1(new_n9706_), .A2(new_n9688_), .B(new_n9707_), .ZN(new_n9708_));
  NAND2_X1   g09626(.A1(new_n9677_), .A2(new_n9676_), .ZN(new_n9709_));
  AOI21_X1   g09627(.A1(new_n9076_), .A2(new_n9075_), .B(new_n9077_), .ZN(new_n9710_));
  NOR3_X1    g09628(.A1(new_n9066_), .A2(new_n9069_), .A3(new_n9072_), .ZN(new_n9711_));
  NOR2_X1    g09629(.A1(new_n9710_), .A2(new_n9711_), .ZN(new_n9712_));
  NOR3_X1    g09630(.A1(new_n9712_), .A2(new_n9056_), .A3(new_n9064_), .ZN(new_n9713_));
  AOI21_X1   g09631(.A1(new_n9709_), .A2(new_n9674_), .B(new_n9713_), .ZN(new_n9714_));
  AOI21_X1   g09632(.A1(new_n9708_), .A2(new_n9689_), .B(new_n9714_), .ZN(new_n9715_));
  NAND3_X1   g09633(.A1(new_n9708_), .A2(new_n9714_), .A3(new_n9689_), .ZN(new_n9716_));
  AOI21_X1   g09634(.A1(new_n9716_), .A2(new_n9696_), .B(new_n9715_), .ZN(new_n9717_));
  NOR2_X1    g09635(.A1(new_n9086_), .A2(new_n9088_), .ZN(new_n9718_));
  XOR2_X1    g09636(.A1(new_n9718_), .A2(new_n9079_), .Z(new_n9719_));
  AOI21_X1   g09637(.A1(new_n9717_), .A2(new_n9703_), .B(new_n9719_), .ZN(new_n9720_));
  INV_X1     g09638(.I(new_n9079_), .ZN(new_n9721_));
  INV_X1     g09639(.I(new_n9718_), .ZN(new_n9722_));
  INV_X1     g09640(.I(new_n9088_), .ZN(new_n9723_));
  NAND3_X1   g09641(.A1(new_n9101_), .A2(new_n9094_), .A3(new_n9102_), .ZN(new_n9724_));
  OAI21_X1   g09642(.A1(new_n9095_), .A2(new_n9096_), .B(new_n9099_), .ZN(new_n9725_));
  NAND3_X1   g09643(.A1(new_n9725_), .A2(new_n9724_), .A3(new_n9723_), .ZN(new_n9726_));
  NAND3_X1   g09644(.A1(new_n9726_), .A2(new_n9721_), .A3(new_n9722_), .ZN(new_n9727_));
  NOR3_X1    g09645(.A1(new_n9103_), .A2(new_n9100_), .A3(new_n9088_), .ZN(new_n9728_));
  OAI21_X1   g09646(.A1(new_n9728_), .A2(new_n9718_), .B(new_n9079_), .ZN(new_n9729_));
  NAND2_X1   g09647(.A1(new_n9729_), .A2(new_n9727_), .ZN(new_n9730_));
  OAI21_X1   g09648(.A1(new_n9720_), .A2(new_n9704_), .B(new_n9730_), .ZN(new_n9731_));
  NAND3_X1   g09649(.A1(new_n9653_), .A2(new_n9637_), .A3(new_n9659_), .ZN(new_n9732_));
  AOI21_X1   g09650(.A1(new_n9732_), .A2(new_n9707_), .B(new_n9660_), .ZN(new_n9733_));
  INV_X1     g09651(.I(new_n9696_), .ZN(new_n9734_));
  AOI21_X1   g09652(.A1(new_n9733_), .A2(new_n9714_), .B(new_n9734_), .ZN(new_n9735_));
  INV_X1     g09653(.I(new_n9703_), .ZN(new_n9736_));
  OAI21_X1   g09654(.A1(new_n9735_), .A2(new_n9715_), .B(new_n9736_), .ZN(new_n9737_));
  NOR3_X1    g09655(.A1(new_n9671_), .A2(new_n9660_), .A3(new_n9680_), .ZN(new_n9738_));
  OAI21_X1   g09656(.A1(new_n9738_), .A2(new_n9734_), .B(new_n9681_), .ZN(new_n9739_));
  XNOR2_X1   g09657(.A1(new_n9718_), .A2(new_n9079_), .ZN(new_n9740_));
  OAI21_X1   g09658(.A1(new_n9739_), .A2(new_n9736_), .B(new_n9740_), .ZN(new_n9741_));
  NOR3_X1    g09659(.A1(new_n9728_), .A2(new_n9079_), .A3(new_n9718_), .ZN(new_n9742_));
  AOI21_X1   g09660(.A1(new_n9726_), .A2(new_n9722_), .B(new_n9721_), .ZN(new_n9743_));
  NOR2_X1    g09661(.A1(new_n9742_), .A2(new_n9743_), .ZN(new_n9744_));
  NAND3_X1   g09662(.A1(new_n9741_), .A2(new_n9744_), .A3(new_n9737_), .ZN(new_n9745_));
  NAND2_X1   g09663(.A1(new_n4100_), .A2(new_n3455_), .ZN(new_n9746_));
  NOR2_X1    g09664(.A1(new_n6704_), .A2(new_n9425_), .ZN(new_n9747_));
  AOI21_X1   g09665(.A1(new_n9747_), .A2(new_n9746_), .B(new_n3414_), .ZN(new_n9748_));
  NAND2_X1   g09666(.A1(new_n5080_), .A2(new_n9748_), .ZN(new_n9749_));
  XOR2_X1    g09667(.A1(new_n9749_), .A2(\a[2] ), .Z(new_n9750_));
  INV_X1     g09668(.I(new_n9750_), .ZN(new_n9751_));
  NAND2_X1   g09669(.A1(new_n9745_), .A2(new_n9751_), .ZN(new_n9752_));
  OAI21_X1   g09670(.A1(new_n8905_), .A2(new_n8902_), .B(new_n9111_), .ZN(new_n9753_));
  INV_X1     g09671(.I(new_n9753_), .ZN(new_n9754_));
  NAND2_X1   g09672(.A1(new_n9754_), .A2(new_n9105_), .ZN(new_n9755_));
  NAND3_X1   g09673(.A1(new_n9753_), .A2(new_n9079_), .A3(new_n9104_), .ZN(new_n9756_));
  AOI21_X1   g09674(.A1(new_n9755_), .A2(new_n9756_), .B(new_n9103_), .ZN(new_n9757_));
  NAND3_X1   g09675(.A1(new_n9755_), .A2(new_n9756_), .A3(new_n9103_), .ZN(new_n9758_));
  INV_X1     g09676(.I(new_n9758_), .ZN(new_n9759_));
  NOR2_X1    g09677(.A1(new_n9759_), .A2(new_n9757_), .ZN(new_n9760_));
  AOI21_X1   g09678(.A1(new_n9752_), .A2(new_n9731_), .B(new_n9760_), .ZN(new_n9761_));
  AOI21_X1   g09679(.A1(new_n9741_), .A2(new_n9737_), .B(new_n9744_), .ZN(new_n9762_));
  AOI21_X1   g09680(.A1(new_n9745_), .A2(new_n9751_), .B(new_n9762_), .ZN(new_n9763_));
  NAND2_X1   g09681(.A1(new_n4091_), .A2(new_n3455_), .ZN(new_n9764_));
  NOR2_X1    g09682(.A1(new_n4320_), .A2(new_n9425_), .ZN(new_n9765_));
  AOI21_X1   g09683(.A1(new_n9764_), .A2(new_n9765_), .B(new_n3414_), .ZN(new_n9766_));
  NAND2_X1   g09684(.A1(new_n5197_), .A2(new_n9766_), .ZN(new_n9767_));
  XOR2_X1    g09685(.A1(new_n9767_), .A2(\a[2] ), .Z(new_n9768_));
  AOI21_X1   g09686(.A1(new_n9763_), .A2(new_n9760_), .B(new_n9768_), .ZN(new_n9769_));
  AOI22_X1   g09687(.A1(new_n6419_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n4328_), .ZN(new_n9770_));
  OAI21_X1   g09688(.A1(new_n9770_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n9771_));
  XNOR2_X1   g09689(.A1(new_n5139_), .A2(new_n9771_), .ZN(new_n9772_));
  INV_X1     g09690(.I(new_n9772_), .ZN(new_n9773_));
  OAI21_X1   g09691(.A1(new_n9769_), .A2(new_n9761_), .B(new_n9773_), .ZN(new_n9774_));
  NAND3_X1   g09692(.A1(new_n9697_), .A2(new_n9681_), .A3(new_n9703_), .ZN(new_n9775_));
  AOI21_X1   g09693(.A1(new_n9775_), .A2(new_n9740_), .B(new_n9704_), .ZN(new_n9776_));
  AOI21_X1   g09694(.A1(new_n9776_), .A2(new_n9744_), .B(new_n9750_), .ZN(new_n9777_));
  INV_X1     g09695(.I(new_n9757_), .ZN(new_n9778_));
  NAND2_X1   g09696(.A1(new_n9778_), .A2(new_n9758_), .ZN(new_n9779_));
  OAI21_X1   g09697(.A1(new_n9777_), .A2(new_n9762_), .B(new_n9779_), .ZN(new_n9780_));
  NOR3_X1    g09698(.A1(new_n9777_), .A2(new_n9779_), .A3(new_n9762_), .ZN(new_n9781_));
  OAI21_X1   g09699(.A1(new_n9781_), .A2(new_n9768_), .B(new_n9780_), .ZN(new_n9782_));
  NOR3_X1    g09700(.A1(new_n9130_), .A2(new_n9134_), .A3(new_n9114_), .ZN(new_n9783_));
  INV_X1     g09701(.I(new_n9114_), .ZN(new_n9784_));
  NAND3_X1   g09702(.A1(new_n9132_), .A2(new_n9133_), .A3(new_n9128_), .ZN(new_n9785_));
  OAI21_X1   g09703(.A1(new_n9125_), .A2(new_n9122_), .B(new_n9129_), .ZN(new_n9786_));
  AOI21_X1   g09704(.A1(new_n9786_), .A2(new_n9785_), .B(new_n9784_), .ZN(new_n9787_));
  OR2_X2     g09705(.A1(new_n9783_), .A2(new_n9787_), .Z(new_n9788_));
  OAI21_X1   g09706(.A1(new_n9782_), .A2(new_n9773_), .B(new_n9788_), .ZN(new_n9789_));
  AOI22_X1   g09707(.A1(new_n4333_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n4082_), .ZN(new_n9790_));
  OAI21_X1   g09708(.A1(new_n9790_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n9791_));
  XNOR2_X1   g09709(.A1(new_n5162_), .A2(new_n9791_), .ZN(new_n9792_));
  AOI21_X1   g09710(.A1(new_n9789_), .A2(new_n9774_), .B(new_n9792_), .ZN(new_n9793_));
  NOR3_X1    g09711(.A1(new_n9720_), .A2(new_n9704_), .A3(new_n9730_), .ZN(new_n9794_));
  OAI21_X1   g09712(.A1(new_n9794_), .A2(new_n9750_), .B(new_n9731_), .ZN(new_n9795_));
  INV_X1     g09713(.I(new_n9768_), .ZN(new_n9796_));
  OAI21_X1   g09714(.A1(new_n9795_), .A2(new_n9779_), .B(new_n9796_), .ZN(new_n9797_));
  AOI21_X1   g09715(.A1(new_n9797_), .A2(new_n9780_), .B(new_n9772_), .ZN(new_n9798_));
  NAND3_X1   g09716(.A1(new_n9797_), .A2(new_n9780_), .A3(new_n9772_), .ZN(new_n9799_));
  AOI21_X1   g09717(.A1(new_n9799_), .A2(new_n9788_), .B(new_n9798_), .ZN(new_n9800_));
  NOR2_X1    g09718(.A1(new_n9131_), .A2(new_n9134_), .ZN(new_n9801_));
  NAND2_X1   g09719(.A1(new_n9142_), .A2(new_n9144_), .ZN(new_n9802_));
  NOR2_X1    g09720(.A1(new_n9801_), .A2(new_n9802_), .ZN(new_n9803_));
  INV_X1     g09721(.I(new_n9802_), .ZN(new_n9804_));
  NOR3_X1    g09722(.A1(new_n9804_), .A2(new_n9131_), .A3(new_n9134_), .ZN(new_n9805_));
  NOR2_X1    g09723(.A1(new_n9805_), .A2(new_n9803_), .ZN(new_n9806_));
  AOI21_X1   g09724(.A1(new_n9800_), .A2(new_n9792_), .B(new_n9806_), .ZN(new_n9807_));
  NAND3_X1   g09725(.A1(new_n9158_), .A2(new_n9152_), .A3(new_n9156_), .ZN(new_n9808_));
  OAI21_X1   g09726(.A1(new_n9153_), .A2(new_n9151_), .B(new_n9159_), .ZN(new_n9809_));
  AOI22_X1   g09727(.A1(new_n9808_), .A2(new_n9809_), .B1(new_n9143_), .B2(new_n9144_), .ZN(new_n9810_));
  AOI21_X1   g09728(.A1(new_n9157_), .A2(new_n9160_), .B(new_n9145_), .ZN(new_n9811_));
  NOR2_X1    g09729(.A1(new_n9811_), .A2(new_n9810_), .ZN(new_n9812_));
  INV_X1     g09730(.I(new_n9812_), .ZN(new_n9813_));
  OAI21_X1   g09731(.A1(new_n9807_), .A2(new_n9793_), .B(new_n9813_), .ZN(new_n9814_));
  NAND3_X1   g09732(.A1(new_n9752_), .A2(new_n9760_), .A3(new_n9731_), .ZN(new_n9815_));
  AOI21_X1   g09733(.A1(new_n9815_), .A2(new_n9796_), .B(new_n9761_), .ZN(new_n9816_));
  NOR2_X1    g09734(.A1(new_n9783_), .A2(new_n9787_), .ZN(new_n9817_));
  AOI21_X1   g09735(.A1(new_n9816_), .A2(new_n9772_), .B(new_n9817_), .ZN(new_n9818_));
  INV_X1     g09736(.I(new_n9792_), .ZN(new_n9819_));
  OAI21_X1   g09737(.A1(new_n9818_), .A2(new_n9798_), .B(new_n9819_), .ZN(new_n9820_));
  NOR3_X1    g09738(.A1(new_n9769_), .A2(new_n9761_), .A3(new_n9773_), .ZN(new_n9821_));
  OAI21_X1   g09739(.A1(new_n9821_), .A2(new_n9817_), .B(new_n9774_), .ZN(new_n9822_));
  INV_X1     g09740(.I(new_n9806_), .ZN(new_n9823_));
  OAI21_X1   g09741(.A1(new_n9822_), .A2(new_n9819_), .B(new_n9823_), .ZN(new_n9824_));
  NAND3_X1   g09742(.A1(new_n9824_), .A2(new_n9820_), .A3(new_n9812_), .ZN(new_n9825_));
  NAND2_X1   g09743(.A1(new_n4071_), .A2(new_n3455_), .ZN(new_n9826_));
  NOR2_X1    g09744(.A1(new_n5917_), .A2(new_n9425_), .ZN(new_n9827_));
  AOI21_X1   g09745(.A1(new_n9826_), .A2(new_n9827_), .B(new_n3414_), .ZN(new_n9828_));
  NAND2_X1   g09746(.A1(new_n4928_), .A2(new_n9828_), .ZN(new_n9829_));
  XOR2_X1    g09747(.A1(new_n9829_), .A2(\a[2] ), .Z(new_n9830_));
  INV_X1     g09748(.I(new_n9830_), .ZN(new_n9831_));
  NAND2_X1   g09749(.A1(new_n9825_), .A2(new_n9831_), .ZN(new_n9832_));
  NAND2_X1   g09750(.A1(new_n4061_), .A2(new_n3455_), .ZN(new_n9833_));
  NOR2_X1    g09751(.A1(new_n4336_), .A2(new_n9425_), .ZN(new_n9834_));
  AOI21_X1   g09752(.A1(new_n9834_), .A2(new_n9833_), .B(new_n3414_), .ZN(new_n9835_));
  NAND2_X1   g09753(.A1(new_n4935_), .A2(new_n9835_), .ZN(new_n9836_));
  XOR2_X1    g09754(.A1(new_n9836_), .A2(\a[2] ), .Z(new_n9837_));
  AOI21_X1   g09755(.A1(new_n9832_), .A2(new_n9814_), .B(new_n9837_), .ZN(new_n9838_));
  AOI21_X1   g09756(.A1(new_n9824_), .A2(new_n9820_), .B(new_n9812_), .ZN(new_n9839_));
  AOI21_X1   g09757(.A1(new_n9825_), .A2(new_n9831_), .B(new_n9839_), .ZN(new_n9840_));
  NOR2_X1    g09758(.A1(new_n9174_), .A2(new_n9172_), .ZN(new_n9841_));
  XNOR2_X1   g09759(.A1(new_n9162_), .A2(new_n9841_), .ZN(new_n9842_));
  AOI21_X1   g09760(.A1(new_n9840_), .A2(new_n9837_), .B(new_n9842_), .ZN(new_n9843_));
  INV_X1     g09761(.I(new_n9841_), .ZN(new_n9844_));
  NOR2_X1    g09762(.A1(new_n9184_), .A2(new_n9174_), .ZN(new_n9845_));
  INV_X1     g09763(.I(new_n9845_), .ZN(new_n9846_));
  AND3_X2    g09764(.A1(new_n9846_), .A2(new_n9162_), .A3(new_n9844_), .Z(new_n9847_));
  AOI21_X1   g09765(.A1(new_n9846_), .A2(new_n9844_), .B(new_n9162_), .ZN(new_n9848_));
  NOR2_X1    g09766(.A1(new_n9847_), .A2(new_n9848_), .ZN(new_n9849_));
  INV_X1     g09767(.I(new_n9849_), .ZN(new_n9850_));
  OAI21_X1   g09768(.A1(new_n9843_), .A2(new_n9838_), .B(new_n9850_), .ZN(new_n9851_));
  NAND3_X1   g09769(.A1(new_n9789_), .A2(new_n9774_), .A3(new_n9792_), .ZN(new_n9852_));
  AOI21_X1   g09770(.A1(new_n9852_), .A2(new_n9823_), .B(new_n9793_), .ZN(new_n9853_));
  AOI21_X1   g09771(.A1(new_n9853_), .A2(new_n9812_), .B(new_n9830_), .ZN(new_n9854_));
  INV_X1     g09772(.I(new_n9837_), .ZN(new_n9855_));
  OAI21_X1   g09773(.A1(new_n9854_), .A2(new_n9839_), .B(new_n9855_), .ZN(new_n9856_));
  NOR3_X1    g09774(.A1(new_n9854_), .A2(new_n9839_), .A3(new_n9855_), .ZN(new_n9857_));
  OAI21_X1   g09775(.A1(new_n9857_), .A2(new_n9842_), .B(new_n9856_), .ZN(new_n9858_));
  NAND2_X1   g09776(.A1(new_n4054_), .A2(new_n3455_), .ZN(new_n9859_));
  NOR2_X1    g09777(.A1(new_n4339_), .A2(new_n9425_), .ZN(new_n9860_));
  AOI21_X1   g09778(.A1(new_n9860_), .A2(new_n9859_), .B(new_n3414_), .ZN(new_n9861_));
  NAND2_X1   g09779(.A1(new_n4652_), .A2(new_n9861_), .ZN(new_n9862_));
  XOR2_X1    g09780(.A1(new_n9862_), .A2(\a[2] ), .Z(new_n9863_));
  INV_X1     g09781(.I(new_n9863_), .ZN(new_n9864_));
  OAI21_X1   g09782(.A1(new_n9858_), .A2(new_n9850_), .B(new_n9864_), .ZN(new_n9865_));
  INV_X1     g09783(.I(new_n9194_), .ZN(new_n9866_));
  NAND2_X1   g09784(.A1(new_n9365_), .A2(new_n9866_), .ZN(new_n9867_));
  XOR2_X1    g09785(.A1(new_n9867_), .A2(new_n9188_), .Z(new_n9868_));
  XOR2_X1    g09786(.A1(new_n9868_), .A2(new_n9191_), .Z(new_n9869_));
  AOI21_X1   g09787(.A1(new_n9865_), .A2(new_n9851_), .B(new_n9869_), .ZN(new_n9870_));
  NOR3_X1    g09788(.A1(new_n9807_), .A2(new_n9813_), .A3(new_n9793_), .ZN(new_n9871_));
  OAI21_X1   g09789(.A1(new_n9871_), .A2(new_n9830_), .B(new_n9814_), .ZN(new_n9872_));
  INV_X1     g09790(.I(new_n9842_), .ZN(new_n9873_));
  OAI21_X1   g09791(.A1(new_n9872_), .A2(new_n9855_), .B(new_n9873_), .ZN(new_n9874_));
  AOI21_X1   g09792(.A1(new_n9874_), .A2(new_n9856_), .B(new_n9849_), .ZN(new_n9875_));
  NAND3_X1   g09793(.A1(new_n9874_), .A2(new_n9856_), .A3(new_n9849_), .ZN(new_n9876_));
  AOI21_X1   g09794(.A1(new_n9876_), .A2(new_n9864_), .B(new_n9875_), .ZN(new_n9877_));
  NAND2_X1   g09795(.A1(new_n4043_), .A2(new_n3455_), .ZN(new_n9878_));
  NOR2_X1    g09796(.A1(new_n4342_), .A2(new_n9425_), .ZN(new_n9879_));
  AOI21_X1   g09797(.A1(new_n9878_), .A2(new_n9879_), .B(new_n3414_), .ZN(new_n9880_));
  NAND2_X1   g09798(.A1(new_n4864_), .A2(new_n9880_), .ZN(new_n9881_));
  XOR2_X1    g09799(.A1(new_n9881_), .A2(\a[2] ), .Z(new_n9882_));
  AOI21_X1   g09800(.A1(new_n9877_), .A2(new_n9869_), .B(new_n9882_), .ZN(new_n9883_));
  AOI22_X1   g09801(.A1(new_n4347_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n4036_), .ZN(new_n9884_));
  OAI21_X1   g09802(.A1(new_n9884_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n9885_));
  XOR2_X1    g09803(.A1(new_n4672_), .A2(new_n9885_), .Z(new_n9886_));
  INV_X1     g09804(.I(new_n9886_), .ZN(new_n9887_));
  OAI21_X1   g09805(.A1(new_n9883_), .A2(new_n9870_), .B(new_n9887_), .ZN(new_n9888_));
  NAND3_X1   g09806(.A1(new_n9832_), .A2(new_n9814_), .A3(new_n9837_), .ZN(new_n9889_));
  AOI21_X1   g09807(.A1(new_n9889_), .A2(new_n9873_), .B(new_n9838_), .ZN(new_n9890_));
  AOI21_X1   g09808(.A1(new_n9890_), .A2(new_n9849_), .B(new_n9863_), .ZN(new_n9891_));
  XNOR2_X1   g09809(.A1(new_n9868_), .A2(new_n9191_), .ZN(new_n9892_));
  OAI21_X1   g09810(.A1(new_n9891_), .A2(new_n9875_), .B(new_n9892_), .ZN(new_n9893_));
  NOR3_X1    g09811(.A1(new_n9843_), .A2(new_n9838_), .A3(new_n9850_), .ZN(new_n9894_));
  OAI21_X1   g09812(.A1(new_n9894_), .A2(new_n9863_), .B(new_n9851_), .ZN(new_n9895_));
  INV_X1     g09813(.I(new_n9882_), .ZN(new_n9896_));
  OAI21_X1   g09814(.A1(new_n9895_), .A2(new_n9892_), .B(new_n9896_), .ZN(new_n9897_));
  NAND3_X1   g09815(.A1(new_n9897_), .A2(new_n9893_), .A3(new_n9886_), .ZN(new_n9898_));
  NAND2_X1   g09816(.A1(new_n9367_), .A2(new_n9366_), .ZN(new_n9899_));
  NAND2_X1   g09817(.A1(new_n9209_), .A2(new_n9211_), .ZN(new_n9900_));
  XNOR2_X1   g09818(.A1(new_n9900_), .A2(new_n9899_), .ZN(new_n9901_));
  INV_X1     g09819(.I(new_n9901_), .ZN(new_n9902_));
  NAND2_X1   g09820(.A1(new_n9898_), .A2(new_n9902_), .ZN(new_n9903_));
  AOI22_X1   g09821(.A1(new_n5935_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n4029_), .ZN(new_n9904_));
  OAI21_X1   g09822(.A1(new_n9904_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n9905_));
  XOR2_X1    g09823(.A1(new_n4687_), .A2(new_n9905_), .Z(new_n9906_));
  AOI21_X1   g09824(.A1(new_n9903_), .A2(new_n9888_), .B(new_n9906_), .ZN(new_n9907_));
  AOI21_X1   g09825(.A1(new_n9897_), .A2(new_n9893_), .B(new_n9886_), .ZN(new_n9908_));
  AOI21_X1   g09826(.A1(new_n9898_), .A2(new_n9902_), .B(new_n9908_), .ZN(new_n9909_));
  NOR2_X1    g09827(.A1(new_n9368_), .A2(new_n9369_), .ZN(new_n9910_));
  NOR2_X1    g09828(.A1(new_n9221_), .A2(new_n9223_), .ZN(new_n9911_));
  XNOR2_X1   g09829(.A1(new_n9911_), .A2(new_n9910_), .ZN(new_n9912_));
  AOI21_X1   g09830(.A1(new_n9909_), .A2(new_n9906_), .B(new_n9912_), .ZN(new_n9913_));
  OAI22_X1   g09831(.A1(new_n4028_), .A2(new_n9405_), .B1(new_n4035_), .B2(new_n9408_), .ZN(new_n9914_));
  OAI21_X1   g09832(.A1(new_n4017_), .A2(new_n3456_), .B(new_n9914_), .ZN(new_n9915_));
  AOI21_X1   g09833(.A1(new_n9915_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n9916_));
  XNOR2_X1   g09834(.A1(new_n4705_), .A2(new_n9916_), .ZN(new_n9917_));
  INV_X1     g09835(.I(new_n9917_), .ZN(new_n9918_));
  OAI21_X1   g09836(.A1(new_n9913_), .A2(new_n9907_), .B(new_n9918_), .ZN(new_n9919_));
  NAND3_X1   g09837(.A1(new_n9865_), .A2(new_n9869_), .A3(new_n9851_), .ZN(new_n9920_));
  AOI21_X1   g09838(.A1(new_n9920_), .A2(new_n9896_), .B(new_n9870_), .ZN(new_n9921_));
  AOI21_X1   g09839(.A1(new_n9921_), .A2(new_n9886_), .B(new_n9901_), .ZN(new_n9922_));
  INV_X1     g09840(.I(new_n9906_), .ZN(new_n9923_));
  OAI21_X1   g09841(.A1(new_n9922_), .A2(new_n9908_), .B(new_n9923_), .ZN(new_n9924_));
  NOR3_X1    g09842(.A1(new_n9922_), .A2(new_n9908_), .A3(new_n9923_), .ZN(new_n9925_));
  OAI21_X1   g09843(.A1(new_n9925_), .A2(new_n9912_), .B(new_n9924_), .ZN(new_n9926_));
  NAND2_X1   g09844(.A1(new_n9370_), .A2(new_n9371_), .ZN(new_n9927_));
  NOR2_X1    g09845(.A1(new_n9375_), .A2(new_n9237_), .ZN(new_n9928_));
  XOR2_X1    g09846(.A1(new_n9928_), .A2(new_n9927_), .Z(new_n9929_));
  INV_X1     g09847(.I(new_n9929_), .ZN(new_n9930_));
  OAI21_X1   g09848(.A1(new_n9926_), .A2(new_n9918_), .B(new_n9930_), .ZN(new_n9931_));
  NAND2_X1   g09849(.A1(new_n4375_), .A2(new_n3455_), .ZN(new_n9932_));
  NOR2_X1    g09850(.A1(new_n4355_), .A2(new_n9425_), .ZN(new_n9933_));
  AOI21_X1   g09851(.A1(new_n9933_), .A2(new_n9932_), .B(new_n3414_), .ZN(new_n9934_));
  NAND2_X1   g09852(.A1(new_n4730_), .A2(new_n9934_), .ZN(new_n9935_));
  XOR2_X1    g09853(.A1(new_n9935_), .A2(\a[2] ), .Z(new_n9936_));
  AOI21_X1   g09854(.A1(new_n9931_), .A2(new_n9919_), .B(new_n9936_), .ZN(new_n9937_));
  NOR3_X1    g09855(.A1(new_n9883_), .A2(new_n9870_), .A3(new_n9887_), .ZN(new_n9938_));
  OAI21_X1   g09856(.A1(new_n9938_), .A2(new_n9901_), .B(new_n9888_), .ZN(new_n9939_));
  INV_X1     g09857(.I(new_n9912_), .ZN(new_n9940_));
  OAI21_X1   g09858(.A1(new_n9939_), .A2(new_n9923_), .B(new_n9940_), .ZN(new_n9941_));
  AOI21_X1   g09859(.A1(new_n9941_), .A2(new_n9924_), .B(new_n9917_), .ZN(new_n9942_));
  NAND3_X1   g09860(.A1(new_n9941_), .A2(new_n9924_), .A3(new_n9917_), .ZN(new_n9943_));
  AOI21_X1   g09861(.A1(new_n9943_), .A2(new_n9930_), .B(new_n9942_), .ZN(new_n9944_));
  NOR2_X1    g09862(.A1(new_n9376_), .A2(new_n9237_), .ZN(new_n9945_));
  NAND3_X1   g09863(.A1(new_n9246_), .A2(new_n9247_), .A3(new_n9239_), .ZN(new_n9946_));
  OAI21_X1   g09864(.A1(new_n9240_), .A2(new_n9241_), .B(new_n9244_), .ZN(new_n9947_));
  NAND2_X1   g09865(.A1(new_n9947_), .A2(new_n9946_), .ZN(new_n9948_));
  XOR2_X1    g09866(.A1(new_n9945_), .A2(new_n9948_), .Z(new_n9949_));
  AOI21_X1   g09867(.A1(new_n9944_), .A2(new_n9936_), .B(new_n9949_), .ZN(new_n9950_));
  NAND3_X1   g09868(.A1(new_n9257_), .A2(new_n9947_), .A3(new_n9259_), .ZN(new_n9951_));
  AND3_X2    g09869(.A1(new_n9951_), .A2(new_n9945_), .A3(new_n9948_), .Z(new_n9952_));
  AOI21_X1   g09870(.A1(new_n9951_), .A2(new_n9948_), .B(new_n9945_), .ZN(new_n9953_));
  NOR2_X1    g09871(.A1(new_n9952_), .A2(new_n9953_), .ZN(new_n9954_));
  INV_X1     g09872(.I(new_n9954_), .ZN(new_n9955_));
  NOR3_X1    g09873(.A1(new_n9379_), .A2(new_n9262_), .A3(new_n9272_), .ZN(new_n9956_));
  NOR2_X1    g09874(.A1(new_n9379_), .A2(new_n9272_), .ZN(new_n9957_));
  NOR2_X1    g09875(.A1(new_n9957_), .A2(new_n9377_), .ZN(new_n9958_));
  OAI21_X1   g09876(.A1(new_n9958_), .A2(new_n9956_), .B(new_n9268_), .ZN(new_n9959_));
  INV_X1     g09877(.I(new_n9959_), .ZN(new_n9960_));
  NOR3_X1    g09878(.A1(new_n9958_), .A2(new_n9956_), .A3(new_n9268_), .ZN(new_n9961_));
  OAI22_X1   g09879(.A1(new_n4397_), .A2(new_n9405_), .B1(new_n4374_), .B2(new_n9408_), .ZN(new_n9962_));
  OAI21_X1   g09880(.A1(new_n4437_), .A2(new_n3456_), .B(new_n9962_), .ZN(new_n9963_));
  AOI21_X1   g09881(.A1(new_n9963_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n9964_));
  XOR2_X1    g09882(.A1(new_n4541_), .A2(new_n9964_), .Z(new_n9965_));
  NOR3_X1    g09883(.A1(new_n9960_), .A2(new_n9961_), .A3(new_n9965_), .ZN(new_n9966_));
  INV_X1     g09884(.I(new_n9961_), .ZN(new_n9967_));
  INV_X1     g09885(.I(new_n9965_), .ZN(new_n9968_));
  AOI21_X1   g09886(.A1(new_n9967_), .A2(new_n9959_), .B(new_n9968_), .ZN(new_n9969_));
  NOR3_X1    g09887(.A1(new_n9969_), .A2(new_n9966_), .A3(new_n9955_), .ZN(new_n9970_));
  OAI22_X1   g09888(.A1(new_n4444_), .A2(new_n9425_), .B1(new_n3456_), .B2(new_n4397_), .ZN(new_n9971_));
  AOI21_X1   g09889(.A1(new_n9971_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n9972_));
  XNOR2_X1   g09890(.A1(new_n4403_), .A2(new_n9972_), .ZN(new_n9973_));
  OAI21_X1   g09891(.A1(new_n9969_), .A2(new_n9966_), .B(new_n9955_), .ZN(new_n9974_));
  AOI21_X1   g09892(.A1(new_n9973_), .A2(new_n9974_), .B(new_n9970_), .ZN(new_n9975_));
  OAI21_X1   g09893(.A1(new_n9950_), .A2(new_n9937_), .B(new_n9975_), .ZN(new_n9976_));
  NOR2_X1    g09894(.A1(new_n9976_), .A2(new_n9382_), .ZN(new_n9977_));
  OAI21_X1   g09895(.A1(new_n9960_), .A2(new_n9961_), .B(new_n9965_), .ZN(new_n9978_));
  AOI22_X1   g09896(.A1(new_n4448_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n4469_), .ZN(new_n9979_));
  OAI21_X1   g09897(.A1(new_n9979_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n9980_));
  XNOR2_X1   g09898(.A1(new_n4477_), .A2(new_n9980_), .ZN(new_n9981_));
  NOR2_X1    g09899(.A1(new_n9978_), .A2(new_n9981_), .ZN(new_n9982_));
  INV_X1     g09900(.I(new_n9982_), .ZN(new_n9983_));
  AOI21_X1   g09901(.A1(new_n9976_), .A2(new_n9382_), .B(new_n9983_), .ZN(new_n9984_));
  NOR2_X1    g09902(.A1(new_n9984_), .A2(new_n9977_), .ZN(new_n9985_));
  NOR3_X1    g09903(.A1(new_n8879_), .A2(new_n8878_), .A3(new_n8881_), .ZN(new_n9986_));
  AOI21_X1   g09904(.A1(new_n8866_), .A2(new_n8869_), .B(new_n8876_), .ZN(new_n9987_));
  NOR2_X1    g09905(.A1(new_n9986_), .A2(new_n9987_), .ZN(new_n9988_));
  NAND3_X1   g09906(.A1(new_n9288_), .A2(new_n9284_), .A3(new_n8877_), .ZN(new_n9989_));
  NAND3_X1   g09907(.A1(new_n9989_), .A2(new_n9275_), .A3(new_n9988_), .ZN(new_n9990_));
  INV_X1     g09908(.I(new_n9990_), .ZN(new_n9991_));
  AOI21_X1   g09909(.A1(new_n9989_), .A2(new_n9275_), .B(new_n9988_), .ZN(new_n9992_));
  NOR2_X1    g09910(.A1(new_n9991_), .A2(new_n9992_), .ZN(new_n9993_));
  INV_X1     g09911(.I(new_n9993_), .ZN(new_n9994_));
  AOI21_X1   g09912(.A1(new_n9280_), .A2(new_n9278_), .B(new_n9283_), .ZN(new_n9995_));
  OAI21_X1   g09913(.A1(new_n9292_), .A2(new_n9995_), .B(new_n9986_), .ZN(new_n9996_));
  AOI21_X1   g09914(.A1(new_n9996_), .A2(new_n9381_), .B(new_n9988_), .ZN(new_n9997_));
  OAI21_X1   g09915(.A1(new_n8851_), .A2(new_n8847_), .B(new_n9301_), .ZN(new_n9998_));
  NOR2_X1    g09916(.A1(new_n9997_), .A2(new_n9998_), .ZN(new_n9999_));
  OAI21_X1   g09917(.A1(new_n8849_), .A2(new_n8850_), .B(new_n8848_), .ZN(new_n10000_));
  NAND3_X1   g09918(.A1(new_n8846_), .A2(new_n8844_), .A3(new_n8705_), .ZN(new_n10001_));
  AOI21_X1   g09919(.A1(new_n10000_), .A2(new_n10001_), .B(new_n9300_), .ZN(new_n10002_));
  NOR2_X1    g09920(.A1(new_n9290_), .A2(new_n10002_), .ZN(new_n10003_));
  OAI21_X1   g09921(.A1(new_n9999_), .A2(new_n10003_), .B(new_n9284_), .ZN(new_n10004_));
  NAND2_X1   g09922(.A1(new_n9290_), .A2(new_n10002_), .ZN(new_n10005_));
  NAND2_X1   g09923(.A1(new_n9997_), .A2(new_n9998_), .ZN(new_n10006_));
  NAND3_X1   g09924(.A1(new_n10006_), .A2(new_n10005_), .A3(new_n9292_), .ZN(new_n10007_));
  NOR2_X1    g09925(.A1(new_n4501_), .A2(new_n9405_), .ZN(new_n10008_));
  NOR2_X1    g09926(.A1(new_n4468_), .A2(new_n9408_), .ZN(new_n10009_));
  OAI22_X1   g09927(.A1(new_n4516_), .A2(new_n3456_), .B1(new_n10008_), .B2(new_n10009_), .ZN(new_n10010_));
  AOI21_X1   g09928(.A1(new_n10010_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n10011_));
  XOR2_X1    g09929(.A1(new_n4524_), .A2(new_n10011_), .Z(new_n10012_));
  NAND3_X1   g09930(.A1(new_n10004_), .A2(new_n10007_), .A3(new_n10012_), .ZN(new_n10013_));
  AOI21_X1   g09931(.A1(new_n10006_), .A2(new_n10005_), .B(new_n9292_), .ZN(new_n10014_));
  NOR3_X1    g09932(.A1(new_n9999_), .A2(new_n10003_), .A3(new_n9284_), .ZN(new_n10015_));
  INV_X1     g09933(.I(new_n10012_), .ZN(new_n10016_));
  OAI21_X1   g09934(.A1(new_n10014_), .A2(new_n10015_), .B(new_n10016_), .ZN(new_n10017_));
  NAND2_X1   g09935(.A1(new_n10017_), .A2(new_n10013_), .ZN(new_n10018_));
  NOR2_X1    g09936(.A1(new_n10018_), .A2(new_n9994_), .ZN(new_n10019_));
  AOI22_X1   g09937(.A1(new_n4473_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n4555_), .ZN(new_n10020_));
  OAI21_X1   g09938(.A1(new_n10020_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n10021_));
  NOR3_X1    g09939(.A1(new_n4583_), .A2(new_n4581_), .A3(new_n10021_), .ZN(new_n10022_));
  OAI21_X1   g09940(.A1(new_n4583_), .A2(new_n4581_), .B(new_n10021_), .ZN(new_n10023_));
  INV_X1     g09941(.I(new_n10023_), .ZN(new_n10024_));
  NOR2_X1    g09942(.A1(new_n10024_), .A2(new_n10022_), .ZN(new_n10025_));
  NAND2_X1   g09943(.A1(new_n10018_), .A2(new_n9994_), .ZN(new_n10026_));
  AOI21_X1   g09944(.A1(new_n10025_), .A2(new_n10026_), .B(new_n10019_), .ZN(new_n10027_));
  INV_X1     g09945(.I(new_n10027_), .ZN(new_n10028_));
  NOR2_X1    g09946(.A1(new_n9985_), .A2(new_n10028_), .ZN(new_n10029_));
  NAND2_X1   g09947(.A1(new_n10029_), .A2(new_n9362_), .ZN(new_n10030_));
  NAND2_X1   g09948(.A1(new_n10004_), .A2(new_n10007_), .ZN(new_n10031_));
  NAND2_X1   g09949(.A1(new_n10031_), .A2(new_n10012_), .ZN(new_n10032_));
  OAI22_X1   g09950(.A1(new_n5552_), .A2(new_n9425_), .B1(new_n3456_), .B2(new_n4563_), .ZN(new_n10033_));
  AOI21_X1   g09951(.A1(new_n10033_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n10034_));
  XOR2_X1    g09952(.A1(new_n4569_), .A2(new_n10034_), .Z(new_n10035_));
  INV_X1     g09953(.I(new_n10035_), .ZN(new_n10036_));
  NOR2_X1    g09954(.A1(new_n10032_), .A2(new_n10036_), .ZN(new_n10037_));
  OAI21_X1   g09955(.A1(new_n10029_), .A2(new_n9362_), .B(new_n10037_), .ZN(new_n10038_));
  INV_X1     g09956(.I(new_n8840_), .ZN(new_n10039_));
  NOR3_X1    g09957(.A1(new_n9324_), .A2(new_n9325_), .A3(new_n9327_), .ZN(new_n10040_));
  AOI21_X1   g09958(.A1(new_n9314_), .A2(new_n9311_), .B(new_n9322_), .ZN(new_n10041_));
  NOR2_X1    g09959(.A1(new_n10041_), .A2(new_n10040_), .ZN(new_n10042_));
  NAND2_X1   g09960(.A1(new_n10042_), .A2(new_n8836_), .ZN(new_n10043_));
  NAND3_X1   g09961(.A1(new_n10043_), .A2(new_n10039_), .A3(new_n9305_), .ZN(new_n10044_));
  INV_X1     g09962(.I(new_n10044_), .ZN(new_n10045_));
  AOI21_X1   g09963(.A1(new_n10043_), .A2(new_n9305_), .B(new_n10039_), .ZN(new_n10046_));
  NOR2_X1    g09964(.A1(new_n10045_), .A2(new_n10046_), .ZN(new_n10047_));
  OAI21_X1   g09965(.A1(new_n10042_), .A2(new_n8836_), .B(new_n9304_), .ZN(new_n10048_));
  AOI21_X1   g09966(.A1(new_n8822_), .A2(new_n8821_), .B(new_n8738_), .ZN(new_n10049_));
  NOR3_X1    g09967(.A1(new_n8818_), .A2(new_n8819_), .A3(new_n8813_), .ZN(new_n10050_));
  INV_X1     g09968(.I(new_n9336_), .ZN(new_n10051_));
  OAI21_X1   g09969(.A1(new_n10050_), .A2(new_n10049_), .B(new_n10051_), .ZN(new_n10052_));
  AOI21_X1   g09970(.A1(new_n10048_), .A2(new_n8840_), .B(new_n10052_), .ZN(new_n10053_));
  AOI21_X1   g09971(.A1(new_n8820_), .A2(new_n8823_), .B(new_n9336_), .ZN(new_n10054_));
  NOR2_X1    g09972(.A1(new_n9330_), .A2(new_n10054_), .ZN(new_n10055_));
  OAI21_X1   g09973(.A1(new_n10053_), .A2(new_n10055_), .B(new_n9323_), .ZN(new_n10056_));
  NAND2_X1   g09974(.A1(new_n9330_), .A2(new_n10054_), .ZN(new_n10057_));
  NAND3_X1   g09975(.A1(new_n10052_), .A2(new_n10048_), .A3(new_n8840_), .ZN(new_n10058_));
  NAND3_X1   g09976(.A1(new_n10058_), .A2(new_n10057_), .A3(new_n10040_), .ZN(new_n10059_));
  NOR3_X1    g09977(.A1(new_n3409_), .A2(new_n451_), .A3(\a[1] ), .ZN(new_n10060_));
  XNOR2_X1   g09978(.A1(new_n4609_), .A2(new_n10060_), .ZN(new_n10061_));
  NAND3_X1   g09979(.A1(new_n10056_), .A2(new_n10059_), .A3(new_n10061_), .ZN(new_n10062_));
  AOI21_X1   g09980(.A1(new_n10058_), .A2(new_n10057_), .B(new_n10040_), .ZN(new_n10063_));
  NOR3_X1    g09981(.A1(new_n10053_), .A2(new_n10055_), .A3(new_n9323_), .ZN(new_n10064_));
  INV_X1     g09982(.I(new_n10061_), .ZN(new_n10065_));
  OAI21_X1   g09983(.A1(new_n10064_), .A2(new_n10063_), .B(new_n10065_), .ZN(new_n10066_));
  NAND3_X1   g09984(.A1(new_n10066_), .A2(new_n10062_), .A3(new_n10047_), .ZN(new_n10067_));
  OAI22_X1   g09985(.A1(new_n4567_), .A2(new_n9425_), .B1(new_n3456_), .B2(new_n4564_), .ZN(new_n10068_));
  AOI21_X1   g09986(.A1(new_n10068_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n10069_));
  XOR2_X1    g09987(.A1(new_n4594_), .A2(new_n10069_), .Z(new_n10070_));
  INV_X1     g09988(.I(new_n10070_), .ZN(new_n10071_));
  AOI21_X1   g09989(.A1(new_n10066_), .A2(new_n10062_), .B(new_n10047_), .ZN(new_n10072_));
  OAI21_X1   g09990(.A1(new_n10071_), .A2(new_n10072_), .B(new_n10067_), .ZN(new_n10073_));
  AOI21_X1   g09991(.A1(new_n10030_), .A2(new_n10038_), .B(new_n10073_), .ZN(new_n10074_));
  NAND2_X1   g09992(.A1(new_n10074_), .A2(new_n9361_), .ZN(new_n10075_));
  NOR2_X1    g09993(.A1(new_n10064_), .A2(new_n10063_), .ZN(new_n10076_));
  NOR2_X1    g09994(.A1(new_n3456_), .A2(new_n9405_), .ZN(new_n10077_));
  AOI21_X1   g09995(.A1(new_n9408_), .A2(new_n10077_), .B(new_n4563_), .ZN(new_n10078_));
  AOI21_X1   g09996(.A1(new_n10078_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n10079_));
  XNOR2_X1   g09997(.A1(new_n5001_), .A2(new_n10079_), .ZN(new_n10080_));
  NOR3_X1    g09998(.A1(new_n10076_), .A2(new_n10065_), .A3(new_n10080_), .ZN(new_n10081_));
  OAI21_X1   g09999(.A1(new_n10074_), .A2(new_n9361_), .B(new_n10081_), .ZN(new_n10082_));
  NAND2_X1   g10000(.A1(new_n9357_), .A2(new_n9339_), .ZN(new_n10083_));
  AOI21_X1   g10001(.A1(new_n8750_), .A2(new_n8757_), .B(new_n8759_), .ZN(new_n10084_));
  INV_X1     g10002(.I(new_n8771_), .ZN(new_n10085_));
  AOI21_X1   g10003(.A1(new_n10085_), .A2(new_n8770_), .B(new_n10084_), .ZN(new_n10086_));
  INV_X1     g10004(.I(new_n8766_), .ZN(new_n10087_));
  AND3_X2    g10005(.A1(new_n10087_), .A2(new_n8764_), .A3(new_n8769_), .Z(new_n10088_));
  AOI21_X1   g10006(.A1(new_n10087_), .A2(new_n8764_), .B(new_n8769_), .ZN(new_n10089_));
  OAI21_X1   g10007(.A1(new_n10088_), .A2(new_n10089_), .B(new_n10084_), .ZN(new_n10090_));
  INV_X1     g10008(.I(new_n10090_), .ZN(new_n10091_));
  AOI22_X1   g10009(.A1(new_n5418_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n4563_), .ZN(new_n10092_));
  OAI21_X1   g10010(.A1(new_n10092_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n10093_));
  XNOR2_X1   g10011(.A1(new_n4594_), .A2(new_n10093_), .ZN(new_n10094_));
  OAI21_X1   g10012(.A1(new_n10091_), .A2(new_n10086_), .B(new_n10094_), .ZN(new_n10095_));
  INV_X1     g10013(.I(new_n8770_), .ZN(new_n10096_));
  OAI21_X1   g10014(.A1(new_n10096_), .A2(new_n8771_), .B(new_n8761_), .ZN(new_n10097_));
  INV_X1     g10015(.I(new_n10094_), .ZN(new_n10098_));
  NAND3_X1   g10016(.A1(new_n10097_), .A2(new_n10090_), .A3(new_n10098_), .ZN(new_n10099_));
  AOI22_X1   g10017(.A1(new_n10095_), .A2(new_n10099_), .B1(new_n10083_), .B2(new_n9358_), .ZN(new_n10100_));
  INV_X1     g10018(.I(new_n10100_), .ZN(new_n10101_));
  NAND3_X1   g10019(.A1(new_n10097_), .A2(new_n10090_), .A3(new_n10094_), .ZN(new_n10102_));
  OAI21_X1   g10020(.A1(new_n10091_), .A2(new_n10086_), .B(new_n10098_), .ZN(new_n10103_));
  NAND2_X1   g10021(.A1(new_n10103_), .A2(new_n10102_), .ZN(new_n10104_));
  NAND3_X1   g10022(.A1(new_n10104_), .A2(new_n10083_), .A3(new_n9358_), .ZN(new_n10105_));
  NOR3_X1    g10023(.A1(new_n3409_), .A2(new_n451_), .A3(\a[1] ), .ZN(new_n10106_));
  XNOR2_X1   g10024(.A1(new_n4610_), .A2(new_n10106_), .ZN(new_n10107_));
  INV_X1     g10025(.I(new_n10107_), .ZN(new_n10108_));
  AOI21_X1   g10026(.A1(new_n10101_), .A2(new_n10105_), .B(new_n10108_), .ZN(new_n10109_));
  AOI21_X1   g10027(.A1(new_n10082_), .A2(new_n10075_), .B(new_n10109_), .ZN(new_n10110_));
  INV_X1     g10028(.I(new_n10110_), .ZN(new_n10111_));
  INV_X1     g10029(.I(new_n10105_), .ZN(new_n10112_));
  NOR3_X1    g10030(.A1(new_n10112_), .A2(new_n10100_), .A3(new_n10107_), .ZN(new_n10113_));
  INV_X1     g10031(.I(new_n10113_), .ZN(new_n10114_));
  OAI21_X1   g10032(.A1(new_n10084_), .A2(new_n10096_), .B(new_n10085_), .ZN(new_n10115_));
  NOR3_X1    g10033(.A1(new_n8795_), .A2(new_n8796_), .A3(new_n8793_), .ZN(new_n10116_));
  AOI21_X1   g10034(.A1(new_n8788_), .A2(new_n8785_), .B(new_n8792_), .ZN(new_n10117_));
  OAI21_X1   g10035(.A1(new_n10116_), .A2(new_n10117_), .B(new_n10115_), .ZN(new_n10118_));
  OAI21_X1   g10036(.A1(new_n8794_), .A2(new_n8797_), .B(new_n8772_), .ZN(new_n10119_));
  NAND2_X1   g10037(.A1(new_n4564_), .A2(new_n5031_), .ZN(new_n10120_));
  NAND2_X1   g10038(.A1(new_n4563_), .A2(new_n5033_), .ZN(new_n10121_));
  AOI22_X1   g10039(.A1(new_n10120_), .A2(new_n10121_), .B1(new_n2898_), .B2(new_n4564_), .ZN(new_n10122_));
  OAI21_X1   g10040(.A1(new_n10122_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n10123_));
  XOR2_X1    g10041(.A1(new_n4609_), .A2(new_n10123_), .Z(new_n10124_));
  INV_X1     g10042(.I(new_n10124_), .ZN(new_n10125_));
  NAND3_X1   g10043(.A1(new_n10118_), .A2(new_n10119_), .A3(new_n10125_), .ZN(new_n10126_));
  NOR2_X1    g10044(.A1(new_n10116_), .A2(new_n10117_), .ZN(new_n10127_));
  NOR2_X1    g10045(.A1(new_n10127_), .A2(new_n8772_), .ZN(new_n10128_));
  INV_X1     g10046(.I(new_n10119_), .ZN(new_n10129_));
  OAI21_X1   g10047(.A1(new_n10129_), .A2(new_n10128_), .B(new_n10124_), .ZN(new_n10130_));
  NAND2_X1   g10048(.A1(new_n10130_), .A2(new_n10126_), .ZN(new_n10131_));
  INV_X1     g10049(.I(new_n9358_), .ZN(new_n10132_));
  NOR3_X1    g10050(.A1(new_n9341_), .A2(new_n9346_), .A3(new_n9354_), .ZN(new_n10133_));
  NOR2_X1    g10051(.A1(new_n9340_), .A2(new_n10133_), .ZN(new_n10134_));
  OAI21_X1   g10052(.A1(new_n10134_), .A2(new_n10132_), .B(new_n10102_), .ZN(new_n10135_));
  AOI21_X1   g10053(.A1(new_n10135_), .A2(new_n10103_), .B(new_n3413_), .ZN(new_n10136_));
  INV_X1     g10054(.I(new_n10103_), .ZN(new_n10137_));
  NOR2_X1    g10055(.A1(new_n10091_), .A2(new_n10086_), .ZN(new_n10138_));
  AOI22_X1   g10056(.A1(new_n10083_), .A2(new_n9358_), .B1(new_n10138_), .B2(new_n10094_), .ZN(new_n10139_));
  NOR3_X1    g10057(.A1(new_n10139_), .A2(new_n3412_), .A3(new_n10137_), .ZN(new_n10140_));
  OAI21_X1   g10058(.A1(new_n10140_), .A2(new_n10136_), .B(new_n10131_), .ZN(new_n10141_));
  INV_X1     g10059(.I(new_n10126_), .ZN(new_n10142_));
  AOI21_X1   g10060(.A1(new_n10118_), .A2(new_n10119_), .B(new_n10125_), .ZN(new_n10143_));
  NOR2_X1    g10061(.A1(new_n10142_), .A2(new_n10143_), .ZN(new_n10144_));
  NOR3_X1    g10062(.A1(new_n10139_), .A2(new_n3413_), .A3(new_n10137_), .ZN(new_n10145_));
  AOI21_X1   g10063(.A1(new_n10135_), .A2(new_n10103_), .B(new_n3412_), .ZN(new_n10146_));
  OAI21_X1   g10064(.A1(new_n10145_), .A2(new_n10146_), .B(new_n10144_), .ZN(new_n10147_));
  NAND2_X1   g10065(.A1(new_n10147_), .A2(new_n10141_), .ZN(new_n10148_));
  NAND3_X1   g10066(.A1(new_n10111_), .A2(new_n10114_), .A3(new_n10148_), .ZN(new_n10149_));
  NOR2_X1    g10067(.A1(new_n10149_), .A2(new_n8812_), .ZN(new_n10150_));
  NOR2_X1    g10068(.A1(new_n10139_), .A2(new_n10137_), .ZN(new_n10151_));
  XOR2_X1    g10069(.A1(new_n10131_), .A2(new_n3413_), .Z(new_n10152_));
  NAND2_X1   g10070(.A1(new_n10152_), .A2(new_n10151_), .ZN(new_n10153_));
  INV_X1     g10071(.I(new_n10153_), .ZN(new_n10154_));
  NAND2_X1   g10072(.A1(new_n10125_), .A2(new_n3413_), .ZN(new_n10155_));
  NAND2_X1   g10073(.A1(new_n10124_), .A2(new_n3412_), .ZN(new_n10156_));
  NAND3_X1   g10074(.A1(new_n10118_), .A2(new_n10119_), .A3(new_n10156_), .ZN(new_n10157_));
  NAND2_X1   g10075(.A1(new_n10157_), .A2(new_n10155_), .ZN(new_n10158_));
  NAND2_X1   g10076(.A1(new_n10154_), .A2(new_n10158_), .ZN(new_n10159_));
  AOI21_X1   g10077(.A1(new_n8812_), .A2(new_n10149_), .B(new_n10159_), .ZN(new_n10160_));
  XOR2_X1    g10078(.A1(new_n7843_), .A2(new_n7841_), .Z(new_n10161_));
  XOR2_X1    g10079(.A1(new_n10161_), .A2(new_n7835_), .Z(new_n10162_));
  XOR2_X1    g10080(.A1(new_n10162_), .A2(new_n7451_), .Z(new_n10163_));
  NOR2_X1    g10081(.A1(new_n8329_), .A2(new_n8333_), .ZN(new_n10164_));
  NAND2_X1   g10082(.A1(new_n8329_), .A2(new_n8333_), .ZN(new_n10165_));
  XOR2_X1    g10083(.A1(new_n8330_), .A2(new_n7828_), .Z(new_n10166_));
  AOI21_X1   g10084(.A1(new_n10166_), .A2(new_n10165_), .B(new_n10164_), .ZN(new_n10167_));
  INV_X1     g10085(.I(new_n10167_), .ZN(new_n10168_));
  NAND3_X1   g10086(.A1(new_n4563_), .A2(new_n2898_), .A3(new_n3042_), .ZN(new_n10169_));
  AOI21_X1   g10087(.A1(new_n10169_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n10170_));
  XNOR2_X1   g10088(.A1(new_n4610_), .A2(new_n10170_), .ZN(new_n10171_));
  INV_X1     g10089(.I(new_n10171_), .ZN(new_n10172_));
  NOR2_X1    g10090(.A1(new_n10168_), .A2(new_n10172_), .ZN(new_n10173_));
  INV_X1     g10091(.I(new_n10173_), .ZN(new_n10174_));
  NOR2_X1    g10092(.A1(new_n10167_), .A2(new_n10171_), .ZN(new_n10175_));
  INV_X1     g10093(.I(new_n10175_), .ZN(new_n10176_));
  AOI21_X1   g10094(.A1(new_n10174_), .A2(new_n10176_), .B(new_n10163_), .ZN(new_n10177_));
  XOR2_X1    g10095(.A1(new_n10162_), .A2(new_n7452_), .Z(new_n10178_));
  XOR2_X1    g10096(.A1(new_n10167_), .A2(new_n10172_), .Z(new_n10179_));
  NOR2_X1    g10097(.A1(new_n10178_), .A2(new_n10179_), .ZN(new_n10180_));
  NOR2_X1    g10098(.A1(new_n10177_), .A2(new_n10180_), .ZN(new_n10181_));
  OAI21_X1   g10099(.A1(new_n8809_), .A2(new_n8805_), .B(new_n8806_), .ZN(new_n10182_));
  INV_X1     g10100(.I(new_n10182_), .ZN(new_n10183_));
  NAND2_X1   g10101(.A1(new_n10181_), .A2(new_n10183_), .ZN(new_n10184_));
  OAI21_X1   g10102(.A1(new_n10160_), .A2(new_n10150_), .B(new_n10184_), .ZN(new_n10185_));
  NOR2_X1    g10103(.A1(new_n10181_), .A2(new_n10183_), .ZN(new_n10186_));
  INV_X1     g10104(.I(new_n10186_), .ZN(new_n10187_));
  XOR2_X1    g10105(.A1(new_n7846_), .A2(new_n2899_), .Z(new_n10188_));
  INV_X1     g10106(.I(new_n10188_), .ZN(new_n10189_));
  OAI21_X1   g10107(.A1(new_n10163_), .A2(new_n10173_), .B(new_n10176_), .ZN(new_n10190_));
  XOR2_X1    g10108(.A1(new_n10190_), .A2(new_n10189_), .Z(new_n10191_));
  NOR2_X1    g10109(.A1(new_n10191_), .A2(new_n7468_), .ZN(new_n10192_));
  XOR2_X1    g10110(.A1(new_n10190_), .A2(new_n10189_), .Z(new_n10193_));
  AOI21_X1   g10111(.A1(new_n10193_), .A2(new_n7468_), .B(new_n10192_), .ZN(new_n10194_));
  INV_X1     g10112(.I(new_n10194_), .ZN(new_n10195_));
  NAND3_X1   g10113(.A1(new_n10185_), .A2(new_n10195_), .A3(new_n10187_), .ZN(new_n10196_));
  XOR2_X1    g10114(.A1(new_n7468_), .A2(new_n10188_), .Z(new_n10197_));
  NOR2_X1    g10115(.A1(new_n10197_), .A2(new_n10190_), .ZN(new_n10198_));
  INV_X1     g10116(.I(new_n10198_), .ZN(new_n10199_));
  NOR2_X1    g10117(.A1(new_n7872_), .A2(new_n7849_), .ZN(new_n10200_));
  OR3_X2     g10118(.A1(new_n10196_), .A2(new_n10199_), .A3(new_n10200_), .Z(new_n10201_));
  NAND2_X1   g10119(.A1(new_n7869_), .A2(new_n7851_), .ZN(new_n10202_));
  NAND2_X1   g10120(.A1(new_n10202_), .A2(new_n7870_), .ZN(new_n10203_));
  INV_X1     g10121(.I(new_n10203_), .ZN(new_n10204_));
  XOR2_X1    g10122(.A1(new_n6791_), .A2(new_n2470_), .Z(new_n10205_));
  XNOR2_X1   g10123(.A1(new_n6767_), .A2(new_n10205_), .ZN(new_n10206_));
  XOR2_X1    g10124(.A1(new_n10206_), .A2(new_n6796_), .Z(new_n10207_));
  NAND2_X1   g10125(.A1(new_n6764_), .A2(new_n6766_), .ZN(new_n10208_));
  XOR2_X1    g10126(.A1(new_n6755_), .A2(new_n6761_), .Z(new_n10209_));
  NOR2_X1    g10127(.A1(new_n6481_), .A2(new_n10209_), .ZN(new_n10210_));
  AOI21_X1   g10128(.A1(new_n6481_), .A2(new_n10208_), .B(new_n10210_), .ZN(new_n10211_));
  INV_X1     g10129(.I(new_n10211_), .ZN(new_n10212_));
  NOR2_X1    g10130(.A1(new_n7859_), .A2(new_n7854_), .ZN(new_n10213_));
  AOI21_X1   g10131(.A1(new_n7854_), .A2(new_n7859_), .B(new_n7861_), .ZN(new_n10214_));
  NOR2_X1    g10132(.A1(new_n10214_), .A2(new_n10213_), .ZN(new_n10215_));
  INV_X1     g10133(.I(new_n10215_), .ZN(new_n10216_));
  NAND3_X1   g10134(.A1(new_n4563_), .A2(new_n2469_), .A3(new_n2718_), .ZN(new_n10217_));
  AOI21_X1   g10135(.A1(new_n10217_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n10218_));
  XNOR2_X1   g10136(.A1(new_n4610_), .A2(new_n10218_), .ZN(new_n10219_));
  INV_X1     g10137(.I(new_n10219_), .ZN(new_n10220_));
  NOR2_X1    g10138(.A1(new_n10216_), .A2(new_n10220_), .ZN(new_n10221_));
  INV_X1     g10139(.I(new_n10221_), .ZN(new_n10222_));
  NOR2_X1    g10140(.A1(new_n10215_), .A2(new_n10219_), .ZN(new_n10223_));
  AOI21_X1   g10141(.A1(new_n10222_), .A2(new_n10212_), .B(new_n10223_), .ZN(new_n10224_));
  XNOR2_X1   g10142(.A1(new_n10207_), .A2(new_n10224_), .ZN(new_n10225_));
  NAND2_X1   g10143(.A1(new_n10225_), .A2(new_n10204_), .ZN(new_n10226_));
  OAI21_X1   g10144(.A1(new_n10221_), .A2(new_n10223_), .B(new_n10212_), .ZN(new_n10227_));
  XOR2_X1    g10145(.A1(new_n10215_), .A2(new_n10220_), .Z(new_n10228_));
  OAI21_X1   g10146(.A1(new_n10212_), .A2(new_n10228_), .B(new_n10227_), .ZN(new_n10229_));
  INV_X1     g10147(.I(new_n10229_), .ZN(new_n10230_));
  OAI21_X1   g10148(.A1(new_n10225_), .A2(new_n10204_), .B(new_n10230_), .ZN(new_n10231_));
  NAND2_X1   g10149(.A1(new_n10231_), .A2(new_n10226_), .ZN(new_n10232_));
  AOI21_X1   g10150(.A1(new_n10201_), .A2(new_n7873_), .B(new_n10232_), .ZN(new_n10233_));
  NAND2_X1   g10151(.A1(new_n10207_), .A2(new_n10224_), .ZN(new_n10234_));
  AOI21_X1   g10152(.A1(new_n6827_), .A2(new_n6799_), .B(new_n10234_), .ZN(new_n10235_));
  AOI21_X1   g10153(.A1(new_n10233_), .A2(new_n10235_), .B(new_n6828_), .ZN(new_n10236_));
  NOR2_X1    g10154(.A1(new_n5972_), .A2(new_n5974_), .ZN(new_n10237_));
  XOR2_X1    g10155(.A1(new_n5965_), .A2(new_n5971_), .Z(new_n10238_));
  NAND2_X1   g10156(.A1(new_n10238_), .A2(new_n5887_), .ZN(new_n10239_));
  OAI21_X1   g10157(.A1(new_n5887_), .A2(new_n10237_), .B(new_n10239_), .ZN(new_n10240_));
  NOR2_X1    g10158(.A1(new_n6807_), .A2(new_n6805_), .ZN(new_n10241_));
  AOI21_X1   g10159(.A1(new_n6805_), .A2(new_n6807_), .B(new_n6813_), .ZN(new_n10242_));
  NOR2_X1    g10160(.A1(new_n10242_), .A2(new_n10241_), .ZN(new_n10243_));
  INV_X1     g10161(.I(new_n10243_), .ZN(new_n10244_));
  NAND3_X1   g10162(.A1(new_n4563_), .A2(new_n805_), .A3(new_n2258_), .ZN(new_n10245_));
  AOI21_X1   g10163(.A1(new_n10245_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n10246_));
  XNOR2_X1   g10164(.A1(new_n4610_), .A2(new_n10246_), .ZN(new_n10247_));
  INV_X1     g10165(.I(new_n10247_), .ZN(new_n10248_));
  NOR2_X1    g10166(.A1(new_n10244_), .A2(new_n10248_), .ZN(new_n10249_));
  NOR2_X1    g10167(.A1(new_n10243_), .A2(new_n10247_), .ZN(new_n10250_));
  OAI21_X1   g10168(.A1(new_n10249_), .A2(new_n10250_), .B(new_n10240_), .ZN(new_n10251_));
  XOR2_X1    g10169(.A1(new_n10243_), .A2(new_n10248_), .Z(new_n10252_));
  OAI21_X1   g10170(.A1(new_n10240_), .A2(new_n10252_), .B(new_n10251_), .ZN(new_n10253_));
  OAI21_X1   g10171(.A1(new_n6802_), .A2(new_n6823_), .B(new_n6825_), .ZN(new_n10254_));
  NOR2_X1    g10172(.A1(new_n10254_), .A2(new_n10253_), .ZN(new_n10255_));
  INV_X1     g10173(.I(new_n10255_), .ZN(new_n10256_));
  NAND2_X1   g10174(.A1(new_n10254_), .A2(new_n10253_), .ZN(new_n10257_));
  NOR2_X1    g10175(.A1(new_n6010_), .A2(new_n6012_), .ZN(new_n10258_));
  NOR2_X1    g10176(.A1(new_n10258_), .A2(new_n5975_), .ZN(new_n10259_));
  XOR2_X1    g10177(.A1(new_n6008_), .A2(new_n806_), .Z(new_n10260_));
  AOI21_X1   g10178(.A1(new_n5975_), .A2(new_n10260_), .B(new_n10259_), .ZN(new_n10261_));
  INV_X1     g10179(.I(new_n10249_), .ZN(new_n10262_));
  AOI21_X1   g10180(.A1(new_n10262_), .A2(new_n10240_), .B(new_n10250_), .ZN(new_n10263_));
  XNOR2_X1   g10181(.A1(new_n10261_), .A2(new_n10263_), .ZN(new_n10264_));
  NAND2_X1   g10182(.A1(new_n10256_), .A2(new_n10257_), .ZN(new_n10265_));
  INV_X1     g10183(.I(new_n10265_), .ZN(new_n10266_));
  NAND2_X1   g10184(.A1(new_n10261_), .A2(new_n10263_), .ZN(new_n10267_));
  AND2_X2    g10185(.A1(new_n6037_), .A2(new_n6013_), .Z(new_n10268_));
  NOR4_X1    g10186(.A1(new_n10236_), .A2(new_n10266_), .A3(new_n10267_), .A4(new_n10268_), .ZN(new_n10269_));
  NOR2_X1    g10187(.A1(new_n10269_), .A2(new_n6038_), .ZN(new_n10270_));
  INV_X1     g10188(.I(new_n10270_), .ZN(new_n10271_));
  INV_X1     g10189(.I(new_n5427_), .ZN(new_n10272_));
  OAI21_X1   g10190(.A1(new_n10272_), .A2(new_n5426_), .B(new_n5349_), .ZN(new_n10273_));
  XOR2_X1    g10191(.A1(new_n5417_), .A2(new_n5424_), .Z(new_n10274_));
  OAI21_X1   g10192(.A1(new_n5349_), .A2(new_n10274_), .B(new_n10273_), .ZN(new_n10275_));
  NOR2_X1    g10193(.A1(new_n6020_), .A2(new_n6018_), .ZN(new_n10276_));
  AOI21_X1   g10194(.A1(new_n6018_), .A2(new_n6020_), .B(new_n6023_), .ZN(new_n10277_));
  NOR2_X1    g10195(.A1(new_n10277_), .A2(new_n10276_), .ZN(new_n10278_));
  INV_X1     g10196(.I(new_n10278_), .ZN(new_n10279_));
  NAND3_X1   g10197(.A1(new_n4563_), .A2(new_n785_), .A3(new_n1851_), .ZN(new_n10280_));
  AOI21_X1   g10198(.A1(new_n10280_), .A2(new_n279_), .B(new_n643_), .ZN(new_n10281_));
  XNOR2_X1   g10199(.A1(new_n4610_), .A2(new_n10281_), .ZN(new_n10282_));
  INV_X1     g10200(.I(new_n10282_), .ZN(new_n10283_));
  NOR2_X1    g10201(.A1(new_n10279_), .A2(new_n10283_), .ZN(new_n10284_));
  NOR2_X1    g10202(.A1(new_n10278_), .A2(new_n10282_), .ZN(new_n10285_));
  OAI21_X1   g10203(.A1(new_n10284_), .A2(new_n10285_), .B(new_n10275_), .ZN(new_n10286_));
  XOR2_X1    g10204(.A1(new_n10278_), .A2(new_n10283_), .Z(new_n10287_));
  OAI21_X1   g10205(.A1(new_n10275_), .A2(new_n10287_), .B(new_n10286_), .ZN(new_n10288_));
  OAI21_X1   g10206(.A1(new_n6015_), .A2(new_n6033_), .B(new_n6035_), .ZN(new_n10289_));
  NOR2_X1    g10207(.A1(new_n10289_), .A2(new_n10288_), .ZN(new_n10290_));
  INV_X1     g10208(.I(new_n10290_), .ZN(new_n10291_));
  NAND2_X1   g10209(.A1(new_n10289_), .A2(new_n10288_), .ZN(new_n10292_));
  NOR2_X1    g10210(.A1(new_n5500_), .A2(new_n5502_), .ZN(new_n10293_));
  XOR2_X1    g10211(.A1(new_n5498_), .A2(new_n644_), .Z(new_n10294_));
  MUX2_X1    g10212(.I0(new_n10294_), .I1(new_n10293_), .S(new_n5428_), .Z(new_n10295_));
  INV_X1     g10213(.I(new_n10284_), .ZN(new_n10296_));
  AOI21_X1   g10214(.A1(new_n10296_), .A2(new_n10275_), .B(new_n10285_), .ZN(new_n10297_));
  XNOR2_X1   g10215(.A1(new_n10297_), .A2(new_n10295_), .ZN(new_n10298_));
  NAND2_X1   g10216(.A1(new_n10291_), .A2(new_n10292_), .ZN(new_n10299_));
  NAND2_X1   g10217(.A1(new_n10271_), .A2(new_n10299_), .ZN(new_n10300_));
  NAND2_X1   g10218(.A1(new_n10297_), .A2(new_n10295_), .ZN(new_n10301_));
  AOI21_X1   g10219(.A1(new_n5503_), .A2(new_n5577_), .B(new_n10301_), .ZN(new_n10302_));
  INV_X1     g10220(.I(new_n10302_), .ZN(new_n10303_));
  OAI21_X1   g10221(.A1(new_n10300_), .A2(new_n10303_), .B(new_n5579_), .ZN(new_n10304_));
  OAI21_X1   g10222(.A1(new_n5505_), .A2(new_n5573_), .B(new_n5575_), .ZN(new_n10305_));
  XOR2_X1    g10223(.A1(new_n5539_), .A2(new_n5544_), .Z(new_n10306_));
  NOR2_X1    g10224(.A1(new_n10306_), .A2(new_n5541_), .ZN(new_n10307_));
  NOR2_X1    g10225(.A1(new_n5539_), .A2(new_n5545_), .ZN(new_n10308_));
  INV_X1     g10226(.I(new_n10308_), .ZN(new_n10309_));
  NOR2_X1    g10227(.A1(new_n5521_), .A2(new_n5507_), .ZN(new_n10310_));
  NOR2_X1    g10228(.A1(new_n10310_), .A2(new_n5522_), .ZN(new_n10311_));
  XOR2_X1    g10229(.A1(new_n4955_), .A2(new_n4657_), .Z(new_n10312_));
  OAI21_X1   g10230(.A1(new_n4957_), .A2(new_n4959_), .B(new_n4950_), .ZN(new_n10313_));
  OAI21_X1   g10231(.A1(new_n4950_), .A2(new_n10312_), .B(new_n10313_), .ZN(new_n10314_));
  AOI22_X1   g10232(.A1(new_n4018_), .A2(new_n4613_), .B1(new_n4375_), .B2(new_n4767_), .ZN(new_n10315_));
  AOI21_X1   g10233(.A1(new_n117_), .A2(new_n4399_), .B(new_n10315_), .ZN(new_n10316_));
  OAI21_X1   g10234(.A1(new_n10316_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n10317_));
  XOR2_X1    g10235(.A1(new_n4403_), .A2(new_n10317_), .Z(new_n10318_));
  AND2_X2    g10236(.A1(new_n10314_), .A2(new_n10318_), .Z(new_n10319_));
  NOR2_X1    g10237(.A1(new_n10314_), .A2(new_n10318_), .ZN(new_n10320_));
  NOR2_X1    g10238(.A1(new_n10319_), .A2(new_n10320_), .ZN(new_n10321_));
  NOR2_X1    g10239(.A1(new_n10321_), .A2(new_n10311_), .ZN(new_n10322_));
  XNOR2_X1   g10240(.A1(new_n10314_), .A2(new_n10318_), .ZN(new_n10323_));
  INV_X1     g10241(.I(new_n10323_), .ZN(new_n10324_));
  AOI21_X1   g10242(.A1(new_n10311_), .A2(new_n10324_), .B(new_n10322_), .ZN(new_n10325_));
  INV_X1     g10243(.I(new_n5532_), .ZN(new_n10326_));
  AOI21_X1   g10244(.A1(new_n10326_), .A2(new_n5525_), .B(new_n5534_), .ZN(new_n10327_));
  OAI22_X1   g10245(.A1(new_n4472_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4501_), .ZN(new_n10328_));
  AOI21_X1   g10246(.A1(new_n10328_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n10329_));
  XOR2_X1    g10247(.A1(new_n4584_), .A2(new_n10329_), .Z(new_n10330_));
  AND2_X2    g10248(.A1(new_n10330_), .A2(new_n10327_), .Z(new_n10331_));
  NOR2_X1    g10249(.A1(new_n10330_), .A2(new_n10327_), .ZN(new_n10332_));
  NOR2_X1    g10250(.A1(new_n10331_), .A2(new_n10332_), .ZN(new_n10333_));
  NOR2_X1    g10251(.A1(new_n10333_), .A2(new_n10325_), .ZN(new_n10334_));
  INV_X1     g10252(.I(new_n10325_), .ZN(new_n10335_));
  XNOR2_X1   g10253(.A1(new_n10330_), .A2(new_n10327_), .ZN(new_n10336_));
  NOR2_X1    g10254(.A1(new_n10336_), .A2(new_n10335_), .ZN(new_n10337_));
  NOR2_X1    g10255(.A1(new_n10334_), .A2(new_n10337_), .ZN(new_n10338_));
  AOI22_X1   g10256(.A1(new_n5418_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n4563_), .ZN(new_n10339_));
  OAI21_X1   g10257(.A1(new_n10339_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n10340_));
  XNOR2_X1   g10258(.A1(new_n4594_), .A2(new_n10340_), .ZN(new_n10341_));
  NOR2_X1    g10259(.A1(new_n10338_), .A2(new_n10341_), .ZN(new_n10342_));
  XOR2_X1    g10260(.A1(new_n10342_), .A2(new_n10309_), .Z(new_n10343_));
  XOR2_X1    g10261(.A1(new_n10343_), .A2(new_n10307_), .Z(new_n10344_));
  OAI21_X1   g10262(.A1(new_n5562_), .A2(new_n5558_), .B(new_n5560_), .ZN(new_n10345_));
  NAND3_X1   g10263(.A1(new_n4563_), .A2(new_n4660_), .A3(new_n1622_), .ZN(new_n10346_));
  AOI21_X1   g10264(.A1(new_n10346_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n10347_));
  XNOR2_X1   g10265(.A1(new_n4610_), .A2(new_n10347_), .ZN(new_n10348_));
  INV_X1     g10266(.I(new_n10348_), .ZN(new_n10349_));
  NOR2_X1    g10267(.A1(new_n10345_), .A2(new_n10349_), .ZN(new_n10350_));
  INV_X1     g10268(.I(new_n10350_), .ZN(new_n10351_));
  NAND2_X1   g10269(.A1(new_n10345_), .A2(new_n10349_), .ZN(new_n10352_));
  AOI21_X1   g10270(.A1(new_n10351_), .A2(new_n10352_), .B(new_n10344_), .ZN(new_n10353_));
  INV_X1     g10271(.I(new_n10344_), .ZN(new_n10354_));
  XOR2_X1    g10272(.A1(new_n10345_), .A2(new_n10348_), .Z(new_n10355_));
  NOR2_X1    g10273(.A1(new_n10354_), .A2(new_n10355_), .ZN(new_n10356_));
  NOR2_X1    g10274(.A1(new_n10356_), .A2(new_n10353_), .ZN(new_n10357_));
  INV_X1     g10275(.I(new_n10357_), .ZN(new_n10358_));
  NOR2_X1    g10276(.A1(new_n10358_), .A2(new_n10305_), .ZN(new_n10359_));
  INV_X1     g10277(.I(new_n10359_), .ZN(new_n10360_));
  NAND2_X1   g10278(.A1(new_n10358_), .A2(new_n10305_), .ZN(new_n10361_));
  INV_X1     g10279(.I(new_n10361_), .ZN(new_n10362_));
  AOI21_X1   g10280(.A1(new_n10304_), .A2(new_n10360_), .B(new_n10362_), .ZN(new_n10363_));
  NOR2_X1    g10281(.A1(new_n10338_), .A2(new_n10309_), .ZN(new_n10364_));
  NOR3_X1    g10282(.A1(new_n10334_), .A2(new_n10337_), .A3(new_n10308_), .ZN(new_n10365_));
  NOR4_X1    g10283(.A1(new_n10365_), .A2(new_n5541_), .A3(new_n10306_), .A4(new_n10341_), .ZN(new_n10366_));
  NOR2_X1    g10284(.A1(new_n10366_), .A2(new_n10364_), .ZN(new_n10367_));
  NOR2_X1    g10285(.A1(new_n10319_), .A2(new_n10311_), .ZN(new_n10368_));
  INV_X1     g10286(.I(new_n4968_), .ZN(new_n10369_));
  XNOR2_X1   g10287(.A1(new_n4963_), .A2(new_n4960_), .ZN(new_n10370_));
  NOR2_X1    g10288(.A1(new_n10370_), .A2(new_n10369_), .ZN(new_n10371_));
  NOR2_X1    g10289(.A1(new_n4969_), .A2(new_n4964_), .ZN(new_n10372_));
  NOR2_X1    g10290(.A1(new_n10372_), .A2(new_n4968_), .ZN(new_n10373_));
  NOR2_X1    g10291(.A1(new_n10373_), .A2(new_n10371_), .ZN(new_n10374_));
  OAI22_X1   g10292(.A1(new_n1973_), .A2(new_n4468_), .B1(new_n4501_), .B2(new_n4902_), .ZN(new_n10375_));
  OAI21_X1   g10293(.A1(new_n4516_), .A2(new_n1239_), .B(new_n10375_), .ZN(new_n10376_));
  AOI21_X1   g10294(.A1(new_n10376_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n10377_));
  XOR2_X1    g10295(.A1(new_n4524_), .A2(new_n10377_), .Z(new_n10378_));
  AND2_X2    g10296(.A1(new_n10374_), .A2(new_n10378_), .Z(new_n10379_));
  NOR2_X1    g10297(.A1(new_n10374_), .A2(new_n10378_), .ZN(new_n10380_));
  OAI22_X1   g10298(.A1(new_n10379_), .A2(new_n10380_), .B1(new_n10320_), .B2(new_n10368_), .ZN(new_n10381_));
  NOR2_X1    g10299(.A1(new_n10368_), .A2(new_n10320_), .ZN(new_n10382_));
  XOR2_X1    g10300(.A1(new_n10374_), .A2(new_n10378_), .Z(new_n10383_));
  NAND2_X1   g10301(.A1(new_n10383_), .A2(new_n10382_), .ZN(new_n10384_));
  INV_X1     g10302(.I(new_n10331_), .ZN(new_n10385_));
  AOI21_X1   g10303(.A1(new_n10385_), .A2(new_n10335_), .B(new_n10332_), .ZN(new_n10386_));
  NAND2_X1   g10304(.A1(new_n4563_), .A2(new_n4722_), .ZN(new_n10387_));
  NAND2_X1   g10305(.A1(new_n4564_), .A2(new_n4720_), .ZN(new_n10388_));
  AOI22_X1   g10306(.A1(new_n10388_), .A2(new_n10387_), .B1(new_n4717_), .B2(new_n4564_), .ZN(new_n10389_));
  OAI21_X1   g10307(.A1(new_n10389_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n10390_));
  XOR2_X1    g10308(.A1(new_n4609_), .A2(new_n10390_), .Z(new_n10391_));
  AND2_X2    g10309(.A1(new_n10386_), .A2(new_n10391_), .Z(new_n10392_));
  INV_X1     g10310(.I(new_n10392_), .ZN(new_n10393_));
  NOR2_X1    g10311(.A1(new_n10386_), .A2(new_n10391_), .ZN(new_n10394_));
  INV_X1     g10312(.I(new_n10394_), .ZN(new_n10395_));
  AOI22_X1   g10313(.A1(new_n10393_), .A2(new_n10395_), .B1(new_n10381_), .B2(new_n10384_), .ZN(new_n10396_));
  NAND2_X1   g10314(.A1(new_n10384_), .A2(new_n10381_), .ZN(new_n10397_));
  XNOR2_X1   g10315(.A1(new_n10386_), .A2(new_n10391_), .ZN(new_n10398_));
  NOR2_X1    g10316(.A1(new_n10398_), .A2(new_n10397_), .ZN(new_n10399_));
  NOR3_X1    g10317(.A1(new_n10396_), .A2(new_n443_), .A3(new_n10399_), .ZN(new_n10400_));
  NOR2_X1    g10318(.A1(new_n10396_), .A2(new_n10399_), .ZN(new_n10401_));
  NOR2_X1    g10319(.A1(new_n10401_), .A2(new_n568_), .ZN(new_n10402_));
  NOR2_X1    g10320(.A1(new_n10402_), .A2(new_n10400_), .ZN(new_n10403_));
  NOR2_X1    g10321(.A1(new_n10403_), .A2(new_n10367_), .ZN(new_n10404_));
  INV_X1     g10322(.I(new_n10367_), .ZN(new_n10405_));
  XOR2_X1    g10323(.A1(new_n10401_), .A2(new_n443_), .Z(new_n10406_));
  NOR2_X1    g10324(.A1(new_n10406_), .A2(new_n10405_), .ZN(new_n10407_));
  OAI21_X1   g10325(.A1(new_n10344_), .A2(new_n10350_), .B(new_n10352_), .ZN(new_n10408_));
  NOR3_X1    g10326(.A1(new_n10407_), .A2(new_n10408_), .A3(new_n10404_), .ZN(new_n10409_));
  NOR2_X1    g10327(.A1(new_n10407_), .A2(new_n10404_), .ZN(new_n10410_));
  INV_X1     g10328(.I(new_n10408_), .ZN(new_n10411_));
  NOR2_X1    g10329(.A1(new_n10410_), .A2(new_n10411_), .ZN(new_n10412_));
  INV_X1     g10330(.I(new_n10412_), .ZN(new_n10413_));
  OAI21_X1   g10331(.A1(new_n10363_), .A2(new_n10409_), .B(new_n10413_), .ZN(new_n10414_));
  AOI21_X1   g10332(.A1(new_n10393_), .A2(new_n10397_), .B(new_n10394_), .ZN(new_n10415_));
  NOR2_X1    g10333(.A1(new_n10379_), .A2(new_n10382_), .ZN(new_n10416_));
  NOR2_X1    g10334(.A1(new_n10416_), .A2(new_n10380_), .ZN(new_n10417_));
  XOR2_X1    g10335(.A1(new_n4970_), .A2(new_n4974_), .Z(new_n10418_));
  INV_X1     g10336(.I(new_n10418_), .ZN(new_n10419_));
  AOI21_X1   g10337(.A1(new_n4977_), .A2(new_n4978_), .B(new_n4922_), .ZN(new_n10420_));
  AOI21_X1   g10338(.A1(new_n10419_), .A2(new_n4922_), .B(new_n10420_), .ZN(new_n10421_));
  INV_X1     g10339(.I(new_n10421_), .ZN(new_n10422_));
  OAI22_X1   g10340(.A1(new_n5552_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n4563_), .ZN(new_n10423_));
  AOI21_X1   g10341(.A1(new_n10423_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n10424_));
  XNOR2_X1   g10342(.A1(new_n4569_), .A2(new_n10424_), .ZN(new_n10425_));
  NOR2_X1    g10343(.A1(new_n10422_), .A2(new_n10425_), .ZN(new_n10426_));
  NAND2_X1   g10344(.A1(new_n10422_), .A2(new_n10425_), .ZN(new_n10427_));
  INV_X1     g10345(.I(new_n10427_), .ZN(new_n10428_));
  NOR2_X1    g10346(.A1(new_n10428_), .A2(new_n10426_), .ZN(new_n10429_));
  XNOR2_X1   g10347(.A1(new_n10429_), .A2(new_n10417_), .ZN(new_n10430_));
  NAND2_X1   g10348(.A1(new_n4722_), .A2(new_n4717_), .ZN(new_n10431_));
  OAI21_X1   g10349(.A1(new_n4720_), .A2(new_n10431_), .B(new_n4564_), .ZN(new_n10432_));
  OAI21_X1   g10350(.A1(new_n10432_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n10433_));
  XOR2_X1    g10351(.A1(new_n5001_), .A2(new_n10433_), .Z(new_n10434_));
  XOR2_X1    g10352(.A1(new_n10430_), .A2(new_n10434_), .Z(new_n10435_));
  NOR2_X1    g10353(.A1(new_n10435_), .A2(new_n10415_), .ZN(new_n10436_));
  INV_X1     g10354(.I(new_n10415_), .ZN(new_n10437_));
  INV_X1     g10355(.I(new_n10434_), .ZN(new_n10438_));
  NOR2_X1    g10356(.A1(new_n10430_), .A2(new_n10438_), .ZN(new_n10439_));
  INV_X1     g10357(.I(new_n10439_), .ZN(new_n10440_));
  NAND2_X1   g10358(.A1(new_n10430_), .A2(new_n10438_), .ZN(new_n10441_));
  AOI21_X1   g10359(.A1(new_n10440_), .A2(new_n10441_), .B(new_n10437_), .ZN(new_n10442_));
  NOR2_X1    g10360(.A1(new_n10436_), .A2(new_n10442_), .ZN(new_n10443_));
  INV_X1     g10361(.I(new_n10400_), .ZN(new_n10444_));
  AOI21_X1   g10362(.A1(new_n10444_), .A2(new_n10405_), .B(new_n10402_), .ZN(new_n10445_));
  INV_X1     g10363(.I(new_n10445_), .ZN(new_n10446_));
  NOR2_X1    g10364(.A1(new_n10443_), .A2(new_n10446_), .ZN(new_n10447_));
  INV_X1     g10365(.I(new_n10447_), .ZN(new_n10448_));
  NOR3_X1    g10366(.A1(new_n10436_), .A2(new_n10442_), .A3(new_n10445_), .ZN(new_n10449_));
  AOI21_X1   g10367(.A1(new_n10414_), .A2(new_n10448_), .B(new_n10449_), .ZN(new_n10450_));
  OAI21_X1   g10368(.A1(new_n10415_), .A2(new_n10439_), .B(new_n10441_), .ZN(new_n10451_));
  OAI21_X1   g10369(.A1(new_n4985_), .A2(new_n4987_), .B(new_n4917_), .ZN(new_n10452_));
  XOR2_X1    g10370(.A1(new_n4980_), .A2(new_n4984_), .Z(new_n10453_));
  NAND2_X1   g10371(.A1(new_n10453_), .A2(new_n4918_), .ZN(new_n10454_));
  NAND2_X1   g10372(.A1(new_n10454_), .A2(new_n10452_), .ZN(new_n10455_));
  INV_X1     g10373(.I(new_n10455_), .ZN(new_n10456_));
  NAND2_X1   g10374(.A1(new_n10429_), .A2(new_n10417_), .ZN(new_n10457_));
  NOR2_X1    g10375(.A1(new_n10457_), .A2(new_n10456_), .ZN(new_n10458_));
  NAND2_X1   g10376(.A1(new_n10457_), .A2(new_n10456_), .ZN(new_n10459_));
  NAND3_X1   g10377(.A1(new_n4563_), .A2(new_n4717_), .A3(new_n4719_), .ZN(new_n10460_));
  AOI21_X1   g10378(.A1(new_n10460_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n10461_));
  XNOR2_X1   g10379(.A1(new_n4610_), .A2(new_n10461_), .ZN(new_n10462_));
  NOR2_X1    g10380(.A1(new_n10427_), .A2(new_n10462_), .ZN(new_n10463_));
  AOI21_X1   g10381(.A1(new_n10459_), .A2(new_n10463_), .B(new_n10458_), .ZN(new_n10464_));
  NOR2_X1    g10382(.A1(new_n4990_), .A2(new_n4992_), .ZN(new_n10465_));
  NOR2_X1    g10383(.A1(new_n10465_), .A2(new_n4914_), .ZN(new_n10466_));
  XOR2_X1    g10384(.A1(new_n4988_), .A2(new_n273_), .Z(new_n10467_));
  AOI21_X1   g10385(.A1(new_n4914_), .A2(new_n10467_), .B(new_n10466_), .ZN(new_n10468_));
  XNOR2_X1   g10386(.A1(new_n10468_), .A2(new_n10464_), .ZN(new_n10469_));
  INV_X1     g10387(.I(new_n10469_), .ZN(new_n10470_));
  NOR2_X1    g10388(.A1(new_n10470_), .A2(new_n10451_), .ZN(new_n10471_));
  NOR2_X1    g10389(.A1(new_n10456_), .A2(new_n10462_), .ZN(new_n10472_));
  XOR2_X1    g10390(.A1(new_n10472_), .A2(new_n10457_), .Z(new_n10473_));
  NOR2_X1    g10391(.A1(new_n10473_), .A2(new_n10428_), .ZN(new_n10474_));
  NAND2_X1   g10392(.A1(new_n10473_), .A2(new_n10428_), .ZN(new_n10475_));
  INV_X1     g10393(.I(new_n10475_), .ZN(new_n10476_));
  NOR2_X1    g10394(.A1(new_n10476_), .A2(new_n10474_), .ZN(new_n10477_));
  NAND2_X1   g10395(.A1(new_n10470_), .A2(new_n10451_), .ZN(new_n10478_));
  AOI21_X1   g10396(.A1(new_n10477_), .A2(new_n10478_), .B(new_n10471_), .ZN(new_n10479_));
  INV_X1     g10397(.I(new_n10479_), .ZN(new_n10480_));
  NAND2_X1   g10398(.A1(new_n10468_), .A2(new_n10464_), .ZN(new_n10481_));
  AOI21_X1   g10399(.A1(new_n4993_), .A2(new_n5014_), .B(new_n10481_), .ZN(new_n10482_));
  INV_X1     g10400(.I(new_n10482_), .ZN(new_n10483_));
  NOR3_X1    g10401(.A1(new_n10450_), .A2(new_n10480_), .A3(new_n10483_), .ZN(new_n10484_));
  INV_X1     g10402(.I(new_n5010_), .ZN(new_n10485_));
  AOI21_X1   g10403(.A1(new_n10485_), .A2(new_n5009_), .B(new_n5011_), .ZN(new_n10486_));
  XOR2_X1    g10404(.A1(new_n4805_), .A2(new_n4850_), .Z(new_n10487_));
  OAI21_X1   g10405(.A1(new_n4846_), .A2(new_n4849_), .B(new_n4810_), .ZN(new_n10488_));
  XOR2_X1    g10406(.A1(new_n4841_), .A2(new_n4844_), .Z(new_n10489_));
  OAI21_X1   g10407(.A1(new_n4810_), .A2(new_n10489_), .B(new_n10488_), .ZN(new_n10490_));
  NOR2_X1    g10408(.A1(new_n10487_), .A2(new_n10486_), .ZN(new_n10491_));
  NOR2_X1    g10409(.A1(new_n10491_), .A2(new_n10490_), .ZN(new_n10492_));
  AOI21_X1   g10410(.A1(new_n10486_), .A2(new_n10487_), .B(new_n10492_), .ZN(new_n10493_));
  OAI21_X1   g10411(.A1(new_n10484_), .A2(new_n5015_), .B(new_n10493_), .ZN(new_n10494_));
  INV_X1     g10412(.I(new_n4792_), .ZN(new_n10495_));
  AOI21_X1   g10413(.A1(new_n10495_), .A2(new_n4780_), .B(new_n4793_), .ZN(new_n10496_));
  OAI22_X1   g10414(.A1(new_n4765_), .A2(new_n4767_), .B1(new_n4563_), .B2(new_n4612_), .ZN(new_n10497_));
  AOI21_X1   g10415(.A1(new_n10497_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n10498_));
  XNOR2_X1   g10416(.A1(new_n5001_), .A2(new_n10498_), .ZN(new_n10499_));
  INV_X1     g10417(.I(new_n10499_), .ZN(new_n10500_));
  INV_X1     g10418(.I(new_n4576_), .ZN(new_n10501_));
  AOI21_X1   g10419(.A1(new_n10501_), .A2(new_n4575_), .B(new_n4491_), .ZN(new_n10502_));
  XNOR2_X1   g10420(.A1(new_n4554_), .A2(new_n4574_), .ZN(new_n10503_));
  NOR2_X1    g10421(.A1(new_n10503_), .A2(new_n4492_), .ZN(new_n10504_));
  NOR3_X1    g10422(.A1(new_n10504_), .A2(new_n10500_), .A3(new_n10502_), .ZN(new_n10505_));
  NOR2_X1    g10423(.A1(new_n10504_), .A2(new_n10502_), .ZN(new_n10506_));
  NOR2_X1    g10424(.A1(new_n10506_), .A2(new_n10499_), .ZN(new_n10507_));
  NOR2_X1    g10425(.A1(new_n10507_), .A2(new_n10505_), .ZN(new_n10508_));
  NOR2_X1    g10426(.A1(new_n10508_), .A2(new_n10496_), .ZN(new_n10509_));
  INV_X1     g10427(.I(new_n10496_), .ZN(new_n10510_));
  XOR2_X1    g10428(.A1(new_n10506_), .A2(new_n10500_), .Z(new_n10511_));
  NOR2_X1    g10429(.A1(new_n10511_), .A2(new_n10510_), .ZN(new_n10512_));
  NOR2_X1    g10430(.A1(new_n10512_), .A2(new_n10509_), .ZN(new_n10513_));
  AOI21_X1   g10431(.A1(new_n4851_), .A2(new_n4801_), .B(new_n10513_), .ZN(new_n10514_));
  INV_X1     g10432(.I(new_n10514_), .ZN(new_n10515_));
  OAI21_X1   g10433(.A1(new_n10494_), .A2(new_n10515_), .B(new_n4853_), .ZN(new_n10516_));
  INV_X1     g10434(.I(new_n4577_), .ZN(new_n10517_));
  OAI21_X1   g10435(.A1(new_n4618_), .A2(new_n4620_), .B(new_n10517_), .ZN(new_n10518_));
  XOR2_X1    g10436(.A1(new_n4605_), .A2(new_n4617_), .Z(new_n10519_));
  OAI21_X1   g10437(.A1(new_n10517_), .A2(new_n10519_), .B(new_n10518_), .ZN(new_n10520_));
  NOR2_X1    g10438(.A1(new_n10505_), .A2(new_n10496_), .ZN(new_n10521_));
  NOR2_X1    g10439(.A1(new_n10521_), .A2(new_n10507_), .ZN(new_n10522_));
  INV_X1     g10440(.I(new_n10522_), .ZN(new_n10523_));
  NOR2_X1    g10441(.A1(new_n10523_), .A2(new_n10520_), .ZN(new_n10524_));
  INV_X1     g10442(.I(new_n10524_), .ZN(new_n10525_));
  NAND2_X1   g10443(.A1(new_n10523_), .A2(new_n10520_), .ZN(new_n10526_));
  XNOR2_X1   g10444(.A1(new_n4647_), .A2(new_n4621_), .ZN(new_n10527_));
  NAND2_X1   g10445(.A1(new_n10525_), .A2(new_n10526_), .ZN(new_n10528_));
  NAND2_X1   g10446(.A1(new_n10516_), .A2(new_n10528_), .ZN(new_n10529_));
  INV_X1     g10447(.I(new_n4632_), .ZN(new_n10530_));
  AOI21_X1   g10448(.A1(new_n4631_), .A2(new_n10530_), .B(new_n4634_), .ZN(new_n10531_));
  OAI22_X1   g10449(.A1(new_n4596_), .A2(new_n4526_), .B1(new_n4529_), .B2(new_n4563_), .ZN(new_n10532_));
  AOI21_X1   g10450(.A1(new_n10532_), .A2(new_n72_), .B(new_n79_), .ZN(new_n10533_));
  XNOR2_X1   g10451(.A1(new_n5001_), .A2(new_n10533_), .ZN(new_n10534_));
  NAND2_X1   g10452(.A1(new_n4518_), .A2(new_n87_), .ZN(new_n10535_));
  AOI22_X1   g10453(.A1(new_n4564_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n4555_), .ZN(new_n10536_));
  AOI21_X1   g10454(.A1(new_n10535_), .A2(new_n10536_), .B(new_n82_), .ZN(new_n10537_));
  NAND2_X1   g10455(.A1(new_n4569_), .A2(new_n10537_), .ZN(new_n10538_));
  NOR3_X1    g10456(.A1(new_n4613_), .A2(new_n117_), .A3(new_n4767_), .ZN(new_n10539_));
  XOR2_X1    g10457(.A1(new_n10539_), .A2(new_n65_), .Z(new_n10540_));
  INV_X1     g10458(.I(new_n10540_), .ZN(new_n10541_));
  NOR2_X1    g10459(.A1(new_n10538_), .A2(new_n10541_), .ZN(new_n10542_));
  INV_X1     g10460(.I(new_n10542_), .ZN(new_n10543_));
  NAND2_X1   g10461(.A1(new_n10538_), .A2(new_n10541_), .ZN(new_n10544_));
  AOI21_X1   g10462(.A1(new_n10543_), .A2(new_n10544_), .B(new_n4628_), .ZN(new_n10545_));
  XOR2_X1    g10463(.A1(new_n10538_), .A2(new_n10540_), .Z(new_n10546_));
  NOR2_X1    g10464(.A1(new_n10546_), .A2(new_n4633_), .ZN(new_n10547_));
  NOR2_X1    g10465(.A1(new_n10547_), .A2(new_n10545_), .ZN(new_n10548_));
  XNOR2_X1   g10466(.A1(new_n10548_), .A2(new_n10534_), .ZN(new_n10549_));
  NOR2_X1    g10467(.A1(new_n10549_), .A2(new_n10531_), .ZN(new_n10550_));
  INV_X1     g10468(.I(new_n10531_), .ZN(new_n10551_));
  AND2_X2    g10469(.A1(new_n10548_), .A2(new_n10534_), .Z(new_n10552_));
  NOR2_X1    g10470(.A1(new_n10548_), .A2(new_n10534_), .ZN(new_n10553_));
  NOR2_X1    g10471(.A1(new_n10552_), .A2(new_n10553_), .ZN(new_n10554_));
  NOR2_X1    g10472(.A1(new_n10551_), .A2(new_n10554_), .ZN(new_n10555_));
  NOR2_X1    g10473(.A1(new_n10555_), .A2(new_n10550_), .ZN(new_n10556_));
  NOR2_X1    g10474(.A1(new_n4638_), .A2(new_n4643_), .ZN(new_n10557_));
  NOR2_X1    g10475(.A1(new_n10557_), .A2(new_n4644_), .ZN(new_n10558_));
  NOR2_X1    g10476(.A1(new_n10558_), .A2(new_n10556_), .ZN(new_n10559_));
  XOR2_X1    g10477(.A1(new_n10529_), .A2(new_n10559_), .Z(new_n10560_));
  NOR2_X1    g10478(.A1(new_n10560_), .A2(new_n4649_), .ZN(new_n10561_));
  NAND2_X1   g10479(.A1(new_n10560_), .A2(new_n4649_), .ZN(new_n10562_));
  INV_X1     g10480(.I(new_n10562_), .ZN(new_n10563_));
  NOR2_X1    g10481(.A1(new_n10563_), .A2(new_n10561_), .ZN(new_n10564_));
  INV_X1     g10482(.I(new_n10516_), .ZN(new_n10565_));
  OAI21_X1   g10483(.A1(new_n10527_), .A2(new_n10526_), .B(new_n10525_), .ZN(new_n10566_));
  NAND2_X1   g10484(.A1(new_n10565_), .A2(new_n10566_), .ZN(new_n10567_));
  INV_X1     g10485(.I(new_n10567_), .ZN(new_n10568_));
  NOR2_X1    g10486(.A1(new_n10565_), .A2(new_n10566_), .ZN(new_n10569_));
  NOR2_X1    g10487(.A1(new_n10568_), .A2(new_n10569_), .ZN(new_n10570_));
  INV_X1     g10488(.I(new_n10570_), .ZN(new_n10571_));
  NOR2_X1    g10489(.A1(new_n10513_), .A2(new_n4801_), .ZN(new_n10572_));
  XNOR2_X1   g10490(.A1(new_n10494_), .A2(new_n10572_), .ZN(new_n10573_));
  NAND2_X1   g10491(.A1(new_n10573_), .A2(new_n4851_), .ZN(new_n10574_));
  INV_X1     g10492(.I(new_n10574_), .ZN(new_n10575_));
  NOR2_X1    g10493(.A1(new_n10573_), .A2(new_n4851_), .ZN(new_n10576_));
  NOR2_X1    g10494(.A1(new_n10575_), .A2(new_n10576_), .ZN(new_n10577_));
  NOR2_X1    g10495(.A1(new_n10450_), .A2(new_n10480_), .ZN(new_n10578_));
  XOR2_X1    g10496(.A1(new_n10578_), .A2(new_n5015_), .Z(new_n10579_));
  NAND2_X1   g10497(.A1(new_n10579_), .A2(new_n10481_), .ZN(new_n10580_));
  INV_X1     g10498(.I(new_n10580_), .ZN(new_n10581_));
  NOR2_X1    g10499(.A1(new_n10579_), .A2(new_n10481_), .ZN(new_n10582_));
  NOR2_X1    g10500(.A1(new_n10581_), .A2(new_n10582_), .ZN(new_n10583_));
  INV_X1     g10501(.I(new_n10583_), .ZN(new_n10584_));
  XOR2_X1    g10502(.A1(new_n10443_), .A2(new_n10446_), .Z(new_n10585_));
  AND2_X2    g10503(.A1(new_n10414_), .A2(new_n10585_), .Z(new_n10586_));
  NOR2_X1    g10504(.A1(new_n10447_), .A2(new_n10449_), .ZN(new_n10587_));
  NOR2_X1    g10505(.A1(new_n10414_), .A2(new_n10587_), .ZN(new_n10588_));
  NOR2_X1    g10506(.A1(new_n10586_), .A2(new_n10588_), .ZN(new_n10589_));
  XOR2_X1    g10507(.A1(new_n10410_), .A2(new_n10408_), .Z(new_n10590_));
  NOR2_X1    g10508(.A1(new_n10363_), .A2(new_n10590_), .ZN(new_n10591_));
  INV_X1     g10509(.I(new_n10363_), .ZN(new_n10592_));
  NOR2_X1    g10510(.A1(new_n10412_), .A2(new_n10409_), .ZN(new_n10593_));
  NOR2_X1    g10511(.A1(new_n10592_), .A2(new_n10593_), .ZN(new_n10594_));
  NOR2_X1    g10512(.A1(new_n10594_), .A2(new_n10591_), .ZN(new_n10595_));
  XNOR2_X1   g10513(.A1(new_n10357_), .A2(new_n10305_), .ZN(new_n10596_));
  AND2_X2    g10514(.A1(new_n10304_), .A2(new_n10596_), .Z(new_n10597_));
  AOI21_X1   g10515(.A1(new_n10360_), .A2(new_n10361_), .B(new_n10304_), .ZN(new_n10598_));
  NOR2_X1    g10516(.A1(new_n10597_), .A2(new_n10598_), .ZN(new_n10599_));
  INV_X1     g10517(.I(new_n10599_), .ZN(new_n10600_));
  INV_X1     g10518(.I(new_n10301_), .ZN(new_n10601_));
  XOR2_X1    g10519(.A1(new_n10300_), .A2(new_n5578_), .Z(new_n10602_));
  NOR2_X1    g10520(.A1(new_n10602_), .A2(new_n10601_), .ZN(new_n10603_));
  NAND2_X1   g10521(.A1(new_n10602_), .A2(new_n10601_), .ZN(new_n10604_));
  INV_X1     g10522(.I(new_n10604_), .ZN(new_n10605_));
  NOR2_X1    g10523(.A1(new_n10605_), .A2(new_n10603_), .ZN(new_n10606_));
  AND2_X2    g10524(.A1(new_n10291_), .A2(new_n10292_), .Z(new_n10607_));
  NOR2_X1    g10525(.A1(new_n10271_), .A2(new_n10607_), .ZN(new_n10608_));
  INV_X1     g10526(.I(new_n10607_), .ZN(new_n10609_));
  NOR2_X1    g10527(.A1(new_n10270_), .A2(new_n10609_), .ZN(new_n10610_));
  NOR2_X1    g10528(.A1(new_n10608_), .A2(new_n10610_), .ZN(new_n10611_));
  INV_X1     g10529(.I(new_n10611_), .ZN(new_n10612_));
  INV_X1     g10530(.I(new_n10267_), .ZN(new_n10613_));
  NOR2_X1    g10531(.A1(new_n10236_), .A2(new_n10266_), .ZN(new_n10614_));
  XNOR2_X1   g10532(.A1(new_n10614_), .A2(new_n6038_), .ZN(new_n10615_));
  NOR2_X1    g10533(.A1(new_n10615_), .A2(new_n10613_), .ZN(new_n10616_));
  NAND2_X1   g10534(.A1(new_n10615_), .A2(new_n10613_), .ZN(new_n10617_));
  INV_X1     g10535(.I(new_n10617_), .ZN(new_n10618_));
  NOR2_X1    g10536(.A1(new_n10618_), .A2(new_n10616_), .ZN(new_n10619_));
  INV_X1     g10537(.I(new_n10619_), .ZN(new_n10620_));
  XOR2_X1    g10538(.A1(new_n10233_), .A2(new_n6828_), .Z(new_n10621_));
  NAND2_X1   g10539(.A1(new_n10621_), .A2(new_n10234_), .ZN(new_n10622_));
  NOR2_X1    g10540(.A1(new_n10621_), .A2(new_n10234_), .ZN(new_n10623_));
  INV_X1     g10541(.I(new_n10623_), .ZN(new_n10624_));
  NAND2_X1   g10542(.A1(new_n10624_), .A2(new_n10622_), .ZN(new_n10625_));
  XOR2_X1    g10543(.A1(new_n10196_), .A2(new_n7873_), .Z(new_n10626_));
  NAND2_X1   g10544(.A1(new_n10626_), .A2(new_n10199_), .ZN(new_n10627_));
  XNOR2_X1   g10545(.A1(new_n10196_), .A2(new_n7873_), .ZN(new_n10628_));
  NAND2_X1   g10546(.A1(new_n10628_), .A2(new_n10198_), .ZN(new_n10629_));
  NAND2_X1   g10547(.A1(new_n10629_), .A2(new_n10627_), .ZN(new_n10630_));
  INV_X1     g10548(.I(new_n10630_), .ZN(new_n10631_));
  NAND2_X1   g10549(.A1(new_n10185_), .A2(new_n10187_), .ZN(new_n10632_));
  XOR2_X1    g10550(.A1(new_n10632_), .A2(new_n10195_), .Z(new_n10633_));
  NOR2_X1    g10551(.A1(new_n10160_), .A2(new_n10150_), .ZN(new_n10634_));
  XOR2_X1    g10552(.A1(new_n10181_), .A2(new_n10182_), .Z(new_n10635_));
  NAND2_X1   g10553(.A1(new_n10187_), .A2(new_n10184_), .ZN(new_n10636_));
  NAND2_X1   g10554(.A1(new_n10634_), .A2(new_n10636_), .ZN(new_n10637_));
  OAI21_X1   g10555(.A1(new_n10634_), .A2(new_n10635_), .B(new_n10637_), .ZN(new_n10638_));
  AOI22_X1   g10556(.A1(new_n8811_), .A2(new_n8808_), .B1(new_n10155_), .B2(new_n10157_), .ZN(new_n10639_));
  NAND2_X1   g10557(.A1(new_n10149_), .A2(new_n10639_), .ZN(new_n10640_));
  NOR2_X1    g10558(.A1(new_n10149_), .A2(new_n10639_), .ZN(new_n10641_));
  INV_X1     g10559(.I(new_n10641_), .ZN(new_n10642_));
  AOI21_X1   g10560(.A1(new_n10642_), .A2(new_n10640_), .B(new_n10154_), .ZN(new_n10643_));
  INV_X1     g10561(.I(new_n10640_), .ZN(new_n10644_));
  NOR3_X1    g10562(.A1(new_n10644_), .A2(new_n10153_), .A3(new_n10641_), .ZN(new_n10645_));
  NOR2_X1    g10563(.A1(new_n10643_), .A2(new_n10645_), .ZN(new_n10646_));
  NOR2_X1    g10564(.A1(new_n10140_), .A2(new_n10136_), .ZN(new_n10647_));
  NOR2_X1    g10565(.A1(new_n10145_), .A2(new_n10146_), .ZN(new_n10648_));
  MUX2_X1    g10566(.I0(new_n10648_), .I1(new_n10647_), .S(new_n10131_), .Z(new_n10649_));
  NAND3_X1   g10567(.A1(new_n10111_), .A2(new_n10649_), .A3(new_n10114_), .ZN(new_n10650_));
  OAI21_X1   g10568(.A1(new_n10110_), .A2(new_n10113_), .B(new_n10148_), .ZN(new_n10651_));
  NAND2_X1   g10569(.A1(new_n10650_), .A2(new_n10651_), .ZN(new_n10652_));
  NAND2_X1   g10570(.A1(new_n10082_), .A2(new_n10075_), .ZN(new_n10653_));
  NOR3_X1    g10571(.A1(new_n10112_), .A2(new_n10100_), .A3(new_n10108_), .ZN(new_n10654_));
  AOI21_X1   g10572(.A1(new_n10101_), .A2(new_n10105_), .B(new_n10107_), .ZN(new_n10655_));
  NOR2_X1    g10573(.A1(new_n10654_), .A2(new_n10655_), .ZN(new_n10656_));
  NOR2_X1    g10574(.A1(new_n10113_), .A2(new_n10109_), .ZN(new_n10657_));
  MUX2_X1    g10575(.I0(new_n10657_), .I1(new_n10656_), .S(new_n10653_), .Z(new_n10658_));
  NOR2_X1    g10576(.A1(new_n10076_), .A2(new_n10065_), .ZN(new_n10659_));
  NAND2_X1   g10577(.A1(new_n10038_), .A2(new_n10030_), .ZN(new_n10660_));
  INV_X1     g10578(.I(new_n10073_), .ZN(new_n10661_));
  NAND2_X1   g10579(.A1(new_n10660_), .A2(new_n10661_), .ZN(new_n10662_));
  INV_X1     g10580(.I(new_n10080_), .ZN(new_n10663_));
  OAI21_X1   g10581(.A1(new_n9356_), .A2(new_n9359_), .B(new_n10663_), .ZN(new_n10664_));
  INV_X1     g10582(.I(new_n10664_), .ZN(new_n10665_));
  NAND2_X1   g10583(.A1(new_n10662_), .A2(new_n10665_), .ZN(new_n10666_));
  NAND2_X1   g10584(.A1(new_n10074_), .A2(new_n10664_), .ZN(new_n10667_));
  AOI21_X1   g10585(.A1(new_n10666_), .A2(new_n10667_), .B(new_n10659_), .ZN(new_n10668_));
  NOR2_X1    g10586(.A1(new_n10074_), .A2(new_n10664_), .ZN(new_n10669_));
  NOR2_X1    g10587(.A1(new_n10662_), .A2(new_n10665_), .ZN(new_n10670_));
  NOR4_X1    g10588(.A1(new_n10670_), .A2(new_n10076_), .A3(new_n10065_), .A4(new_n10669_), .ZN(new_n10671_));
  NOR2_X1    g10589(.A1(new_n10671_), .A2(new_n10668_), .ZN(new_n10672_));
  NAND2_X1   g10590(.A1(new_n10066_), .A2(new_n10062_), .ZN(new_n10673_));
  NOR2_X1    g10591(.A1(new_n10047_), .A2(new_n10070_), .ZN(new_n10674_));
  INV_X1     g10592(.I(new_n10674_), .ZN(new_n10675_));
  OAI21_X1   g10593(.A1(new_n10045_), .A2(new_n10046_), .B(new_n10070_), .ZN(new_n10676_));
  INV_X1     g10594(.I(new_n10046_), .ZN(new_n10677_));
  NAND3_X1   g10595(.A1(new_n10677_), .A2(new_n10044_), .A3(new_n10071_), .ZN(new_n10678_));
  NAND2_X1   g10596(.A1(new_n10678_), .A2(new_n10676_), .ZN(new_n10679_));
  NAND3_X1   g10597(.A1(new_n10673_), .A2(new_n10675_), .A3(new_n10679_), .ZN(new_n10680_));
  NOR3_X1    g10598(.A1(new_n10064_), .A2(new_n10063_), .A3(new_n10065_), .ZN(new_n10681_));
  AOI21_X1   g10599(.A1(new_n10056_), .A2(new_n10059_), .B(new_n10061_), .ZN(new_n10682_));
  OAI21_X1   g10600(.A1(new_n10681_), .A2(new_n10682_), .B(new_n10679_), .ZN(new_n10683_));
  NAND2_X1   g10601(.A1(new_n10683_), .A2(new_n10674_), .ZN(new_n10684_));
  NAND2_X1   g10602(.A1(new_n10684_), .A2(new_n10680_), .ZN(new_n10685_));
  NAND3_X1   g10603(.A1(new_n10685_), .A2(new_n10030_), .A3(new_n10038_), .ZN(new_n10686_));
  NOR2_X1    g10604(.A1(new_n10683_), .A2(new_n10674_), .ZN(new_n10687_));
  AOI21_X1   g10605(.A1(new_n10673_), .A2(new_n10679_), .B(new_n10675_), .ZN(new_n10688_));
  NOR2_X1    g10606(.A1(new_n10687_), .A2(new_n10688_), .ZN(new_n10689_));
  NAND2_X1   g10607(.A1(new_n10689_), .A2(new_n10660_), .ZN(new_n10690_));
  NAND2_X1   g10608(.A1(new_n10690_), .A2(new_n10686_), .ZN(new_n10691_));
  NAND2_X1   g10609(.A1(new_n10047_), .A2(new_n10070_), .ZN(new_n10692_));
  AOI22_X1   g10610(.A1(new_n10038_), .A2(new_n10030_), .B1(new_n10675_), .B2(new_n10692_), .ZN(new_n10693_));
  NAND3_X1   g10611(.A1(new_n10038_), .A2(new_n10030_), .A3(new_n10679_), .ZN(new_n10694_));
  INV_X1     g10612(.I(new_n10694_), .ZN(new_n10695_));
  NOR2_X1    g10613(.A1(new_n10695_), .A2(new_n10693_), .ZN(new_n10696_));
  INV_X1     g10614(.I(new_n10032_), .ZN(new_n10697_));
  NAND2_X1   g10615(.A1(new_n9362_), .A2(new_n10035_), .ZN(new_n10698_));
  INV_X1     g10616(.I(new_n10698_), .ZN(new_n10699_));
  OAI21_X1   g10617(.A1(new_n9985_), .A2(new_n10028_), .B(new_n10699_), .ZN(new_n10700_));
  INV_X1     g10618(.I(new_n9382_), .ZN(new_n10701_));
  NAND3_X1   g10619(.A1(new_n9903_), .A2(new_n9888_), .A3(new_n9906_), .ZN(new_n10702_));
  AOI21_X1   g10620(.A1(new_n10702_), .A2(new_n9940_), .B(new_n9907_), .ZN(new_n10703_));
  AOI21_X1   g10621(.A1(new_n10703_), .A2(new_n9917_), .B(new_n9929_), .ZN(new_n10704_));
  INV_X1     g10622(.I(new_n9936_), .ZN(new_n10705_));
  OAI21_X1   g10623(.A1(new_n10704_), .A2(new_n9942_), .B(new_n10705_), .ZN(new_n10706_));
  NOR3_X1    g10624(.A1(new_n9913_), .A2(new_n9907_), .A3(new_n9918_), .ZN(new_n10707_));
  OAI21_X1   g10625(.A1(new_n10707_), .A2(new_n9929_), .B(new_n9919_), .ZN(new_n10708_));
  INV_X1     g10626(.I(new_n9949_), .ZN(new_n10709_));
  OAI21_X1   g10627(.A1(new_n10708_), .A2(new_n10705_), .B(new_n10709_), .ZN(new_n10710_));
  NAND3_X1   g10628(.A1(new_n9967_), .A2(new_n9959_), .A3(new_n9968_), .ZN(new_n10711_));
  NAND3_X1   g10629(.A1(new_n9978_), .A2(new_n10711_), .A3(new_n9954_), .ZN(new_n10712_));
  INV_X1     g10630(.I(new_n9973_), .ZN(new_n10713_));
  AOI21_X1   g10631(.A1(new_n9978_), .A2(new_n10711_), .B(new_n9954_), .ZN(new_n10714_));
  OAI21_X1   g10632(.A1(new_n10713_), .A2(new_n10714_), .B(new_n10712_), .ZN(new_n10715_));
  AOI21_X1   g10633(.A1(new_n10710_), .A2(new_n10706_), .B(new_n10715_), .ZN(new_n10716_));
  NAND2_X1   g10634(.A1(new_n10716_), .A2(new_n10701_), .ZN(new_n10717_));
  OAI21_X1   g10635(.A1(new_n10716_), .A2(new_n10701_), .B(new_n9982_), .ZN(new_n10718_));
  NAND2_X1   g10636(.A1(new_n10718_), .A2(new_n10717_), .ZN(new_n10719_));
  NAND3_X1   g10637(.A1(new_n10719_), .A2(new_n10027_), .A3(new_n10698_), .ZN(new_n10720_));
  AOI21_X1   g10638(.A1(new_n10700_), .A2(new_n10720_), .B(new_n10697_), .ZN(new_n10721_));
  AOI21_X1   g10639(.A1(new_n10719_), .A2(new_n10027_), .B(new_n10698_), .ZN(new_n10722_));
  NOR3_X1    g10640(.A1(new_n9985_), .A2(new_n10028_), .A3(new_n10699_), .ZN(new_n10723_));
  NOR3_X1    g10641(.A1(new_n10723_), .A2(new_n10722_), .A3(new_n10032_), .ZN(new_n10724_));
  NOR2_X1    g10642(.A1(new_n10724_), .A2(new_n10721_), .ZN(new_n10725_));
  NOR2_X1    g10643(.A1(new_n9993_), .A2(new_n10025_), .ZN(new_n10726_));
  INV_X1     g10644(.I(new_n10726_), .ZN(new_n10727_));
  OAI21_X1   g10645(.A1(new_n9991_), .A2(new_n9992_), .B(new_n10025_), .ZN(new_n10728_));
  INV_X1     g10646(.I(new_n9992_), .ZN(new_n10729_));
  INV_X1     g10647(.I(new_n10022_), .ZN(new_n10730_));
  NAND2_X1   g10648(.A1(new_n10730_), .A2(new_n10023_), .ZN(new_n10731_));
  NAND3_X1   g10649(.A1(new_n10731_), .A2(new_n10729_), .A3(new_n9990_), .ZN(new_n10732_));
  NAND2_X1   g10650(.A1(new_n10728_), .A2(new_n10732_), .ZN(new_n10733_));
  NAND3_X1   g10651(.A1(new_n10018_), .A2(new_n10727_), .A3(new_n10733_), .ZN(new_n10734_));
  NOR3_X1    g10652(.A1(new_n10014_), .A2(new_n10015_), .A3(new_n10016_), .ZN(new_n10735_));
  AOI21_X1   g10653(.A1(new_n10004_), .A2(new_n10007_), .B(new_n10012_), .ZN(new_n10736_));
  OAI21_X1   g10654(.A1(new_n10735_), .A2(new_n10736_), .B(new_n10733_), .ZN(new_n10737_));
  NAND2_X1   g10655(.A1(new_n10737_), .A2(new_n10726_), .ZN(new_n10738_));
  NAND2_X1   g10656(.A1(new_n10738_), .A2(new_n10734_), .ZN(new_n10739_));
  NAND3_X1   g10657(.A1(new_n10718_), .A2(new_n10717_), .A3(new_n10739_), .ZN(new_n10740_));
  NOR2_X1    g10658(.A1(new_n10737_), .A2(new_n10726_), .ZN(new_n10741_));
  AOI21_X1   g10659(.A1(new_n10018_), .A2(new_n10733_), .B(new_n10727_), .ZN(new_n10742_));
  NOR2_X1    g10660(.A1(new_n10741_), .A2(new_n10742_), .ZN(new_n10743_));
  OAI21_X1   g10661(.A1(new_n9984_), .A2(new_n9977_), .B(new_n10743_), .ZN(new_n10744_));
  NAND2_X1   g10662(.A1(new_n10744_), .A2(new_n10740_), .ZN(new_n10745_));
  NAND3_X1   g10663(.A1(new_n9931_), .A2(new_n9919_), .A3(new_n9936_), .ZN(new_n10746_));
  AOI21_X1   g10664(.A1(new_n10746_), .A2(new_n10709_), .B(new_n9937_), .ZN(new_n10747_));
  NAND2_X1   g10665(.A1(new_n9978_), .A2(new_n10711_), .ZN(new_n10748_));
  NAND2_X1   g10666(.A1(new_n9955_), .A2(new_n10713_), .ZN(new_n10749_));
  XOR2_X1    g10667(.A1(new_n9954_), .A2(new_n9973_), .Z(new_n10750_));
  NAND3_X1   g10668(.A1(new_n10748_), .A2(new_n10749_), .A3(new_n10750_), .ZN(new_n10751_));
  NAND2_X1   g10669(.A1(new_n10748_), .A2(new_n10750_), .ZN(new_n10752_));
  NAND3_X1   g10670(.A1(new_n10752_), .A2(new_n9955_), .A3(new_n10713_), .ZN(new_n10753_));
  NAND2_X1   g10671(.A1(new_n10753_), .A2(new_n10751_), .ZN(new_n10754_));
  XOR2_X1    g10672(.A1(new_n10754_), .A2(new_n10747_), .Z(new_n10755_));
  NAND2_X1   g10673(.A1(new_n9993_), .A2(new_n10025_), .ZN(new_n10756_));
  NAND2_X1   g10674(.A1(new_n10727_), .A2(new_n10756_), .ZN(new_n10757_));
  INV_X1     g10675(.I(new_n10757_), .ZN(new_n10758_));
  AOI21_X1   g10676(.A1(new_n10718_), .A2(new_n10717_), .B(new_n10758_), .ZN(new_n10759_));
  INV_X1     g10677(.I(new_n10733_), .ZN(new_n10760_));
  NOR3_X1    g10678(.A1(new_n9984_), .A2(new_n9977_), .A3(new_n10760_), .ZN(new_n10761_));
  NOR2_X1    g10679(.A1(new_n10761_), .A2(new_n10759_), .ZN(new_n10762_));
  NOR2_X1    g10680(.A1(new_n9382_), .A2(new_n9981_), .ZN(new_n10763_));
  OAI21_X1   g10681(.A1(new_n10747_), .A2(new_n10715_), .B(new_n10763_), .ZN(new_n10764_));
  NAND2_X1   g10682(.A1(new_n10710_), .A2(new_n10706_), .ZN(new_n10765_));
  INV_X1     g10683(.I(new_n10763_), .ZN(new_n10766_));
  NAND3_X1   g10684(.A1(new_n10765_), .A2(new_n9975_), .A3(new_n10766_), .ZN(new_n10767_));
  AOI21_X1   g10685(.A1(new_n10767_), .A2(new_n10764_), .B(new_n9969_), .ZN(new_n10768_));
  NOR2_X1    g10686(.A1(new_n10716_), .A2(new_n10766_), .ZN(new_n10769_));
  NOR3_X1    g10687(.A1(new_n10747_), .A2(new_n10715_), .A3(new_n10763_), .ZN(new_n10770_));
  NOR3_X1    g10688(.A1(new_n10769_), .A2(new_n10770_), .A3(new_n9978_), .ZN(new_n10771_));
  NOR2_X1    g10689(.A1(new_n10771_), .A2(new_n10768_), .ZN(new_n10772_));
  NOR3_X1    g10690(.A1(new_n10762_), .A2(new_n10745_), .A3(new_n10755_), .ZN(new_n10773_));
  INV_X1     g10691(.I(new_n10773_), .ZN(new_n10774_));
  NOR3_X1    g10692(.A1(new_n9984_), .A2(new_n9977_), .A3(new_n10743_), .ZN(new_n10775_));
  AOI21_X1   g10693(.A1(new_n10718_), .A2(new_n10717_), .B(new_n10739_), .ZN(new_n10776_));
  NOR2_X1    g10694(.A1(new_n10775_), .A2(new_n10776_), .ZN(new_n10777_));
  NAND2_X1   g10695(.A1(new_n10754_), .A2(new_n10747_), .ZN(new_n10778_));
  NAND3_X1   g10696(.A1(new_n10765_), .A2(new_n10751_), .A3(new_n10753_), .ZN(new_n10779_));
  NAND2_X1   g10697(.A1(new_n10779_), .A2(new_n10778_), .ZN(new_n10780_));
  OAI21_X1   g10698(.A1(new_n10769_), .A2(new_n10770_), .B(new_n9978_), .ZN(new_n10781_));
  NAND3_X1   g10699(.A1(new_n10767_), .A2(new_n10764_), .A3(new_n9969_), .ZN(new_n10782_));
  NAND2_X1   g10700(.A1(new_n10781_), .A2(new_n10782_), .ZN(new_n10783_));
  NAND3_X1   g10701(.A1(new_n10745_), .A2(new_n10783_), .A3(new_n10755_), .ZN(new_n10784_));
  OAI21_X1   g10702(.A1(new_n10777_), .A2(new_n10772_), .B(new_n10780_), .ZN(new_n10785_));
  AOI21_X1   g10703(.A1(new_n10785_), .A2(new_n10784_), .B(new_n10762_), .ZN(new_n10786_));
  NOR3_X1    g10704(.A1(new_n10786_), .A2(new_n10777_), .A3(new_n10780_), .ZN(new_n10787_));
  NOR4_X1    g10705(.A1(new_n10691_), .A2(new_n10696_), .A3(new_n10725_), .A4(new_n10774_), .ZN(new_n10788_));
  INV_X1     g10706(.I(new_n10788_), .ZN(new_n10789_));
  NOR2_X1    g10707(.A1(new_n10689_), .A2(new_n10660_), .ZN(new_n10790_));
  AOI21_X1   g10708(.A1(new_n10030_), .A2(new_n10038_), .B(new_n10685_), .ZN(new_n10791_));
  NOR2_X1    g10709(.A1(new_n10791_), .A2(new_n10790_), .ZN(new_n10792_));
  INV_X1     g10710(.I(new_n10693_), .ZN(new_n10793_));
  NAND2_X1   g10711(.A1(new_n10793_), .A2(new_n10694_), .ZN(new_n10794_));
  NOR2_X1    g10712(.A1(new_n10777_), .A2(new_n10755_), .ZN(new_n10795_));
  NOR2_X1    g10713(.A1(new_n10786_), .A2(new_n10795_), .ZN(new_n10796_));
  NAND3_X1   g10714(.A1(new_n10796_), .A2(new_n10725_), .A3(new_n10745_), .ZN(new_n10797_));
  NOR3_X1    g10715(.A1(new_n10696_), .A2(new_n10725_), .A3(new_n10774_), .ZN(new_n10798_));
  NOR4_X1    g10716(.A1(new_n10798_), .A2(new_n10792_), .A3(new_n10794_), .A4(new_n10797_), .ZN(new_n10799_));
  NOR4_X1    g10717(.A1(new_n10652_), .A2(new_n10658_), .A3(new_n10672_), .A4(new_n10789_), .ZN(new_n10800_));
  NOR2_X1    g10718(.A1(new_n10662_), .A2(new_n9360_), .ZN(new_n10801_));
  INV_X1     g10719(.I(new_n10081_), .ZN(new_n10802_));
  AOI21_X1   g10720(.A1(new_n10662_), .A2(new_n9360_), .B(new_n10802_), .ZN(new_n10803_));
  OAI22_X1   g10721(.A1(new_n10803_), .A2(new_n10801_), .B1(new_n10654_), .B2(new_n10655_), .ZN(new_n10804_));
  OAI21_X1   g10722(.A1(new_n10653_), .A2(new_n10657_), .B(new_n10804_), .ZN(new_n10805_));
  NOR2_X1    g10723(.A1(new_n10797_), .A2(new_n10794_), .ZN(new_n10806_));
  OAI21_X1   g10724(.A1(new_n10723_), .A2(new_n10722_), .B(new_n10032_), .ZN(new_n10807_));
  NAND3_X1   g10725(.A1(new_n10700_), .A2(new_n10720_), .A3(new_n10697_), .ZN(new_n10808_));
  NAND2_X1   g10726(.A1(new_n10807_), .A2(new_n10808_), .ZN(new_n10809_));
  NAND3_X1   g10727(.A1(new_n10794_), .A2(new_n10809_), .A3(new_n10773_), .ZN(new_n10810_));
  NAND3_X1   g10728(.A1(new_n10806_), .A2(new_n10691_), .A3(new_n10810_), .ZN(new_n10811_));
  AOI21_X1   g10729(.A1(new_n10811_), .A2(new_n10672_), .B(new_n10788_), .ZN(new_n10812_));
  NAND2_X1   g10730(.A1(new_n10812_), .A2(new_n10672_), .ZN(new_n10813_));
  NOR2_X1    g10731(.A1(new_n10813_), .A2(new_n10805_), .ZN(new_n10814_));
  OAI22_X1   g10732(.A1(new_n10670_), .A2(new_n10669_), .B1(new_n10076_), .B2(new_n10065_), .ZN(new_n10815_));
  NAND3_X1   g10733(.A1(new_n10666_), .A2(new_n10659_), .A3(new_n10667_), .ZN(new_n10816_));
  NAND2_X1   g10734(.A1(new_n10815_), .A2(new_n10816_), .ZN(new_n10817_));
  OAI21_X1   g10735(.A1(new_n10799_), .A2(new_n10817_), .B(new_n10789_), .ZN(new_n10818_));
  NOR2_X1    g10736(.A1(new_n10658_), .A2(new_n10672_), .ZN(new_n10819_));
  NAND2_X1   g10737(.A1(new_n10819_), .A2(new_n10818_), .ZN(new_n10820_));
  NAND3_X1   g10738(.A1(new_n10814_), .A2(new_n10652_), .A3(new_n10820_), .ZN(new_n10821_));
  AOI21_X1   g10739(.A1(new_n10646_), .A2(new_n10821_), .B(new_n10800_), .ZN(new_n10822_));
  NAND2_X1   g10740(.A1(new_n10822_), .A2(new_n10646_), .ZN(new_n10823_));
  NOR2_X1    g10741(.A1(new_n10823_), .A2(new_n10638_), .ZN(new_n10824_));
  NOR2_X1    g10742(.A1(new_n10824_), .A2(new_n10633_), .ZN(new_n10825_));
  OAI21_X1   g10743(.A1(new_n10644_), .A2(new_n10641_), .B(new_n10153_), .ZN(new_n10826_));
  NAND3_X1   g10744(.A1(new_n10642_), .A2(new_n10154_), .A3(new_n10640_), .ZN(new_n10827_));
  NAND2_X1   g10745(.A1(new_n10826_), .A2(new_n10827_), .ZN(new_n10828_));
  NAND2_X1   g10746(.A1(new_n10638_), .A2(new_n10828_), .ZN(new_n10829_));
  NOR2_X1    g10747(.A1(new_n10829_), .A2(new_n10822_), .ZN(new_n10830_));
  OAI21_X1   g10748(.A1(new_n10825_), .A2(new_n10830_), .B(new_n10633_), .ZN(new_n10831_));
  INV_X1     g10749(.I(new_n10831_), .ZN(new_n10832_));
  XOR2_X1    g10750(.A1(new_n10632_), .A2(new_n10194_), .Z(new_n10833_));
  NOR2_X1    g10751(.A1(new_n10825_), .A2(new_n10830_), .ZN(new_n10834_));
  NAND2_X1   g10752(.A1(new_n10834_), .A2(new_n10833_), .ZN(new_n10835_));
  OAI21_X1   g10753(.A1(new_n10832_), .A2(new_n10835_), .B(new_n10631_), .ZN(new_n10836_));
  XOR2_X1    g10754(.A1(new_n10203_), .A2(new_n10230_), .Z(new_n10837_));
  AOI21_X1   g10755(.A1(new_n10201_), .A2(new_n7873_), .B(new_n10837_), .ZN(new_n10838_));
  INV_X1     g10756(.I(new_n10838_), .ZN(new_n10839_));
  NAND2_X1   g10757(.A1(new_n10201_), .A2(new_n7873_), .ZN(new_n10840_));
  XOR2_X1    g10758(.A1(new_n10203_), .A2(new_n10229_), .Z(new_n10841_));
  OR2_X2     g10759(.A1(new_n10840_), .A2(new_n10841_), .Z(new_n10842_));
  NAND2_X1   g10760(.A1(new_n10842_), .A2(new_n10839_), .ZN(new_n10843_));
  INV_X1     g10761(.I(new_n10843_), .ZN(new_n10844_));
  INV_X1     g10762(.I(new_n10824_), .ZN(new_n10845_));
  NAND2_X1   g10763(.A1(new_n10831_), .A2(new_n10630_), .ZN(new_n10847_));
  NAND2_X1   g10764(.A1(new_n10844_), .A2(new_n10847_), .ZN(new_n10848_));
  NAND2_X1   g10765(.A1(new_n10848_), .A2(new_n10836_), .ZN(new_n10849_));
  NAND2_X1   g10766(.A1(new_n10203_), .A2(new_n10229_), .ZN(new_n10850_));
  NOR2_X1    g10767(.A1(new_n10837_), .A2(new_n10225_), .ZN(new_n10851_));
  XOR2_X1    g10768(.A1(new_n10851_), .A2(new_n10850_), .Z(new_n10852_));
  NOR2_X1    g10769(.A1(new_n10840_), .A2(new_n10852_), .ZN(new_n10853_));
  NAND2_X1   g10770(.A1(new_n10840_), .A2(new_n10852_), .ZN(new_n10854_));
  INV_X1     g10771(.I(new_n10854_), .ZN(new_n10855_));
  NOR2_X1    g10772(.A1(new_n10855_), .A2(new_n10853_), .ZN(new_n10856_));
  INV_X1     g10773(.I(new_n10856_), .ZN(new_n10857_));
  NOR2_X1    g10774(.A1(new_n10857_), .A2(new_n10843_), .ZN(new_n10858_));
  INV_X1     g10775(.I(new_n10858_), .ZN(new_n10859_));
  OAI21_X1   g10776(.A1(new_n10849_), .A2(new_n10859_), .B(new_n10625_), .ZN(new_n10860_));
  NOR2_X1    g10777(.A1(new_n10844_), .A2(new_n10856_), .ZN(new_n10861_));
  NAND2_X1   g10778(.A1(new_n10849_), .A2(new_n10861_), .ZN(new_n10862_));
  AOI21_X1   g10779(.A1(new_n10860_), .A2(new_n10862_), .B(new_n10625_), .ZN(new_n10863_));
  INV_X1     g10780(.I(new_n10236_), .ZN(new_n10864_));
  AOI21_X1   g10781(.A1(new_n10256_), .A2(new_n10257_), .B(new_n10864_), .ZN(new_n10865_));
  NAND2_X1   g10782(.A1(new_n10256_), .A2(new_n10257_), .ZN(new_n10866_));
  NOR2_X1    g10783(.A1(new_n10236_), .A2(new_n10866_), .ZN(new_n10867_));
  NOR2_X1    g10784(.A1(new_n10865_), .A2(new_n10867_), .ZN(new_n10868_));
  INV_X1     g10785(.I(new_n10622_), .ZN(new_n10869_));
  NOR2_X1    g10786(.A1(new_n10869_), .A2(new_n10623_), .ZN(new_n10870_));
  NOR3_X1    g10787(.A1(new_n10849_), .A2(new_n10870_), .A3(new_n10859_), .ZN(new_n10871_));
  INV_X1     g10788(.I(new_n10871_), .ZN(new_n10872_));
  AOI21_X1   g10789(.A1(new_n10868_), .A2(new_n10872_), .B(new_n10863_), .ZN(new_n10873_));
  INV_X1     g10790(.I(new_n10873_), .ZN(new_n10874_));
  INV_X1     g10791(.I(new_n10868_), .ZN(new_n10875_));
  NAND2_X1   g10792(.A1(new_n10264_), .A2(new_n10256_), .ZN(new_n10876_));
  NAND2_X1   g10793(.A1(new_n10876_), .A2(new_n10866_), .ZN(new_n10877_));
  NOR2_X1    g10794(.A1(new_n10864_), .A2(new_n10877_), .ZN(new_n10878_));
  NAND2_X1   g10795(.A1(new_n10864_), .A2(new_n10877_), .ZN(new_n10879_));
  INV_X1     g10796(.I(new_n10879_), .ZN(new_n10880_));
  NOR2_X1    g10797(.A1(new_n10880_), .A2(new_n10878_), .ZN(new_n10881_));
  INV_X1     g10798(.I(new_n10881_), .ZN(new_n10882_));
  NOR2_X1    g10799(.A1(new_n10882_), .A2(new_n10875_), .ZN(new_n10883_));
  NAND2_X1   g10800(.A1(new_n10873_), .A2(new_n10883_), .ZN(new_n10884_));
  NOR2_X1    g10801(.A1(new_n10881_), .A2(new_n10868_), .ZN(new_n10885_));
  AOI22_X1   g10802(.A1(new_n10884_), .A2(new_n10620_), .B1(new_n10874_), .B2(new_n10885_), .ZN(new_n10886_));
  NOR2_X1    g10803(.A1(new_n10886_), .A2(new_n10620_), .ZN(new_n10887_));
  NAND2_X1   g10804(.A1(new_n10886_), .A2(new_n10620_), .ZN(new_n10888_));
  AOI21_X1   g10805(.A1(new_n10611_), .A2(new_n10888_), .B(new_n10887_), .ZN(new_n10889_));
  INV_X1     g10806(.I(new_n10889_), .ZN(new_n10890_));
  NAND2_X1   g10807(.A1(new_n10291_), .A2(new_n10298_), .ZN(new_n10891_));
  NAND2_X1   g10808(.A1(new_n10609_), .A2(new_n10891_), .ZN(new_n10892_));
  NOR2_X1    g10809(.A1(new_n10271_), .A2(new_n10892_), .ZN(new_n10893_));
  NAND2_X1   g10810(.A1(new_n10271_), .A2(new_n10892_), .ZN(new_n10894_));
  INV_X1     g10811(.I(new_n10894_), .ZN(new_n10895_));
  NOR2_X1    g10812(.A1(new_n10895_), .A2(new_n10893_), .ZN(new_n10896_));
  INV_X1     g10813(.I(new_n10896_), .ZN(new_n10897_));
  NAND4_X1   g10814(.A1(new_n10890_), .A2(new_n10606_), .A3(new_n10612_), .A4(new_n10897_), .ZN(new_n10898_));
  NOR2_X1    g10815(.A1(new_n10897_), .A2(new_n10612_), .ZN(new_n10899_));
  INV_X1     g10816(.I(new_n10899_), .ZN(new_n10900_));
  NOR2_X1    g10817(.A1(new_n10896_), .A2(new_n10611_), .ZN(new_n10901_));
  NOR3_X1    g10818(.A1(new_n10890_), .A2(new_n10606_), .A3(new_n10900_), .ZN(new_n10902_));
  OAI21_X1   g10819(.A1(new_n10600_), .A2(new_n10902_), .B(new_n10898_), .ZN(new_n10903_));
  NOR2_X1    g10820(.A1(new_n10903_), .A2(new_n10600_), .ZN(new_n10904_));
  AOI21_X1   g10821(.A1(new_n10904_), .A2(new_n10595_), .B(new_n10589_), .ZN(new_n10905_));
  NOR3_X1    g10822(.A1(new_n10898_), .A2(new_n10595_), .A3(new_n10599_), .ZN(new_n10906_));
  OAI21_X1   g10823(.A1(new_n10905_), .A2(new_n10906_), .B(new_n10589_), .ZN(new_n10907_));
  XOR2_X1    g10824(.A1(new_n10477_), .A2(new_n10451_), .Z(new_n10908_));
  NOR2_X1    g10825(.A1(new_n10450_), .A2(new_n10908_), .ZN(new_n10909_));
  INV_X1     g10826(.I(new_n10450_), .ZN(new_n10910_));
  XNOR2_X1   g10827(.A1(new_n10477_), .A2(new_n10451_), .ZN(new_n10911_));
  NOR2_X1    g10828(.A1(new_n10910_), .A2(new_n10911_), .ZN(new_n10912_));
  NOR2_X1    g10829(.A1(new_n10912_), .A2(new_n10909_), .ZN(new_n10913_));
  INV_X1     g10830(.I(new_n10913_), .ZN(new_n10914_));
  NOR3_X1    g10831(.A1(new_n10905_), .A2(new_n10589_), .A3(new_n10906_), .ZN(new_n10915_));
  OAI21_X1   g10832(.A1(new_n10914_), .A2(new_n10915_), .B(new_n10907_), .ZN(new_n10916_));
  OAI21_X1   g10833(.A1(new_n10476_), .A2(new_n10474_), .B(new_n10451_), .ZN(new_n10917_));
  NOR2_X1    g10834(.A1(new_n10908_), .A2(new_n10469_), .ZN(new_n10918_));
  XOR2_X1    g10835(.A1(new_n10918_), .A2(new_n10917_), .Z(new_n10919_));
  NOR2_X1    g10836(.A1(new_n10910_), .A2(new_n10919_), .ZN(new_n10920_));
  NAND2_X1   g10837(.A1(new_n10910_), .A2(new_n10919_), .ZN(new_n10921_));
  INV_X1     g10838(.I(new_n10921_), .ZN(new_n10922_));
  NOR2_X1    g10839(.A1(new_n10922_), .A2(new_n10920_), .ZN(new_n10923_));
  INV_X1     g10840(.I(new_n10923_), .ZN(new_n10924_));
  NOR2_X1    g10841(.A1(new_n10924_), .A2(new_n10914_), .ZN(new_n10925_));
  INV_X1     g10842(.I(new_n10925_), .ZN(new_n10926_));
  OAI21_X1   g10843(.A1(new_n10916_), .A2(new_n10926_), .B(new_n10584_), .ZN(new_n10927_));
  NOR2_X1    g10844(.A1(new_n10923_), .A2(new_n10913_), .ZN(new_n10928_));
  NAND2_X1   g10845(.A1(new_n10916_), .A2(new_n10928_), .ZN(new_n10929_));
  AOI21_X1   g10846(.A1(new_n10927_), .A2(new_n10929_), .B(new_n10584_), .ZN(new_n10930_));
  NOR2_X1    g10847(.A1(new_n10484_), .A2(new_n5015_), .ZN(new_n10931_));
  XOR2_X1    g10848(.A1(new_n10490_), .A2(new_n10486_), .Z(new_n10932_));
  NOR2_X1    g10849(.A1(new_n10931_), .A2(new_n10932_), .ZN(new_n10933_));
  INV_X1     g10850(.I(new_n10933_), .ZN(new_n10934_));
  XOR2_X1    g10851(.A1(new_n10490_), .A2(new_n10486_), .Z(new_n10935_));
  NAND2_X1   g10852(.A1(new_n10931_), .A2(new_n10935_), .ZN(new_n10936_));
  NAND2_X1   g10853(.A1(new_n10934_), .A2(new_n10936_), .ZN(new_n10937_));
  INV_X1     g10854(.I(new_n10937_), .ZN(new_n10938_));
  INV_X1     g10855(.I(new_n10916_), .ZN(new_n10939_));
  NAND3_X1   g10856(.A1(new_n10939_), .A2(new_n10584_), .A3(new_n10925_), .ZN(new_n10940_));
  AOI21_X1   g10857(.A1(new_n10938_), .A2(new_n10940_), .B(new_n10930_), .ZN(new_n10941_));
  INV_X1     g10858(.I(new_n10486_), .ZN(new_n10942_));
  NAND2_X1   g10859(.A1(new_n10490_), .A2(new_n10942_), .ZN(new_n10943_));
  NOR2_X1    g10860(.A1(new_n10487_), .A2(new_n10932_), .ZN(new_n10944_));
  XNOR2_X1   g10861(.A1(new_n10944_), .A2(new_n10943_), .ZN(new_n10945_));
  NAND2_X1   g10862(.A1(new_n10931_), .A2(new_n10945_), .ZN(new_n10946_));
  NOR2_X1    g10863(.A1(new_n10931_), .A2(new_n10945_), .ZN(new_n10947_));
  INV_X1     g10864(.I(new_n10947_), .ZN(new_n10948_));
  NAND2_X1   g10865(.A1(new_n10948_), .A2(new_n10946_), .ZN(new_n10949_));
  NOR2_X1    g10866(.A1(new_n10949_), .A2(new_n10937_), .ZN(new_n10950_));
  AOI21_X1   g10867(.A1(new_n10941_), .A2(new_n10950_), .B(new_n10577_), .ZN(new_n10951_));
  INV_X1     g10868(.I(new_n10949_), .ZN(new_n10952_));
  NOR2_X1    g10869(.A1(new_n10938_), .A2(new_n10952_), .ZN(new_n10953_));
  INV_X1     g10870(.I(new_n10953_), .ZN(new_n10954_));
  NOR2_X1    g10871(.A1(new_n10941_), .A2(new_n10954_), .ZN(new_n10955_));
  NOR2_X1    g10872(.A1(new_n10951_), .A2(new_n10955_), .ZN(new_n10956_));
  INV_X1     g10873(.I(new_n10956_), .ZN(new_n10957_));
  INV_X1     g10874(.I(new_n10577_), .ZN(new_n10958_));
  AOI21_X1   g10875(.A1(new_n10525_), .A2(new_n10526_), .B(new_n10516_), .ZN(new_n10959_));
  AND3_X2    g10876(.A1(new_n10516_), .A2(new_n10525_), .A3(new_n10526_), .Z(new_n10960_));
  NOR2_X1    g10877(.A1(new_n10960_), .A2(new_n10959_), .ZN(new_n10961_));
  INV_X1     g10878(.I(new_n10961_), .ZN(new_n10962_));
  NOR2_X1    g10879(.A1(new_n10958_), .A2(new_n10962_), .ZN(new_n10963_));
  NAND2_X1   g10880(.A1(new_n10956_), .A2(new_n10963_), .ZN(new_n10964_));
  NOR2_X1    g10881(.A1(new_n10577_), .A2(new_n10961_), .ZN(new_n10965_));
  AOI22_X1   g10882(.A1(new_n10964_), .A2(new_n10571_), .B1(new_n10957_), .B2(new_n10965_), .ZN(new_n10966_));
  NAND2_X1   g10883(.A1(new_n10966_), .A2(new_n10570_), .ZN(new_n10967_));
  NOR2_X1    g10884(.A1(new_n10966_), .A2(new_n10570_), .ZN(new_n10968_));
  INV_X1     g10885(.I(new_n10968_), .ZN(new_n10969_));
  AOI21_X1   g10886(.A1(new_n10969_), .A2(new_n10967_), .B(new_n10564_), .ZN(new_n10970_));
  INV_X1     g10887(.I(new_n10564_), .ZN(new_n10971_));
  NOR4_X1    g10888(.A1(new_n10956_), .A2(new_n10571_), .A3(new_n10577_), .A4(new_n10961_), .ZN(new_n10972_));
  INV_X1     g10889(.I(new_n10972_), .ZN(new_n10973_));
  NAND3_X1   g10890(.A1(new_n10956_), .A2(new_n10571_), .A3(new_n10963_), .ZN(new_n10974_));
  AOI21_X1   g10891(.A1(new_n10973_), .A2(new_n10974_), .B(new_n10971_), .ZN(new_n10975_));
  NOR2_X1    g10892(.A1(new_n10970_), .A2(new_n10975_), .ZN(new_n10976_));
  OAI22_X1   g10893(.A1(new_n10570_), .A2(new_n9405_), .B1(new_n9408_), .B2(new_n10961_), .ZN(new_n10977_));
  OAI21_X1   g10894(.A1(new_n10564_), .A2(new_n3456_), .B(new_n10977_), .ZN(new_n10978_));
  AOI21_X1   g10895(.A1(new_n10978_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n10979_));
  XOR2_X1    g10896(.A1(new_n10976_), .A2(new_n10979_), .Z(new_n10980_));
  INV_X1     g10897(.I(new_n10980_), .ZN(new_n10981_));
  XNOR2_X1   g10898(.A1(new_n10896_), .A2(new_n10611_), .ZN(new_n10982_));
  OAI21_X1   g10899(.A1(new_n10899_), .A2(new_n10901_), .B(new_n10889_), .ZN(new_n10983_));
  OAI21_X1   g10900(.A1(new_n10889_), .A2(new_n10982_), .B(new_n10983_), .ZN(new_n10984_));
  NOR2_X1    g10901(.A1(new_n10619_), .A2(new_n10611_), .ZN(new_n10985_));
  INV_X1     g10902(.I(new_n10985_), .ZN(new_n10986_));
  AOI22_X1   g10903(.A1(new_n10986_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n10897_), .ZN(new_n10987_));
  OAI21_X1   g10904(.A1(new_n10987_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n10988_));
  XOR2_X1    g10905(.A1(new_n10984_), .A2(new_n10988_), .Z(new_n10989_));
  NOR2_X1    g10906(.A1(new_n10780_), .A2(new_n1120_), .ZN(new_n10990_));
  OAI21_X1   g10907(.A1(new_n10775_), .A2(new_n10776_), .B(new_n10755_), .ZN(new_n10991_));
  NAND3_X1   g10908(.A1(new_n10744_), .A2(new_n10740_), .A3(new_n10780_), .ZN(new_n10992_));
  OAI21_X1   g10909(.A1(new_n9984_), .A2(new_n9977_), .B(new_n10757_), .ZN(new_n10993_));
  NAND3_X1   g10910(.A1(new_n10718_), .A2(new_n10717_), .A3(new_n10733_), .ZN(new_n10994_));
  NAND4_X1   g10911(.A1(new_n10744_), .A2(new_n10993_), .A3(new_n10740_), .A4(new_n10994_), .ZN(new_n10995_));
  NAND4_X1   g10912(.A1(new_n10995_), .A2(new_n10991_), .A3(new_n10992_), .A4(new_n10772_), .ZN(new_n10996_));
  AOI21_X1   g10913(.A1(new_n10744_), .A2(new_n10740_), .B(new_n10780_), .ZN(new_n10997_));
  NOR3_X1    g10914(.A1(new_n10775_), .A2(new_n10776_), .A3(new_n10755_), .ZN(new_n10998_));
  NOR4_X1    g10915(.A1(new_n10775_), .A2(new_n10761_), .A3(new_n10776_), .A4(new_n10759_), .ZN(new_n10999_));
  OAI22_X1   g10916(.A1(new_n10999_), .A2(new_n10783_), .B1(new_n10998_), .B2(new_n10997_), .ZN(new_n11000_));
  NAND2_X1   g10917(.A1(new_n11000_), .A2(new_n10996_), .ZN(new_n11001_));
  NAND2_X1   g10918(.A1(new_n10993_), .A2(new_n10994_), .ZN(new_n11002_));
  NAND2_X1   g10919(.A1(new_n11002_), .A2(new_n10783_), .ZN(new_n11003_));
  AOI22_X1   g10920(.A1(new_n11003_), .A2(new_n5783_), .B1(new_n247_), .B2(new_n10745_), .ZN(new_n11004_));
  OAI21_X1   g10921(.A1(new_n11004_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n11005_));
  XOR2_X1    g10922(.A1(new_n11005_), .A2(new_n11001_), .Z(new_n11006_));
  NOR2_X1    g10923(.A1(new_n11006_), .A2(new_n10990_), .ZN(new_n11007_));
  NAND3_X1   g10924(.A1(new_n10783_), .A2(new_n1239_), .A3(new_n10780_), .ZN(new_n11008_));
  NAND2_X1   g10925(.A1(new_n10783_), .A2(new_n10780_), .ZN(new_n11009_));
  AOI21_X1   g10926(.A1(new_n11009_), .A2(new_n247_), .B(new_n11002_), .ZN(new_n11010_));
  OAI22_X1   g10927(.A1(new_n10772_), .A2(new_n4902_), .B1(new_n1973_), .B2(new_n10755_), .ZN(new_n11011_));
  OAI21_X1   g10928(.A1(new_n1239_), .A2(new_n10762_), .B(new_n11011_), .ZN(new_n11012_));
  AOI21_X1   g10929(.A1(new_n11008_), .A2(new_n11010_), .B(new_n11012_), .ZN(new_n11013_));
  XOR2_X1    g10930(.A1(new_n11013_), .A2(\a[23] ), .Z(new_n11014_));
  NAND2_X1   g10931(.A1(new_n10772_), .A2(new_n10780_), .ZN(new_n11015_));
  NAND2_X1   g10932(.A1(new_n10783_), .A2(new_n10755_), .ZN(new_n11016_));
  NAND2_X1   g10933(.A1(new_n11015_), .A2(new_n11016_), .ZN(new_n11017_));
  NOR2_X1    g10934(.A1(new_n10772_), .A2(new_n1973_), .ZN(new_n11018_));
  OAI21_X1   g10935(.A1(new_n10755_), .A2(new_n1239_), .B(new_n68_), .ZN(new_n11019_));
  OAI21_X1   g10936(.A1(new_n11018_), .A2(new_n11019_), .B(new_n247_), .ZN(new_n11020_));
  XOR2_X1    g10937(.A1(new_n11020_), .A2(new_n11017_), .Z(new_n11021_));
  NOR2_X1    g10938(.A1(new_n10780_), .A2(new_n1121_), .ZN(new_n11022_));
  NOR2_X1    g10939(.A1(new_n11022_), .A2(new_n68_), .ZN(new_n11023_));
  AND2_X2    g10940(.A1(new_n11021_), .A2(new_n11023_), .Z(new_n11024_));
  NAND2_X1   g10941(.A1(new_n11014_), .A2(new_n11024_), .ZN(new_n11025_));
  NAND2_X1   g10942(.A1(new_n11006_), .A2(new_n10990_), .ZN(new_n11026_));
  AOI21_X1   g10943(.A1(new_n11025_), .A2(new_n11026_), .B(new_n11007_), .ZN(new_n11027_));
  NOR2_X1    g10944(.A1(new_n10783_), .A2(new_n10755_), .ZN(new_n11028_));
  NOR2_X1    g10945(.A1(new_n10772_), .A2(new_n10780_), .ZN(new_n11029_));
  NOR2_X1    g10946(.A1(new_n11029_), .A2(new_n11028_), .ZN(new_n11030_));
  NAND2_X1   g10947(.A1(new_n10783_), .A2(new_n4613_), .ZN(new_n11031_));
  AOI21_X1   g10948(.A1(new_n10780_), .A2(new_n117_), .B(\a[26] ), .ZN(new_n11032_));
  AOI21_X1   g10949(.A1(new_n11031_), .A2(new_n11032_), .B(new_n1128_), .ZN(new_n11033_));
  XOR2_X1    g10950(.A1(new_n11030_), .A2(new_n11033_), .Z(new_n11034_));
  NOR2_X1    g10951(.A1(new_n10990_), .A2(new_n65_), .ZN(new_n11035_));
  INV_X1     g10952(.I(new_n11035_), .ZN(new_n11036_));
  XOR2_X1    g10953(.A1(new_n11034_), .A2(new_n11036_), .Z(new_n11037_));
  INV_X1     g10954(.I(new_n11037_), .ZN(new_n11038_));
  OAI21_X1   g10955(.A1(new_n10787_), .A2(new_n10773_), .B(new_n10809_), .ZN(new_n11039_));
  AOI21_X1   g10956(.A1(new_n11002_), .A2(new_n10780_), .B(new_n10745_), .ZN(new_n11040_));
  NOR3_X1    g10957(.A1(new_n10777_), .A2(new_n10772_), .A3(new_n10780_), .ZN(new_n11041_));
  AOI21_X1   g10958(.A1(new_n10745_), .A2(new_n10783_), .B(new_n10755_), .ZN(new_n11042_));
  OAI21_X1   g10959(.A1(new_n11041_), .A2(new_n11042_), .B(new_n11002_), .ZN(new_n11043_));
  AOI21_X1   g10960(.A1(new_n11043_), .A2(new_n10755_), .B(new_n10777_), .ZN(new_n11044_));
  OAI21_X1   g10961(.A1(new_n11044_), .A2(new_n11040_), .B(new_n10725_), .ZN(new_n11045_));
  NAND2_X1   g10962(.A1(new_n11045_), .A2(new_n11039_), .ZN(new_n11046_));
  NOR2_X1    g10963(.A1(new_n10762_), .A2(new_n10777_), .ZN(new_n11047_));
  OAI22_X1   g10964(.A1(new_n10725_), .A2(new_n1239_), .B1(new_n4981_), .B2(new_n11047_), .ZN(new_n11048_));
  AOI21_X1   g10965(.A1(new_n11048_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n11049_));
  XNOR2_X1   g10966(.A1(new_n11046_), .A2(new_n11049_), .ZN(new_n11050_));
  NAND2_X1   g10967(.A1(new_n11050_), .A2(new_n11038_), .ZN(new_n11051_));
  INV_X1     g10968(.I(new_n11051_), .ZN(new_n11052_));
  XOR2_X1    g10969(.A1(new_n11046_), .A2(new_n11049_), .Z(new_n11053_));
  NAND2_X1   g10970(.A1(new_n11053_), .A2(new_n11037_), .ZN(new_n11054_));
  OAI21_X1   g10971(.A1(new_n11052_), .A2(new_n11027_), .B(new_n11054_), .ZN(new_n11055_));
  AOI21_X1   g10972(.A1(new_n10796_), .A2(new_n10745_), .B(new_n10809_), .ZN(new_n11056_));
  NOR2_X1    g10973(.A1(new_n10725_), .A2(new_n10773_), .ZN(new_n11057_));
  OAI21_X1   g10974(.A1(new_n11056_), .A2(new_n11057_), .B(new_n10794_), .ZN(new_n11058_));
  INV_X1     g10975(.I(new_n10795_), .ZN(new_n11059_));
  NAND2_X1   g10976(.A1(new_n11043_), .A2(new_n11059_), .ZN(new_n11060_));
  NOR3_X1    g10977(.A1(new_n11060_), .A2(new_n10809_), .A3(new_n10777_), .ZN(new_n11061_));
  NOR2_X1    g10978(.A1(new_n10725_), .A2(new_n10774_), .ZN(new_n11062_));
  OAI21_X1   g10979(.A1(new_n11061_), .A2(new_n11062_), .B(new_n10696_), .ZN(new_n11063_));
  NAND2_X1   g10980(.A1(new_n11063_), .A2(new_n11058_), .ZN(new_n11064_));
  NAND2_X1   g10981(.A1(new_n10809_), .A2(new_n10745_), .ZN(new_n11065_));
  AOI22_X1   g10982(.A1(new_n10794_), .A2(new_n247_), .B1(new_n5783_), .B2(new_n11065_), .ZN(new_n11066_));
  OAI21_X1   g10983(.A1(new_n11066_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n11067_));
  XOR2_X1    g10984(.A1(new_n11064_), .A2(new_n11067_), .Z(new_n11068_));
  NAND3_X1   g10985(.A1(new_n10783_), .A2(new_n1128_), .A3(new_n10780_), .ZN(new_n11069_));
  AOI21_X1   g10986(.A1(new_n11009_), .A2(new_n117_), .B(new_n11002_), .ZN(new_n11070_));
  OAI22_X1   g10987(.A1(new_n10772_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10755_), .ZN(new_n11071_));
  OAI21_X1   g10988(.A1(new_n1128_), .A2(new_n10762_), .B(new_n11071_), .ZN(new_n11072_));
  AOI21_X1   g10989(.A1(new_n11069_), .A2(new_n11070_), .B(new_n11072_), .ZN(new_n11073_));
  XOR2_X1    g10990(.A1(new_n11073_), .A2(\a[26] ), .Z(new_n11074_));
  NAND2_X1   g10991(.A1(new_n11034_), .A2(new_n11035_), .ZN(new_n11075_));
  XOR2_X1    g10992(.A1(new_n11074_), .A2(new_n11075_), .Z(new_n11076_));
  XNOR2_X1   g10993(.A1(new_n11068_), .A2(new_n11076_), .ZN(new_n11077_));
  NAND2_X1   g10994(.A1(new_n11077_), .A2(new_n11055_), .ZN(new_n11078_));
  INV_X1     g10995(.I(new_n11076_), .ZN(new_n11079_));
  NOR2_X1    g10996(.A1(new_n11079_), .A2(new_n11068_), .ZN(new_n11080_));
  NAND2_X1   g10997(.A1(new_n11079_), .A2(new_n11068_), .ZN(new_n11081_));
  INV_X1     g10998(.I(new_n11081_), .ZN(new_n11082_));
  NOR2_X1    g10999(.A1(new_n11082_), .A2(new_n11080_), .ZN(new_n11083_));
  OAI21_X1   g11000(.A1(new_n11055_), .A2(new_n11083_), .B(new_n11078_), .ZN(new_n11084_));
  AOI22_X1   g11001(.A1(new_n11003_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n10745_), .ZN(new_n11085_));
  OAI21_X1   g11002(.A1(new_n11085_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n11086_));
  XOR2_X1    g11003(.A1(new_n11086_), .A2(new_n11001_), .Z(new_n11087_));
  NOR2_X1    g11004(.A1(new_n11087_), .A2(new_n11022_), .ZN(new_n11088_));
  NAND3_X1   g11005(.A1(new_n10783_), .A2(new_n5398_), .A3(new_n10780_), .ZN(new_n11089_));
  AOI21_X1   g11006(.A1(new_n11009_), .A2(new_n4717_), .B(new_n11002_), .ZN(new_n11090_));
  OAI22_X1   g11007(.A1(new_n10772_), .A2(new_n5335_), .B1(new_n4719_), .B2(new_n10755_), .ZN(new_n11091_));
  OAI21_X1   g11008(.A1(new_n5398_), .A2(new_n10762_), .B(new_n11091_), .ZN(new_n11092_));
  AOI21_X1   g11009(.A1(new_n11089_), .A2(new_n11090_), .B(new_n11092_), .ZN(new_n11093_));
  XOR2_X1    g11010(.A1(new_n11093_), .A2(\a[20] ), .Z(new_n11094_));
  NOR2_X1    g11011(.A1(new_n10772_), .A2(new_n4719_), .ZN(new_n11095_));
  OAI21_X1   g11012(.A1(new_n10755_), .A2(new_n5398_), .B(new_n90_), .ZN(new_n11096_));
  OAI21_X1   g11013(.A1(new_n11095_), .A2(new_n11096_), .B(new_n4717_), .ZN(new_n11097_));
  XOR2_X1    g11014(.A1(new_n11097_), .A2(new_n11017_), .Z(new_n11098_));
  NOR2_X1    g11015(.A1(new_n10780_), .A2(new_n1467_), .ZN(new_n11099_));
  NOR2_X1    g11016(.A1(new_n11099_), .A2(new_n90_), .ZN(new_n11100_));
  AND2_X2    g11017(.A1(new_n11098_), .A2(new_n11100_), .Z(new_n11101_));
  NAND2_X1   g11018(.A1(new_n11094_), .A2(new_n11101_), .ZN(new_n11102_));
  NAND2_X1   g11019(.A1(new_n11087_), .A2(new_n11022_), .ZN(new_n11103_));
  AOI21_X1   g11020(.A1(new_n11102_), .A2(new_n11103_), .B(new_n11088_), .ZN(new_n11104_));
  XNOR2_X1   g11021(.A1(new_n11021_), .A2(new_n11023_), .ZN(new_n11105_));
  OAI22_X1   g11022(.A1(new_n10725_), .A2(new_n5398_), .B1(new_n5336_), .B2(new_n11047_), .ZN(new_n11106_));
  AOI21_X1   g11023(.A1(new_n11106_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n11107_));
  XOR2_X1    g11024(.A1(new_n11046_), .A2(new_n11107_), .Z(new_n11108_));
  NOR2_X1    g11025(.A1(new_n11108_), .A2(new_n11105_), .ZN(new_n11109_));
  NAND2_X1   g11026(.A1(new_n11108_), .A2(new_n11105_), .ZN(new_n11110_));
  OAI21_X1   g11027(.A1(new_n11104_), .A2(new_n11109_), .B(new_n11110_), .ZN(new_n11111_));
  XNOR2_X1   g11028(.A1(new_n11014_), .A2(new_n11024_), .ZN(new_n11112_));
  AOI22_X1   g11029(.A1(new_n10794_), .A2(new_n4717_), .B1(new_n5337_), .B2(new_n11065_), .ZN(new_n11113_));
  OAI21_X1   g11030(.A1(new_n11113_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n11114_));
  XNOR2_X1   g11031(.A1(new_n11064_), .A2(new_n11114_), .ZN(new_n11115_));
  NOR2_X1    g11032(.A1(new_n11115_), .A2(new_n11112_), .ZN(new_n11116_));
  INV_X1     g11033(.I(new_n11116_), .ZN(new_n11117_));
  NAND2_X1   g11034(.A1(new_n11115_), .A2(new_n11112_), .ZN(new_n11118_));
  INV_X1     g11035(.I(new_n11118_), .ZN(new_n11119_));
  AOI21_X1   g11036(.A1(new_n11111_), .A2(new_n11117_), .B(new_n11119_), .ZN(new_n11120_));
  XNOR2_X1   g11037(.A1(new_n11006_), .A2(new_n10990_), .ZN(new_n11121_));
  INV_X1     g11038(.I(new_n11007_), .ZN(new_n11122_));
  AOI22_X1   g11039(.A1(new_n11122_), .A2(new_n11026_), .B1(new_n11014_), .B2(new_n11024_), .ZN(new_n11123_));
  INV_X1     g11040(.I(new_n11123_), .ZN(new_n11124_));
  OAI21_X1   g11041(.A1(new_n11121_), .A2(new_n11025_), .B(new_n11124_), .ZN(new_n11125_));
  OAI21_X1   g11042(.A1(new_n11060_), .A2(new_n10777_), .B(new_n10725_), .ZN(new_n11126_));
  INV_X1     g11043(.I(new_n11057_), .ZN(new_n11127_));
  NAND2_X1   g11044(.A1(new_n11126_), .A2(new_n11127_), .ZN(new_n11128_));
  NOR2_X1    g11045(.A1(new_n10787_), .A2(new_n10809_), .ZN(new_n11129_));
  NOR3_X1    g11046(.A1(new_n11129_), .A2(new_n10792_), .A3(new_n10773_), .ZN(new_n11130_));
  NAND3_X1   g11047(.A1(new_n11043_), .A2(new_n10745_), .A3(new_n10755_), .ZN(new_n11131_));
  NAND2_X1   g11048(.A1(new_n11131_), .A2(new_n10725_), .ZN(new_n11132_));
  AOI21_X1   g11049(.A1(new_n11132_), .A2(new_n10774_), .B(new_n10691_), .ZN(new_n11133_));
  OAI21_X1   g11050(.A1(new_n11130_), .A2(new_n11133_), .B(new_n11128_), .ZN(new_n11134_));
  NOR2_X1    g11051(.A1(new_n11134_), .A2(new_n10794_), .ZN(new_n11135_));
  NAND3_X1   g11052(.A1(new_n11132_), .A2(new_n10691_), .A3(new_n10774_), .ZN(new_n11136_));
  OAI21_X1   g11053(.A1(new_n11129_), .A2(new_n10773_), .B(new_n10792_), .ZN(new_n11137_));
  NAND2_X1   g11054(.A1(new_n11137_), .A2(new_n11136_), .ZN(new_n11138_));
  AOI21_X1   g11055(.A1(new_n11138_), .A2(new_n11128_), .B(new_n10696_), .ZN(new_n11139_));
  NOR2_X1    g11056(.A1(new_n11135_), .A2(new_n11139_), .ZN(new_n11140_));
  NAND2_X1   g11057(.A1(new_n10794_), .A2(new_n10809_), .ZN(new_n11141_));
  AOI22_X1   g11058(.A1(new_n11141_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n10691_), .ZN(new_n11142_));
  OAI21_X1   g11059(.A1(new_n11142_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n11143_));
  XOR2_X1    g11060(.A1(new_n11140_), .A2(new_n11143_), .Z(new_n11144_));
  NOR2_X1    g11061(.A1(new_n11144_), .A2(new_n11125_), .ZN(new_n11145_));
  NOR2_X1    g11062(.A1(new_n11120_), .A2(new_n11145_), .ZN(new_n11146_));
  AND2_X2    g11063(.A1(new_n11144_), .A2(new_n11125_), .Z(new_n11147_));
  XOR2_X1    g11064(.A1(new_n11053_), .A2(new_n11037_), .Z(new_n11148_));
  INV_X1     g11065(.I(new_n11148_), .ZN(new_n11149_));
  NAND2_X1   g11066(.A1(new_n11051_), .A2(new_n11054_), .ZN(new_n11150_));
  NAND2_X1   g11067(.A1(new_n11150_), .A2(new_n11027_), .ZN(new_n11151_));
  OAI21_X1   g11068(.A1(new_n11149_), .A2(new_n11027_), .B(new_n11151_), .ZN(new_n11152_));
  OAI21_X1   g11069(.A1(new_n10799_), .A2(new_n10788_), .B(new_n10817_), .ZN(new_n11153_));
  AOI21_X1   g11070(.A1(new_n11061_), .A2(new_n10696_), .B(new_n10792_), .ZN(new_n11154_));
  NOR3_X1    g11071(.A1(new_n11154_), .A2(new_n10691_), .A3(new_n10798_), .ZN(new_n11155_));
  AOI21_X1   g11072(.A1(new_n10806_), .A2(new_n10810_), .B(new_n10792_), .ZN(new_n11156_));
  OAI21_X1   g11073(.A1(new_n11155_), .A2(new_n11156_), .B(new_n10672_), .ZN(new_n11157_));
  NAND2_X1   g11074(.A1(new_n11157_), .A2(new_n11153_), .ZN(new_n11158_));
  NOR2_X1    g11075(.A1(new_n10792_), .A2(new_n10696_), .ZN(new_n11159_));
  OAI22_X1   g11076(.A1(new_n10672_), .A2(new_n5398_), .B1(new_n5336_), .B2(new_n11159_), .ZN(new_n11160_));
  AOI21_X1   g11077(.A1(new_n11160_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n11161_));
  XNOR2_X1   g11078(.A1(new_n11158_), .A2(new_n11161_), .ZN(new_n11162_));
  NOR2_X1    g11079(.A1(new_n11152_), .A2(new_n11162_), .ZN(new_n11163_));
  NAND2_X1   g11080(.A1(new_n11152_), .A2(new_n11162_), .ZN(new_n11164_));
  INV_X1     g11081(.I(new_n11164_), .ZN(new_n11165_));
  NOR4_X1    g11082(.A1(new_n11165_), .A2(new_n11146_), .A3(new_n11147_), .A4(new_n11163_), .ZN(new_n11166_));
  NAND2_X1   g11083(.A1(new_n11166_), .A2(new_n11084_), .ZN(new_n11167_));
  NAND2_X1   g11084(.A1(new_n10818_), .A2(new_n10672_), .ZN(new_n11168_));
  NOR2_X1    g11085(.A1(new_n10672_), .A2(new_n10788_), .ZN(new_n11169_));
  INV_X1     g11086(.I(new_n11169_), .ZN(new_n11170_));
  AOI21_X1   g11087(.A1(new_n11168_), .A2(new_n11170_), .B(new_n10658_), .ZN(new_n11171_));
  NOR2_X1    g11088(.A1(new_n10672_), .A2(new_n10789_), .ZN(new_n11172_));
  INV_X1     g11089(.I(new_n11172_), .ZN(new_n11173_));
  AOI21_X1   g11090(.A1(new_n10813_), .A2(new_n11173_), .B(new_n10805_), .ZN(new_n11174_));
  NOR2_X1    g11091(.A1(new_n11174_), .A2(new_n11171_), .ZN(new_n11175_));
  NOR2_X1    g11092(.A1(new_n10672_), .A2(new_n10792_), .ZN(new_n11176_));
  OAI22_X1   g11093(.A1(new_n11176_), .A2(new_n5336_), .B1(new_n10658_), .B2(new_n5398_), .ZN(new_n11177_));
  AOI21_X1   g11094(.A1(new_n11177_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n11178_));
  XOR2_X1    g11095(.A1(new_n11175_), .A2(new_n11178_), .Z(new_n11179_));
  NOR2_X1    g11096(.A1(new_n11164_), .A2(new_n11179_), .ZN(new_n11180_));
  OAI21_X1   g11097(.A1(new_n11166_), .A2(new_n11084_), .B(new_n11180_), .ZN(new_n11181_));
  NAND2_X1   g11098(.A1(new_n11181_), .A2(new_n11167_), .ZN(new_n11182_));
  AOI21_X1   g11099(.A1(new_n11055_), .A2(new_n11081_), .B(new_n11080_), .ZN(new_n11183_));
  INV_X1     g11100(.I(new_n11183_), .ZN(new_n11184_));
  NAND3_X1   g11101(.A1(new_n11074_), .A2(new_n11034_), .A3(new_n11035_), .ZN(new_n11185_));
  NOR4_X1    g11102(.A1(new_n10999_), .A2(new_n10997_), .A3(new_n10998_), .A4(new_n10783_), .ZN(new_n11186_));
  AOI22_X1   g11103(.A1(new_n10995_), .A2(new_n10772_), .B1(new_n10991_), .B2(new_n10992_), .ZN(new_n11187_));
  NOR2_X1    g11104(.A1(new_n11186_), .A2(new_n11187_), .ZN(new_n11188_));
  OAI21_X1   g11105(.A1(new_n4781_), .A2(new_n10762_), .B(new_n11031_), .ZN(new_n11189_));
  OAI21_X1   g11106(.A1(new_n1128_), .A2(new_n10777_), .B(new_n11189_), .ZN(new_n11190_));
  AOI21_X1   g11107(.A1(new_n11190_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n11191_));
  XOR2_X1    g11108(.A1(new_n11191_), .A2(new_n11188_), .Z(new_n11192_));
  NOR2_X1    g11109(.A1(new_n10780_), .A2(new_n918_), .ZN(new_n11193_));
  XNOR2_X1   g11110(.A1(new_n11192_), .A2(new_n11193_), .ZN(new_n11194_));
  NOR2_X1    g11111(.A1(new_n11192_), .A2(new_n11193_), .ZN(new_n11195_));
  NAND2_X1   g11112(.A1(new_n11192_), .A2(new_n11193_), .ZN(new_n11196_));
  INV_X1     g11113(.I(new_n11196_), .ZN(new_n11197_));
  OAI21_X1   g11114(.A1(new_n11197_), .A2(new_n11195_), .B(new_n11185_), .ZN(new_n11198_));
  OAI21_X1   g11115(.A1(new_n11185_), .A2(new_n11194_), .B(new_n11198_), .ZN(new_n11199_));
  AOI22_X1   g11116(.A1(new_n11141_), .A2(new_n5783_), .B1(new_n247_), .B2(new_n10691_), .ZN(new_n11200_));
  OAI21_X1   g11117(.A1(new_n11200_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n11201_));
  XOR2_X1    g11118(.A1(new_n11140_), .A2(new_n11201_), .Z(new_n11202_));
  XOR2_X1    g11119(.A1(new_n11202_), .A2(new_n11199_), .Z(new_n11203_));
  NAND2_X1   g11120(.A1(new_n11203_), .A2(new_n11184_), .ZN(new_n11204_));
  NOR2_X1    g11121(.A1(new_n11202_), .A2(new_n11199_), .ZN(new_n11205_));
  AND2_X2    g11122(.A1(new_n11202_), .A2(new_n11199_), .Z(new_n11206_));
  OAI21_X1   g11123(.A1(new_n11206_), .A2(new_n11205_), .B(new_n11183_), .ZN(new_n11207_));
  NAND2_X1   g11124(.A1(new_n11204_), .A2(new_n11207_), .ZN(new_n11208_));
  INV_X1     g11125(.I(new_n11208_), .ZN(new_n11209_));
  NOR2_X1    g11126(.A1(new_n10812_), .A2(new_n10817_), .ZN(new_n11210_));
  NOR2_X1    g11127(.A1(new_n11210_), .A2(new_n11169_), .ZN(new_n11211_));
  NOR3_X1    g11128(.A1(new_n10148_), .A2(new_n10110_), .A3(new_n10113_), .ZN(new_n11212_));
  AOI21_X1   g11129(.A1(new_n10111_), .A2(new_n10114_), .B(new_n10649_), .ZN(new_n11213_));
  NOR2_X1    g11130(.A1(new_n11213_), .A2(new_n11212_), .ZN(new_n11214_));
  NOR2_X1    g11131(.A1(new_n11214_), .A2(new_n10818_), .ZN(new_n11215_));
  NOR2_X1    g11132(.A1(new_n10812_), .A2(new_n10652_), .ZN(new_n11216_));
  NOR2_X1    g11133(.A1(new_n11216_), .A2(new_n11215_), .ZN(new_n11217_));
  NOR3_X1    g11134(.A1(new_n11217_), .A2(new_n11211_), .A3(new_n10805_), .ZN(new_n11218_));
  NAND2_X1   g11135(.A1(new_n11168_), .A2(new_n11170_), .ZN(new_n11219_));
  NAND2_X1   g11136(.A1(new_n10812_), .A2(new_n10652_), .ZN(new_n11220_));
  NAND2_X1   g11137(.A1(new_n11214_), .A2(new_n10818_), .ZN(new_n11221_));
  NAND2_X1   g11138(.A1(new_n11220_), .A2(new_n11221_), .ZN(new_n11222_));
  AOI21_X1   g11139(.A1(new_n11222_), .A2(new_n11219_), .B(new_n10658_), .ZN(new_n11223_));
  NOR2_X1    g11140(.A1(new_n11218_), .A2(new_n11223_), .ZN(new_n11224_));
  OAI22_X1   g11141(.A1(new_n10819_), .A2(new_n5336_), .B1(new_n11214_), .B2(new_n5398_), .ZN(new_n11225_));
  AOI21_X1   g11142(.A1(new_n11225_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n11226_));
  XOR2_X1    g11143(.A1(new_n11224_), .A2(new_n11226_), .Z(new_n11227_));
  INV_X1     g11144(.I(new_n11227_), .ZN(new_n11228_));
  NOR2_X1    g11145(.A1(new_n11209_), .A2(new_n11228_), .ZN(new_n11229_));
  NOR2_X1    g11146(.A1(new_n11208_), .A2(new_n11227_), .ZN(new_n11230_));
  OAI21_X1   g11147(.A1(new_n11229_), .A2(new_n11230_), .B(new_n11182_), .ZN(new_n11231_));
  XOR2_X1    g11148(.A1(new_n11208_), .A2(new_n11227_), .Z(new_n11232_));
  NAND3_X1   g11149(.A1(new_n11232_), .A2(new_n11167_), .A3(new_n11181_), .ZN(new_n11233_));
  AND2_X2    g11150(.A1(new_n11233_), .A2(new_n11231_), .Z(new_n11234_));
  INV_X1     g11151(.I(new_n11234_), .ZN(new_n11235_));
  INV_X1     g11152(.I(new_n10800_), .ZN(new_n11236_));
  AOI21_X1   g11153(.A1(new_n11236_), .A2(new_n10821_), .B(new_n10646_), .ZN(new_n11237_));
  INV_X1     g11154(.I(new_n11237_), .ZN(new_n11238_));
  OAI21_X1   g11155(.A1(new_n10814_), .A2(new_n11214_), .B(new_n10820_), .ZN(new_n11239_));
  NOR2_X1    g11156(.A1(new_n11239_), .A2(new_n10652_), .ZN(new_n11240_));
  NOR2_X1    g11157(.A1(new_n10818_), .A2(new_n10817_), .ZN(new_n11241_));
  NAND2_X1   g11158(.A1(new_n11241_), .A2(new_n10658_), .ZN(new_n11242_));
  AOI22_X1   g11159(.A1(new_n11242_), .A2(new_n10652_), .B1(new_n10818_), .B2(new_n10819_), .ZN(new_n11243_));
  NOR2_X1    g11160(.A1(new_n11243_), .A2(new_n11214_), .ZN(new_n11244_));
  OAI21_X1   g11161(.A1(new_n11244_), .A2(new_n11240_), .B(new_n10646_), .ZN(new_n11245_));
  NAND2_X1   g11162(.A1(new_n11245_), .A2(new_n11238_), .ZN(new_n11246_));
  AOI21_X1   g11163(.A1(new_n10652_), .A2(new_n10805_), .B(new_n5420_), .ZN(new_n11247_));
  NOR2_X1    g11164(.A1(new_n10646_), .A2(new_n1620_), .ZN(new_n11248_));
  OAI21_X1   g11165(.A1(new_n11248_), .A2(new_n11247_), .B(new_n126_), .ZN(new_n11249_));
  NAND2_X1   g11166(.A1(new_n11249_), .A2(new_n4660_), .ZN(new_n11250_));
  XOR2_X1    g11167(.A1(new_n11246_), .A2(new_n11250_), .Z(new_n11251_));
  NOR2_X1    g11168(.A1(new_n11146_), .A2(new_n11147_), .ZN(new_n11252_));
  NOR2_X1    g11169(.A1(new_n11165_), .A2(new_n11163_), .ZN(new_n11253_));
  XNOR2_X1   g11170(.A1(new_n11253_), .A2(new_n11252_), .ZN(new_n11254_));
  INV_X1     g11171(.I(new_n11179_), .ZN(new_n11255_));
  NAND2_X1   g11172(.A1(new_n11084_), .A2(new_n11255_), .ZN(new_n11256_));
  XNOR2_X1   g11173(.A1(new_n11166_), .A2(new_n11256_), .ZN(new_n11257_));
  XOR2_X1    g11174(.A1(new_n11257_), .A2(new_n11164_), .Z(new_n11258_));
  INV_X1     g11175(.I(new_n11258_), .ZN(new_n11259_));
  NOR2_X1    g11176(.A1(new_n10822_), .A2(new_n10828_), .ZN(new_n11260_));
  NOR2_X1    g11177(.A1(new_n10646_), .A2(new_n10800_), .ZN(new_n11262_));
  OAI21_X1   g11178(.A1(new_n11260_), .A2(new_n11262_), .B(new_n10638_), .ZN(new_n11263_));
  INV_X1     g11179(.I(new_n10638_), .ZN(new_n11264_));
  NAND2_X1   g11180(.A1(new_n10828_), .A2(new_n10800_), .ZN(new_n11265_));
  NAND2_X1   g11181(.A1(new_n10823_), .A2(new_n11265_), .ZN(new_n11266_));
  NAND2_X1   g11182(.A1(new_n11266_), .A2(new_n11264_), .ZN(new_n11267_));
  NAND2_X1   g11183(.A1(new_n11267_), .A2(new_n11263_), .ZN(new_n11268_));
  NAND2_X1   g11184(.A1(new_n10828_), .A2(new_n10652_), .ZN(new_n11269_));
  AOI22_X1   g11185(.A1(new_n10638_), .A2(new_n4660_), .B1(new_n5421_), .B2(new_n11269_), .ZN(new_n11270_));
  NOR2_X1    g11186(.A1(new_n11270_), .A2(\a[17] ), .ZN(new_n11271_));
  NOR2_X1    g11187(.A1(new_n11271_), .A2(new_n1620_), .ZN(new_n11272_));
  XNOR2_X1   g11188(.A1(new_n11268_), .A2(new_n11272_), .ZN(new_n11273_));
  INV_X1     g11189(.I(new_n11273_), .ZN(new_n11274_));
  NOR2_X1    g11190(.A1(new_n11259_), .A2(new_n11274_), .ZN(new_n11275_));
  NOR2_X1    g11191(.A1(new_n11258_), .A2(new_n11273_), .ZN(new_n11276_));
  NOR2_X1    g11192(.A1(new_n11275_), .A2(new_n11276_), .ZN(new_n11277_));
  OAI21_X1   g11193(.A1(new_n11277_), .A2(new_n11254_), .B(new_n11251_), .ZN(new_n11278_));
  INV_X1     g11194(.I(new_n11120_), .ZN(new_n11279_));
  XOR2_X1    g11195(.A1(new_n11144_), .A2(new_n11125_), .Z(new_n11280_));
  NAND2_X1   g11196(.A1(new_n11280_), .A2(new_n11279_), .ZN(new_n11281_));
  OAI21_X1   g11197(.A1(new_n11147_), .A2(new_n11145_), .B(new_n11120_), .ZN(new_n11282_));
  NAND2_X1   g11198(.A1(new_n11281_), .A2(new_n11282_), .ZN(new_n11283_));
  INV_X1     g11199(.I(new_n11283_), .ZN(new_n11284_));
  AOI22_X1   g11200(.A1(new_n11003_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n10745_), .ZN(new_n11285_));
  OAI21_X1   g11201(.A1(new_n11285_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n11286_));
  XOR2_X1    g11202(.A1(new_n11286_), .A2(new_n11001_), .Z(new_n11287_));
  NOR2_X1    g11203(.A1(new_n11287_), .A2(new_n11099_), .ZN(new_n11288_));
  INV_X1     g11204(.I(new_n11288_), .ZN(new_n11289_));
  NAND3_X1   g11205(.A1(new_n10783_), .A2(new_n1620_), .A3(new_n10780_), .ZN(new_n11290_));
  AOI21_X1   g11206(.A1(new_n11009_), .A2(new_n4660_), .B(new_n11002_), .ZN(new_n11291_));
  OAI22_X1   g11207(.A1(new_n10772_), .A2(new_n5419_), .B1(new_n1622_), .B2(new_n10755_), .ZN(new_n11292_));
  OAI21_X1   g11208(.A1(new_n1620_), .A2(new_n10762_), .B(new_n11292_), .ZN(new_n11293_));
  AOI21_X1   g11209(.A1(new_n11290_), .A2(new_n11291_), .B(new_n11293_), .ZN(new_n11294_));
  XOR2_X1    g11210(.A1(new_n11294_), .A2(\a[17] ), .Z(new_n11295_));
  INV_X1     g11211(.I(new_n11295_), .ZN(new_n11296_));
  NAND2_X1   g11212(.A1(new_n10783_), .A2(new_n4661_), .ZN(new_n11297_));
  AOI21_X1   g11213(.A1(new_n10780_), .A2(new_n4660_), .B(\a[17] ), .ZN(new_n11298_));
  AOI21_X1   g11214(.A1(new_n11297_), .A2(new_n11298_), .B(new_n1620_), .ZN(new_n11299_));
  XOR2_X1    g11215(.A1(new_n11299_), .A2(new_n11017_), .Z(new_n11300_));
  NOR2_X1    g11216(.A1(new_n10780_), .A2(new_n1468_), .ZN(new_n11301_));
  NOR2_X1    g11217(.A1(new_n11301_), .A2(new_n126_), .ZN(new_n11302_));
  INV_X1     g11218(.I(new_n11302_), .ZN(new_n11303_));
  NOR2_X1    g11219(.A1(new_n11300_), .A2(new_n11303_), .ZN(new_n11304_));
  INV_X1     g11220(.I(new_n11304_), .ZN(new_n11305_));
  NOR2_X1    g11221(.A1(new_n11296_), .A2(new_n11305_), .ZN(new_n11306_));
  AND2_X2    g11222(.A1(new_n11287_), .A2(new_n11099_), .Z(new_n11307_));
  OAI21_X1   g11223(.A1(new_n11306_), .A2(new_n11307_), .B(new_n11289_), .ZN(new_n11308_));
  XNOR2_X1   g11224(.A1(new_n11098_), .A2(new_n11100_), .ZN(new_n11309_));
  OAI22_X1   g11225(.A1(new_n10725_), .A2(new_n1620_), .B1(new_n5420_), .B2(new_n11047_), .ZN(new_n11310_));
  AOI21_X1   g11226(.A1(new_n11310_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n11311_));
  XOR2_X1    g11227(.A1(new_n11046_), .A2(new_n11311_), .Z(new_n11312_));
  NOR2_X1    g11228(.A1(new_n11312_), .A2(new_n11309_), .ZN(new_n11313_));
  INV_X1     g11229(.I(new_n11313_), .ZN(new_n11314_));
  NAND2_X1   g11230(.A1(new_n11312_), .A2(new_n11309_), .ZN(new_n11315_));
  INV_X1     g11231(.I(new_n11315_), .ZN(new_n11316_));
  AOI21_X1   g11232(.A1(new_n11308_), .A2(new_n11314_), .B(new_n11316_), .ZN(new_n11317_));
  XNOR2_X1   g11233(.A1(new_n11094_), .A2(new_n11101_), .ZN(new_n11318_));
  AOI22_X1   g11234(.A1(new_n10794_), .A2(new_n4660_), .B1(new_n5421_), .B2(new_n11065_), .ZN(new_n11319_));
  OAI21_X1   g11235(.A1(new_n11319_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n11320_));
  XOR2_X1    g11236(.A1(new_n11064_), .A2(new_n11320_), .Z(new_n11321_));
  INV_X1     g11237(.I(new_n11321_), .ZN(new_n11322_));
  NOR2_X1    g11238(.A1(new_n11322_), .A2(new_n11318_), .ZN(new_n11323_));
  NAND2_X1   g11239(.A1(new_n11322_), .A2(new_n11318_), .ZN(new_n11324_));
  OAI21_X1   g11240(.A1(new_n11317_), .A2(new_n11323_), .B(new_n11324_), .ZN(new_n11325_));
  XNOR2_X1   g11241(.A1(new_n11087_), .A2(new_n11022_), .ZN(new_n11326_));
  NOR2_X1    g11242(.A1(new_n11326_), .A2(new_n11102_), .ZN(new_n11327_));
  INV_X1     g11243(.I(new_n11088_), .ZN(new_n11328_));
  NAND2_X1   g11244(.A1(new_n11328_), .A2(new_n11103_), .ZN(new_n11329_));
  AOI21_X1   g11245(.A1(new_n11102_), .A2(new_n11329_), .B(new_n11327_), .ZN(new_n11330_));
  NAND3_X1   g11246(.A1(new_n11138_), .A2(new_n10696_), .A3(new_n11128_), .ZN(new_n11331_));
  NAND2_X1   g11247(.A1(new_n11134_), .A2(new_n10794_), .ZN(new_n11332_));
  NAND2_X1   g11248(.A1(new_n11332_), .A2(new_n11331_), .ZN(new_n11333_));
  AOI22_X1   g11249(.A1(new_n11141_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n10691_), .ZN(new_n11334_));
  OAI21_X1   g11250(.A1(new_n11334_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n11335_));
  XOR2_X1    g11251(.A1(new_n11333_), .A2(new_n11335_), .Z(new_n11336_));
  NAND2_X1   g11252(.A1(new_n11336_), .A2(new_n11330_), .ZN(new_n11337_));
  NAND2_X1   g11253(.A1(new_n11325_), .A2(new_n11337_), .ZN(new_n11338_));
  OR2_X2     g11254(.A1(new_n11336_), .A2(new_n11330_), .Z(new_n11339_));
  NAND2_X1   g11255(.A1(new_n11338_), .A2(new_n11339_), .ZN(new_n11340_));
  XNOR2_X1   g11256(.A1(new_n11108_), .A2(new_n11105_), .ZN(new_n11341_));
  INV_X1     g11257(.I(new_n11109_), .ZN(new_n11342_));
  NAND2_X1   g11258(.A1(new_n11342_), .A2(new_n11110_), .ZN(new_n11343_));
  NAND2_X1   g11259(.A1(new_n11343_), .A2(new_n11104_), .ZN(new_n11344_));
  OAI21_X1   g11260(.A1(new_n11104_), .A2(new_n11341_), .B(new_n11344_), .ZN(new_n11345_));
  OAI22_X1   g11261(.A1(new_n10672_), .A2(new_n1620_), .B1(new_n5420_), .B2(new_n11159_), .ZN(new_n11346_));
  AOI21_X1   g11262(.A1(new_n11346_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n11347_));
  XNOR2_X1   g11263(.A1(new_n11158_), .A2(new_n11347_), .ZN(new_n11348_));
  NAND2_X1   g11264(.A1(new_n11345_), .A2(new_n11348_), .ZN(new_n11349_));
  NAND2_X1   g11265(.A1(new_n11340_), .A2(new_n11349_), .ZN(new_n11350_));
  OR2_X2     g11266(.A1(new_n11345_), .A2(new_n11348_), .Z(new_n11351_));
  XOR2_X1    g11267(.A1(new_n11115_), .A2(new_n11112_), .Z(new_n11352_));
  NAND2_X1   g11268(.A1(new_n11352_), .A2(new_n11111_), .ZN(new_n11353_));
  NOR2_X1    g11269(.A1(new_n11119_), .A2(new_n11116_), .ZN(new_n11354_));
  OAI21_X1   g11270(.A1(new_n11111_), .A2(new_n11354_), .B(new_n11353_), .ZN(new_n11355_));
  OAI22_X1   g11271(.A1(new_n11176_), .A2(new_n5420_), .B1(new_n10658_), .B2(new_n1620_), .ZN(new_n11356_));
  AOI21_X1   g11272(.A1(new_n11356_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n11357_));
  XOR2_X1    g11273(.A1(new_n11175_), .A2(new_n11357_), .Z(new_n11358_));
  NOR2_X1    g11274(.A1(new_n11355_), .A2(new_n11358_), .ZN(new_n11359_));
  NAND2_X1   g11275(.A1(new_n11355_), .A2(new_n11358_), .ZN(new_n11360_));
  INV_X1     g11276(.I(new_n11360_), .ZN(new_n11361_));
  NOR2_X1    g11277(.A1(new_n11361_), .A2(new_n11359_), .ZN(new_n11362_));
  NAND3_X1   g11278(.A1(new_n11362_), .A2(new_n11350_), .A3(new_n11351_), .ZN(new_n11363_));
  NOR2_X1    g11279(.A1(new_n11363_), .A2(new_n11284_), .ZN(new_n11364_));
  NAND2_X1   g11280(.A1(new_n11363_), .A2(new_n11284_), .ZN(new_n11365_));
  OAI22_X1   g11281(.A1(new_n10819_), .A2(new_n5420_), .B1(new_n11214_), .B2(new_n1620_), .ZN(new_n11366_));
  AOI21_X1   g11282(.A1(new_n11366_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n11367_));
  XOR2_X1    g11283(.A1(new_n11224_), .A2(new_n11367_), .Z(new_n11368_));
  NOR2_X1    g11284(.A1(new_n11360_), .A2(new_n11368_), .ZN(new_n11369_));
  AOI21_X1   g11285(.A1(new_n11365_), .A2(new_n11369_), .B(new_n11364_), .ZN(new_n11370_));
  AOI21_X1   g11286(.A1(new_n11277_), .A2(new_n11254_), .B(new_n11370_), .ZN(new_n11371_));
  NAND3_X1   g11287(.A1(new_n11371_), .A2(new_n11278_), .A3(new_n11235_), .ZN(new_n11372_));
  AOI21_X1   g11288(.A1(new_n11371_), .A2(new_n11278_), .B(new_n11235_), .ZN(new_n11373_));
  NOR2_X1    g11289(.A1(new_n11260_), .A2(new_n11262_), .ZN(new_n11374_));
  INV_X1     g11290(.I(new_n10822_), .ZN(new_n11375_));
  NOR2_X1    g11291(.A1(new_n10633_), .A2(new_n11375_), .ZN(new_n11376_));
  NOR2_X1    g11292(.A1(new_n10833_), .A2(new_n10822_), .ZN(new_n11377_));
  NOR2_X1    g11293(.A1(new_n11376_), .A2(new_n11377_), .ZN(new_n11378_));
  NOR3_X1    g11294(.A1(new_n11378_), .A2(new_n11374_), .A3(new_n10638_), .ZN(new_n11379_));
  INV_X1     g11295(.I(new_n11374_), .ZN(new_n11380_));
  NAND2_X1   g11296(.A1(new_n10833_), .A2(new_n10822_), .ZN(new_n11381_));
  NAND2_X1   g11297(.A1(new_n10633_), .A2(new_n11375_), .ZN(new_n11382_));
  NAND2_X1   g11298(.A1(new_n11382_), .A2(new_n11381_), .ZN(new_n11383_));
  AOI21_X1   g11299(.A1(new_n11383_), .A2(new_n11380_), .B(new_n11264_), .ZN(new_n11384_));
  NOR2_X1    g11300(.A1(new_n11379_), .A2(new_n11384_), .ZN(new_n11385_));
  INV_X1     g11301(.I(new_n10829_), .ZN(new_n11386_));
  OAI22_X1   g11302(.A1(new_n11386_), .A2(new_n5420_), .B1(new_n1620_), .B2(new_n10633_), .ZN(new_n11387_));
  AOI21_X1   g11303(.A1(new_n11387_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n11388_));
  XOR2_X1    g11304(.A1(new_n11385_), .A2(new_n11388_), .Z(new_n11389_));
  INV_X1     g11305(.I(new_n11389_), .ZN(new_n11390_));
  NAND2_X1   g11306(.A1(new_n11275_), .A2(new_n11390_), .ZN(new_n11391_));
  OAI21_X1   g11307(.A1(new_n11373_), .A2(new_n11391_), .B(new_n11372_), .ZN(new_n11392_));
  INV_X1     g11308(.I(new_n11229_), .ZN(new_n11393_));
  AOI21_X1   g11309(.A1(new_n11393_), .A2(new_n11182_), .B(new_n11230_), .ZN(new_n11394_));
  INV_X1     g11310(.I(new_n11394_), .ZN(new_n11395_));
  NOR2_X1    g11311(.A1(new_n11205_), .A2(new_n11183_), .ZN(new_n11396_));
  NOR2_X1    g11312(.A1(new_n11396_), .A2(new_n11206_), .ZN(new_n11397_));
  AOI21_X1   g11313(.A1(new_n11185_), .A2(new_n11196_), .B(new_n11195_), .ZN(new_n11398_));
  INV_X1     g11314(.I(new_n11398_), .ZN(new_n11399_));
  OAI22_X1   g11315(.A1(new_n4612_), .A2(new_n10762_), .B1(new_n10777_), .B2(new_n4781_), .ZN(new_n11400_));
  OAI21_X1   g11316(.A1(new_n10725_), .A2(new_n1128_), .B(new_n11400_), .ZN(new_n11401_));
  AOI21_X1   g11317(.A1(new_n11401_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n11402_));
  XOR2_X1    g11318(.A1(new_n11046_), .A2(new_n11402_), .Z(new_n11403_));
  NAND2_X1   g11319(.A1(new_n10783_), .A2(new_n4570_), .ZN(new_n11404_));
  AOI21_X1   g11320(.A1(new_n10780_), .A2(new_n101_), .B(\a[29] ), .ZN(new_n11405_));
  AOI21_X1   g11321(.A1(new_n11404_), .A2(new_n11405_), .B(new_n79_), .ZN(new_n11406_));
  XOR2_X1    g11322(.A1(new_n11030_), .A2(new_n11406_), .Z(new_n11407_));
  NOR2_X1    g11323(.A1(new_n11193_), .A2(new_n72_), .ZN(new_n11408_));
  INV_X1     g11324(.I(new_n11408_), .ZN(new_n11409_));
  XOR2_X1    g11325(.A1(new_n11407_), .A2(new_n11409_), .Z(new_n11410_));
  XOR2_X1    g11326(.A1(new_n11403_), .A2(new_n11410_), .Z(new_n11411_));
  NAND2_X1   g11327(.A1(new_n11411_), .A2(new_n11399_), .ZN(new_n11412_));
  AND2_X2    g11328(.A1(new_n11403_), .A2(new_n11410_), .Z(new_n11413_));
  NOR2_X1    g11329(.A1(new_n11403_), .A2(new_n11410_), .ZN(new_n11414_));
  OAI21_X1   g11330(.A1(new_n11413_), .A2(new_n11414_), .B(new_n11398_), .ZN(new_n11415_));
  NAND2_X1   g11331(.A1(new_n11412_), .A2(new_n11415_), .ZN(new_n11416_));
  OAI22_X1   g11332(.A1(new_n10672_), .A2(new_n1239_), .B1(new_n4981_), .B2(new_n11159_), .ZN(new_n11417_));
  AOI21_X1   g11333(.A1(new_n11417_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n11418_));
  XNOR2_X1   g11334(.A1(new_n11158_), .A2(new_n11418_), .ZN(new_n11419_));
  NOR2_X1    g11335(.A1(new_n11416_), .A2(new_n11419_), .ZN(new_n11420_));
  NAND2_X1   g11336(.A1(new_n11416_), .A2(new_n11419_), .ZN(new_n11421_));
  INV_X1     g11337(.I(new_n11421_), .ZN(new_n11422_));
  NOR2_X1    g11338(.A1(new_n11422_), .A2(new_n11420_), .ZN(new_n11423_));
  INV_X1     g11339(.I(new_n11423_), .ZN(new_n11424_));
  NAND2_X1   g11340(.A1(new_n11424_), .A2(new_n11397_), .ZN(new_n11425_));
  INV_X1     g11341(.I(new_n11425_), .ZN(new_n11426_));
  NOR2_X1    g11342(.A1(new_n11424_), .A2(new_n11397_), .ZN(new_n11427_));
  AOI21_X1   g11343(.A1(new_n10652_), .A2(new_n10805_), .B(new_n5336_), .ZN(new_n11428_));
  NOR2_X1    g11344(.A1(new_n10646_), .A2(new_n5398_), .ZN(new_n11429_));
  OAI21_X1   g11345(.A1(new_n11429_), .A2(new_n11428_), .B(new_n90_), .ZN(new_n11430_));
  NAND2_X1   g11346(.A1(new_n11430_), .A2(new_n4717_), .ZN(new_n11431_));
  XOR2_X1    g11347(.A1(new_n11246_), .A2(new_n11431_), .Z(new_n11432_));
  INV_X1     g11348(.I(new_n11432_), .ZN(new_n11433_));
  NOR3_X1    g11349(.A1(new_n11426_), .A2(new_n11427_), .A3(new_n11433_), .ZN(new_n11434_));
  NOR2_X1    g11350(.A1(new_n11426_), .A2(new_n11427_), .ZN(new_n11435_));
  NOR2_X1    g11351(.A1(new_n11435_), .A2(new_n11432_), .ZN(new_n11436_));
  OAI21_X1   g11352(.A1(new_n11434_), .A2(new_n11436_), .B(new_n11395_), .ZN(new_n11437_));
  XOR2_X1    g11353(.A1(new_n11435_), .A2(new_n11433_), .Z(new_n11438_));
  OR2_X2     g11354(.A1(new_n11438_), .A2(new_n11395_), .Z(new_n11439_));
  NAND2_X1   g11355(.A1(new_n11439_), .A2(new_n11437_), .ZN(new_n11440_));
  NAND2_X1   g11356(.A1(new_n10834_), .A2(new_n10633_), .ZN(new_n11441_));
  OAI21_X1   g11357(.A1(new_n10845_), .A2(new_n10830_), .B(new_n10833_), .ZN(new_n11442_));
  AOI21_X1   g11358(.A1(new_n11441_), .A2(new_n11442_), .B(new_n10631_), .ZN(new_n11443_));
  AOI21_X1   g11359(.A1(new_n10835_), .A2(new_n10831_), .B(new_n10630_), .ZN(new_n11444_));
  NOR2_X1    g11360(.A1(new_n11444_), .A2(new_n11443_), .ZN(new_n11445_));
  NAND2_X1   g11361(.A1(new_n10833_), .A2(new_n10638_), .ZN(new_n11446_));
  AOI22_X1   g11362(.A1(new_n10630_), .A2(new_n4660_), .B1(new_n5421_), .B2(new_n11446_), .ZN(new_n11447_));
  NOR2_X1    g11363(.A1(new_n11447_), .A2(\a[17] ), .ZN(new_n11448_));
  NOR2_X1    g11364(.A1(new_n11448_), .A2(new_n1620_), .ZN(new_n11449_));
  XOR2_X1    g11365(.A1(new_n11445_), .A2(new_n11449_), .Z(new_n11450_));
  INV_X1     g11366(.I(new_n11450_), .ZN(new_n11451_));
  XOR2_X1    g11367(.A1(new_n11440_), .A2(new_n11451_), .Z(new_n11452_));
  INV_X1     g11368(.I(new_n11452_), .ZN(new_n11453_));
  INV_X1     g11369(.I(new_n11440_), .ZN(new_n11454_));
  NOR2_X1    g11370(.A1(new_n11454_), .A2(new_n11451_), .ZN(new_n11455_));
  NOR2_X1    g11371(.A1(new_n11440_), .A2(new_n11450_), .ZN(new_n11456_));
  NOR2_X1    g11372(.A1(new_n11455_), .A2(new_n11456_), .ZN(new_n11457_));
  NOR2_X1    g11373(.A1(new_n11392_), .A2(new_n11457_), .ZN(new_n11458_));
  AOI21_X1   g11374(.A1(new_n11392_), .A2(new_n11453_), .B(new_n11458_), .ZN(new_n11459_));
  NOR2_X1    g11375(.A1(new_n11284_), .A2(new_n11368_), .ZN(new_n11460_));
  XNOR2_X1   g11376(.A1(new_n11363_), .A2(new_n11460_), .ZN(new_n11461_));
  XOR2_X1    g11377(.A1(new_n11461_), .A2(new_n11360_), .Z(new_n11462_));
  INV_X1     g11378(.I(new_n11462_), .ZN(new_n11463_));
  AOI21_X1   g11379(.A1(new_n10652_), .A2(new_n10805_), .B(new_n5967_), .ZN(new_n11464_));
  NOR2_X1    g11380(.A1(new_n10646_), .A2(new_n643_), .ZN(new_n11465_));
  OAI21_X1   g11381(.A1(new_n11465_), .A2(new_n11464_), .B(new_n279_), .ZN(new_n11466_));
  NAND2_X1   g11382(.A1(new_n11466_), .A2(new_n785_), .ZN(new_n11467_));
  XOR2_X1    g11383(.A1(new_n11246_), .A2(new_n11467_), .Z(new_n11468_));
  XOR2_X1    g11384(.A1(new_n11345_), .A2(new_n11348_), .Z(new_n11469_));
  NAND2_X1   g11385(.A1(new_n11469_), .A2(new_n11340_), .ZN(new_n11470_));
  AOI21_X1   g11386(.A1(new_n11351_), .A2(new_n11349_), .B(new_n11340_), .ZN(new_n11471_));
  INV_X1     g11387(.I(new_n11471_), .ZN(new_n11472_));
  NAND2_X1   g11388(.A1(new_n11472_), .A2(new_n11470_), .ZN(new_n11473_));
  INV_X1     g11389(.I(new_n11473_), .ZN(new_n11474_));
  NAND2_X1   g11390(.A1(new_n11350_), .A2(new_n11351_), .ZN(new_n11475_));
  XNOR2_X1   g11391(.A1(new_n11362_), .A2(new_n11475_), .ZN(new_n11476_));
  AOI22_X1   g11392(.A1(new_n10638_), .A2(new_n785_), .B1(new_n5968_), .B2(new_n11269_), .ZN(new_n11477_));
  OAI21_X1   g11393(.A1(new_n11477_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n11478_));
  XOR2_X1    g11394(.A1(new_n11268_), .A2(new_n11478_), .Z(new_n11479_));
  AND2_X2    g11395(.A1(new_n11476_), .A2(new_n11479_), .Z(new_n11480_));
  NOR2_X1    g11396(.A1(new_n11476_), .A2(new_n11479_), .ZN(new_n11481_));
  NOR2_X1    g11397(.A1(new_n11480_), .A2(new_n11481_), .ZN(new_n11482_));
  OAI21_X1   g11398(.A1(new_n11482_), .A2(new_n11474_), .B(new_n11468_), .ZN(new_n11483_));
  XOR2_X1    g11399(.A1(new_n11336_), .A2(new_n11330_), .Z(new_n11484_));
  AOI21_X1   g11400(.A1(new_n11339_), .A2(new_n11337_), .B(new_n11325_), .ZN(new_n11485_));
  AOI21_X1   g11401(.A1(new_n11325_), .A2(new_n11484_), .B(new_n11485_), .ZN(new_n11486_));
  INV_X1     g11402(.I(new_n11301_), .ZN(new_n11487_));
  AOI22_X1   g11403(.A1(new_n11003_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n10745_), .ZN(new_n11488_));
  OAI21_X1   g11404(.A1(new_n11488_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n11489_));
  XOR2_X1    g11405(.A1(new_n11489_), .A2(new_n11001_), .Z(new_n11490_));
  INV_X1     g11406(.I(new_n11490_), .ZN(new_n11491_));
  NAND2_X1   g11407(.A1(new_n11491_), .A2(new_n11487_), .ZN(new_n11492_));
  NAND3_X1   g11408(.A1(new_n10783_), .A2(new_n643_), .A3(new_n10780_), .ZN(new_n11493_));
  AOI21_X1   g11409(.A1(new_n11009_), .A2(new_n785_), .B(new_n11002_), .ZN(new_n11494_));
  OAI22_X1   g11410(.A1(new_n10772_), .A2(new_n5966_), .B1(new_n1851_), .B2(new_n10755_), .ZN(new_n11495_));
  OAI21_X1   g11411(.A1(new_n643_), .A2(new_n10762_), .B(new_n11495_), .ZN(new_n11496_));
  AOI21_X1   g11412(.A1(new_n11493_), .A2(new_n11494_), .B(new_n11496_), .ZN(new_n11497_));
  XOR2_X1    g11413(.A1(new_n11497_), .A2(new_n279_), .Z(new_n11498_));
  NOR2_X1    g11414(.A1(new_n10772_), .A2(new_n1851_), .ZN(new_n11499_));
  OAI21_X1   g11415(.A1(new_n10755_), .A2(new_n643_), .B(new_n279_), .ZN(new_n11500_));
  OAI21_X1   g11416(.A1(new_n11499_), .A2(new_n11500_), .B(new_n785_), .ZN(new_n11501_));
  XOR2_X1    g11417(.A1(new_n11501_), .A2(new_n11017_), .Z(new_n11502_));
  NOR2_X1    g11418(.A1(new_n10780_), .A2(new_n1733_), .ZN(new_n11503_));
  NOR2_X1    g11419(.A1(new_n11503_), .A2(new_n279_), .ZN(new_n11504_));
  NAND2_X1   g11420(.A1(new_n11502_), .A2(new_n11504_), .ZN(new_n11505_));
  NOR2_X1    g11421(.A1(new_n11498_), .A2(new_n11505_), .ZN(new_n11506_));
  NOR2_X1    g11422(.A1(new_n11491_), .A2(new_n11487_), .ZN(new_n11507_));
  OAI21_X1   g11423(.A1(new_n11506_), .A2(new_n11507_), .B(new_n11492_), .ZN(new_n11508_));
  XOR2_X1    g11424(.A1(new_n11300_), .A2(new_n11303_), .Z(new_n11509_));
  INV_X1     g11425(.I(new_n11509_), .ZN(new_n11510_));
  OAI22_X1   g11426(.A1(new_n10725_), .A2(new_n643_), .B1(new_n5967_), .B2(new_n11047_), .ZN(new_n11511_));
  AOI21_X1   g11427(.A1(new_n11511_), .A2(new_n279_), .B(new_n643_), .ZN(new_n11512_));
  XOR2_X1    g11428(.A1(new_n11046_), .A2(new_n11512_), .Z(new_n11513_));
  OR2_X2     g11429(.A1(new_n11513_), .A2(new_n11510_), .Z(new_n11514_));
  NAND2_X1   g11430(.A1(new_n11514_), .A2(new_n11508_), .ZN(new_n11515_));
  NAND2_X1   g11431(.A1(new_n11513_), .A2(new_n11510_), .ZN(new_n11516_));
  NAND2_X1   g11432(.A1(new_n11515_), .A2(new_n11516_), .ZN(new_n11517_));
  AOI22_X1   g11433(.A1(new_n10794_), .A2(new_n785_), .B1(new_n5968_), .B2(new_n11065_), .ZN(new_n11518_));
  OAI21_X1   g11434(.A1(new_n11518_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n11519_));
  XOR2_X1    g11435(.A1(new_n11064_), .A2(new_n11519_), .Z(new_n11520_));
  INV_X1     g11436(.I(new_n11520_), .ZN(new_n11521_));
  NAND2_X1   g11437(.A1(new_n11517_), .A2(new_n11521_), .ZN(new_n11522_));
  NOR2_X1    g11438(.A1(new_n11295_), .A2(new_n11304_), .ZN(new_n11523_));
  OAI22_X1   g11439(.A1(new_n11517_), .A2(new_n11521_), .B1(new_n11306_), .B2(new_n11523_), .ZN(new_n11524_));
  AND2_X2    g11440(.A1(new_n11524_), .A2(new_n11522_), .Z(new_n11525_));
  XNOR2_X1   g11441(.A1(new_n11287_), .A2(new_n11099_), .ZN(new_n11526_));
  NOR2_X1    g11442(.A1(new_n11307_), .A2(new_n11288_), .ZN(new_n11527_));
  MUX2_X1    g11443(.I0(new_n11527_), .I1(new_n11526_), .S(new_n11306_), .Z(new_n11528_));
  AOI22_X1   g11444(.A1(new_n11141_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n10691_), .ZN(new_n11529_));
  OAI21_X1   g11445(.A1(new_n11529_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n11530_));
  XOR2_X1    g11446(.A1(new_n11333_), .A2(new_n11530_), .Z(new_n11531_));
  NAND2_X1   g11447(.A1(new_n11531_), .A2(new_n11528_), .ZN(new_n11532_));
  INV_X1     g11448(.I(new_n11532_), .ZN(new_n11533_));
  NOR2_X1    g11449(.A1(new_n11531_), .A2(new_n11528_), .ZN(new_n11534_));
  INV_X1     g11450(.I(new_n11534_), .ZN(new_n11535_));
  OAI21_X1   g11451(.A1(new_n11525_), .A2(new_n11533_), .B(new_n11535_), .ZN(new_n11536_));
  INV_X1     g11452(.I(new_n11308_), .ZN(new_n11537_));
  XNOR2_X1   g11453(.A1(new_n11312_), .A2(new_n11309_), .ZN(new_n11538_));
  NOR2_X1    g11454(.A1(new_n11538_), .A2(new_n11537_), .ZN(new_n11539_));
  AOI21_X1   g11455(.A1(new_n11314_), .A2(new_n11315_), .B(new_n11308_), .ZN(new_n11540_));
  NOR2_X1    g11456(.A1(new_n11539_), .A2(new_n11540_), .ZN(new_n11541_));
  OAI22_X1   g11457(.A1(new_n10672_), .A2(new_n643_), .B1(new_n5967_), .B2(new_n11159_), .ZN(new_n11542_));
  AOI21_X1   g11458(.A1(new_n11542_), .A2(new_n279_), .B(new_n643_), .ZN(new_n11543_));
  XNOR2_X1   g11459(.A1(new_n11158_), .A2(new_n11543_), .ZN(new_n11544_));
  INV_X1     g11460(.I(new_n11544_), .ZN(new_n11545_));
  NOR2_X1    g11461(.A1(new_n11541_), .A2(new_n11545_), .ZN(new_n11546_));
  INV_X1     g11462(.I(new_n11546_), .ZN(new_n11547_));
  AND2_X2    g11463(.A1(new_n11536_), .A2(new_n11547_), .Z(new_n11548_));
  NOR3_X1    g11464(.A1(new_n11539_), .A2(new_n11540_), .A3(new_n11544_), .ZN(new_n11549_));
  NOR2_X1    g11465(.A1(new_n11548_), .A2(new_n11549_), .ZN(new_n11550_));
  XOR2_X1    g11466(.A1(new_n11321_), .A2(new_n11318_), .Z(new_n11551_));
  INV_X1     g11467(.I(new_n11324_), .ZN(new_n11552_));
  OAI21_X1   g11468(.A1(new_n11552_), .A2(new_n11323_), .B(new_n11317_), .ZN(new_n11553_));
  OAI21_X1   g11469(.A1(new_n11317_), .A2(new_n11551_), .B(new_n11553_), .ZN(new_n11554_));
  OAI22_X1   g11470(.A1(new_n11176_), .A2(new_n5967_), .B1(new_n10658_), .B2(new_n643_), .ZN(new_n11555_));
  AOI21_X1   g11471(.A1(new_n11555_), .A2(new_n279_), .B(new_n643_), .ZN(new_n11556_));
  XOR2_X1    g11472(.A1(new_n11175_), .A2(new_n11556_), .Z(new_n11557_));
  NOR2_X1    g11473(.A1(new_n11554_), .A2(new_n11557_), .ZN(new_n11558_));
  NAND2_X1   g11474(.A1(new_n11554_), .A2(new_n11557_), .ZN(new_n11559_));
  INV_X1     g11475(.I(new_n11559_), .ZN(new_n11560_));
  NOR2_X1    g11476(.A1(new_n11560_), .A2(new_n11558_), .ZN(new_n11561_));
  NAND2_X1   g11477(.A1(new_n11550_), .A2(new_n11561_), .ZN(new_n11562_));
  NOR2_X1    g11478(.A1(new_n11562_), .A2(new_n11486_), .ZN(new_n11563_));
  OAI22_X1   g11479(.A1(new_n10819_), .A2(new_n5967_), .B1(new_n11214_), .B2(new_n643_), .ZN(new_n11564_));
  AOI21_X1   g11480(.A1(new_n11564_), .A2(new_n279_), .B(new_n643_), .ZN(new_n11565_));
  XOR2_X1    g11481(.A1(new_n11224_), .A2(new_n11565_), .Z(new_n11566_));
  OR2_X2     g11482(.A1(new_n11559_), .A2(new_n11566_), .Z(new_n11567_));
  AOI21_X1   g11483(.A1(new_n11562_), .A2(new_n11486_), .B(new_n11567_), .ZN(new_n11568_));
  OR2_X2     g11484(.A1(new_n11568_), .A2(new_n11563_), .Z(new_n11569_));
  INV_X1     g11485(.I(new_n11569_), .ZN(new_n11570_));
  AOI21_X1   g11486(.A1(new_n11474_), .A2(new_n11482_), .B(new_n11570_), .ZN(new_n11571_));
  NAND3_X1   g11487(.A1(new_n11571_), .A2(new_n11463_), .A3(new_n11483_), .ZN(new_n11572_));
  INV_X1     g11488(.I(new_n11572_), .ZN(new_n11573_));
  NAND2_X1   g11489(.A1(new_n11571_), .A2(new_n11483_), .ZN(new_n11574_));
  NAND2_X1   g11490(.A1(new_n11574_), .A2(new_n11462_), .ZN(new_n11575_));
  INV_X1     g11491(.I(new_n11480_), .ZN(new_n11576_));
  OAI22_X1   g11492(.A1(new_n11386_), .A2(new_n5967_), .B1(new_n643_), .B2(new_n10633_), .ZN(new_n11577_));
  AOI21_X1   g11493(.A1(new_n11577_), .A2(new_n279_), .B(new_n643_), .ZN(new_n11578_));
  XOR2_X1    g11494(.A1(new_n11385_), .A2(new_n11578_), .Z(new_n11579_));
  NOR2_X1    g11495(.A1(new_n11576_), .A2(new_n11579_), .ZN(new_n11580_));
  AOI21_X1   g11496(.A1(new_n11575_), .A2(new_n11580_), .B(new_n11573_), .ZN(new_n11581_));
  AOI22_X1   g11497(.A1(new_n10630_), .A2(new_n785_), .B1(new_n5968_), .B2(new_n11446_), .ZN(new_n11582_));
  NOR2_X1    g11498(.A1(new_n11582_), .A2(\a[14] ), .ZN(new_n11583_));
  NOR2_X1    g11499(.A1(new_n11583_), .A2(new_n643_), .ZN(new_n11584_));
  XOR2_X1    g11500(.A1(new_n11445_), .A2(new_n11584_), .Z(new_n11585_));
  NOR2_X1    g11501(.A1(new_n11581_), .A2(new_n11585_), .ZN(new_n11586_));
  INV_X1     g11502(.I(new_n11370_), .ZN(new_n11587_));
  NAND2_X1   g11503(.A1(new_n11254_), .A2(new_n11251_), .ZN(new_n11588_));
  NOR2_X1    g11504(.A1(new_n11254_), .A2(new_n11251_), .ZN(new_n11589_));
  INV_X1     g11505(.I(new_n11589_), .ZN(new_n11590_));
  AND2_X2    g11506(.A1(new_n11590_), .A2(new_n11588_), .Z(new_n11591_));
  XOR2_X1    g11507(.A1(new_n11591_), .A2(new_n11587_), .Z(new_n11592_));
  AOI21_X1   g11508(.A1(new_n11581_), .A2(new_n11585_), .B(new_n11592_), .ZN(new_n11593_));
  XNOR2_X1   g11509(.A1(new_n11254_), .A2(new_n11251_), .ZN(new_n11594_));
  OR3_X2     g11510(.A1(new_n11277_), .A2(new_n11589_), .A3(new_n11594_), .Z(new_n11595_));
  NOR2_X1    g11511(.A1(new_n11254_), .A2(new_n11251_), .ZN(new_n11596_));
  INV_X1     g11512(.I(new_n11596_), .ZN(new_n11597_));
  NAND2_X1   g11513(.A1(new_n11595_), .A2(new_n11597_), .ZN(new_n11598_));
  NAND2_X1   g11514(.A1(new_n11598_), .A2(new_n11370_), .ZN(new_n11599_));
  INV_X1     g11515(.I(new_n11599_), .ZN(new_n11600_));
  NOR2_X1    g11516(.A1(new_n11598_), .A2(new_n11370_), .ZN(new_n11601_));
  NOR3_X1    g11517(.A1(new_n10832_), .A2(new_n10835_), .A3(new_n10630_), .ZN(new_n11602_));
  NOR2_X1    g11518(.A1(new_n10631_), .A2(new_n10831_), .ZN(new_n11603_));
  OAI21_X1   g11519(.A1(new_n11602_), .A2(new_n11603_), .B(new_n10843_), .ZN(new_n11604_));
  NAND2_X1   g11520(.A1(new_n10836_), .A2(new_n10847_), .ZN(new_n11605_));
  NAND2_X1   g11521(.A1(new_n11605_), .A2(new_n10844_), .ZN(new_n11606_));
  NAND2_X1   g11522(.A1(new_n11606_), .A2(new_n11604_), .ZN(new_n11607_));
  NAND2_X1   g11523(.A1(new_n10630_), .A2(new_n10833_), .ZN(new_n11608_));
  AOI22_X1   g11524(.A1(new_n785_), .A2(new_n10843_), .B1(new_n11608_), .B2(new_n5968_), .ZN(new_n11609_));
  OAI21_X1   g11525(.A1(new_n11609_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n11610_));
  XOR2_X1    g11526(.A1(new_n11607_), .A2(new_n11610_), .Z(new_n11611_));
  OAI21_X1   g11527(.A1(new_n11600_), .A2(new_n11601_), .B(new_n11611_), .ZN(new_n11612_));
  OAI21_X1   g11528(.A1(new_n11586_), .A2(new_n11593_), .B(new_n11612_), .ZN(new_n11613_));
  INV_X1     g11529(.I(new_n11601_), .ZN(new_n11614_));
  NAND2_X1   g11530(.A1(new_n11614_), .A2(new_n11599_), .ZN(new_n11615_));
  NOR2_X1    g11531(.A1(new_n11615_), .A2(new_n11611_), .ZN(new_n11616_));
  INV_X1     g11532(.I(new_n11616_), .ZN(new_n11617_));
  NAND2_X1   g11533(.A1(new_n11371_), .A2(new_n11278_), .ZN(new_n11618_));
  NOR2_X1    g11534(.A1(new_n11234_), .A2(new_n11389_), .ZN(new_n11619_));
  NAND2_X1   g11535(.A1(new_n11618_), .A2(new_n11619_), .ZN(new_n11620_));
  INV_X1     g11536(.I(new_n11619_), .ZN(new_n11621_));
  NAND3_X1   g11537(.A1(new_n11371_), .A2(new_n11278_), .A3(new_n11621_), .ZN(new_n11622_));
  AOI21_X1   g11538(.A1(new_n11620_), .A2(new_n11622_), .B(new_n11275_), .ZN(new_n11623_));
  INV_X1     g11539(.I(new_n11623_), .ZN(new_n11624_));
  NAND3_X1   g11540(.A1(new_n11620_), .A2(new_n11275_), .A3(new_n11622_), .ZN(new_n11625_));
  INV_X1     g11541(.I(new_n10849_), .ZN(new_n11626_));
  XOR2_X1    g11542(.A1(new_n10856_), .A2(new_n10843_), .Z(new_n11627_));
  NOR2_X1    g11543(.A1(new_n11626_), .A2(new_n11627_), .ZN(new_n11628_));
  INV_X1     g11544(.I(new_n10861_), .ZN(new_n11629_));
  AOI21_X1   g11545(.A1(new_n10859_), .A2(new_n11629_), .B(new_n10849_), .ZN(new_n11630_));
  NOR2_X1    g11546(.A1(new_n11628_), .A2(new_n11630_), .ZN(new_n11631_));
  NAND2_X1   g11547(.A1(new_n10843_), .A2(new_n10630_), .ZN(new_n11632_));
  AOI22_X1   g11548(.A1(new_n11632_), .A2(new_n5968_), .B1(new_n10857_), .B2(new_n785_), .ZN(new_n11633_));
  OAI21_X1   g11549(.A1(new_n11633_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n11634_));
  XNOR2_X1   g11550(.A1(new_n11631_), .A2(new_n11634_), .ZN(new_n11635_));
  INV_X1     g11551(.I(new_n11635_), .ZN(new_n11636_));
  NAND3_X1   g11552(.A1(new_n11624_), .A2(new_n11625_), .A3(new_n11636_), .ZN(new_n11637_));
  INV_X1     g11553(.I(new_n11625_), .ZN(new_n11638_));
  OAI21_X1   g11554(.A1(new_n11638_), .A2(new_n11623_), .B(new_n11635_), .ZN(new_n11639_));
  NAND4_X1   g11555(.A1(new_n11617_), .A2(new_n11613_), .A3(new_n11637_), .A4(new_n11639_), .ZN(new_n11640_));
  NOR2_X1    g11556(.A1(new_n11640_), .A2(new_n11459_), .ZN(new_n11641_));
  NAND2_X1   g11557(.A1(new_n10625_), .A2(new_n10856_), .ZN(new_n11642_));
  NAND2_X1   g11558(.A1(new_n10870_), .A2(new_n10857_), .ZN(new_n11643_));
  AOI21_X1   g11559(.A1(new_n11642_), .A2(new_n11643_), .B(new_n11627_), .ZN(new_n11644_));
  NAND2_X1   g11560(.A1(new_n11644_), .A2(new_n11626_), .ZN(new_n11645_));
  INV_X1     g11561(.I(new_n11645_), .ZN(new_n11646_));
  NOR2_X1    g11562(.A1(new_n11644_), .A2(new_n11626_), .ZN(new_n11647_));
  NOR2_X1    g11563(.A1(new_n11646_), .A2(new_n11647_), .ZN(new_n11648_));
  OAI22_X1   g11564(.A1(new_n10870_), .A2(new_n643_), .B1(new_n5967_), .B2(new_n10861_), .ZN(new_n11649_));
  AOI21_X1   g11565(.A1(new_n11649_), .A2(new_n279_), .B(new_n643_), .ZN(new_n11650_));
  XOR2_X1    g11566(.A1(new_n11648_), .A2(new_n11650_), .Z(new_n11651_));
  NOR2_X1    g11567(.A1(new_n11639_), .A2(new_n11651_), .ZN(new_n11652_));
  INV_X1     g11568(.I(new_n11652_), .ZN(new_n11653_));
  AOI21_X1   g11569(.A1(new_n11640_), .A2(new_n11459_), .B(new_n11653_), .ZN(new_n11654_));
  NOR2_X1    g11570(.A1(new_n11654_), .A2(new_n11641_), .ZN(new_n11655_));
  INV_X1     g11571(.I(new_n11655_), .ZN(new_n11656_));
  INV_X1     g11572(.I(new_n11455_), .ZN(new_n11657_));
  AOI21_X1   g11573(.A1(new_n11392_), .A2(new_n11657_), .B(new_n11456_), .ZN(new_n11658_));
  NAND2_X1   g11574(.A1(new_n11423_), .A2(new_n11397_), .ZN(new_n11659_));
  NOR2_X1    g11575(.A1(new_n11398_), .A2(new_n11414_), .ZN(new_n11660_));
  NOR2_X1    g11576(.A1(new_n11660_), .A2(new_n11413_), .ZN(new_n11661_));
  OAI22_X1   g11577(.A1(new_n10725_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10777_), .ZN(new_n11662_));
  OAI21_X1   g11578(.A1(new_n10696_), .A2(new_n1128_), .B(new_n11662_), .ZN(new_n11663_));
  AOI21_X1   g11579(.A1(new_n11663_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n11664_));
  XOR2_X1    g11580(.A1(new_n11064_), .A2(new_n11664_), .Z(new_n11665_));
  NAND3_X1   g11581(.A1(new_n10783_), .A2(new_n79_), .A3(new_n10780_), .ZN(new_n11666_));
  AOI21_X1   g11582(.A1(new_n11009_), .A2(new_n101_), .B(new_n11002_), .ZN(new_n11667_));
  OAI22_X1   g11583(.A1(new_n10772_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10755_), .ZN(new_n11668_));
  OAI21_X1   g11584(.A1(new_n79_), .A2(new_n10762_), .B(new_n11668_), .ZN(new_n11669_));
  AOI21_X1   g11585(.A1(new_n11666_), .A2(new_n11667_), .B(new_n11669_), .ZN(new_n11670_));
  XOR2_X1    g11586(.A1(new_n11670_), .A2(\a[29] ), .Z(new_n11671_));
  NAND2_X1   g11587(.A1(new_n11407_), .A2(new_n11408_), .ZN(new_n11672_));
  XOR2_X1    g11588(.A1(new_n11671_), .A2(new_n11672_), .Z(new_n11673_));
  XNOR2_X1   g11589(.A1(new_n11665_), .A2(new_n11673_), .ZN(new_n11674_));
  NOR2_X1    g11590(.A1(new_n11674_), .A2(new_n11661_), .ZN(new_n11675_));
  INV_X1     g11591(.I(new_n11661_), .ZN(new_n11676_));
  NAND2_X1   g11592(.A1(new_n11665_), .A2(new_n11673_), .ZN(new_n11677_));
  NOR2_X1    g11593(.A1(new_n11665_), .A2(new_n11673_), .ZN(new_n11678_));
  INV_X1     g11594(.I(new_n11678_), .ZN(new_n11679_));
  AOI21_X1   g11595(.A1(new_n11677_), .A2(new_n11679_), .B(new_n11676_), .ZN(new_n11680_));
  NOR2_X1    g11596(.A1(new_n11680_), .A2(new_n11675_), .ZN(new_n11681_));
  OAI22_X1   g11597(.A1(new_n11176_), .A2(new_n4981_), .B1(new_n10658_), .B2(new_n1239_), .ZN(new_n11682_));
  AOI21_X1   g11598(.A1(new_n11682_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n11683_));
  XOR2_X1    g11599(.A1(new_n11175_), .A2(new_n11683_), .Z(new_n11684_));
  NOR2_X1    g11600(.A1(new_n11681_), .A2(new_n11684_), .ZN(new_n11685_));
  XOR2_X1    g11601(.A1(new_n11659_), .A2(new_n11685_), .Z(new_n11686_));
  XOR2_X1    g11602(.A1(new_n11686_), .A2(new_n11421_), .Z(new_n11687_));
  AOI22_X1   g11603(.A1(new_n10638_), .A2(new_n4717_), .B1(new_n5337_), .B2(new_n11269_), .ZN(new_n11688_));
  NOR2_X1    g11604(.A1(new_n11688_), .A2(\a[20] ), .ZN(new_n11689_));
  NOR2_X1    g11605(.A1(new_n11689_), .A2(new_n5398_), .ZN(new_n11690_));
  XNOR2_X1   g11606(.A1(new_n11268_), .A2(new_n11690_), .ZN(new_n11691_));
  INV_X1     g11607(.I(new_n11691_), .ZN(new_n11692_));
  NOR2_X1    g11608(.A1(new_n11687_), .A2(new_n11692_), .ZN(new_n11693_));
  XOR2_X1    g11609(.A1(new_n11686_), .A2(new_n11422_), .Z(new_n11694_));
  NOR2_X1    g11610(.A1(new_n11694_), .A2(new_n11691_), .ZN(new_n11695_));
  NOR2_X1    g11611(.A1(new_n11693_), .A2(new_n11695_), .ZN(new_n11696_));
  NOR3_X1    g11612(.A1(new_n11696_), .A2(new_n11436_), .A3(new_n11438_), .ZN(new_n11697_));
  NOR2_X1    g11613(.A1(new_n11435_), .A2(new_n11432_), .ZN(new_n11698_));
  OAI21_X1   g11614(.A1(new_n11697_), .A2(new_n11698_), .B(new_n11394_), .ZN(new_n11699_));
  NOR3_X1    g11615(.A1(new_n11697_), .A2(new_n11394_), .A3(new_n11698_), .ZN(new_n11700_));
  INV_X1     g11616(.I(new_n11700_), .ZN(new_n11701_));
  AOI22_X1   g11617(.A1(new_n4660_), .A2(new_n10843_), .B1(new_n11608_), .B2(new_n5421_), .ZN(new_n11702_));
  OAI21_X1   g11618(.A1(new_n11702_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n11703_));
  XOR2_X1    g11619(.A1(new_n11607_), .A2(new_n11703_), .Z(new_n11704_));
  INV_X1     g11620(.I(new_n11704_), .ZN(new_n11705_));
  AOI21_X1   g11621(.A1(new_n11701_), .A2(new_n11699_), .B(new_n11705_), .ZN(new_n11706_));
  INV_X1     g11622(.I(new_n11706_), .ZN(new_n11707_));
  INV_X1     g11623(.I(new_n11699_), .ZN(new_n11708_));
  NOR3_X1    g11624(.A1(new_n11708_), .A2(new_n11700_), .A3(new_n11704_), .ZN(new_n11709_));
  INV_X1     g11625(.I(new_n11709_), .ZN(new_n11710_));
  AOI21_X1   g11626(.A1(new_n11707_), .A2(new_n11710_), .B(new_n11658_), .ZN(new_n11711_));
  NOR3_X1    g11627(.A1(new_n11708_), .A2(new_n11700_), .A3(new_n11705_), .ZN(new_n11712_));
  AOI21_X1   g11628(.A1(new_n11701_), .A2(new_n11699_), .B(new_n11704_), .ZN(new_n11713_));
  OAI21_X1   g11629(.A1(new_n11712_), .A2(new_n11713_), .B(new_n11658_), .ZN(new_n11714_));
  INV_X1     g11630(.I(new_n11714_), .ZN(new_n11715_));
  NAND3_X1   g11631(.A1(new_n10860_), .A2(new_n10862_), .A3(new_n10870_), .ZN(new_n11716_));
  AOI21_X1   g11632(.A1(new_n11626_), .A2(new_n10858_), .B(new_n10870_), .ZN(new_n11717_));
  INV_X1     g11633(.I(new_n11717_), .ZN(new_n11718_));
  AOI21_X1   g11634(.A1(new_n11718_), .A2(new_n11716_), .B(new_n10868_), .ZN(new_n11719_));
  NOR2_X1    g11635(.A1(new_n10863_), .A2(new_n10871_), .ZN(new_n11720_));
  NOR2_X1    g11636(.A1(new_n11720_), .A2(new_n10875_), .ZN(new_n11721_));
  NOR2_X1    g11637(.A1(new_n11721_), .A2(new_n11719_), .ZN(new_n11722_));
  NOR2_X1    g11638(.A1(new_n10870_), .A2(new_n10856_), .ZN(new_n11723_));
  INV_X1     g11639(.I(new_n11723_), .ZN(new_n11724_));
  AOI22_X1   g11640(.A1(new_n11724_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n10875_), .ZN(new_n11725_));
  OAI21_X1   g11641(.A1(new_n11725_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n11726_));
  XNOR2_X1   g11642(.A1(new_n11722_), .A2(new_n11726_), .ZN(new_n11727_));
  INV_X1     g11643(.I(new_n11727_), .ZN(new_n11728_));
  NOR3_X1    g11644(.A1(new_n11715_), .A2(new_n11711_), .A3(new_n11728_), .ZN(new_n11729_));
  OAI21_X1   g11645(.A1(new_n11715_), .A2(new_n11711_), .B(new_n11728_), .ZN(new_n11730_));
  INV_X1     g11646(.I(new_n11730_), .ZN(new_n11731_));
  NOR2_X1    g11647(.A1(new_n11731_), .A2(new_n11729_), .ZN(new_n11732_));
  OAI21_X1   g11648(.A1(new_n11658_), .A2(new_n11706_), .B(new_n11710_), .ZN(new_n11733_));
  INV_X1     g11649(.I(new_n11733_), .ZN(new_n11734_));
  INV_X1     g11650(.I(new_n11693_), .ZN(new_n11735_));
  OAI21_X1   g11651(.A1(new_n11696_), .A2(new_n11435_), .B(new_n11432_), .ZN(new_n11736_));
  AOI21_X1   g11652(.A1(new_n11696_), .A2(new_n11435_), .B(new_n11394_), .ZN(new_n11737_));
  INV_X1     g11653(.I(new_n11659_), .ZN(new_n11738_));
  INV_X1     g11654(.I(new_n11681_), .ZN(new_n11739_));
  NAND2_X1   g11655(.A1(new_n11738_), .A2(new_n11739_), .ZN(new_n11740_));
  NOR2_X1    g11656(.A1(new_n11421_), .A2(new_n11684_), .ZN(new_n11741_));
  OAI21_X1   g11657(.A1(new_n11738_), .A2(new_n11739_), .B(new_n11741_), .ZN(new_n11742_));
  NAND2_X1   g11658(.A1(new_n11742_), .A2(new_n11740_), .ZN(new_n11743_));
  OAI21_X1   g11659(.A1(new_n11661_), .A2(new_n11678_), .B(new_n11677_), .ZN(new_n11744_));
  AOI22_X1   g11660(.A1(new_n10794_), .A2(new_n4767_), .B1(new_n4613_), .B2(new_n10809_), .ZN(new_n11745_));
  AOI21_X1   g11661(.A1(new_n117_), .A2(new_n10691_), .B(new_n11745_), .ZN(new_n11746_));
  OAI21_X1   g11662(.A1(new_n11746_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n11747_));
  XOR2_X1    g11663(.A1(new_n11333_), .A2(new_n11747_), .Z(new_n11748_));
  NAND3_X1   g11664(.A1(new_n11671_), .A2(new_n11407_), .A3(new_n11408_), .ZN(new_n11749_));
  OAI21_X1   g11665(.A1(new_n4527_), .A2(new_n10762_), .B(new_n11404_), .ZN(new_n11750_));
  OAI21_X1   g11666(.A1(new_n79_), .A2(new_n10777_), .B(new_n11750_), .ZN(new_n11751_));
  AOI21_X1   g11667(.A1(new_n11751_), .A2(new_n72_), .B(new_n79_), .ZN(new_n11752_));
  XOR2_X1    g11668(.A1(new_n11752_), .A2(new_n11188_), .Z(new_n11753_));
  NOR2_X1    g11669(.A1(new_n10780_), .A2(new_n935_), .ZN(new_n11754_));
  NOR2_X1    g11670(.A1(new_n11753_), .A2(new_n11754_), .ZN(new_n11755_));
  INV_X1     g11671(.I(new_n11755_), .ZN(new_n11756_));
  NAND2_X1   g11672(.A1(new_n11753_), .A2(new_n11754_), .ZN(new_n11757_));
  AOI21_X1   g11673(.A1(new_n11756_), .A2(new_n11757_), .B(new_n11749_), .ZN(new_n11758_));
  INV_X1     g11674(.I(new_n11749_), .ZN(new_n11759_));
  XNOR2_X1   g11675(.A1(new_n11753_), .A2(new_n11754_), .ZN(new_n11760_));
  NOR2_X1    g11676(.A1(new_n11760_), .A2(new_n11759_), .ZN(new_n11761_));
  NOR2_X1    g11677(.A1(new_n11761_), .A2(new_n11758_), .ZN(new_n11762_));
  XNOR2_X1   g11678(.A1(new_n11762_), .A2(new_n11748_), .ZN(new_n11763_));
  INV_X1     g11679(.I(new_n11748_), .ZN(new_n11764_));
  NAND2_X1   g11680(.A1(new_n11764_), .A2(new_n11762_), .ZN(new_n11765_));
  OAI21_X1   g11681(.A1(new_n11758_), .A2(new_n11761_), .B(new_n11748_), .ZN(new_n11766_));
  NAND2_X1   g11682(.A1(new_n11765_), .A2(new_n11766_), .ZN(new_n11767_));
  MUX2_X1    g11683(.I0(new_n11767_), .I1(new_n11763_), .S(new_n11744_), .Z(new_n11768_));
  OAI22_X1   g11684(.A1(new_n10819_), .A2(new_n4981_), .B1(new_n11214_), .B2(new_n1239_), .ZN(new_n11769_));
  AOI21_X1   g11685(.A1(new_n11769_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n11770_));
  XOR2_X1    g11686(.A1(new_n11224_), .A2(new_n11770_), .Z(new_n11771_));
  INV_X1     g11687(.I(new_n11771_), .ZN(new_n11772_));
  XOR2_X1    g11688(.A1(new_n11768_), .A2(new_n11772_), .Z(new_n11773_));
  INV_X1     g11689(.I(new_n11773_), .ZN(new_n11774_));
  XOR2_X1    g11690(.A1(new_n11768_), .A2(new_n11771_), .Z(new_n11775_));
  NOR2_X1    g11691(.A1(new_n11743_), .A2(new_n11775_), .ZN(new_n11776_));
  AOI21_X1   g11692(.A1(new_n11743_), .A2(new_n11774_), .B(new_n11776_), .ZN(new_n11777_));
  OAI22_X1   g11693(.A1(new_n11386_), .A2(new_n5336_), .B1(new_n5398_), .B2(new_n10633_), .ZN(new_n11778_));
  AOI21_X1   g11694(.A1(new_n11778_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n11779_));
  XOR2_X1    g11695(.A1(new_n11385_), .A2(new_n11779_), .Z(new_n11780_));
  NOR2_X1    g11696(.A1(new_n11777_), .A2(new_n11780_), .ZN(new_n11781_));
  INV_X1     g11697(.I(new_n11781_), .ZN(new_n11782_));
  AOI21_X1   g11698(.A1(new_n11737_), .A2(new_n11736_), .B(new_n11782_), .ZN(new_n11783_));
  NAND2_X1   g11699(.A1(new_n11737_), .A2(new_n11736_), .ZN(new_n11784_));
  NOR2_X1    g11700(.A1(new_n11784_), .A2(new_n11781_), .ZN(new_n11785_));
  OAI21_X1   g11701(.A1(new_n11785_), .A2(new_n11783_), .B(new_n11735_), .ZN(new_n11786_));
  NOR3_X1    g11702(.A1(new_n11785_), .A2(new_n11735_), .A3(new_n11783_), .ZN(new_n11787_));
  INV_X1     g11703(.I(new_n11787_), .ZN(new_n11788_));
  AOI22_X1   g11704(.A1(new_n11632_), .A2(new_n5421_), .B1(new_n10857_), .B2(new_n4660_), .ZN(new_n11789_));
  OAI21_X1   g11705(.A1(new_n11789_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n11790_));
  XNOR2_X1   g11706(.A1(new_n11631_), .A2(new_n11790_), .ZN(new_n11791_));
  NAND3_X1   g11707(.A1(new_n11788_), .A2(new_n11786_), .A3(new_n11791_), .ZN(new_n11792_));
  INV_X1     g11708(.I(new_n11786_), .ZN(new_n11793_));
  INV_X1     g11709(.I(new_n11791_), .ZN(new_n11794_));
  OAI21_X1   g11710(.A1(new_n11793_), .A2(new_n11787_), .B(new_n11794_), .ZN(new_n11795_));
  NAND2_X1   g11711(.A1(new_n11795_), .A2(new_n11792_), .ZN(new_n11796_));
  XOR2_X1    g11712(.A1(new_n11796_), .A2(new_n11734_), .Z(new_n11797_));
  XNOR2_X1   g11713(.A1(new_n10881_), .A2(new_n10868_), .ZN(new_n11798_));
  INV_X1     g11714(.I(new_n11798_), .ZN(new_n11799_));
  NAND2_X1   g11715(.A1(new_n10874_), .A2(new_n11799_), .ZN(new_n11800_));
  OAI21_X1   g11716(.A1(new_n10883_), .A2(new_n10885_), .B(new_n10873_), .ZN(new_n11801_));
  NAND2_X1   g11717(.A1(new_n11800_), .A2(new_n11801_), .ZN(new_n11802_));
  NOR2_X1    g11718(.A1(new_n10870_), .A2(new_n10868_), .ZN(new_n11803_));
  OAI22_X1   g11719(.A1(new_n11803_), .A2(new_n5967_), .B1(new_n643_), .B2(new_n10881_), .ZN(new_n11804_));
  AOI21_X1   g11720(.A1(new_n11804_), .A2(new_n279_), .B(new_n643_), .ZN(new_n11805_));
  XNOR2_X1   g11721(.A1(new_n11802_), .A2(new_n11805_), .ZN(new_n11806_));
  NOR2_X1    g11722(.A1(new_n11797_), .A2(new_n11806_), .ZN(new_n11807_));
  AND2_X2    g11723(.A1(new_n11795_), .A2(new_n11792_), .Z(new_n11808_));
  NAND2_X1   g11724(.A1(new_n11808_), .A2(new_n11734_), .ZN(new_n11809_));
  NAND2_X1   g11725(.A1(new_n11796_), .A2(new_n11733_), .ZN(new_n11810_));
  INV_X1     g11726(.I(new_n11806_), .ZN(new_n11811_));
  AOI21_X1   g11727(.A1(new_n11809_), .A2(new_n11810_), .B(new_n11811_), .ZN(new_n11812_));
  NOR3_X1    g11728(.A1(new_n11807_), .A2(new_n11729_), .A3(new_n11812_), .ZN(new_n11813_));
  NOR3_X1    g11729(.A1(new_n11813_), .A2(new_n11656_), .A3(new_n11732_), .ZN(new_n11814_));
  INV_X1     g11730(.I(new_n11814_), .ZN(new_n11815_));
  OAI21_X1   g11731(.A1(new_n11813_), .A2(new_n11732_), .B(new_n11656_), .ZN(new_n11816_));
  NAND2_X1   g11732(.A1(new_n11815_), .A2(new_n11816_), .ZN(new_n11817_));
  NAND2_X1   g11733(.A1(new_n11817_), .A2(new_n10989_), .ZN(new_n11818_));
  NOR2_X1    g11734(.A1(new_n11459_), .A2(new_n11651_), .ZN(new_n11819_));
  NAND2_X1   g11735(.A1(new_n11640_), .A2(new_n11819_), .ZN(new_n11820_));
  NAND2_X1   g11736(.A1(new_n11575_), .A2(new_n11580_), .ZN(new_n11821_));
  NAND2_X1   g11737(.A1(new_n11821_), .A2(new_n11572_), .ZN(new_n11822_));
  INV_X1     g11738(.I(new_n11585_), .ZN(new_n11823_));
  NAND2_X1   g11739(.A1(new_n11822_), .A2(new_n11823_), .ZN(new_n11824_));
  INV_X1     g11740(.I(new_n11592_), .ZN(new_n11825_));
  OAI21_X1   g11741(.A1(new_n11822_), .A2(new_n11823_), .B(new_n11825_), .ZN(new_n11826_));
  INV_X1     g11742(.I(new_n11611_), .ZN(new_n11827_));
  AOI21_X1   g11743(.A1(new_n11614_), .A2(new_n11599_), .B(new_n11827_), .ZN(new_n11828_));
  AOI21_X1   g11744(.A1(new_n11826_), .A2(new_n11824_), .B(new_n11828_), .ZN(new_n11829_));
  NAND2_X1   g11745(.A1(new_n11637_), .A2(new_n11639_), .ZN(new_n11830_));
  NOR3_X1    g11746(.A1(new_n11830_), .A2(new_n11829_), .A3(new_n11616_), .ZN(new_n11831_));
  OAI21_X1   g11747(.A1(new_n11459_), .A2(new_n11651_), .B(new_n11831_), .ZN(new_n11832_));
  NAND2_X1   g11748(.A1(new_n11832_), .A2(new_n11820_), .ZN(new_n11833_));
  NAND2_X1   g11749(.A1(new_n11833_), .A2(new_n11639_), .ZN(new_n11834_));
  NAND2_X1   g11750(.A1(new_n11624_), .A2(new_n11625_), .ZN(new_n11835_));
  NAND4_X1   g11751(.A1(new_n11832_), .A2(new_n11835_), .A3(new_n11635_), .A4(new_n11820_), .ZN(new_n11836_));
  NAND2_X1   g11752(.A1(new_n11834_), .A2(new_n11836_), .ZN(new_n11837_));
  INV_X1     g11753(.I(new_n11837_), .ZN(new_n11838_));
  NAND2_X1   g11754(.A1(new_n11581_), .A2(new_n11823_), .ZN(new_n11839_));
  NAND2_X1   g11755(.A1(new_n11822_), .A2(new_n11585_), .ZN(new_n11840_));
  AOI21_X1   g11756(.A1(new_n11840_), .A2(new_n11839_), .B(new_n11587_), .ZN(new_n11841_));
  NOR2_X1    g11757(.A1(new_n11822_), .A2(new_n11585_), .ZN(new_n11842_));
  NOR2_X1    g11758(.A1(new_n11581_), .A2(new_n11823_), .ZN(new_n11843_));
  NOR3_X1    g11759(.A1(new_n11842_), .A2(new_n11370_), .A3(new_n11843_), .ZN(new_n11844_));
  OAI21_X1   g11760(.A1(new_n11844_), .A2(new_n11841_), .B(new_n11591_), .ZN(new_n11845_));
  INV_X1     g11761(.I(new_n11591_), .ZN(new_n11846_));
  OAI21_X1   g11762(.A1(new_n11842_), .A2(new_n11843_), .B(new_n11370_), .ZN(new_n11847_));
  NAND3_X1   g11763(.A1(new_n11840_), .A2(new_n11587_), .A3(new_n11839_), .ZN(new_n11848_));
  NAND3_X1   g11764(.A1(new_n11847_), .A2(new_n11848_), .A3(new_n11846_), .ZN(new_n11849_));
  NAND2_X1   g11765(.A1(new_n11845_), .A2(new_n11849_), .ZN(new_n11850_));
  NOR2_X1    g11766(.A1(new_n11486_), .A2(new_n11566_), .ZN(new_n11851_));
  NAND2_X1   g11767(.A1(new_n11562_), .A2(new_n11851_), .ZN(new_n11852_));
  NOR2_X1    g11768(.A1(new_n11562_), .A2(new_n11851_), .ZN(new_n11853_));
  INV_X1     g11769(.I(new_n11853_), .ZN(new_n11854_));
  AOI21_X1   g11770(.A1(new_n11854_), .A2(new_n11852_), .B(new_n11560_), .ZN(new_n11855_));
  AND3_X2    g11771(.A1(new_n11854_), .A2(new_n11560_), .A3(new_n11852_), .Z(new_n11856_));
  NOR2_X1    g11772(.A1(new_n11856_), .A2(new_n11855_), .ZN(new_n11857_));
  AOI21_X1   g11773(.A1(new_n10652_), .A2(new_n10805_), .B(new_n6757_), .ZN(new_n11858_));
  NOR2_X1    g11774(.A1(new_n10646_), .A2(new_n1078_), .ZN(new_n11859_));
  OAI21_X1   g11775(.A1(new_n11859_), .A2(new_n11858_), .B(new_n294_), .ZN(new_n11860_));
  NAND2_X1   g11776(.A1(new_n11860_), .A2(new_n805_), .ZN(new_n11861_));
  XOR2_X1    g11777(.A1(new_n11246_), .A2(new_n11861_), .Z(new_n11862_));
  XOR2_X1    g11778(.A1(new_n11541_), .A2(new_n11545_), .Z(new_n11863_));
  NAND2_X1   g11779(.A1(new_n11536_), .A2(new_n11863_), .ZN(new_n11864_));
  NOR2_X1    g11780(.A1(new_n11546_), .A2(new_n11549_), .ZN(new_n11865_));
  OR2_X2     g11781(.A1(new_n11536_), .A2(new_n11865_), .Z(new_n11866_));
  NAND2_X1   g11782(.A1(new_n11866_), .A2(new_n11864_), .ZN(new_n11867_));
  INV_X1     g11783(.I(new_n11867_), .ZN(new_n11868_));
  INV_X1     g11784(.I(new_n11562_), .ZN(new_n11869_));
  NOR2_X1    g11785(.A1(new_n11550_), .A2(new_n11561_), .ZN(new_n11870_));
  AOI22_X1   g11786(.A1(new_n10638_), .A2(new_n805_), .B1(new_n6758_), .B2(new_n11269_), .ZN(new_n11871_));
  NOR2_X1    g11787(.A1(new_n11871_), .A2(\a[11] ), .ZN(new_n11872_));
  NOR2_X1    g11788(.A1(new_n11872_), .A2(new_n1078_), .ZN(new_n11873_));
  XNOR2_X1   g11789(.A1(new_n11268_), .A2(new_n11873_), .ZN(new_n11874_));
  INV_X1     g11790(.I(new_n11874_), .ZN(new_n11875_));
  NOR3_X1    g11791(.A1(new_n11869_), .A2(new_n11870_), .A3(new_n11875_), .ZN(new_n11876_));
  INV_X1     g11792(.I(new_n11870_), .ZN(new_n11877_));
  AOI21_X1   g11793(.A1(new_n11877_), .A2(new_n11562_), .B(new_n11874_), .ZN(new_n11878_));
  NOR2_X1    g11794(.A1(new_n11878_), .A2(new_n11876_), .ZN(new_n11879_));
  OAI21_X1   g11795(.A1(new_n11879_), .A2(new_n11868_), .B(new_n11862_), .ZN(new_n11880_));
  INV_X1     g11796(.I(new_n11880_), .ZN(new_n11881_));
  OR2_X2     g11797(.A1(new_n11878_), .A2(new_n11876_), .Z(new_n11882_));
  XNOR2_X1   g11798(.A1(new_n11531_), .A2(new_n11528_), .ZN(new_n11883_));
  NOR2_X1    g11799(.A1(new_n11525_), .A2(new_n11883_), .ZN(new_n11884_));
  NAND2_X1   g11800(.A1(new_n11524_), .A2(new_n11522_), .ZN(new_n11885_));
  AOI21_X1   g11801(.A1(new_n11532_), .A2(new_n11535_), .B(new_n11885_), .ZN(new_n11886_));
  NOR2_X1    g11802(.A1(new_n11884_), .A2(new_n11886_), .ZN(new_n11887_));
  AOI22_X1   g11803(.A1(new_n11003_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n10745_), .ZN(new_n11888_));
  OAI21_X1   g11804(.A1(new_n11888_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n11889_));
  XOR2_X1    g11805(.A1(new_n11889_), .A2(new_n11001_), .Z(new_n11890_));
  NOR2_X1    g11806(.A1(new_n11890_), .A2(new_n11503_), .ZN(new_n11891_));
  INV_X1     g11807(.I(new_n11891_), .ZN(new_n11892_));
  NAND3_X1   g11808(.A1(new_n10783_), .A2(new_n1078_), .A3(new_n10780_), .ZN(new_n11893_));
  AOI21_X1   g11809(.A1(new_n11009_), .A2(new_n805_), .B(new_n11002_), .ZN(new_n11894_));
  OAI22_X1   g11810(.A1(new_n10772_), .A2(new_n6756_), .B1(new_n2258_), .B2(new_n10755_), .ZN(new_n11895_));
  OAI21_X1   g11811(.A1(new_n1078_), .A2(new_n10762_), .B(new_n11895_), .ZN(new_n11896_));
  AOI21_X1   g11812(.A1(new_n11893_), .A2(new_n11894_), .B(new_n11896_), .ZN(new_n11897_));
  XOR2_X1    g11813(.A1(new_n11897_), .A2(\a[11] ), .Z(new_n11898_));
  AOI21_X1   g11814(.A1(new_n10780_), .A2(new_n805_), .B(\a[11] ), .ZN(new_n11899_));
  OAI21_X1   g11815(.A1(new_n10772_), .A2(new_n2258_), .B(new_n11899_), .ZN(new_n11900_));
  AND3_X2    g11816(.A1(new_n11030_), .A2(new_n805_), .A3(new_n11900_), .Z(new_n11901_));
  AOI21_X1   g11817(.A1(new_n805_), .A2(new_n11900_), .B(new_n11030_), .ZN(new_n11902_));
  NOR2_X1    g11818(.A1(new_n10780_), .A2(new_n2573_), .ZN(new_n11903_));
  NOR2_X1    g11819(.A1(new_n11903_), .A2(new_n294_), .ZN(new_n11904_));
  INV_X1     g11820(.I(new_n11904_), .ZN(new_n11905_));
  NOR3_X1    g11821(.A1(new_n11901_), .A2(new_n11902_), .A3(new_n11905_), .ZN(new_n11906_));
  NAND2_X1   g11822(.A1(new_n11898_), .A2(new_n11906_), .ZN(new_n11907_));
  NAND2_X1   g11823(.A1(new_n11890_), .A2(new_n11503_), .ZN(new_n11908_));
  NAND2_X1   g11824(.A1(new_n11907_), .A2(new_n11908_), .ZN(new_n11909_));
  NAND2_X1   g11825(.A1(new_n11909_), .A2(new_n11892_), .ZN(new_n11910_));
  XNOR2_X1   g11826(.A1(new_n11502_), .A2(new_n11504_), .ZN(new_n11911_));
  INV_X1     g11827(.I(new_n11911_), .ZN(new_n11912_));
  OAI22_X1   g11828(.A1(new_n10725_), .A2(new_n1078_), .B1(new_n6757_), .B2(new_n11047_), .ZN(new_n11913_));
  AOI21_X1   g11829(.A1(new_n11913_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n11914_));
  XNOR2_X1   g11830(.A1(new_n11046_), .A2(new_n11914_), .ZN(new_n11915_));
  NAND2_X1   g11831(.A1(new_n11915_), .A2(new_n11912_), .ZN(new_n11916_));
  NAND2_X1   g11832(.A1(new_n11916_), .A2(new_n11910_), .ZN(new_n11917_));
  XOR2_X1    g11833(.A1(new_n11046_), .A2(new_n11914_), .Z(new_n11918_));
  NAND2_X1   g11834(.A1(new_n11918_), .A2(new_n11911_), .ZN(new_n11919_));
  AND2_X2    g11835(.A1(new_n11917_), .A2(new_n11919_), .Z(new_n11920_));
  AOI22_X1   g11836(.A1(new_n10794_), .A2(new_n805_), .B1(new_n6758_), .B2(new_n11065_), .ZN(new_n11921_));
  OAI21_X1   g11837(.A1(new_n11921_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n11922_));
  XOR2_X1    g11838(.A1(new_n11064_), .A2(new_n11922_), .Z(new_n11923_));
  NOR2_X1    g11839(.A1(new_n11920_), .A2(new_n11923_), .ZN(new_n11924_));
  INV_X1     g11840(.I(new_n11506_), .ZN(new_n11925_));
  NAND2_X1   g11841(.A1(new_n11498_), .A2(new_n11505_), .ZN(new_n11926_));
  AOI22_X1   g11842(.A1(new_n11920_), .A2(new_n11923_), .B1(new_n11925_), .B2(new_n11926_), .ZN(new_n11927_));
  NOR2_X1    g11843(.A1(new_n11927_), .A2(new_n11924_), .ZN(new_n11928_));
  XOR2_X1    g11844(.A1(new_n11490_), .A2(new_n11487_), .Z(new_n11929_));
  NOR2_X1    g11845(.A1(new_n11929_), .A2(new_n11925_), .ZN(new_n11930_));
  INV_X1     g11846(.I(new_n11507_), .ZN(new_n11931_));
  AOI21_X1   g11847(.A1(new_n11931_), .A2(new_n11492_), .B(new_n11506_), .ZN(new_n11932_));
  NOR2_X1    g11848(.A1(new_n11932_), .A2(new_n11930_), .ZN(new_n11933_));
  INV_X1     g11849(.I(new_n11933_), .ZN(new_n11934_));
  AOI22_X1   g11850(.A1(new_n11141_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n10691_), .ZN(new_n11935_));
  OAI21_X1   g11851(.A1(new_n11935_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n11936_));
  XOR2_X1    g11852(.A1(new_n11333_), .A2(new_n11936_), .Z(new_n11937_));
  INV_X1     g11853(.I(new_n11937_), .ZN(new_n11938_));
  NOR2_X1    g11854(.A1(new_n11938_), .A2(new_n11934_), .ZN(new_n11939_));
  NAND2_X1   g11855(.A1(new_n11938_), .A2(new_n11934_), .ZN(new_n11940_));
  OAI21_X1   g11856(.A1(new_n11928_), .A2(new_n11939_), .B(new_n11940_), .ZN(new_n11941_));
  XOR2_X1    g11857(.A1(new_n11513_), .A2(new_n11510_), .Z(new_n11942_));
  AND2_X2    g11858(.A1(new_n11942_), .A2(new_n11508_), .Z(new_n11943_));
  AOI21_X1   g11859(.A1(new_n11514_), .A2(new_n11516_), .B(new_n11508_), .ZN(new_n11944_));
  OR2_X2     g11860(.A1(new_n11943_), .A2(new_n11944_), .Z(new_n11945_));
  OAI22_X1   g11861(.A1(new_n10672_), .A2(new_n1078_), .B1(new_n6757_), .B2(new_n11159_), .ZN(new_n11946_));
  AOI21_X1   g11862(.A1(new_n11946_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n11947_));
  XOR2_X1    g11863(.A1(new_n11158_), .A2(new_n11947_), .Z(new_n11948_));
  INV_X1     g11864(.I(new_n11948_), .ZN(new_n11949_));
  NAND2_X1   g11865(.A1(new_n11945_), .A2(new_n11949_), .ZN(new_n11950_));
  NOR2_X1    g11866(.A1(new_n11943_), .A2(new_n11944_), .ZN(new_n11951_));
  NAND2_X1   g11867(.A1(new_n11951_), .A2(new_n11948_), .ZN(new_n11952_));
  INV_X1     g11868(.I(new_n11952_), .ZN(new_n11953_));
  AOI21_X1   g11869(.A1(new_n11941_), .A2(new_n11950_), .B(new_n11953_), .ZN(new_n11954_));
  XOR2_X1    g11870(.A1(new_n11517_), .A2(new_n11295_), .Z(new_n11955_));
  NOR2_X1    g11871(.A1(new_n11955_), .A2(new_n11521_), .ZN(new_n11956_));
  XOR2_X1    g11872(.A1(new_n11517_), .A2(new_n11296_), .Z(new_n11957_));
  NOR2_X1    g11873(.A1(new_n11957_), .A2(new_n11520_), .ZN(new_n11958_));
  OAI21_X1   g11874(.A1(new_n11956_), .A2(new_n11958_), .B(new_n11305_), .ZN(new_n11959_));
  NAND2_X1   g11875(.A1(new_n11957_), .A2(new_n11520_), .ZN(new_n11960_));
  NAND2_X1   g11876(.A1(new_n11955_), .A2(new_n11521_), .ZN(new_n11961_));
  NAND3_X1   g11877(.A1(new_n11960_), .A2(new_n11961_), .A3(new_n11304_), .ZN(new_n11962_));
  OAI22_X1   g11878(.A1(new_n11176_), .A2(new_n6757_), .B1(new_n10658_), .B2(new_n1078_), .ZN(new_n11963_));
  AOI21_X1   g11879(.A1(new_n11963_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n11964_));
  XOR2_X1    g11880(.A1(new_n11175_), .A2(new_n11964_), .Z(new_n11965_));
  INV_X1     g11881(.I(new_n11965_), .ZN(new_n11966_));
  NAND3_X1   g11882(.A1(new_n11959_), .A2(new_n11962_), .A3(new_n11966_), .ZN(new_n11967_));
  AOI21_X1   g11883(.A1(new_n11960_), .A2(new_n11961_), .B(new_n11304_), .ZN(new_n11968_));
  NOR3_X1    g11884(.A1(new_n11956_), .A2(new_n11958_), .A3(new_n11305_), .ZN(new_n11969_));
  OAI21_X1   g11885(.A1(new_n11968_), .A2(new_n11969_), .B(new_n11965_), .ZN(new_n11970_));
  NAND3_X1   g11886(.A1(new_n11970_), .A2(new_n11967_), .A3(new_n11954_), .ZN(new_n11971_));
  NOR2_X1    g11887(.A1(new_n11971_), .A2(new_n11887_), .ZN(new_n11972_));
  AOI21_X1   g11888(.A1(new_n11959_), .A2(new_n11962_), .B(new_n11966_), .ZN(new_n11973_));
  OAI22_X1   g11889(.A1(new_n10819_), .A2(new_n6757_), .B1(new_n11214_), .B2(new_n1078_), .ZN(new_n11974_));
  AOI21_X1   g11890(.A1(new_n11974_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n11975_));
  XOR2_X1    g11891(.A1(new_n11224_), .A2(new_n11975_), .Z(new_n11976_));
  INV_X1     g11892(.I(new_n11976_), .ZN(new_n11977_));
  NAND2_X1   g11893(.A1(new_n11973_), .A2(new_n11977_), .ZN(new_n11978_));
  AOI21_X1   g11894(.A1(new_n11971_), .A2(new_n11887_), .B(new_n11978_), .ZN(new_n11979_));
  NOR2_X1    g11895(.A1(new_n11979_), .A2(new_n11972_), .ZN(new_n11980_));
  INV_X1     g11896(.I(new_n11980_), .ZN(new_n11981_));
  OAI21_X1   g11897(.A1(new_n11882_), .A2(new_n11867_), .B(new_n11981_), .ZN(new_n11982_));
  OR3_X2     g11898(.A1(new_n11881_), .A2(new_n11982_), .A3(new_n11857_), .Z(new_n11983_));
  OAI21_X1   g11899(.A1(new_n11881_), .A2(new_n11982_), .B(new_n11857_), .ZN(new_n11984_));
  NAND3_X1   g11900(.A1(new_n11383_), .A2(new_n11380_), .A3(new_n11264_), .ZN(new_n11985_));
  OAI21_X1   g11901(.A1(new_n11378_), .A2(new_n11374_), .B(new_n10638_), .ZN(new_n11986_));
  NAND2_X1   g11902(.A1(new_n11986_), .A2(new_n11985_), .ZN(new_n11987_));
  OAI22_X1   g11903(.A1(new_n11386_), .A2(new_n6757_), .B1(new_n1078_), .B2(new_n10633_), .ZN(new_n11988_));
  AOI21_X1   g11904(.A1(new_n11988_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n11989_));
  XOR2_X1    g11905(.A1(new_n11987_), .A2(new_n11989_), .Z(new_n11990_));
  NAND2_X1   g11906(.A1(new_n11876_), .A2(new_n11990_), .ZN(new_n11991_));
  INV_X1     g11907(.I(new_n11991_), .ZN(new_n11992_));
  NAND2_X1   g11908(.A1(new_n11984_), .A2(new_n11992_), .ZN(new_n11993_));
  NAND2_X1   g11909(.A1(new_n11993_), .A2(new_n11983_), .ZN(new_n11994_));
  AOI22_X1   g11910(.A1(new_n10630_), .A2(new_n805_), .B1(new_n6758_), .B2(new_n11446_), .ZN(new_n11995_));
  NOR2_X1    g11911(.A1(new_n11995_), .A2(\a[11] ), .ZN(new_n11996_));
  NOR2_X1    g11912(.A1(new_n11996_), .A2(new_n1078_), .ZN(new_n11997_));
  XOR2_X1    g11913(.A1(new_n11445_), .A2(new_n11997_), .Z(new_n11998_));
  INV_X1     g11914(.I(new_n11998_), .ZN(new_n11999_));
  NAND2_X1   g11915(.A1(new_n11994_), .A2(new_n11999_), .ZN(new_n12000_));
  NAND2_X1   g11916(.A1(new_n11474_), .A2(new_n11468_), .ZN(new_n12001_));
  INV_X1     g11917(.I(new_n11468_), .ZN(new_n12002_));
  NAND2_X1   g11918(.A1(new_n11473_), .A2(new_n12002_), .ZN(new_n12003_));
  AND2_X2    g11919(.A1(new_n12001_), .A2(new_n12003_), .Z(new_n12004_));
  INV_X1     g11920(.I(new_n12004_), .ZN(new_n12005_));
  XOR2_X1    g11921(.A1(new_n11569_), .A2(new_n12005_), .Z(new_n12006_));
  OAI21_X1   g11922(.A1(new_n11994_), .A2(new_n11999_), .B(new_n12006_), .ZN(new_n12007_));
  NAND2_X1   g11923(.A1(new_n12007_), .A2(new_n12000_), .ZN(new_n12008_));
  XOR2_X1    g11924(.A1(new_n11473_), .A2(new_n11468_), .Z(new_n12009_));
  NOR2_X1    g11925(.A1(new_n11482_), .A2(new_n12009_), .ZN(new_n12010_));
  XOR2_X1    g11926(.A1(new_n12010_), .A2(new_n12003_), .Z(new_n12011_));
  OR2_X2     g11927(.A1(new_n12011_), .A2(new_n11569_), .Z(new_n12012_));
  NAND2_X1   g11928(.A1(new_n12011_), .A2(new_n11569_), .ZN(new_n12013_));
  NAND2_X1   g11929(.A1(new_n12012_), .A2(new_n12013_), .ZN(new_n12014_));
  AOI22_X1   g11930(.A1(new_n805_), .A2(new_n10843_), .B1(new_n11608_), .B2(new_n6758_), .ZN(new_n12015_));
  OAI21_X1   g11931(.A1(new_n12015_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n12016_));
  XOR2_X1    g11932(.A1(new_n11607_), .A2(new_n12016_), .Z(new_n12017_));
  NAND2_X1   g11933(.A1(new_n12014_), .A2(new_n12017_), .ZN(new_n12018_));
  NAND2_X1   g11934(.A1(new_n12008_), .A2(new_n12018_), .ZN(new_n12019_));
  NOR2_X1    g11935(.A1(new_n12014_), .A2(new_n12017_), .ZN(new_n12020_));
  INV_X1     g11936(.I(new_n12020_), .ZN(new_n12021_));
  NAND2_X1   g11937(.A1(new_n12019_), .A2(new_n12021_), .ZN(new_n12022_));
  INV_X1     g11938(.I(new_n11579_), .ZN(new_n12023_));
  NAND3_X1   g11939(.A1(new_n11574_), .A2(new_n11463_), .A3(new_n12023_), .ZN(new_n12024_));
  NAND2_X1   g11940(.A1(new_n11463_), .A2(new_n12023_), .ZN(new_n12025_));
  NAND3_X1   g11941(.A1(new_n11571_), .A2(new_n12025_), .A3(new_n11483_), .ZN(new_n12026_));
  NAND2_X1   g11942(.A1(new_n12024_), .A2(new_n12026_), .ZN(new_n12027_));
  NAND2_X1   g11943(.A1(new_n12027_), .A2(new_n11576_), .ZN(new_n12028_));
  NAND3_X1   g11944(.A1(new_n12024_), .A2(new_n11480_), .A3(new_n12026_), .ZN(new_n12029_));
  AOI22_X1   g11945(.A1(new_n11632_), .A2(new_n6758_), .B1(new_n10857_), .B2(new_n805_), .ZN(new_n12030_));
  OAI21_X1   g11946(.A1(new_n12030_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n12031_));
  XNOR2_X1   g11947(.A1(new_n11631_), .A2(new_n12031_), .ZN(new_n12032_));
  INV_X1     g11948(.I(new_n12032_), .ZN(new_n12033_));
  NAND3_X1   g11949(.A1(new_n12028_), .A2(new_n12029_), .A3(new_n12033_), .ZN(new_n12034_));
  NAND2_X1   g11950(.A1(new_n12028_), .A2(new_n12029_), .ZN(new_n12035_));
  NAND2_X1   g11951(.A1(new_n12035_), .A2(new_n12032_), .ZN(new_n12036_));
  NAND2_X1   g11952(.A1(new_n12036_), .A2(new_n12034_), .ZN(new_n12037_));
  NOR2_X1    g11953(.A1(new_n12022_), .A2(new_n12037_), .ZN(new_n12038_));
  NAND2_X1   g11954(.A1(new_n11850_), .A2(new_n12038_), .ZN(new_n12039_));
  OAI22_X1   g11955(.A1(new_n10870_), .A2(new_n1078_), .B1(new_n6757_), .B2(new_n10861_), .ZN(new_n12040_));
  AOI21_X1   g11956(.A1(new_n12040_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n12041_));
  XOR2_X1    g11957(.A1(new_n11648_), .A2(new_n12041_), .Z(new_n12042_));
  NOR2_X1    g11958(.A1(new_n12036_), .A2(new_n12042_), .ZN(new_n12043_));
  OAI21_X1   g11959(.A1(new_n11850_), .A2(new_n12038_), .B(new_n12043_), .ZN(new_n12044_));
  NOR2_X1    g11960(.A1(new_n11593_), .A2(new_n11586_), .ZN(new_n12045_));
  AOI21_X1   g11961(.A1(new_n11617_), .A2(new_n11612_), .B(new_n12045_), .ZN(new_n12046_));
  NAND3_X1   g11962(.A1(new_n11614_), .A2(new_n11599_), .A3(new_n11611_), .ZN(new_n12047_));
  NAND2_X1   g11963(.A1(new_n11615_), .A2(new_n11827_), .ZN(new_n12048_));
  NAND2_X1   g11964(.A1(new_n12048_), .A2(new_n12047_), .ZN(new_n12049_));
  AOI21_X1   g11965(.A1(new_n12045_), .A2(new_n12049_), .B(new_n12046_), .ZN(new_n12050_));
  AOI22_X1   g11966(.A1(new_n11724_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n10875_), .ZN(new_n12051_));
  OAI21_X1   g11967(.A1(new_n12051_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n12052_));
  XNOR2_X1   g11968(.A1(new_n11722_), .A2(new_n12052_), .ZN(new_n12053_));
  AOI22_X1   g11969(.A1(new_n12044_), .A2(new_n12039_), .B1(new_n12050_), .B2(new_n12053_), .ZN(new_n12054_));
  NOR2_X1    g11970(.A1(new_n12050_), .A2(new_n12053_), .ZN(new_n12055_));
  NOR2_X1    g11971(.A1(new_n12054_), .A2(new_n12055_), .ZN(new_n12056_));
  NAND2_X1   g11972(.A1(new_n11617_), .A2(new_n11613_), .ZN(new_n12057_));
  OAI22_X1   g11973(.A1(new_n11803_), .A2(new_n6757_), .B1(new_n1078_), .B2(new_n10881_), .ZN(new_n12058_));
  AOI21_X1   g11974(.A1(new_n12058_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n12059_));
  XNOR2_X1   g11975(.A1(new_n11802_), .A2(new_n12059_), .ZN(new_n12060_));
  XOR2_X1    g11976(.A1(new_n11830_), .A2(new_n12060_), .Z(new_n12061_));
  XOR2_X1    g11977(.A1(new_n11830_), .A2(new_n12060_), .Z(new_n12062_));
  NOR2_X1    g11978(.A1(new_n12062_), .A2(new_n12057_), .ZN(new_n12063_));
  AOI21_X1   g11979(.A1(new_n12057_), .A2(new_n12061_), .B(new_n12063_), .ZN(new_n12064_));
  NAND2_X1   g11980(.A1(new_n12056_), .A2(new_n12064_), .ZN(new_n12065_));
  NOR2_X1    g11981(.A1(new_n12065_), .A2(new_n11838_), .ZN(new_n12066_));
  XOR2_X1    g11982(.A1(new_n12057_), .A2(new_n11830_), .Z(new_n12067_));
  NAND2_X1   g11983(.A1(new_n12067_), .A2(new_n12060_), .ZN(new_n12068_));
  XOR2_X1    g11984(.A1(new_n10619_), .A2(new_n10881_), .Z(new_n12069_));
  NAND2_X1   g11985(.A1(new_n12069_), .A2(new_n11799_), .ZN(new_n12070_));
  NOR2_X1    g11986(.A1(new_n12070_), .A2(new_n10874_), .ZN(new_n12071_));
  NAND2_X1   g11987(.A1(new_n12070_), .A2(new_n10874_), .ZN(new_n12072_));
  INV_X1     g11988(.I(new_n12072_), .ZN(new_n12073_));
  NOR2_X1    g11989(.A1(new_n12073_), .A2(new_n12071_), .ZN(new_n12074_));
  OAI22_X1   g11990(.A1(new_n10619_), .A2(new_n1078_), .B1(new_n6757_), .B2(new_n10885_), .ZN(new_n12075_));
  AOI21_X1   g11991(.A1(new_n12075_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n12076_));
  XOR2_X1    g11992(.A1(new_n12074_), .A2(new_n12076_), .Z(new_n12077_));
  NOR2_X1    g11993(.A1(new_n12068_), .A2(new_n12077_), .ZN(new_n12078_));
  INV_X1     g11994(.I(new_n12078_), .ZN(new_n12079_));
  AOI21_X1   g11995(.A1(new_n12065_), .A2(new_n11838_), .B(new_n12079_), .ZN(new_n12080_));
  NOR2_X1    g11996(.A1(new_n12080_), .A2(new_n12066_), .ZN(new_n12081_));
  OAI21_X1   g11997(.A1(new_n11729_), .A2(new_n11731_), .B(new_n11655_), .ZN(new_n12082_));
  NAND2_X1   g11998(.A1(new_n11656_), .A2(new_n11732_), .ZN(new_n12083_));
  NAND2_X1   g11999(.A1(new_n12083_), .A2(new_n12082_), .ZN(new_n12084_));
  NAND2_X1   g12000(.A1(new_n10886_), .A2(new_n10619_), .ZN(new_n12085_));
  OR2_X2     g12001(.A1(new_n10886_), .A2(new_n10619_), .Z(new_n12086_));
  AOI21_X1   g12002(.A1(new_n12086_), .A2(new_n12085_), .B(new_n10611_), .ZN(new_n12087_));
  INV_X1     g12003(.I(new_n10887_), .ZN(new_n12088_));
  AOI21_X1   g12004(.A1(new_n12088_), .A2(new_n10888_), .B(new_n10612_), .ZN(new_n12089_));
  NOR2_X1    g12005(.A1(new_n12089_), .A2(new_n12087_), .ZN(new_n12090_));
  NOR2_X1    g12006(.A1(new_n10619_), .A2(new_n10881_), .ZN(new_n12091_));
  OAI22_X1   g12007(.A1(new_n12091_), .A2(new_n6757_), .B1(new_n1078_), .B2(new_n10611_), .ZN(new_n12092_));
  AOI21_X1   g12008(.A1(new_n12092_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n12093_));
  XOR2_X1    g12009(.A1(new_n12090_), .A2(new_n12093_), .Z(new_n12094_));
  NOR2_X1    g12010(.A1(new_n12084_), .A2(new_n12094_), .ZN(new_n12095_));
  INV_X1     g12011(.I(new_n12094_), .ZN(new_n12096_));
  AOI21_X1   g12012(.A1(new_n12083_), .A2(new_n12082_), .B(new_n12096_), .ZN(new_n12097_));
  INV_X1     g12013(.I(new_n10989_), .ZN(new_n12098_));
  NOR2_X1    g12014(.A1(new_n11817_), .A2(new_n12098_), .ZN(new_n12099_));
  INV_X1     g12015(.I(new_n11816_), .ZN(new_n12100_));
  NOR2_X1    g12016(.A1(new_n12100_), .A2(new_n11814_), .ZN(new_n12101_));
  NOR2_X1    g12017(.A1(new_n12101_), .A2(new_n10989_), .ZN(new_n12102_));
  NOR2_X1    g12018(.A1(new_n12095_), .A2(new_n12097_), .ZN(new_n12104_));
  NOR2_X1    g12019(.A1(new_n12081_), .A2(new_n12104_), .ZN(new_n12105_));
  NAND2_X1   g12020(.A1(new_n11797_), .A2(new_n11806_), .ZN(new_n12106_));
  OAI22_X1   g12021(.A1(new_n11654_), .A2(new_n11641_), .B1(new_n11729_), .B2(new_n11731_), .ZN(new_n12108_));
  NAND2_X1   g12022(.A1(new_n11788_), .A2(new_n11786_), .ZN(new_n12109_));
  NAND2_X1   g12023(.A1(new_n12109_), .A2(new_n11791_), .ZN(new_n12110_));
  NOR2_X1    g12024(.A1(new_n11784_), .A2(new_n11777_), .ZN(new_n12111_));
  NAND2_X1   g12025(.A1(new_n11784_), .A2(new_n11777_), .ZN(new_n12112_));
  NOR2_X1    g12026(.A1(new_n11735_), .A2(new_n11780_), .ZN(new_n12113_));
  AOI21_X1   g12027(.A1(new_n12112_), .A2(new_n12113_), .B(new_n12111_), .ZN(new_n12114_));
  NAND2_X1   g12028(.A1(new_n11768_), .A2(new_n11772_), .ZN(new_n12115_));
  NAND2_X1   g12029(.A1(new_n11766_), .A2(new_n11744_), .ZN(new_n12116_));
  NAND2_X1   g12030(.A1(new_n12116_), .A2(new_n11765_), .ZN(new_n12117_));
  AOI21_X1   g12031(.A1(new_n11749_), .A2(new_n11757_), .B(new_n11755_), .ZN(new_n12118_));
  OAI22_X1   g12032(.A1(new_n4527_), .A2(new_n10777_), .B1(new_n10762_), .B2(new_n4529_), .ZN(new_n12119_));
  OAI21_X1   g12033(.A1(new_n10725_), .A2(new_n79_), .B(new_n12119_), .ZN(new_n12120_));
  AOI21_X1   g12034(.A1(new_n12120_), .A2(new_n72_), .B(new_n79_), .ZN(new_n12121_));
  XNOR2_X1   g12035(.A1(new_n11046_), .A2(new_n12121_), .ZN(new_n12122_));
  NAND2_X1   g12036(.A1(new_n10780_), .A2(new_n962_), .ZN(new_n12123_));
  NAND2_X1   g12037(.A1(new_n10783_), .A2(new_n4406_), .ZN(new_n12124_));
  AOI22_X1   g12038(.A1(new_n11030_), .A2(new_n961_), .B1(new_n12123_), .B2(new_n12124_), .ZN(new_n12125_));
  NAND2_X1   g12039(.A1(new_n12122_), .A2(new_n12125_), .ZN(new_n12126_));
  NOR2_X1    g12040(.A1(new_n12122_), .A2(new_n12125_), .ZN(new_n12127_));
  INV_X1     g12041(.I(new_n12127_), .ZN(new_n12128_));
  AOI21_X1   g12042(.A1(new_n12128_), .A2(new_n12126_), .B(new_n12118_), .ZN(new_n12129_));
  INV_X1     g12043(.I(new_n12118_), .ZN(new_n12130_));
  XNOR2_X1   g12044(.A1(new_n12122_), .A2(new_n12125_), .ZN(new_n12131_));
  NOR2_X1    g12045(.A1(new_n12131_), .A2(new_n12130_), .ZN(new_n12132_));
  NOR2_X1    g12046(.A1(new_n12132_), .A2(new_n12129_), .ZN(new_n12133_));
  OAI22_X1   g12047(.A1(new_n10792_), .A2(new_n4781_), .B1(new_n10696_), .B2(new_n4612_), .ZN(new_n12134_));
  OAI21_X1   g12048(.A1(new_n10672_), .A2(new_n1128_), .B(new_n12134_), .ZN(new_n12135_));
  AOI21_X1   g12049(.A1(new_n12135_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n12136_));
  XNOR2_X1   g12050(.A1(new_n11158_), .A2(new_n12136_), .ZN(new_n12137_));
  NAND2_X1   g12051(.A1(new_n12133_), .A2(new_n12137_), .ZN(new_n12138_));
  INV_X1     g12052(.I(new_n12137_), .ZN(new_n12139_));
  OAI21_X1   g12053(.A1(new_n12129_), .A2(new_n12132_), .B(new_n12139_), .ZN(new_n12140_));
  NAND2_X1   g12054(.A1(new_n12138_), .A2(new_n12140_), .ZN(new_n12141_));
  XOR2_X1    g12055(.A1(new_n12133_), .A2(new_n12139_), .Z(new_n12142_));
  NOR2_X1    g12056(.A1(new_n12142_), .A2(new_n12117_), .ZN(new_n12143_));
  AOI21_X1   g12057(.A1(new_n12117_), .A2(new_n12141_), .B(new_n12143_), .ZN(new_n12144_));
  NAND2_X1   g12058(.A1(new_n10652_), .A2(new_n10805_), .ZN(new_n12145_));
  AOI22_X1   g12059(.A1(new_n10828_), .A2(new_n247_), .B1(new_n5783_), .B2(new_n12145_), .ZN(new_n12146_));
  OAI21_X1   g12060(.A1(new_n12146_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n12147_));
  XOR2_X1    g12061(.A1(new_n11246_), .A2(new_n12147_), .Z(new_n12148_));
  AND2_X2    g12062(.A1(new_n12144_), .A2(new_n12148_), .Z(new_n12149_));
  NOR2_X1    g12063(.A1(new_n12144_), .A2(new_n12148_), .ZN(new_n12150_));
  NOR2_X1    g12064(.A1(new_n12149_), .A2(new_n12150_), .ZN(new_n12151_));
  NOR2_X1    g12065(.A1(new_n12151_), .A2(new_n11775_), .ZN(new_n12152_));
  XOR2_X1    g12066(.A1(new_n12152_), .A2(new_n12115_), .Z(new_n12153_));
  NOR2_X1    g12067(.A1(new_n12153_), .A2(new_n11743_), .ZN(new_n12154_));
  INV_X1     g12068(.I(new_n12154_), .ZN(new_n12155_));
  NAND2_X1   g12069(.A1(new_n12153_), .A2(new_n11743_), .ZN(new_n12156_));
  AOI22_X1   g12070(.A1(new_n10630_), .A2(new_n4717_), .B1(new_n5337_), .B2(new_n11446_), .ZN(new_n12157_));
  NOR2_X1    g12071(.A1(new_n12157_), .A2(\a[20] ), .ZN(new_n12158_));
  NOR2_X1    g12072(.A1(new_n12158_), .A2(new_n5398_), .ZN(new_n12159_));
  XOR2_X1    g12073(.A1(new_n11445_), .A2(new_n12159_), .Z(new_n12160_));
  INV_X1     g12074(.I(new_n12160_), .ZN(new_n12161_));
  AOI21_X1   g12075(.A1(new_n12155_), .A2(new_n12156_), .B(new_n12161_), .ZN(new_n12162_));
  INV_X1     g12076(.I(new_n12156_), .ZN(new_n12163_));
  NOR3_X1    g12077(.A1(new_n12163_), .A2(new_n12154_), .A3(new_n12160_), .ZN(new_n12164_));
  NOR2_X1    g12078(.A1(new_n12162_), .A2(new_n12164_), .ZN(new_n12165_));
  NOR2_X1    g12079(.A1(new_n12114_), .A2(new_n12165_), .ZN(new_n12166_));
  INV_X1     g12080(.I(new_n12111_), .ZN(new_n12167_));
  NAND2_X1   g12081(.A1(new_n12112_), .A2(new_n12113_), .ZN(new_n12168_));
  NAND2_X1   g12082(.A1(new_n12168_), .A2(new_n12167_), .ZN(new_n12169_));
  NOR3_X1    g12083(.A1(new_n12163_), .A2(new_n12154_), .A3(new_n12161_), .ZN(new_n12170_));
  AOI21_X1   g12084(.A1(new_n12155_), .A2(new_n12156_), .B(new_n12160_), .ZN(new_n12171_));
  NOR2_X1    g12085(.A1(new_n12171_), .A2(new_n12170_), .ZN(new_n12172_));
  NOR2_X1    g12086(.A1(new_n12169_), .A2(new_n12172_), .ZN(new_n12173_));
  OAI22_X1   g12087(.A1(new_n10870_), .A2(new_n1620_), .B1(new_n5420_), .B2(new_n10861_), .ZN(new_n12174_));
  AOI21_X1   g12088(.A1(new_n12174_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n12175_));
  XOR2_X1    g12089(.A1(new_n11648_), .A2(new_n12175_), .Z(new_n12176_));
  INV_X1     g12090(.I(new_n12176_), .ZN(new_n12177_));
  OAI21_X1   g12091(.A1(new_n12173_), .A2(new_n12166_), .B(new_n12177_), .ZN(new_n12178_));
  AOI21_X1   g12092(.A1(new_n11796_), .A2(new_n11734_), .B(new_n12178_), .ZN(new_n12179_));
  NAND3_X1   g12093(.A1(new_n11796_), .A2(new_n12178_), .A3(new_n11734_), .ZN(new_n12180_));
  INV_X1     g12094(.I(new_n12180_), .ZN(new_n12181_));
  OAI21_X1   g12095(.A1(new_n12181_), .A2(new_n12179_), .B(new_n12110_), .ZN(new_n12182_));
  INV_X1     g12096(.I(new_n12110_), .ZN(new_n12183_));
  INV_X1     g12097(.I(new_n12179_), .ZN(new_n12184_));
  NAND3_X1   g12098(.A1(new_n12184_), .A2(new_n12180_), .A3(new_n12183_), .ZN(new_n12185_));
  NAND2_X1   g12099(.A1(new_n12185_), .A2(new_n12182_), .ZN(new_n12186_));
  OAI22_X1   g12100(.A1(new_n10619_), .A2(new_n643_), .B1(new_n5967_), .B2(new_n10885_), .ZN(new_n12187_));
  AOI21_X1   g12101(.A1(new_n12187_), .A2(new_n279_), .B(new_n643_), .ZN(new_n12188_));
  XOR2_X1    g12102(.A1(new_n12074_), .A2(new_n12188_), .Z(new_n12189_));
  INV_X1     g12103(.I(new_n12189_), .ZN(new_n12190_));
  NAND3_X1   g12104(.A1(new_n12186_), .A2(new_n12108_), .A3(new_n12190_), .ZN(new_n12191_));
  INV_X1     g12105(.I(new_n11459_), .ZN(new_n12192_));
  NAND2_X1   g12106(.A1(new_n11831_), .A2(new_n12192_), .ZN(new_n12193_));
  OAI21_X1   g12107(.A1(new_n11831_), .A2(new_n12192_), .B(new_n11652_), .ZN(new_n12194_));
  INV_X1     g12108(.I(new_n11729_), .ZN(new_n12195_));
  AOI22_X1   g12109(.A1(new_n12194_), .A2(new_n12193_), .B1(new_n12195_), .B2(new_n11730_), .ZN(new_n12196_));
  AOI21_X1   g12110(.A1(new_n12184_), .A2(new_n12180_), .B(new_n12183_), .ZN(new_n12197_));
  NOR3_X1    g12111(.A1(new_n12181_), .A2(new_n12179_), .A3(new_n12110_), .ZN(new_n12198_));
  NOR2_X1    g12112(.A1(new_n12197_), .A2(new_n12198_), .ZN(new_n12199_));
  OAI21_X1   g12113(.A1(new_n12199_), .A2(new_n12189_), .B(new_n12196_), .ZN(new_n12200_));
  NAND2_X1   g12114(.A1(new_n12200_), .A2(new_n12191_), .ZN(new_n12201_));
  NAND2_X1   g12115(.A1(new_n12201_), .A2(new_n12106_), .ZN(new_n12202_));
  NAND3_X1   g12116(.A1(new_n12200_), .A2(new_n12191_), .A3(new_n11812_), .ZN(new_n12203_));
  INV_X1     g12117(.I(new_n10606_), .ZN(new_n12204_));
  NAND2_X1   g12118(.A1(new_n12204_), .A2(new_n10896_), .ZN(new_n12205_));
  NAND2_X1   g12119(.A1(new_n10606_), .A2(new_n10897_), .ZN(new_n12206_));
  AOI21_X1   g12120(.A1(new_n12205_), .A2(new_n12206_), .B(new_n10982_), .ZN(new_n12207_));
  NAND2_X1   g12121(.A1(new_n10889_), .A2(new_n12207_), .ZN(new_n12208_));
  INV_X1     g12122(.I(new_n12208_), .ZN(new_n12209_));
  NOR2_X1    g12123(.A1(new_n10889_), .A2(new_n12207_), .ZN(new_n12210_));
  NOR2_X1    g12124(.A1(new_n12209_), .A2(new_n12210_), .ZN(new_n12211_));
  OAI22_X1   g12125(.A1(new_n10606_), .A2(new_n1078_), .B1(new_n6757_), .B2(new_n10901_), .ZN(new_n12212_));
  AOI21_X1   g12126(.A1(new_n12212_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n12213_));
  XOR2_X1    g12127(.A1(new_n12211_), .A2(new_n12213_), .Z(new_n12214_));
  AOI21_X1   g12128(.A1(new_n12202_), .A2(new_n12203_), .B(new_n12214_), .ZN(new_n12215_));
  INV_X1     g12129(.I(new_n12215_), .ZN(new_n12216_));
  NOR2_X1    g12130(.A1(new_n12105_), .A2(new_n12216_), .ZN(new_n12217_));
  NAND2_X1   g12131(.A1(new_n12061_), .A2(new_n12057_), .ZN(new_n12218_));
  OAI21_X1   g12132(.A1(new_n12057_), .A2(new_n12062_), .B(new_n12218_), .ZN(new_n12219_));
  NOR3_X1    g12133(.A1(new_n12219_), .A2(new_n12054_), .A3(new_n12055_), .ZN(new_n12220_));
  NAND2_X1   g12134(.A1(new_n12220_), .A2(new_n11837_), .ZN(new_n12221_));
  OAI21_X1   g12135(.A1(new_n12220_), .A2(new_n11837_), .B(new_n12078_), .ZN(new_n12222_));
  NAND2_X1   g12136(.A1(new_n12222_), .A2(new_n12221_), .ZN(new_n12223_));
  OAI21_X1   g12137(.A1(new_n12095_), .A2(new_n12097_), .B(new_n12223_), .ZN(new_n12224_));
  NOR2_X1    g12138(.A1(new_n12224_), .A2(new_n12215_), .ZN(new_n12225_));
  OAI21_X1   g12139(.A1(new_n12217_), .A2(new_n12225_), .B(new_n11818_), .ZN(new_n12226_));
  NOR2_X1    g12140(.A1(new_n12101_), .A2(new_n12098_), .ZN(new_n12227_));
  NAND2_X1   g12141(.A1(new_n12224_), .A2(new_n12215_), .ZN(new_n12228_));
  NAND2_X1   g12142(.A1(new_n12105_), .A2(new_n12216_), .ZN(new_n12229_));
  NAND3_X1   g12143(.A1(new_n12229_), .A2(new_n12228_), .A3(new_n12227_), .ZN(new_n12230_));
  NAND2_X1   g12144(.A1(new_n12226_), .A2(new_n12230_), .ZN(new_n12231_));
  AOI21_X1   g12145(.A1(new_n11834_), .A2(new_n11836_), .B(new_n12077_), .ZN(new_n12232_));
  INV_X1     g12146(.I(new_n12232_), .ZN(new_n12233_));
  NOR2_X1    g12147(.A1(new_n12233_), .A2(new_n12220_), .ZN(new_n12234_));
  NOR2_X1    g12148(.A1(new_n12065_), .A2(new_n12232_), .ZN(new_n12235_));
  OAI21_X1   g12149(.A1(new_n12235_), .A2(new_n12234_), .B(new_n12068_), .ZN(new_n12236_));
  INV_X1     g12150(.I(new_n12068_), .ZN(new_n12237_));
  NAND2_X1   g12151(.A1(new_n12065_), .A2(new_n12232_), .ZN(new_n12238_));
  NAND2_X1   g12152(.A1(new_n12233_), .A2(new_n12220_), .ZN(new_n12239_));
  NAND3_X1   g12153(.A1(new_n12238_), .A2(new_n12239_), .A3(new_n12237_), .ZN(new_n12240_));
  NAND2_X1   g12154(.A1(new_n12236_), .A2(new_n12240_), .ZN(new_n12241_));
  AOI21_X1   g12155(.A1(new_n12028_), .A2(new_n12029_), .B(new_n12033_), .ZN(new_n12242_));
  INV_X1     g12156(.I(new_n12034_), .ZN(new_n12243_));
  NOR2_X1    g12157(.A1(new_n12243_), .A2(new_n12242_), .ZN(new_n12244_));
  NAND3_X1   g12158(.A1(new_n12244_), .A2(new_n12019_), .A3(new_n12021_), .ZN(new_n12245_));
  INV_X1     g12159(.I(new_n12042_), .ZN(new_n12246_));
  NAND3_X1   g12160(.A1(new_n11850_), .A2(new_n12245_), .A3(new_n12246_), .ZN(new_n12247_));
  AOI21_X1   g12161(.A1(new_n11847_), .A2(new_n11848_), .B(new_n11846_), .ZN(new_n12248_));
  NOR3_X1    g12162(.A1(new_n11844_), .A2(new_n11841_), .A3(new_n11591_), .ZN(new_n12249_));
  NOR2_X1    g12163(.A1(new_n12249_), .A2(new_n12248_), .ZN(new_n12250_));
  OAI21_X1   g12164(.A1(new_n12250_), .A2(new_n12042_), .B(new_n12038_), .ZN(new_n12251_));
  AOI21_X1   g12165(.A1(new_n12251_), .A2(new_n12247_), .B(new_n12242_), .ZN(new_n12252_));
  NOR3_X1    g12166(.A1(new_n12250_), .A2(new_n12038_), .A3(new_n12042_), .ZN(new_n12253_));
  AOI21_X1   g12167(.A1(new_n11850_), .A2(new_n12246_), .B(new_n12245_), .ZN(new_n12254_));
  NOR3_X1    g12168(.A1(new_n12253_), .A2(new_n12254_), .A3(new_n12036_), .ZN(new_n12255_));
  NOR2_X1    g12169(.A1(new_n12255_), .A2(new_n12252_), .ZN(new_n12256_));
  NAND3_X1   g12170(.A1(new_n11993_), .A2(new_n11983_), .A3(new_n11999_), .ZN(new_n12257_));
  AOI21_X1   g12171(.A1(new_n11879_), .A2(new_n11868_), .B(new_n11980_), .ZN(new_n12258_));
  NAND2_X1   g12172(.A1(new_n12258_), .A2(new_n11880_), .ZN(new_n12259_));
  NOR2_X1    g12173(.A1(new_n12259_), .A2(new_n11857_), .ZN(new_n12260_));
  AOI21_X1   g12174(.A1(new_n12259_), .A2(new_n11857_), .B(new_n11991_), .ZN(new_n12261_));
  OAI21_X1   g12175(.A1(new_n12261_), .A2(new_n12260_), .B(new_n11998_), .ZN(new_n12262_));
  AOI21_X1   g12176(.A1(new_n12257_), .A2(new_n12262_), .B(new_n11569_), .ZN(new_n12263_));
  NOR3_X1    g12177(.A1(new_n12261_), .A2(new_n12260_), .A3(new_n11998_), .ZN(new_n12264_));
  INV_X1     g12178(.I(new_n12262_), .ZN(new_n12265_));
  NOR3_X1    g12179(.A1(new_n12265_), .A2(new_n11570_), .A3(new_n12264_), .ZN(new_n12266_));
  OAI21_X1   g12180(.A1(new_n12266_), .A2(new_n12263_), .B(new_n12004_), .ZN(new_n12267_));
  OAI21_X1   g12181(.A1(new_n12265_), .A2(new_n12264_), .B(new_n11570_), .ZN(new_n12268_));
  NAND3_X1   g12182(.A1(new_n12257_), .A2(new_n11569_), .A3(new_n12262_), .ZN(new_n12269_));
  NAND3_X1   g12183(.A1(new_n12268_), .A2(new_n12269_), .A3(new_n12005_), .ZN(new_n12270_));
  NAND2_X1   g12184(.A1(new_n12267_), .A2(new_n12270_), .ZN(new_n12271_));
  INV_X1     g12185(.I(new_n11954_), .ZN(new_n12272_));
  NOR3_X1    g12186(.A1(new_n11968_), .A2(new_n11969_), .A3(new_n11965_), .ZN(new_n12273_));
  NOR3_X1    g12187(.A1(new_n12273_), .A2(new_n11973_), .A3(new_n12272_), .ZN(new_n12274_));
  NOR2_X1    g12188(.A1(new_n11887_), .A2(new_n11976_), .ZN(new_n12275_));
  INV_X1     g12189(.I(new_n12275_), .ZN(new_n12276_));
  NOR2_X1    g12190(.A1(new_n12274_), .A2(new_n12276_), .ZN(new_n12277_));
  NOR2_X1    g12191(.A1(new_n11971_), .A2(new_n12275_), .ZN(new_n12278_));
  OAI21_X1   g12192(.A1(new_n12277_), .A2(new_n12278_), .B(new_n11970_), .ZN(new_n12279_));
  NAND2_X1   g12193(.A1(new_n11971_), .A2(new_n12275_), .ZN(new_n12280_));
  NAND2_X1   g12194(.A1(new_n12274_), .A2(new_n12276_), .ZN(new_n12281_));
  NAND3_X1   g12195(.A1(new_n12281_), .A2(new_n12280_), .A3(new_n11973_), .ZN(new_n12282_));
  NAND2_X1   g12196(.A1(new_n12279_), .A2(new_n12282_), .ZN(new_n12283_));
  INV_X1     g12197(.I(new_n11923_), .ZN(new_n12284_));
  NAND2_X1   g12198(.A1(new_n11920_), .A2(new_n11498_), .ZN(new_n12285_));
  INV_X1     g12199(.I(new_n11498_), .ZN(new_n12286_));
  NAND2_X1   g12200(.A1(new_n11917_), .A2(new_n11919_), .ZN(new_n12287_));
  NAND2_X1   g12201(.A1(new_n12287_), .A2(new_n12286_), .ZN(new_n12288_));
  AOI21_X1   g12202(.A1(new_n12285_), .A2(new_n12288_), .B(new_n12284_), .ZN(new_n12289_));
  NAND3_X1   g12203(.A1(new_n12285_), .A2(new_n12284_), .A3(new_n12288_), .ZN(new_n12290_));
  INV_X1     g12204(.I(new_n12290_), .ZN(new_n12291_));
  OAI21_X1   g12205(.A1(new_n12291_), .A2(new_n12289_), .B(new_n11505_), .ZN(new_n12292_));
  INV_X1     g12206(.I(new_n11505_), .ZN(new_n12293_));
  NAND2_X1   g12207(.A1(new_n12285_), .A2(new_n12288_), .ZN(new_n12294_));
  NAND2_X1   g12208(.A1(new_n12294_), .A2(new_n11923_), .ZN(new_n12295_));
  NAND3_X1   g12209(.A1(new_n12295_), .A2(new_n12290_), .A3(new_n12293_), .ZN(new_n12296_));
  NAND2_X1   g12210(.A1(new_n12292_), .A2(new_n12296_), .ZN(new_n12297_));
  XOR2_X1    g12211(.A1(new_n11890_), .A2(new_n11503_), .Z(new_n12298_));
  NAND3_X1   g12212(.A1(new_n12298_), .A2(new_n11898_), .A3(new_n11906_), .ZN(new_n12299_));
  NAND2_X1   g12213(.A1(new_n11892_), .A2(new_n11908_), .ZN(new_n12300_));
  NAND2_X1   g12214(.A1(new_n12300_), .A2(new_n11907_), .ZN(new_n12301_));
  NAND2_X1   g12215(.A1(new_n12301_), .A2(new_n12299_), .ZN(new_n12302_));
  AOI22_X1   g12216(.A1(new_n11141_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n10691_), .ZN(new_n12303_));
  OAI21_X1   g12217(.A1(new_n12303_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n12304_));
  INV_X1     g12218(.I(new_n12304_), .ZN(new_n12305_));
  NAND2_X1   g12219(.A1(new_n11140_), .A2(new_n12305_), .ZN(new_n12306_));
  NAND2_X1   g12220(.A1(new_n11333_), .A2(new_n12304_), .ZN(new_n12307_));
  NAND2_X1   g12221(.A1(new_n12306_), .A2(new_n12307_), .ZN(new_n12308_));
  NAND2_X1   g12222(.A1(new_n11915_), .A2(new_n11911_), .ZN(new_n12309_));
  NAND2_X1   g12223(.A1(new_n11918_), .A2(new_n11912_), .ZN(new_n12310_));
  AOI22_X1   g12224(.A1(new_n12309_), .A2(new_n12310_), .B1(new_n11892_), .B2(new_n11909_), .ZN(new_n12311_));
  AOI21_X1   g12225(.A1(new_n11916_), .A2(new_n11919_), .B(new_n11910_), .ZN(new_n12312_));
  NOR2_X1    g12226(.A1(new_n12311_), .A2(new_n12312_), .ZN(new_n12313_));
  INV_X1     g12227(.I(new_n11159_), .ZN(new_n12314_));
  AOI22_X1   g12228(.A1(new_n10817_), .A2(new_n2469_), .B1(new_n12314_), .B2(new_n7838_), .ZN(new_n12315_));
  OAI21_X1   g12229(.A1(new_n12315_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n12316_));
  XOR2_X1    g12230(.A1(new_n11158_), .A2(new_n12316_), .Z(new_n12317_));
  INV_X1     g12231(.I(new_n12317_), .ZN(new_n12318_));
  NAND2_X1   g12232(.A1(new_n12318_), .A2(new_n12313_), .ZN(new_n12319_));
  OAI21_X1   g12233(.A1(new_n12311_), .A2(new_n12312_), .B(new_n12317_), .ZN(new_n12320_));
  NAND2_X1   g12234(.A1(new_n12319_), .A2(new_n12320_), .ZN(new_n12321_));
  AOI21_X1   g12235(.A1(new_n12321_), .A2(new_n12308_), .B(new_n12302_), .ZN(new_n12322_));
  OAI22_X1   g12236(.A1(new_n10725_), .A2(new_n2495_), .B1(new_n7837_), .B2(new_n11047_), .ZN(new_n12323_));
  AOI21_X1   g12237(.A1(new_n12323_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12324_));
  XOR2_X1    g12238(.A1(new_n11046_), .A2(new_n12324_), .Z(new_n12325_));
  NOR3_X1    g12239(.A1(new_n11901_), .A2(new_n11902_), .A3(new_n11904_), .ZN(new_n12326_));
  NOR2_X1    g12240(.A1(new_n11901_), .A2(new_n11902_), .ZN(new_n12327_));
  NOR2_X1    g12241(.A1(new_n12327_), .A2(new_n11905_), .ZN(new_n12328_));
  NOR2_X1    g12242(.A1(new_n12328_), .A2(new_n12326_), .ZN(new_n12329_));
  INV_X1     g12243(.I(new_n12329_), .ZN(new_n12330_));
  INV_X1     g12244(.I(new_n11903_), .ZN(new_n12331_));
  NOR2_X1    g12245(.A1(new_n11009_), .A2(new_n2469_), .ZN(new_n12332_));
  NAND2_X1   g12246(.A1(new_n11009_), .A2(new_n2469_), .ZN(new_n12333_));
  NAND2_X1   g12247(.A1(new_n12333_), .A2(new_n10762_), .ZN(new_n12334_));
  NOR2_X1    g12248(.A1(new_n12334_), .A2(new_n12332_), .ZN(new_n12335_));
  NAND2_X1   g12249(.A1(new_n10780_), .A2(new_n5108_), .ZN(new_n12336_));
  NAND2_X1   g12250(.A1(new_n10783_), .A2(new_n5110_), .ZN(new_n12337_));
  AOI22_X1   g12251(.A1(new_n12337_), .A2(new_n12336_), .B1(new_n11002_), .B2(new_n2469_), .ZN(new_n12338_));
  INV_X1     g12252(.I(new_n12338_), .ZN(new_n12339_));
  OAI21_X1   g12253(.A1(new_n12335_), .A2(new_n12339_), .B(new_n498_), .ZN(new_n12340_));
  NOR3_X1    g12254(.A1(new_n12335_), .A2(new_n498_), .A3(new_n12339_), .ZN(new_n12341_));
  INV_X1     g12255(.I(new_n12341_), .ZN(new_n12342_));
  NAND2_X1   g12256(.A1(new_n12342_), .A2(new_n12340_), .ZN(new_n12343_));
  NAND2_X1   g12257(.A1(new_n10783_), .A2(new_n5108_), .ZN(new_n12344_));
  AOI21_X1   g12258(.A1(new_n10780_), .A2(new_n2469_), .B(\a[8] ), .ZN(new_n12345_));
  AOI21_X1   g12259(.A1(new_n12344_), .A2(new_n12345_), .B(new_n2495_), .ZN(new_n12346_));
  NAND2_X1   g12260(.A1(new_n11030_), .A2(new_n12346_), .ZN(new_n12347_));
  NOR2_X1    g12261(.A1(new_n11030_), .A2(new_n12346_), .ZN(new_n12348_));
  INV_X1     g12262(.I(new_n12348_), .ZN(new_n12349_));
  NAND2_X1   g12263(.A1(new_n12349_), .A2(new_n12347_), .ZN(new_n12350_));
  NOR2_X1    g12264(.A1(new_n10780_), .A2(new_n2583_), .ZN(new_n12351_));
  NOR2_X1    g12265(.A1(new_n12351_), .A2(new_n498_), .ZN(new_n12352_));
  INV_X1     g12266(.I(new_n12352_), .ZN(new_n12353_));
  NOR2_X1    g12267(.A1(new_n12350_), .A2(new_n12353_), .ZN(new_n12354_));
  INV_X1     g12268(.I(new_n12354_), .ZN(new_n12355_));
  NOR3_X1    g12269(.A1(new_n12355_), .A2(new_n12343_), .A3(new_n12331_), .ZN(new_n12356_));
  INV_X1     g12270(.I(new_n12340_), .ZN(new_n12357_));
  NOR2_X1    g12271(.A1(new_n12357_), .A2(new_n12341_), .ZN(new_n12358_));
  AOI21_X1   g12272(.A1(new_n12358_), .A2(new_n12354_), .B(new_n11903_), .ZN(new_n12359_));
  AOI22_X1   g12273(.A1(new_n11003_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n10745_), .ZN(new_n12360_));
  NOR2_X1    g12274(.A1(new_n12360_), .A2(\a[8] ), .ZN(new_n12361_));
  NOR2_X1    g12275(.A1(new_n12361_), .A2(new_n2495_), .ZN(new_n12362_));
  XOR2_X1    g12276(.A1(new_n12362_), .A2(new_n11188_), .Z(new_n12363_));
  NAND2_X1   g12277(.A1(new_n12325_), .A2(new_n12330_), .ZN(new_n12364_));
  AOI22_X1   g12278(.A1(new_n10794_), .A2(new_n2469_), .B1(new_n7838_), .B2(new_n11065_), .ZN(new_n12365_));
  OAI21_X1   g12279(.A1(new_n12365_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n12366_));
  XOR2_X1    g12280(.A1(new_n11064_), .A2(new_n12366_), .Z(new_n12367_));
  NOR2_X1    g12281(.A1(new_n12367_), .A2(new_n12364_), .ZN(new_n12368_));
  XOR2_X1    g12282(.A1(new_n11897_), .A2(new_n294_), .Z(new_n12369_));
  INV_X1     g12283(.I(new_n11906_), .ZN(new_n12370_));
  NAND2_X1   g12284(.A1(new_n12369_), .A2(new_n12370_), .ZN(new_n12371_));
  AOI22_X1   g12285(.A1(new_n12367_), .A2(new_n12364_), .B1(new_n11907_), .B2(new_n12371_), .ZN(new_n12372_));
  NOR2_X1    g12286(.A1(new_n12372_), .A2(new_n12368_), .ZN(new_n12373_));
  INV_X1     g12287(.I(new_n12373_), .ZN(new_n12374_));
  OAI21_X1   g12288(.A1(new_n12321_), .A2(new_n12308_), .B(new_n12374_), .ZN(new_n12375_));
  NOR2_X1    g12289(.A1(new_n12322_), .A2(new_n12375_), .ZN(new_n12376_));
  NAND2_X1   g12290(.A1(new_n12297_), .A2(new_n12376_), .ZN(new_n12377_));
  OAI22_X1   g12291(.A1(new_n11176_), .A2(new_n7837_), .B1(new_n10658_), .B2(new_n2495_), .ZN(new_n12378_));
  AOI21_X1   g12292(.A1(new_n12378_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12379_));
  XOR2_X1    g12293(.A1(new_n11175_), .A2(new_n12379_), .Z(new_n12380_));
  NOR2_X1    g12294(.A1(new_n12380_), .A2(new_n12320_), .ZN(new_n12381_));
  OAI21_X1   g12295(.A1(new_n12297_), .A2(new_n12376_), .B(new_n12381_), .ZN(new_n12382_));
  NOR2_X1    g12296(.A1(new_n11938_), .A2(new_n11933_), .ZN(new_n12383_));
  NOR2_X1    g12297(.A1(new_n11937_), .A2(new_n11934_), .ZN(new_n12384_));
  OAI22_X1   g12298(.A1(new_n11927_), .A2(new_n11924_), .B1(new_n12383_), .B2(new_n12384_), .ZN(new_n12385_));
  NOR2_X1    g12299(.A1(new_n11937_), .A2(new_n11933_), .ZN(new_n12386_));
  OAI21_X1   g12300(.A1(new_n11939_), .A2(new_n12386_), .B(new_n11928_), .ZN(new_n12387_));
  NAND2_X1   g12301(.A1(new_n12387_), .A2(new_n12385_), .ZN(new_n12388_));
  OAI22_X1   g12302(.A1(new_n10819_), .A2(new_n7837_), .B1(new_n11214_), .B2(new_n2495_), .ZN(new_n12389_));
  AOI21_X1   g12303(.A1(new_n12389_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12390_));
  XOR2_X1    g12304(.A1(new_n11224_), .A2(new_n12390_), .Z(new_n12391_));
  AOI22_X1   g12305(.A1(new_n12382_), .A2(new_n12377_), .B1(new_n12388_), .B2(new_n12391_), .ZN(new_n12392_));
  INV_X1     g12306(.I(new_n12391_), .ZN(new_n12393_));
  NAND3_X1   g12307(.A1(new_n12387_), .A2(new_n12385_), .A3(new_n12393_), .ZN(new_n12394_));
  INV_X1     g12308(.I(new_n12394_), .ZN(new_n12395_));
  XOR2_X1    g12309(.A1(new_n11951_), .A2(new_n11948_), .Z(new_n12396_));
  AND2_X2    g12310(.A1(new_n12396_), .A2(new_n11941_), .Z(new_n12397_));
  AOI21_X1   g12311(.A1(new_n11950_), .A2(new_n11952_), .B(new_n11941_), .ZN(new_n12398_));
  NOR2_X1    g12312(.A1(new_n12397_), .A2(new_n12398_), .ZN(new_n12399_));
  AOI21_X1   g12313(.A1(new_n10652_), .A2(new_n10805_), .B(new_n7837_), .ZN(new_n12400_));
  NOR2_X1    g12314(.A1(new_n10646_), .A2(new_n2495_), .ZN(new_n12401_));
  OAI21_X1   g12315(.A1(new_n12401_), .A2(new_n12400_), .B(new_n498_), .ZN(new_n12402_));
  NAND2_X1   g12316(.A1(new_n12402_), .A2(new_n2469_), .ZN(new_n12403_));
  XOR2_X1    g12317(.A1(new_n11246_), .A2(new_n12403_), .Z(new_n12404_));
  INV_X1     g12318(.I(new_n12404_), .ZN(new_n12405_));
  OAI22_X1   g12319(.A1(new_n12392_), .A2(new_n12395_), .B1(new_n12399_), .B2(new_n12405_), .ZN(new_n12406_));
  INV_X1     g12320(.I(new_n12406_), .ZN(new_n12407_));
  INV_X1     g12321(.I(new_n12399_), .ZN(new_n12408_));
  NOR2_X1    g12322(.A1(new_n12408_), .A2(new_n12404_), .ZN(new_n12409_));
  OAI21_X1   g12323(.A1(new_n12273_), .A2(new_n11973_), .B(new_n12272_), .ZN(new_n12410_));
  AOI22_X1   g12324(.A1(new_n10638_), .A2(new_n2469_), .B1(new_n7838_), .B2(new_n11269_), .ZN(new_n12411_));
  NOR2_X1    g12325(.A1(new_n12411_), .A2(\a[8] ), .ZN(new_n12412_));
  NOR2_X1    g12326(.A1(new_n12412_), .A2(new_n2495_), .ZN(new_n12413_));
  XNOR2_X1   g12327(.A1(new_n11268_), .A2(new_n12413_), .ZN(new_n12414_));
  NAND3_X1   g12328(.A1(new_n12410_), .A2(new_n11971_), .A3(new_n12414_), .ZN(new_n12415_));
  AOI21_X1   g12329(.A1(new_n11970_), .A2(new_n11967_), .B(new_n11954_), .ZN(new_n12416_));
  INV_X1     g12330(.I(new_n12414_), .ZN(new_n12417_));
  OAI21_X1   g12331(.A1(new_n12274_), .A2(new_n12416_), .B(new_n12417_), .ZN(new_n12418_));
  NAND2_X1   g12332(.A1(new_n12418_), .A2(new_n12415_), .ZN(new_n12419_));
  NOR3_X1    g12333(.A1(new_n12407_), .A2(new_n12419_), .A3(new_n12409_), .ZN(new_n12420_));
  NAND2_X1   g12334(.A1(new_n12420_), .A2(new_n12283_), .ZN(new_n12421_));
  NOR3_X1    g12335(.A1(new_n12417_), .A2(new_n12274_), .A3(new_n12416_), .ZN(new_n12422_));
  OAI22_X1   g12336(.A1(new_n11386_), .A2(new_n7837_), .B1(new_n2495_), .B2(new_n10633_), .ZN(new_n12423_));
  AOI21_X1   g12337(.A1(new_n12423_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12424_));
  XOR2_X1    g12338(.A1(new_n11987_), .A2(new_n12424_), .Z(new_n12425_));
  NAND2_X1   g12339(.A1(new_n12422_), .A2(new_n12425_), .ZN(new_n12426_));
  INV_X1     g12340(.I(new_n12426_), .ZN(new_n12427_));
  OAI21_X1   g12341(.A1(new_n12420_), .A2(new_n12283_), .B(new_n12427_), .ZN(new_n12428_));
  AOI22_X1   g12342(.A1(new_n10630_), .A2(new_n2469_), .B1(new_n7838_), .B2(new_n11446_), .ZN(new_n12429_));
  NOR2_X1    g12343(.A1(new_n12429_), .A2(\a[8] ), .ZN(new_n12430_));
  NOR2_X1    g12344(.A1(new_n12430_), .A2(new_n2495_), .ZN(new_n12431_));
  XOR2_X1    g12345(.A1(new_n11445_), .A2(new_n12431_), .Z(new_n12432_));
  AOI21_X1   g12346(.A1(new_n12428_), .A2(new_n12421_), .B(new_n12432_), .ZN(new_n12433_));
  AND2_X2    g12347(.A1(new_n12279_), .A2(new_n12282_), .Z(new_n12434_));
  INV_X1     g12348(.I(new_n12409_), .ZN(new_n12435_));
  AOI21_X1   g12349(.A1(new_n12410_), .A2(new_n11971_), .B(new_n12414_), .ZN(new_n12436_));
  NOR2_X1    g12350(.A1(new_n12422_), .A2(new_n12436_), .ZN(new_n12437_));
  NAND3_X1   g12351(.A1(new_n12437_), .A2(new_n12406_), .A3(new_n12435_), .ZN(new_n12438_));
  NOR2_X1    g12352(.A1(new_n12434_), .A2(new_n12438_), .ZN(new_n12439_));
  AOI21_X1   g12353(.A1(new_n12434_), .A2(new_n12438_), .B(new_n12426_), .ZN(new_n12440_));
  INV_X1     g12354(.I(new_n12432_), .ZN(new_n12441_));
  NOR3_X1    g12355(.A1(new_n12440_), .A2(new_n12439_), .A3(new_n12441_), .ZN(new_n12442_));
  NAND2_X1   g12356(.A1(new_n11868_), .A2(new_n11862_), .ZN(new_n12443_));
  NOR2_X1    g12357(.A1(new_n11868_), .A2(new_n11862_), .ZN(new_n12444_));
  INV_X1     g12358(.I(new_n12444_), .ZN(new_n12445_));
  NAND2_X1   g12359(.A1(new_n12445_), .A2(new_n12443_), .ZN(new_n12446_));
  XOR2_X1    g12360(.A1(new_n12446_), .A2(new_n11980_), .Z(new_n12447_));
  NOR2_X1    g12361(.A1(new_n12442_), .A2(new_n12447_), .ZN(new_n12448_));
  NOR2_X1    g12362(.A1(new_n12448_), .A2(new_n12433_), .ZN(new_n12449_));
  INV_X1     g12363(.I(new_n12449_), .ZN(new_n12450_));
  XOR2_X1    g12364(.A1(new_n11867_), .A2(new_n11862_), .Z(new_n12451_));
  NOR3_X1    g12365(.A1(new_n11879_), .A2(new_n12444_), .A3(new_n12451_), .ZN(new_n12452_));
  NOR2_X1    g12366(.A1(new_n11868_), .A2(new_n11862_), .ZN(new_n12453_));
  NOR2_X1    g12367(.A1(new_n12452_), .A2(new_n12453_), .ZN(new_n12454_));
  NOR2_X1    g12368(.A1(new_n12454_), .A2(new_n11981_), .ZN(new_n12455_));
  INV_X1     g12369(.I(new_n12455_), .ZN(new_n12456_));
  NAND2_X1   g12370(.A1(new_n12454_), .A2(new_n11981_), .ZN(new_n12457_));
  NAND2_X1   g12371(.A1(new_n12456_), .A2(new_n12457_), .ZN(new_n12458_));
  AOI22_X1   g12372(.A1(new_n2469_), .A2(new_n10843_), .B1(new_n11608_), .B2(new_n7838_), .ZN(new_n12459_));
  OAI21_X1   g12373(.A1(new_n12459_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n12460_));
  XOR2_X1    g12374(.A1(new_n11607_), .A2(new_n12460_), .Z(new_n12461_));
  NAND2_X1   g12375(.A1(new_n12458_), .A2(new_n12461_), .ZN(new_n12462_));
  NAND2_X1   g12376(.A1(new_n12462_), .A2(new_n12450_), .ZN(new_n12463_));
  INV_X1     g12377(.I(new_n12457_), .ZN(new_n12464_));
  NOR2_X1    g12378(.A1(new_n12464_), .A2(new_n12455_), .ZN(new_n12465_));
  INV_X1     g12379(.I(new_n12461_), .ZN(new_n12466_));
  NAND2_X1   g12380(.A1(new_n12465_), .A2(new_n12466_), .ZN(new_n12467_));
  INV_X1     g12381(.I(new_n11876_), .ZN(new_n12468_));
  OAI21_X1   g12382(.A1(new_n11856_), .A2(new_n11855_), .B(new_n11990_), .ZN(new_n12469_));
  AOI21_X1   g12383(.A1(new_n11880_), .A2(new_n12258_), .B(new_n12469_), .ZN(new_n12470_));
  INV_X1     g12384(.I(new_n12469_), .ZN(new_n12471_));
  NOR2_X1    g12385(.A1(new_n12471_), .A2(new_n12259_), .ZN(new_n12472_));
  OAI21_X1   g12386(.A1(new_n12472_), .A2(new_n12470_), .B(new_n12468_), .ZN(new_n12473_));
  NOR3_X1    g12387(.A1(new_n12472_), .A2(new_n12468_), .A3(new_n12470_), .ZN(new_n12474_));
  INV_X1     g12388(.I(new_n12474_), .ZN(new_n12475_));
  AOI22_X1   g12389(.A1(new_n11632_), .A2(new_n7838_), .B1(new_n10857_), .B2(new_n2469_), .ZN(new_n12476_));
  OAI21_X1   g12390(.A1(new_n12476_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n12477_));
  XNOR2_X1   g12391(.A1(new_n11631_), .A2(new_n12477_), .ZN(new_n12478_));
  INV_X1     g12392(.I(new_n12478_), .ZN(new_n12479_));
  NAND3_X1   g12393(.A1(new_n12475_), .A2(new_n12473_), .A3(new_n12479_), .ZN(new_n12480_));
  INV_X1     g12394(.I(new_n12473_), .ZN(new_n12481_));
  OAI21_X1   g12395(.A1(new_n12481_), .A2(new_n12474_), .B(new_n12478_), .ZN(new_n12482_));
  NAND4_X1   g12396(.A1(new_n12463_), .A2(new_n12482_), .A3(new_n12480_), .A4(new_n12467_), .ZN(new_n12483_));
  INV_X1     g12397(.I(new_n12483_), .ZN(new_n12484_));
  NAND2_X1   g12398(.A1(new_n12484_), .A2(new_n12271_), .ZN(new_n12485_));
  OAI22_X1   g12399(.A1(new_n10870_), .A2(new_n2495_), .B1(new_n7837_), .B2(new_n10861_), .ZN(new_n12486_));
  AOI21_X1   g12400(.A1(new_n12486_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12487_));
  XOR2_X1    g12401(.A1(new_n11648_), .A2(new_n12487_), .Z(new_n12488_));
  NOR2_X1    g12402(.A1(new_n12482_), .A2(new_n12488_), .ZN(new_n12489_));
  OAI21_X1   g12403(.A1(new_n12484_), .A2(new_n12271_), .B(new_n12489_), .ZN(new_n12490_));
  NAND2_X1   g12404(.A1(new_n12490_), .A2(new_n12485_), .ZN(new_n12491_));
  INV_X1     g12405(.I(new_n12018_), .ZN(new_n12492_));
  OAI21_X1   g12406(.A1(new_n12492_), .A2(new_n12020_), .B(new_n12008_), .ZN(new_n12493_));
  INV_X1     g12407(.I(new_n12493_), .ZN(new_n12494_));
  NAND3_X1   g12408(.A1(new_n12012_), .A2(new_n12013_), .A3(new_n12017_), .ZN(new_n12495_));
  INV_X1     g12409(.I(new_n12017_), .ZN(new_n12496_));
  NAND2_X1   g12410(.A1(new_n12014_), .A2(new_n12496_), .ZN(new_n12497_));
  AOI21_X1   g12411(.A1(new_n12495_), .A2(new_n12497_), .B(new_n12008_), .ZN(new_n12498_));
  AOI22_X1   g12412(.A1(new_n11724_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n10875_), .ZN(new_n12499_));
  OAI21_X1   g12413(.A1(new_n12499_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n12500_));
  XNOR2_X1   g12414(.A1(new_n11722_), .A2(new_n12500_), .ZN(new_n12501_));
  INV_X1     g12415(.I(new_n12501_), .ZN(new_n12502_));
  NOR3_X1    g12416(.A1(new_n12494_), .A2(new_n12498_), .A3(new_n12502_), .ZN(new_n12503_));
  INV_X1     g12417(.I(new_n12503_), .ZN(new_n12504_));
  NAND2_X1   g12418(.A1(new_n12504_), .A2(new_n12491_), .ZN(new_n12505_));
  NOR2_X1    g12419(.A1(new_n12494_), .A2(new_n12498_), .ZN(new_n12506_));
  NOR2_X1    g12420(.A1(new_n12506_), .A2(new_n12501_), .ZN(new_n12507_));
  INV_X1     g12421(.I(new_n12507_), .ZN(new_n12508_));
  INV_X1     g12422(.I(new_n12022_), .ZN(new_n12509_));
  OAI22_X1   g12423(.A1(new_n11803_), .A2(new_n7837_), .B1(new_n2495_), .B2(new_n10881_), .ZN(new_n12510_));
  AOI21_X1   g12424(.A1(new_n12510_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12511_));
  XNOR2_X1   g12425(.A1(new_n11802_), .A2(new_n12511_), .ZN(new_n12512_));
  NAND2_X1   g12426(.A1(new_n12244_), .A2(new_n12512_), .ZN(new_n12513_));
  INV_X1     g12427(.I(new_n12512_), .ZN(new_n12514_));
  NAND2_X1   g12428(.A1(new_n12037_), .A2(new_n12514_), .ZN(new_n12515_));
  AOI21_X1   g12429(.A1(new_n12513_), .A2(new_n12515_), .B(new_n12509_), .ZN(new_n12516_));
  NOR2_X1    g12430(.A1(new_n12037_), .A2(new_n12512_), .ZN(new_n12517_));
  NOR2_X1    g12431(.A1(new_n12244_), .A2(new_n12514_), .ZN(new_n12518_));
  OAI21_X1   g12432(.A1(new_n12517_), .A2(new_n12518_), .B(new_n12509_), .ZN(new_n12519_));
  INV_X1     g12433(.I(new_n12519_), .ZN(new_n12520_));
  NOR2_X1    g12434(.A1(new_n12520_), .A2(new_n12516_), .ZN(new_n12521_));
  NAND3_X1   g12435(.A1(new_n12521_), .A2(new_n12505_), .A3(new_n12508_), .ZN(new_n12522_));
  NOR2_X1    g12436(.A1(new_n12522_), .A2(new_n12256_), .ZN(new_n12523_));
  NAND2_X1   g12437(.A1(new_n12522_), .A2(new_n12256_), .ZN(new_n12524_));
  XOR2_X1    g12438(.A1(new_n12022_), .A2(new_n12037_), .Z(new_n12525_));
  NAND2_X1   g12439(.A1(new_n12525_), .A2(new_n12512_), .ZN(new_n12526_));
  OAI22_X1   g12440(.A1(new_n10619_), .A2(new_n2495_), .B1(new_n7837_), .B2(new_n10885_), .ZN(new_n12527_));
  AOI21_X1   g12441(.A1(new_n12527_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12528_));
  XOR2_X1    g12442(.A1(new_n12074_), .A2(new_n12528_), .Z(new_n12529_));
  NOR2_X1    g12443(.A1(new_n12526_), .A2(new_n12529_), .ZN(new_n12530_));
  AOI21_X1   g12444(.A1(new_n12524_), .A2(new_n12530_), .B(new_n12523_), .ZN(new_n12531_));
  NAND2_X1   g12445(.A1(new_n12044_), .A2(new_n12039_), .ZN(new_n12532_));
  XOR2_X1    g12446(.A1(new_n12050_), .A2(new_n12053_), .Z(new_n12533_));
  NAND2_X1   g12447(.A1(new_n12533_), .A2(new_n12532_), .ZN(new_n12534_));
  NAND2_X1   g12448(.A1(new_n12050_), .A2(new_n12053_), .ZN(new_n12535_));
  INV_X1     g12449(.I(new_n12055_), .ZN(new_n12536_));
  NAND2_X1   g12450(.A1(new_n12536_), .A2(new_n12535_), .ZN(new_n12537_));
  NAND3_X1   g12451(.A1(new_n12537_), .A2(new_n12039_), .A3(new_n12044_), .ZN(new_n12538_));
  OAI22_X1   g12452(.A1(new_n12091_), .A2(new_n7837_), .B1(new_n2495_), .B2(new_n10611_), .ZN(new_n12539_));
  AOI21_X1   g12453(.A1(new_n12539_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12540_));
  XOR2_X1    g12454(.A1(new_n12090_), .A2(new_n12540_), .Z(new_n12541_));
  INV_X1     g12455(.I(new_n12541_), .ZN(new_n12542_));
  AOI21_X1   g12456(.A1(new_n12538_), .A2(new_n12534_), .B(new_n12542_), .ZN(new_n12543_));
  NOR2_X1    g12457(.A1(new_n12531_), .A2(new_n12543_), .ZN(new_n12544_));
  NAND3_X1   g12458(.A1(new_n12538_), .A2(new_n12534_), .A3(new_n12542_), .ZN(new_n12545_));
  INV_X1     g12459(.I(new_n12545_), .ZN(new_n12546_));
  INV_X1     g12460(.I(new_n12056_), .ZN(new_n12547_));
  AOI22_X1   g12461(.A1(new_n10986_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n10897_), .ZN(new_n12548_));
  OAI21_X1   g12462(.A1(new_n12548_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n12549_));
  XOR2_X1    g12463(.A1(new_n10984_), .A2(new_n12549_), .Z(new_n12550_));
  XOR2_X1    g12464(.A1(new_n12219_), .A2(new_n12550_), .Z(new_n12551_));
  NAND2_X1   g12465(.A1(new_n12551_), .A2(new_n12547_), .ZN(new_n12552_));
  XOR2_X1    g12466(.A1(new_n12219_), .A2(new_n12550_), .Z(new_n12553_));
  OAI21_X1   g12467(.A1(new_n12547_), .A2(new_n12553_), .B(new_n12552_), .ZN(new_n12554_));
  NOR3_X1    g12468(.A1(new_n12554_), .A2(new_n12544_), .A3(new_n12546_), .ZN(new_n12555_));
  NAND2_X1   g12469(.A1(new_n12555_), .A2(new_n12241_), .ZN(new_n12556_));
  NOR2_X1    g12470(.A1(new_n12056_), .A2(new_n12219_), .ZN(new_n12557_));
  NOR2_X1    g12471(.A1(new_n12547_), .A2(new_n12064_), .ZN(new_n12558_));
  OAI21_X1   g12472(.A1(new_n12558_), .A2(new_n12557_), .B(new_n12550_), .ZN(new_n12559_));
  OAI22_X1   g12473(.A1(new_n10606_), .A2(new_n2495_), .B1(new_n7837_), .B2(new_n10901_), .ZN(new_n12560_));
  AOI21_X1   g12474(.A1(new_n12560_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12561_));
  XOR2_X1    g12475(.A1(new_n12211_), .A2(new_n12561_), .Z(new_n12562_));
  NOR2_X1    g12476(.A1(new_n12559_), .A2(new_n12562_), .ZN(new_n12563_));
  OAI21_X1   g12477(.A1(new_n12555_), .A2(new_n12241_), .B(new_n12563_), .ZN(new_n12564_));
  NOR2_X1    g12478(.A1(new_n12095_), .A2(new_n12097_), .ZN(new_n12565_));
  NAND2_X1   g12479(.A1(new_n12081_), .A2(new_n12565_), .ZN(new_n12566_));
  INV_X1     g12480(.I(new_n12565_), .ZN(new_n12567_));
  NAND2_X1   g12481(.A1(new_n12567_), .A2(new_n12223_), .ZN(new_n12568_));
  NAND2_X1   g12482(.A1(new_n10889_), .A2(new_n10899_), .ZN(new_n12569_));
  AOI22_X1   g12483(.A1(new_n12569_), .A2(new_n12204_), .B1(new_n10890_), .B2(new_n10901_), .ZN(new_n12570_));
  NAND2_X1   g12484(.A1(new_n12570_), .A2(new_n10606_), .ZN(new_n12571_));
  OAI21_X1   g12485(.A1(new_n10890_), .A2(new_n10900_), .B(new_n12204_), .ZN(new_n12572_));
  AOI21_X1   g12486(.A1(new_n12571_), .A2(new_n12572_), .B(new_n10599_), .ZN(new_n12573_));
  INV_X1     g12487(.I(new_n10902_), .ZN(new_n12574_));
  AOI21_X1   g12488(.A1(new_n12574_), .A2(new_n10898_), .B(new_n10600_), .ZN(new_n12575_));
  NOR2_X1    g12489(.A1(new_n12573_), .A2(new_n12575_), .ZN(new_n12576_));
  NOR2_X1    g12490(.A1(new_n10606_), .A2(new_n10896_), .ZN(new_n12577_));
  INV_X1     g12491(.I(new_n12577_), .ZN(new_n12578_));
  AOI22_X1   g12492(.A1(new_n12578_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n10600_), .ZN(new_n12579_));
  OAI21_X1   g12493(.A1(new_n12579_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n12580_));
  XNOR2_X1   g12494(.A1(new_n12576_), .A2(new_n12580_), .ZN(new_n12581_));
  NAND3_X1   g12495(.A1(new_n12566_), .A2(new_n12568_), .A3(new_n12581_), .ZN(new_n12582_));
  NOR2_X1    g12496(.A1(new_n12567_), .A2(new_n12223_), .ZN(new_n12583_));
  INV_X1     g12497(.I(new_n12568_), .ZN(new_n12584_));
  INV_X1     g12498(.I(new_n12581_), .ZN(new_n12585_));
  OAI21_X1   g12499(.A1(new_n12584_), .A2(new_n12583_), .B(new_n12585_), .ZN(new_n12586_));
  NOR3_X1    g12500(.A1(new_n12102_), .A2(new_n12099_), .A3(new_n12097_), .ZN(new_n12587_));
  NOR3_X1    g12501(.A1(new_n12587_), .A2(new_n12223_), .A3(new_n12565_), .ZN(new_n12588_));
  INV_X1     g12502(.I(new_n12097_), .ZN(new_n12589_));
  NAND2_X1   g12503(.A1(new_n12101_), .A2(new_n10989_), .ZN(new_n12590_));
  NAND2_X1   g12504(.A1(new_n11817_), .A2(new_n12098_), .ZN(new_n12591_));
  NAND3_X1   g12505(.A1(new_n12590_), .A2(new_n12591_), .A3(new_n12589_), .ZN(new_n12592_));
  AOI21_X1   g12506(.A1(new_n12592_), .A2(new_n12567_), .B(new_n12081_), .ZN(new_n12593_));
  NAND2_X1   g12507(.A1(new_n10903_), .A2(new_n10599_), .ZN(new_n12594_));
  NAND2_X1   g12508(.A1(new_n10898_), .A2(new_n10600_), .ZN(new_n12595_));
  AOI21_X1   g12509(.A1(new_n12594_), .A2(new_n12595_), .B(new_n10595_), .ZN(new_n12596_));
  NOR2_X1    g12510(.A1(new_n10898_), .A2(new_n10599_), .ZN(new_n12597_));
  OAI21_X1   g12511(.A1(new_n10904_), .A2(new_n12597_), .B(new_n10595_), .ZN(new_n12598_));
  INV_X1     g12512(.I(new_n12598_), .ZN(new_n12599_));
  NOR2_X1    g12513(.A1(new_n12599_), .A2(new_n12596_), .ZN(new_n12600_));
  NOR2_X1    g12514(.A1(new_n10606_), .A2(new_n10599_), .ZN(new_n12601_));
  OAI22_X1   g12515(.A1(new_n12601_), .A2(new_n7837_), .B1(new_n2495_), .B2(new_n10595_), .ZN(new_n12602_));
  AOI21_X1   g12516(.A1(new_n12602_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12603_));
  XOR2_X1    g12517(.A1(new_n12600_), .A2(new_n12603_), .Z(new_n12604_));
  NOR3_X1    g12518(.A1(new_n12588_), .A2(new_n12593_), .A3(new_n12604_), .ZN(new_n12605_));
  INV_X1     g12519(.I(new_n12588_), .ZN(new_n12606_));
  OAI21_X1   g12520(.A1(new_n12587_), .A2(new_n12565_), .B(new_n12223_), .ZN(new_n12607_));
  INV_X1     g12521(.I(new_n12604_), .ZN(new_n12608_));
  AOI21_X1   g12522(.A1(new_n12606_), .A2(new_n12607_), .B(new_n12608_), .ZN(new_n12609_));
  AOI22_X1   g12523(.A1(new_n12564_), .A2(new_n12556_), .B1(new_n12582_), .B2(new_n12586_), .ZN(new_n12611_));
  NAND2_X1   g12524(.A1(new_n12611_), .A2(new_n12231_), .ZN(new_n12612_));
  OAI21_X1   g12525(.A1(new_n12588_), .A2(new_n12593_), .B(new_n12604_), .ZN(new_n12613_));
  INV_X1     g12526(.I(new_n10595_), .ZN(new_n12614_));
  NAND2_X1   g12527(.A1(new_n12594_), .A2(new_n12595_), .ZN(new_n12615_));
  INV_X1     g12528(.I(new_n10589_), .ZN(new_n12616_));
  XOR2_X1    g12529(.A1(new_n10903_), .A2(new_n12616_), .Z(new_n12617_));
  NAND2_X1   g12530(.A1(new_n12617_), .A2(new_n12615_), .ZN(new_n12618_));
  NOR2_X1    g12531(.A1(new_n12618_), .A2(new_n12614_), .ZN(new_n12619_));
  NAND2_X1   g12532(.A1(new_n12618_), .A2(new_n12614_), .ZN(new_n12620_));
  INV_X1     g12533(.I(new_n12620_), .ZN(new_n12621_));
  NOR2_X1    g12534(.A1(new_n12621_), .A2(new_n12619_), .ZN(new_n12622_));
  NOR2_X1    g12535(.A1(new_n10595_), .A2(new_n10599_), .ZN(new_n12623_));
  OAI22_X1   g12536(.A1(new_n10589_), .A2(new_n2495_), .B1(new_n12623_), .B2(new_n7837_), .ZN(new_n12624_));
  AOI21_X1   g12537(.A1(new_n12624_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12625_));
  XOR2_X1    g12538(.A1(new_n12622_), .A2(new_n12625_), .Z(new_n12626_));
  NOR2_X1    g12539(.A1(new_n12613_), .A2(new_n12626_), .ZN(new_n12627_));
  OAI21_X1   g12540(.A1(new_n12611_), .A2(new_n12231_), .B(new_n12627_), .ZN(new_n12628_));
  NAND2_X1   g12541(.A1(new_n12628_), .A2(new_n12612_), .ZN(new_n12629_));
  NAND2_X1   g12542(.A1(new_n12202_), .A2(new_n12203_), .ZN(new_n12630_));
  INV_X1     g12543(.I(new_n12630_), .ZN(new_n12631_));
  NOR2_X1    g12544(.A1(new_n12224_), .A2(new_n12631_), .ZN(new_n12632_));
  INV_X1     g12545(.I(new_n12214_), .ZN(new_n12633_));
  NAND2_X1   g12546(.A1(new_n12227_), .A2(new_n12633_), .ZN(new_n12634_));
  AOI21_X1   g12547(.A1(new_n12224_), .A2(new_n12631_), .B(new_n12634_), .ZN(new_n12635_));
  NOR2_X1    g12548(.A1(new_n12635_), .A2(new_n12632_), .ZN(new_n12636_));
  NAND2_X1   g12549(.A1(new_n12186_), .A2(new_n12196_), .ZN(new_n12637_));
  NOR2_X1    g12550(.A1(new_n12186_), .A2(new_n12196_), .ZN(new_n12638_));
  NAND2_X1   g12551(.A1(new_n11812_), .A2(new_n12190_), .ZN(new_n12639_));
  OAI21_X1   g12552(.A1(new_n12638_), .A2(new_n12639_), .B(new_n12637_), .ZN(new_n12640_));
  NOR2_X1    g12553(.A1(new_n12173_), .A2(new_n12166_), .ZN(new_n12641_));
  NOR3_X1    g12554(.A1(new_n11808_), .A2(new_n11733_), .A3(new_n12641_), .ZN(new_n12642_));
  NAND2_X1   g12555(.A1(new_n11796_), .A2(new_n11734_), .ZN(new_n12643_));
  NOR2_X1    g12556(.A1(new_n12110_), .A2(new_n12176_), .ZN(new_n12644_));
  INV_X1     g12557(.I(new_n12644_), .ZN(new_n12645_));
  AOI21_X1   g12558(.A1(new_n12643_), .A2(new_n12641_), .B(new_n12645_), .ZN(new_n12646_));
  INV_X1     g12559(.I(new_n12164_), .ZN(new_n12647_));
  OAI21_X1   g12560(.A1(new_n12114_), .A2(new_n12162_), .B(new_n12647_), .ZN(new_n12648_));
  INV_X1     g12561(.I(new_n12149_), .ZN(new_n12649_));
  INV_X1     g12562(.I(new_n12151_), .ZN(new_n12650_));
  AOI21_X1   g12563(.A1(new_n12650_), .A2(new_n11768_), .B(new_n11772_), .ZN(new_n12651_));
  OAI21_X1   g12564(.A1(new_n12650_), .A2(new_n11768_), .B(new_n11743_), .ZN(new_n12652_));
  NOR2_X1    g12565(.A1(new_n12651_), .A2(new_n12652_), .ZN(new_n12653_));
  NAND2_X1   g12566(.A1(new_n12117_), .A2(new_n12138_), .ZN(new_n12654_));
  NAND2_X1   g12567(.A1(new_n12654_), .A2(new_n12140_), .ZN(new_n12655_));
  AOI21_X1   g12568(.A1(new_n12130_), .A2(new_n12126_), .B(new_n12127_), .ZN(new_n12656_));
  OAI22_X1   g12569(.A1(new_n10725_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10777_), .ZN(new_n12657_));
  OAI21_X1   g12570(.A1(new_n10696_), .A2(new_n79_), .B(new_n12657_), .ZN(new_n12658_));
  AOI21_X1   g12571(.A1(new_n12658_), .A2(new_n72_), .B(new_n79_), .ZN(new_n12659_));
  XOR2_X1    g12572(.A1(new_n11064_), .A2(new_n12659_), .Z(new_n12660_));
  AOI22_X1   g12573(.A1(new_n10783_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n10780_), .ZN(new_n12661_));
  AOI21_X1   g12574(.A1(new_n962_), .A2(new_n11002_), .B(new_n12661_), .ZN(new_n12662_));
  OR2_X2     g12575(.A1(new_n12662_), .A2(new_n11009_), .Z(new_n12663_));
  AOI21_X1   g12576(.A1(new_n12662_), .A2(new_n11009_), .B(new_n11002_), .ZN(new_n12664_));
  AOI21_X1   g12577(.A1(new_n12663_), .A2(new_n12664_), .B(new_n82_), .ZN(new_n12665_));
  XNOR2_X1   g12578(.A1(new_n12665_), .A2(new_n12125_), .ZN(new_n12666_));
  XOR2_X1    g12579(.A1(new_n12660_), .A2(new_n12666_), .Z(new_n12667_));
  INV_X1     g12580(.I(new_n12666_), .ZN(new_n12668_));
  NOR2_X1    g12581(.A1(new_n12660_), .A2(new_n12668_), .ZN(new_n12669_));
  NAND2_X1   g12582(.A1(new_n12660_), .A2(new_n12668_), .ZN(new_n12670_));
  INV_X1     g12583(.I(new_n12670_), .ZN(new_n12671_));
  OAI21_X1   g12584(.A1(new_n12671_), .A2(new_n12669_), .B(new_n12656_), .ZN(new_n12672_));
  OAI21_X1   g12585(.A1(new_n12656_), .A2(new_n12667_), .B(new_n12672_), .ZN(new_n12673_));
  OAI22_X1   g12586(.A1(new_n10672_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10792_), .ZN(new_n12674_));
  OAI21_X1   g12587(.A1(new_n1128_), .A2(new_n10658_), .B(new_n12674_), .ZN(new_n12675_));
  AOI21_X1   g12588(.A1(new_n12675_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n12676_));
  XOR2_X1    g12589(.A1(new_n11175_), .A2(new_n12676_), .Z(new_n12677_));
  INV_X1     g12590(.I(new_n12677_), .ZN(new_n12678_));
  XOR2_X1    g12591(.A1(new_n12673_), .A2(new_n12678_), .Z(new_n12679_));
  NAND2_X1   g12592(.A1(new_n12679_), .A2(new_n12655_), .ZN(new_n12680_));
  INV_X1     g12593(.I(new_n12655_), .ZN(new_n12681_));
  NOR2_X1    g12594(.A1(new_n12673_), .A2(new_n12678_), .ZN(new_n12682_));
  NAND2_X1   g12595(.A1(new_n12673_), .A2(new_n12678_), .ZN(new_n12683_));
  INV_X1     g12596(.I(new_n12683_), .ZN(new_n12684_));
  OAI21_X1   g12597(.A1(new_n12682_), .A2(new_n12684_), .B(new_n12681_), .ZN(new_n12685_));
  NAND2_X1   g12598(.A1(new_n12685_), .A2(new_n12680_), .ZN(new_n12686_));
  AOI22_X1   g12599(.A1(new_n10638_), .A2(new_n247_), .B1(new_n5783_), .B2(new_n11269_), .ZN(new_n12687_));
  NOR2_X1    g12600(.A1(new_n12687_), .A2(\a[23] ), .ZN(new_n12688_));
  NOR2_X1    g12601(.A1(new_n12688_), .A2(new_n1239_), .ZN(new_n12689_));
  XNOR2_X1   g12602(.A1(new_n11268_), .A2(new_n12689_), .ZN(new_n12690_));
  INV_X1     g12603(.I(new_n12690_), .ZN(new_n12691_));
  NAND2_X1   g12604(.A1(new_n12686_), .A2(new_n12691_), .ZN(new_n12692_));
  NOR2_X1    g12605(.A1(new_n12653_), .A2(new_n12692_), .ZN(new_n12693_));
  NAND2_X1   g12606(.A1(new_n12653_), .A2(new_n12692_), .ZN(new_n12694_));
  INV_X1     g12607(.I(new_n12694_), .ZN(new_n12695_));
  OAI21_X1   g12608(.A1(new_n12695_), .A2(new_n12693_), .B(new_n12649_), .ZN(new_n12696_));
  INV_X1     g12609(.I(new_n12693_), .ZN(new_n12697_));
  NAND3_X1   g12610(.A1(new_n12697_), .A2(new_n12149_), .A3(new_n12694_), .ZN(new_n12698_));
  AOI22_X1   g12611(.A1(new_n4717_), .A2(new_n10843_), .B1(new_n11608_), .B2(new_n5337_), .ZN(new_n12699_));
  OAI21_X1   g12612(.A1(new_n12699_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n12700_));
  XOR2_X1    g12613(.A1(new_n11607_), .A2(new_n12700_), .Z(new_n12701_));
  INV_X1     g12614(.I(new_n12701_), .ZN(new_n12702_));
  AOI21_X1   g12615(.A1(new_n12696_), .A2(new_n12698_), .B(new_n12702_), .ZN(new_n12703_));
  AOI21_X1   g12616(.A1(new_n12697_), .A2(new_n12694_), .B(new_n12149_), .ZN(new_n12704_));
  INV_X1     g12617(.I(new_n12698_), .ZN(new_n12705_));
  NOR3_X1    g12618(.A1(new_n12705_), .A2(new_n12704_), .A3(new_n12701_), .ZN(new_n12706_));
  OAI21_X1   g12619(.A1(new_n12703_), .A2(new_n12706_), .B(new_n12648_), .ZN(new_n12707_));
  INV_X1     g12620(.I(new_n12707_), .ZN(new_n12708_));
  NOR3_X1    g12621(.A1(new_n12705_), .A2(new_n12704_), .A3(new_n12702_), .ZN(new_n12709_));
  AOI21_X1   g12622(.A1(new_n12696_), .A2(new_n12698_), .B(new_n12701_), .ZN(new_n12710_));
  NOR2_X1    g12623(.A1(new_n12709_), .A2(new_n12710_), .ZN(new_n12711_));
  NOR2_X1    g12624(.A1(new_n12711_), .A2(new_n12648_), .ZN(new_n12712_));
  AOI22_X1   g12625(.A1(new_n11724_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n10875_), .ZN(new_n12713_));
  OAI21_X1   g12626(.A1(new_n12713_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n12714_));
  XNOR2_X1   g12627(.A1(new_n11722_), .A2(new_n12714_), .ZN(new_n12715_));
  INV_X1     g12628(.I(new_n12715_), .ZN(new_n12716_));
  NOR3_X1    g12629(.A1(new_n12708_), .A2(new_n12712_), .A3(new_n12716_), .ZN(new_n12717_));
  INV_X1     g12630(.I(new_n12712_), .ZN(new_n12718_));
  AOI21_X1   g12631(.A1(new_n12718_), .A2(new_n12707_), .B(new_n12715_), .ZN(new_n12719_));
  NOR2_X1    g12632(.A1(new_n12717_), .A2(new_n12719_), .ZN(new_n12720_));
  NOR3_X1    g12633(.A1(new_n12646_), .A2(new_n12720_), .A3(new_n12642_), .ZN(new_n12721_));
  NAND2_X1   g12634(.A1(new_n12643_), .A2(new_n12641_), .ZN(new_n12722_));
  AOI21_X1   g12635(.A1(new_n12722_), .A2(new_n12644_), .B(new_n12642_), .ZN(new_n12723_));
  NAND3_X1   g12636(.A1(new_n12718_), .A2(new_n12707_), .A3(new_n12715_), .ZN(new_n12724_));
  OAI21_X1   g12637(.A1(new_n12708_), .A2(new_n12712_), .B(new_n12716_), .ZN(new_n12725_));
  NAND2_X1   g12638(.A1(new_n12725_), .A2(new_n12724_), .ZN(new_n12726_));
  NOR2_X1    g12639(.A1(new_n12723_), .A2(new_n12726_), .ZN(new_n12727_));
  OAI22_X1   g12640(.A1(new_n12091_), .A2(new_n5967_), .B1(new_n643_), .B2(new_n10611_), .ZN(new_n12728_));
  AOI21_X1   g12641(.A1(new_n12728_), .A2(new_n279_), .B(new_n643_), .ZN(new_n12729_));
  XOR2_X1    g12642(.A1(new_n12090_), .A2(new_n12729_), .Z(new_n12730_));
  OAI21_X1   g12643(.A1(new_n12727_), .A2(new_n12721_), .B(new_n12730_), .ZN(new_n12731_));
  NOR3_X1    g12644(.A1(new_n12727_), .A2(new_n12721_), .A3(new_n12730_), .ZN(new_n12732_));
  INV_X1     g12645(.I(new_n12732_), .ZN(new_n12733_));
  NAND2_X1   g12646(.A1(new_n12733_), .A2(new_n12731_), .ZN(new_n12734_));
  NAND2_X1   g12647(.A1(new_n12734_), .A2(new_n12640_), .ZN(new_n12735_));
  INV_X1     g12648(.I(new_n12640_), .ZN(new_n12736_));
  INV_X1     g12649(.I(new_n12721_), .ZN(new_n12737_));
  INV_X1     g12650(.I(new_n12727_), .ZN(new_n12738_));
  NAND2_X1   g12651(.A1(new_n12738_), .A2(new_n12737_), .ZN(new_n12739_));
  XOR2_X1    g12652(.A1(new_n12739_), .A2(new_n12730_), .Z(new_n12740_));
  NAND2_X1   g12653(.A1(new_n12740_), .A2(new_n12736_), .ZN(new_n12741_));
  AOI22_X1   g12654(.A1(new_n12578_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n10600_), .ZN(new_n12742_));
  OAI21_X1   g12655(.A1(new_n12742_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n12743_));
  XNOR2_X1   g12656(.A1(new_n12576_), .A2(new_n12743_), .ZN(new_n12744_));
  NAND3_X1   g12657(.A1(new_n12741_), .A2(new_n12735_), .A3(new_n12744_), .ZN(new_n12745_));
  INV_X1     g12658(.I(new_n12735_), .ZN(new_n12746_));
  XNOR2_X1   g12659(.A1(new_n12739_), .A2(new_n12730_), .ZN(new_n12747_));
  NOR2_X1    g12660(.A1(new_n12747_), .A2(new_n12640_), .ZN(new_n12748_));
  INV_X1     g12661(.I(new_n12744_), .ZN(new_n12749_));
  OAI21_X1   g12662(.A1(new_n12748_), .A2(new_n12746_), .B(new_n12749_), .ZN(new_n12750_));
  NAND2_X1   g12663(.A1(new_n12750_), .A2(new_n12745_), .ZN(new_n12751_));
  NAND2_X1   g12664(.A1(new_n12636_), .A2(new_n12751_), .ZN(new_n12752_));
  NAND2_X1   g12665(.A1(new_n12105_), .A2(new_n12630_), .ZN(new_n12753_));
  NOR2_X1    g12666(.A1(new_n11818_), .A2(new_n12214_), .ZN(new_n12754_));
  OAI21_X1   g12667(.A1(new_n12105_), .A2(new_n12630_), .B(new_n12754_), .ZN(new_n12755_));
  NAND2_X1   g12668(.A1(new_n12755_), .A2(new_n12753_), .ZN(new_n12756_));
  NOR3_X1    g12669(.A1(new_n12748_), .A2(new_n12746_), .A3(new_n12749_), .ZN(new_n12757_));
  AOI21_X1   g12670(.A1(new_n12741_), .A2(new_n12735_), .B(new_n12744_), .ZN(new_n12758_));
  NOR2_X1    g12671(.A1(new_n12757_), .A2(new_n12758_), .ZN(new_n12759_));
  NAND2_X1   g12672(.A1(new_n12756_), .A2(new_n12759_), .ZN(new_n12760_));
  NOR2_X1    g12673(.A1(new_n10905_), .A2(new_n10906_), .ZN(new_n12761_));
  NAND2_X1   g12674(.A1(new_n12761_), .A2(new_n10589_), .ZN(new_n12762_));
  OAI21_X1   g12675(.A1(new_n10905_), .A2(new_n10906_), .B(new_n12616_), .ZN(new_n12763_));
  AOI21_X1   g12676(.A1(new_n12762_), .A2(new_n12763_), .B(new_n10913_), .ZN(new_n12764_));
  INV_X1     g12677(.I(new_n10915_), .ZN(new_n12765_));
  AOI21_X1   g12678(.A1(new_n12765_), .A2(new_n10907_), .B(new_n10914_), .ZN(new_n12766_));
  NOR2_X1    g12679(.A1(new_n12766_), .A2(new_n12764_), .ZN(new_n12767_));
  NOR2_X1    g12680(.A1(new_n10589_), .A2(new_n10595_), .ZN(new_n12768_));
  OAI22_X1   g12681(.A1(new_n10913_), .A2(new_n2495_), .B1(new_n12768_), .B2(new_n7837_), .ZN(new_n12769_));
  AOI21_X1   g12682(.A1(new_n12769_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n12770_));
  XOR2_X1    g12683(.A1(new_n12767_), .A2(new_n12770_), .Z(new_n12771_));
  INV_X1     g12684(.I(new_n12771_), .ZN(new_n12772_));
  NAND3_X1   g12685(.A1(new_n12760_), .A2(new_n12752_), .A3(new_n12772_), .ZN(new_n12773_));
  INV_X1     g12686(.I(new_n12773_), .ZN(new_n12774_));
  AOI21_X1   g12687(.A1(new_n12760_), .A2(new_n12752_), .B(new_n12772_), .ZN(new_n12775_));
  NOR2_X1    g12688(.A1(new_n12774_), .A2(new_n12775_), .ZN(new_n12776_));
  NOR2_X1    g12689(.A1(new_n12199_), .A2(new_n12108_), .ZN(new_n12777_));
  AOI21_X1   g12690(.A1(new_n12199_), .A2(new_n12108_), .B(new_n12639_), .ZN(new_n12778_));
  OAI21_X1   g12691(.A1(new_n12778_), .A2(new_n12777_), .B(new_n12731_), .ZN(new_n12779_));
  NAND2_X1   g12692(.A1(new_n12779_), .A2(new_n12733_), .ZN(new_n12780_));
  INV_X1     g12693(.I(new_n12703_), .ZN(new_n12781_));
  AOI21_X1   g12694(.A1(new_n12648_), .A2(new_n12781_), .B(new_n12706_), .ZN(new_n12782_));
  INV_X1     g12695(.I(new_n12686_), .ZN(new_n12783_));
  AOI21_X1   g12696(.A1(new_n12783_), .A2(new_n12649_), .B(new_n12690_), .ZN(new_n12784_));
  AOI22_X1   g12697(.A1(new_n12653_), .A2(new_n12784_), .B1(new_n12149_), .B2(new_n12686_), .ZN(new_n12785_));
  OAI22_X1   g12698(.A1(new_n11386_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n10633_), .ZN(new_n12786_));
  AOI21_X1   g12699(.A1(new_n12786_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n12787_));
  XOR2_X1    g12700(.A1(new_n11385_), .A2(new_n12787_), .Z(new_n12788_));
  OAI21_X1   g12701(.A1(new_n12656_), .A2(new_n12669_), .B(new_n12670_), .ZN(new_n12789_));
  INV_X1     g12702(.I(new_n12789_), .ZN(new_n12790_));
  AOI22_X1   g12703(.A1(new_n10794_), .A2(new_n4526_), .B1(new_n4570_), .B2(new_n10809_), .ZN(new_n12791_));
  AOI21_X1   g12704(.A1(new_n101_), .A2(new_n10691_), .B(new_n12791_), .ZN(new_n12792_));
  OAI21_X1   g12705(.A1(new_n12792_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n12793_));
  XOR2_X1    g12706(.A1(new_n11333_), .A2(new_n12793_), .Z(new_n12794_));
  NAND2_X1   g12707(.A1(new_n12665_), .A2(new_n12125_), .ZN(new_n12795_));
  NOR2_X1    g12708(.A1(new_n10762_), .A2(new_n88_), .ZN(new_n12796_));
  OAI21_X1   g12709(.A1(new_n511_), .A2(new_n10777_), .B(new_n12124_), .ZN(new_n12797_));
  OAI21_X1   g12710(.A1(new_n12797_), .A2(new_n12796_), .B(new_n961_), .ZN(new_n12798_));
  NOR2_X1    g12711(.A1(new_n12798_), .A2(new_n11188_), .ZN(new_n12799_));
  XOR2_X1    g12712(.A1(new_n12795_), .A2(new_n12799_), .Z(new_n12800_));
  XNOR2_X1   g12713(.A1(new_n12794_), .A2(new_n12800_), .ZN(new_n12801_));
  NAND2_X1   g12714(.A1(new_n12794_), .A2(new_n12800_), .ZN(new_n12802_));
  INV_X1     g12715(.I(new_n12802_), .ZN(new_n12803_));
  NOR2_X1    g12716(.A1(new_n12794_), .A2(new_n12800_), .ZN(new_n12804_));
  OAI21_X1   g12717(.A1(new_n12803_), .A2(new_n12804_), .B(new_n12790_), .ZN(new_n12805_));
  OAI21_X1   g12718(.A1(new_n12790_), .A2(new_n12801_), .B(new_n12805_), .ZN(new_n12806_));
  AOI22_X1   g12719(.A1(new_n10805_), .A2(new_n4767_), .B1(new_n4613_), .B2(new_n10817_), .ZN(new_n12807_));
  NOR2_X1    g12720(.A1(new_n11214_), .A2(new_n1128_), .ZN(new_n12808_));
  OAI21_X1   g12721(.A1(new_n12808_), .A2(new_n12807_), .B(new_n65_), .ZN(new_n12809_));
  NAND2_X1   g12722(.A1(new_n12809_), .A2(new_n117_), .ZN(new_n12810_));
  XNOR2_X1   g12723(.A1(new_n11224_), .A2(new_n12810_), .ZN(new_n12811_));
  XNOR2_X1   g12724(.A1(new_n12806_), .A2(new_n12811_), .ZN(new_n12812_));
  NAND2_X1   g12725(.A1(new_n12812_), .A2(new_n12679_), .ZN(new_n12813_));
  XOR2_X1    g12726(.A1(new_n12813_), .A2(new_n12683_), .Z(new_n12814_));
  NAND2_X1   g12727(.A1(new_n12814_), .A2(new_n12681_), .ZN(new_n12815_));
  INV_X1     g12728(.I(new_n12815_), .ZN(new_n12816_));
  NOR2_X1    g12729(.A1(new_n12814_), .A2(new_n12681_), .ZN(new_n12817_));
  NOR3_X1    g12730(.A1(new_n12816_), .A2(new_n12788_), .A3(new_n12817_), .ZN(new_n12818_));
  INV_X1     g12731(.I(new_n12788_), .ZN(new_n12819_));
  INV_X1     g12732(.I(new_n12817_), .ZN(new_n12820_));
  AOI21_X1   g12733(.A1(new_n12820_), .A2(new_n12815_), .B(new_n12819_), .ZN(new_n12821_));
  NOR2_X1    g12734(.A1(new_n12821_), .A2(new_n12818_), .ZN(new_n12822_));
  NOR2_X1    g12735(.A1(new_n12822_), .A2(new_n12785_), .ZN(new_n12823_));
  NOR3_X1    g12736(.A1(new_n12816_), .A2(new_n12819_), .A3(new_n12817_), .ZN(new_n12824_));
  AOI21_X1   g12737(.A1(new_n12820_), .A2(new_n12815_), .B(new_n12788_), .ZN(new_n12825_));
  OAI21_X1   g12738(.A1(new_n12824_), .A2(new_n12825_), .B(new_n12785_), .ZN(new_n12826_));
  INV_X1     g12739(.I(new_n12826_), .ZN(new_n12827_));
  AOI22_X1   g12740(.A1(new_n11632_), .A2(new_n5337_), .B1(new_n10857_), .B2(new_n4717_), .ZN(new_n12828_));
  OAI21_X1   g12741(.A1(new_n12828_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n12829_));
  XNOR2_X1   g12742(.A1(new_n11631_), .A2(new_n12829_), .ZN(new_n12830_));
  NOR3_X1    g12743(.A1(new_n12823_), .A2(new_n12827_), .A3(new_n12830_), .ZN(new_n12831_));
  OR2_X2     g12744(.A1(new_n12651_), .A2(new_n12652_), .Z(new_n12832_));
  INV_X1     g12745(.I(new_n12784_), .ZN(new_n12833_));
  OAI22_X1   g12746(.A1(new_n12832_), .A2(new_n12833_), .B1(new_n12649_), .B2(new_n12783_), .ZN(new_n12834_));
  OAI21_X1   g12747(.A1(new_n12818_), .A2(new_n12821_), .B(new_n12834_), .ZN(new_n12835_));
  INV_X1     g12748(.I(new_n12830_), .ZN(new_n12836_));
  AOI21_X1   g12749(.A1(new_n12835_), .A2(new_n12826_), .B(new_n12836_), .ZN(new_n12837_));
  NOR2_X1    g12750(.A1(new_n12831_), .A2(new_n12837_), .ZN(new_n12838_));
  NAND2_X1   g12751(.A1(new_n12782_), .A2(new_n12838_), .ZN(new_n12839_));
  NOR2_X1    g12752(.A1(new_n12782_), .A2(new_n12838_), .ZN(new_n12840_));
  INV_X1     g12753(.I(new_n12840_), .ZN(new_n12841_));
  OAI22_X1   g12754(.A1(new_n11803_), .A2(new_n5420_), .B1(new_n1620_), .B2(new_n10881_), .ZN(new_n12842_));
  AOI21_X1   g12755(.A1(new_n12842_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n12843_));
  XNOR2_X1   g12756(.A1(new_n11802_), .A2(new_n12843_), .ZN(new_n12844_));
  NAND3_X1   g12757(.A1(new_n12841_), .A2(new_n12839_), .A3(new_n12844_), .ZN(new_n12845_));
  INV_X1     g12758(.I(new_n12839_), .ZN(new_n12846_));
  INV_X1     g12759(.I(new_n12844_), .ZN(new_n12847_));
  OAI21_X1   g12760(.A1(new_n12846_), .A2(new_n12840_), .B(new_n12847_), .ZN(new_n12848_));
  NAND3_X1   g12761(.A1(new_n12848_), .A2(new_n12845_), .A3(new_n12724_), .ZN(new_n12849_));
  NAND3_X1   g12762(.A1(new_n12849_), .A2(new_n12723_), .A3(new_n12726_), .ZN(new_n12850_));
  INV_X1     g12763(.I(new_n12642_), .ZN(new_n12851_));
  NAND2_X1   g12764(.A1(new_n12722_), .A2(new_n12644_), .ZN(new_n12852_));
  NAND2_X1   g12765(.A1(new_n12852_), .A2(new_n12851_), .ZN(new_n12853_));
  NOR3_X1    g12766(.A1(new_n12846_), .A2(new_n12840_), .A3(new_n12847_), .ZN(new_n12854_));
  AOI21_X1   g12767(.A1(new_n12841_), .A2(new_n12839_), .B(new_n12844_), .ZN(new_n12855_));
  NOR3_X1    g12768(.A1(new_n12855_), .A2(new_n12854_), .A3(new_n12717_), .ZN(new_n12856_));
  OAI21_X1   g12769(.A1(new_n12856_), .A2(new_n12720_), .B(new_n12853_), .ZN(new_n12857_));
  AOI22_X1   g12770(.A1(new_n10986_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n10897_), .ZN(new_n12858_));
  OAI21_X1   g12771(.A1(new_n12858_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n12859_));
  XOR2_X1    g12772(.A1(new_n10984_), .A2(new_n12859_), .Z(new_n12860_));
  INV_X1     g12773(.I(new_n12860_), .ZN(new_n12861_));
  NAND3_X1   g12774(.A1(new_n12857_), .A2(new_n12850_), .A3(new_n12861_), .ZN(new_n12862_));
  NOR3_X1    g12775(.A1(new_n12853_), .A2(new_n12856_), .A3(new_n12720_), .ZN(new_n12863_));
  AOI21_X1   g12776(.A1(new_n12849_), .A2(new_n12726_), .B(new_n12723_), .ZN(new_n12864_));
  OAI21_X1   g12777(.A1(new_n12863_), .A2(new_n12864_), .B(new_n12860_), .ZN(new_n12865_));
  NAND2_X1   g12778(.A1(new_n12862_), .A2(new_n12865_), .ZN(new_n12866_));
  NOR2_X1    g12779(.A1(new_n12780_), .A2(new_n12866_), .ZN(new_n12867_));
  AOI21_X1   g12780(.A1(new_n12640_), .A2(new_n12731_), .B(new_n12732_), .ZN(new_n12868_));
  NOR3_X1    g12781(.A1(new_n12863_), .A2(new_n12864_), .A3(new_n12860_), .ZN(new_n12869_));
  AOI21_X1   g12782(.A1(new_n12857_), .A2(new_n12850_), .B(new_n12861_), .ZN(new_n12870_));
  NOR2_X1    g12783(.A1(new_n12870_), .A2(new_n12869_), .ZN(new_n12871_));
  NOR2_X1    g12784(.A1(new_n12868_), .A2(new_n12871_), .ZN(new_n12872_));
  OAI22_X1   g12785(.A1(new_n12601_), .A2(new_n6757_), .B1(new_n1078_), .B2(new_n10595_), .ZN(new_n12873_));
  AOI21_X1   g12786(.A1(new_n12873_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n12874_));
  XOR2_X1    g12787(.A1(new_n12600_), .A2(new_n12874_), .Z(new_n12875_));
  INV_X1     g12788(.I(new_n12875_), .ZN(new_n12876_));
  NOR3_X1    g12789(.A1(new_n12872_), .A2(new_n12867_), .A3(new_n12876_), .ZN(new_n12877_));
  OAI21_X1   g12790(.A1(new_n12867_), .A2(new_n12872_), .B(new_n12876_), .ZN(new_n12878_));
  INV_X1     g12791(.I(new_n12878_), .ZN(new_n12879_));
  NOR3_X1    g12792(.A1(new_n12879_), .A2(new_n12757_), .A3(new_n12877_), .ZN(new_n12880_));
  NOR3_X1    g12793(.A1(new_n12880_), .A2(new_n12756_), .A3(new_n12759_), .ZN(new_n12881_));
  INV_X1     g12794(.I(new_n12877_), .ZN(new_n12882_));
  NAND3_X1   g12795(.A1(new_n12882_), .A2(new_n12745_), .A3(new_n12878_), .ZN(new_n12883_));
  AOI21_X1   g12796(.A1(new_n12883_), .A2(new_n12751_), .B(new_n12636_), .ZN(new_n12884_));
  XNOR2_X1   g12797(.A1(new_n10923_), .A2(new_n10913_), .ZN(new_n12885_));
  INV_X1     g12798(.I(new_n12885_), .ZN(new_n12886_));
  INV_X1     g12799(.I(new_n10928_), .ZN(new_n12887_));
  AOI21_X1   g12800(.A1(new_n10926_), .A2(new_n12887_), .B(new_n10916_), .ZN(new_n12888_));
  AOI21_X1   g12801(.A1(new_n10916_), .A2(new_n12886_), .B(new_n12888_), .ZN(new_n12889_));
  NOR2_X1    g12802(.A1(new_n10913_), .A2(new_n10589_), .ZN(new_n12890_));
  INV_X1     g12803(.I(new_n12890_), .ZN(new_n12891_));
  AOI22_X1   g12804(.A1(new_n12891_), .A2(new_n7838_), .B1(new_n10924_), .B2(new_n2469_), .ZN(new_n12892_));
  OAI21_X1   g12805(.A1(new_n12892_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n12893_));
  XNOR2_X1   g12806(.A1(new_n12889_), .A2(new_n12893_), .ZN(new_n12894_));
  NOR3_X1    g12807(.A1(new_n12884_), .A2(new_n12881_), .A3(new_n12894_), .ZN(new_n12895_));
  NAND3_X1   g12808(.A1(new_n12883_), .A2(new_n12636_), .A3(new_n12751_), .ZN(new_n12896_));
  OAI21_X1   g12809(.A1(new_n12880_), .A2(new_n12759_), .B(new_n12756_), .ZN(new_n12897_));
  INV_X1     g12810(.I(new_n12894_), .ZN(new_n12898_));
  AOI21_X1   g12811(.A1(new_n12897_), .A2(new_n12896_), .B(new_n12898_), .ZN(new_n12899_));
  NOR3_X1    g12812(.A1(new_n12895_), .A2(new_n12899_), .A3(new_n12775_), .ZN(new_n12900_));
  NOR3_X1    g12813(.A1(new_n12900_), .A2(new_n12776_), .A3(new_n12629_), .ZN(new_n12901_));
  INV_X1     g12814(.I(new_n12629_), .ZN(new_n12902_));
  NOR2_X1    g12815(.A1(new_n12900_), .A2(new_n12776_), .ZN(new_n12903_));
  NOR2_X1    g12816(.A1(new_n12903_), .A2(new_n12902_), .ZN(new_n12904_));
  XNOR2_X1   g12817(.A1(new_n10937_), .A2(new_n10949_), .ZN(new_n12905_));
  OAI21_X1   g12818(.A1(new_n10950_), .A2(new_n10953_), .B(new_n10941_), .ZN(new_n12906_));
  OAI21_X1   g12819(.A1(new_n10941_), .A2(new_n12905_), .B(new_n12906_), .ZN(new_n12907_));
  NOR2_X1    g12820(.A1(new_n10583_), .A2(new_n10938_), .ZN(new_n12908_));
  INV_X1     g12821(.I(new_n12908_), .ZN(new_n12909_));
  AOI22_X1   g12822(.A1(new_n12909_), .A2(new_n8832_), .B1(new_n10949_), .B2(new_n2898_), .ZN(new_n12910_));
  OAI21_X1   g12823(.A1(new_n12910_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n12911_));
  XOR2_X1    g12824(.A1(new_n12907_), .A2(new_n12911_), .Z(new_n12912_));
  INV_X1     g12825(.I(new_n12912_), .ZN(new_n12913_));
  NOR3_X1    g12826(.A1(new_n12904_), .A2(new_n12901_), .A3(new_n12913_), .ZN(new_n12914_));
  INV_X1     g12827(.I(new_n12914_), .ZN(new_n12915_));
  NAND2_X1   g12828(.A1(new_n12564_), .A2(new_n12556_), .ZN(new_n12916_));
  AND2_X2    g12829(.A1(new_n12586_), .A2(new_n12582_), .Z(new_n12917_));
  NOR2_X1    g12830(.A1(new_n12917_), .A2(new_n12916_), .ZN(new_n12918_));
  AND2_X2    g12831(.A1(new_n12564_), .A2(new_n12556_), .Z(new_n12919_));
  NAND2_X1   g12832(.A1(new_n12586_), .A2(new_n12582_), .ZN(new_n12920_));
  NOR2_X1    g12833(.A1(new_n12919_), .A2(new_n12920_), .ZN(new_n12921_));
  OAI22_X1   g12834(.A1(new_n10913_), .A2(new_n3040_), .B1(new_n12768_), .B2(new_n8831_), .ZN(new_n12922_));
  AOI21_X1   g12835(.A1(new_n12922_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n12923_));
  XOR2_X1    g12836(.A1(new_n12767_), .A2(new_n12923_), .Z(new_n12924_));
  NOR3_X1    g12837(.A1(new_n12921_), .A2(new_n12918_), .A3(new_n12924_), .ZN(new_n12925_));
  NAND2_X1   g12838(.A1(new_n12919_), .A2(new_n12920_), .ZN(new_n12926_));
  NAND2_X1   g12839(.A1(new_n12917_), .A2(new_n12916_), .ZN(new_n12927_));
  INV_X1     g12840(.I(new_n12924_), .ZN(new_n12928_));
  AOI21_X1   g12841(.A1(new_n12926_), .A2(new_n12927_), .B(new_n12928_), .ZN(new_n12929_));
  OR2_X2     g12842(.A1(new_n12925_), .A2(new_n12929_), .Z(new_n12930_));
  NOR2_X1    g12843(.A1(new_n12544_), .A2(new_n12546_), .ZN(new_n12931_));
  INV_X1     g12844(.I(new_n12554_), .ZN(new_n12932_));
  NOR2_X1    g12845(.A1(new_n12932_), .A2(new_n12931_), .ZN(new_n12933_));
  NAND2_X1   g12846(.A1(new_n12538_), .A2(new_n12534_), .ZN(new_n12934_));
  NAND2_X1   g12847(.A1(new_n12934_), .A2(new_n12541_), .ZN(new_n12935_));
  AOI21_X1   g12848(.A1(new_n12935_), .A2(new_n12545_), .B(new_n12531_), .ZN(new_n12936_));
  INV_X1     g12849(.I(new_n12531_), .ZN(new_n12937_));
  NOR2_X1    g12850(.A1(new_n12934_), .A2(new_n12542_), .ZN(new_n12938_));
  AOI21_X1   g12851(.A1(new_n12538_), .A2(new_n12534_), .B(new_n12541_), .ZN(new_n12939_));
  NOR2_X1    g12852(.A1(new_n12938_), .A2(new_n12939_), .ZN(new_n12940_));
  NOR2_X1    g12853(.A1(new_n12940_), .A2(new_n12937_), .ZN(new_n12941_));
  NOR2_X1    g12854(.A1(new_n12941_), .A2(new_n12936_), .ZN(new_n12942_));
  INV_X1     g12855(.I(new_n12526_), .ZN(new_n12943_));
  OAI21_X1   g12856(.A1(new_n12253_), .A2(new_n12254_), .B(new_n12036_), .ZN(new_n12944_));
  NAND3_X1   g12857(.A1(new_n12251_), .A2(new_n12247_), .A3(new_n12242_), .ZN(new_n12945_));
  AOI21_X1   g12858(.A1(new_n12944_), .A2(new_n12945_), .B(new_n12529_), .ZN(new_n12946_));
  NAND2_X1   g12859(.A1(new_n12522_), .A2(new_n12946_), .ZN(new_n12947_));
  NAND2_X1   g12860(.A1(new_n12505_), .A2(new_n12508_), .ZN(new_n12948_));
  NAND2_X1   g12861(.A1(new_n12513_), .A2(new_n12515_), .ZN(new_n12949_));
  NAND2_X1   g12862(.A1(new_n12949_), .A2(new_n12022_), .ZN(new_n12950_));
  NAND2_X1   g12863(.A1(new_n12950_), .A2(new_n12519_), .ZN(new_n12951_));
  NOR2_X1    g12864(.A1(new_n12948_), .A2(new_n12951_), .ZN(new_n12952_));
  OAI21_X1   g12865(.A1(new_n12256_), .A2(new_n12529_), .B(new_n12952_), .ZN(new_n12953_));
  AOI21_X1   g12866(.A1(new_n12953_), .A2(new_n12947_), .B(new_n12943_), .ZN(new_n12954_));
  NOR3_X1    g12867(.A1(new_n12952_), .A2(new_n12256_), .A3(new_n12529_), .ZN(new_n12955_));
  NOR2_X1    g12868(.A1(new_n12522_), .A2(new_n12946_), .ZN(new_n12956_));
  NOR3_X1    g12869(.A1(new_n12955_), .A2(new_n12956_), .A3(new_n12526_), .ZN(new_n12957_));
  NOR2_X1    g12870(.A1(new_n12954_), .A2(new_n12957_), .ZN(new_n12958_));
  INV_X1     g12871(.I(new_n12446_), .ZN(new_n12959_));
  NAND3_X1   g12872(.A1(new_n12428_), .A2(new_n12421_), .A3(new_n12441_), .ZN(new_n12960_));
  OAI21_X1   g12873(.A1(new_n12440_), .A2(new_n12439_), .B(new_n12432_), .ZN(new_n12961_));
  AOI21_X1   g12874(.A1(new_n12961_), .A2(new_n12960_), .B(new_n11981_), .ZN(new_n12962_));
  NOR3_X1    g12875(.A1(new_n12440_), .A2(new_n12439_), .A3(new_n12432_), .ZN(new_n12963_));
  AOI21_X1   g12876(.A1(new_n12428_), .A2(new_n12421_), .B(new_n12441_), .ZN(new_n12964_));
  NOR3_X1    g12877(.A1(new_n12963_), .A2(new_n12964_), .A3(new_n11980_), .ZN(new_n12965_));
  OAI21_X1   g12878(.A1(new_n12965_), .A2(new_n12962_), .B(new_n12959_), .ZN(new_n12966_));
  OAI21_X1   g12879(.A1(new_n12963_), .A2(new_n12964_), .B(new_n11980_), .ZN(new_n12967_));
  NAND3_X1   g12880(.A1(new_n12961_), .A2(new_n12960_), .A3(new_n11981_), .ZN(new_n12968_));
  NAND3_X1   g12881(.A1(new_n12967_), .A2(new_n12968_), .A3(new_n12446_), .ZN(new_n12969_));
  NAND2_X1   g12882(.A1(new_n12966_), .A2(new_n12969_), .ZN(new_n12970_));
  NAND2_X1   g12883(.A1(new_n12382_), .A2(new_n12377_), .ZN(new_n12971_));
  NAND2_X1   g12884(.A1(new_n12388_), .A2(new_n12391_), .ZN(new_n12972_));
  NAND2_X1   g12885(.A1(new_n12972_), .A2(new_n12394_), .ZN(new_n12973_));
  NAND2_X1   g12886(.A1(new_n12971_), .A2(new_n12973_), .ZN(new_n12974_));
  NAND3_X1   g12887(.A1(new_n12387_), .A2(new_n12385_), .A3(new_n12391_), .ZN(new_n12975_));
  NAND2_X1   g12888(.A1(new_n12388_), .A2(new_n12393_), .ZN(new_n12976_));
  NAND2_X1   g12889(.A1(new_n12976_), .A2(new_n12975_), .ZN(new_n12977_));
  NAND3_X1   g12890(.A1(new_n12977_), .A2(new_n12377_), .A3(new_n12382_), .ZN(new_n12978_));
  NAND2_X1   g12891(.A1(new_n12974_), .A2(new_n12978_), .ZN(new_n12979_));
  INV_X1     g12892(.I(new_n12979_), .ZN(new_n12980_));
  INV_X1     g12893(.I(new_n12367_), .ZN(new_n12981_));
  NAND2_X1   g12894(.A1(new_n12364_), .A2(new_n12369_), .ZN(new_n12982_));
  INV_X1     g12895(.I(new_n12324_), .ZN(new_n12983_));
  NOR2_X1    g12896(.A1(new_n11046_), .A2(new_n12983_), .ZN(new_n12984_));
  AOI21_X1   g12897(.A1(new_n11039_), .A2(new_n11045_), .B(new_n12324_), .ZN(new_n12985_));
  NOR2_X1    g12898(.A1(new_n12984_), .A2(new_n12985_), .ZN(new_n12986_));
  NOR2_X1    g12899(.A1(new_n12986_), .A2(new_n12329_), .ZN(new_n12987_));
  NAND2_X1   g12900(.A1(new_n12987_), .A2(new_n11898_), .ZN(new_n12988_));
  AOI21_X1   g12901(.A1(new_n12982_), .A2(new_n12988_), .B(new_n12981_), .ZN(new_n12989_));
  NOR2_X1    g12902(.A1(new_n12987_), .A2(new_n11898_), .ZN(new_n12990_));
  INV_X1     g12903(.I(new_n12988_), .ZN(new_n12991_));
  NOR3_X1    g12904(.A1(new_n12991_), .A2(new_n12367_), .A3(new_n12990_), .ZN(new_n12992_));
  OAI21_X1   g12905(.A1(new_n12992_), .A2(new_n12989_), .B(new_n12370_), .ZN(new_n12993_));
  OAI21_X1   g12906(.A1(new_n12991_), .A2(new_n12990_), .B(new_n12367_), .ZN(new_n12994_));
  NAND3_X1   g12907(.A1(new_n12982_), .A2(new_n12981_), .A3(new_n12988_), .ZN(new_n12995_));
  NAND3_X1   g12908(.A1(new_n12994_), .A2(new_n12995_), .A3(new_n11906_), .ZN(new_n12996_));
  NAND2_X1   g12909(.A1(new_n12993_), .A2(new_n12996_), .ZN(new_n12997_));
  NOR2_X1    g12910(.A1(new_n12986_), .A2(new_n12329_), .ZN(new_n12998_));
  NAND3_X1   g12911(.A1(new_n12358_), .A2(new_n11903_), .A3(new_n12354_), .ZN(new_n12999_));
  OAI21_X1   g12912(.A1(new_n12355_), .A2(new_n12343_), .B(new_n12331_), .ZN(new_n13000_));
  NAND3_X1   g12913(.A1(new_n13000_), .A2(new_n12999_), .A3(new_n12363_), .ZN(new_n13001_));
  NAND2_X1   g12914(.A1(new_n13001_), .A2(new_n12998_), .ZN(new_n13002_));
  NAND2_X1   g12915(.A1(new_n12325_), .A2(new_n12330_), .ZN(new_n13003_));
  INV_X1     g12916(.I(new_n12363_), .ZN(new_n13004_));
  NOR3_X1    g12917(.A1(new_n12356_), .A2(new_n12359_), .A3(new_n13004_), .ZN(new_n13005_));
  NAND2_X1   g12918(.A1(new_n13003_), .A2(new_n13005_), .ZN(new_n13006_));
  AOI21_X1   g12919(.A1(new_n13006_), .A2(new_n13002_), .B(new_n12356_), .ZN(new_n13007_));
  NOR2_X1    g12920(.A1(new_n12998_), .A2(new_n12999_), .ZN(new_n13008_));
  AOI22_X1   g12921(.A1(new_n10817_), .A2(new_n2898_), .B1(new_n12314_), .B2(new_n8832_), .ZN(new_n13009_));
  OAI21_X1   g12922(.A1(new_n13009_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n13010_));
  NOR2_X1    g12923(.A1(new_n11158_), .A2(new_n13010_), .ZN(new_n13011_));
  OAI22_X1   g12924(.A1(new_n10672_), .A2(new_n3040_), .B1(new_n8831_), .B2(new_n11159_), .ZN(new_n13012_));
  AOI21_X1   g12925(.A1(new_n13012_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13013_));
  AOI21_X1   g12926(.A1(new_n11153_), .A2(new_n11157_), .B(new_n13013_), .ZN(new_n13014_));
  NOR2_X1    g12927(.A1(new_n13014_), .A2(new_n13011_), .ZN(new_n13015_));
  NOR3_X1    g12928(.A1(new_n13007_), .A2(new_n13015_), .A3(new_n13008_), .ZN(new_n13016_));
  NOR2_X1    g12929(.A1(new_n13003_), .A2(new_n13005_), .ZN(new_n13017_));
  NOR2_X1    g12930(.A1(new_n13001_), .A2(new_n12998_), .ZN(new_n13018_));
  OAI21_X1   g12931(.A1(new_n13017_), .A2(new_n13018_), .B(new_n12999_), .ZN(new_n13019_));
  INV_X1     g12932(.I(new_n13008_), .ZN(new_n13020_));
  NAND3_X1   g12933(.A1(new_n13013_), .A2(new_n11157_), .A3(new_n11153_), .ZN(new_n13021_));
  NAND2_X1   g12934(.A1(new_n11158_), .A2(new_n13010_), .ZN(new_n13022_));
  NAND2_X1   g12935(.A1(new_n13022_), .A2(new_n13021_), .ZN(new_n13023_));
  AOI21_X1   g12936(.A1(new_n13019_), .A2(new_n13020_), .B(new_n13023_), .ZN(new_n13024_));
  NAND2_X1   g12937(.A1(new_n11003_), .A2(new_n8832_), .ZN(new_n13025_));
  NAND2_X1   g12938(.A1(new_n10745_), .A2(new_n2898_), .ZN(new_n13026_));
  AOI21_X1   g12939(.A1(new_n13025_), .A2(new_n13026_), .B(\a[5] ), .ZN(new_n13027_));
  NOR2_X1    g12940(.A1(new_n13027_), .A2(new_n3040_), .ZN(new_n13028_));
  NAND2_X1   g12941(.A1(new_n13028_), .A2(new_n11188_), .ZN(new_n13029_));
  INV_X1     g12942(.I(new_n13029_), .ZN(new_n13030_));
  NOR2_X1    g12943(.A1(new_n13028_), .A2(new_n11188_), .ZN(new_n13031_));
  NOR2_X1    g12944(.A1(new_n13030_), .A2(new_n13031_), .ZN(new_n13032_));
  NOR2_X1    g12945(.A1(new_n13032_), .A2(new_n12351_), .ZN(new_n13033_));
  NOR2_X1    g12946(.A1(new_n11009_), .A2(new_n2898_), .ZN(new_n13034_));
  AOI21_X1   g12947(.A1(new_n10783_), .A2(new_n10780_), .B(new_n3040_), .ZN(new_n13035_));
  NOR3_X1    g12948(.A1(new_n13034_), .A2(new_n11002_), .A3(new_n13035_), .ZN(new_n13036_));
  OAI22_X1   g12949(.A1(new_n10772_), .A2(new_n8830_), .B1(new_n3042_), .B2(new_n10755_), .ZN(new_n13037_));
  OAI21_X1   g12950(.A1(new_n3040_), .A2(new_n10762_), .B(new_n13037_), .ZN(new_n13038_));
  NOR2_X1    g12951(.A1(new_n13036_), .A2(new_n13038_), .ZN(new_n13039_));
  NOR2_X1    g12952(.A1(new_n13039_), .A2(\a[5] ), .ZN(new_n13040_));
  OR2_X2     g12953(.A1(new_n13036_), .A2(new_n13038_), .Z(new_n13041_));
  NOR2_X1    g12954(.A1(new_n13041_), .A2(new_n452_), .ZN(new_n13042_));
  NOR2_X1    g12955(.A1(new_n13042_), .A2(new_n13040_), .ZN(new_n13043_));
  NOR2_X1    g12956(.A1(new_n10772_), .A2(new_n3042_), .ZN(new_n13044_));
  OAI21_X1   g12957(.A1(new_n10755_), .A2(new_n3040_), .B(new_n452_), .ZN(new_n13045_));
  OAI21_X1   g12958(.A1(new_n13044_), .A2(new_n13045_), .B(new_n2898_), .ZN(new_n13046_));
  NOR2_X1    g12959(.A1(new_n13046_), .A2(new_n11017_), .ZN(new_n13047_));
  INV_X1     g12960(.I(new_n13047_), .ZN(new_n13048_));
  NAND2_X1   g12961(.A1(new_n13046_), .A2(new_n11017_), .ZN(new_n13049_));
  NAND2_X1   g12962(.A1(new_n13048_), .A2(new_n13049_), .ZN(new_n13050_));
  NOR2_X1    g12963(.A1(new_n10780_), .A2(new_n3419_), .ZN(new_n13051_));
  NOR2_X1    g12964(.A1(new_n13051_), .A2(new_n452_), .ZN(new_n13052_));
  INV_X1     g12965(.I(new_n13052_), .ZN(new_n13053_));
  NOR2_X1    g12966(.A1(new_n13050_), .A2(new_n13053_), .ZN(new_n13054_));
  NAND2_X1   g12967(.A1(new_n13043_), .A2(new_n13054_), .ZN(new_n13055_));
  NAND2_X1   g12968(.A1(new_n13032_), .A2(new_n12351_), .ZN(new_n13056_));
  AOI21_X1   g12969(.A1(new_n13055_), .A2(new_n13056_), .B(new_n13033_), .ZN(new_n13057_));
  NOR2_X1    g12970(.A1(new_n12350_), .A2(new_n12352_), .ZN(new_n13058_));
  AOI21_X1   g12971(.A1(new_n12349_), .A2(new_n12347_), .B(new_n12353_), .ZN(new_n13059_));
  NOR2_X1    g12972(.A1(new_n13058_), .A2(new_n13059_), .ZN(new_n13060_));
  INV_X1     g12973(.I(new_n13060_), .ZN(new_n13061_));
  OAI22_X1   g12974(.A1(new_n10725_), .A2(new_n3040_), .B1(new_n8831_), .B2(new_n11047_), .ZN(new_n13062_));
  AOI21_X1   g12975(.A1(new_n13062_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13063_));
  NAND3_X1   g12976(.A1(new_n11045_), .A2(new_n13063_), .A3(new_n11039_), .ZN(new_n13064_));
  INV_X1     g12977(.I(new_n13063_), .ZN(new_n13065_));
  NAND2_X1   g12978(.A1(new_n11046_), .A2(new_n13065_), .ZN(new_n13066_));
  NAND3_X1   g12979(.A1(new_n13061_), .A2(new_n13066_), .A3(new_n13064_), .ZN(new_n13067_));
  INV_X1     g12980(.I(new_n13067_), .ZN(new_n13068_));
  NAND2_X1   g12981(.A1(new_n13066_), .A2(new_n13064_), .ZN(new_n13069_));
  NAND2_X1   g12982(.A1(new_n13069_), .A2(new_n13060_), .ZN(new_n13070_));
  OAI21_X1   g12983(.A1(new_n13068_), .A2(new_n13057_), .B(new_n13070_), .ZN(new_n13071_));
  XOR2_X1    g12984(.A1(new_n12358_), .A2(new_n12354_), .Z(new_n13072_));
  AOI22_X1   g12985(.A1(new_n10794_), .A2(new_n2898_), .B1(new_n8832_), .B2(new_n11065_), .ZN(new_n13073_));
  OAI21_X1   g12986(.A1(new_n13073_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n13074_));
  XOR2_X1    g12987(.A1(new_n11064_), .A2(new_n13074_), .Z(new_n13075_));
  NAND2_X1   g12988(.A1(new_n13075_), .A2(new_n13072_), .ZN(new_n13076_));
  NOR2_X1    g12989(.A1(new_n13075_), .A2(new_n13072_), .ZN(new_n13077_));
  AOI21_X1   g12990(.A1(new_n13071_), .A2(new_n13076_), .B(new_n13077_), .ZN(new_n13078_));
  OAI21_X1   g12991(.A1(new_n12356_), .A2(new_n12359_), .B(new_n13004_), .ZN(new_n13079_));
  NAND2_X1   g12992(.A1(new_n13079_), .A2(new_n13001_), .ZN(new_n13080_));
  NOR2_X1    g12993(.A1(new_n10696_), .A2(new_n10725_), .ZN(new_n13081_));
  OAI22_X1   g12994(.A1(new_n13081_), .A2(new_n8831_), .B1(new_n3040_), .B2(new_n10792_), .ZN(new_n13082_));
  AOI21_X1   g12995(.A1(new_n13082_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13083_));
  INV_X1     g12996(.I(new_n13083_), .ZN(new_n13084_));
  NOR2_X1    g12997(.A1(new_n11333_), .A2(new_n13084_), .ZN(new_n13085_));
  NOR2_X1    g12998(.A1(new_n11140_), .A2(new_n13083_), .ZN(new_n13086_));
  NOR3_X1    g12999(.A1(new_n13080_), .A2(new_n13086_), .A3(new_n13085_), .ZN(new_n13087_));
  NOR2_X1    g13000(.A1(new_n13078_), .A2(new_n13087_), .ZN(new_n13088_));
  OAI21_X1   g13001(.A1(new_n13085_), .A2(new_n13086_), .B(new_n13080_), .ZN(new_n13089_));
  INV_X1     g13002(.I(new_n13089_), .ZN(new_n13090_));
  NOR4_X1    g13003(.A1(new_n13016_), .A2(new_n13088_), .A3(new_n13024_), .A4(new_n13090_), .ZN(new_n13091_));
  NAND2_X1   g13004(.A1(new_n13091_), .A2(new_n12997_), .ZN(new_n13092_));
  OAI21_X1   g13005(.A1(new_n13007_), .A2(new_n13008_), .B(new_n13015_), .ZN(new_n13093_));
  NAND2_X1   g13006(.A1(new_n10817_), .A2(new_n10691_), .ZN(new_n13094_));
  AOI22_X1   g13007(.A1(new_n13094_), .A2(new_n8832_), .B1(new_n10805_), .B2(new_n2898_), .ZN(new_n13095_));
  OAI21_X1   g13008(.A1(new_n13095_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n13096_));
  NOR3_X1    g13009(.A1(new_n11174_), .A2(new_n13096_), .A3(new_n11171_), .ZN(new_n13097_));
  INV_X1     g13010(.I(new_n13096_), .ZN(new_n13098_));
  NOR2_X1    g13011(.A1(new_n11175_), .A2(new_n13098_), .ZN(new_n13099_));
  NOR2_X1    g13012(.A1(new_n13099_), .A2(new_n13097_), .ZN(new_n13100_));
  NOR2_X1    g13013(.A1(new_n13100_), .A2(new_n13093_), .ZN(new_n13101_));
  OAI21_X1   g13014(.A1(new_n13091_), .A2(new_n12997_), .B(new_n13101_), .ZN(new_n13102_));
  NAND2_X1   g13015(.A1(new_n13102_), .A2(new_n13092_), .ZN(new_n13103_));
  INV_X1     g13016(.I(new_n12302_), .ZN(new_n13104_));
  NOR2_X1    g13017(.A1(new_n13104_), .A2(new_n12308_), .ZN(new_n13105_));
  INV_X1     g13018(.I(new_n13105_), .ZN(new_n13106_));
  NAND2_X1   g13019(.A1(new_n13104_), .A2(new_n12308_), .ZN(new_n13107_));
  AOI21_X1   g13020(.A1(new_n13107_), .A2(new_n13106_), .B(new_n12373_), .ZN(new_n13108_));
  NAND3_X1   g13021(.A1(new_n13104_), .A2(new_n12306_), .A3(new_n12307_), .ZN(new_n13109_));
  NAND2_X1   g13022(.A1(new_n12308_), .A2(new_n12302_), .ZN(new_n13110_));
  AOI21_X1   g13023(.A1(new_n13109_), .A2(new_n13110_), .B(new_n12374_), .ZN(new_n13111_));
  NOR2_X1    g13024(.A1(new_n13108_), .A2(new_n13111_), .ZN(new_n13112_));
  OAI22_X1   g13025(.A1(new_n10819_), .A2(new_n8831_), .B1(new_n11214_), .B2(new_n3040_), .ZN(new_n13113_));
  AOI21_X1   g13026(.A1(new_n13113_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13114_));
  XOR2_X1    g13027(.A1(new_n11224_), .A2(new_n13114_), .Z(new_n13115_));
  INV_X1     g13028(.I(new_n13115_), .ZN(new_n13116_));
  OAI21_X1   g13029(.A1(new_n13112_), .A2(new_n13116_), .B(new_n13103_), .ZN(new_n13117_));
  INV_X1     g13030(.I(new_n13112_), .ZN(new_n13118_));
  NOR2_X1    g13031(.A1(new_n13118_), .A2(new_n13115_), .ZN(new_n13119_));
  INV_X1     g13032(.I(new_n13119_), .ZN(new_n13120_));
  NAND2_X1   g13033(.A1(new_n13120_), .A2(new_n13117_), .ZN(new_n13121_));
  NAND2_X1   g13034(.A1(new_n13106_), .A2(new_n13107_), .ZN(new_n13122_));
  NAND3_X1   g13035(.A1(new_n12321_), .A2(new_n13122_), .A3(new_n13110_), .ZN(new_n13123_));
  NAND2_X1   g13036(.A1(new_n12308_), .A2(new_n12302_), .ZN(new_n13125_));
  AOI21_X1   g13037(.A1(new_n13123_), .A2(new_n13125_), .B(new_n12374_), .ZN(new_n13126_));
  NAND3_X1   g13038(.A1(new_n13123_), .A2(new_n12374_), .A3(new_n13125_), .ZN(new_n13127_));
  INV_X1     g13039(.I(new_n13127_), .ZN(new_n13128_));
  AOI22_X1   g13040(.A1(new_n10828_), .A2(new_n2898_), .B1(new_n8832_), .B2(new_n12145_), .ZN(new_n13129_));
  NOR2_X1    g13041(.A1(new_n13129_), .A2(\a[5] ), .ZN(new_n13130_));
  NOR3_X1    g13042(.A1(new_n11246_), .A2(new_n3040_), .A3(new_n13130_), .ZN(new_n13131_));
  NAND2_X1   g13043(.A1(new_n11243_), .A2(new_n11214_), .ZN(new_n13132_));
  NAND2_X1   g13044(.A1(new_n11239_), .A2(new_n10652_), .ZN(new_n13133_));
  AOI21_X1   g13045(.A1(new_n13132_), .A2(new_n13133_), .B(new_n10828_), .ZN(new_n13134_));
  NOR2_X1    g13046(.A1(new_n13134_), .A2(new_n11237_), .ZN(new_n13135_));
  NOR2_X1    g13047(.A1(new_n13130_), .A2(new_n3040_), .ZN(new_n13136_));
  NOR2_X1    g13048(.A1(new_n13136_), .A2(new_n13135_), .ZN(new_n13137_));
  NOR2_X1    g13049(.A1(new_n13131_), .A2(new_n13137_), .ZN(new_n13138_));
  OAI21_X1   g13050(.A1(new_n13128_), .A2(new_n13126_), .B(new_n13138_), .ZN(new_n13139_));
  INV_X1     g13051(.I(new_n13126_), .ZN(new_n13140_));
  OR2_X2     g13052(.A1(new_n13131_), .A2(new_n13137_), .Z(new_n13141_));
  NAND3_X1   g13053(.A1(new_n13140_), .A2(new_n13141_), .A3(new_n13127_), .ZN(new_n13142_));
  INV_X1     g13054(.I(new_n13142_), .ZN(new_n13143_));
  AOI21_X1   g13055(.A1(new_n13121_), .A2(new_n13139_), .B(new_n13143_), .ZN(new_n13144_));
  AOI21_X1   g13056(.A1(new_n12295_), .A2(new_n12290_), .B(new_n12293_), .ZN(new_n13145_));
  NOR3_X1    g13057(.A1(new_n12291_), .A2(new_n11505_), .A3(new_n12289_), .ZN(new_n13146_));
  NOR2_X1    g13058(.A1(new_n13146_), .A2(new_n13145_), .ZN(new_n13147_));
  NOR3_X1    g13059(.A1(new_n13147_), .A2(new_n12376_), .A3(new_n12380_), .ZN(new_n13148_));
  INV_X1     g13060(.I(new_n12376_), .ZN(new_n13149_));
  AOI21_X1   g13061(.A1(new_n12292_), .A2(new_n12296_), .B(new_n12380_), .ZN(new_n13150_));
  NOR2_X1    g13062(.A1(new_n13150_), .A2(new_n13149_), .ZN(new_n13151_));
  OAI21_X1   g13063(.A1(new_n13148_), .A2(new_n13151_), .B(new_n12320_), .ZN(new_n13152_));
  INV_X1     g13064(.I(new_n12320_), .ZN(new_n13153_));
  NAND2_X1   g13065(.A1(new_n13150_), .A2(new_n13149_), .ZN(new_n13154_));
  OAI21_X1   g13066(.A1(new_n13147_), .A2(new_n12380_), .B(new_n12376_), .ZN(new_n13155_));
  NAND3_X1   g13067(.A1(new_n13155_), .A2(new_n13154_), .A3(new_n13153_), .ZN(new_n13156_));
  AOI22_X1   g13068(.A1(new_n10638_), .A2(new_n2898_), .B1(new_n8832_), .B2(new_n11269_), .ZN(new_n13157_));
  NOR2_X1    g13069(.A1(new_n13157_), .A2(\a[5] ), .ZN(new_n13158_));
  NOR2_X1    g13070(.A1(new_n13158_), .A2(new_n3040_), .ZN(new_n13159_));
  XNOR2_X1   g13071(.A1(new_n11268_), .A2(new_n13159_), .ZN(new_n13160_));
  NAND3_X1   g13072(.A1(new_n13152_), .A2(new_n13156_), .A3(new_n13160_), .ZN(new_n13161_));
  AOI21_X1   g13073(.A1(new_n13155_), .A2(new_n13154_), .B(new_n13153_), .ZN(new_n13162_));
  NOR3_X1    g13074(.A1(new_n13148_), .A2(new_n13151_), .A3(new_n12320_), .ZN(new_n13163_));
  INV_X1     g13075(.I(new_n13160_), .ZN(new_n13164_));
  OAI21_X1   g13076(.A1(new_n13162_), .A2(new_n13163_), .B(new_n13164_), .ZN(new_n13165_));
  NAND3_X1   g13077(.A1(new_n13165_), .A2(new_n13161_), .A3(new_n13144_), .ZN(new_n13166_));
  NOR2_X1    g13078(.A1(new_n13166_), .A2(new_n12980_), .ZN(new_n13167_));
  NOR3_X1    g13079(.A1(new_n13162_), .A2(new_n13163_), .A3(new_n13164_), .ZN(new_n13168_));
  OAI22_X1   g13080(.A1(new_n11386_), .A2(new_n8831_), .B1(new_n3040_), .B2(new_n10633_), .ZN(new_n13169_));
  AOI21_X1   g13081(.A1(new_n13169_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13170_));
  XOR2_X1    g13082(.A1(new_n11987_), .A2(new_n13170_), .Z(new_n13171_));
  NAND2_X1   g13083(.A1(new_n13168_), .A2(new_n13171_), .ZN(new_n13172_));
  AOI21_X1   g13084(.A1(new_n13166_), .A2(new_n12980_), .B(new_n13172_), .ZN(new_n13173_));
  NOR2_X1    g13085(.A1(new_n13173_), .A2(new_n13167_), .ZN(new_n13174_));
  NAND2_X1   g13086(.A1(new_n12971_), .A2(new_n12972_), .ZN(new_n13175_));
  XOR2_X1    g13087(.A1(new_n12399_), .A2(new_n12404_), .Z(new_n13176_));
  AOI21_X1   g13088(.A1(new_n13175_), .A2(new_n12394_), .B(new_n13176_), .ZN(new_n13177_));
  NAND2_X1   g13089(.A1(new_n13175_), .A2(new_n12394_), .ZN(new_n13178_));
  NOR2_X1    g13090(.A1(new_n12399_), .A2(new_n12405_), .ZN(new_n13179_));
  NOR2_X1    g13091(.A1(new_n12409_), .A2(new_n13179_), .ZN(new_n13180_));
  NOR2_X1    g13092(.A1(new_n13180_), .A2(new_n13178_), .ZN(new_n13181_));
  NOR2_X1    g13093(.A1(new_n13177_), .A2(new_n13181_), .ZN(new_n13182_));
  NAND2_X1   g13094(.A1(new_n11446_), .A2(new_n8832_), .ZN(new_n13183_));
  OAI21_X1   g13095(.A1(new_n10631_), .A2(new_n3040_), .B(new_n13183_), .ZN(new_n13184_));
  AOI21_X1   g13096(.A1(new_n13184_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13185_));
  XOR2_X1    g13097(.A1(new_n11445_), .A2(new_n13185_), .Z(new_n13186_));
  INV_X1     g13098(.I(new_n13186_), .ZN(new_n13187_));
  NOR2_X1    g13099(.A1(new_n13182_), .A2(new_n13187_), .ZN(new_n13188_));
  NOR2_X1    g13100(.A1(new_n13188_), .A2(new_n13174_), .ZN(new_n13189_));
  NOR3_X1    g13101(.A1(new_n13177_), .A2(new_n13181_), .A3(new_n13186_), .ZN(new_n13190_));
  NOR2_X1    g13102(.A1(new_n13189_), .A2(new_n13190_), .ZN(new_n13191_));
  NOR2_X1    g13103(.A1(new_n12407_), .A2(new_n12409_), .ZN(new_n13192_));
  NAND2_X1   g13104(.A1(new_n13192_), .A2(new_n12419_), .ZN(new_n13193_));
  NOR2_X1    g13105(.A1(new_n13192_), .A2(new_n12419_), .ZN(new_n13194_));
  INV_X1     g13106(.I(new_n13194_), .ZN(new_n13195_));
  AOI22_X1   g13107(.A1(new_n2898_), .A2(new_n10843_), .B1(new_n11608_), .B2(new_n8832_), .ZN(new_n13196_));
  OAI21_X1   g13108(.A1(new_n13196_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n13197_));
  XOR2_X1    g13109(.A1(new_n11607_), .A2(new_n13197_), .Z(new_n13198_));
  INV_X1     g13110(.I(new_n13198_), .ZN(new_n13199_));
  NAND3_X1   g13111(.A1(new_n13195_), .A2(new_n13199_), .A3(new_n13193_), .ZN(new_n13200_));
  INV_X1     g13112(.I(new_n13193_), .ZN(new_n13201_));
  OAI21_X1   g13113(.A1(new_n13201_), .A2(new_n13194_), .B(new_n13198_), .ZN(new_n13202_));
  NAND2_X1   g13114(.A1(new_n12283_), .A2(new_n12425_), .ZN(new_n13203_));
  NOR2_X1    g13115(.A1(new_n13203_), .A2(new_n12420_), .ZN(new_n13204_));
  AOI21_X1   g13116(.A1(new_n12283_), .A2(new_n12425_), .B(new_n12438_), .ZN(new_n13205_));
  OAI21_X1   g13117(.A1(new_n13204_), .A2(new_n13205_), .B(new_n12415_), .ZN(new_n13206_));
  NAND3_X1   g13118(.A1(new_n12438_), .A2(new_n12283_), .A3(new_n12425_), .ZN(new_n13207_));
  NAND2_X1   g13119(.A1(new_n13203_), .A2(new_n12420_), .ZN(new_n13208_));
  NAND3_X1   g13120(.A1(new_n13208_), .A2(new_n13207_), .A3(new_n12422_), .ZN(new_n13209_));
  INV_X1     g13121(.I(new_n11631_), .ZN(new_n13210_));
  AOI22_X1   g13122(.A1(new_n11632_), .A2(new_n8832_), .B1(new_n10857_), .B2(new_n2898_), .ZN(new_n13211_));
  OAI21_X1   g13123(.A1(new_n13211_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n13212_));
  NOR2_X1    g13124(.A1(new_n13210_), .A2(new_n13212_), .ZN(new_n13213_));
  INV_X1     g13125(.I(new_n13212_), .ZN(new_n13214_));
  NOR2_X1    g13126(.A1(new_n11631_), .A2(new_n13214_), .ZN(new_n13215_));
  NOR2_X1    g13127(.A1(new_n13213_), .A2(new_n13215_), .ZN(new_n13216_));
  INV_X1     g13128(.I(new_n13216_), .ZN(new_n13217_));
  NAND3_X1   g13129(.A1(new_n13217_), .A2(new_n13206_), .A3(new_n13209_), .ZN(new_n13218_));
  INV_X1     g13130(.I(new_n13218_), .ZN(new_n13219_));
  AOI21_X1   g13131(.A1(new_n13206_), .A2(new_n13209_), .B(new_n13217_), .ZN(new_n13220_));
  AOI21_X1   g13132(.A1(new_n13200_), .A2(new_n13202_), .B(new_n13191_), .ZN(new_n13222_));
  NOR2_X1    g13133(.A1(new_n12970_), .A2(new_n13222_), .ZN(new_n13223_));
  INV_X1     g13134(.I(new_n11647_), .ZN(new_n13224_));
  NAND2_X1   g13135(.A1(new_n13224_), .A2(new_n11645_), .ZN(new_n13225_));
  OAI22_X1   g13136(.A1(new_n10870_), .A2(new_n3040_), .B1(new_n8831_), .B2(new_n10861_), .ZN(new_n13226_));
  AOI21_X1   g13137(.A1(new_n13226_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13227_));
  XOR2_X1    g13138(.A1(new_n13225_), .A2(new_n13227_), .Z(new_n13228_));
  NAND2_X1   g13139(.A1(new_n13220_), .A2(new_n13228_), .ZN(new_n13229_));
  NOR2_X1    g13140(.A1(new_n13223_), .A2(new_n13229_), .ZN(new_n13230_));
  AOI21_X1   g13141(.A1(new_n12970_), .A2(new_n13222_), .B(new_n13230_), .ZN(new_n13231_));
  AOI21_X1   g13142(.A1(new_n12467_), .A2(new_n12462_), .B(new_n12449_), .ZN(new_n13232_));
  NAND2_X1   g13143(.A1(new_n12465_), .A2(new_n12461_), .ZN(new_n13233_));
  NAND2_X1   g13144(.A1(new_n12458_), .A2(new_n12466_), .ZN(new_n13234_));
  AOI21_X1   g13145(.A1(new_n13233_), .A2(new_n13234_), .B(new_n12450_), .ZN(new_n13235_));
  AOI22_X1   g13146(.A1(new_n11724_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n10875_), .ZN(new_n13236_));
  OAI21_X1   g13147(.A1(new_n13236_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n13237_));
  XOR2_X1    g13148(.A1(new_n11722_), .A2(new_n13237_), .Z(new_n13238_));
  NOR3_X1    g13149(.A1(new_n13235_), .A2(new_n13232_), .A3(new_n13238_), .ZN(new_n13239_));
  OAI21_X1   g13150(.A1(new_n13235_), .A2(new_n13232_), .B(new_n13238_), .ZN(new_n13240_));
  OAI21_X1   g13151(.A1(new_n13231_), .A2(new_n13239_), .B(new_n13240_), .ZN(new_n13241_));
  INV_X1     g13152(.I(new_n11803_), .ZN(new_n13242_));
  AOI22_X1   g13153(.A1(new_n13242_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n10882_), .ZN(new_n13243_));
  OAI21_X1   g13154(.A1(new_n13243_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n13244_));
  NOR2_X1    g13155(.A1(new_n11802_), .A2(new_n13244_), .ZN(new_n13245_));
  AND2_X2    g13156(.A1(new_n11802_), .A2(new_n13244_), .Z(new_n13246_));
  NOR2_X1    g13157(.A1(new_n13246_), .A2(new_n13245_), .ZN(new_n13247_));
  INV_X1     g13158(.I(new_n13247_), .ZN(new_n13248_));
  NAND2_X1   g13159(.A1(new_n13241_), .A2(new_n13248_), .ZN(new_n13249_));
  INV_X1     g13160(.I(new_n13249_), .ZN(new_n13250_));
  INV_X1     g13161(.I(new_n13241_), .ZN(new_n13251_));
  NAND2_X1   g13162(.A1(new_n12463_), .A2(new_n12467_), .ZN(new_n13252_));
  NAND2_X1   g13163(.A1(new_n12482_), .A2(new_n12480_), .ZN(new_n13253_));
  XNOR2_X1   g13164(.A1(new_n13252_), .A2(new_n13253_), .ZN(new_n13254_));
  AOI21_X1   g13165(.A1(new_n13251_), .A2(new_n13247_), .B(new_n13254_), .ZN(new_n13255_));
  INV_X1     g13166(.I(new_n12482_), .ZN(new_n13256_));
  INV_X1     g13167(.I(new_n12488_), .ZN(new_n13257_));
  NAND3_X1   g13168(.A1(new_n12271_), .A2(new_n12483_), .A3(new_n13257_), .ZN(new_n13258_));
  AOI21_X1   g13169(.A1(new_n12268_), .A2(new_n12269_), .B(new_n12005_), .ZN(new_n13259_));
  NOR3_X1    g13170(.A1(new_n12266_), .A2(new_n12263_), .A3(new_n12004_), .ZN(new_n13260_));
  OAI21_X1   g13171(.A1(new_n13260_), .A2(new_n13259_), .B(new_n13257_), .ZN(new_n13261_));
  NAND2_X1   g13172(.A1(new_n13261_), .A2(new_n12484_), .ZN(new_n13262_));
  AOI21_X1   g13173(.A1(new_n13262_), .A2(new_n13258_), .B(new_n13256_), .ZN(new_n13263_));
  NOR2_X1    g13174(.A1(new_n13261_), .A2(new_n12484_), .ZN(new_n13264_));
  AOI21_X1   g13175(.A1(new_n12271_), .A2(new_n13257_), .B(new_n12483_), .ZN(new_n13265_));
  NOR3_X1    g13176(.A1(new_n13264_), .A2(new_n13265_), .A3(new_n12482_), .ZN(new_n13266_));
  OAI22_X1   g13177(.A1(new_n10619_), .A2(new_n3040_), .B1(new_n8831_), .B2(new_n10885_), .ZN(new_n13267_));
  AOI21_X1   g13178(.A1(new_n13267_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13268_));
  XOR2_X1    g13179(.A1(new_n12074_), .A2(new_n13268_), .Z(new_n13269_));
  OAI21_X1   g13180(.A1(new_n13266_), .A2(new_n13263_), .B(new_n13269_), .ZN(new_n13270_));
  OAI21_X1   g13181(.A1(new_n13250_), .A2(new_n13255_), .B(new_n13270_), .ZN(new_n13271_));
  OAI21_X1   g13182(.A1(new_n13264_), .A2(new_n13265_), .B(new_n12482_), .ZN(new_n13272_));
  NAND3_X1   g13183(.A1(new_n13262_), .A2(new_n13258_), .A3(new_n13256_), .ZN(new_n13273_));
  INV_X1     g13184(.I(new_n13269_), .ZN(new_n13274_));
  NAND3_X1   g13185(.A1(new_n13272_), .A2(new_n13273_), .A3(new_n13274_), .ZN(new_n13275_));
  NAND2_X1   g13186(.A1(new_n13271_), .A2(new_n13275_), .ZN(new_n13276_));
  OAI21_X1   g13187(.A1(new_n12494_), .A2(new_n12498_), .B(new_n12501_), .ZN(new_n13277_));
  NAND2_X1   g13188(.A1(new_n12506_), .A2(new_n12502_), .ZN(new_n13278_));
  AOI22_X1   g13189(.A1(new_n13278_), .A2(new_n13277_), .B1(new_n12485_), .B2(new_n12490_), .ZN(new_n13279_));
  NOR2_X1    g13190(.A1(new_n12507_), .A2(new_n12503_), .ZN(new_n13280_));
  NOR2_X1    g13191(.A1(new_n13280_), .A2(new_n12491_), .ZN(new_n13281_));
  OAI22_X1   g13192(.A1(new_n12091_), .A2(new_n8831_), .B1(new_n3040_), .B2(new_n10611_), .ZN(new_n13282_));
  AOI21_X1   g13193(.A1(new_n13282_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13283_));
  XOR2_X1    g13194(.A1(new_n12090_), .A2(new_n13283_), .Z(new_n13284_));
  NOR3_X1    g13195(.A1(new_n13281_), .A2(new_n13279_), .A3(new_n13284_), .ZN(new_n13285_));
  OAI21_X1   g13196(.A1(new_n13281_), .A2(new_n13279_), .B(new_n13284_), .ZN(new_n13286_));
  INV_X1     g13197(.I(new_n13286_), .ZN(new_n13287_));
  AOI22_X1   g13198(.A1(new_n10986_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n10897_), .ZN(new_n13288_));
  OAI21_X1   g13199(.A1(new_n13288_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n13289_));
  NOR2_X1    g13200(.A1(new_n10984_), .A2(new_n13289_), .ZN(new_n13290_));
  NOR2_X1    g13201(.A1(new_n10889_), .A2(new_n10982_), .ZN(new_n13291_));
  INV_X1     g13202(.I(new_n10983_), .ZN(new_n13292_));
  NOR2_X1    g13203(.A1(new_n13292_), .A2(new_n13291_), .ZN(new_n13293_));
  INV_X1     g13204(.I(new_n13289_), .ZN(new_n13294_));
  NOR2_X1    g13205(.A1(new_n13293_), .A2(new_n13294_), .ZN(new_n13295_));
  NOR2_X1    g13206(.A1(new_n13295_), .A2(new_n13290_), .ZN(new_n13296_));
  INV_X1     g13207(.I(new_n13296_), .ZN(new_n13297_));
  NOR2_X1    g13208(.A1(new_n12951_), .A2(new_n13297_), .ZN(new_n13298_));
  NOR2_X1    g13209(.A1(new_n12521_), .A2(new_n13296_), .ZN(new_n13299_));
  OAI21_X1   g13210(.A1(new_n13299_), .A2(new_n13298_), .B(new_n12948_), .ZN(new_n13300_));
  INV_X1     g13211(.I(new_n13300_), .ZN(new_n13301_));
  NAND2_X1   g13212(.A1(new_n12521_), .A2(new_n13297_), .ZN(new_n13302_));
  NAND2_X1   g13213(.A1(new_n12951_), .A2(new_n13296_), .ZN(new_n13303_));
  AOI21_X1   g13214(.A1(new_n13302_), .A2(new_n13303_), .B(new_n12948_), .ZN(new_n13304_));
  OAI21_X1   g13215(.A1(new_n13287_), .A2(new_n13285_), .B(new_n13276_), .ZN(new_n13306_));
  NOR2_X1    g13216(.A1(new_n12958_), .A2(new_n13306_), .ZN(new_n13307_));
  XOR2_X1    g13217(.A1(new_n12948_), .A2(new_n12951_), .Z(new_n13308_));
  OAI22_X1   g13218(.A1(new_n10606_), .A2(new_n3040_), .B1(new_n8831_), .B2(new_n10901_), .ZN(new_n13309_));
  AOI21_X1   g13219(.A1(new_n13309_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13310_));
  XOR2_X1    g13220(.A1(new_n12211_), .A2(new_n13310_), .Z(new_n13311_));
  INV_X1     g13221(.I(new_n13311_), .ZN(new_n13312_));
  NAND3_X1   g13222(.A1(new_n13308_), .A2(new_n13296_), .A3(new_n13312_), .ZN(new_n13313_));
  AOI21_X1   g13223(.A1(new_n12958_), .A2(new_n13306_), .B(new_n13313_), .ZN(new_n13314_));
  AOI22_X1   g13224(.A1(new_n12578_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n10600_), .ZN(new_n13315_));
  OAI21_X1   g13225(.A1(new_n13315_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n13316_));
  XNOR2_X1   g13226(.A1(new_n12576_), .A2(new_n13316_), .ZN(new_n13317_));
  INV_X1     g13227(.I(new_n13317_), .ZN(new_n13318_));
  NOR3_X1    g13228(.A1(new_n13314_), .A2(new_n13307_), .A3(new_n13318_), .ZN(new_n13319_));
  OAI21_X1   g13229(.A1(new_n13314_), .A2(new_n13307_), .B(new_n13318_), .ZN(new_n13320_));
  OAI21_X1   g13230(.A1(new_n12942_), .A2(new_n13319_), .B(new_n13320_), .ZN(new_n13321_));
  OAI22_X1   g13231(.A1(new_n12601_), .A2(new_n8831_), .B1(new_n3040_), .B2(new_n10595_), .ZN(new_n13322_));
  AOI21_X1   g13232(.A1(new_n13322_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13323_));
  XOR2_X1    g13233(.A1(new_n12600_), .A2(new_n13323_), .Z(new_n13324_));
  INV_X1     g13234(.I(new_n13324_), .ZN(new_n13325_));
  OAI22_X1   g13235(.A1(new_n13321_), .A2(new_n13325_), .B1(new_n12555_), .B2(new_n12933_), .ZN(new_n13326_));
  NAND2_X1   g13236(.A1(new_n13321_), .A2(new_n13325_), .ZN(new_n13327_));
  OAI22_X1   g13237(.A1(new_n10589_), .A2(new_n3040_), .B1(new_n12623_), .B2(new_n8831_), .ZN(new_n13328_));
  AOI21_X1   g13238(.A1(new_n13328_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13329_));
  XOR2_X1    g13239(.A1(new_n12622_), .A2(new_n13329_), .Z(new_n13330_));
  AOI21_X1   g13240(.A1(new_n13326_), .A2(new_n13327_), .B(new_n13330_), .ZN(new_n13331_));
  INV_X1     g13241(.I(new_n13331_), .ZN(new_n13332_));
  INV_X1     g13242(.I(new_n12559_), .ZN(new_n13333_));
  INV_X1     g13243(.I(new_n12562_), .ZN(new_n13334_));
  NAND2_X1   g13244(.A1(new_n12241_), .A2(new_n13334_), .ZN(new_n13335_));
  OR2_X2     g13245(.A1(new_n12555_), .A2(new_n13335_), .Z(new_n13336_));
  NAND2_X1   g13246(.A1(new_n13335_), .A2(new_n12555_), .ZN(new_n13337_));
  AOI21_X1   g13247(.A1(new_n13336_), .A2(new_n13337_), .B(new_n13333_), .ZN(new_n13338_));
  NAND3_X1   g13248(.A1(new_n13336_), .A2(new_n13333_), .A3(new_n13337_), .ZN(new_n13339_));
  INV_X1     g13249(.I(new_n13339_), .ZN(new_n13340_));
  NOR2_X1    g13250(.A1(new_n13340_), .A2(new_n13338_), .ZN(new_n13341_));
  NAND3_X1   g13251(.A1(new_n13326_), .A2(new_n13327_), .A3(new_n13330_), .ZN(new_n13342_));
  NAND2_X1   g13252(.A1(new_n13342_), .A2(new_n13341_), .ZN(new_n13343_));
  NAND2_X1   g13253(.A1(new_n13343_), .A2(new_n13332_), .ZN(new_n13344_));
  OAI21_X1   g13254(.A1(new_n12921_), .A2(new_n12918_), .B(new_n12924_), .ZN(new_n13345_));
  AOI22_X1   g13255(.A1(new_n12891_), .A2(new_n8832_), .B1(new_n10924_), .B2(new_n2898_), .ZN(new_n13346_));
  OAI21_X1   g13256(.A1(new_n13346_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n13347_));
  XNOR2_X1   g13257(.A1(new_n12889_), .A2(new_n13347_), .ZN(new_n13348_));
  NAND3_X1   g13258(.A1(new_n12606_), .A2(new_n12607_), .A3(new_n12608_), .ZN(new_n13349_));
  NAND3_X1   g13259(.A1(new_n13349_), .A2(new_n12582_), .A3(new_n12613_), .ZN(new_n13350_));
  NAND3_X1   g13260(.A1(new_n13350_), .A2(new_n12919_), .A3(new_n12920_), .ZN(new_n13351_));
  INV_X1     g13261(.I(new_n12582_), .ZN(new_n13352_));
  NOR3_X1    g13262(.A1(new_n12609_), .A2(new_n12605_), .A3(new_n13352_), .ZN(new_n13353_));
  OAI21_X1   g13263(.A1(new_n13353_), .A2(new_n12917_), .B(new_n12916_), .ZN(new_n13354_));
  NAND3_X1   g13264(.A1(new_n13354_), .A2(new_n13351_), .A3(new_n13348_), .ZN(new_n13355_));
  INV_X1     g13265(.I(new_n13348_), .ZN(new_n13356_));
  NOR3_X1    g13266(.A1(new_n13353_), .A2(new_n12916_), .A3(new_n12917_), .ZN(new_n13357_));
  AOI21_X1   g13267(.A1(new_n13350_), .A2(new_n12920_), .B(new_n12919_), .ZN(new_n13358_));
  OAI21_X1   g13268(.A1(new_n13358_), .A2(new_n13357_), .B(new_n13356_), .ZN(new_n13359_));
  AOI21_X1   g13269(.A1(new_n13359_), .A2(new_n13355_), .B(new_n13345_), .ZN(new_n13360_));
  OAI21_X1   g13270(.A1(new_n13344_), .A2(new_n13360_), .B(new_n12930_), .ZN(new_n13361_));
  AOI21_X1   g13271(.A1(new_n13354_), .A2(new_n13351_), .B(new_n13356_), .ZN(new_n13362_));
  INV_X1     g13272(.I(new_n13362_), .ZN(new_n13363_));
  AOI21_X1   g13273(.A1(new_n12226_), .A2(new_n12230_), .B(new_n12626_), .ZN(new_n13364_));
  INV_X1     g13274(.I(new_n13364_), .ZN(new_n13365_));
  NOR2_X1    g13275(.A1(new_n13365_), .A2(new_n12611_), .ZN(new_n13366_));
  INV_X1     g13276(.I(new_n13366_), .ZN(new_n13367_));
  NAND2_X1   g13277(.A1(new_n13365_), .A2(new_n12611_), .ZN(new_n13368_));
  AOI21_X1   g13278(.A1(new_n13367_), .A2(new_n13368_), .B(new_n12609_), .ZN(new_n13369_));
  INV_X1     g13279(.I(new_n13368_), .ZN(new_n13370_));
  NOR3_X1    g13280(.A1(new_n13370_), .A2(new_n12613_), .A3(new_n13366_), .ZN(new_n13371_));
  NOR2_X1    g13281(.A1(new_n10583_), .A2(new_n10924_), .ZN(new_n13372_));
  NOR2_X1    g13282(.A1(new_n10584_), .A2(new_n10923_), .ZN(new_n13373_));
  OAI21_X1   g13283(.A1(new_n13373_), .A2(new_n13372_), .B(new_n12886_), .ZN(new_n13374_));
  NOR2_X1    g13284(.A1(new_n10916_), .A2(new_n13374_), .ZN(new_n13375_));
  INV_X1     g13285(.I(new_n13375_), .ZN(new_n13376_));
  NAND2_X1   g13286(.A1(new_n10916_), .A2(new_n13374_), .ZN(new_n13377_));
  NAND2_X1   g13287(.A1(new_n13376_), .A2(new_n13377_), .ZN(new_n13378_));
  OAI22_X1   g13288(.A1(new_n10583_), .A2(new_n3040_), .B1(new_n8831_), .B2(new_n10928_), .ZN(new_n13379_));
  AOI21_X1   g13289(.A1(new_n13379_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13380_));
  XNOR2_X1   g13290(.A1(new_n13378_), .A2(new_n13380_), .ZN(new_n13381_));
  INV_X1     g13291(.I(new_n13381_), .ZN(new_n13382_));
  OR3_X2     g13292(.A1(new_n13369_), .A2(new_n13371_), .A3(new_n13382_), .Z(new_n13383_));
  NAND3_X1   g13293(.A1(new_n13361_), .A2(new_n13383_), .A3(new_n13363_), .ZN(new_n13384_));
  OAI21_X1   g13294(.A1(new_n13369_), .A2(new_n13371_), .B(new_n13382_), .ZN(new_n13385_));
  NOR3_X1    g13295(.A1(new_n12629_), .A2(new_n12774_), .A3(new_n12775_), .ZN(new_n13386_));
  INV_X1     g13296(.I(new_n13386_), .ZN(new_n13387_));
  OAI21_X1   g13297(.A1(new_n12774_), .A2(new_n12775_), .B(new_n12629_), .ZN(new_n13388_));
  NAND3_X1   g13298(.A1(new_n10927_), .A2(new_n10929_), .A3(new_n10583_), .ZN(new_n13389_));
  OAI21_X1   g13299(.A1(new_n10916_), .A2(new_n10926_), .B(new_n10584_), .ZN(new_n13390_));
  AOI21_X1   g13300(.A1(new_n13389_), .A2(new_n13390_), .B(new_n10938_), .ZN(new_n13391_));
  INV_X1     g13301(.I(new_n10930_), .ZN(new_n13392_));
  AOI21_X1   g13302(.A1(new_n13392_), .A2(new_n10940_), .B(new_n10937_), .ZN(new_n13393_));
  NOR2_X1    g13303(.A1(new_n13393_), .A2(new_n13391_), .ZN(new_n13394_));
  NOR2_X1    g13304(.A1(new_n10583_), .A2(new_n10923_), .ZN(new_n13395_));
  OAI22_X1   g13305(.A1(new_n13395_), .A2(new_n8831_), .B1(new_n3040_), .B2(new_n10938_), .ZN(new_n13396_));
  AOI21_X1   g13306(.A1(new_n13396_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13397_));
  XOR2_X1    g13307(.A1(new_n13394_), .A2(new_n13397_), .Z(new_n13398_));
  NAND3_X1   g13308(.A1(new_n13387_), .A2(new_n13388_), .A3(new_n13398_), .ZN(new_n13399_));
  NOR2_X1    g13309(.A1(new_n12902_), .A2(new_n12776_), .ZN(new_n13400_));
  INV_X1     g13310(.I(new_n13398_), .ZN(new_n13401_));
  OAI21_X1   g13311(.A1(new_n13400_), .A2(new_n13386_), .B(new_n13401_), .ZN(new_n13402_));
  OAI21_X1   g13312(.A1(new_n12904_), .A2(new_n12901_), .B(new_n12913_), .ZN(new_n13403_));
  AOI22_X1   g13313(.A1(new_n13384_), .A2(new_n13385_), .B1(new_n13399_), .B2(new_n13402_), .ZN(new_n13405_));
  NOR2_X1    g13314(.A1(new_n12756_), .A2(new_n12759_), .ZN(new_n13406_));
  NOR2_X1    g13315(.A1(new_n12636_), .A2(new_n12751_), .ZN(new_n13407_));
  OAI21_X1   g13316(.A1(new_n13406_), .A2(new_n13407_), .B(new_n12771_), .ZN(new_n13408_));
  AOI22_X1   g13317(.A1(new_n12628_), .A2(new_n12612_), .B1(new_n12773_), .B2(new_n13408_), .ZN(new_n13410_));
  INV_X1     g13318(.I(new_n13410_), .ZN(new_n13411_));
  AOI22_X1   g13319(.A1(new_n12755_), .A2(new_n12753_), .B1(new_n12750_), .B2(new_n12745_), .ZN(new_n13413_));
  NAND4_X1   g13320(.A1(new_n12779_), .A2(new_n12733_), .A3(new_n12862_), .A4(new_n12865_), .ZN(new_n13414_));
  AOI22_X1   g13321(.A1(new_n12852_), .A2(new_n12851_), .B1(new_n12724_), .B2(new_n12725_), .ZN(new_n13416_));
  NAND3_X1   g13322(.A1(new_n12820_), .A2(new_n12788_), .A3(new_n12815_), .ZN(new_n13417_));
  AOI21_X1   g13323(.A1(new_n12834_), .A2(new_n13417_), .B(new_n12825_), .ZN(new_n13418_));
  AOI22_X1   g13324(.A1(new_n10630_), .A2(new_n247_), .B1(new_n5783_), .B2(new_n11446_), .ZN(new_n13419_));
  NOR2_X1    g13325(.A1(new_n13419_), .A2(\a[23] ), .ZN(new_n13420_));
  NOR2_X1    g13326(.A1(new_n13420_), .A2(new_n1239_), .ZN(new_n13421_));
  XOR2_X1    g13327(.A1(new_n11445_), .A2(new_n13421_), .Z(new_n13422_));
  AND2_X2    g13328(.A1(new_n12806_), .A2(new_n12811_), .Z(new_n13423_));
  AOI21_X1   g13329(.A1(new_n12812_), .A2(new_n12673_), .B(new_n12678_), .ZN(new_n13424_));
  OAI21_X1   g13330(.A1(new_n12812_), .A2(new_n12673_), .B(new_n12655_), .ZN(new_n13425_));
  NOR2_X1    g13331(.A1(new_n13424_), .A2(new_n13425_), .ZN(new_n13426_));
  AOI21_X1   g13332(.A1(new_n12789_), .A2(new_n12802_), .B(new_n12804_), .ZN(new_n13427_));
  OAI22_X1   g13333(.A1(new_n10792_), .A2(new_n4527_), .B1(new_n10696_), .B2(new_n4529_), .ZN(new_n13428_));
  OAI21_X1   g13334(.A1(new_n10672_), .A2(new_n79_), .B(new_n13428_), .ZN(new_n13429_));
  AOI21_X1   g13335(.A1(new_n13429_), .A2(new_n72_), .B(new_n79_), .ZN(new_n13430_));
  XNOR2_X1   g13336(.A1(new_n11158_), .A2(new_n13430_), .ZN(new_n13431_));
  NOR3_X1    g13337(.A1(new_n12795_), .A2(new_n11188_), .A3(new_n12798_), .ZN(new_n13432_));
  NAND2_X1   g13338(.A1(new_n10809_), .A2(new_n962_), .ZN(new_n13433_));
  AOI22_X1   g13339(.A1(new_n87_), .A2(new_n10745_), .B1(new_n11002_), .B2(new_n4406_), .ZN(new_n13434_));
  AOI21_X1   g13340(.A1(new_n13433_), .A2(new_n13434_), .B(new_n82_), .ZN(new_n13435_));
  NAND2_X1   g13341(.A1(new_n11046_), .A2(new_n13435_), .ZN(new_n13436_));
  XOR2_X1    g13342(.A1(new_n13432_), .A2(new_n13436_), .Z(new_n13437_));
  INV_X1     g13343(.I(new_n13437_), .ZN(new_n13438_));
  XOR2_X1    g13344(.A1(new_n13431_), .A2(new_n13438_), .Z(new_n13439_));
  AND2_X2    g13345(.A1(new_n13431_), .A2(new_n13437_), .Z(new_n13440_));
  NOR2_X1    g13346(.A1(new_n13431_), .A2(new_n13437_), .ZN(new_n13441_));
  NOR2_X1    g13347(.A1(new_n13440_), .A2(new_n13441_), .ZN(new_n13442_));
  MUX2_X1    g13348(.I0(new_n13439_), .I1(new_n13442_), .S(new_n13427_), .Z(new_n13443_));
  AOI22_X1   g13349(.A1(new_n10652_), .A2(new_n4767_), .B1(new_n4613_), .B2(new_n10805_), .ZN(new_n13444_));
  NOR2_X1    g13350(.A1(new_n10646_), .A2(new_n1128_), .ZN(new_n13445_));
  OAI21_X1   g13351(.A1(new_n13445_), .A2(new_n13444_), .B(new_n65_), .ZN(new_n13446_));
  NAND2_X1   g13352(.A1(new_n13446_), .A2(new_n117_), .ZN(new_n13447_));
  XOR2_X1    g13353(.A1(new_n11246_), .A2(new_n13447_), .Z(new_n13448_));
  NOR2_X1    g13354(.A1(new_n13448_), .A2(new_n13443_), .ZN(new_n13449_));
  INV_X1     g13355(.I(new_n13449_), .ZN(new_n13450_));
  NOR2_X1    g13356(.A1(new_n13426_), .A2(new_n13450_), .ZN(new_n13451_));
  INV_X1     g13357(.I(new_n13451_), .ZN(new_n13452_));
  NAND2_X1   g13358(.A1(new_n13426_), .A2(new_n13450_), .ZN(new_n13453_));
  AOI21_X1   g13359(.A1(new_n13452_), .A2(new_n13453_), .B(new_n13423_), .ZN(new_n13454_));
  NAND3_X1   g13360(.A1(new_n13452_), .A2(new_n13423_), .A3(new_n13453_), .ZN(new_n13455_));
  INV_X1     g13361(.I(new_n13455_), .ZN(new_n13456_));
  NOR3_X1    g13362(.A1(new_n13456_), .A2(new_n13422_), .A3(new_n13454_), .ZN(new_n13457_));
  INV_X1     g13363(.I(new_n13457_), .ZN(new_n13458_));
  OAI21_X1   g13364(.A1(new_n13456_), .A2(new_n13454_), .B(new_n13422_), .ZN(new_n13459_));
  AOI21_X1   g13365(.A1(new_n13458_), .A2(new_n13459_), .B(new_n13418_), .ZN(new_n13460_));
  OAI21_X1   g13366(.A1(new_n12816_), .A2(new_n12817_), .B(new_n12819_), .ZN(new_n13461_));
  OAI21_X1   g13367(.A1(new_n12785_), .A2(new_n12824_), .B(new_n13461_), .ZN(new_n13462_));
  INV_X1     g13368(.I(new_n13454_), .ZN(new_n13463_));
  NAND3_X1   g13369(.A1(new_n13463_), .A2(new_n13455_), .A3(new_n13422_), .ZN(new_n13464_));
  INV_X1     g13370(.I(new_n13422_), .ZN(new_n13465_));
  OAI21_X1   g13371(.A1(new_n13456_), .A2(new_n13454_), .B(new_n13465_), .ZN(new_n13466_));
  AOI21_X1   g13372(.A1(new_n13464_), .A2(new_n13466_), .B(new_n13462_), .ZN(new_n13467_));
  NOR2_X1    g13373(.A1(new_n13460_), .A2(new_n13467_), .ZN(new_n13468_));
  OAI22_X1   g13374(.A1(new_n10870_), .A2(new_n5398_), .B1(new_n5336_), .B2(new_n10861_), .ZN(new_n13469_));
  AOI21_X1   g13375(.A1(new_n13469_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n13470_));
  XOR2_X1    g13376(.A1(new_n11648_), .A2(new_n13470_), .Z(new_n13471_));
  NOR2_X1    g13377(.A1(new_n13468_), .A2(new_n13471_), .ZN(new_n13472_));
  NAND2_X1   g13378(.A1(new_n12839_), .A2(new_n13472_), .ZN(new_n13473_));
  OR2_X2     g13379(.A1(new_n13460_), .A2(new_n13467_), .Z(new_n13474_));
  INV_X1     g13380(.I(new_n13471_), .ZN(new_n13475_));
  NAND2_X1   g13381(.A1(new_n13474_), .A2(new_n13475_), .ZN(new_n13476_));
  NAND3_X1   g13382(.A1(new_n13476_), .A2(new_n12782_), .A3(new_n12838_), .ZN(new_n13477_));
  AOI21_X1   g13383(.A1(new_n13473_), .A2(new_n13477_), .B(new_n12837_), .ZN(new_n13478_));
  INV_X1     g13384(.I(new_n12837_), .ZN(new_n13479_));
  AOI21_X1   g13385(.A1(new_n12782_), .A2(new_n12838_), .B(new_n13476_), .ZN(new_n13480_));
  NOR2_X1    g13386(.A1(new_n12839_), .A2(new_n13472_), .ZN(new_n13481_));
  NOR3_X1    g13387(.A1(new_n13480_), .A2(new_n13481_), .A3(new_n13479_), .ZN(new_n13482_));
  OAI22_X1   g13388(.A1(new_n10619_), .A2(new_n1620_), .B1(new_n5420_), .B2(new_n10885_), .ZN(new_n13483_));
  AOI21_X1   g13389(.A1(new_n13483_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n13484_));
  XOR2_X1    g13390(.A1(new_n12074_), .A2(new_n13484_), .Z(new_n13485_));
  INV_X1     g13391(.I(new_n13485_), .ZN(new_n13486_));
  OAI21_X1   g13392(.A1(new_n13482_), .A2(new_n13478_), .B(new_n13486_), .ZN(new_n13487_));
  NOR2_X1    g13393(.A1(new_n13416_), .A2(new_n13487_), .ZN(new_n13488_));
  OAI22_X1   g13394(.A1(new_n12646_), .A2(new_n12642_), .B1(new_n12717_), .B2(new_n12719_), .ZN(new_n13489_));
  OAI21_X1   g13395(.A1(new_n13480_), .A2(new_n13481_), .B(new_n13479_), .ZN(new_n13490_));
  NAND3_X1   g13396(.A1(new_n13473_), .A2(new_n13477_), .A3(new_n12837_), .ZN(new_n13491_));
  AOI21_X1   g13397(.A1(new_n13490_), .A2(new_n13491_), .B(new_n13485_), .ZN(new_n13492_));
  NOR2_X1    g13398(.A1(new_n13489_), .A2(new_n13492_), .ZN(new_n13493_));
  OAI21_X1   g13399(.A1(new_n13488_), .A2(new_n13493_), .B(new_n12845_), .ZN(new_n13494_));
  NAND2_X1   g13400(.A1(new_n13489_), .A2(new_n13492_), .ZN(new_n13495_));
  NAND2_X1   g13401(.A1(new_n13416_), .A2(new_n13487_), .ZN(new_n13496_));
  NAND3_X1   g13402(.A1(new_n13496_), .A2(new_n13495_), .A3(new_n12854_), .ZN(new_n13497_));
  OAI22_X1   g13403(.A1(new_n10606_), .A2(new_n643_), .B1(new_n5967_), .B2(new_n10901_), .ZN(new_n13498_));
  AOI21_X1   g13404(.A1(new_n13498_), .A2(new_n279_), .B(new_n643_), .ZN(new_n13499_));
  XOR2_X1    g13405(.A1(new_n12211_), .A2(new_n13499_), .Z(new_n13500_));
  AOI21_X1   g13406(.A1(new_n13494_), .A2(new_n13497_), .B(new_n13500_), .ZN(new_n13501_));
  NAND2_X1   g13407(.A1(new_n13414_), .A2(new_n13501_), .ZN(new_n13502_));
  INV_X1     g13408(.I(new_n13502_), .ZN(new_n13503_));
  NOR2_X1    g13409(.A1(new_n13414_), .A2(new_n13501_), .ZN(new_n13504_));
  OAI21_X1   g13410(.A1(new_n13503_), .A2(new_n13504_), .B(new_n12865_), .ZN(new_n13505_));
  INV_X1     g13411(.I(new_n13501_), .ZN(new_n13506_));
  NAND2_X1   g13412(.A1(new_n12867_), .A2(new_n13506_), .ZN(new_n13507_));
  NAND3_X1   g13413(.A1(new_n13507_), .A2(new_n12870_), .A3(new_n13502_), .ZN(new_n13508_));
  NAND2_X1   g13414(.A1(new_n13505_), .A2(new_n13508_), .ZN(new_n13509_));
  OAI22_X1   g13415(.A1(new_n10589_), .A2(new_n1078_), .B1(new_n12623_), .B2(new_n6757_), .ZN(new_n13510_));
  AOI21_X1   g13416(.A1(new_n13510_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n13511_));
  XOR2_X1    g13417(.A1(new_n12622_), .A2(new_n13511_), .Z(new_n13512_));
  INV_X1     g13418(.I(new_n13512_), .ZN(new_n13513_));
  NAND2_X1   g13419(.A1(new_n13509_), .A2(new_n13513_), .ZN(new_n13514_));
  NOR2_X1    g13420(.A1(new_n13514_), .A2(new_n13413_), .ZN(new_n13515_));
  OAI22_X1   g13421(.A1(new_n12635_), .A2(new_n12632_), .B1(new_n12757_), .B2(new_n12758_), .ZN(new_n13516_));
  AOI21_X1   g13422(.A1(new_n13509_), .A2(new_n13513_), .B(new_n13516_), .ZN(new_n13517_));
  OAI21_X1   g13423(.A1(new_n13515_), .A2(new_n13517_), .B(new_n12882_), .ZN(new_n13518_));
  NAND3_X1   g13424(.A1(new_n13516_), .A2(new_n13509_), .A3(new_n13513_), .ZN(new_n13519_));
  NAND2_X1   g13425(.A1(new_n13514_), .A2(new_n13413_), .ZN(new_n13520_));
  NAND3_X1   g13426(.A1(new_n13520_), .A2(new_n13519_), .A3(new_n12877_), .ZN(new_n13521_));
  NAND2_X1   g13427(.A1(new_n13518_), .A2(new_n13521_), .ZN(new_n13522_));
  OAI22_X1   g13428(.A1(new_n10583_), .A2(new_n2495_), .B1(new_n7837_), .B2(new_n10928_), .ZN(new_n13523_));
  AOI21_X1   g13429(.A1(new_n13523_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n13524_));
  XNOR2_X1   g13430(.A1(new_n13378_), .A2(new_n13524_), .ZN(new_n13525_));
  INV_X1     g13431(.I(new_n13525_), .ZN(new_n13526_));
  NAND3_X1   g13432(.A1(new_n13411_), .A2(new_n13522_), .A3(new_n13526_), .ZN(new_n13527_));
  NAND2_X1   g13433(.A1(new_n13522_), .A2(new_n13526_), .ZN(new_n13528_));
  NAND2_X1   g13434(.A1(new_n13528_), .A2(new_n13410_), .ZN(new_n13529_));
  AOI21_X1   g13435(.A1(new_n13527_), .A2(new_n13529_), .B(new_n12899_), .ZN(new_n13530_));
  OAI21_X1   g13436(.A1(new_n12884_), .A2(new_n12881_), .B(new_n12894_), .ZN(new_n13531_));
  NOR2_X1    g13437(.A1(new_n13528_), .A2(new_n13410_), .ZN(new_n13532_));
  AOI21_X1   g13438(.A1(new_n13522_), .A2(new_n13526_), .B(new_n13411_), .ZN(new_n13533_));
  NOR3_X1    g13439(.A1(new_n13533_), .A2(new_n13532_), .A3(new_n13531_), .ZN(new_n13534_));
  NOR2_X1    g13440(.A1(new_n13534_), .A2(new_n13530_), .ZN(new_n13535_));
  INV_X1     g13441(.I(new_n10941_), .ZN(new_n13536_));
  INV_X1     g13442(.I(new_n12905_), .ZN(new_n13537_));
  NOR2_X1    g13443(.A1(new_n10577_), .A2(new_n10937_), .ZN(new_n13538_));
  NOR2_X1    g13444(.A1(new_n10958_), .A2(new_n10938_), .ZN(new_n13539_));
  OAI21_X1   g13445(.A1(new_n13539_), .A2(new_n13538_), .B(new_n13537_), .ZN(new_n13540_));
  NOR2_X1    g13446(.A1(new_n13536_), .A2(new_n13540_), .ZN(new_n13541_));
  NAND2_X1   g13447(.A1(new_n13536_), .A2(new_n13540_), .ZN(new_n13542_));
  INV_X1     g13448(.I(new_n13542_), .ZN(new_n13543_));
  NOR2_X1    g13449(.A1(new_n13543_), .A2(new_n13541_), .ZN(new_n13544_));
  OAI22_X1   g13450(.A1(new_n3042_), .A2(new_n10938_), .B1(new_n10952_), .B2(new_n8830_), .ZN(new_n13545_));
  OAI21_X1   g13451(.A1(new_n10577_), .A2(new_n3040_), .B(new_n13545_), .ZN(new_n13546_));
  AOI21_X1   g13452(.A1(new_n13546_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n13547_));
  XOR2_X1    g13453(.A1(new_n13544_), .A2(new_n13547_), .Z(new_n13548_));
  NOR3_X1    g13454(.A1(new_n13405_), .A2(new_n13535_), .A3(new_n13548_), .ZN(new_n13549_));
  NOR2_X1    g13455(.A1(new_n12925_), .A2(new_n12929_), .ZN(new_n13550_));
  AOI21_X1   g13456(.A1(new_n13341_), .A2(new_n13342_), .B(new_n13331_), .ZN(new_n13551_));
  NOR3_X1    g13457(.A1(new_n13358_), .A2(new_n13357_), .A3(new_n13356_), .ZN(new_n13552_));
  AOI21_X1   g13458(.A1(new_n13354_), .A2(new_n13351_), .B(new_n13348_), .ZN(new_n13553_));
  OAI21_X1   g13459(.A1(new_n13552_), .A2(new_n13553_), .B(new_n12929_), .ZN(new_n13554_));
  AOI21_X1   g13460(.A1(new_n13554_), .A2(new_n13551_), .B(new_n13550_), .ZN(new_n13555_));
  NOR3_X1    g13461(.A1(new_n13369_), .A2(new_n13371_), .A3(new_n13382_), .ZN(new_n13556_));
  NOR3_X1    g13462(.A1(new_n13555_), .A2(new_n13362_), .A3(new_n13556_), .ZN(new_n13557_));
  INV_X1     g13463(.I(new_n13385_), .ZN(new_n13558_));
  NAND2_X1   g13464(.A1(new_n13399_), .A2(new_n13402_), .ZN(new_n13559_));
  OAI21_X1   g13465(.A1(new_n13557_), .A2(new_n13558_), .B(new_n13559_), .ZN(new_n13560_));
  NOR2_X1    g13466(.A1(new_n13535_), .A2(new_n13548_), .ZN(new_n13561_));
  NOR2_X1    g13467(.A1(new_n13561_), .A2(new_n13560_), .ZN(new_n13562_));
  OAI21_X1   g13468(.A1(new_n13549_), .A2(new_n13562_), .B(new_n12915_), .ZN(new_n13563_));
  NAND2_X1   g13469(.A1(new_n13561_), .A2(new_n13560_), .ZN(new_n13564_));
  OAI21_X1   g13470(.A1(new_n13535_), .A2(new_n13548_), .B(new_n13405_), .ZN(new_n13565_));
  NAND3_X1   g13471(.A1(new_n13565_), .A2(new_n12914_), .A3(new_n13564_), .ZN(new_n13566_));
  AOI21_X1   g13472(.A1(new_n13566_), .A2(new_n13563_), .B(new_n10981_), .ZN(new_n13567_));
  NAND3_X1   g13473(.A1(new_n13140_), .A2(new_n13127_), .A3(new_n13138_), .ZN(new_n13568_));
  OAI21_X1   g13474(.A1(new_n13128_), .A2(new_n13126_), .B(new_n13141_), .ZN(new_n13569_));
  NAND2_X1   g13475(.A1(new_n13569_), .A2(new_n13568_), .ZN(new_n13570_));
  NAND2_X1   g13476(.A1(new_n13570_), .A2(new_n13121_), .ZN(new_n13571_));
  INV_X1     g13477(.I(new_n13121_), .ZN(new_n13572_));
  NAND2_X1   g13478(.A1(new_n13142_), .A2(new_n13139_), .ZN(new_n13573_));
  NAND2_X1   g13479(.A1(new_n13572_), .A2(new_n13573_), .ZN(new_n13574_));
  NAND2_X1   g13480(.A1(new_n13574_), .A2(new_n13571_), .ZN(new_n13575_));
  INV_X1     g13481(.I(new_n12351_), .ZN(new_n13576_));
  INV_X1     g13482(.I(new_n13031_), .ZN(new_n13577_));
  NAND2_X1   g13483(.A1(new_n13577_), .A2(new_n13029_), .ZN(new_n13578_));
  NAND2_X1   g13484(.A1(new_n13578_), .A2(new_n13576_), .ZN(new_n13579_));
  INV_X1     g13485(.I(new_n13049_), .ZN(new_n13580_));
  NOR2_X1    g13486(.A1(new_n13580_), .A2(new_n13047_), .ZN(new_n13581_));
  NAND2_X1   g13487(.A1(new_n13581_), .A2(new_n13052_), .ZN(new_n13582_));
  NOR3_X1    g13488(.A1(new_n13582_), .A2(new_n13042_), .A3(new_n13040_), .ZN(new_n13583_));
  NOR2_X1    g13489(.A1(new_n13578_), .A2(new_n13576_), .ZN(new_n13584_));
  OAI21_X1   g13490(.A1(new_n13583_), .A2(new_n13584_), .B(new_n13579_), .ZN(new_n13585_));
  NAND3_X1   g13491(.A1(new_n13066_), .A2(new_n13060_), .A3(new_n13064_), .ZN(new_n13586_));
  NAND2_X1   g13492(.A1(new_n13069_), .A2(new_n13061_), .ZN(new_n13587_));
  NAND2_X1   g13493(.A1(new_n13587_), .A2(new_n13586_), .ZN(new_n13588_));
  NAND2_X1   g13494(.A1(new_n13588_), .A2(new_n13585_), .ZN(new_n13589_));
  AOI21_X1   g13495(.A1(new_n13064_), .A2(new_n13066_), .B(new_n13061_), .ZN(new_n13590_));
  OAI21_X1   g13496(.A1(new_n13068_), .A2(new_n13590_), .B(new_n13057_), .ZN(new_n13591_));
  NAND2_X1   g13497(.A1(new_n13589_), .A2(new_n13591_), .ZN(new_n13592_));
  NOR3_X1    g13498(.A1(new_n13054_), .A2(new_n13042_), .A3(new_n13040_), .ZN(new_n13593_));
  NAND2_X1   g13499(.A1(new_n13041_), .A2(new_n452_), .ZN(new_n13594_));
  NAND2_X1   g13500(.A1(new_n13039_), .A2(\a[5] ), .ZN(new_n13595_));
  AOI21_X1   g13501(.A1(new_n13594_), .A2(new_n13595_), .B(new_n13582_), .ZN(new_n13596_));
  NOR2_X1    g13502(.A1(new_n13596_), .A2(new_n13593_), .ZN(new_n13597_));
  NOR2_X1    g13503(.A1(new_n10755_), .A2(new_n9408_), .ZN(new_n13598_));
  AOI21_X1   g13504(.A1(new_n10781_), .A2(new_n10782_), .B(new_n9405_), .ZN(new_n13599_));
  OAI21_X1   g13505(.A1(new_n13599_), .A2(new_n13598_), .B(\a[2] ), .ZN(new_n13600_));
  AOI21_X1   g13506(.A1(new_n13600_), .A2(new_n3456_), .B(new_n10762_), .ZN(new_n13601_));
  NAND3_X1   g13507(.A1(new_n10762_), .A2(new_n10780_), .A3(new_n10783_), .ZN(new_n13602_));
  NAND2_X1   g13508(.A1(new_n11009_), .A2(new_n11002_), .ZN(new_n13603_));
  AOI21_X1   g13509(.A1(new_n13603_), .A2(new_n13602_), .B(new_n3412_), .ZN(new_n13604_));
  NOR2_X1    g13510(.A1(new_n11017_), .A2(new_n3412_), .ZN(new_n13605_));
  NAND2_X1   g13511(.A1(new_n10783_), .A2(new_n9416_), .ZN(new_n13606_));
  OAI21_X1   g13512(.A1(new_n10755_), .A2(new_n451_), .B(new_n9406_), .ZN(new_n13607_));
  NAND3_X1   g13513(.A1(new_n13606_), .A2(\a[0] ), .A3(new_n13607_), .ZN(new_n13608_));
  NOR4_X1    g13514(.A1(new_n13604_), .A2(new_n13605_), .A3(new_n13601_), .A4(new_n13608_), .ZN(new_n13609_));
  NAND2_X1   g13515(.A1(new_n13609_), .A2(new_n13051_), .ZN(new_n13610_));
  NOR2_X1    g13516(.A1(new_n10777_), .A2(new_n3456_), .ZN(new_n13611_));
  INV_X1     g13517(.I(new_n13611_), .ZN(new_n13612_));
  AOI21_X1   g13518(.A1(new_n11002_), .A2(new_n10783_), .B(new_n9425_), .ZN(new_n13613_));
  AOI21_X1   g13519(.A1(new_n13612_), .A2(new_n13613_), .B(new_n3414_), .ZN(new_n13614_));
  AOI21_X1   g13520(.A1(new_n11001_), .A2(new_n13614_), .B(new_n451_), .ZN(new_n13615_));
  INV_X1     g13521(.I(new_n13613_), .ZN(new_n13616_));
  OAI21_X1   g13522(.A1(new_n13616_), .A2(new_n13611_), .B(new_n3411_), .ZN(new_n13617_));
  NOR3_X1    g13523(.A1(new_n11188_), .A2(new_n13617_), .A3(\a[2] ), .ZN(new_n13618_));
  OAI22_X1   g13524(.A1(new_n13618_), .A2(new_n13615_), .B1(new_n13609_), .B2(new_n13051_), .ZN(new_n13619_));
  NAND2_X1   g13525(.A1(new_n13619_), .A2(new_n13610_), .ZN(new_n13620_));
  OAI21_X1   g13526(.A1(new_n10762_), .A2(new_n10777_), .B(new_n9433_), .ZN(new_n13621_));
  OAI21_X1   g13527(.A1(new_n10725_), .A2(new_n3456_), .B(new_n13621_), .ZN(new_n13622_));
  AOI21_X1   g13528(.A1(new_n13622_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n13623_));
  NAND3_X1   g13529(.A1(new_n11039_), .A2(new_n11045_), .A3(new_n13623_), .ZN(new_n13624_));
  AOI21_X1   g13530(.A1(new_n11131_), .A2(new_n10774_), .B(new_n10725_), .ZN(new_n13625_));
  INV_X1     g13531(.I(new_n11040_), .ZN(new_n13626_));
  OAI21_X1   g13532(.A1(new_n10786_), .A2(new_n10780_), .B(new_n10745_), .ZN(new_n13627_));
  AOI21_X1   g13533(.A1(new_n13627_), .A2(new_n13626_), .B(new_n10809_), .ZN(new_n13628_));
  INV_X1     g13534(.I(new_n13621_), .ZN(new_n13629_));
  AOI21_X1   g13535(.A1(new_n10807_), .A2(new_n10808_), .B(new_n3456_), .ZN(new_n13630_));
  OAI21_X1   g13536(.A1(new_n13630_), .A2(new_n13629_), .B(new_n451_), .ZN(new_n13631_));
  NAND2_X1   g13537(.A1(new_n13631_), .A2(new_n3411_), .ZN(new_n13632_));
  OAI21_X1   g13538(.A1(new_n13628_), .A2(new_n13625_), .B(new_n13632_), .ZN(new_n13633_));
  NAND2_X1   g13539(.A1(new_n13633_), .A2(new_n13624_), .ZN(new_n13634_));
  NAND2_X1   g13540(.A1(new_n13634_), .A2(new_n13620_), .ZN(new_n13635_));
  NAND2_X1   g13541(.A1(new_n13050_), .A2(new_n13053_), .ZN(new_n13636_));
  NAND2_X1   g13542(.A1(new_n13582_), .A2(new_n13636_), .ZN(new_n13637_));
  OAI21_X1   g13543(.A1(new_n13634_), .A2(new_n13620_), .B(new_n13637_), .ZN(new_n13638_));
  AOI21_X1   g13544(.A1(new_n13638_), .A2(new_n13635_), .B(new_n13597_), .ZN(new_n13639_));
  NAND3_X1   g13545(.A1(new_n13638_), .A2(new_n13635_), .A3(new_n13597_), .ZN(new_n13640_));
  INV_X1     g13546(.I(new_n11062_), .ZN(new_n13641_));
  AOI21_X1   g13547(.A1(new_n10797_), .A2(new_n13641_), .B(new_n10794_), .ZN(new_n13642_));
  AOI21_X1   g13548(.A1(new_n11128_), .A2(new_n10794_), .B(new_n13642_), .ZN(new_n13643_));
  NAND2_X1   g13549(.A1(new_n10794_), .A2(new_n3455_), .ZN(new_n13644_));
  AOI21_X1   g13550(.A1(new_n10809_), .A2(new_n10745_), .B(new_n9425_), .ZN(new_n13645_));
  AOI21_X1   g13551(.A1(new_n13644_), .A2(new_n13645_), .B(new_n3414_), .ZN(new_n13646_));
  INV_X1     g13552(.I(new_n13646_), .ZN(new_n13647_));
  OAI21_X1   g13553(.A1(new_n13643_), .A2(new_n13647_), .B(\a[2] ), .ZN(new_n13648_));
  NAND3_X1   g13554(.A1(new_n11064_), .A2(new_n451_), .A3(new_n13646_), .ZN(new_n13649_));
  NAND2_X1   g13555(.A1(new_n13648_), .A2(new_n13649_), .ZN(new_n13650_));
  AOI21_X1   g13556(.A1(new_n13640_), .A2(new_n13650_), .B(new_n13639_), .ZN(new_n13651_));
  AOI22_X1   g13557(.A1(new_n11141_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n10691_), .ZN(new_n13652_));
  OAI21_X1   g13558(.A1(new_n13652_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n13653_));
  NOR3_X1    g13559(.A1(new_n11135_), .A2(new_n11139_), .A3(new_n13653_), .ZN(new_n13654_));
  OAI22_X1   g13560(.A1(new_n13081_), .A2(new_n9425_), .B1(new_n3456_), .B2(new_n10792_), .ZN(new_n13655_));
  AOI21_X1   g13561(.A1(new_n13655_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n13656_));
  AOI21_X1   g13562(.A1(new_n11332_), .A2(new_n11331_), .B(new_n13656_), .ZN(new_n13657_));
  NOR2_X1    g13563(.A1(new_n13654_), .A2(new_n13657_), .ZN(new_n13658_));
  NOR2_X1    g13564(.A1(new_n13651_), .A2(new_n13658_), .ZN(new_n13659_));
  NOR2_X1    g13565(.A1(new_n13583_), .A2(new_n12351_), .ZN(new_n13660_));
  NAND2_X1   g13566(.A1(new_n13583_), .A2(new_n12351_), .ZN(new_n13661_));
  INV_X1     g13567(.I(new_n13661_), .ZN(new_n13662_));
  NOR3_X1    g13568(.A1(new_n13662_), .A2(new_n13660_), .A3(new_n13032_), .ZN(new_n13663_));
  NAND2_X1   g13569(.A1(new_n13055_), .A2(new_n13576_), .ZN(new_n13664_));
  AOI21_X1   g13570(.A1(new_n13664_), .A2(new_n13661_), .B(new_n13578_), .ZN(new_n13665_));
  NOR2_X1    g13571(.A1(new_n13663_), .A2(new_n13665_), .ZN(new_n13666_));
  AOI21_X1   g13572(.A1(new_n13651_), .A2(new_n13658_), .B(new_n13666_), .ZN(new_n13667_));
  OAI21_X1   g13573(.A1(new_n13667_), .A2(new_n13659_), .B(new_n13592_), .ZN(new_n13668_));
  NOR3_X1    g13574(.A1(new_n13667_), .A2(new_n13659_), .A3(new_n13592_), .ZN(new_n13669_));
  NAND2_X1   g13575(.A1(new_n10817_), .A2(new_n3455_), .ZN(new_n13670_));
  NOR2_X1    g13576(.A1(new_n11159_), .A2(new_n9425_), .ZN(new_n13671_));
  AOI21_X1   g13577(.A1(new_n13670_), .A2(new_n13671_), .B(new_n3414_), .ZN(new_n13672_));
  AOI21_X1   g13578(.A1(new_n11158_), .A2(new_n13672_), .B(new_n451_), .ZN(new_n13673_));
  AND3_X2    g13579(.A1(new_n11158_), .A2(new_n451_), .A3(new_n13672_), .Z(new_n13674_));
  NOR2_X1    g13580(.A1(new_n13674_), .A2(new_n13673_), .ZN(new_n13675_));
  OAI21_X1   g13581(.A1(new_n13669_), .A2(new_n13675_), .B(new_n13668_), .ZN(new_n13676_));
  XNOR2_X1   g13582(.A1(new_n11064_), .A2(new_n13074_), .ZN(new_n13677_));
  NOR2_X1    g13583(.A1(new_n13677_), .A2(new_n13072_), .ZN(new_n13678_));
  XOR2_X1    g13584(.A1(new_n12343_), .A2(new_n12354_), .Z(new_n13679_));
  NOR2_X1    g13585(.A1(new_n13075_), .A2(new_n13679_), .ZN(new_n13680_));
  OAI21_X1   g13586(.A1(new_n13678_), .A2(new_n13680_), .B(new_n13071_), .ZN(new_n13681_));
  INV_X1     g13587(.I(new_n13681_), .ZN(new_n13682_));
  AOI21_X1   g13588(.A1(new_n13585_), .A2(new_n13067_), .B(new_n13590_), .ZN(new_n13683_));
  NOR2_X1    g13589(.A1(new_n13677_), .A2(new_n13679_), .ZN(new_n13684_));
  OAI21_X1   g13590(.A1(new_n13684_), .A2(new_n13077_), .B(new_n13683_), .ZN(new_n13685_));
  INV_X1     g13591(.I(new_n13685_), .ZN(new_n13686_));
  OAI21_X1   g13592(.A1(new_n11210_), .A2(new_n11169_), .B(new_n10805_), .ZN(new_n13687_));
  OAI21_X1   g13593(.A1(new_n11241_), .A2(new_n11172_), .B(new_n10658_), .ZN(new_n13688_));
  OAI22_X1   g13594(.A1(new_n11176_), .A2(new_n9425_), .B1(new_n10658_), .B2(new_n3456_), .ZN(new_n13689_));
  AOI21_X1   g13595(.A1(new_n13689_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n13690_));
  NAND3_X1   g13596(.A1(new_n13687_), .A2(new_n13690_), .A3(new_n13688_), .ZN(new_n13691_));
  AOI22_X1   g13597(.A1(new_n13094_), .A2(new_n9433_), .B1(new_n10805_), .B2(new_n3455_), .ZN(new_n13692_));
  OAI21_X1   g13598(.A1(new_n13692_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n13693_));
  OAI21_X1   g13599(.A1(new_n11171_), .A2(new_n11174_), .B(new_n13693_), .ZN(new_n13694_));
  AND2_X2    g13600(.A1(new_n13694_), .A2(new_n13691_), .Z(new_n13695_));
  OAI21_X1   g13601(.A1(new_n13682_), .A2(new_n13686_), .B(new_n13695_), .ZN(new_n13696_));
  NAND2_X1   g13602(.A1(new_n13694_), .A2(new_n13691_), .ZN(new_n13697_));
  NAND3_X1   g13603(.A1(new_n13697_), .A2(new_n13681_), .A3(new_n13685_), .ZN(new_n13698_));
  INV_X1     g13604(.I(new_n13698_), .ZN(new_n13699_));
  AOI21_X1   g13605(.A1(new_n13676_), .A2(new_n13696_), .B(new_n13699_), .ZN(new_n13700_));
  NAND2_X1   g13606(.A1(new_n11140_), .A2(new_n13083_), .ZN(new_n13701_));
  NAND2_X1   g13607(.A1(new_n11333_), .A2(new_n13084_), .ZN(new_n13702_));
  NAND3_X1   g13608(.A1(new_n13080_), .A2(new_n13701_), .A3(new_n13702_), .ZN(new_n13703_));
  AND2_X2    g13609(.A1(new_n13079_), .A2(new_n13001_), .Z(new_n13704_));
  OAI21_X1   g13610(.A1(new_n13085_), .A2(new_n13086_), .B(new_n13704_), .ZN(new_n13705_));
  AOI21_X1   g13611(.A1(new_n13705_), .A2(new_n13703_), .B(new_n13078_), .ZN(new_n13706_));
  NAND2_X1   g13612(.A1(new_n13677_), .A2(new_n13679_), .ZN(new_n13707_));
  OAI21_X1   g13613(.A1(new_n13683_), .A2(new_n13684_), .B(new_n13707_), .ZN(new_n13708_));
  NAND3_X1   g13614(.A1(new_n13704_), .A2(new_n13701_), .A3(new_n13702_), .ZN(new_n13709_));
  AOI21_X1   g13615(.A1(new_n13709_), .A2(new_n13089_), .B(new_n13708_), .ZN(new_n13710_));
  NOR2_X1    g13616(.A1(new_n13710_), .A2(new_n13706_), .ZN(new_n13711_));
  NAND2_X1   g13617(.A1(new_n10805_), .A2(new_n10817_), .ZN(new_n13712_));
  AOI22_X1   g13618(.A1(new_n13712_), .A2(new_n9433_), .B1(new_n10652_), .B2(new_n3455_), .ZN(new_n13713_));
  NOR2_X1    g13619(.A1(new_n13713_), .A2(\a[2] ), .ZN(new_n13714_));
  NOR4_X1    g13620(.A1(new_n11218_), .A2(new_n11223_), .A3(new_n3414_), .A4(new_n13714_), .ZN(new_n13715_));
  NAND3_X1   g13621(.A1(new_n11222_), .A2(new_n11219_), .A3(new_n10658_), .ZN(new_n13716_));
  OAI21_X1   g13622(.A1(new_n11217_), .A2(new_n11211_), .B(new_n10805_), .ZN(new_n13717_));
  OAI22_X1   g13623(.A1(new_n10819_), .A2(new_n9425_), .B1(new_n11214_), .B2(new_n3456_), .ZN(new_n13718_));
  AOI21_X1   g13624(.A1(new_n13718_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n13719_));
  AOI21_X1   g13625(.A1(new_n13717_), .A2(new_n13716_), .B(new_n13719_), .ZN(new_n13720_));
  NOR3_X1    g13626(.A1(new_n13711_), .A2(new_n13715_), .A3(new_n13720_), .ZN(new_n13721_));
  NOR2_X1    g13627(.A1(new_n13715_), .A2(new_n13720_), .ZN(new_n13722_));
  NOR3_X1    g13628(.A1(new_n13722_), .A2(new_n13710_), .A3(new_n13706_), .ZN(new_n13723_));
  INV_X1     g13629(.I(new_n13723_), .ZN(new_n13724_));
  OAI21_X1   g13630(.A1(new_n13700_), .A2(new_n13721_), .B(new_n13724_), .ZN(new_n13725_));
  AOI21_X1   g13631(.A1(new_n10652_), .A2(new_n10805_), .B(new_n9425_), .ZN(new_n13726_));
  INV_X1     g13632(.I(new_n13726_), .ZN(new_n13727_));
  NAND2_X1   g13633(.A1(new_n10828_), .A2(new_n3455_), .ZN(new_n13728_));
  AOI21_X1   g13634(.A1(new_n13728_), .A2(new_n13727_), .B(\a[2] ), .ZN(new_n13729_));
  NOR4_X1    g13635(.A1(new_n13134_), .A2(new_n13729_), .A3(new_n11237_), .A4(new_n3414_), .ZN(new_n13730_));
  NOR2_X1    g13636(.A1(new_n13729_), .A2(new_n3414_), .ZN(new_n13731_));
  NOR2_X1    g13637(.A1(new_n13135_), .A2(new_n13731_), .ZN(new_n13732_));
  OR2_X2     g13638(.A1(new_n13732_), .A2(new_n13730_), .Z(new_n13733_));
  NAND2_X1   g13639(.A1(new_n13725_), .A2(new_n13733_), .ZN(new_n13734_));
  NAND3_X1   g13640(.A1(new_n13019_), .A2(new_n13023_), .A3(new_n13020_), .ZN(new_n13735_));
  NAND2_X1   g13641(.A1(new_n13093_), .A2(new_n13735_), .ZN(new_n13736_));
  NAND2_X1   g13642(.A1(new_n13708_), .A2(new_n13709_), .ZN(new_n13737_));
  NAND2_X1   g13643(.A1(new_n13737_), .A2(new_n13089_), .ZN(new_n13738_));
  XOR2_X1    g13644(.A1(new_n13738_), .A2(new_n13736_), .Z(new_n13739_));
  OAI21_X1   g13645(.A1(new_n13725_), .A2(new_n13733_), .B(new_n13739_), .ZN(new_n13740_));
  NAND4_X1   g13646(.A1(new_n13737_), .A2(new_n13093_), .A3(new_n13735_), .A4(new_n13089_), .ZN(new_n13741_));
  AOI21_X1   g13647(.A1(new_n12993_), .A2(new_n12996_), .B(new_n13100_), .ZN(new_n13742_));
  NAND2_X1   g13648(.A1(new_n13742_), .A2(new_n13741_), .ZN(new_n13743_));
  AOI21_X1   g13649(.A1(new_n12994_), .A2(new_n12995_), .B(new_n11906_), .ZN(new_n13744_));
  NOR3_X1    g13650(.A1(new_n12992_), .A2(new_n12989_), .A3(new_n12370_), .ZN(new_n13745_));
  OAI22_X1   g13651(.A1(new_n13745_), .A2(new_n13744_), .B1(new_n13097_), .B2(new_n13099_), .ZN(new_n13746_));
  NAND2_X1   g13652(.A1(new_n13746_), .A2(new_n13091_), .ZN(new_n13747_));
  AOI21_X1   g13653(.A1(new_n13747_), .A2(new_n13743_), .B(new_n13024_), .ZN(new_n13748_));
  NOR2_X1    g13654(.A1(new_n13746_), .A2(new_n13091_), .ZN(new_n13749_));
  NOR2_X1    g13655(.A1(new_n13742_), .A2(new_n13741_), .ZN(new_n13750_));
  NOR3_X1    g13656(.A1(new_n13749_), .A2(new_n13750_), .A3(new_n13093_), .ZN(new_n13751_));
  NOR2_X1    g13657(.A1(new_n13748_), .A2(new_n13751_), .ZN(new_n13752_));
  AOI21_X1   g13658(.A1(new_n13740_), .A2(new_n13734_), .B(new_n13752_), .ZN(new_n13753_));
  NAND3_X1   g13659(.A1(new_n13740_), .A2(new_n13734_), .A3(new_n13752_), .ZN(new_n13754_));
  NAND2_X1   g13660(.A1(new_n10638_), .A2(new_n3455_), .ZN(new_n13755_));
  AOI21_X1   g13661(.A1(new_n10828_), .A2(new_n10652_), .B(new_n9425_), .ZN(new_n13756_));
  AOI21_X1   g13662(.A1(new_n13755_), .A2(new_n13756_), .B(new_n3414_), .ZN(new_n13757_));
  AOI21_X1   g13663(.A1(new_n11268_), .A2(new_n13757_), .B(new_n451_), .ZN(new_n13758_));
  INV_X1     g13664(.I(new_n13758_), .ZN(new_n13759_));
  NAND3_X1   g13665(.A1(new_n11268_), .A2(new_n451_), .A3(new_n13757_), .ZN(new_n13760_));
  NAND2_X1   g13666(.A1(new_n13759_), .A2(new_n13760_), .ZN(new_n13761_));
  AOI21_X1   g13667(.A1(new_n13754_), .A2(new_n13761_), .B(new_n13753_), .ZN(new_n13762_));
  NOR2_X1    g13668(.A1(new_n13118_), .A2(new_n13116_), .ZN(new_n13763_));
  NOR2_X1    g13669(.A1(new_n13112_), .A2(new_n13115_), .ZN(new_n13764_));
  OAI21_X1   g13670(.A1(new_n13763_), .A2(new_n13764_), .B(new_n13103_), .ZN(new_n13765_));
  NOR2_X1    g13671(.A1(new_n13116_), .A2(new_n13112_), .ZN(new_n13766_));
  NOR2_X1    g13672(.A1(new_n13119_), .A2(new_n13766_), .ZN(new_n13767_));
  OAI21_X1   g13673(.A1(new_n13103_), .A2(new_n13767_), .B(new_n13765_), .ZN(new_n13768_));
  INV_X1     g13674(.I(new_n13768_), .ZN(new_n13769_));
  NOR2_X1    g13675(.A1(new_n13762_), .A2(new_n13769_), .ZN(new_n13770_));
  NOR2_X1    g13676(.A1(new_n10633_), .A2(new_n3456_), .ZN(new_n13771_));
  NAND2_X1   g13677(.A1(new_n10829_), .A2(new_n9433_), .ZN(new_n13772_));
  OAI21_X1   g13678(.A1(new_n13771_), .A2(new_n13772_), .B(new_n3411_), .ZN(new_n13773_));
  INV_X1     g13679(.I(new_n13773_), .ZN(new_n13774_));
  AOI21_X1   g13680(.A1(new_n11987_), .A2(new_n13774_), .B(new_n451_), .ZN(new_n13775_));
  NOR3_X1    g13681(.A1(new_n11385_), .A2(\a[2] ), .A3(new_n13773_), .ZN(new_n13776_));
  NOR2_X1    g13682(.A1(new_n13776_), .A2(new_n13775_), .ZN(new_n13777_));
  AOI21_X1   g13683(.A1(new_n13762_), .A2(new_n13769_), .B(new_n13777_), .ZN(new_n13778_));
  OAI21_X1   g13684(.A1(new_n13778_), .A2(new_n13770_), .B(new_n13575_), .ZN(new_n13779_));
  NOR3_X1    g13685(.A1(new_n13778_), .A2(new_n13770_), .A3(new_n13575_), .ZN(new_n13780_));
  NAND2_X1   g13686(.A1(new_n10630_), .A2(new_n3455_), .ZN(new_n13781_));
  NAND3_X1   g13687(.A1(new_n13781_), .A2(new_n9433_), .A3(new_n11446_), .ZN(new_n13782_));
  NAND2_X1   g13688(.A1(new_n13782_), .A2(new_n3411_), .ZN(new_n13783_));
  OAI21_X1   g13689(.A1(new_n11445_), .A2(new_n13783_), .B(\a[2] ), .ZN(new_n13784_));
  OR3_X2     g13690(.A1(new_n11445_), .A2(\a[2] ), .A3(new_n13783_), .Z(new_n13785_));
  NAND2_X1   g13691(.A1(new_n13785_), .A2(new_n13784_), .ZN(new_n13786_));
  INV_X1     g13692(.I(new_n13786_), .ZN(new_n13787_));
  OAI21_X1   g13693(.A1(new_n13780_), .A2(new_n13787_), .B(new_n13779_), .ZN(new_n13788_));
  NAND2_X1   g13694(.A1(new_n11608_), .A2(new_n9433_), .ZN(new_n13789_));
  OAI21_X1   g13695(.A1(new_n3456_), .A2(new_n10844_), .B(new_n13789_), .ZN(new_n13790_));
  AOI21_X1   g13696(.A1(new_n13790_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n13791_));
  INV_X1     g13697(.I(new_n13791_), .ZN(new_n13792_));
  NOR2_X1    g13698(.A1(new_n11607_), .A2(new_n13792_), .ZN(new_n13793_));
  AOI21_X1   g13699(.A1(new_n11606_), .A2(new_n11604_), .B(new_n13791_), .ZN(new_n13794_));
  NOR2_X1    g13700(.A1(new_n13793_), .A2(new_n13794_), .ZN(new_n13795_));
  INV_X1     g13701(.I(new_n13795_), .ZN(new_n13796_));
  NAND2_X1   g13702(.A1(new_n13788_), .A2(new_n13796_), .ZN(new_n13797_));
  NAND2_X1   g13703(.A1(new_n13121_), .A2(new_n13139_), .ZN(new_n13798_));
  NAND2_X1   g13704(.A1(new_n13798_), .A2(new_n13142_), .ZN(new_n13799_));
  AOI21_X1   g13705(.A1(new_n13165_), .A2(new_n13161_), .B(new_n13799_), .ZN(new_n13800_));
  AOI21_X1   g13706(.A1(new_n13152_), .A2(new_n13156_), .B(new_n13160_), .ZN(new_n13801_));
  NOR3_X1    g13707(.A1(new_n13168_), .A2(new_n13801_), .A3(new_n13144_), .ZN(new_n13802_));
  NOR2_X1    g13708(.A1(new_n13802_), .A2(new_n13800_), .ZN(new_n13803_));
  INV_X1     g13709(.I(new_n13803_), .ZN(new_n13804_));
  OAI21_X1   g13710(.A1(new_n13788_), .A2(new_n13796_), .B(new_n13804_), .ZN(new_n13805_));
  AOI22_X1   g13711(.A1(new_n11632_), .A2(new_n9433_), .B1(new_n10857_), .B2(new_n3455_), .ZN(new_n13806_));
  OAI21_X1   g13712(.A1(new_n13806_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n13807_));
  XNOR2_X1   g13713(.A1(new_n11631_), .A2(new_n13807_), .ZN(new_n13808_));
  AOI21_X1   g13714(.A1(new_n13805_), .A2(new_n13797_), .B(new_n13808_), .ZN(new_n13809_));
  NAND3_X1   g13715(.A1(new_n13805_), .A2(new_n13797_), .A3(new_n13808_), .ZN(new_n13810_));
  NAND2_X1   g13716(.A1(new_n13166_), .A2(new_n13161_), .ZN(new_n13811_));
  XNOR2_X1   g13717(.A1(new_n12979_), .A2(new_n13171_), .ZN(new_n13812_));
  XNOR2_X1   g13718(.A1(new_n13812_), .A2(new_n13811_), .ZN(new_n13813_));
  AOI21_X1   g13719(.A1(new_n13810_), .A2(new_n13813_), .B(new_n13809_), .ZN(new_n13814_));
  NOR3_X1    g13720(.A1(new_n13187_), .A2(new_n13177_), .A3(new_n13181_), .ZN(new_n13815_));
  NOR2_X1    g13721(.A1(new_n13182_), .A2(new_n13186_), .ZN(new_n13816_));
  NOR2_X1    g13722(.A1(new_n13816_), .A2(new_n13815_), .ZN(new_n13817_));
  NOR2_X1    g13723(.A1(new_n13188_), .A2(new_n13190_), .ZN(new_n13818_));
  MUX2_X1    g13724(.I0(new_n13817_), .I1(new_n13818_), .S(new_n13174_), .Z(new_n13819_));
  NOR2_X1    g13725(.A1(new_n13814_), .A2(new_n13819_), .ZN(new_n13820_));
  NOR2_X1    g13726(.A1(new_n13225_), .A2(new_n3414_), .ZN(new_n13821_));
  AOI22_X1   g13727(.A1(new_n10625_), .A2(new_n3455_), .B1(new_n11629_), .B2(new_n9433_), .ZN(new_n13822_));
  INV_X1     g13728(.I(new_n13822_), .ZN(new_n13823_));
  NOR3_X1    g13729(.A1(new_n13821_), .A2(new_n451_), .A3(new_n13823_), .ZN(new_n13824_));
  NAND2_X1   g13730(.A1(new_n11648_), .A2(new_n3411_), .ZN(new_n13825_));
  AOI21_X1   g13731(.A1(new_n13825_), .A2(new_n13822_), .B(\a[2] ), .ZN(new_n13826_));
  NOR2_X1    g13732(.A1(new_n13824_), .A2(new_n13826_), .ZN(new_n13827_));
  AOI21_X1   g13733(.A1(new_n13814_), .A2(new_n13819_), .B(new_n13827_), .ZN(new_n13828_));
  NAND2_X1   g13734(.A1(new_n10875_), .A2(new_n3455_), .ZN(new_n13829_));
  NOR2_X1    g13735(.A1(new_n11723_), .A2(new_n9425_), .ZN(new_n13830_));
  AOI21_X1   g13736(.A1(new_n13830_), .A2(new_n13829_), .B(new_n3414_), .ZN(new_n13831_));
  INV_X1     g13737(.I(new_n13831_), .ZN(new_n13832_));
  NOR2_X1    g13738(.A1(new_n11722_), .A2(new_n13832_), .ZN(new_n13833_));
  NOR2_X1    g13739(.A1(new_n13833_), .A2(new_n451_), .ZN(new_n13834_));
  NOR3_X1    g13740(.A1(new_n11722_), .A2(\a[2] ), .A3(new_n13832_), .ZN(new_n13835_));
  NOR2_X1    g13741(.A1(new_n13834_), .A2(new_n13835_), .ZN(new_n13836_));
  INV_X1     g13742(.I(new_n13836_), .ZN(new_n13837_));
  OAI21_X1   g13743(.A1(new_n13828_), .A2(new_n13820_), .B(new_n13837_), .ZN(new_n13838_));
  NOR3_X1    g13744(.A1(new_n13828_), .A2(new_n13820_), .A3(new_n13837_), .ZN(new_n13839_));
  INV_X1     g13745(.I(new_n13191_), .ZN(new_n13840_));
  NOR3_X1    g13746(.A1(new_n13201_), .A2(new_n13194_), .A3(new_n13198_), .ZN(new_n13841_));
  AOI21_X1   g13747(.A1(new_n13195_), .A2(new_n13193_), .B(new_n13199_), .ZN(new_n13842_));
  NOR2_X1    g13748(.A1(new_n13842_), .A2(new_n13841_), .ZN(new_n13843_));
  NOR2_X1    g13749(.A1(new_n13840_), .A2(new_n13843_), .ZN(new_n13844_));
  NAND2_X1   g13750(.A1(new_n13202_), .A2(new_n13200_), .ZN(new_n13845_));
  NOR2_X1    g13751(.A1(new_n13845_), .A2(new_n13191_), .ZN(new_n13846_));
  NOR2_X1    g13752(.A1(new_n13844_), .A2(new_n13846_), .ZN(new_n13847_));
  OAI21_X1   g13753(.A1(new_n13839_), .A2(new_n13847_), .B(new_n13838_), .ZN(new_n13848_));
  NAND2_X1   g13754(.A1(new_n13206_), .A2(new_n13209_), .ZN(new_n13849_));
  NAND2_X1   g13755(.A1(new_n13849_), .A2(new_n13216_), .ZN(new_n13850_));
  NAND3_X1   g13756(.A1(new_n13850_), .A2(new_n13202_), .A3(new_n13218_), .ZN(new_n13851_));
  NAND3_X1   g13757(.A1(new_n13851_), .A2(new_n13191_), .A3(new_n13845_), .ZN(new_n13852_));
  AOI21_X1   g13758(.A1(new_n13851_), .A2(new_n13845_), .B(new_n13191_), .ZN(new_n13853_));
  INV_X1     g13759(.I(new_n13853_), .ZN(new_n13854_));
  NAND2_X1   g13760(.A1(new_n13854_), .A2(new_n13852_), .ZN(new_n13855_));
  NAND2_X1   g13761(.A1(new_n13848_), .A2(new_n13855_), .ZN(new_n13856_));
  NAND2_X1   g13762(.A1(new_n10882_), .A2(new_n3455_), .ZN(new_n13857_));
  NOR2_X1    g13763(.A1(new_n11803_), .A2(new_n9425_), .ZN(new_n13858_));
  AOI21_X1   g13764(.A1(new_n13858_), .A2(new_n13857_), .B(new_n3414_), .ZN(new_n13859_));
  NAND2_X1   g13765(.A1(new_n11802_), .A2(new_n13859_), .ZN(new_n13860_));
  XOR2_X1    g13766(.A1(new_n13860_), .A2(\a[2] ), .Z(new_n13861_));
  INV_X1     g13767(.I(new_n13861_), .ZN(new_n13862_));
  OAI21_X1   g13768(.A1(new_n13848_), .A2(new_n13855_), .B(new_n13862_), .ZN(new_n13863_));
  INV_X1     g13769(.I(new_n13222_), .ZN(new_n13864_));
  NAND3_X1   g13770(.A1(new_n12970_), .A2(new_n13864_), .A3(new_n13228_), .ZN(new_n13865_));
  AOI21_X1   g13771(.A1(new_n12967_), .A2(new_n12968_), .B(new_n12446_), .ZN(new_n13866_));
  NOR3_X1    g13772(.A1(new_n12965_), .A2(new_n12962_), .A3(new_n12959_), .ZN(new_n13867_));
  OAI21_X1   g13773(.A1(new_n13867_), .A2(new_n13866_), .B(new_n13228_), .ZN(new_n13868_));
  NAND2_X1   g13774(.A1(new_n13868_), .A2(new_n13222_), .ZN(new_n13869_));
  AOI21_X1   g13775(.A1(new_n13869_), .A2(new_n13865_), .B(new_n13220_), .ZN(new_n13870_));
  NOR2_X1    g13776(.A1(new_n13868_), .A2(new_n13222_), .ZN(new_n13871_));
  AOI21_X1   g13777(.A1(new_n12970_), .A2(new_n13228_), .B(new_n13864_), .ZN(new_n13872_));
  NOR3_X1    g13778(.A1(new_n13871_), .A2(new_n13872_), .A3(new_n13850_), .ZN(new_n13873_));
  NOR2_X1    g13779(.A1(new_n13873_), .A2(new_n13870_), .ZN(new_n13874_));
  AOI21_X1   g13780(.A1(new_n13863_), .A2(new_n13856_), .B(new_n13874_), .ZN(new_n13875_));
  NAND3_X1   g13781(.A1(new_n13863_), .A2(new_n13856_), .A3(new_n13874_), .ZN(new_n13876_));
  INV_X1     g13782(.I(new_n12074_), .ZN(new_n13877_));
  NAND2_X1   g13783(.A1(new_n10620_), .A2(new_n3455_), .ZN(new_n13878_));
  NOR2_X1    g13784(.A1(new_n10885_), .A2(new_n9425_), .ZN(new_n13879_));
  AOI21_X1   g13785(.A1(new_n13878_), .A2(new_n13879_), .B(new_n3414_), .ZN(new_n13880_));
  NAND2_X1   g13786(.A1(new_n13877_), .A2(new_n13880_), .ZN(new_n13881_));
  XOR2_X1    g13787(.A1(new_n13881_), .A2(\a[2] ), .Z(new_n13882_));
  INV_X1     g13788(.I(new_n13882_), .ZN(new_n13883_));
  AOI21_X1   g13789(.A1(new_n13876_), .A2(new_n13883_), .B(new_n13875_), .ZN(new_n13884_));
  INV_X1     g13790(.I(new_n13238_), .ZN(new_n13885_));
  OAI21_X1   g13791(.A1(new_n13235_), .A2(new_n13232_), .B(new_n13885_), .ZN(new_n13886_));
  INV_X1     g13792(.I(new_n13886_), .ZN(new_n13887_));
  NOR3_X1    g13793(.A1(new_n13235_), .A2(new_n13232_), .A3(new_n13885_), .ZN(new_n13888_));
  NOR2_X1    g13794(.A1(new_n13887_), .A2(new_n13888_), .ZN(new_n13889_));
  INV_X1     g13795(.I(new_n13240_), .ZN(new_n13890_));
  NOR2_X1    g13796(.A1(new_n13890_), .A2(new_n13239_), .ZN(new_n13891_));
  MUX2_X1    g13797(.I0(new_n13889_), .I1(new_n13891_), .S(new_n13231_), .Z(new_n13892_));
  NOR2_X1    g13798(.A1(new_n13884_), .A2(new_n13892_), .ZN(new_n13893_));
  INV_X1     g13799(.I(new_n12090_), .ZN(new_n13894_));
  NOR2_X1    g13800(.A1(new_n13894_), .A2(new_n3414_), .ZN(new_n13895_));
  OAI22_X1   g13801(.A1(new_n12091_), .A2(new_n9425_), .B1(new_n3456_), .B2(new_n10611_), .ZN(new_n13896_));
  NOR3_X1    g13802(.A1(new_n13895_), .A2(new_n451_), .A3(new_n13896_), .ZN(new_n13897_));
  NOR2_X1    g13803(.A1(new_n13895_), .A2(new_n13896_), .ZN(new_n13898_));
  NOR2_X1    g13804(.A1(new_n13898_), .A2(\a[2] ), .ZN(new_n13899_));
  NOR2_X1    g13805(.A1(new_n13899_), .A2(new_n13897_), .ZN(new_n13900_));
  AOI21_X1   g13806(.A1(new_n13884_), .A2(new_n13892_), .B(new_n13900_), .ZN(new_n13901_));
  OAI22_X1   g13807(.A1(new_n10985_), .A2(new_n9425_), .B1(new_n3456_), .B2(new_n10896_), .ZN(new_n13902_));
  AOI21_X1   g13808(.A1(new_n13902_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n13903_));
  XOR2_X1    g13809(.A1(new_n10984_), .A2(new_n13903_), .Z(new_n13904_));
  OAI21_X1   g13810(.A1(new_n13901_), .A2(new_n13893_), .B(new_n13904_), .ZN(new_n13905_));
  NOR3_X1    g13811(.A1(new_n13901_), .A2(new_n13893_), .A3(new_n13904_), .ZN(new_n13906_));
  NOR2_X1    g13812(.A1(new_n13253_), .A2(new_n13248_), .ZN(new_n13907_));
  AOI21_X1   g13813(.A1(new_n12482_), .A2(new_n12480_), .B(new_n13247_), .ZN(new_n13908_));
  OAI21_X1   g13814(.A1(new_n13907_), .A2(new_n13908_), .B(new_n13252_), .ZN(new_n13909_));
  XOR2_X1    g13815(.A1(new_n13253_), .A2(new_n13247_), .Z(new_n13910_));
  OAI21_X1   g13816(.A1(new_n13910_), .A2(new_n13252_), .B(new_n13909_), .ZN(new_n13911_));
  XNOR2_X1   g13817(.A1(new_n13911_), .A2(new_n13241_), .ZN(new_n13912_));
  OAI21_X1   g13818(.A1(new_n13906_), .A2(new_n13912_), .B(new_n13905_), .ZN(new_n13913_));
  NOR2_X1    g13819(.A1(new_n13255_), .A2(new_n13250_), .ZN(new_n13914_));
  NAND3_X1   g13820(.A1(new_n13272_), .A2(new_n13273_), .A3(new_n13269_), .ZN(new_n13915_));
  OAI21_X1   g13821(.A1(new_n13266_), .A2(new_n13263_), .B(new_n13274_), .ZN(new_n13916_));
  NAND2_X1   g13822(.A1(new_n13916_), .A2(new_n13915_), .ZN(new_n13917_));
  NAND2_X1   g13823(.A1(new_n13270_), .A2(new_n13275_), .ZN(new_n13918_));
  MUX2_X1    g13824(.I0(new_n13917_), .I1(new_n13918_), .S(new_n13914_), .Z(new_n13919_));
  NAND2_X1   g13825(.A1(new_n13913_), .A2(new_n13919_), .ZN(new_n13920_));
  OAI22_X1   g13826(.A1(new_n10606_), .A2(new_n3456_), .B1(new_n9425_), .B2(new_n10901_), .ZN(new_n13921_));
  AOI21_X1   g13827(.A1(new_n12211_), .A2(new_n3411_), .B(new_n13921_), .ZN(new_n13922_));
  XOR2_X1    g13828(.A1(new_n13922_), .A2(\a[2] ), .Z(new_n13923_));
  INV_X1     g13829(.I(new_n13923_), .ZN(new_n13924_));
  OAI21_X1   g13830(.A1(new_n13913_), .A2(new_n13919_), .B(new_n13924_), .ZN(new_n13925_));
  NOR2_X1    g13831(.A1(new_n10599_), .A2(new_n3456_), .ZN(new_n13926_));
  NOR3_X1    g13832(.A1(new_n12577_), .A2(new_n9425_), .A3(new_n13926_), .ZN(new_n13927_));
  NOR3_X1    g13833(.A1(new_n12576_), .A2(new_n3414_), .A3(new_n13927_), .ZN(new_n13928_));
  XOR2_X1    g13834(.A1(new_n13928_), .A2(new_n451_), .Z(new_n13929_));
  AOI21_X1   g13835(.A1(new_n13925_), .A2(new_n13920_), .B(new_n13929_), .ZN(new_n13930_));
  NAND3_X1   g13836(.A1(new_n13925_), .A2(new_n13920_), .A3(new_n13929_), .ZN(new_n13931_));
  INV_X1     g13837(.I(new_n13276_), .ZN(new_n13932_));
  INV_X1     g13838(.I(new_n13285_), .ZN(new_n13933_));
  NAND2_X1   g13839(.A1(new_n13933_), .A2(new_n13286_), .ZN(new_n13934_));
  NOR2_X1    g13840(.A1(new_n13934_), .A2(new_n13932_), .ZN(new_n13935_));
  NOR2_X1    g13841(.A1(new_n13287_), .A2(new_n13285_), .ZN(new_n13936_));
  NOR2_X1    g13842(.A1(new_n13936_), .A2(new_n13276_), .ZN(new_n13937_));
  NOR2_X1    g13843(.A1(new_n13937_), .A2(new_n13935_), .ZN(new_n13938_));
  INV_X1     g13844(.I(new_n13938_), .ZN(new_n13939_));
  AOI21_X1   g13845(.A1(new_n13931_), .A2(new_n13939_), .B(new_n13930_), .ZN(new_n13940_));
  INV_X1     g13846(.I(new_n13304_), .ZN(new_n13941_));
  NAND3_X1   g13847(.A1(new_n13941_), .A2(new_n13300_), .A3(new_n13286_), .ZN(new_n13942_));
  NAND3_X1   g13848(.A1(new_n13942_), .A2(new_n13932_), .A3(new_n13934_), .ZN(new_n13943_));
  NOR3_X1    g13849(.A1(new_n13301_), .A2(new_n13304_), .A3(new_n13287_), .ZN(new_n13944_));
  OAI21_X1   g13850(.A1(new_n13944_), .A2(new_n13936_), .B(new_n13276_), .ZN(new_n13945_));
  AND2_X2    g13851(.A1(new_n13945_), .A2(new_n13943_), .Z(new_n13946_));
  NOR2_X1    g13852(.A1(new_n13940_), .A2(new_n13946_), .ZN(new_n13947_));
  INV_X1     g13853(.I(new_n12596_), .ZN(new_n13948_));
  NAND2_X1   g13854(.A1(new_n13948_), .A2(new_n12598_), .ZN(new_n13949_));
  NAND2_X1   g13855(.A1(new_n12614_), .A2(new_n3455_), .ZN(new_n13950_));
  NOR2_X1    g13856(.A1(new_n12601_), .A2(new_n9425_), .ZN(new_n13951_));
  AOI21_X1   g13857(.A1(new_n13951_), .A2(new_n13950_), .B(new_n3414_), .ZN(new_n13952_));
  NAND2_X1   g13858(.A1(new_n13949_), .A2(new_n13952_), .ZN(new_n13953_));
  XOR2_X1    g13859(.A1(new_n13953_), .A2(\a[2] ), .Z(new_n13954_));
  AOI21_X1   g13860(.A1(new_n13940_), .A2(new_n13946_), .B(new_n13954_), .ZN(new_n13955_));
  NAND2_X1   g13861(.A1(new_n13308_), .A2(new_n13296_), .ZN(new_n13956_));
  INV_X1     g13862(.I(new_n13306_), .ZN(new_n13957_));
  NOR3_X1    g13863(.A1(new_n12958_), .A2(new_n13957_), .A3(new_n13311_), .ZN(new_n13958_));
  OAI21_X1   g13864(.A1(new_n12955_), .A2(new_n12956_), .B(new_n12526_), .ZN(new_n13959_));
  NAND3_X1   g13865(.A1(new_n12953_), .A2(new_n12947_), .A3(new_n12943_), .ZN(new_n13960_));
  NAND2_X1   g13866(.A1(new_n13960_), .A2(new_n13959_), .ZN(new_n13961_));
  AOI21_X1   g13867(.A1(new_n13961_), .A2(new_n13312_), .B(new_n13306_), .ZN(new_n13962_));
  OAI21_X1   g13868(.A1(new_n13958_), .A2(new_n13962_), .B(new_n13956_), .ZN(new_n13963_));
  INV_X1     g13869(.I(new_n13956_), .ZN(new_n13964_));
  NAND3_X1   g13870(.A1(new_n13961_), .A2(new_n13306_), .A3(new_n13312_), .ZN(new_n13965_));
  OAI21_X1   g13871(.A1(new_n12958_), .A2(new_n13311_), .B(new_n13957_), .ZN(new_n13966_));
  NAND3_X1   g13872(.A1(new_n13966_), .A2(new_n13965_), .A3(new_n13964_), .ZN(new_n13967_));
  NAND2_X1   g13873(.A1(new_n13963_), .A2(new_n13967_), .ZN(new_n13968_));
  OAI21_X1   g13874(.A1(new_n13955_), .A2(new_n13947_), .B(new_n13968_), .ZN(new_n13969_));
  NOR3_X1    g13875(.A1(new_n13955_), .A2(new_n13947_), .A3(new_n13968_), .ZN(new_n13970_));
  INV_X1     g13876(.I(new_n12619_), .ZN(new_n13971_));
  NAND2_X1   g13877(.A1(new_n13971_), .A2(new_n12620_), .ZN(new_n13972_));
  NAND2_X1   g13878(.A1(new_n12616_), .A2(new_n3455_), .ZN(new_n13973_));
  NOR2_X1    g13879(.A1(new_n12623_), .A2(new_n9425_), .ZN(new_n13974_));
  AOI21_X1   g13880(.A1(new_n13973_), .A2(new_n13974_), .B(new_n3414_), .ZN(new_n13975_));
  NAND2_X1   g13881(.A1(new_n13972_), .A2(new_n13975_), .ZN(new_n13976_));
  XOR2_X1    g13882(.A1(new_n13976_), .A2(\a[2] ), .Z(new_n13977_));
  OAI21_X1   g13883(.A1(new_n13970_), .A2(new_n13977_), .B(new_n13969_), .ZN(new_n13978_));
  OAI22_X1   g13884(.A1(new_n10913_), .A2(new_n3456_), .B1(new_n12768_), .B2(new_n9425_), .ZN(new_n13979_));
  AOI21_X1   g13885(.A1(new_n13979_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n13980_));
  XOR2_X1    g13886(.A1(new_n12767_), .A2(new_n13980_), .Z(new_n13981_));
  INV_X1     g13887(.I(new_n13981_), .ZN(new_n13982_));
  NAND2_X1   g13888(.A1(new_n13978_), .A2(new_n13982_), .ZN(new_n13983_));
  OR2_X2     g13889(.A1(new_n13314_), .A2(new_n13307_), .Z(new_n13984_));
  NAND2_X1   g13890(.A1(new_n12942_), .A2(new_n13317_), .ZN(new_n13985_));
  OAI21_X1   g13891(.A1(new_n12941_), .A2(new_n12936_), .B(new_n13318_), .ZN(new_n13986_));
  NAND2_X1   g13892(.A1(new_n13985_), .A2(new_n13986_), .ZN(new_n13987_));
  XOR2_X1    g13893(.A1(new_n13987_), .A2(new_n13984_), .Z(new_n13988_));
  OAI21_X1   g13894(.A1(new_n13978_), .A2(new_n13982_), .B(new_n13988_), .ZN(new_n13989_));
  OAI22_X1   g13895(.A1(new_n12890_), .A2(new_n9425_), .B1(new_n10923_), .B2(new_n3456_), .ZN(new_n13990_));
  AOI21_X1   g13896(.A1(new_n13990_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n13991_));
  XOR2_X1    g13897(.A1(new_n12889_), .A2(new_n13991_), .Z(new_n13992_));
  AOI21_X1   g13898(.A1(new_n13989_), .A2(new_n13983_), .B(new_n13992_), .ZN(new_n13993_));
  NAND3_X1   g13899(.A1(new_n13989_), .A2(new_n13983_), .A3(new_n13992_), .ZN(new_n13994_));
  NOR2_X1    g13900(.A1(new_n12933_), .A2(new_n12555_), .ZN(new_n13995_));
  XOR2_X1    g13901(.A1(new_n13995_), .A2(new_n13325_), .Z(new_n13996_));
  XNOR2_X1   g13902(.A1(new_n13996_), .A2(new_n13321_), .ZN(new_n13997_));
  INV_X1     g13903(.I(new_n13997_), .ZN(new_n13998_));
  AOI21_X1   g13904(.A1(new_n13994_), .A2(new_n13998_), .B(new_n13993_), .ZN(new_n13999_));
  OAI22_X1   g13905(.A1(new_n10583_), .A2(new_n3456_), .B1(new_n9425_), .B2(new_n10928_), .ZN(new_n14000_));
  AOI21_X1   g13906(.A1(new_n14000_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n14001_));
  XNOR2_X1   g13907(.A1(new_n13378_), .A2(new_n14001_), .ZN(new_n14002_));
  NOR2_X1    g13908(.A1(new_n13999_), .A2(new_n14002_), .ZN(new_n14003_));
  INV_X1     g13909(.I(new_n13326_), .ZN(new_n14004_));
  INV_X1     g13910(.I(new_n13327_), .ZN(new_n14005_));
  NOR2_X1    g13911(.A1(new_n14004_), .A2(new_n14005_), .ZN(new_n14006_));
  INV_X1     g13912(.I(new_n13330_), .ZN(new_n14007_));
  INV_X1     g13913(.I(new_n13338_), .ZN(new_n14008_));
  NAND3_X1   g13914(.A1(new_n14008_), .A2(new_n14007_), .A3(new_n13339_), .ZN(new_n14009_));
  OAI21_X1   g13915(.A1(new_n13340_), .A2(new_n13338_), .B(new_n13330_), .ZN(new_n14010_));
  NAND2_X1   g13916(.A1(new_n14009_), .A2(new_n14010_), .ZN(new_n14011_));
  XOR2_X1    g13917(.A1(new_n14011_), .A2(new_n14006_), .Z(new_n14012_));
  AOI21_X1   g13918(.A1(new_n13999_), .A2(new_n14002_), .B(new_n14012_), .ZN(new_n14013_));
  INV_X1     g13919(.I(new_n13394_), .ZN(new_n14014_));
  NAND2_X1   g13920(.A1(new_n10937_), .A2(new_n3455_), .ZN(new_n14015_));
  NOR2_X1    g13921(.A1(new_n13395_), .A2(new_n9425_), .ZN(new_n14016_));
  AOI21_X1   g13922(.A1(new_n14016_), .A2(new_n14015_), .B(new_n3414_), .ZN(new_n14017_));
  NAND2_X1   g13923(.A1(new_n14014_), .A2(new_n14017_), .ZN(new_n14018_));
  XOR2_X1    g13924(.A1(new_n14018_), .A2(\a[2] ), .Z(new_n14019_));
  INV_X1     g13925(.I(new_n14019_), .ZN(new_n14020_));
  OAI21_X1   g13926(.A1(new_n14013_), .A2(new_n14003_), .B(new_n14020_), .ZN(new_n14021_));
  NOR3_X1    g13927(.A1(new_n14013_), .A2(new_n14003_), .A3(new_n14020_), .ZN(new_n14022_));
  XNOR2_X1   g13928(.A1(new_n13551_), .A2(new_n13550_), .ZN(new_n14023_));
  OAI21_X1   g13929(.A1(new_n14022_), .A2(new_n14023_), .B(new_n14021_), .ZN(new_n14024_));
  NAND3_X1   g13930(.A1(new_n13359_), .A2(new_n13355_), .A3(new_n13345_), .ZN(new_n14025_));
  AND3_X2    g13931(.A1(new_n13344_), .A2(new_n13550_), .A3(new_n14025_), .Z(new_n14026_));
  AOI21_X1   g13932(.A1(new_n13344_), .A2(new_n14025_), .B(new_n13550_), .ZN(new_n14027_));
  NOR2_X1    g13933(.A1(new_n14026_), .A2(new_n14027_), .ZN(new_n14028_));
  INV_X1     g13934(.I(new_n14028_), .ZN(new_n14029_));
  NAND2_X1   g13935(.A1(new_n14024_), .A2(new_n14029_), .ZN(new_n14030_));
  NAND2_X1   g13936(.A1(new_n10949_), .A2(new_n3455_), .ZN(new_n14031_));
  NOR2_X1    g13937(.A1(new_n12908_), .A2(new_n9425_), .ZN(new_n14032_));
  AOI21_X1   g13938(.A1(new_n14032_), .A2(new_n14031_), .B(new_n3414_), .ZN(new_n14033_));
  NAND2_X1   g13939(.A1(new_n12907_), .A2(new_n14033_), .ZN(new_n14034_));
  XOR2_X1    g13940(.A1(new_n14034_), .A2(\a[2] ), .Z(new_n14035_));
  INV_X1     g13941(.I(new_n14035_), .ZN(new_n14036_));
  OAI21_X1   g13942(.A1(new_n14024_), .A2(new_n14029_), .B(new_n14036_), .ZN(new_n14037_));
  OAI22_X1   g13943(.A1(new_n9405_), .A2(new_n10952_), .B1(new_n10938_), .B2(new_n9408_), .ZN(new_n14038_));
  OAI21_X1   g13944(.A1(new_n10577_), .A2(new_n3456_), .B(new_n14038_), .ZN(new_n14039_));
  AOI21_X1   g13945(.A1(new_n14039_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n14040_));
  XOR2_X1    g13946(.A1(new_n13544_), .A2(new_n14040_), .Z(new_n14041_));
  AOI21_X1   g13947(.A1(new_n14037_), .A2(new_n14030_), .B(new_n14041_), .ZN(new_n14042_));
  NAND3_X1   g13948(.A1(new_n14037_), .A2(new_n14030_), .A3(new_n14041_), .ZN(new_n14043_));
  NOR2_X1    g13949(.A1(new_n13555_), .A2(new_n13362_), .ZN(new_n14044_));
  NAND2_X1   g13950(.A1(new_n13383_), .A2(new_n13385_), .ZN(new_n14045_));
  XNOR2_X1   g13951(.A1(new_n14044_), .A2(new_n14045_), .ZN(new_n14046_));
  INV_X1     g13952(.I(new_n14046_), .ZN(new_n14047_));
  AOI21_X1   g13953(.A1(new_n14043_), .A2(new_n14047_), .B(new_n14042_), .ZN(new_n14048_));
  NOR2_X1    g13954(.A1(new_n10963_), .A2(new_n10965_), .ZN(new_n14049_));
  NOR2_X1    g13955(.A1(new_n10956_), .A2(new_n14049_), .ZN(new_n14050_));
  XOR2_X1    g13956(.A1(new_n10577_), .A2(new_n10962_), .Z(new_n14051_));
  NOR2_X1    g13957(.A1(new_n10957_), .A2(new_n14051_), .ZN(new_n14052_));
  NOR2_X1    g13958(.A1(new_n14052_), .A2(new_n14050_), .ZN(new_n14053_));
  NOR2_X1    g13959(.A1(new_n10577_), .A2(new_n10952_), .ZN(new_n14054_));
  OAI22_X1   g13960(.A1(new_n14054_), .A2(new_n9425_), .B1(new_n3456_), .B2(new_n10961_), .ZN(new_n14055_));
  AOI21_X1   g13961(.A1(new_n14055_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n14056_));
  XOR2_X1    g13962(.A1(new_n14053_), .A2(new_n14056_), .Z(new_n14057_));
  NOR2_X1    g13963(.A1(new_n14048_), .A2(new_n14057_), .ZN(new_n14058_));
  NOR2_X1    g13964(.A1(new_n13557_), .A2(new_n13558_), .ZN(new_n14059_));
  NAND2_X1   g13965(.A1(new_n13399_), .A2(new_n13402_), .ZN(new_n14060_));
  XOR2_X1    g13966(.A1(new_n14059_), .A2(new_n14060_), .Z(new_n14061_));
  AOI21_X1   g13967(.A1(new_n14048_), .A2(new_n14057_), .B(new_n14061_), .ZN(new_n14062_));
  NAND3_X1   g13968(.A1(new_n12915_), .A2(new_n13403_), .A3(new_n13399_), .ZN(new_n14063_));
  NAND3_X1   g13969(.A1(new_n14059_), .A2(new_n14063_), .A3(new_n14060_), .ZN(new_n14064_));
  INV_X1     g13970(.I(new_n14059_), .ZN(new_n14065_));
  NAND2_X1   g13971(.A1(new_n14063_), .A2(new_n14060_), .ZN(new_n14066_));
  NAND2_X1   g13972(.A1(new_n14066_), .A2(new_n14065_), .ZN(new_n14067_));
  NAND2_X1   g13973(.A1(new_n14067_), .A2(new_n14064_), .ZN(new_n14068_));
  AOI21_X1   g13974(.A1(new_n13565_), .A2(new_n13564_), .B(new_n12914_), .ZN(new_n14069_));
  NOR3_X1    g13975(.A1(new_n13549_), .A2(new_n12915_), .A3(new_n13562_), .ZN(new_n14070_));
  NOR3_X1    g13976(.A1(new_n14069_), .A2(new_n14070_), .A3(new_n10980_), .ZN(new_n14071_));
  NOR3_X1    g13977(.A1(new_n14071_), .A2(new_n13567_), .A3(new_n14068_), .ZN(new_n14072_));
  INV_X1     g13978(.I(new_n14051_), .ZN(new_n14073_));
  NOR2_X1    g13979(.A1(new_n10962_), .A2(new_n10570_), .ZN(new_n14074_));
  NOR2_X1    g13980(.A1(new_n10571_), .A2(new_n10961_), .ZN(new_n14075_));
  OAI21_X1   g13981(.A1(new_n14074_), .A2(new_n14075_), .B(new_n14073_), .ZN(new_n14076_));
  XOR2_X1    g13982(.A1(new_n10956_), .A2(new_n14076_), .Z(new_n14077_));
  OAI22_X1   g13983(.A1(new_n10965_), .A2(new_n9425_), .B1(new_n3456_), .B2(new_n10570_), .ZN(new_n14078_));
  AOI21_X1   g13984(.A1(new_n14078_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n14079_));
  XNOR2_X1   g13985(.A1(new_n14077_), .A2(new_n14079_), .ZN(new_n14080_));
  OAI21_X1   g13986(.A1(new_n14071_), .A2(new_n13567_), .B(new_n14068_), .ZN(new_n14081_));
  AOI21_X1   g13987(.A1(new_n14080_), .A2(new_n14081_), .B(new_n14072_), .ZN(new_n14082_));
  OAI21_X1   g13988(.A1(new_n14062_), .A2(new_n14058_), .B(new_n14082_), .ZN(new_n14083_));
  NOR2_X1    g13989(.A1(new_n13560_), .A2(new_n13535_), .ZN(new_n14084_));
  INV_X1     g13990(.I(new_n13548_), .ZN(new_n14085_));
  NAND2_X1   g13991(.A1(new_n12914_), .A2(new_n14085_), .ZN(new_n14086_));
  AOI21_X1   g13992(.A1(new_n13560_), .A2(new_n13535_), .B(new_n14086_), .ZN(new_n14087_));
  NOR2_X1    g13993(.A1(new_n14087_), .A2(new_n14084_), .ZN(new_n14088_));
  NAND2_X1   g13994(.A1(new_n13522_), .A2(new_n12899_), .ZN(new_n14089_));
  NAND3_X1   g13995(.A1(new_n13518_), .A2(new_n13521_), .A3(new_n13531_), .ZN(new_n14090_));
  NAND3_X1   g13996(.A1(new_n14090_), .A2(new_n13410_), .A3(new_n13526_), .ZN(new_n14091_));
  NAND2_X1   g13997(.A1(new_n14091_), .A2(new_n14089_), .ZN(new_n14092_));
  AOI21_X1   g13998(.A1(new_n13494_), .A2(new_n13497_), .B(new_n12865_), .ZN(new_n14093_));
  AOI21_X1   g13999(.A1(new_n13496_), .A2(new_n13495_), .B(new_n12854_), .ZN(new_n14094_));
  NOR3_X1    g14000(.A1(new_n13488_), .A2(new_n13493_), .A3(new_n12845_), .ZN(new_n14095_));
  NOR3_X1    g14001(.A1(new_n14094_), .A2(new_n14095_), .A3(new_n12870_), .ZN(new_n14096_));
  NOR3_X1    g14002(.A1(new_n13414_), .A2(new_n14096_), .A3(new_n13500_), .ZN(new_n14097_));
  NAND2_X1   g14003(.A1(new_n13474_), .A2(new_n12837_), .ZN(new_n14098_));
  AOI21_X1   g14004(.A1(new_n13468_), .A2(new_n13479_), .B(new_n13471_), .ZN(new_n14099_));
  NAND3_X1   g14005(.A1(new_n12782_), .A2(new_n14099_), .A3(new_n12838_), .ZN(new_n14100_));
  NAND2_X1   g14006(.A1(new_n14100_), .A2(new_n14098_), .ZN(new_n14101_));
  INV_X1     g14007(.I(new_n13464_), .ZN(new_n14102_));
  OAI21_X1   g14008(.A1(new_n13418_), .A2(new_n14102_), .B(new_n13466_), .ZN(new_n14103_));
  AOI22_X1   g14009(.A1(new_n247_), .A2(new_n10843_), .B1(new_n11608_), .B2(new_n5783_), .ZN(new_n14104_));
  OAI21_X1   g14010(.A1(new_n14104_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n14105_));
  XOR2_X1    g14011(.A1(new_n11607_), .A2(new_n14105_), .Z(new_n14106_));
  INV_X1     g14012(.I(new_n14106_), .ZN(new_n14107_));
  INV_X1     g14013(.I(new_n13423_), .ZN(new_n14108_));
  AOI21_X1   g14014(.A1(new_n14108_), .A2(new_n13443_), .B(new_n13448_), .ZN(new_n14109_));
  NAND2_X1   g14015(.A1(new_n13426_), .A2(new_n14109_), .ZN(new_n14110_));
  OAI21_X1   g14016(.A1(new_n14108_), .A2(new_n13443_), .B(new_n14110_), .ZN(new_n14111_));
  NOR2_X1    g14017(.A1(new_n13427_), .A2(new_n13440_), .ZN(new_n14112_));
  NOR2_X1    g14018(.A1(new_n14112_), .A2(new_n13441_), .ZN(new_n14113_));
  OAI22_X1   g14019(.A1(new_n10672_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10792_), .ZN(new_n14114_));
  OAI21_X1   g14020(.A1(new_n79_), .A2(new_n10658_), .B(new_n14114_), .ZN(new_n14115_));
  AOI21_X1   g14021(.A1(new_n14115_), .A2(new_n72_), .B(new_n79_), .ZN(new_n14116_));
  XOR2_X1    g14022(.A1(new_n11175_), .A2(new_n14116_), .Z(new_n14117_));
  NAND3_X1   g14023(.A1(new_n13432_), .A2(new_n11046_), .A3(new_n13435_), .ZN(new_n14118_));
  NAND2_X1   g14024(.A1(new_n10794_), .A2(new_n962_), .ZN(new_n14119_));
  AOI22_X1   g14025(.A1(new_n10809_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n10745_), .ZN(new_n14120_));
  AOI21_X1   g14026(.A1(new_n14119_), .A2(new_n14120_), .B(new_n82_), .ZN(new_n14121_));
  NAND2_X1   g14027(.A1(new_n11064_), .A2(new_n14121_), .ZN(new_n14122_));
  XNOR2_X1   g14028(.A1(new_n14118_), .A2(new_n14122_), .ZN(new_n14123_));
  INV_X1     g14029(.I(new_n14123_), .ZN(new_n14124_));
  XOR2_X1    g14030(.A1(new_n14117_), .A2(new_n14124_), .Z(new_n14125_));
  NOR2_X1    g14031(.A1(new_n14113_), .A2(new_n14125_), .ZN(new_n14126_));
  INV_X1     g14032(.I(new_n14113_), .ZN(new_n14127_));
  AND2_X2    g14033(.A1(new_n14117_), .A2(new_n14123_), .Z(new_n14128_));
  NOR2_X1    g14034(.A1(new_n14117_), .A2(new_n14123_), .ZN(new_n14129_));
  NOR2_X1    g14035(.A1(new_n14128_), .A2(new_n14129_), .ZN(new_n14130_));
  NOR2_X1    g14036(.A1(new_n14127_), .A2(new_n14130_), .ZN(new_n14131_));
  NOR2_X1    g14037(.A1(new_n14131_), .A2(new_n14126_), .ZN(new_n14132_));
  OAI22_X1   g14038(.A1(new_n10646_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n11214_), .ZN(new_n14133_));
  OAI21_X1   g14039(.A1(new_n1128_), .A2(new_n11264_), .B(new_n14133_), .ZN(new_n14134_));
  AOI21_X1   g14040(.A1(new_n14134_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n14135_));
  XNOR2_X1   g14041(.A1(new_n11268_), .A2(new_n14135_), .ZN(new_n14136_));
  XNOR2_X1   g14042(.A1(new_n14132_), .A2(new_n14136_), .ZN(new_n14137_));
  INV_X1     g14043(.I(new_n14137_), .ZN(new_n14138_));
  NAND2_X1   g14044(.A1(new_n14111_), .A2(new_n14138_), .ZN(new_n14139_));
  INV_X1     g14045(.I(new_n14132_), .ZN(new_n14140_));
  INV_X1     g14046(.I(new_n14136_), .ZN(new_n14141_));
  NOR2_X1    g14047(.A1(new_n14140_), .A2(new_n14141_), .ZN(new_n14142_));
  NOR2_X1    g14048(.A1(new_n14132_), .A2(new_n14136_), .ZN(new_n14143_));
  NOR2_X1    g14049(.A1(new_n14142_), .A2(new_n14143_), .ZN(new_n14144_));
  NOR2_X1    g14050(.A1(new_n14111_), .A2(new_n14144_), .ZN(new_n14145_));
  INV_X1     g14051(.I(new_n14145_), .ZN(new_n14146_));
  NAND2_X1   g14052(.A1(new_n14146_), .A2(new_n14139_), .ZN(new_n14147_));
  XOR2_X1    g14053(.A1(new_n14147_), .A2(new_n14107_), .Z(new_n14148_));
  NAND2_X1   g14054(.A1(new_n14148_), .A2(new_n14103_), .ZN(new_n14149_));
  AOI21_X1   g14055(.A1(new_n13463_), .A2(new_n13455_), .B(new_n13422_), .ZN(new_n14150_));
  AOI21_X1   g14056(.A1(new_n13462_), .A2(new_n13464_), .B(new_n14150_), .ZN(new_n14151_));
  NAND3_X1   g14057(.A1(new_n14146_), .A2(new_n14106_), .A3(new_n14139_), .ZN(new_n14152_));
  INV_X1     g14058(.I(new_n14152_), .ZN(new_n14153_));
  AOI21_X1   g14059(.A1(new_n14146_), .A2(new_n14139_), .B(new_n14106_), .ZN(new_n14154_));
  OAI21_X1   g14060(.A1(new_n14153_), .A2(new_n14154_), .B(new_n14151_), .ZN(new_n14155_));
  AOI22_X1   g14061(.A1(new_n11724_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n10875_), .ZN(new_n14156_));
  OAI21_X1   g14062(.A1(new_n14156_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n14157_));
  XNOR2_X1   g14063(.A1(new_n11722_), .A2(new_n14157_), .ZN(new_n14158_));
  INV_X1     g14064(.I(new_n14158_), .ZN(new_n14159_));
  AOI21_X1   g14065(.A1(new_n14149_), .A2(new_n14155_), .B(new_n14159_), .ZN(new_n14160_));
  NAND2_X1   g14066(.A1(new_n14149_), .A2(new_n14155_), .ZN(new_n14161_));
  NOR2_X1    g14067(.A1(new_n14161_), .A2(new_n14158_), .ZN(new_n14162_));
  OAI21_X1   g14068(.A1(new_n14160_), .A2(new_n14162_), .B(new_n14101_), .ZN(new_n14163_));
  INV_X1     g14069(.I(new_n14163_), .ZN(new_n14164_));
  NAND3_X1   g14070(.A1(new_n14149_), .A2(new_n14155_), .A3(new_n14158_), .ZN(new_n14165_));
  NAND2_X1   g14071(.A1(new_n14161_), .A2(new_n14159_), .ZN(new_n14166_));
  AOI21_X1   g14072(.A1(new_n14165_), .A2(new_n14166_), .B(new_n14101_), .ZN(new_n14167_));
  OAI22_X1   g14073(.A1(new_n12091_), .A2(new_n5420_), .B1(new_n1620_), .B2(new_n10611_), .ZN(new_n14168_));
  AOI21_X1   g14074(.A1(new_n14168_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n14169_));
  XOR2_X1    g14075(.A1(new_n12090_), .A2(new_n14169_), .Z(new_n14170_));
  INV_X1     g14076(.I(new_n14170_), .ZN(new_n14171_));
  NOR3_X1    g14077(.A1(new_n14164_), .A2(new_n14171_), .A3(new_n14167_), .ZN(new_n14172_));
  INV_X1     g14078(.I(new_n14167_), .ZN(new_n14173_));
  AOI21_X1   g14079(.A1(new_n14173_), .A2(new_n14163_), .B(new_n14170_), .ZN(new_n14174_));
  NOR2_X1    g14080(.A1(new_n14174_), .A2(new_n14172_), .ZN(new_n14175_));
  NOR2_X1    g14081(.A1(new_n13482_), .A2(new_n13478_), .ZN(new_n14176_));
  NAND3_X1   g14082(.A1(new_n13490_), .A2(new_n13491_), .A3(new_n12845_), .ZN(new_n14177_));
  NAND2_X1   g14083(.A1(new_n14177_), .A2(new_n13486_), .ZN(new_n14178_));
  OAI22_X1   g14084(.A1(new_n14178_), .A2(new_n13489_), .B1(new_n12845_), .B2(new_n14176_), .ZN(new_n14179_));
  NAND2_X1   g14085(.A1(new_n14175_), .A2(new_n14179_), .ZN(new_n14180_));
  NAND3_X1   g14086(.A1(new_n14173_), .A2(new_n14163_), .A3(new_n14170_), .ZN(new_n14181_));
  OAI21_X1   g14087(.A1(new_n14164_), .A2(new_n14167_), .B(new_n14171_), .ZN(new_n14182_));
  NAND2_X1   g14088(.A1(new_n14182_), .A2(new_n14181_), .ZN(new_n14183_));
  NOR2_X1    g14089(.A1(new_n14176_), .A2(new_n12845_), .ZN(new_n14184_));
  NOR2_X1    g14090(.A1(new_n14178_), .A2(new_n13489_), .ZN(new_n14185_));
  NOR2_X1    g14091(.A1(new_n14185_), .A2(new_n14184_), .ZN(new_n14186_));
  NAND2_X1   g14092(.A1(new_n14186_), .A2(new_n14183_), .ZN(new_n14187_));
  INV_X1     g14093(.I(new_n12576_), .ZN(new_n14188_));
  AOI22_X1   g14094(.A1(new_n12578_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n10600_), .ZN(new_n14189_));
  OAI21_X1   g14095(.A1(new_n14189_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n14190_));
  NOR2_X1    g14096(.A1(new_n14188_), .A2(new_n14190_), .ZN(new_n14191_));
  INV_X1     g14097(.I(new_n14190_), .ZN(new_n14192_));
  NOR2_X1    g14098(.A1(new_n12576_), .A2(new_n14192_), .ZN(new_n14193_));
  NOR2_X1    g14099(.A1(new_n14191_), .A2(new_n14193_), .ZN(new_n14194_));
  INV_X1     g14100(.I(new_n14194_), .ZN(new_n14195_));
  AOI21_X1   g14101(.A1(new_n14187_), .A2(new_n14180_), .B(new_n14195_), .ZN(new_n14196_));
  NOR2_X1    g14102(.A1(new_n14186_), .A2(new_n14183_), .ZN(new_n14197_));
  NOR2_X1    g14103(.A1(new_n14175_), .A2(new_n14179_), .ZN(new_n14198_));
  NOR3_X1    g14104(.A1(new_n14197_), .A2(new_n14198_), .A3(new_n14194_), .ZN(new_n14199_));
  OAI22_X1   g14105(.A1(new_n14097_), .A2(new_n14093_), .B1(new_n14199_), .B2(new_n14196_), .ZN(new_n14200_));
  NOR2_X1    g14106(.A1(new_n14097_), .A2(new_n14093_), .ZN(new_n14201_));
  NAND3_X1   g14107(.A1(new_n14187_), .A2(new_n14180_), .A3(new_n14194_), .ZN(new_n14202_));
  OAI21_X1   g14108(.A1(new_n14197_), .A2(new_n14198_), .B(new_n14195_), .ZN(new_n14203_));
  NAND2_X1   g14109(.A1(new_n14203_), .A2(new_n14202_), .ZN(new_n14204_));
  NAND2_X1   g14110(.A1(new_n14201_), .A2(new_n14204_), .ZN(new_n14205_));
  OAI22_X1   g14111(.A1(new_n10913_), .A2(new_n1078_), .B1(new_n12768_), .B2(new_n6757_), .ZN(new_n14206_));
  AOI21_X1   g14112(.A1(new_n14206_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n14207_));
  XOR2_X1    g14113(.A1(new_n12767_), .A2(new_n14207_), .Z(new_n14208_));
  NAND3_X1   g14114(.A1(new_n14205_), .A2(new_n14200_), .A3(new_n14208_), .ZN(new_n14209_));
  AOI21_X1   g14115(.A1(new_n14205_), .A2(new_n14200_), .B(new_n14208_), .ZN(new_n14210_));
  INV_X1     g14116(.I(new_n14210_), .ZN(new_n14211_));
  NAND2_X1   g14117(.A1(new_n14211_), .A2(new_n14209_), .ZN(new_n14212_));
  AOI21_X1   g14118(.A1(new_n13505_), .A2(new_n13508_), .B(new_n12882_), .ZN(new_n14213_));
  AOI21_X1   g14119(.A1(new_n13507_), .A2(new_n13502_), .B(new_n12870_), .ZN(new_n14214_));
  NOR3_X1    g14120(.A1(new_n13503_), .A2(new_n12865_), .A3(new_n13504_), .ZN(new_n14215_));
  NOR3_X1    g14121(.A1(new_n14215_), .A2(new_n14214_), .A3(new_n12877_), .ZN(new_n14216_));
  NOR2_X1    g14122(.A1(new_n14216_), .A2(new_n13512_), .ZN(new_n14217_));
  AOI21_X1   g14123(.A1(new_n14217_), .A2(new_n13413_), .B(new_n14213_), .ZN(new_n14218_));
  NOR2_X1    g14124(.A1(new_n14218_), .A2(new_n14212_), .ZN(new_n14219_));
  INV_X1     g14125(.I(new_n14209_), .ZN(new_n14220_));
  NOR2_X1    g14126(.A1(new_n14220_), .A2(new_n14210_), .ZN(new_n14221_));
  NAND2_X1   g14127(.A1(new_n13509_), .A2(new_n12877_), .ZN(new_n14222_));
  OAI21_X1   g14128(.A1(new_n13509_), .A2(new_n12877_), .B(new_n13513_), .ZN(new_n14223_));
  OAI21_X1   g14129(.A1(new_n14223_), .A2(new_n13516_), .B(new_n14222_), .ZN(new_n14224_));
  NOR2_X1    g14130(.A1(new_n14224_), .A2(new_n14221_), .ZN(new_n14225_));
  OAI22_X1   g14131(.A1(new_n13395_), .A2(new_n7837_), .B1(new_n2495_), .B2(new_n10938_), .ZN(new_n14226_));
  AOI21_X1   g14132(.A1(new_n14226_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n14227_));
  XOR2_X1    g14133(.A1(new_n13394_), .A2(new_n14227_), .Z(new_n14228_));
  NOR3_X1    g14134(.A1(new_n14219_), .A2(new_n14225_), .A3(new_n14228_), .ZN(new_n14229_));
  INV_X1     g14135(.I(new_n14229_), .ZN(new_n14230_));
  OAI21_X1   g14136(.A1(new_n14219_), .A2(new_n14225_), .B(new_n14228_), .ZN(new_n14231_));
  NAND2_X1   g14137(.A1(new_n14230_), .A2(new_n14231_), .ZN(new_n14232_));
  NOR2_X1    g14138(.A1(new_n14092_), .A2(new_n14232_), .ZN(new_n14233_));
  NAND2_X1   g14139(.A1(new_n14092_), .A2(new_n14232_), .ZN(new_n14234_));
  INV_X1     g14140(.I(new_n14234_), .ZN(new_n14235_));
  OAI22_X1   g14141(.A1(new_n14054_), .A2(new_n8831_), .B1(new_n3040_), .B2(new_n10961_), .ZN(new_n14236_));
  AOI21_X1   g14142(.A1(new_n14236_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n14237_));
  XOR2_X1    g14143(.A1(new_n14053_), .A2(new_n14237_), .Z(new_n14238_));
  INV_X1     g14144(.I(new_n14238_), .ZN(new_n14239_));
  NOR3_X1    g14145(.A1(new_n14235_), .A2(new_n14233_), .A3(new_n14239_), .ZN(new_n14240_));
  INV_X1     g14146(.I(new_n14233_), .ZN(new_n14241_));
  AOI21_X1   g14147(.A1(new_n14241_), .A2(new_n14234_), .B(new_n14238_), .ZN(new_n14242_));
  NOR2_X1    g14148(.A1(new_n14242_), .A2(new_n14240_), .ZN(new_n14243_));
  INV_X1     g14149(.I(new_n14243_), .ZN(new_n14244_));
  XOR2_X1    g14150(.A1(new_n14088_), .A2(new_n14244_), .Z(new_n14245_));
  AOI21_X1   g14151(.A1(new_n10564_), .A2(new_n10974_), .B(new_n10972_), .ZN(new_n14246_));
  INV_X1     g14152(.I(new_n14246_), .ZN(new_n14247_));
  INV_X1     g14153(.I(new_n10556_), .ZN(new_n14248_));
  OAI22_X1   g14154(.A1(new_n4649_), .A2(new_n14248_), .B1(new_n4644_), .B2(new_n10557_), .ZN(new_n14249_));
  OAI22_X1   g14155(.A1(new_n10529_), .A2(new_n14249_), .B1(new_n4648_), .B2(new_n10556_), .ZN(new_n14250_));
  INV_X1     g14156(.I(new_n10552_), .ZN(new_n14251_));
  AOI21_X1   g14157(.A1(new_n10551_), .A2(new_n14251_), .B(new_n10553_), .ZN(new_n14252_));
  NOR3_X1    g14158(.A1(new_n4564_), .A2(new_n79_), .A3(new_n4570_), .ZN(new_n14253_));
  OAI21_X1   g14159(.A1(new_n14253_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n14254_));
  XOR2_X1    g14160(.A1(new_n4610_), .A2(new_n14254_), .Z(new_n14255_));
  NOR2_X1    g14161(.A1(new_n4516_), .A2(new_n92_), .ZN(new_n14256_));
  INV_X1     g14162(.I(new_n14256_), .ZN(new_n14257_));
  NOR2_X1    g14163(.A1(new_n4564_), .A2(new_n511_), .ZN(new_n14258_));
  AOI21_X1   g14164(.A1(new_n87_), .A2(new_n4564_), .B(new_n14258_), .ZN(new_n14259_));
  AOI21_X1   g14165(.A1(new_n14257_), .A2(new_n14259_), .B(new_n82_), .ZN(new_n14260_));
  OAI21_X1   g14166(.A1(new_n4593_), .A2(new_n4591_), .B(new_n14260_), .ZN(new_n14261_));
  INV_X1     g14167(.I(new_n14261_), .ZN(new_n14262_));
  NAND2_X1   g14168(.A1(new_n10544_), .A2(new_n4633_), .ZN(new_n14263_));
  NAND2_X1   g14169(.A1(new_n14263_), .A2(new_n10543_), .ZN(new_n14264_));
  XOR2_X1    g14170(.A1(new_n14264_), .A2(new_n14262_), .Z(new_n14265_));
  NOR2_X1    g14171(.A1(new_n14264_), .A2(new_n14261_), .ZN(new_n14266_));
  NAND2_X1   g14172(.A1(new_n14264_), .A2(new_n14261_), .ZN(new_n14267_));
  INV_X1     g14173(.I(new_n14267_), .ZN(new_n14268_));
  OAI21_X1   g14174(.A1(new_n14268_), .A2(new_n14266_), .B(new_n14255_), .ZN(new_n14269_));
  OAI21_X1   g14175(.A1(new_n14255_), .A2(new_n14265_), .B(new_n14269_), .ZN(new_n14270_));
  XOR2_X1    g14176(.A1(new_n14252_), .A2(new_n14270_), .Z(new_n14271_));
  NAND2_X1   g14177(.A1(new_n14250_), .A2(new_n14271_), .ZN(new_n14272_));
  XOR2_X1    g14178(.A1(new_n14252_), .A2(new_n14270_), .Z(new_n14273_));
  OAI21_X1   g14179(.A1(new_n14250_), .A2(new_n14273_), .B(new_n14272_), .ZN(new_n14274_));
  NOR2_X1    g14180(.A1(new_n10971_), .A2(new_n14274_), .ZN(new_n14275_));
  INV_X1     g14181(.I(new_n14274_), .ZN(new_n14276_));
  NOR2_X1    g14182(.A1(new_n10564_), .A2(new_n14276_), .ZN(new_n14277_));
  OAI21_X1   g14183(.A1(new_n14275_), .A2(new_n14277_), .B(new_n14247_), .ZN(new_n14278_));
  XOR2_X1    g14184(.A1(new_n10564_), .A2(new_n14274_), .Z(new_n14279_));
  OAI21_X1   g14185(.A1(new_n14247_), .A2(new_n14279_), .B(new_n14278_), .ZN(new_n14280_));
  NAND2_X1   g14186(.A1(new_n10971_), .A2(new_n10571_), .ZN(new_n14281_));
  AOI22_X1   g14187(.A1(new_n14281_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n14274_), .ZN(new_n14282_));
  OAI21_X1   g14188(.A1(new_n14282_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n14283_));
  XOR2_X1    g14189(.A1(new_n14280_), .A2(new_n14283_), .Z(new_n14284_));
  NOR2_X1    g14190(.A1(new_n14245_), .A2(new_n14284_), .ZN(new_n14285_));
  NAND2_X1   g14191(.A1(new_n14083_), .A2(new_n14285_), .ZN(new_n14286_));
  AOI21_X1   g14192(.A1(new_n13070_), .A2(new_n13067_), .B(new_n13585_), .ZN(new_n14287_));
  AOI21_X1   g14193(.A1(new_n13585_), .A2(new_n13588_), .B(new_n14287_), .ZN(new_n14288_));
  NAND3_X1   g14194(.A1(new_n13582_), .A2(new_n13594_), .A3(new_n13595_), .ZN(new_n14289_));
  OAI21_X1   g14195(.A1(new_n13040_), .A2(new_n13042_), .B(new_n13054_), .ZN(new_n14290_));
  NAND2_X1   g14196(.A1(new_n14290_), .A2(new_n14289_), .ZN(new_n14291_));
  INV_X1     g14197(.I(new_n13051_), .ZN(new_n14292_));
  INV_X1     g14198(.I(new_n13601_), .ZN(new_n14293_));
  NOR2_X1    g14199(.A1(new_n11009_), .A2(new_n11002_), .ZN(new_n14294_));
  AOI21_X1   g14200(.A1(new_n10780_), .A2(new_n10783_), .B(new_n10762_), .ZN(new_n14295_));
  OAI21_X1   g14201(.A1(new_n14294_), .A2(new_n14295_), .B(new_n3413_), .ZN(new_n14296_));
  AOI21_X1   g14202(.A1(new_n11030_), .A2(new_n3413_), .B(new_n13608_), .ZN(new_n14297_));
  NAND3_X1   g14203(.A1(new_n14297_), .A2(new_n14293_), .A3(new_n14296_), .ZN(new_n14298_));
  NOR2_X1    g14204(.A1(new_n14298_), .A2(new_n14292_), .ZN(new_n14299_));
  OAI21_X1   g14205(.A1(new_n11188_), .A2(new_n13617_), .B(\a[2] ), .ZN(new_n14300_));
  NAND3_X1   g14206(.A1(new_n11001_), .A2(new_n13614_), .A3(new_n451_), .ZN(new_n14301_));
  AOI22_X1   g14207(.A1(new_n14300_), .A2(new_n14301_), .B1(new_n14298_), .B2(new_n14292_), .ZN(new_n14302_));
  NOR2_X1    g14208(.A1(new_n14302_), .A2(new_n14299_), .ZN(new_n14303_));
  NOR3_X1    g14209(.A1(new_n13628_), .A2(new_n13625_), .A3(new_n13632_), .ZN(new_n14304_));
  AOI21_X1   g14210(.A1(new_n11045_), .A2(new_n11039_), .B(new_n13623_), .ZN(new_n14305_));
  NOR2_X1    g14211(.A1(new_n14305_), .A2(new_n14304_), .ZN(new_n14306_));
  NOR2_X1    g14212(.A1(new_n14306_), .A2(new_n14303_), .ZN(new_n14307_));
  NOR2_X1    g14213(.A1(new_n13581_), .A2(new_n13052_), .ZN(new_n14308_));
  NOR2_X1    g14214(.A1(new_n14308_), .A2(new_n13054_), .ZN(new_n14309_));
  AOI21_X1   g14215(.A1(new_n14306_), .A2(new_n14303_), .B(new_n14309_), .ZN(new_n14310_));
  NOR3_X1    g14216(.A1(new_n14310_), .A2(new_n14307_), .A3(new_n14291_), .ZN(new_n14311_));
  AOI21_X1   g14217(.A1(new_n11064_), .A2(new_n13646_), .B(new_n451_), .ZN(new_n14312_));
  NOR3_X1    g14218(.A1(new_n13643_), .A2(new_n13647_), .A3(\a[2] ), .ZN(new_n14313_));
  NOR2_X1    g14219(.A1(new_n14313_), .A2(new_n14312_), .ZN(new_n14314_));
  NOR2_X1    g14220(.A1(new_n14311_), .A2(new_n14314_), .ZN(new_n14315_));
  NAND3_X1   g14221(.A1(new_n11332_), .A2(new_n11331_), .A3(new_n13656_), .ZN(new_n14316_));
  OAI21_X1   g14222(.A1(new_n11135_), .A2(new_n11139_), .B(new_n13653_), .ZN(new_n14317_));
  NAND2_X1   g14223(.A1(new_n14317_), .A2(new_n14316_), .ZN(new_n14318_));
  OAI21_X1   g14224(.A1(new_n14315_), .A2(new_n13639_), .B(new_n14318_), .ZN(new_n14319_));
  OAI21_X1   g14225(.A1(new_n14310_), .A2(new_n14307_), .B(new_n14291_), .ZN(new_n14320_));
  OAI21_X1   g14226(.A1(new_n14311_), .A2(new_n14314_), .B(new_n14320_), .ZN(new_n14321_));
  NAND3_X1   g14227(.A1(new_n13664_), .A2(new_n13661_), .A3(new_n13578_), .ZN(new_n14322_));
  OAI21_X1   g14228(.A1(new_n13662_), .A2(new_n13660_), .B(new_n13032_), .ZN(new_n14323_));
  NAND2_X1   g14229(.A1(new_n14323_), .A2(new_n14322_), .ZN(new_n14324_));
  OAI21_X1   g14230(.A1(new_n14321_), .A2(new_n14318_), .B(new_n14324_), .ZN(new_n14325_));
  NAND3_X1   g14231(.A1(new_n14325_), .A2(new_n14288_), .A3(new_n14319_), .ZN(new_n14326_));
  INV_X1     g14232(.I(new_n13675_), .ZN(new_n14327_));
  NAND2_X1   g14233(.A1(new_n14326_), .A2(new_n14327_), .ZN(new_n14328_));
  AOI21_X1   g14234(.A1(new_n13681_), .A2(new_n13685_), .B(new_n13697_), .ZN(new_n14329_));
  AOI21_X1   g14235(.A1(new_n14328_), .A2(new_n13668_), .B(new_n14329_), .ZN(new_n14330_));
  OAI21_X1   g14236(.A1(new_n13706_), .A2(new_n13710_), .B(new_n13722_), .ZN(new_n14331_));
  OAI21_X1   g14237(.A1(new_n14330_), .A2(new_n13699_), .B(new_n14331_), .ZN(new_n14332_));
  NOR2_X1    g14238(.A1(new_n13732_), .A2(new_n13730_), .ZN(new_n14333_));
  AOI21_X1   g14239(.A1(new_n14332_), .A2(new_n13724_), .B(new_n14333_), .ZN(new_n14334_));
  NAND3_X1   g14240(.A1(new_n14332_), .A2(new_n13724_), .A3(new_n14333_), .ZN(new_n14335_));
  AOI21_X1   g14241(.A1(new_n14335_), .A2(new_n13739_), .B(new_n14334_), .ZN(new_n14336_));
  AND3_X2    g14242(.A1(new_n11268_), .A2(new_n451_), .A3(new_n13757_), .Z(new_n14337_));
  NOR2_X1    g14243(.A1(new_n14337_), .A2(new_n13758_), .ZN(new_n14338_));
  AOI21_X1   g14244(.A1(new_n14336_), .A2(new_n13752_), .B(new_n14338_), .ZN(new_n14339_));
  OAI21_X1   g14245(.A1(new_n14339_), .A2(new_n13753_), .B(new_n13768_), .ZN(new_n14340_));
  NOR3_X1    g14246(.A1(new_n14339_), .A2(new_n13753_), .A3(new_n13768_), .ZN(new_n14341_));
  OAI21_X1   g14247(.A1(new_n14341_), .A2(new_n13777_), .B(new_n14340_), .ZN(new_n14342_));
  OAI21_X1   g14248(.A1(new_n14342_), .A2(new_n13575_), .B(new_n13786_), .ZN(new_n14343_));
  AOI21_X1   g14249(.A1(new_n14343_), .A2(new_n13779_), .B(new_n13795_), .ZN(new_n14344_));
  NAND3_X1   g14250(.A1(new_n14343_), .A2(new_n13779_), .A3(new_n13795_), .ZN(new_n14345_));
  AOI21_X1   g14251(.A1(new_n14345_), .A2(new_n13804_), .B(new_n14344_), .ZN(new_n14346_));
  XOR2_X1    g14252(.A1(new_n13812_), .A2(new_n13811_), .Z(new_n14347_));
  AOI21_X1   g14253(.A1(new_n14346_), .A2(new_n13808_), .B(new_n14347_), .ZN(new_n14348_));
  OAI21_X1   g14254(.A1(new_n13188_), .A2(new_n13190_), .B(new_n13174_), .ZN(new_n14349_));
  OAI21_X1   g14255(.A1(new_n13174_), .A2(new_n13817_), .B(new_n14349_), .ZN(new_n14350_));
  OAI21_X1   g14256(.A1(new_n14348_), .A2(new_n13809_), .B(new_n14350_), .ZN(new_n14351_));
  NOR3_X1    g14257(.A1(new_n14348_), .A2(new_n13809_), .A3(new_n14350_), .ZN(new_n14352_));
  OAI21_X1   g14258(.A1(new_n14352_), .A2(new_n13827_), .B(new_n14351_), .ZN(new_n14353_));
  INV_X1     g14259(.I(new_n13847_), .ZN(new_n14354_));
  OAI21_X1   g14260(.A1(new_n14353_), .A2(new_n13837_), .B(new_n14354_), .ZN(new_n14355_));
  NOR3_X1    g14261(.A1(new_n13219_), .A2(new_n13842_), .A3(new_n13220_), .ZN(new_n14356_));
  NOR3_X1    g14262(.A1(new_n14356_), .A2(new_n13840_), .A3(new_n13843_), .ZN(new_n14357_));
  NOR2_X1    g14263(.A1(new_n14357_), .A2(new_n13853_), .ZN(new_n14358_));
  AOI21_X1   g14264(.A1(new_n14355_), .A2(new_n13838_), .B(new_n14358_), .ZN(new_n14359_));
  NAND3_X1   g14265(.A1(new_n14355_), .A2(new_n13838_), .A3(new_n14358_), .ZN(new_n14360_));
  AOI21_X1   g14266(.A1(new_n14360_), .A2(new_n13862_), .B(new_n14359_), .ZN(new_n14361_));
  AOI21_X1   g14267(.A1(new_n14361_), .A2(new_n13874_), .B(new_n13882_), .ZN(new_n14362_));
  INV_X1     g14268(.I(new_n13888_), .ZN(new_n14363_));
  NAND2_X1   g14269(.A1(new_n14363_), .A2(new_n13886_), .ZN(new_n14364_));
  INV_X1     g14270(.I(new_n13239_), .ZN(new_n14365_));
  NAND2_X1   g14271(.A1(new_n14365_), .A2(new_n13240_), .ZN(new_n14366_));
  MUX2_X1    g14272(.I0(new_n14364_), .I1(new_n14366_), .S(new_n13231_), .Z(new_n14367_));
  OAI21_X1   g14273(.A1(new_n14362_), .A2(new_n13875_), .B(new_n14367_), .ZN(new_n14368_));
  NOR3_X1    g14274(.A1(new_n14362_), .A2(new_n13875_), .A3(new_n14367_), .ZN(new_n14369_));
  OAI21_X1   g14275(.A1(new_n14369_), .A2(new_n13900_), .B(new_n14368_), .ZN(new_n14370_));
  INV_X1     g14276(.I(new_n13912_), .ZN(new_n14371_));
  OAI21_X1   g14277(.A1(new_n14370_), .A2(new_n13904_), .B(new_n14371_), .ZN(new_n14372_));
  INV_X1     g14278(.I(new_n13254_), .ZN(new_n14373_));
  OAI21_X1   g14279(.A1(new_n13241_), .A2(new_n13248_), .B(new_n14373_), .ZN(new_n14374_));
  AOI22_X1   g14280(.A1(new_n13915_), .A2(new_n13916_), .B1(new_n14374_), .B2(new_n13249_), .ZN(new_n14375_));
  AOI21_X1   g14281(.A1(new_n13914_), .A2(new_n13918_), .B(new_n14375_), .ZN(new_n14376_));
  AOI21_X1   g14282(.A1(new_n14372_), .A2(new_n13905_), .B(new_n14376_), .ZN(new_n14377_));
  NAND3_X1   g14283(.A1(new_n14372_), .A2(new_n14376_), .A3(new_n13905_), .ZN(new_n14378_));
  AOI21_X1   g14284(.A1(new_n14378_), .A2(new_n13924_), .B(new_n14377_), .ZN(new_n14379_));
  AOI21_X1   g14285(.A1(new_n14379_), .A2(new_n13929_), .B(new_n13938_), .ZN(new_n14380_));
  NAND2_X1   g14286(.A1(new_n13945_), .A2(new_n13943_), .ZN(new_n14381_));
  OAI21_X1   g14287(.A1(new_n14380_), .A2(new_n13930_), .B(new_n14381_), .ZN(new_n14382_));
  NOR3_X1    g14288(.A1(new_n14380_), .A2(new_n13930_), .A3(new_n14381_), .ZN(new_n14383_));
  OAI21_X1   g14289(.A1(new_n14383_), .A2(new_n13954_), .B(new_n14382_), .ZN(new_n14384_));
  INV_X1     g14290(.I(new_n13977_), .ZN(new_n14385_));
  OAI21_X1   g14291(.A1(new_n14384_), .A2(new_n13968_), .B(new_n14385_), .ZN(new_n14386_));
  AOI21_X1   g14292(.A1(new_n14386_), .A2(new_n13969_), .B(new_n13981_), .ZN(new_n14387_));
  NAND3_X1   g14293(.A1(new_n14386_), .A2(new_n13969_), .A3(new_n13981_), .ZN(new_n14388_));
  AOI21_X1   g14294(.A1(new_n14388_), .A2(new_n13988_), .B(new_n14387_), .ZN(new_n14389_));
  AOI21_X1   g14295(.A1(new_n14389_), .A2(new_n13992_), .B(new_n13997_), .ZN(new_n14390_));
  INV_X1     g14296(.I(new_n14002_), .ZN(new_n14391_));
  OAI21_X1   g14297(.A1(new_n14390_), .A2(new_n13993_), .B(new_n14391_), .ZN(new_n14392_));
  NOR3_X1    g14298(.A1(new_n14390_), .A2(new_n13993_), .A3(new_n14391_), .ZN(new_n14393_));
  OAI21_X1   g14299(.A1(new_n14393_), .A2(new_n14012_), .B(new_n14392_), .ZN(new_n14394_));
  INV_X1     g14300(.I(new_n14023_), .ZN(new_n14395_));
  OAI21_X1   g14301(.A1(new_n14394_), .A2(new_n14020_), .B(new_n14395_), .ZN(new_n14396_));
  AOI21_X1   g14302(.A1(new_n14396_), .A2(new_n14021_), .B(new_n14028_), .ZN(new_n14397_));
  NAND3_X1   g14303(.A1(new_n14396_), .A2(new_n14021_), .A3(new_n14028_), .ZN(new_n14398_));
  AOI21_X1   g14304(.A1(new_n14398_), .A2(new_n14036_), .B(new_n14397_), .ZN(new_n14399_));
  AOI21_X1   g14305(.A1(new_n14399_), .A2(new_n14041_), .B(new_n14046_), .ZN(new_n14400_));
  INV_X1     g14306(.I(new_n14057_), .ZN(new_n14401_));
  OAI21_X1   g14307(.A1(new_n14400_), .A2(new_n14042_), .B(new_n14401_), .ZN(new_n14402_));
  NOR3_X1    g14308(.A1(new_n14400_), .A2(new_n14042_), .A3(new_n14401_), .ZN(new_n14403_));
  OAI21_X1   g14309(.A1(new_n14403_), .A2(new_n14061_), .B(new_n14402_), .ZN(new_n14404_));
  INV_X1     g14310(.I(new_n14285_), .ZN(new_n14405_));
  NAND3_X1   g14311(.A1(new_n14404_), .A2(new_n14082_), .A3(new_n14405_), .ZN(new_n14406_));
  AOI21_X1   g14312(.A1(new_n14286_), .A2(new_n14406_), .B(new_n13567_), .ZN(new_n14407_));
  OAI21_X1   g14313(.A1(new_n14069_), .A2(new_n14070_), .B(new_n10980_), .ZN(new_n14408_));
  AOI21_X1   g14314(.A1(new_n14404_), .A2(new_n14082_), .B(new_n14405_), .ZN(new_n14409_));
  NOR2_X1    g14315(.A1(new_n14083_), .A2(new_n14285_), .ZN(new_n14410_));
  NOR3_X1    g14316(.A1(new_n14410_), .A2(new_n14409_), .A3(new_n14408_), .ZN(new_n14411_));
  NOR2_X1    g14317(.A1(new_n14411_), .A2(new_n14407_), .ZN(new_n14412_));
  NAND3_X1   g14318(.A1(new_n13566_), .A2(new_n13563_), .A3(new_n10981_), .ZN(new_n14413_));
  NAND2_X1   g14319(.A1(new_n14408_), .A2(new_n14413_), .ZN(new_n14414_));
  INV_X1     g14320(.I(new_n14068_), .ZN(new_n14415_));
  NOR2_X1    g14321(.A1(new_n14415_), .A2(new_n14080_), .ZN(new_n14416_));
  INV_X1     g14322(.I(new_n14416_), .ZN(new_n14417_));
  INV_X1     g14323(.I(new_n14080_), .ZN(new_n14418_));
  XOR2_X1    g14324(.A1(new_n14068_), .A2(new_n14418_), .Z(new_n14419_));
  AND3_X2    g14325(.A1(new_n14417_), .A2(new_n14414_), .A3(new_n14419_), .Z(new_n14420_));
  AOI21_X1   g14326(.A1(new_n14419_), .A2(new_n14414_), .B(new_n14417_), .ZN(new_n14421_));
  NOR2_X1    g14327(.A1(new_n14420_), .A2(new_n14421_), .ZN(new_n14422_));
  XNOR2_X1   g14328(.A1(new_n14404_), .A2(new_n14422_), .ZN(new_n14423_));
  XOR2_X1    g14329(.A1(new_n14412_), .A2(new_n14423_), .Z(\result[0] ));
  NOR2_X1    g14330(.A1(new_n14245_), .A2(new_n14408_), .ZN(new_n14425_));
  INV_X1     g14331(.I(new_n14425_), .ZN(new_n14426_));
  AOI21_X1   g14332(.A1(new_n14245_), .A2(new_n14408_), .B(new_n14284_), .ZN(new_n14427_));
  INV_X1     g14333(.I(new_n14427_), .ZN(new_n14428_));
  OAI21_X1   g14334(.A1(new_n14083_), .A2(new_n14428_), .B(new_n14426_), .ZN(new_n14429_));
  INV_X1     g14335(.I(new_n14240_), .ZN(new_n14430_));
  INV_X1     g14336(.I(new_n14092_), .ZN(new_n14431_));
  INV_X1     g14337(.I(new_n14231_), .ZN(new_n14432_));
  INV_X1     g14338(.I(new_n14199_), .ZN(new_n14433_));
  NOR2_X1    g14339(.A1(new_n14197_), .A2(new_n14198_), .ZN(new_n14434_));
  OAI22_X1   g14340(.A1(new_n14097_), .A2(new_n14093_), .B1(new_n14434_), .B2(new_n14195_), .ZN(new_n14435_));
  AOI21_X1   g14341(.A1(new_n14100_), .A2(new_n14098_), .B(new_n14160_), .ZN(new_n14436_));
  INV_X1     g14342(.I(new_n14154_), .ZN(new_n14437_));
  OAI21_X1   g14343(.A1(new_n14151_), .A2(new_n14153_), .B(new_n14437_), .ZN(new_n14438_));
  AOI22_X1   g14344(.A1(new_n11632_), .A2(new_n5783_), .B1(new_n10857_), .B2(new_n247_), .ZN(new_n14439_));
  OAI21_X1   g14345(.A1(new_n14439_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n14440_));
  XNOR2_X1   g14346(.A1(new_n11631_), .A2(new_n14440_), .ZN(new_n14441_));
  INV_X1     g14347(.I(new_n14441_), .ZN(new_n14442_));
  INV_X1     g14348(.I(new_n14111_), .ZN(new_n14443_));
  NOR2_X1    g14349(.A1(new_n14113_), .A2(new_n14128_), .ZN(new_n14444_));
  NOR2_X1    g14350(.A1(new_n14444_), .A2(new_n14129_), .ZN(new_n14445_));
  NOR2_X1    g14351(.A1(new_n14118_), .A2(new_n14122_), .ZN(new_n14446_));
  NAND2_X1   g14352(.A1(new_n10794_), .A2(new_n87_), .ZN(new_n14447_));
  AOI22_X1   g14353(.A1(new_n10691_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n10809_), .ZN(new_n14448_));
  AOI21_X1   g14354(.A1(new_n14448_), .A2(new_n14447_), .B(new_n82_), .ZN(new_n14449_));
  NAND2_X1   g14355(.A1(new_n11333_), .A2(new_n14449_), .ZN(new_n14450_));
  XNOR2_X1   g14356(.A1(new_n14450_), .A2(new_n14446_), .ZN(new_n14451_));
  AOI22_X1   g14357(.A1(new_n10805_), .A2(new_n4526_), .B1(new_n4570_), .B2(new_n10817_), .ZN(new_n14452_));
  NOR2_X1    g14358(.A1(new_n11214_), .A2(new_n79_), .ZN(new_n14453_));
  OAI21_X1   g14359(.A1(new_n14453_), .A2(new_n14452_), .B(new_n72_), .ZN(new_n14454_));
  NAND2_X1   g14360(.A1(new_n14454_), .A2(new_n101_), .ZN(new_n14455_));
  XOR2_X1    g14361(.A1(new_n11224_), .A2(new_n14455_), .Z(new_n14456_));
  XNOR2_X1   g14362(.A1(new_n14456_), .A2(new_n14451_), .ZN(new_n14457_));
  NOR2_X1    g14363(.A1(new_n14456_), .A2(new_n14451_), .ZN(new_n14458_));
  INV_X1     g14364(.I(new_n14458_), .ZN(new_n14459_));
  NAND2_X1   g14365(.A1(new_n14456_), .A2(new_n14451_), .ZN(new_n14460_));
  NAND2_X1   g14366(.A1(new_n14459_), .A2(new_n14460_), .ZN(new_n14461_));
  NAND2_X1   g14367(.A1(new_n14445_), .A2(new_n14461_), .ZN(new_n14462_));
  OAI21_X1   g14368(.A1(new_n14445_), .A2(new_n14457_), .B(new_n14462_), .ZN(new_n14463_));
  OAI22_X1   g14369(.A1(new_n11264_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10646_), .ZN(new_n14464_));
  OAI21_X1   g14370(.A1(new_n1128_), .A2(new_n10633_), .B(new_n14464_), .ZN(new_n14465_));
  AOI21_X1   g14371(.A1(new_n14465_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n14466_));
  XOR2_X1    g14372(.A1(new_n11385_), .A2(new_n14466_), .Z(new_n14467_));
  NOR2_X1    g14373(.A1(new_n14467_), .A2(new_n14463_), .ZN(new_n14468_));
  NAND2_X1   g14374(.A1(new_n14467_), .A2(new_n14463_), .ZN(new_n14469_));
  INV_X1     g14375(.I(new_n14469_), .ZN(new_n14470_));
  NOR2_X1    g14376(.A1(new_n14470_), .A2(new_n14468_), .ZN(new_n14471_));
  NOR3_X1    g14377(.A1(new_n14471_), .A2(new_n14137_), .A3(new_n14143_), .ZN(new_n14472_));
  NOR2_X1    g14378(.A1(new_n14132_), .A2(new_n14136_), .ZN(new_n14473_));
  OAI21_X1   g14379(.A1(new_n14472_), .A2(new_n14473_), .B(new_n14443_), .ZN(new_n14474_));
  INV_X1     g14380(.I(new_n14474_), .ZN(new_n14475_));
  NOR3_X1    g14381(.A1(new_n14472_), .A2(new_n14443_), .A3(new_n14473_), .ZN(new_n14476_));
  NOR3_X1    g14382(.A1(new_n14475_), .A2(new_n14442_), .A3(new_n14476_), .ZN(new_n14477_));
  INV_X1     g14383(.I(new_n14476_), .ZN(new_n14478_));
  AOI21_X1   g14384(.A1(new_n14478_), .A2(new_n14474_), .B(new_n14441_), .ZN(new_n14479_));
  NOR2_X1    g14385(.A1(new_n14477_), .A2(new_n14479_), .ZN(new_n14480_));
  NOR2_X1    g14386(.A1(new_n14438_), .A2(new_n14480_), .ZN(new_n14481_));
  AOI21_X1   g14387(.A1(new_n14103_), .A2(new_n14152_), .B(new_n14154_), .ZN(new_n14482_));
  INV_X1     g14388(.I(new_n14480_), .ZN(new_n14483_));
  NOR2_X1    g14389(.A1(new_n14483_), .A2(new_n14482_), .ZN(new_n14484_));
  OAI22_X1   g14390(.A1(new_n11803_), .A2(new_n5336_), .B1(new_n5398_), .B2(new_n10881_), .ZN(new_n14485_));
  AOI21_X1   g14391(.A1(new_n14485_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n14486_));
  XOR2_X1    g14392(.A1(new_n11802_), .A2(new_n14486_), .Z(new_n14487_));
  INV_X1     g14393(.I(new_n14487_), .ZN(new_n14488_));
  NOR3_X1    g14394(.A1(new_n14484_), .A2(new_n14481_), .A3(new_n14488_), .ZN(new_n14489_));
  NAND2_X1   g14395(.A1(new_n14483_), .A2(new_n14482_), .ZN(new_n14490_));
  NAND2_X1   g14396(.A1(new_n14438_), .A2(new_n14480_), .ZN(new_n14491_));
  AOI21_X1   g14397(.A1(new_n14490_), .A2(new_n14491_), .B(new_n14487_), .ZN(new_n14492_));
  NOR4_X1    g14398(.A1(new_n14436_), .A2(new_n14162_), .A3(new_n14489_), .A4(new_n14492_), .ZN(new_n14493_));
  NOR2_X1    g14399(.A1(new_n14436_), .A2(new_n14162_), .ZN(new_n14494_));
  NOR2_X1    g14400(.A1(new_n14489_), .A2(new_n14492_), .ZN(new_n14495_));
  NOR2_X1    g14401(.A1(new_n14494_), .A2(new_n14495_), .ZN(new_n14496_));
  AOI22_X1   g14402(.A1(new_n10986_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n10897_), .ZN(new_n14497_));
  OAI21_X1   g14403(.A1(new_n14497_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n14498_));
  XOR2_X1    g14404(.A1(new_n10984_), .A2(new_n14498_), .Z(new_n14499_));
  INV_X1     g14405(.I(new_n14499_), .ZN(new_n14500_));
  NOR3_X1    g14406(.A1(new_n14496_), .A2(new_n14500_), .A3(new_n14493_), .ZN(new_n14501_));
  OAI21_X1   g14407(.A1(new_n14496_), .A2(new_n14493_), .B(new_n14500_), .ZN(new_n14502_));
  INV_X1     g14408(.I(new_n14502_), .ZN(new_n14503_));
  NOR3_X1    g14409(.A1(new_n14503_), .A2(new_n14501_), .A3(new_n14172_), .ZN(new_n14504_));
  NOR3_X1    g14410(.A1(new_n14504_), .A2(new_n14186_), .A3(new_n14183_), .ZN(new_n14505_));
  NOR2_X1    g14411(.A1(new_n14496_), .A2(new_n14493_), .ZN(new_n14506_));
  NAND2_X1   g14412(.A1(new_n14506_), .A2(new_n14499_), .ZN(new_n14507_));
  NAND3_X1   g14413(.A1(new_n14507_), .A2(new_n14502_), .A3(new_n14181_), .ZN(new_n14508_));
  AOI21_X1   g14414(.A1(new_n14508_), .A2(new_n14179_), .B(new_n14175_), .ZN(new_n14509_));
  OAI22_X1   g14415(.A1(new_n12601_), .A2(new_n5967_), .B1(new_n643_), .B2(new_n10595_), .ZN(new_n14510_));
  AOI21_X1   g14416(.A1(new_n14510_), .A2(new_n279_), .B(new_n643_), .ZN(new_n14511_));
  INV_X1     g14417(.I(new_n14511_), .ZN(new_n14512_));
  NOR2_X1    g14418(.A1(new_n13949_), .A2(new_n14512_), .ZN(new_n14513_));
  NOR2_X1    g14419(.A1(new_n12600_), .A2(new_n14511_), .ZN(new_n14514_));
  NOR2_X1    g14420(.A1(new_n14514_), .A2(new_n14513_), .ZN(new_n14515_));
  NOR3_X1    g14421(.A1(new_n14505_), .A2(new_n14509_), .A3(new_n14515_), .ZN(new_n14516_));
  NAND3_X1   g14422(.A1(new_n14508_), .A2(new_n14175_), .A3(new_n14179_), .ZN(new_n14517_));
  OAI21_X1   g14423(.A1(new_n14504_), .A2(new_n14186_), .B(new_n14183_), .ZN(new_n14518_));
  INV_X1     g14424(.I(new_n14515_), .ZN(new_n14519_));
  AOI21_X1   g14425(.A1(new_n14518_), .A2(new_n14517_), .B(new_n14519_), .ZN(new_n14520_));
  NOR2_X1    g14426(.A1(new_n14516_), .A2(new_n14520_), .ZN(new_n14521_));
  NAND3_X1   g14427(.A1(new_n14435_), .A2(new_n14521_), .A3(new_n14433_), .ZN(new_n14522_));
  INV_X1     g14428(.I(new_n14093_), .ZN(new_n14523_));
  INV_X1     g14429(.I(new_n13500_), .ZN(new_n14524_));
  NAND3_X1   g14430(.A1(new_n13494_), .A2(new_n13497_), .A3(new_n12865_), .ZN(new_n14525_));
  NAND4_X1   g14431(.A1(new_n12868_), .A2(new_n14525_), .A3(new_n12871_), .A4(new_n14524_), .ZN(new_n14526_));
  AOI21_X1   g14432(.A1(new_n14526_), .A2(new_n14523_), .B(new_n14196_), .ZN(new_n14527_));
  OAI22_X1   g14433(.A1(new_n14527_), .A2(new_n14199_), .B1(new_n14516_), .B2(new_n14520_), .ZN(new_n14528_));
  NAND2_X1   g14434(.A1(new_n10916_), .A2(new_n12886_), .ZN(new_n14529_));
  INV_X1     g14435(.I(new_n12888_), .ZN(new_n14530_));
  NAND2_X1   g14436(.A1(new_n14530_), .A2(new_n14529_), .ZN(new_n14531_));
  AOI22_X1   g14437(.A1(new_n12891_), .A2(new_n6758_), .B1(new_n10924_), .B2(new_n805_), .ZN(new_n14532_));
  OAI21_X1   g14438(.A1(new_n14532_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n14533_));
  NOR2_X1    g14439(.A1(new_n14531_), .A2(new_n14533_), .ZN(new_n14534_));
  INV_X1     g14440(.I(new_n14533_), .ZN(new_n14535_));
  NOR2_X1    g14441(.A1(new_n12889_), .A2(new_n14535_), .ZN(new_n14536_));
  NOR2_X1    g14442(.A1(new_n14534_), .A2(new_n14536_), .ZN(new_n14537_));
  NAND3_X1   g14443(.A1(new_n14522_), .A2(new_n14528_), .A3(new_n14537_), .ZN(new_n14538_));
  NOR4_X1    g14444(.A1(new_n14527_), .A2(new_n14199_), .A3(new_n14516_), .A4(new_n14520_), .ZN(new_n14539_));
  AOI21_X1   g14445(.A1(new_n14433_), .A2(new_n14435_), .B(new_n14521_), .ZN(new_n14540_));
  INV_X1     g14446(.I(new_n14537_), .ZN(new_n14541_));
  OAI21_X1   g14447(.A1(new_n14540_), .A2(new_n14539_), .B(new_n14541_), .ZN(new_n14542_));
  NAND3_X1   g14448(.A1(new_n14542_), .A2(new_n14538_), .A3(new_n14209_), .ZN(new_n14543_));
  NAND3_X1   g14449(.A1(new_n14543_), .A2(new_n14224_), .A3(new_n14221_), .ZN(new_n14544_));
  INV_X1     g14450(.I(new_n14544_), .ZN(new_n14545_));
  AOI21_X1   g14451(.A1(new_n14543_), .A2(new_n14224_), .B(new_n14221_), .ZN(new_n14546_));
  AOI22_X1   g14452(.A1(new_n12909_), .A2(new_n7838_), .B1(new_n10949_), .B2(new_n2469_), .ZN(new_n14547_));
  OAI21_X1   g14453(.A1(new_n14547_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n14548_));
  XOR2_X1    g14454(.A1(new_n12907_), .A2(new_n14548_), .Z(new_n14549_));
  NOR3_X1    g14455(.A1(new_n14545_), .A2(new_n14546_), .A3(new_n14549_), .ZN(new_n14550_));
  INV_X1     g14456(.I(new_n14546_), .ZN(new_n14551_));
  INV_X1     g14457(.I(new_n14549_), .ZN(new_n14552_));
  AOI21_X1   g14458(.A1(new_n14551_), .A2(new_n14544_), .B(new_n14552_), .ZN(new_n14553_));
  NOR3_X1    g14459(.A1(new_n14553_), .A2(new_n14550_), .A3(new_n14432_), .ZN(new_n14554_));
  INV_X1     g14460(.I(new_n14554_), .ZN(new_n14555_));
  NAND3_X1   g14461(.A1(new_n14555_), .A2(new_n14232_), .A3(new_n14431_), .ZN(new_n14556_));
  INV_X1     g14462(.I(new_n14232_), .ZN(new_n14557_));
  OAI21_X1   g14463(.A1(new_n14557_), .A2(new_n14554_), .B(new_n14092_), .ZN(new_n14558_));
  OAI22_X1   g14464(.A1(new_n10965_), .A2(new_n8831_), .B1(new_n3040_), .B2(new_n10570_), .ZN(new_n14559_));
  AOI21_X1   g14465(.A1(new_n14559_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n14560_));
  XNOR2_X1   g14466(.A1(new_n14077_), .A2(new_n14560_), .ZN(new_n14561_));
  NAND3_X1   g14467(.A1(new_n14556_), .A2(new_n14558_), .A3(new_n14561_), .ZN(new_n14562_));
  NOR3_X1    g14468(.A1(new_n14557_), .A2(new_n14554_), .A3(new_n14092_), .ZN(new_n14563_));
  AOI21_X1   g14469(.A1(new_n14555_), .A2(new_n14232_), .B(new_n14431_), .ZN(new_n14564_));
  INV_X1     g14470(.I(new_n14561_), .ZN(new_n14565_));
  OAI21_X1   g14471(.A1(new_n14564_), .A2(new_n14563_), .B(new_n14565_), .ZN(new_n14566_));
  AND2_X2    g14472(.A1(new_n14566_), .A2(new_n14562_), .Z(new_n14567_));
  NAND2_X1   g14473(.A1(new_n14567_), .A2(new_n14430_), .ZN(new_n14568_));
  NAND3_X1   g14474(.A1(new_n14568_), .A2(new_n14088_), .A3(new_n14244_), .ZN(new_n14569_));
  AND3_X2    g14475(.A1(new_n14430_), .A2(new_n14562_), .A3(new_n14566_), .Z(new_n14570_));
  OAI22_X1   g14476(.A1(new_n14570_), .A2(new_n14243_), .B1(new_n14084_), .B2(new_n14087_), .ZN(new_n14571_));
  NAND2_X1   g14477(.A1(new_n14569_), .A2(new_n14571_), .ZN(new_n14572_));
  INV_X1     g14478(.I(new_n14572_), .ZN(new_n14573_));
  INV_X1     g14479(.I(new_n14275_), .ZN(new_n14574_));
  OAI21_X1   g14480(.A1(new_n14246_), .A2(new_n14277_), .B(new_n14574_), .ZN(new_n14575_));
  INV_X1     g14481(.I(new_n14252_), .ZN(new_n14576_));
  NAND2_X1   g14482(.A1(new_n14576_), .A2(new_n14270_), .ZN(new_n14577_));
  INV_X1     g14483(.I(new_n14273_), .ZN(new_n14578_));
  OAI21_X1   g14484(.A1(new_n14255_), .A2(new_n14266_), .B(new_n14267_), .ZN(new_n14579_));
  INV_X1     g14485(.I(new_n4545_), .ZN(new_n14580_));
  NOR3_X1    g14486(.A1(new_n14580_), .A2(new_n83_), .A3(new_n960_), .ZN(new_n14581_));
  AOI21_X1   g14487(.A1(new_n4609_), .A2(new_n14581_), .B(new_n80_), .ZN(new_n14582_));
  NAND2_X1   g14488(.A1(new_n4609_), .A2(new_n14581_), .ZN(new_n14583_));
  NOR2_X1    g14489(.A1(new_n14583_), .A2(new_n102_), .ZN(new_n14584_));
  OAI21_X1   g14490(.A1(new_n14584_), .A2(new_n14582_), .B(new_n14261_), .ZN(new_n14585_));
  XOR2_X1    g14491(.A1(new_n14583_), .A2(new_n80_), .Z(new_n14586_));
  OAI21_X1   g14492(.A1(new_n14261_), .A2(new_n14586_), .B(new_n14585_), .ZN(new_n14587_));
  XOR2_X1    g14493(.A1(new_n14579_), .A2(new_n14587_), .Z(new_n14588_));
  NAND2_X1   g14494(.A1(new_n14578_), .A2(new_n14588_), .ZN(new_n14589_));
  XNOR2_X1   g14495(.A1(new_n14589_), .A2(new_n14577_), .ZN(new_n14590_));
  NOR2_X1    g14496(.A1(new_n14250_), .A2(new_n14590_), .ZN(new_n14591_));
  NAND2_X1   g14497(.A1(new_n14250_), .A2(new_n14590_), .ZN(new_n14592_));
  INV_X1     g14498(.I(new_n14592_), .ZN(new_n14593_));
  NOR2_X1    g14499(.A1(new_n14593_), .A2(new_n14591_), .ZN(new_n14594_));
  XOR2_X1    g14500(.A1(new_n14594_), .A2(new_n14274_), .Z(new_n14595_));
  INV_X1     g14501(.I(new_n14595_), .ZN(new_n14596_));
  NAND2_X1   g14502(.A1(new_n14276_), .A2(new_n14594_), .ZN(new_n14597_));
  NOR2_X1    g14503(.A1(new_n14276_), .A2(new_n14594_), .ZN(new_n14598_));
  INV_X1     g14504(.I(new_n14598_), .ZN(new_n14599_));
  AOI21_X1   g14505(.A1(new_n14597_), .A2(new_n14599_), .B(new_n14575_), .ZN(new_n14600_));
  AOI21_X1   g14506(.A1(new_n14575_), .A2(new_n14596_), .B(new_n14600_), .ZN(new_n14601_));
  INV_X1     g14507(.I(new_n14277_), .ZN(new_n14602_));
  INV_X1     g14508(.I(new_n14594_), .ZN(new_n14603_));
  AOI22_X1   g14509(.A1(new_n14602_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n14603_), .ZN(new_n14604_));
  OAI21_X1   g14510(.A1(new_n14604_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n14605_));
  XNOR2_X1   g14511(.A1(new_n14601_), .A2(new_n14605_), .ZN(new_n14606_));
  NAND2_X1   g14512(.A1(new_n14573_), .A2(new_n14606_), .ZN(new_n14607_));
  INV_X1     g14513(.I(new_n14606_), .ZN(new_n14608_));
  NAND2_X1   g14514(.A1(new_n14572_), .A2(new_n14608_), .ZN(new_n14609_));
  NAND2_X1   g14515(.A1(new_n14607_), .A2(new_n14609_), .ZN(new_n14610_));
  NAND2_X1   g14516(.A1(new_n14429_), .A2(new_n14610_), .ZN(new_n14611_));
  XOR2_X1    g14517(.A1(new_n14423_), .A2(new_n14611_), .Z(new_n14612_));
  XOR2_X1    g14518(.A1(new_n14612_), .A2(new_n14412_), .Z(\result[1] ));
  INV_X1     g14519(.I(new_n14610_), .ZN(new_n14614_));
  OAI21_X1   g14520(.A1(new_n14411_), .A2(new_n14407_), .B(new_n14614_), .ZN(new_n14615_));
  OAI21_X1   g14521(.A1(new_n14410_), .A2(new_n14409_), .B(new_n14408_), .ZN(new_n14616_));
  NAND3_X1   g14522(.A1(new_n14286_), .A2(new_n14406_), .A3(new_n13567_), .ZN(new_n14617_));
  NAND3_X1   g14523(.A1(new_n14616_), .A2(new_n14617_), .A3(new_n14610_), .ZN(new_n14618_));
  NAND2_X1   g14524(.A1(new_n14423_), .A2(new_n14429_), .ZN(new_n14619_));
  AOI21_X1   g14525(.A1(new_n14615_), .A2(new_n14618_), .B(new_n14619_), .ZN(new_n14620_));
  AOI21_X1   g14526(.A1(new_n13139_), .A2(new_n13142_), .B(new_n13121_), .ZN(new_n14621_));
  AOI21_X1   g14527(.A1(new_n13121_), .A2(new_n13570_), .B(new_n14621_), .ZN(new_n14622_));
  AOI21_X1   g14528(.A1(new_n14325_), .A2(new_n14319_), .B(new_n14288_), .ZN(new_n14623_));
  AOI21_X1   g14529(.A1(new_n14326_), .A2(new_n14327_), .B(new_n14623_), .ZN(new_n14624_));
  OAI21_X1   g14530(.A1(new_n14624_), .A2(new_n14329_), .B(new_n13698_), .ZN(new_n14625_));
  AOI21_X1   g14531(.A1(new_n14625_), .A2(new_n14331_), .B(new_n13723_), .ZN(new_n14626_));
  XNOR2_X1   g14532(.A1(new_n13738_), .A2(new_n13736_), .ZN(new_n14627_));
  AOI21_X1   g14533(.A1(new_n14626_), .A2(new_n14333_), .B(new_n14627_), .ZN(new_n14628_));
  OAI21_X1   g14534(.A1(new_n13749_), .A2(new_n13750_), .B(new_n13093_), .ZN(new_n14629_));
  NAND3_X1   g14535(.A1(new_n13747_), .A2(new_n13743_), .A3(new_n13024_), .ZN(new_n14630_));
  NAND2_X1   g14536(.A1(new_n14629_), .A2(new_n14630_), .ZN(new_n14631_));
  OAI21_X1   g14537(.A1(new_n14628_), .A2(new_n14334_), .B(new_n14631_), .ZN(new_n14632_));
  NOR3_X1    g14538(.A1(new_n14628_), .A2(new_n14334_), .A3(new_n14631_), .ZN(new_n14633_));
  OAI21_X1   g14539(.A1(new_n14633_), .A2(new_n14338_), .B(new_n14632_), .ZN(new_n14634_));
  OAI21_X1   g14540(.A1(new_n11385_), .A2(new_n13773_), .B(\a[2] ), .ZN(new_n14635_));
  NAND3_X1   g14541(.A1(new_n11987_), .A2(new_n451_), .A3(new_n13774_), .ZN(new_n14636_));
  NAND2_X1   g14542(.A1(new_n14635_), .A2(new_n14636_), .ZN(new_n14637_));
  OAI21_X1   g14543(.A1(new_n14634_), .A2(new_n13768_), .B(new_n14637_), .ZN(new_n14638_));
  AOI21_X1   g14544(.A1(new_n14638_), .A2(new_n14340_), .B(new_n14622_), .ZN(new_n14639_));
  NAND3_X1   g14545(.A1(new_n14638_), .A2(new_n14622_), .A3(new_n14340_), .ZN(new_n14640_));
  AOI21_X1   g14546(.A1(new_n14640_), .A2(new_n13786_), .B(new_n14639_), .ZN(new_n14641_));
  AOI21_X1   g14547(.A1(new_n14641_), .A2(new_n13795_), .B(new_n13803_), .ZN(new_n14642_));
  XOR2_X1    g14548(.A1(new_n11631_), .A2(new_n13807_), .Z(new_n14643_));
  OAI21_X1   g14549(.A1(new_n14642_), .A2(new_n14344_), .B(new_n14643_), .ZN(new_n14644_));
  NOR3_X1    g14550(.A1(new_n14642_), .A2(new_n14344_), .A3(new_n14643_), .ZN(new_n14645_));
  OAI21_X1   g14551(.A1(new_n14645_), .A2(new_n14347_), .B(new_n14644_), .ZN(new_n14646_));
  NAND3_X1   g14552(.A1(new_n13825_), .A2(\a[2] ), .A3(new_n13822_), .ZN(new_n14647_));
  OAI21_X1   g14553(.A1(new_n13821_), .A2(new_n13823_), .B(new_n451_), .ZN(new_n14648_));
  NAND2_X1   g14554(.A1(new_n14648_), .A2(new_n14647_), .ZN(new_n14649_));
  OAI21_X1   g14555(.A1(new_n14646_), .A2(new_n14350_), .B(new_n14649_), .ZN(new_n14650_));
  AOI21_X1   g14556(.A1(new_n14650_), .A2(new_n14351_), .B(new_n13836_), .ZN(new_n14651_));
  NAND3_X1   g14557(.A1(new_n14650_), .A2(new_n14351_), .A3(new_n13836_), .ZN(new_n14652_));
  AOI21_X1   g14558(.A1(new_n14652_), .A2(new_n14354_), .B(new_n14651_), .ZN(new_n14653_));
  AOI21_X1   g14559(.A1(new_n14653_), .A2(new_n14358_), .B(new_n13861_), .ZN(new_n14654_));
  OAI21_X1   g14560(.A1(new_n13871_), .A2(new_n13872_), .B(new_n13850_), .ZN(new_n14655_));
  NAND3_X1   g14561(.A1(new_n13869_), .A2(new_n13865_), .A3(new_n13220_), .ZN(new_n14656_));
  NAND2_X1   g14562(.A1(new_n14655_), .A2(new_n14656_), .ZN(new_n14657_));
  OAI21_X1   g14563(.A1(new_n14654_), .A2(new_n14359_), .B(new_n14657_), .ZN(new_n14658_));
  NOR3_X1    g14564(.A1(new_n14654_), .A2(new_n14359_), .A3(new_n14657_), .ZN(new_n14659_));
  OAI21_X1   g14565(.A1(new_n14659_), .A2(new_n13882_), .B(new_n14658_), .ZN(new_n14660_));
  INV_X1     g14566(.I(new_n13900_), .ZN(new_n14661_));
  OAI21_X1   g14567(.A1(new_n14660_), .A2(new_n14367_), .B(new_n14661_), .ZN(new_n14662_));
  INV_X1     g14568(.I(new_n13904_), .ZN(new_n14663_));
  AOI21_X1   g14569(.A1(new_n14662_), .A2(new_n14368_), .B(new_n14663_), .ZN(new_n14664_));
  NAND3_X1   g14570(.A1(new_n14662_), .A2(new_n14368_), .A3(new_n14663_), .ZN(new_n14665_));
  AOI21_X1   g14571(.A1(new_n14665_), .A2(new_n14371_), .B(new_n14664_), .ZN(new_n14666_));
  AOI21_X1   g14572(.A1(new_n14666_), .A2(new_n14376_), .B(new_n13923_), .ZN(new_n14667_));
  INV_X1     g14573(.I(new_n13929_), .ZN(new_n14668_));
  OAI21_X1   g14574(.A1(new_n14667_), .A2(new_n14377_), .B(new_n14668_), .ZN(new_n14669_));
  NOR3_X1    g14575(.A1(new_n14667_), .A2(new_n14377_), .A3(new_n14668_), .ZN(new_n14670_));
  OAI21_X1   g14576(.A1(new_n14670_), .A2(new_n13938_), .B(new_n14669_), .ZN(new_n14671_));
  INV_X1     g14577(.I(new_n13954_), .ZN(new_n14672_));
  OAI21_X1   g14578(.A1(new_n14671_), .A2(new_n14381_), .B(new_n14672_), .ZN(new_n14673_));
  AOI21_X1   g14579(.A1(new_n13966_), .A2(new_n13965_), .B(new_n13964_), .ZN(new_n14674_));
  NOR3_X1    g14580(.A1(new_n13958_), .A2(new_n13962_), .A3(new_n13956_), .ZN(new_n14675_));
  NOR2_X1    g14581(.A1(new_n14675_), .A2(new_n14674_), .ZN(new_n14676_));
  AOI21_X1   g14582(.A1(new_n14673_), .A2(new_n14382_), .B(new_n14676_), .ZN(new_n14677_));
  NAND3_X1   g14583(.A1(new_n14673_), .A2(new_n14382_), .A3(new_n14676_), .ZN(new_n14678_));
  AOI21_X1   g14584(.A1(new_n14678_), .A2(new_n14385_), .B(new_n14677_), .ZN(new_n14679_));
  XNOR2_X1   g14585(.A1(new_n13987_), .A2(new_n13984_), .ZN(new_n14680_));
  AOI21_X1   g14586(.A1(new_n14679_), .A2(new_n13981_), .B(new_n14680_), .ZN(new_n14681_));
  INV_X1     g14587(.I(new_n13992_), .ZN(new_n14682_));
  OAI21_X1   g14588(.A1(new_n14681_), .A2(new_n14387_), .B(new_n14682_), .ZN(new_n14683_));
  NOR3_X1    g14589(.A1(new_n14681_), .A2(new_n14387_), .A3(new_n14682_), .ZN(new_n14684_));
  OAI21_X1   g14590(.A1(new_n14684_), .A2(new_n13997_), .B(new_n14683_), .ZN(new_n14685_));
  XNOR2_X1   g14591(.A1(new_n14011_), .A2(new_n14006_), .ZN(new_n14686_));
  OAI21_X1   g14592(.A1(new_n14685_), .A2(new_n14391_), .B(new_n14686_), .ZN(new_n14687_));
  AOI21_X1   g14593(.A1(new_n14687_), .A2(new_n14392_), .B(new_n14019_), .ZN(new_n14688_));
  NAND3_X1   g14594(.A1(new_n14687_), .A2(new_n14392_), .A3(new_n14019_), .ZN(new_n14689_));
  AOI21_X1   g14595(.A1(new_n14689_), .A2(new_n14395_), .B(new_n14688_), .ZN(new_n14690_));
  AOI21_X1   g14596(.A1(new_n14690_), .A2(new_n14028_), .B(new_n14035_), .ZN(new_n14691_));
  INV_X1     g14597(.I(new_n14041_), .ZN(new_n14692_));
  OAI21_X1   g14598(.A1(new_n14691_), .A2(new_n14397_), .B(new_n14692_), .ZN(new_n14693_));
  NOR3_X1    g14599(.A1(new_n14691_), .A2(new_n14397_), .A3(new_n14692_), .ZN(new_n14694_));
  OAI21_X1   g14600(.A1(new_n14694_), .A2(new_n14046_), .B(new_n14693_), .ZN(new_n14695_));
  INV_X1     g14601(.I(new_n14061_), .ZN(new_n14696_));
  OAI21_X1   g14602(.A1(new_n14695_), .A2(new_n14401_), .B(new_n14696_), .ZN(new_n14697_));
  NAND3_X1   g14603(.A1(new_n14408_), .A2(new_n14413_), .A3(new_n14415_), .ZN(new_n14698_));
  AOI21_X1   g14604(.A1(new_n14408_), .A2(new_n14413_), .B(new_n14415_), .ZN(new_n14699_));
  OAI21_X1   g14605(.A1(new_n14418_), .A2(new_n14699_), .B(new_n14698_), .ZN(new_n14700_));
  AOI21_X1   g14606(.A1(new_n14697_), .A2(new_n14402_), .B(new_n14700_), .ZN(new_n14701_));
  AOI21_X1   g14607(.A1(new_n14701_), .A2(new_n14427_), .B(new_n14425_), .ZN(new_n14702_));
  INV_X1     g14608(.I(new_n13535_), .ZN(new_n14703_));
  NAND2_X1   g14609(.A1(new_n13405_), .A2(new_n14703_), .ZN(new_n14704_));
  INV_X1     g14610(.I(new_n14086_), .ZN(new_n14705_));
  OAI21_X1   g14611(.A1(new_n13405_), .A2(new_n14703_), .B(new_n14705_), .ZN(new_n14706_));
  NOR2_X1    g14612(.A1(new_n14242_), .A2(new_n14240_), .ZN(new_n14707_));
  AOI21_X1   g14613(.A1(new_n14706_), .A2(new_n14704_), .B(new_n14707_), .ZN(new_n14708_));
  AOI22_X1   g14614(.A1(new_n14091_), .A2(new_n14089_), .B1(new_n14230_), .B2(new_n14231_), .ZN(new_n14710_));
  INV_X1     g14615(.I(new_n14710_), .ZN(new_n14711_));
  NOR3_X1    g14616(.A1(new_n14540_), .A2(new_n14539_), .A3(new_n14541_), .ZN(new_n14712_));
  AOI21_X1   g14617(.A1(new_n14522_), .A2(new_n14528_), .B(new_n14537_), .ZN(new_n14713_));
  OAI21_X1   g14618(.A1(new_n14712_), .A2(new_n14713_), .B(new_n14220_), .ZN(new_n14714_));
  AOI21_X1   g14619(.A1(new_n14714_), .A2(new_n14218_), .B(new_n14221_), .ZN(new_n14715_));
  OAI21_X1   g14620(.A1(new_n14503_), .A2(new_n14501_), .B(new_n14172_), .ZN(new_n14716_));
  AOI21_X1   g14621(.A1(new_n14716_), .A2(new_n14186_), .B(new_n14175_), .ZN(new_n14717_));
  NAND2_X1   g14622(.A1(new_n14494_), .A2(new_n14495_), .ZN(new_n14718_));
  INV_X1     g14623(.I(new_n14468_), .ZN(new_n14719_));
  NAND2_X1   g14624(.A1(new_n14719_), .A2(new_n14469_), .ZN(new_n14720_));
  AOI21_X1   g14625(.A1(new_n14720_), .A2(new_n14140_), .B(new_n14141_), .ZN(new_n14721_));
  OAI21_X1   g14626(.A1(new_n14720_), .A2(new_n14140_), .B(new_n14111_), .ZN(new_n14722_));
  NOR2_X1    g14627(.A1(new_n14722_), .A2(new_n14721_), .ZN(new_n14723_));
  OAI21_X1   g14628(.A1(new_n14445_), .A2(new_n14458_), .B(new_n14460_), .ZN(new_n14724_));
  NOR3_X1    g14629(.A1(new_n14450_), .A2(new_n14118_), .A3(new_n14122_), .ZN(new_n14725_));
  AOI22_X1   g14630(.A1(new_n10691_), .A2(new_n87_), .B1(new_n10794_), .B2(new_n4406_), .ZN(new_n14726_));
  OAI21_X1   g14631(.A1(new_n10672_), .A2(new_n511_), .B(new_n14726_), .ZN(new_n14727_));
  AND3_X2    g14632(.A1(new_n11158_), .A2(new_n961_), .A3(new_n14727_), .Z(new_n14728_));
  XNOR2_X1   g14633(.A1(new_n14725_), .A2(new_n14728_), .ZN(new_n14729_));
  INV_X1     g14634(.I(new_n14729_), .ZN(new_n14730_));
  AOI22_X1   g14635(.A1(new_n10652_), .A2(new_n4526_), .B1(new_n4570_), .B2(new_n10805_), .ZN(new_n14731_));
  NOR2_X1    g14636(.A1(new_n10646_), .A2(new_n79_), .ZN(new_n14732_));
  OAI21_X1   g14637(.A1(new_n14732_), .A2(new_n14731_), .B(new_n72_), .ZN(new_n14733_));
  NAND2_X1   g14638(.A1(new_n14733_), .A2(new_n101_), .ZN(new_n14734_));
  XOR2_X1    g14639(.A1(new_n11246_), .A2(new_n14734_), .Z(new_n14735_));
  XOR2_X1    g14640(.A1(new_n14735_), .A2(new_n14730_), .Z(new_n14736_));
  AND2_X2    g14641(.A1(new_n14735_), .A2(new_n14729_), .Z(new_n14737_));
  NOR2_X1    g14642(.A1(new_n14735_), .A2(new_n14729_), .ZN(new_n14738_));
  NOR2_X1    g14643(.A1(new_n14737_), .A2(new_n14738_), .ZN(new_n14739_));
  MUX2_X1    g14644(.I0(new_n14739_), .I1(new_n14736_), .S(new_n14724_), .Z(new_n14740_));
  OAI22_X1   g14645(.A1(new_n10633_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n11264_), .ZN(new_n14741_));
  OAI21_X1   g14646(.A1(new_n10631_), .A2(new_n1128_), .B(new_n14741_), .ZN(new_n14742_));
  AOI21_X1   g14647(.A1(new_n14742_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n14743_));
  XOR2_X1    g14648(.A1(new_n11445_), .A2(new_n14743_), .Z(new_n14744_));
  NOR2_X1    g14649(.A1(new_n14744_), .A2(new_n14740_), .ZN(new_n14745_));
  INV_X1     g14650(.I(new_n14745_), .ZN(new_n14746_));
  NOR2_X1    g14651(.A1(new_n14723_), .A2(new_n14746_), .ZN(new_n14747_));
  NAND2_X1   g14652(.A1(new_n14723_), .A2(new_n14746_), .ZN(new_n14748_));
  INV_X1     g14653(.I(new_n14748_), .ZN(new_n14749_));
  OAI21_X1   g14654(.A1(new_n14749_), .A2(new_n14747_), .B(new_n14469_), .ZN(new_n14750_));
  INV_X1     g14655(.I(new_n14747_), .ZN(new_n14751_));
  NAND3_X1   g14656(.A1(new_n14751_), .A2(new_n14748_), .A3(new_n14470_), .ZN(new_n14752_));
  OAI22_X1   g14657(.A1(new_n10870_), .A2(new_n1239_), .B1(new_n4981_), .B2(new_n10861_), .ZN(new_n14753_));
  AOI21_X1   g14658(.A1(new_n14753_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n14754_));
  XOR2_X1    g14659(.A1(new_n11648_), .A2(new_n14754_), .Z(new_n14755_));
  AOI21_X1   g14660(.A1(new_n14750_), .A2(new_n14752_), .B(new_n14755_), .ZN(new_n14756_));
  OAI21_X1   g14661(.A1(new_n14438_), .A2(new_n14483_), .B(new_n14756_), .ZN(new_n14757_));
  AOI21_X1   g14662(.A1(new_n14751_), .A2(new_n14748_), .B(new_n14470_), .ZN(new_n14758_));
  NOR3_X1    g14663(.A1(new_n14749_), .A2(new_n14469_), .A3(new_n14747_), .ZN(new_n14759_));
  INV_X1     g14664(.I(new_n14755_), .ZN(new_n14760_));
  OAI21_X1   g14665(.A1(new_n14758_), .A2(new_n14759_), .B(new_n14760_), .ZN(new_n14761_));
  NAND3_X1   g14666(.A1(new_n14761_), .A2(new_n14482_), .A3(new_n14480_), .ZN(new_n14762_));
  AOI21_X1   g14667(.A1(new_n14757_), .A2(new_n14762_), .B(new_n14477_), .ZN(new_n14763_));
  INV_X1     g14668(.I(new_n14763_), .ZN(new_n14764_));
  NAND3_X1   g14669(.A1(new_n14757_), .A2(new_n14762_), .A3(new_n14477_), .ZN(new_n14765_));
  OAI22_X1   g14670(.A1(new_n10619_), .A2(new_n5398_), .B1(new_n5336_), .B2(new_n10885_), .ZN(new_n14766_));
  AOI21_X1   g14671(.A1(new_n14766_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n14767_));
  XOR2_X1    g14672(.A1(new_n12074_), .A2(new_n14767_), .Z(new_n14768_));
  AOI21_X1   g14673(.A1(new_n14764_), .A2(new_n14765_), .B(new_n14768_), .ZN(new_n14769_));
  NAND2_X1   g14674(.A1(new_n14718_), .A2(new_n14769_), .ZN(new_n14770_));
  INV_X1     g14675(.I(new_n14477_), .ZN(new_n14771_));
  AOI21_X1   g14676(.A1(new_n14482_), .A2(new_n14480_), .B(new_n14761_), .ZN(new_n14772_));
  NOR3_X1    g14677(.A1(new_n14756_), .A2(new_n14438_), .A3(new_n14483_), .ZN(new_n14773_));
  NOR3_X1    g14678(.A1(new_n14772_), .A2(new_n14771_), .A3(new_n14773_), .ZN(new_n14774_));
  INV_X1     g14679(.I(new_n14768_), .ZN(new_n14775_));
  OAI21_X1   g14680(.A1(new_n14774_), .A2(new_n14763_), .B(new_n14775_), .ZN(new_n14776_));
  NAND2_X1   g14681(.A1(new_n14493_), .A2(new_n14776_), .ZN(new_n14777_));
  AOI21_X1   g14682(.A1(new_n14770_), .A2(new_n14777_), .B(new_n14492_), .ZN(new_n14778_));
  NAND3_X1   g14683(.A1(new_n14770_), .A2(new_n14777_), .A3(new_n14492_), .ZN(new_n14779_));
  INV_X1     g14684(.I(new_n14779_), .ZN(new_n14780_));
  OAI22_X1   g14685(.A1(new_n10606_), .A2(new_n1620_), .B1(new_n5420_), .B2(new_n10901_), .ZN(new_n14781_));
  AOI21_X1   g14686(.A1(new_n14781_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n14782_));
  XOR2_X1    g14687(.A1(new_n12211_), .A2(new_n14782_), .Z(new_n14783_));
  INV_X1     g14688(.I(new_n14783_), .ZN(new_n14784_));
  OAI21_X1   g14689(.A1(new_n14780_), .A2(new_n14778_), .B(new_n14784_), .ZN(new_n14785_));
  NOR2_X1    g14690(.A1(new_n14717_), .A2(new_n14785_), .ZN(new_n14786_));
  AOI21_X1   g14691(.A1(new_n14507_), .A2(new_n14502_), .B(new_n14181_), .ZN(new_n14787_));
  OAI21_X1   g14692(.A1(new_n14787_), .A2(new_n14179_), .B(new_n14183_), .ZN(new_n14788_));
  INV_X1     g14693(.I(new_n14492_), .ZN(new_n14789_));
  NOR2_X1    g14694(.A1(new_n14493_), .A2(new_n14776_), .ZN(new_n14790_));
  NOR2_X1    g14695(.A1(new_n14718_), .A2(new_n14769_), .ZN(new_n14791_));
  OAI21_X1   g14696(.A1(new_n14791_), .A2(new_n14790_), .B(new_n14789_), .ZN(new_n14792_));
  AOI21_X1   g14697(.A1(new_n14792_), .A2(new_n14779_), .B(new_n14783_), .ZN(new_n14793_));
  NOR2_X1    g14698(.A1(new_n14788_), .A2(new_n14793_), .ZN(new_n14794_));
  OAI21_X1   g14699(.A1(new_n14786_), .A2(new_n14794_), .B(new_n14507_), .ZN(new_n14795_));
  NAND2_X1   g14700(.A1(new_n14788_), .A2(new_n14793_), .ZN(new_n14796_));
  NAND2_X1   g14701(.A1(new_n14717_), .A2(new_n14785_), .ZN(new_n14797_));
  NAND3_X1   g14702(.A1(new_n14797_), .A2(new_n14796_), .A3(new_n14501_), .ZN(new_n14798_));
  OAI22_X1   g14703(.A1(new_n10589_), .A2(new_n643_), .B1(new_n12623_), .B2(new_n5967_), .ZN(new_n14799_));
  AOI21_X1   g14704(.A1(new_n14799_), .A2(new_n279_), .B(new_n643_), .ZN(new_n14800_));
  XOR2_X1    g14705(.A1(new_n12622_), .A2(new_n14800_), .Z(new_n14801_));
  AOI21_X1   g14706(.A1(new_n14795_), .A2(new_n14798_), .B(new_n14801_), .ZN(new_n14802_));
  NAND2_X1   g14707(.A1(new_n14522_), .A2(new_n14802_), .ZN(new_n14803_));
  AOI21_X1   g14708(.A1(new_n14797_), .A2(new_n14796_), .B(new_n14501_), .ZN(new_n14804_));
  NOR3_X1    g14709(.A1(new_n14786_), .A2(new_n14794_), .A3(new_n14507_), .ZN(new_n14805_));
  INV_X1     g14710(.I(new_n14801_), .ZN(new_n14806_));
  OAI21_X1   g14711(.A1(new_n14804_), .A2(new_n14805_), .B(new_n14806_), .ZN(new_n14807_));
  NAND2_X1   g14712(.A1(new_n14807_), .A2(new_n14539_), .ZN(new_n14808_));
  AOI21_X1   g14713(.A1(new_n14808_), .A2(new_n14803_), .B(new_n14520_), .ZN(new_n14809_));
  INV_X1     g14714(.I(new_n14520_), .ZN(new_n14810_));
  NOR2_X1    g14715(.A1(new_n14807_), .A2(new_n14539_), .ZN(new_n14811_));
  NOR2_X1    g14716(.A1(new_n14522_), .A2(new_n14802_), .ZN(new_n14812_));
  NOR3_X1    g14717(.A1(new_n14811_), .A2(new_n14812_), .A3(new_n14810_), .ZN(new_n14813_));
  OAI22_X1   g14718(.A1(new_n10583_), .A2(new_n1078_), .B1(new_n6757_), .B2(new_n10928_), .ZN(new_n14814_));
  AOI21_X1   g14719(.A1(new_n14814_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n14815_));
  XNOR2_X1   g14720(.A1(new_n13378_), .A2(new_n14815_), .ZN(new_n14816_));
  INV_X1     g14721(.I(new_n14816_), .ZN(new_n14817_));
  OAI21_X1   g14722(.A1(new_n14809_), .A2(new_n14813_), .B(new_n14817_), .ZN(new_n14818_));
  NOR2_X1    g14723(.A1(new_n14715_), .A2(new_n14818_), .ZN(new_n14819_));
  AOI21_X1   g14724(.A1(new_n14542_), .A2(new_n14538_), .B(new_n14209_), .ZN(new_n14820_));
  OAI21_X1   g14725(.A1(new_n14820_), .A2(new_n14224_), .B(new_n14212_), .ZN(new_n14821_));
  OAI21_X1   g14726(.A1(new_n14811_), .A2(new_n14812_), .B(new_n14810_), .ZN(new_n14822_));
  NAND3_X1   g14727(.A1(new_n14808_), .A2(new_n14803_), .A3(new_n14520_), .ZN(new_n14823_));
  AOI21_X1   g14728(.A1(new_n14822_), .A2(new_n14823_), .B(new_n14816_), .ZN(new_n14824_));
  NOR2_X1    g14729(.A1(new_n14821_), .A2(new_n14824_), .ZN(new_n14825_));
  OAI21_X1   g14730(.A1(new_n14819_), .A2(new_n14825_), .B(new_n14538_), .ZN(new_n14826_));
  NAND2_X1   g14731(.A1(new_n14821_), .A2(new_n14824_), .ZN(new_n14827_));
  NAND2_X1   g14732(.A1(new_n14715_), .A2(new_n14818_), .ZN(new_n14828_));
  NAND3_X1   g14733(.A1(new_n14828_), .A2(new_n14827_), .A3(new_n14712_), .ZN(new_n14829_));
  NAND2_X1   g14734(.A1(new_n14826_), .A2(new_n14829_), .ZN(new_n14830_));
  OAI22_X1   g14735(.A1(new_n2718_), .A2(new_n10938_), .B1(new_n10952_), .B2(new_n7836_), .ZN(new_n14831_));
  OAI21_X1   g14736(.A1(new_n10577_), .A2(new_n2495_), .B(new_n14831_), .ZN(new_n14832_));
  AOI21_X1   g14737(.A1(new_n14832_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n14833_));
  XOR2_X1    g14738(.A1(new_n13544_), .A2(new_n14833_), .Z(new_n14834_));
  INV_X1     g14739(.I(new_n14834_), .ZN(new_n14835_));
  NAND3_X1   g14740(.A1(new_n14711_), .A2(new_n14830_), .A3(new_n14835_), .ZN(new_n14836_));
  NAND2_X1   g14741(.A1(new_n14830_), .A2(new_n14835_), .ZN(new_n14837_));
  NAND2_X1   g14742(.A1(new_n14837_), .A2(new_n14710_), .ZN(new_n14838_));
  AOI21_X1   g14743(.A1(new_n14838_), .A2(new_n14836_), .B(new_n14553_), .ZN(new_n14839_));
  OAI21_X1   g14744(.A1(new_n14545_), .A2(new_n14546_), .B(new_n14549_), .ZN(new_n14840_));
  NOR2_X1    g14745(.A1(new_n14837_), .A2(new_n14710_), .ZN(new_n14841_));
  AOI21_X1   g14746(.A1(new_n14830_), .A2(new_n14835_), .B(new_n14711_), .ZN(new_n14842_));
  NOR3_X1    g14747(.A1(new_n14842_), .A2(new_n14841_), .A3(new_n14840_), .ZN(new_n14843_));
  OAI22_X1   g14748(.A1(new_n10570_), .A2(new_n8830_), .B1(new_n3042_), .B2(new_n10961_), .ZN(new_n14844_));
  OAI21_X1   g14749(.A1(new_n10564_), .A2(new_n3040_), .B(new_n14844_), .ZN(new_n14845_));
  AOI21_X1   g14750(.A1(new_n14845_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n14846_));
  XOR2_X1    g14751(.A1(new_n10976_), .A2(new_n14846_), .Z(new_n14847_));
  INV_X1     g14752(.I(new_n14847_), .ZN(new_n14848_));
  OAI21_X1   g14753(.A1(new_n14843_), .A2(new_n14839_), .B(new_n14848_), .ZN(new_n14849_));
  NOR2_X1    g14754(.A1(new_n14708_), .A2(new_n14849_), .ZN(new_n14850_));
  OAI22_X1   g14755(.A1(new_n14087_), .A2(new_n14084_), .B1(new_n14240_), .B2(new_n14242_), .ZN(new_n14851_));
  OAI21_X1   g14756(.A1(new_n14842_), .A2(new_n14841_), .B(new_n14840_), .ZN(new_n14852_));
  NAND3_X1   g14757(.A1(new_n14838_), .A2(new_n14836_), .A3(new_n14553_), .ZN(new_n14853_));
  AOI21_X1   g14758(.A1(new_n14852_), .A2(new_n14853_), .B(new_n14847_), .ZN(new_n14854_));
  NOR2_X1    g14759(.A1(new_n14851_), .A2(new_n14854_), .ZN(new_n14855_));
  OAI21_X1   g14760(.A1(new_n14850_), .A2(new_n14855_), .B(new_n14562_), .ZN(new_n14856_));
  NOR3_X1    g14761(.A1(new_n14564_), .A2(new_n14563_), .A3(new_n14565_), .ZN(new_n14857_));
  NAND2_X1   g14762(.A1(new_n14851_), .A2(new_n14854_), .ZN(new_n14858_));
  NAND2_X1   g14763(.A1(new_n14708_), .A2(new_n14849_), .ZN(new_n14859_));
  NAND3_X1   g14764(.A1(new_n14859_), .A2(new_n14858_), .A3(new_n14857_), .ZN(new_n14860_));
  NOR2_X1    g14765(.A1(new_n14579_), .A2(new_n14587_), .ZN(new_n14861_));
  NOR2_X1    g14766(.A1(new_n14588_), .A2(new_n14270_), .ZN(new_n14862_));
  NAND2_X1   g14767(.A1(new_n14588_), .A2(new_n14270_), .ZN(new_n14863_));
  AOI21_X1   g14768(.A1(new_n14252_), .A2(new_n14863_), .B(new_n14862_), .ZN(new_n14864_));
  NAND2_X1   g14769(.A1(new_n14250_), .A2(new_n14864_), .ZN(new_n14865_));
  NOR2_X1    g14770(.A1(new_n14582_), .A2(new_n14262_), .ZN(new_n14866_));
  NOR2_X1    g14771(.A1(new_n14866_), .A2(new_n14584_), .ZN(new_n14867_));
  NAND2_X1   g14772(.A1(new_n4564_), .A2(new_n4406_), .ZN(new_n14868_));
  NOR2_X1    g14773(.A1(new_n14258_), .A2(new_n87_), .ZN(new_n14869_));
  AOI21_X1   g14774(.A1(new_n14869_), .A2(new_n14868_), .B(new_n82_), .ZN(new_n14870_));
  NAND2_X1   g14775(.A1(new_n5001_), .A2(new_n14870_), .ZN(new_n14871_));
  XOR2_X1    g14776(.A1(new_n4526_), .A2(\a[29] ), .Z(new_n14872_));
  XOR2_X1    g14777(.A1(new_n14871_), .A2(new_n14872_), .Z(new_n14873_));
  NOR2_X1    g14778(.A1(new_n14873_), .A2(new_n14261_), .ZN(new_n14874_));
  INV_X1     g14779(.I(new_n14872_), .ZN(new_n14875_));
  NOR2_X1    g14780(.A1(new_n14871_), .A2(new_n14875_), .ZN(new_n14876_));
  INV_X1     g14781(.I(new_n14876_), .ZN(new_n14877_));
  NAND2_X1   g14782(.A1(new_n14871_), .A2(new_n14875_), .ZN(new_n14878_));
  AOI21_X1   g14783(.A1(new_n14877_), .A2(new_n14878_), .B(new_n14262_), .ZN(new_n14879_));
  NOR2_X1    g14784(.A1(new_n14874_), .A2(new_n14879_), .ZN(new_n14880_));
  NOR2_X1    g14785(.A1(new_n14880_), .A2(new_n14867_), .ZN(new_n14881_));
  XOR2_X1    g14786(.A1(new_n14865_), .A2(new_n14881_), .Z(new_n14882_));
  NOR2_X1    g14787(.A1(new_n14882_), .A2(new_n14861_), .ZN(new_n14883_));
  NAND2_X1   g14788(.A1(new_n14882_), .A2(new_n14861_), .ZN(new_n14884_));
  INV_X1     g14789(.I(new_n14884_), .ZN(new_n14885_));
  NOR2_X1    g14790(.A1(new_n14885_), .A2(new_n14883_), .ZN(new_n14886_));
  NOR2_X1    g14791(.A1(new_n14886_), .A2(new_n14274_), .ZN(new_n14887_));
  INV_X1     g14792(.I(new_n14886_), .ZN(new_n14888_));
  NOR2_X1    g14793(.A1(new_n14888_), .A2(new_n14276_), .ZN(new_n14889_));
  OAI21_X1   g14794(.A1(new_n14889_), .A2(new_n14887_), .B(new_n14596_), .ZN(new_n14890_));
  XOR2_X1    g14795(.A1(new_n14575_), .A2(new_n14890_), .Z(new_n14891_));
  OAI22_X1   g14796(.A1(new_n14276_), .A2(new_n9408_), .B1(new_n9405_), .B2(new_n14594_), .ZN(new_n14892_));
  OAI21_X1   g14797(.A1(new_n14886_), .A2(new_n3456_), .B(new_n14892_), .ZN(new_n14893_));
  AOI21_X1   g14798(.A1(new_n14893_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n14894_));
  XOR2_X1    g14799(.A1(new_n14891_), .A2(new_n14894_), .Z(new_n14895_));
  NAND3_X1   g14800(.A1(new_n14856_), .A2(new_n14860_), .A3(new_n14895_), .ZN(new_n14896_));
  AOI21_X1   g14801(.A1(new_n14859_), .A2(new_n14858_), .B(new_n14857_), .ZN(new_n14897_));
  NOR3_X1    g14802(.A1(new_n14850_), .A2(new_n14855_), .A3(new_n14562_), .ZN(new_n14898_));
  INV_X1     g14803(.I(new_n14895_), .ZN(new_n14899_));
  OAI21_X1   g14804(.A1(new_n14898_), .A2(new_n14897_), .B(new_n14899_), .ZN(new_n14900_));
  NAND2_X1   g14805(.A1(new_n14900_), .A2(new_n14896_), .ZN(new_n14901_));
  XOR2_X1    g14806(.A1(new_n14572_), .A2(new_n14608_), .Z(new_n14902_));
  NAND3_X1   g14807(.A1(new_n14902_), .A2(new_n14609_), .A3(new_n14901_), .ZN(new_n14903_));
  NOR2_X1    g14808(.A1(new_n14898_), .A2(new_n14897_), .ZN(new_n14904_));
  NAND2_X1   g14809(.A1(new_n14572_), .A2(new_n14608_), .ZN(new_n14905_));
  AND2_X2    g14810(.A1(new_n14903_), .A2(new_n14905_), .Z(new_n14906_));
  XOR2_X1    g14811(.A1(new_n14906_), .A2(new_n14702_), .Z(new_n14907_));
  XOR2_X1    g14812(.A1(new_n14620_), .A2(new_n14907_), .Z(\result[2] ));
  AOI21_X1   g14813(.A1(new_n14616_), .A2(new_n14617_), .B(new_n14610_), .ZN(new_n14909_));
  NOR3_X1    g14814(.A1(new_n14411_), .A2(new_n14407_), .A3(new_n14614_), .ZN(new_n14910_));
  XOR2_X1    g14815(.A1(new_n14404_), .A2(new_n14422_), .Z(new_n14911_));
  NOR2_X1    g14816(.A1(new_n14911_), .A2(new_n14702_), .ZN(new_n14912_));
  OAI21_X1   g14817(.A1(new_n14910_), .A2(new_n14909_), .B(new_n14912_), .ZN(new_n14913_));
  XOR2_X1    g14818(.A1(new_n14906_), .A2(new_n14429_), .Z(new_n14914_));
  NOR2_X1    g14819(.A1(new_n14904_), .A2(new_n14899_), .ZN(new_n14915_));
  INV_X1     g14820(.I(new_n14915_), .ZN(new_n14916_));
  NAND3_X1   g14821(.A1(new_n14573_), .A2(new_n14900_), .A3(new_n14896_), .ZN(new_n14917_));
  INV_X1     g14822(.I(new_n14917_), .ZN(new_n14918_));
  AOI21_X1   g14823(.A1(new_n14900_), .A2(new_n14896_), .B(new_n14573_), .ZN(new_n14919_));
  NOR2_X1    g14824(.A1(new_n14919_), .A2(new_n14608_), .ZN(new_n14920_));
  NOR2_X1    g14825(.A1(new_n14920_), .A2(new_n14918_), .ZN(new_n14921_));
  AOI21_X1   g14826(.A1(new_n14852_), .A2(new_n14853_), .B(new_n14562_), .ZN(new_n14922_));
  NOR3_X1    g14827(.A1(new_n14843_), .A2(new_n14839_), .A3(new_n14857_), .ZN(new_n14923_));
  NOR2_X1    g14828(.A1(new_n14923_), .A2(new_n14847_), .ZN(new_n14924_));
  AOI21_X1   g14829(.A1(new_n14924_), .A2(new_n14708_), .B(new_n14922_), .ZN(new_n14925_));
  NAND2_X1   g14830(.A1(new_n14830_), .A2(new_n14553_), .ZN(new_n14926_));
  NAND3_X1   g14831(.A1(new_n14826_), .A2(new_n14829_), .A3(new_n14840_), .ZN(new_n14927_));
  NAND3_X1   g14832(.A1(new_n14927_), .A2(new_n14710_), .A3(new_n14835_), .ZN(new_n14928_));
  NAND2_X1   g14833(.A1(new_n14928_), .A2(new_n14926_), .ZN(new_n14929_));
  NAND2_X1   g14834(.A1(new_n14795_), .A2(new_n14798_), .ZN(new_n14930_));
  NAND2_X1   g14835(.A1(new_n14930_), .A2(new_n14520_), .ZN(new_n14931_));
  NAND3_X1   g14836(.A1(new_n14795_), .A2(new_n14798_), .A3(new_n14810_), .ZN(new_n14932_));
  NAND3_X1   g14837(.A1(new_n14539_), .A2(new_n14932_), .A3(new_n14806_), .ZN(new_n14933_));
  NAND2_X1   g14838(.A1(new_n14933_), .A2(new_n14931_), .ZN(new_n14934_));
  NAND2_X1   g14839(.A1(new_n14764_), .A2(new_n14765_), .ZN(new_n14935_));
  NOR3_X1    g14840(.A1(new_n14774_), .A2(new_n14763_), .A3(new_n14492_), .ZN(new_n14936_));
  NOR2_X1    g14841(.A1(new_n14936_), .A2(new_n14768_), .ZN(new_n14937_));
  AOI22_X1   g14842(.A1(new_n14937_), .A2(new_n14493_), .B1(new_n14492_), .B2(new_n14935_), .ZN(new_n14938_));
  INV_X1     g14843(.I(new_n14938_), .ZN(new_n14939_));
  OAI21_X1   g14844(.A1(new_n14758_), .A2(new_n14759_), .B(new_n14477_), .ZN(new_n14940_));
  NAND3_X1   g14845(.A1(new_n14750_), .A2(new_n14752_), .A3(new_n14771_), .ZN(new_n14941_));
  NAND4_X1   g14846(.A1(new_n14941_), .A2(new_n14482_), .A3(new_n14480_), .A4(new_n14760_), .ZN(new_n14942_));
  NAND2_X1   g14847(.A1(new_n14942_), .A2(new_n14940_), .ZN(new_n14943_));
  NOR2_X1    g14848(.A1(new_n14469_), .A2(new_n14740_), .ZN(new_n14944_));
  AOI21_X1   g14849(.A1(new_n14740_), .A2(new_n14469_), .B(new_n14744_), .ZN(new_n14945_));
  AND2_X2    g14850(.A1(new_n14723_), .A2(new_n14945_), .Z(new_n14946_));
  INV_X1     g14851(.I(new_n14737_), .ZN(new_n14947_));
  AOI21_X1   g14852(.A1(new_n14947_), .A2(new_n14724_), .B(new_n14738_), .ZN(new_n14948_));
  INV_X1     g14853(.I(new_n14948_), .ZN(new_n14949_));
  NAND2_X1   g14854(.A1(new_n14725_), .A2(new_n14728_), .ZN(new_n14950_));
  NAND2_X1   g14855(.A1(new_n10805_), .A2(new_n962_), .ZN(new_n14951_));
  AOI22_X1   g14856(.A1(new_n10817_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n10691_), .ZN(new_n14952_));
  AOI21_X1   g14857(.A1(new_n14951_), .A2(new_n14952_), .B(new_n82_), .ZN(new_n14953_));
  OAI21_X1   g14858(.A1(new_n11174_), .A2(new_n11171_), .B(new_n14953_), .ZN(new_n14954_));
  XNOR2_X1   g14859(.A1(new_n14950_), .A2(new_n14954_), .ZN(new_n14955_));
  INV_X1     g14860(.I(new_n14955_), .ZN(new_n14956_));
  OAI22_X1   g14861(.A1(new_n10646_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n11214_), .ZN(new_n14957_));
  OAI21_X1   g14862(.A1(new_n79_), .A2(new_n11264_), .B(new_n14957_), .ZN(new_n14958_));
  AOI21_X1   g14863(.A1(new_n14958_), .A2(new_n72_), .B(new_n79_), .ZN(new_n14959_));
  XOR2_X1    g14864(.A1(new_n11268_), .A2(new_n14959_), .Z(new_n14960_));
  XOR2_X1    g14865(.A1(new_n14960_), .A2(new_n14956_), .Z(new_n14961_));
  NAND2_X1   g14866(.A1(new_n14949_), .A2(new_n14961_), .ZN(new_n14962_));
  NOR2_X1    g14867(.A1(new_n14960_), .A2(new_n14956_), .ZN(new_n14963_));
  NAND2_X1   g14868(.A1(new_n14960_), .A2(new_n14956_), .ZN(new_n14964_));
  INV_X1     g14869(.I(new_n14964_), .ZN(new_n14965_));
  OAI21_X1   g14870(.A1(new_n14963_), .A2(new_n14965_), .B(new_n14948_), .ZN(new_n14966_));
  NAND2_X1   g14871(.A1(new_n14962_), .A2(new_n14966_), .ZN(new_n14967_));
  OAI22_X1   g14872(.A1(new_n10631_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10633_), .ZN(new_n14968_));
  OAI21_X1   g14873(.A1(new_n10844_), .A2(new_n1128_), .B(new_n14968_), .ZN(new_n14969_));
  AOI21_X1   g14874(.A1(new_n14969_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n14970_));
  XNOR2_X1   g14875(.A1(new_n11607_), .A2(new_n14970_), .ZN(new_n14971_));
  NAND2_X1   g14876(.A1(new_n14971_), .A2(new_n14967_), .ZN(new_n14972_));
  INV_X1     g14877(.I(new_n14972_), .ZN(new_n14973_));
  NOR2_X1    g14878(.A1(new_n14971_), .A2(new_n14967_), .ZN(new_n14974_));
  OAI22_X1   g14879(.A1(new_n14946_), .A2(new_n14944_), .B1(new_n14973_), .B2(new_n14974_), .ZN(new_n14975_));
  NOR2_X1    g14880(.A1(new_n14946_), .A2(new_n14944_), .ZN(new_n14976_));
  INV_X1     g14881(.I(new_n14971_), .ZN(new_n14977_));
  NOR2_X1    g14882(.A1(new_n14977_), .A2(new_n14967_), .ZN(new_n14978_));
  NAND2_X1   g14883(.A1(new_n14977_), .A2(new_n14967_), .ZN(new_n14979_));
  INV_X1     g14884(.I(new_n14979_), .ZN(new_n14980_));
  OAI21_X1   g14885(.A1(new_n14978_), .A2(new_n14980_), .B(new_n14976_), .ZN(new_n14981_));
  OAI22_X1   g14886(.A1(new_n11723_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n10868_), .ZN(new_n14982_));
  AOI21_X1   g14887(.A1(new_n14982_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n14983_));
  XOR2_X1    g14888(.A1(new_n11722_), .A2(new_n14983_), .Z(new_n14984_));
  NAND3_X1   g14889(.A1(new_n14981_), .A2(new_n14975_), .A3(new_n14984_), .ZN(new_n14985_));
  INV_X1     g14890(.I(new_n14985_), .ZN(new_n14986_));
  AOI21_X1   g14891(.A1(new_n14981_), .A2(new_n14975_), .B(new_n14984_), .ZN(new_n14987_));
  NOR2_X1    g14892(.A1(new_n14986_), .A2(new_n14987_), .ZN(new_n14988_));
  NOR2_X1    g14893(.A1(new_n14988_), .A2(new_n14943_), .ZN(new_n14989_));
  INV_X1     g14894(.I(new_n14989_), .ZN(new_n14990_));
  NAND2_X1   g14895(.A1(new_n14988_), .A2(new_n14943_), .ZN(new_n14991_));
  OAI22_X1   g14896(.A1(new_n12091_), .A2(new_n5336_), .B1(new_n5398_), .B2(new_n10611_), .ZN(new_n14992_));
  AOI21_X1   g14897(.A1(new_n14992_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n14993_));
  AND2_X2    g14898(.A1(new_n12090_), .A2(new_n14993_), .Z(new_n14994_));
  NOR2_X1    g14899(.A1(new_n12090_), .A2(new_n14993_), .ZN(new_n14995_));
  NOR2_X1    g14900(.A1(new_n14994_), .A2(new_n14995_), .ZN(new_n14996_));
  INV_X1     g14901(.I(new_n14996_), .ZN(new_n14997_));
  NAND3_X1   g14902(.A1(new_n14990_), .A2(new_n14991_), .A3(new_n14997_), .ZN(new_n14998_));
  INV_X1     g14903(.I(new_n14991_), .ZN(new_n14999_));
  OAI21_X1   g14904(.A1(new_n14999_), .A2(new_n14989_), .B(new_n14996_), .ZN(new_n15000_));
  NAND2_X1   g14905(.A1(new_n15000_), .A2(new_n14998_), .ZN(new_n15001_));
  NOR2_X1    g14906(.A1(new_n14939_), .A2(new_n15001_), .ZN(new_n15002_));
  NOR3_X1    g14907(.A1(new_n14999_), .A2(new_n14989_), .A3(new_n14996_), .ZN(new_n15003_));
  AOI21_X1   g14908(.A1(new_n14990_), .A2(new_n14991_), .B(new_n14997_), .ZN(new_n15004_));
  NOR2_X1    g14909(.A1(new_n15004_), .A2(new_n15003_), .ZN(new_n15005_));
  NOR2_X1    g14910(.A1(new_n15005_), .A2(new_n14938_), .ZN(new_n15006_));
  AOI22_X1   g14911(.A1(new_n12578_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n10600_), .ZN(new_n15007_));
  OAI21_X1   g14912(.A1(new_n15007_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n15008_));
  XNOR2_X1   g14913(.A1(new_n12576_), .A2(new_n15008_), .ZN(new_n15009_));
  INV_X1     g14914(.I(new_n15009_), .ZN(new_n15010_));
  NOR3_X1    g14915(.A1(new_n15002_), .A2(new_n15006_), .A3(new_n15010_), .ZN(new_n15011_));
  NAND2_X1   g14916(.A1(new_n15005_), .A2(new_n14938_), .ZN(new_n15012_));
  NAND2_X1   g14917(.A1(new_n14939_), .A2(new_n15001_), .ZN(new_n15013_));
  AOI21_X1   g14918(.A1(new_n15013_), .A2(new_n15012_), .B(new_n15009_), .ZN(new_n15014_));
  NOR2_X1    g14919(.A1(new_n15011_), .A2(new_n15014_), .ZN(new_n15015_));
  NOR2_X1    g14920(.A1(new_n14780_), .A2(new_n14778_), .ZN(new_n15016_));
  NAND3_X1   g14921(.A1(new_n14792_), .A2(new_n14779_), .A3(new_n14507_), .ZN(new_n15017_));
  NAND2_X1   g14922(.A1(new_n15017_), .A2(new_n14784_), .ZN(new_n15018_));
  OAI22_X1   g14923(.A1(new_n15018_), .A2(new_n14788_), .B1(new_n14507_), .B2(new_n15016_), .ZN(new_n15019_));
  NAND2_X1   g14924(.A1(new_n15019_), .A2(new_n15015_), .ZN(new_n15020_));
  NAND3_X1   g14925(.A1(new_n15013_), .A2(new_n15012_), .A3(new_n15009_), .ZN(new_n15021_));
  OAI21_X1   g14926(.A1(new_n15002_), .A2(new_n15006_), .B(new_n15010_), .ZN(new_n15022_));
  NAND2_X1   g14927(.A1(new_n15022_), .A2(new_n15021_), .ZN(new_n15023_));
  AOI21_X1   g14928(.A1(new_n14792_), .A2(new_n14779_), .B(new_n14507_), .ZN(new_n15024_));
  INV_X1     g14929(.I(new_n15018_), .ZN(new_n15025_));
  AOI21_X1   g14930(.A1(new_n15025_), .A2(new_n14717_), .B(new_n15024_), .ZN(new_n15026_));
  NAND2_X1   g14931(.A1(new_n15026_), .A2(new_n15023_), .ZN(new_n15027_));
  OAI22_X1   g14932(.A1(new_n10913_), .A2(new_n643_), .B1(new_n12768_), .B2(new_n5967_), .ZN(new_n15028_));
  AOI21_X1   g14933(.A1(new_n15028_), .A2(new_n279_), .B(new_n643_), .ZN(new_n15029_));
  XOR2_X1    g14934(.A1(new_n12767_), .A2(new_n15029_), .Z(new_n15030_));
  INV_X1     g14935(.I(new_n15030_), .ZN(new_n15031_));
  NAND3_X1   g14936(.A1(new_n15027_), .A2(new_n15031_), .A3(new_n15020_), .ZN(new_n15032_));
  NOR2_X1    g14937(.A1(new_n15026_), .A2(new_n15023_), .ZN(new_n15033_));
  NOR2_X1    g14938(.A1(new_n15019_), .A2(new_n15015_), .ZN(new_n15034_));
  OAI21_X1   g14939(.A1(new_n15033_), .A2(new_n15034_), .B(new_n15030_), .ZN(new_n15035_));
  NAND2_X1   g14940(.A1(new_n15035_), .A2(new_n15032_), .ZN(new_n15036_));
  NOR2_X1    g14941(.A1(new_n14934_), .A2(new_n15036_), .ZN(new_n15037_));
  NOR3_X1    g14942(.A1(new_n14804_), .A2(new_n14805_), .A3(new_n14520_), .ZN(new_n15038_));
  NOR2_X1    g14943(.A1(new_n15038_), .A2(new_n14801_), .ZN(new_n15039_));
  AOI22_X1   g14944(.A1(new_n15039_), .A2(new_n14539_), .B1(new_n14520_), .B2(new_n14930_), .ZN(new_n15040_));
  NOR3_X1    g14945(.A1(new_n15033_), .A2(new_n15030_), .A3(new_n15034_), .ZN(new_n15041_));
  AOI21_X1   g14946(.A1(new_n15027_), .A2(new_n15020_), .B(new_n15031_), .ZN(new_n15042_));
  NOR2_X1    g14947(.A1(new_n15041_), .A2(new_n15042_), .ZN(new_n15043_));
  NOR2_X1    g14948(.A1(new_n15040_), .A2(new_n15043_), .ZN(new_n15044_));
  INV_X1     g14949(.I(new_n13395_), .ZN(new_n15045_));
  AOI22_X1   g14950(.A1(new_n15045_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n10937_), .ZN(new_n15046_));
  OAI21_X1   g14951(.A1(new_n15046_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n15047_));
  NOR2_X1    g14952(.A1(new_n14014_), .A2(new_n15047_), .ZN(new_n15048_));
  INV_X1     g14953(.I(new_n15047_), .ZN(new_n15049_));
  NOR2_X1    g14954(.A1(new_n13394_), .A2(new_n15049_), .ZN(new_n15050_));
  NOR2_X1    g14955(.A1(new_n15048_), .A2(new_n15050_), .ZN(new_n15051_));
  INV_X1     g14956(.I(new_n15051_), .ZN(new_n15052_));
  NOR3_X1    g14957(.A1(new_n15044_), .A2(new_n15037_), .A3(new_n15052_), .ZN(new_n15053_));
  NAND3_X1   g14958(.A1(new_n15043_), .A2(new_n14931_), .A3(new_n14933_), .ZN(new_n15054_));
  NAND2_X1   g14959(.A1(new_n14934_), .A2(new_n15036_), .ZN(new_n15055_));
  AOI21_X1   g14960(.A1(new_n15055_), .A2(new_n15054_), .B(new_n15051_), .ZN(new_n15056_));
  NOR2_X1    g14961(.A1(new_n15053_), .A2(new_n15056_), .ZN(new_n15057_));
  AOI21_X1   g14962(.A1(new_n14822_), .A2(new_n14823_), .B(new_n14538_), .ZN(new_n15058_));
  INV_X1     g14963(.I(new_n15058_), .ZN(new_n15059_));
  NAND3_X1   g14964(.A1(new_n14822_), .A2(new_n14823_), .A3(new_n14538_), .ZN(new_n15060_));
  NAND2_X1   g14965(.A1(new_n15060_), .A2(new_n14817_), .ZN(new_n15061_));
  OAI21_X1   g14966(.A1(new_n15061_), .A2(new_n14821_), .B(new_n15059_), .ZN(new_n15062_));
  NAND2_X1   g14967(.A1(new_n15062_), .A2(new_n15057_), .ZN(new_n15063_));
  NAND3_X1   g14968(.A1(new_n15055_), .A2(new_n15054_), .A3(new_n15051_), .ZN(new_n15064_));
  OAI21_X1   g14969(.A1(new_n15044_), .A2(new_n15037_), .B(new_n15052_), .ZN(new_n15065_));
  NAND2_X1   g14970(.A1(new_n15065_), .A2(new_n15064_), .ZN(new_n15066_));
  NOR3_X1    g14971(.A1(new_n14809_), .A2(new_n14813_), .A3(new_n14712_), .ZN(new_n15067_));
  NOR2_X1    g14972(.A1(new_n15067_), .A2(new_n14816_), .ZN(new_n15068_));
  AOI21_X1   g14973(.A1(new_n15068_), .A2(new_n14715_), .B(new_n15058_), .ZN(new_n15069_));
  NAND2_X1   g14974(.A1(new_n15069_), .A2(new_n15066_), .ZN(new_n15070_));
  INV_X1     g14975(.I(new_n14053_), .ZN(new_n15071_));
  INV_X1     g14976(.I(new_n14054_), .ZN(new_n15072_));
  AOI22_X1   g14977(.A1(new_n15072_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n10962_), .ZN(new_n15073_));
  OAI21_X1   g14978(.A1(new_n15073_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n15074_));
  NOR2_X1    g14979(.A1(new_n15071_), .A2(new_n15074_), .ZN(new_n15075_));
  INV_X1     g14980(.I(new_n15074_), .ZN(new_n15076_));
  NOR2_X1    g14981(.A1(new_n14053_), .A2(new_n15076_), .ZN(new_n15077_));
  NOR2_X1    g14982(.A1(new_n15075_), .A2(new_n15077_), .ZN(new_n15078_));
  INV_X1     g14983(.I(new_n15078_), .ZN(new_n15079_));
  NAND3_X1   g14984(.A1(new_n15063_), .A2(new_n15070_), .A3(new_n15079_), .ZN(new_n15080_));
  NOR2_X1    g14985(.A1(new_n15069_), .A2(new_n15066_), .ZN(new_n15081_));
  NOR2_X1    g14986(.A1(new_n15062_), .A2(new_n15057_), .ZN(new_n15082_));
  OAI21_X1   g14987(.A1(new_n15082_), .A2(new_n15081_), .B(new_n15078_), .ZN(new_n15083_));
  NAND2_X1   g14988(.A1(new_n15083_), .A2(new_n15080_), .ZN(new_n15084_));
  NOR2_X1    g14989(.A1(new_n14929_), .A2(new_n15084_), .ZN(new_n15085_));
  INV_X1     g14990(.I(new_n15085_), .ZN(new_n15086_));
  NAND2_X1   g14991(.A1(new_n14929_), .A2(new_n15084_), .ZN(new_n15087_));
  AOI22_X1   g14992(.A1(new_n14281_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n14274_), .ZN(new_n15088_));
  OAI21_X1   g14993(.A1(new_n15088_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n15089_));
  XOR2_X1    g14994(.A1(new_n14280_), .A2(new_n15089_), .Z(new_n15090_));
  NAND3_X1   g14995(.A1(new_n15086_), .A2(new_n15087_), .A3(new_n15090_), .ZN(new_n15091_));
  INV_X1     g14996(.I(new_n15087_), .ZN(new_n15092_));
  INV_X1     g14997(.I(new_n15090_), .ZN(new_n15093_));
  OAI21_X1   g14998(.A1(new_n15092_), .A2(new_n15085_), .B(new_n15093_), .ZN(new_n15094_));
  NAND2_X1   g14999(.A1(new_n15094_), .A2(new_n15091_), .ZN(new_n15095_));
  XOR2_X1    g15000(.A1(new_n14925_), .A2(new_n15095_), .Z(new_n15096_));
  INV_X1     g15001(.I(new_n14861_), .ZN(new_n15097_));
  AOI21_X1   g15002(.A1(new_n14867_), .A2(new_n14880_), .B(new_n15097_), .ZN(new_n15098_));
  NAND3_X1   g15003(.A1(new_n14250_), .A2(new_n14864_), .A3(new_n15098_), .ZN(new_n15099_));
  INV_X1     g15004(.I(new_n15099_), .ZN(new_n15100_));
  NOR2_X1    g15005(.A1(new_n15100_), .A2(new_n14881_), .ZN(new_n15101_));
  NOR3_X1    g15006(.A1(new_n92_), .A2(new_n83_), .A3(new_n960_), .ZN(new_n15102_));
  NAND2_X1   g15007(.A1(new_n4610_), .A2(new_n15102_), .ZN(new_n15103_));
  INV_X1     g15008(.I(new_n15103_), .ZN(new_n15104_));
  NAND2_X1   g15009(.A1(new_n14878_), .A2(new_n14262_), .ZN(new_n15105_));
  NAND2_X1   g15010(.A1(new_n15105_), .A2(new_n14877_), .ZN(new_n15106_));
  XOR2_X1    g15011(.A1(new_n15106_), .A2(new_n15104_), .Z(new_n15107_));
  NOR2_X1    g15012(.A1(new_n15101_), .A2(new_n15107_), .ZN(new_n15108_));
  INV_X1     g15013(.I(new_n15101_), .ZN(new_n15109_));
  NOR2_X1    g15014(.A1(new_n15106_), .A2(new_n15103_), .ZN(new_n15110_));
  INV_X1     g15015(.I(new_n15110_), .ZN(new_n15111_));
  NAND2_X1   g15016(.A1(new_n15106_), .A2(new_n15103_), .ZN(new_n15112_));
  AOI21_X1   g15017(.A1(new_n15111_), .A2(new_n15112_), .B(new_n15109_), .ZN(new_n15113_));
  NOR2_X1    g15018(.A1(new_n15113_), .A2(new_n15108_), .ZN(new_n15114_));
  INV_X1     g15019(.I(new_n15114_), .ZN(new_n15115_));
  NOR2_X1    g15020(.A1(new_n14575_), .A2(new_n14597_), .ZN(new_n15116_));
  NAND2_X1   g15021(.A1(new_n14575_), .A2(new_n14598_), .ZN(new_n15117_));
  OAI21_X1   g15022(.A1(new_n14886_), .A2(new_n15116_), .B(new_n15117_), .ZN(new_n15118_));
  NOR2_X1    g15023(.A1(new_n15118_), .A2(new_n14888_), .ZN(new_n15119_));
  AOI21_X1   g15024(.A1(new_n15116_), .A2(new_n15117_), .B(new_n14886_), .ZN(new_n15120_));
  OR2_X2     g15025(.A1(new_n15119_), .A2(new_n15120_), .Z(new_n15121_));
  NAND2_X1   g15026(.A1(new_n15118_), .A2(new_n14886_), .ZN(new_n15122_));
  NAND3_X1   g15027(.A1(new_n15116_), .A2(new_n15117_), .A3(new_n14888_), .ZN(new_n15123_));
  AOI21_X1   g15028(.A1(new_n15122_), .A2(new_n15123_), .B(new_n15115_), .ZN(new_n15124_));
  AOI21_X1   g15029(.A1(new_n15121_), .A2(new_n15115_), .B(new_n15124_), .ZN(new_n15125_));
  NOR2_X1    g15030(.A1(new_n14886_), .A2(new_n14594_), .ZN(new_n15126_));
  INV_X1     g15031(.I(new_n15126_), .ZN(new_n15127_));
  AOI22_X1   g15032(.A1(new_n15127_), .A2(new_n9433_), .B1(new_n3455_), .B2(new_n15115_), .ZN(new_n15128_));
  OAI21_X1   g15033(.A1(new_n15128_), .A2(\a[2] ), .B(new_n3411_), .ZN(new_n15129_));
  XNOR2_X1   g15034(.A1(new_n15125_), .A2(new_n15129_), .ZN(new_n15130_));
  NOR2_X1    g15035(.A1(new_n15096_), .A2(new_n15130_), .ZN(new_n15131_));
  INV_X1     g15036(.I(new_n15131_), .ZN(new_n15132_));
  AOI21_X1   g15037(.A1(new_n14429_), .A2(new_n14921_), .B(new_n15132_), .ZN(new_n15133_));
  OAI21_X1   g15038(.A1(new_n14919_), .A2(new_n14608_), .B(new_n14917_), .ZN(new_n15134_));
  NOR3_X1    g15039(.A1(new_n14702_), .A2(new_n15134_), .A3(new_n15131_), .ZN(new_n15135_));
  OAI21_X1   g15040(.A1(new_n15135_), .A2(new_n15133_), .B(new_n14916_), .ZN(new_n15136_));
  OAI21_X1   g15041(.A1(new_n14702_), .A2(new_n15134_), .B(new_n15131_), .ZN(new_n15137_));
  NAND3_X1   g15042(.A1(new_n14429_), .A2(new_n14921_), .A3(new_n15132_), .ZN(new_n15138_));
  NAND3_X1   g15043(.A1(new_n15137_), .A2(new_n15138_), .A3(new_n14915_), .ZN(new_n15139_));
  NAND2_X1   g15044(.A1(new_n15136_), .A2(new_n15139_), .ZN(new_n15140_));
  OAI21_X1   g15045(.A1(new_n14913_), .A2(new_n14914_), .B(new_n15140_), .ZN(new_n15141_));
  AOI21_X1   g15046(.A1(new_n15137_), .A2(new_n15138_), .B(new_n14915_), .ZN(new_n15142_));
  NOR3_X1    g15047(.A1(new_n15135_), .A2(new_n15133_), .A3(new_n14916_), .ZN(new_n15143_));
  NOR2_X1    g15048(.A1(new_n15143_), .A2(new_n15142_), .ZN(new_n15144_));
  NAND3_X1   g15049(.A1(new_n15144_), .A2(new_n14620_), .A3(new_n14907_), .ZN(new_n15145_));
  NAND2_X1   g15050(.A1(new_n15141_), .A2(new_n15145_), .ZN(\result[3] ));
  NAND2_X1   g15051(.A1(new_n14620_), .A2(new_n14907_), .ZN(new_n15147_));
  NAND3_X1   g15052(.A1(new_n14404_), .A2(new_n14082_), .A3(new_n14427_), .ZN(new_n15148_));
  AOI21_X1   g15053(.A1(new_n15148_), .A2(new_n14426_), .B(new_n15134_), .ZN(new_n15149_));
  NOR2_X1    g15054(.A1(new_n14916_), .A2(new_n15096_), .ZN(new_n15150_));
  AOI21_X1   g15055(.A1(new_n14916_), .A2(new_n15096_), .B(new_n15130_), .ZN(new_n15151_));
  AOI21_X1   g15056(.A1(new_n15149_), .A2(new_n15151_), .B(new_n15150_), .ZN(new_n15152_));
  INV_X1     g15057(.I(new_n14922_), .ZN(new_n15153_));
  NAND3_X1   g15058(.A1(new_n14852_), .A2(new_n14853_), .A3(new_n14562_), .ZN(new_n15154_));
  NAND3_X1   g15059(.A1(new_n14708_), .A2(new_n14848_), .A3(new_n15154_), .ZN(new_n15155_));
  NAND2_X1   g15060(.A1(new_n15155_), .A2(new_n15153_), .ZN(new_n15156_));
  INV_X1     g15061(.I(new_n15095_), .ZN(new_n15157_));
  INV_X1     g15062(.I(new_n15091_), .ZN(new_n15158_));
  INV_X1     g15063(.I(new_n15084_), .ZN(new_n15159_));
  INV_X1     g15064(.I(new_n15083_), .ZN(new_n15160_));
  INV_X1     g15065(.I(new_n14943_), .ZN(new_n15161_));
  INV_X1     g15066(.I(new_n14987_), .ZN(new_n15162_));
  NAND2_X1   g15067(.A1(new_n15162_), .A2(new_n14985_), .ZN(new_n15163_));
  INV_X1     g15068(.I(new_n14974_), .ZN(new_n15164_));
  OAI21_X1   g15069(.A1(new_n14946_), .A2(new_n14944_), .B(new_n14972_), .ZN(new_n15165_));
  NOR2_X1    g15070(.A1(new_n14950_), .A2(new_n14954_), .ZN(new_n15166_));
  NAND2_X1   g15071(.A1(new_n10652_), .A2(new_n962_), .ZN(new_n15167_));
  AOI22_X1   g15072(.A1(new_n10805_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n10817_), .ZN(new_n15168_));
  AOI21_X1   g15073(.A1(new_n15167_), .A2(new_n15168_), .B(new_n82_), .ZN(new_n15169_));
  OAI21_X1   g15074(.A1(new_n11218_), .A2(new_n11223_), .B(new_n15169_), .ZN(new_n15170_));
  XOR2_X1    g15075(.A1(new_n15166_), .A2(new_n15170_), .Z(new_n15171_));
  INV_X1     g15076(.I(new_n15171_), .ZN(new_n15172_));
  OAI22_X1   g15077(.A1(new_n11264_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10646_), .ZN(new_n15173_));
  OAI21_X1   g15078(.A1(new_n79_), .A2(new_n10633_), .B(new_n15173_), .ZN(new_n15174_));
  AOI21_X1   g15079(.A1(new_n15174_), .A2(new_n72_), .B(new_n79_), .ZN(new_n15175_));
  XOR2_X1    g15080(.A1(new_n11987_), .A2(new_n15175_), .Z(new_n15176_));
  XOR2_X1    g15081(.A1(new_n15176_), .A2(new_n15172_), .Z(new_n15177_));
  NAND3_X1   g15082(.A1(new_n15177_), .A2(new_n14961_), .A3(new_n14964_), .ZN(new_n15178_));
  NAND2_X1   g15083(.A1(new_n14960_), .A2(new_n14956_), .ZN(new_n15180_));
  NAND2_X1   g15084(.A1(new_n15178_), .A2(new_n15180_), .ZN(new_n15181_));
  NAND2_X1   g15085(.A1(new_n15181_), .A2(new_n14948_), .ZN(new_n15182_));
  NOR2_X1    g15086(.A1(new_n15181_), .A2(new_n14948_), .ZN(new_n15183_));
  INV_X1     g15087(.I(new_n15183_), .ZN(new_n15184_));
  OAI22_X1   g15088(.A1(new_n10844_), .A2(new_n4781_), .B1(new_n10631_), .B2(new_n4612_), .ZN(new_n15185_));
  OAI21_X1   g15089(.A1(new_n1128_), .A2(new_n10856_), .B(new_n15185_), .ZN(new_n15186_));
  AOI21_X1   g15090(.A1(new_n15186_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n15187_));
  XOR2_X1    g15091(.A1(new_n11631_), .A2(new_n15187_), .Z(new_n15188_));
  INV_X1     g15092(.I(new_n15188_), .ZN(new_n15189_));
  NAND3_X1   g15093(.A1(new_n15184_), .A2(new_n15182_), .A3(new_n15189_), .ZN(new_n15190_));
  INV_X1     g15094(.I(new_n15182_), .ZN(new_n15191_));
  OAI21_X1   g15095(.A1(new_n15191_), .A2(new_n15183_), .B(new_n15188_), .ZN(new_n15192_));
  NAND2_X1   g15096(.A1(new_n15192_), .A2(new_n15190_), .ZN(new_n15193_));
  INV_X1     g15097(.I(new_n15193_), .ZN(new_n15194_));
  NAND3_X1   g15098(.A1(new_n15194_), .A2(new_n15165_), .A3(new_n15164_), .ZN(new_n15195_));
  INV_X1     g15099(.I(new_n15165_), .ZN(new_n15196_));
  OAI21_X1   g15100(.A1(new_n15196_), .A2(new_n14974_), .B(new_n15193_), .ZN(new_n15197_));
  AOI22_X1   g15101(.A1(new_n13242_), .A2(new_n5783_), .B1(new_n247_), .B2(new_n10882_), .ZN(new_n15198_));
  OAI21_X1   g15102(.A1(new_n15198_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n15199_));
  NOR2_X1    g15103(.A1(new_n11802_), .A2(new_n15199_), .ZN(new_n15200_));
  AND2_X2    g15104(.A1(new_n11802_), .A2(new_n15199_), .Z(new_n15201_));
  NOR2_X1    g15105(.A1(new_n15201_), .A2(new_n15200_), .ZN(new_n15202_));
  NAND3_X1   g15106(.A1(new_n15195_), .A2(new_n15197_), .A3(new_n15202_), .ZN(new_n15203_));
  NOR3_X1    g15107(.A1(new_n15196_), .A2(new_n15193_), .A3(new_n14974_), .ZN(new_n15204_));
  AOI21_X1   g15108(.A1(new_n15164_), .A2(new_n15165_), .B(new_n15194_), .ZN(new_n15205_));
  INV_X1     g15109(.I(new_n15202_), .ZN(new_n15206_));
  OAI21_X1   g15110(.A1(new_n15205_), .A2(new_n15204_), .B(new_n15206_), .ZN(new_n15207_));
  NAND3_X1   g15111(.A1(new_n15207_), .A2(new_n15203_), .A3(new_n14985_), .ZN(new_n15208_));
  NAND3_X1   g15112(.A1(new_n15208_), .A2(new_n15161_), .A3(new_n15163_), .ZN(new_n15209_));
  NOR3_X1    g15113(.A1(new_n15205_), .A2(new_n15204_), .A3(new_n15206_), .ZN(new_n15210_));
  AOI21_X1   g15114(.A1(new_n15195_), .A2(new_n15197_), .B(new_n15202_), .ZN(new_n15211_));
  NOR3_X1    g15115(.A1(new_n15210_), .A2(new_n15211_), .A3(new_n14986_), .ZN(new_n15212_));
  OAI21_X1   g15116(.A1(new_n15212_), .A2(new_n14988_), .B(new_n14943_), .ZN(new_n15213_));
  AOI22_X1   g15117(.A1(new_n10986_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n10897_), .ZN(new_n15214_));
  OAI21_X1   g15118(.A1(new_n15214_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n15215_));
  NOR2_X1    g15119(.A1(new_n10984_), .A2(new_n15215_), .ZN(new_n15216_));
  INV_X1     g15120(.I(new_n15215_), .ZN(new_n15217_));
  NOR2_X1    g15121(.A1(new_n13293_), .A2(new_n15217_), .ZN(new_n15218_));
  NOR2_X1    g15122(.A1(new_n15218_), .A2(new_n15216_), .ZN(new_n15219_));
  INV_X1     g15123(.I(new_n15219_), .ZN(new_n15220_));
  NAND3_X1   g15124(.A1(new_n15213_), .A2(new_n15209_), .A3(new_n15220_), .ZN(new_n15221_));
  NOR3_X1    g15125(.A1(new_n15212_), .A2(new_n14943_), .A3(new_n14988_), .ZN(new_n15222_));
  AOI21_X1   g15126(.A1(new_n15208_), .A2(new_n15163_), .B(new_n15161_), .ZN(new_n15223_));
  OAI21_X1   g15127(.A1(new_n15222_), .A2(new_n15223_), .B(new_n15219_), .ZN(new_n15224_));
  NAND3_X1   g15128(.A1(new_n15224_), .A2(new_n15221_), .A3(new_n15000_), .ZN(new_n15225_));
  NAND3_X1   g15129(.A1(new_n15225_), .A2(new_n14938_), .A3(new_n15001_), .ZN(new_n15226_));
  NOR3_X1    g15130(.A1(new_n15222_), .A2(new_n15223_), .A3(new_n15219_), .ZN(new_n15227_));
  AOI21_X1   g15131(.A1(new_n15213_), .A2(new_n15209_), .B(new_n15220_), .ZN(new_n15228_));
  NOR3_X1    g15132(.A1(new_n15227_), .A2(new_n15228_), .A3(new_n15004_), .ZN(new_n15229_));
  OAI21_X1   g15133(.A1(new_n15229_), .A2(new_n15005_), .B(new_n14939_), .ZN(new_n15230_));
  OAI22_X1   g15134(.A1(new_n12601_), .A2(new_n5420_), .B1(new_n1620_), .B2(new_n10595_), .ZN(new_n15231_));
  AOI21_X1   g15135(.A1(new_n15231_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n15232_));
  XOR2_X1    g15136(.A1(new_n12600_), .A2(new_n15232_), .Z(new_n15233_));
  NAND3_X1   g15137(.A1(new_n15230_), .A2(new_n15226_), .A3(new_n15233_), .ZN(new_n15234_));
  NOR3_X1    g15138(.A1(new_n15229_), .A2(new_n14939_), .A3(new_n15005_), .ZN(new_n15235_));
  AOI21_X1   g15139(.A1(new_n15225_), .A2(new_n15001_), .B(new_n14938_), .ZN(new_n15236_));
  XOR2_X1    g15140(.A1(new_n13949_), .A2(new_n15232_), .Z(new_n15237_));
  OAI21_X1   g15141(.A1(new_n15235_), .A2(new_n15236_), .B(new_n15237_), .ZN(new_n15238_));
  NAND3_X1   g15142(.A1(new_n15234_), .A2(new_n15238_), .A3(new_n15021_), .ZN(new_n15239_));
  NAND3_X1   g15143(.A1(new_n15239_), .A2(new_n15019_), .A3(new_n15015_), .ZN(new_n15240_));
  NOR3_X1    g15144(.A1(new_n15235_), .A2(new_n15236_), .A3(new_n15237_), .ZN(new_n15241_));
  AOI21_X1   g15145(.A1(new_n15230_), .A2(new_n15226_), .B(new_n15233_), .ZN(new_n15242_));
  NOR3_X1    g15146(.A1(new_n15242_), .A2(new_n15241_), .A3(new_n15011_), .ZN(new_n15243_));
  OAI21_X1   g15147(.A1(new_n15026_), .A2(new_n15243_), .B(new_n15023_), .ZN(new_n15244_));
  AOI22_X1   g15148(.A1(new_n12891_), .A2(new_n5968_), .B1(new_n10924_), .B2(new_n785_), .ZN(new_n15245_));
  OAI21_X1   g15149(.A1(new_n15245_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n15246_));
  XOR2_X1    g15150(.A1(new_n12889_), .A2(new_n15246_), .Z(new_n15247_));
  NAND3_X1   g15151(.A1(new_n15244_), .A2(new_n15240_), .A3(new_n15247_), .ZN(new_n15248_));
  NOR3_X1    g15152(.A1(new_n15026_), .A2(new_n15243_), .A3(new_n15023_), .ZN(new_n15249_));
  AOI21_X1   g15153(.A1(new_n15239_), .A2(new_n15019_), .B(new_n15015_), .ZN(new_n15250_));
  XNOR2_X1   g15154(.A1(new_n12889_), .A2(new_n15246_), .ZN(new_n15251_));
  OAI21_X1   g15155(.A1(new_n15249_), .A2(new_n15250_), .B(new_n15251_), .ZN(new_n15252_));
  NAND3_X1   g15156(.A1(new_n15252_), .A2(new_n15248_), .A3(new_n15035_), .ZN(new_n15253_));
  NAND3_X1   g15157(.A1(new_n15040_), .A2(new_n15253_), .A3(new_n15036_), .ZN(new_n15254_));
  NOR3_X1    g15158(.A1(new_n15249_), .A2(new_n15251_), .A3(new_n15250_), .ZN(new_n15255_));
  AOI21_X1   g15159(.A1(new_n15244_), .A2(new_n15240_), .B(new_n15247_), .ZN(new_n15256_));
  NOR3_X1    g15160(.A1(new_n15255_), .A2(new_n15256_), .A3(new_n15042_), .ZN(new_n15257_));
  OAI21_X1   g15161(.A1(new_n15257_), .A2(new_n15043_), .B(new_n14934_), .ZN(new_n15258_));
  AOI22_X1   g15162(.A1(new_n12909_), .A2(new_n6758_), .B1(new_n10949_), .B2(new_n805_), .ZN(new_n15259_));
  OAI21_X1   g15163(.A1(new_n15259_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n15260_));
  XOR2_X1    g15164(.A1(new_n12907_), .A2(new_n15260_), .Z(new_n15261_));
  NAND3_X1   g15165(.A1(new_n15258_), .A2(new_n15254_), .A3(new_n15261_), .ZN(new_n15262_));
  NOR3_X1    g15166(.A1(new_n15257_), .A2(new_n14934_), .A3(new_n15043_), .ZN(new_n15263_));
  AOI22_X1   g15167(.A1(new_n15253_), .A2(new_n15036_), .B1(new_n14931_), .B2(new_n14933_), .ZN(new_n15264_));
  XNOR2_X1   g15168(.A1(new_n12907_), .A2(new_n15260_), .ZN(new_n15265_));
  OAI21_X1   g15169(.A1(new_n15264_), .A2(new_n15263_), .B(new_n15265_), .ZN(new_n15266_));
  NAND3_X1   g15170(.A1(new_n15262_), .A2(new_n15266_), .A3(new_n15064_), .ZN(new_n15267_));
  NAND3_X1   g15171(.A1(new_n15267_), .A2(new_n15062_), .A3(new_n15057_), .ZN(new_n15268_));
  INV_X1     g15172(.I(new_n15268_), .ZN(new_n15269_));
  AOI21_X1   g15173(.A1(new_n15267_), .A2(new_n15062_), .B(new_n15057_), .ZN(new_n15270_));
  INV_X1     g15174(.I(new_n10965_), .ZN(new_n15271_));
  AOI22_X1   g15175(.A1(new_n15271_), .A2(new_n7838_), .B1(new_n10571_), .B2(new_n2469_), .ZN(new_n15272_));
  OAI21_X1   g15176(.A1(new_n15272_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n15273_));
  INV_X1     g15177(.I(new_n15273_), .ZN(new_n15274_));
  XOR2_X1    g15178(.A1(new_n14077_), .A2(new_n15274_), .Z(new_n15275_));
  INV_X1     g15179(.I(new_n15275_), .ZN(new_n15276_));
  NOR3_X1    g15180(.A1(new_n15269_), .A2(new_n15270_), .A3(new_n15276_), .ZN(new_n15277_));
  NAND2_X1   g15181(.A1(new_n15267_), .A2(new_n15062_), .ZN(new_n15278_));
  NAND2_X1   g15182(.A1(new_n15278_), .A2(new_n15066_), .ZN(new_n15279_));
  AOI21_X1   g15183(.A1(new_n15279_), .A2(new_n15268_), .B(new_n15275_), .ZN(new_n15280_));
  NOR3_X1    g15184(.A1(new_n15280_), .A2(new_n15277_), .A3(new_n15160_), .ZN(new_n15281_));
  NOR3_X1    g15185(.A1(new_n15281_), .A2(new_n15159_), .A3(new_n14929_), .ZN(new_n15282_));
  OAI21_X1   g15186(.A1(new_n15281_), .A2(new_n15159_), .B(new_n14929_), .ZN(new_n15283_));
  INV_X1     g15187(.I(new_n15283_), .ZN(new_n15284_));
  AOI22_X1   g15188(.A1(new_n14602_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n14603_), .ZN(new_n15285_));
  OAI21_X1   g15189(.A1(new_n15285_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n15286_));
  XNOR2_X1   g15190(.A1(new_n14601_), .A2(new_n15286_), .ZN(new_n15287_));
  INV_X1     g15191(.I(new_n15287_), .ZN(new_n15288_));
  NOR3_X1    g15192(.A1(new_n15284_), .A2(new_n15282_), .A3(new_n15288_), .ZN(new_n15289_));
  INV_X1     g15193(.I(new_n15282_), .ZN(new_n15290_));
  AOI21_X1   g15194(.A1(new_n15290_), .A2(new_n15283_), .B(new_n15287_), .ZN(new_n15291_));
  NOR3_X1    g15195(.A1(new_n15291_), .A2(new_n15289_), .A3(new_n15158_), .ZN(new_n15292_));
  NOR3_X1    g15196(.A1(new_n15292_), .A2(new_n15156_), .A3(new_n15157_), .ZN(new_n15293_));
  NAND3_X1   g15197(.A1(new_n15290_), .A2(new_n15283_), .A3(new_n15287_), .ZN(new_n15294_));
  OAI21_X1   g15198(.A1(new_n15284_), .A2(new_n15282_), .B(new_n15288_), .ZN(new_n15295_));
  NAND3_X1   g15199(.A1(new_n15295_), .A2(new_n15294_), .A3(new_n15091_), .ZN(new_n15296_));
  AOI21_X1   g15200(.A1(new_n15296_), .A2(new_n15095_), .B(new_n14925_), .ZN(new_n15297_));
  NOR2_X1    g15201(.A1(new_n15293_), .A2(new_n15297_), .ZN(new_n15298_));
  NAND2_X1   g15202(.A1(new_n15123_), .A2(new_n15114_), .ZN(new_n15299_));
  NAND2_X1   g15203(.A1(new_n15122_), .A2(new_n15299_), .ZN(new_n15300_));
  AOI21_X1   g15204(.A1(new_n14262_), .A2(new_n14878_), .B(new_n14876_), .ZN(new_n15301_));
  NOR2_X1    g15205(.A1(new_n15109_), .A2(new_n15301_), .ZN(new_n15302_));
  NAND2_X1   g15206(.A1(new_n15109_), .A2(new_n15301_), .ZN(new_n15303_));
  INV_X1     g15207(.I(new_n15303_), .ZN(new_n15304_));
  NOR2_X1    g15208(.A1(new_n15304_), .A2(new_n15302_), .ZN(new_n15305_));
  XNOR2_X1   g15209(.A1(new_n15305_), .A2(new_n15114_), .ZN(new_n15306_));
  INV_X1     g15210(.I(new_n15306_), .ZN(new_n15307_));
  NAND2_X1   g15211(.A1(new_n15300_), .A2(new_n15307_), .ZN(new_n15308_));
  INV_X1     g15212(.I(new_n15300_), .ZN(new_n15309_));
  XNOR2_X1   g15213(.A1(new_n15305_), .A2(new_n15114_), .ZN(new_n15310_));
  NAND2_X1   g15214(.A1(new_n15309_), .A2(new_n15310_), .ZN(new_n15311_));
  NAND2_X1   g15215(.A1(new_n15311_), .A2(new_n15308_), .ZN(new_n15312_));
  NOR2_X1    g15216(.A1(new_n14886_), .A2(new_n15114_), .ZN(new_n15313_));
  OAI22_X1   g15217(.A1(new_n15313_), .A2(new_n9425_), .B1(new_n3456_), .B2(new_n15305_), .ZN(new_n15314_));
  AOI21_X1   g15218(.A1(new_n15314_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n15315_));
  XNOR2_X1   g15219(.A1(new_n15312_), .A2(new_n15315_), .ZN(new_n15316_));
  NAND2_X1   g15220(.A1(new_n15298_), .A2(new_n15316_), .ZN(new_n15317_));
  NAND3_X1   g15221(.A1(new_n15296_), .A2(new_n14925_), .A3(new_n15095_), .ZN(new_n15318_));
  OAI21_X1   g15222(.A1(new_n15292_), .A2(new_n15157_), .B(new_n15156_), .ZN(new_n15319_));
  NAND2_X1   g15223(.A1(new_n15319_), .A2(new_n15318_), .ZN(new_n15320_));
  INV_X1     g15224(.I(new_n15316_), .ZN(new_n15321_));
  NAND2_X1   g15225(.A1(new_n15320_), .A2(new_n15321_), .ZN(new_n15322_));
  AOI21_X1   g15226(.A1(new_n15317_), .A2(new_n15322_), .B(new_n15152_), .ZN(new_n15323_));
  INV_X1     g15227(.I(new_n15323_), .ZN(new_n15324_));
  XOR2_X1    g15228(.A1(new_n15147_), .A2(new_n15324_), .Z(new_n15325_));
  XOR2_X1    g15229(.A1(new_n15325_), .A2(new_n15140_), .Z(\result[4] ));
  AOI21_X1   g15230(.A1(new_n15141_), .A2(new_n15145_), .B(new_n15324_), .ZN(new_n15327_));
  AND2_X2    g15231(.A1(new_n15094_), .A2(new_n15091_), .Z(new_n15329_));
  NOR3_X1    g15232(.A1(new_n15264_), .A2(new_n15263_), .A3(new_n15265_), .ZN(new_n15330_));
  AOI21_X1   g15233(.A1(new_n15262_), .A2(new_n15266_), .B(new_n15064_), .ZN(new_n15331_));
  OAI21_X1   g15234(.A1(new_n15331_), .A2(new_n15062_), .B(new_n15066_), .ZN(new_n15332_));
  OAI21_X1   g15235(.A1(new_n15242_), .A2(new_n15241_), .B(new_n15011_), .ZN(new_n15333_));
  AOI21_X1   g15236(.A1(new_n15026_), .A2(new_n15333_), .B(new_n15015_), .ZN(new_n15334_));
  AOI21_X1   g15237(.A1(new_n14998_), .A2(new_n15000_), .B(new_n14938_), .ZN(new_n15336_));
  NAND2_X1   g15238(.A1(new_n10828_), .A2(new_n962_), .ZN(new_n15337_));
  AOI22_X1   g15239(.A1(new_n10652_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n10805_), .ZN(new_n15338_));
  AOI21_X1   g15240(.A1(new_n15337_), .A2(new_n15338_), .B(new_n82_), .ZN(new_n15339_));
  NAND2_X1   g15241(.A1(new_n11246_), .A2(new_n15339_), .ZN(new_n15340_));
  NOR3_X1    g15242(.A1(new_n15170_), .A2(new_n14950_), .A3(new_n14954_), .ZN(new_n15341_));
  XOR2_X1    g15243(.A1(new_n15340_), .A2(new_n15341_), .Z(new_n15342_));
  OAI22_X1   g15244(.A1(new_n10633_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n11264_), .ZN(new_n15343_));
  OAI21_X1   g15245(.A1(new_n10631_), .A2(new_n79_), .B(new_n15343_), .ZN(new_n15344_));
  AOI21_X1   g15246(.A1(new_n15344_), .A2(new_n72_), .B(new_n79_), .ZN(new_n15345_));
  XOR2_X1    g15247(.A1(new_n11445_), .A2(new_n15345_), .Z(new_n15346_));
  XNOR2_X1   g15248(.A1(new_n15346_), .A2(new_n15342_), .ZN(new_n15347_));
  AOI21_X1   g15249(.A1(new_n15177_), .A2(new_n14960_), .B(new_n14956_), .ZN(new_n15348_));
  OAI21_X1   g15250(.A1(new_n15177_), .A2(new_n14960_), .B(new_n14949_), .ZN(new_n15349_));
  OAI22_X1   g15251(.A1(new_n15348_), .A2(new_n15349_), .B1(new_n15172_), .B2(new_n15176_), .ZN(new_n15350_));
  NOR2_X1    g15252(.A1(new_n15350_), .A2(new_n15347_), .ZN(new_n15351_));
  NAND2_X1   g15253(.A1(new_n15350_), .A2(new_n15347_), .ZN(new_n15352_));
  INV_X1     g15254(.I(new_n15352_), .ZN(new_n15353_));
  OAI22_X1   g15255(.A1(new_n10844_), .A2(new_n4612_), .B1(new_n4781_), .B2(new_n10856_), .ZN(new_n15354_));
  OAI21_X1   g15256(.A1(new_n10870_), .A2(new_n1128_), .B(new_n15354_), .ZN(new_n15355_));
  AOI21_X1   g15257(.A1(new_n15355_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n15356_));
  XOR2_X1    g15258(.A1(new_n11648_), .A2(new_n15356_), .Z(new_n15357_));
  NOR3_X1    g15259(.A1(new_n15353_), .A2(new_n15351_), .A3(new_n15357_), .ZN(new_n15358_));
  OAI21_X1   g15260(.A1(new_n15353_), .A2(new_n15351_), .B(new_n15357_), .ZN(new_n15359_));
  INV_X1     g15261(.I(new_n15359_), .ZN(new_n15360_));
  NOR2_X1    g15262(.A1(new_n15360_), .A2(new_n15358_), .ZN(new_n15361_));
  INV_X1     g15263(.I(new_n15361_), .ZN(new_n15362_));
  NAND3_X1   g15264(.A1(new_n15362_), .A2(new_n15195_), .A3(new_n15192_), .ZN(new_n15363_));
  NAND2_X1   g15265(.A1(new_n15195_), .A2(new_n15192_), .ZN(new_n15364_));
  NAND2_X1   g15266(.A1(new_n15364_), .A2(new_n15361_), .ZN(new_n15365_));
  OAI22_X1   g15267(.A1(new_n10619_), .A2(new_n1239_), .B1(new_n4981_), .B2(new_n10885_), .ZN(new_n15366_));
  AOI21_X1   g15268(.A1(new_n15366_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n15367_));
  AND2_X2    g15269(.A1(new_n12074_), .A2(new_n15367_), .Z(new_n15368_));
  NOR2_X1    g15270(.A1(new_n12074_), .A2(new_n15367_), .ZN(new_n15369_));
  NOR2_X1    g15271(.A1(new_n15368_), .A2(new_n15369_), .ZN(new_n15370_));
  NAND3_X1   g15272(.A1(new_n15365_), .A2(new_n15363_), .A3(new_n15370_), .ZN(new_n15371_));
  INV_X1     g15273(.I(new_n15363_), .ZN(new_n15372_));
  AOI21_X1   g15274(.A1(new_n15192_), .A2(new_n15195_), .B(new_n15362_), .ZN(new_n15373_));
  INV_X1     g15275(.I(new_n15370_), .ZN(new_n15374_));
  OAI21_X1   g15276(.A1(new_n15372_), .A2(new_n15373_), .B(new_n15374_), .ZN(new_n15375_));
  NAND2_X1   g15277(.A1(new_n15375_), .A2(new_n15371_), .ZN(new_n15376_));
  OAI21_X1   g15278(.A1(new_n14986_), .A2(new_n14987_), .B(new_n14943_), .ZN(new_n15378_));
  NAND2_X1   g15279(.A1(new_n15378_), .A2(new_n15203_), .ZN(new_n15379_));
  NAND2_X1   g15280(.A1(new_n15376_), .A2(new_n15379_), .ZN(new_n15380_));
  NAND4_X1   g15281(.A1(new_n15375_), .A2(new_n15371_), .A3(new_n15378_), .A4(new_n15203_), .ZN(new_n15381_));
  OAI22_X1   g15282(.A1(new_n10606_), .A2(new_n5398_), .B1(new_n5336_), .B2(new_n10901_), .ZN(new_n15382_));
  AOI21_X1   g15283(.A1(new_n15382_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n15383_));
  AND2_X2    g15284(.A1(new_n12211_), .A2(new_n15383_), .Z(new_n15384_));
  NOR2_X1    g15285(.A1(new_n12211_), .A2(new_n15383_), .ZN(new_n15385_));
  NOR2_X1    g15286(.A1(new_n15384_), .A2(new_n15385_), .ZN(new_n15386_));
  INV_X1     g15287(.I(new_n15386_), .ZN(new_n15387_));
  NAND3_X1   g15288(.A1(new_n15380_), .A2(new_n15387_), .A3(new_n15381_), .ZN(new_n15388_));
  AOI22_X1   g15289(.A1(new_n15162_), .A2(new_n14985_), .B1(new_n14940_), .B2(new_n14942_), .ZN(new_n15389_));
  NOR2_X1    g15290(.A1(new_n15389_), .A2(new_n15210_), .ZN(new_n15390_));
  AOI21_X1   g15291(.A1(new_n15371_), .A2(new_n15375_), .B(new_n15390_), .ZN(new_n15391_));
  NOR3_X1    g15292(.A1(new_n15372_), .A2(new_n15373_), .A3(new_n15374_), .ZN(new_n15392_));
  AOI21_X1   g15293(.A1(new_n15365_), .A2(new_n15363_), .B(new_n15370_), .ZN(new_n15393_));
  NOR4_X1    g15294(.A1(new_n15392_), .A2(new_n15393_), .A3(new_n15210_), .A4(new_n15389_), .ZN(new_n15394_));
  OAI21_X1   g15295(.A1(new_n15391_), .A2(new_n15394_), .B(new_n15386_), .ZN(new_n15395_));
  NAND2_X1   g15296(.A1(new_n15388_), .A2(new_n15395_), .ZN(new_n15396_));
  NAND2_X1   g15297(.A1(new_n15396_), .A2(new_n15224_), .ZN(new_n15397_));
  NOR3_X1    g15298(.A1(new_n15391_), .A2(new_n15394_), .A3(new_n15386_), .ZN(new_n15398_));
  AOI21_X1   g15299(.A1(new_n15380_), .A2(new_n15381_), .B(new_n15387_), .ZN(new_n15399_));
  NOR2_X1    g15300(.A1(new_n15399_), .A2(new_n15398_), .ZN(new_n15400_));
  OAI21_X1   g15301(.A1(new_n15336_), .A2(new_n15228_), .B(new_n15400_), .ZN(new_n15401_));
  OAI21_X1   g15302(.A1(new_n15336_), .A2(new_n15397_), .B(new_n15401_), .ZN(new_n15402_));
  OAI22_X1   g15303(.A1(new_n10589_), .A2(new_n1620_), .B1(new_n12623_), .B2(new_n5420_), .ZN(new_n15403_));
  AOI21_X1   g15304(.A1(new_n15403_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n15404_));
  INV_X1     g15305(.I(new_n15404_), .ZN(new_n15405_));
  NOR2_X1    g15306(.A1(new_n13972_), .A2(new_n15405_), .ZN(new_n15406_));
  NOR2_X1    g15307(.A1(new_n12622_), .A2(new_n15404_), .ZN(new_n15407_));
  NOR2_X1    g15308(.A1(new_n15407_), .A2(new_n15406_), .ZN(new_n15408_));
  INV_X1     g15309(.I(new_n15408_), .ZN(new_n15409_));
  NAND2_X1   g15310(.A1(new_n15402_), .A2(new_n15409_), .ZN(new_n15410_));
  NOR2_X1    g15311(.A1(new_n15334_), .A2(new_n15410_), .ZN(new_n15411_));
  AOI21_X1   g15312(.A1(new_n15234_), .A2(new_n15238_), .B(new_n15021_), .ZN(new_n15412_));
  OAI21_X1   g15313(.A1(new_n15412_), .A2(new_n15019_), .B(new_n15023_), .ZN(new_n15413_));
  NOR2_X1    g15314(.A1(new_n15397_), .A2(new_n15336_), .ZN(new_n15414_));
  NOR2_X1    g15315(.A1(new_n15336_), .A2(new_n15228_), .ZN(new_n15415_));
  NOR2_X1    g15316(.A1(new_n15415_), .A2(new_n15396_), .ZN(new_n15416_));
  NOR2_X1    g15317(.A1(new_n15414_), .A2(new_n15416_), .ZN(new_n15417_));
  NOR2_X1    g15318(.A1(new_n15417_), .A2(new_n15408_), .ZN(new_n15418_));
  NOR2_X1    g15319(.A1(new_n15413_), .A2(new_n15418_), .ZN(new_n15419_));
  OAI21_X1   g15320(.A1(new_n15411_), .A2(new_n15419_), .B(new_n15234_), .ZN(new_n15420_));
  NAND2_X1   g15321(.A1(new_n15413_), .A2(new_n15418_), .ZN(new_n15421_));
  NAND2_X1   g15322(.A1(new_n15334_), .A2(new_n15410_), .ZN(new_n15422_));
  NAND3_X1   g15323(.A1(new_n15422_), .A2(new_n15421_), .A3(new_n15241_), .ZN(new_n15423_));
  AOI22_X1   g15324(.A1(new_n10584_), .A2(new_n785_), .B1(new_n5968_), .B2(new_n12887_), .ZN(new_n15424_));
  OAI21_X1   g15325(.A1(new_n15424_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n15425_));
  NOR2_X1    g15326(.A1(new_n13378_), .A2(new_n15425_), .ZN(new_n15426_));
  AND2_X2    g15327(.A1(new_n13378_), .A2(new_n15425_), .Z(new_n15427_));
  NOR2_X1    g15328(.A1(new_n15427_), .A2(new_n15426_), .ZN(new_n15428_));
  INV_X1     g15329(.I(new_n15428_), .ZN(new_n15429_));
  NAND3_X1   g15330(.A1(new_n15420_), .A2(new_n15423_), .A3(new_n15429_), .ZN(new_n15430_));
  AOI21_X1   g15331(.A1(new_n15422_), .A2(new_n15421_), .B(new_n15241_), .ZN(new_n15431_));
  NOR3_X1    g15332(.A1(new_n15411_), .A2(new_n15419_), .A3(new_n15234_), .ZN(new_n15432_));
  OAI21_X1   g15333(.A1(new_n15432_), .A2(new_n15431_), .B(new_n15428_), .ZN(new_n15433_));
  NOR2_X1    g15334(.A1(new_n15041_), .A2(new_n15042_), .ZN(new_n15435_));
  OAI21_X1   g15335(.A1(new_n15040_), .A2(new_n15435_), .B(new_n15252_), .ZN(new_n15436_));
  AOI21_X1   g15336(.A1(new_n15430_), .A2(new_n15433_), .B(new_n15436_), .ZN(new_n15437_));
  NOR3_X1    g15337(.A1(new_n15432_), .A2(new_n15431_), .A3(new_n15428_), .ZN(new_n15438_));
  AOI21_X1   g15338(.A1(new_n15420_), .A2(new_n15423_), .B(new_n15429_), .ZN(new_n15439_));
  NAND2_X1   g15339(.A1(new_n15035_), .A2(new_n15032_), .ZN(new_n15440_));
  AOI21_X1   g15340(.A1(new_n14934_), .A2(new_n15440_), .B(new_n15256_), .ZN(new_n15441_));
  NOR3_X1    g15341(.A1(new_n15438_), .A2(new_n15441_), .A3(new_n15439_), .ZN(new_n15442_));
  NOR2_X1    g15342(.A1(new_n15437_), .A2(new_n15442_), .ZN(new_n15443_));
  INV_X1     g15343(.I(new_n13544_), .ZN(new_n15444_));
  AOI22_X1   g15344(.A1(new_n5247_), .A2(new_n10937_), .B1(new_n10949_), .B2(new_n5249_), .ZN(new_n15445_));
  AOI21_X1   g15345(.A1(new_n10958_), .A2(new_n805_), .B(new_n15445_), .ZN(new_n15446_));
  OAI21_X1   g15346(.A1(new_n15446_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n15447_));
  NOR2_X1    g15347(.A1(new_n15444_), .A2(new_n15447_), .ZN(new_n15448_));
  INV_X1     g15348(.I(new_n15447_), .ZN(new_n15449_));
  NOR2_X1    g15349(.A1(new_n13544_), .A2(new_n15449_), .ZN(new_n15450_));
  NOR2_X1    g15350(.A1(new_n15448_), .A2(new_n15450_), .ZN(new_n15451_));
  NOR2_X1    g15351(.A1(new_n15443_), .A2(new_n15451_), .ZN(new_n15452_));
  NAND2_X1   g15352(.A1(new_n15332_), .A2(new_n15452_), .ZN(new_n15453_));
  AOI21_X1   g15353(.A1(new_n15258_), .A2(new_n15254_), .B(new_n15261_), .ZN(new_n15454_));
  OAI21_X1   g15354(.A1(new_n15454_), .A2(new_n15330_), .B(new_n15053_), .ZN(new_n15455_));
  AOI21_X1   g15355(.A1(new_n15455_), .A2(new_n15069_), .B(new_n15057_), .ZN(new_n15456_));
  OAI21_X1   g15356(.A1(new_n15438_), .A2(new_n15439_), .B(new_n15441_), .ZN(new_n15457_));
  NAND3_X1   g15357(.A1(new_n15436_), .A2(new_n15433_), .A3(new_n15430_), .ZN(new_n15458_));
  NAND2_X1   g15358(.A1(new_n15457_), .A2(new_n15458_), .ZN(new_n15459_));
  INV_X1     g15359(.I(new_n15451_), .ZN(new_n15460_));
  NAND2_X1   g15360(.A1(new_n15459_), .A2(new_n15460_), .ZN(new_n15461_));
  NAND2_X1   g15361(.A1(new_n15456_), .A2(new_n15461_), .ZN(new_n15462_));
  AOI21_X1   g15362(.A1(new_n15453_), .A2(new_n15462_), .B(new_n15330_), .ZN(new_n15463_));
  NOR2_X1    g15363(.A1(new_n15456_), .A2(new_n15461_), .ZN(new_n15464_));
  NOR2_X1    g15364(.A1(new_n15332_), .A2(new_n15452_), .ZN(new_n15465_));
  NOR3_X1    g15365(.A1(new_n15465_), .A2(new_n15464_), .A3(new_n15262_), .ZN(new_n15466_));
  NOR2_X1    g15366(.A1(new_n10570_), .A2(new_n7836_), .ZN(new_n15467_));
  NOR2_X1    g15367(.A1(new_n10961_), .A2(new_n2718_), .ZN(new_n15468_));
  OAI22_X1   g15368(.A1(new_n10564_), .A2(new_n2495_), .B1(new_n15467_), .B2(new_n15468_), .ZN(new_n15469_));
  AOI21_X1   g15369(.A1(new_n15469_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n15470_));
  NAND2_X1   g15370(.A1(new_n10976_), .A2(new_n15470_), .ZN(new_n15471_));
  INV_X1     g15371(.I(new_n15471_), .ZN(new_n15472_));
  NOR2_X1    g15372(.A1(new_n10976_), .A2(new_n15470_), .ZN(new_n15473_));
  NOR2_X1    g15373(.A1(new_n15472_), .A2(new_n15473_), .ZN(new_n15474_));
  NOR3_X1    g15374(.A1(new_n15463_), .A2(new_n15466_), .A3(new_n15474_), .ZN(new_n15475_));
  OAI21_X1   g15375(.A1(new_n15465_), .A2(new_n15464_), .B(new_n15262_), .ZN(new_n15476_));
  NAND3_X1   g15376(.A1(new_n15453_), .A2(new_n15462_), .A3(new_n15330_), .ZN(new_n15477_));
  INV_X1     g15377(.I(new_n15473_), .ZN(new_n15478_));
  NAND2_X1   g15378(.A1(new_n15478_), .A2(new_n15471_), .ZN(new_n15479_));
  AOI21_X1   g15379(.A1(new_n15476_), .A2(new_n15477_), .B(new_n15479_), .ZN(new_n15480_));
  NAND2_X1   g15380(.A1(new_n15083_), .A2(new_n15080_), .ZN(new_n15481_));
  AOI21_X1   g15381(.A1(new_n14929_), .A2(new_n15481_), .B(new_n15280_), .ZN(new_n15482_));
  OAI21_X1   g15382(.A1(new_n15475_), .A2(new_n15480_), .B(new_n15482_), .ZN(new_n15483_));
  NAND3_X1   g15383(.A1(new_n15476_), .A2(new_n15477_), .A3(new_n15479_), .ZN(new_n15484_));
  OAI21_X1   g15384(.A1(new_n15463_), .A2(new_n15466_), .B(new_n15474_), .ZN(new_n15485_));
  INV_X1     g15385(.I(new_n15482_), .ZN(new_n15486_));
  NAND3_X1   g15386(.A1(new_n15486_), .A2(new_n15484_), .A3(new_n15485_), .ZN(new_n15487_));
  OAI22_X1   g15387(.A1(new_n14276_), .A2(new_n3042_), .B1(new_n8830_), .B2(new_n14594_), .ZN(new_n15488_));
  OAI21_X1   g15388(.A1(new_n14886_), .A2(new_n3040_), .B(new_n15488_), .ZN(new_n15489_));
  AOI21_X1   g15389(.A1(new_n15489_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n15490_));
  XOR2_X1    g15390(.A1(new_n14891_), .A2(new_n15490_), .Z(new_n15491_));
  AOI21_X1   g15391(.A1(new_n15487_), .A2(new_n15483_), .B(new_n15491_), .ZN(new_n15492_));
  OAI21_X1   g15392(.A1(new_n15329_), .A2(new_n14925_), .B(new_n15492_), .ZN(new_n15493_));
  NAND2_X1   g15393(.A1(new_n15094_), .A2(new_n15091_), .ZN(new_n15494_));
  INV_X1     g15394(.I(new_n15492_), .ZN(new_n15495_));
  NAND3_X1   g15395(.A1(new_n15495_), .A2(new_n15156_), .A3(new_n15494_), .ZN(new_n15496_));
  AOI21_X1   g15396(.A1(new_n15496_), .A2(new_n15493_), .B(new_n15289_), .ZN(new_n15497_));
  AOI22_X1   g15397(.A1(new_n15155_), .A2(new_n15153_), .B1(new_n15091_), .B2(new_n15094_), .ZN(new_n15498_));
  NOR2_X1    g15398(.A1(new_n15498_), .A2(new_n15495_), .ZN(new_n15499_));
  NOR3_X1    g15399(.A1(new_n15329_), .A2(new_n14925_), .A3(new_n15492_), .ZN(new_n15500_));
  NOR3_X1    g15400(.A1(new_n15499_), .A2(new_n15294_), .A3(new_n15500_), .ZN(new_n15501_));
  INV_X1     g15401(.I(new_n15112_), .ZN(new_n15502_));
  INV_X1     g15402(.I(new_n14881_), .ZN(new_n15503_));
  AOI21_X1   g15403(.A1(new_n15099_), .A2(new_n15503_), .B(new_n15110_), .ZN(new_n15504_));
  AOI21_X1   g15404(.A1(new_n84_), .A2(new_n83_), .B(new_n72_), .ZN(new_n15505_));
  NOR2_X1    g15405(.A1(new_n15103_), .A2(new_n15505_), .ZN(new_n15506_));
  INV_X1     g15406(.I(new_n15506_), .ZN(new_n15507_));
  NOR3_X1    g15407(.A1(new_n15504_), .A2(new_n15502_), .A3(new_n15507_), .ZN(new_n15508_));
  OAI21_X1   g15408(.A1(new_n15504_), .A2(new_n15502_), .B(new_n15507_), .ZN(new_n15509_));
  INV_X1     g15409(.I(new_n15509_), .ZN(new_n15510_));
  NOR2_X1    g15410(.A1(new_n15510_), .A2(new_n15508_), .ZN(new_n15511_));
  NOR2_X1    g15411(.A1(new_n15115_), .A2(new_n15511_), .ZN(new_n15512_));
  OAI21_X1   g15412(.A1(new_n15100_), .A2(new_n14881_), .B(new_n15111_), .ZN(new_n15513_));
  NAND3_X1   g15413(.A1(new_n15513_), .A2(new_n15112_), .A3(new_n15506_), .ZN(new_n15514_));
  NAND2_X1   g15414(.A1(new_n15514_), .A2(new_n15509_), .ZN(new_n15515_));
  NOR2_X1    g15415(.A1(new_n15114_), .A2(new_n15515_), .ZN(new_n15516_));
  OAI21_X1   g15416(.A1(new_n15512_), .A2(new_n15516_), .B(new_n15307_), .ZN(new_n15517_));
  XOR2_X1    g15417(.A1(new_n15300_), .A2(new_n15517_), .Z(new_n15518_));
  OAI22_X1   g15418(.A1(new_n15305_), .A2(new_n9405_), .B1(new_n15114_), .B2(new_n9408_), .ZN(new_n15519_));
  OAI21_X1   g15419(.A1(new_n3456_), .A2(new_n15515_), .B(new_n15519_), .ZN(new_n15520_));
  AOI21_X1   g15420(.A1(new_n15520_), .A2(new_n451_), .B(new_n3414_), .ZN(new_n15521_));
  XOR2_X1    g15421(.A1(new_n15518_), .A2(new_n15521_), .Z(new_n15522_));
  INV_X1     g15422(.I(new_n15522_), .ZN(new_n15523_));
  NOR3_X1    g15423(.A1(new_n15501_), .A2(new_n15497_), .A3(new_n15523_), .ZN(new_n15524_));
  OAI21_X1   g15424(.A1(new_n15499_), .A2(new_n15500_), .B(new_n15294_), .ZN(new_n15525_));
  NAND3_X1   g15425(.A1(new_n15496_), .A2(new_n15493_), .A3(new_n15289_), .ZN(new_n15526_));
  AOI21_X1   g15426(.A1(new_n15525_), .A2(new_n15526_), .B(new_n15522_), .ZN(new_n15527_));
  NOR2_X1    g15427(.A1(new_n15298_), .A2(new_n15321_), .ZN(new_n15528_));
  NOR2_X1    g15428(.A1(new_n15320_), .A2(new_n15316_), .ZN(new_n15529_));
  OAI22_X1   g15429(.A1(new_n15524_), .A2(new_n15527_), .B1(new_n15528_), .B2(new_n15529_), .ZN(new_n15530_));
  XNOR2_X1   g15430(.A1(new_n15530_), .A2(new_n15322_), .ZN(new_n15531_));
  XOR2_X1    g15431(.A1(new_n15531_), .A2(new_n15152_), .Z(new_n15532_));
  XOR2_X1    g15432(.A1(new_n15327_), .A2(new_n15532_), .Z(\result[5] ));
  AOI21_X1   g15433(.A1(new_n14620_), .A2(new_n14907_), .B(new_n15144_), .ZN(new_n15534_));
  NOR3_X1    g15434(.A1(new_n14913_), .A2(new_n15140_), .A3(new_n14914_), .ZN(new_n15535_));
  OAI21_X1   g15435(.A1(new_n15534_), .A2(new_n15535_), .B(new_n15323_), .ZN(new_n15536_));
  INV_X1     g15436(.I(new_n15150_), .ZN(new_n15537_));
  NAND3_X1   g15437(.A1(new_n14429_), .A2(new_n14921_), .A3(new_n15151_), .ZN(new_n15538_));
  NAND2_X1   g15438(.A1(new_n15538_), .A2(new_n15537_), .ZN(new_n15539_));
  XOR2_X1    g15439(.A1(new_n15531_), .A2(new_n15539_), .Z(new_n15540_));
  AOI21_X1   g15440(.A1(new_n15525_), .A2(new_n15526_), .B(new_n15523_), .ZN(new_n15541_));
  INV_X1     g15441(.I(new_n15541_), .ZN(new_n15542_));
  NOR3_X1    g15442(.A1(new_n15524_), .A2(new_n15527_), .A3(new_n15320_), .ZN(new_n15543_));
  OAI21_X1   g15443(.A1(new_n15524_), .A2(new_n15527_), .B(new_n15320_), .ZN(new_n15544_));
  AOI21_X1   g15444(.A1(new_n15316_), .A2(new_n15544_), .B(new_n15543_), .ZN(new_n15545_));
  INV_X1     g15445(.I(new_n15498_), .ZN(new_n15546_));
  NAND2_X1   g15446(.A1(new_n15487_), .A2(new_n15483_), .ZN(new_n15547_));
  NAND2_X1   g15447(.A1(new_n15289_), .A2(new_n15547_), .ZN(new_n15548_));
  INV_X1     g15448(.I(new_n15491_), .ZN(new_n15549_));
  OAI21_X1   g15449(.A1(new_n15289_), .A2(new_n15547_), .B(new_n15549_), .ZN(new_n15550_));
  OAI21_X1   g15450(.A1(new_n15546_), .A2(new_n15550_), .B(new_n15548_), .ZN(new_n15551_));
  NAND2_X1   g15451(.A1(new_n15459_), .A2(new_n15330_), .ZN(new_n15552_));
  AOI21_X1   g15452(.A1(new_n15443_), .A2(new_n15262_), .B(new_n15451_), .ZN(new_n15553_));
  NAND2_X1   g15453(.A1(new_n15456_), .A2(new_n15553_), .ZN(new_n15554_));
  AOI21_X1   g15454(.A1(new_n15417_), .A2(new_n15234_), .B(new_n15408_), .ZN(new_n15555_));
  AOI22_X1   g15455(.A1(new_n15334_), .A2(new_n15555_), .B1(new_n15241_), .B2(new_n15402_), .ZN(new_n15556_));
  NAND3_X1   g15456(.A1(new_n15379_), .A2(new_n15371_), .A3(new_n15375_), .ZN(new_n15557_));
  NAND2_X1   g15457(.A1(new_n15346_), .A2(new_n15342_), .ZN(new_n15558_));
  INV_X1     g15458(.I(new_n15558_), .ZN(new_n15559_));
  INV_X1     g15459(.I(new_n15350_), .ZN(new_n15560_));
  NOR2_X1    g15460(.A1(new_n15560_), .A2(new_n15347_), .ZN(new_n15561_));
  NAND3_X1   g15461(.A1(new_n11246_), .A2(new_n15339_), .A3(new_n15341_), .ZN(new_n15562_));
  INV_X1     g15462(.I(new_n15562_), .ZN(new_n15563_));
  OAI22_X1   g15463(.A1(new_n10631_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10633_), .ZN(new_n15564_));
  OAI21_X1   g15464(.A1(new_n10844_), .A2(new_n79_), .B(new_n15564_), .ZN(new_n15565_));
  AOI21_X1   g15465(.A1(new_n15565_), .A2(new_n72_), .B(new_n79_), .ZN(new_n15566_));
  XNOR2_X1   g15466(.A1(new_n11607_), .A2(new_n15566_), .ZN(new_n15567_));
  NOR3_X1    g15467(.A1(new_n15561_), .A2(new_n15563_), .A3(new_n15567_), .ZN(new_n15568_));
  NOR2_X1    g15468(.A1(new_n15567_), .A2(new_n15563_), .ZN(new_n15569_));
  NOR3_X1    g15469(.A1(new_n15560_), .A2(new_n15347_), .A3(new_n15569_), .ZN(new_n15570_));
  NOR2_X1    g15470(.A1(new_n15568_), .A2(new_n15570_), .ZN(new_n15571_));
  NOR2_X1    g15471(.A1(new_n15571_), .A2(new_n15559_), .ZN(new_n15572_));
  NAND2_X1   g15472(.A1(new_n15571_), .A2(new_n15559_), .ZN(new_n15573_));
  INV_X1     g15473(.I(new_n15573_), .ZN(new_n15574_));
  AOI22_X1   g15474(.A1(new_n10625_), .A2(new_n4767_), .B1(new_n4613_), .B2(new_n10857_), .ZN(new_n15575_));
  AOI21_X1   g15475(.A1(new_n117_), .A2(new_n10875_), .B(new_n15575_), .ZN(new_n15576_));
  OAI21_X1   g15476(.A1(new_n15576_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n15577_));
  XNOR2_X1   g15477(.A1(new_n11722_), .A2(new_n15577_), .ZN(new_n15578_));
  INV_X1     g15478(.I(new_n15578_), .ZN(new_n15579_));
  OAI21_X1   g15479(.A1(new_n15574_), .A2(new_n15572_), .B(new_n15579_), .ZN(new_n15580_));
  NOR2_X1    g15480(.A1(new_n15373_), .A2(new_n15580_), .ZN(new_n15581_));
  INV_X1     g15481(.I(new_n15572_), .ZN(new_n15582_));
  AOI21_X1   g15482(.A1(new_n15582_), .A2(new_n15573_), .B(new_n15578_), .ZN(new_n15583_));
  NOR2_X1    g15483(.A1(new_n15365_), .A2(new_n15583_), .ZN(new_n15584_));
  OAI21_X1   g15484(.A1(new_n15584_), .A2(new_n15581_), .B(new_n15359_), .ZN(new_n15585_));
  NAND2_X1   g15485(.A1(new_n15365_), .A2(new_n15583_), .ZN(new_n15586_));
  NAND2_X1   g15486(.A1(new_n15373_), .A2(new_n15580_), .ZN(new_n15587_));
  NAND3_X1   g15487(.A1(new_n15586_), .A2(new_n15587_), .A3(new_n15360_), .ZN(new_n15588_));
  OAI22_X1   g15488(.A1(new_n12091_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n10611_), .ZN(new_n15589_));
  AOI21_X1   g15489(.A1(new_n15589_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n15590_));
  XOR2_X1    g15490(.A1(new_n12090_), .A2(new_n15590_), .Z(new_n15591_));
  AOI21_X1   g15491(.A1(new_n15585_), .A2(new_n15588_), .B(new_n15591_), .ZN(new_n15592_));
  NAND2_X1   g15492(.A1(new_n15592_), .A2(new_n15557_), .ZN(new_n15593_));
  NOR2_X1    g15493(.A1(new_n15376_), .A2(new_n15390_), .ZN(new_n15594_));
  AOI21_X1   g15494(.A1(new_n15586_), .A2(new_n15587_), .B(new_n15360_), .ZN(new_n15595_));
  NOR3_X1    g15495(.A1(new_n15584_), .A2(new_n15581_), .A3(new_n15359_), .ZN(new_n15596_));
  INV_X1     g15496(.I(new_n15591_), .ZN(new_n15597_));
  OAI21_X1   g15497(.A1(new_n15596_), .A2(new_n15595_), .B(new_n15597_), .ZN(new_n15598_));
  NAND2_X1   g15498(.A1(new_n15598_), .A2(new_n15594_), .ZN(new_n15599_));
  AOI21_X1   g15499(.A1(new_n15599_), .A2(new_n15593_), .B(new_n15392_), .ZN(new_n15600_));
  NOR2_X1    g15500(.A1(new_n15598_), .A2(new_n15594_), .ZN(new_n15601_));
  NOR2_X1    g15501(.A1(new_n15592_), .A2(new_n15557_), .ZN(new_n15602_));
  NOR3_X1    g15502(.A1(new_n15601_), .A2(new_n15602_), .A3(new_n15371_), .ZN(new_n15603_));
  AOI22_X1   g15503(.A1(new_n12578_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n10600_), .ZN(new_n15604_));
  OAI21_X1   g15504(.A1(new_n15604_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n15605_));
  NOR2_X1    g15505(.A1(new_n14188_), .A2(new_n15605_), .ZN(new_n15606_));
  INV_X1     g15506(.I(new_n15605_), .ZN(new_n15607_));
  NOR2_X1    g15507(.A1(new_n12576_), .A2(new_n15607_), .ZN(new_n15608_));
  OAI22_X1   g15508(.A1(new_n15600_), .A2(new_n15603_), .B1(new_n15606_), .B2(new_n15608_), .ZN(new_n15609_));
  NOR2_X1    g15509(.A1(new_n15609_), .A2(new_n15416_), .ZN(new_n15610_));
  OAI21_X1   g15510(.A1(new_n15601_), .A2(new_n15602_), .B(new_n15371_), .ZN(new_n15611_));
  NAND3_X1   g15511(.A1(new_n15599_), .A2(new_n15593_), .A3(new_n15392_), .ZN(new_n15612_));
  NOR2_X1    g15512(.A1(new_n15606_), .A2(new_n15608_), .ZN(new_n15613_));
  AOI21_X1   g15513(.A1(new_n15611_), .A2(new_n15612_), .B(new_n15613_), .ZN(new_n15614_));
  NOR2_X1    g15514(.A1(new_n15614_), .A2(new_n15401_), .ZN(new_n15615_));
  OAI21_X1   g15515(.A1(new_n15610_), .A2(new_n15615_), .B(new_n15395_), .ZN(new_n15616_));
  NAND2_X1   g15516(.A1(new_n15614_), .A2(new_n15401_), .ZN(new_n15617_));
  NAND2_X1   g15517(.A1(new_n15609_), .A2(new_n15416_), .ZN(new_n15618_));
  NAND3_X1   g15518(.A1(new_n15618_), .A2(new_n15617_), .A3(new_n15399_), .ZN(new_n15619_));
  OAI22_X1   g15519(.A1(new_n10913_), .A2(new_n1620_), .B1(new_n12768_), .B2(new_n5420_), .ZN(new_n15620_));
  AOI21_X1   g15520(.A1(new_n15620_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n15621_));
  XOR2_X1    g15521(.A1(new_n12767_), .A2(new_n15621_), .Z(new_n15622_));
  NAND3_X1   g15522(.A1(new_n15616_), .A2(new_n15619_), .A3(new_n15622_), .ZN(new_n15623_));
  AOI21_X1   g15523(.A1(new_n15618_), .A2(new_n15617_), .B(new_n15399_), .ZN(new_n15624_));
  NOR3_X1    g15524(.A1(new_n15610_), .A2(new_n15615_), .A3(new_n15395_), .ZN(new_n15625_));
  INV_X1     g15525(.I(new_n15622_), .ZN(new_n15626_));
  OAI21_X1   g15526(.A1(new_n15625_), .A2(new_n15624_), .B(new_n15626_), .ZN(new_n15627_));
  AOI21_X1   g15527(.A1(new_n15623_), .A2(new_n15627_), .B(new_n15556_), .ZN(new_n15628_));
  OAI21_X1   g15528(.A1(new_n15402_), .A2(new_n15241_), .B(new_n15409_), .ZN(new_n15629_));
  OAI22_X1   g15529(.A1(new_n15629_), .A2(new_n15413_), .B1(new_n15234_), .B2(new_n15417_), .ZN(new_n15630_));
  OAI21_X1   g15530(.A1(new_n15625_), .A2(new_n15624_), .B(new_n15622_), .ZN(new_n15631_));
  NAND3_X1   g15531(.A1(new_n15616_), .A2(new_n15619_), .A3(new_n15626_), .ZN(new_n15632_));
  AOI21_X1   g15532(.A1(new_n15631_), .A2(new_n15632_), .B(new_n15630_), .ZN(new_n15633_));
  AOI22_X1   g15533(.A1(new_n15045_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n10937_), .ZN(new_n15634_));
  OAI21_X1   g15534(.A1(new_n15634_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n15635_));
  XNOR2_X1   g15535(.A1(new_n13394_), .A2(new_n15635_), .ZN(new_n15636_));
  INV_X1     g15536(.I(new_n15636_), .ZN(new_n15637_));
  OAI21_X1   g15537(.A1(new_n15628_), .A2(new_n15633_), .B(new_n15637_), .ZN(new_n15638_));
  NOR2_X1    g15538(.A1(new_n15442_), .A2(new_n15638_), .ZN(new_n15639_));
  NAND2_X1   g15539(.A1(new_n15627_), .A2(new_n15623_), .ZN(new_n15640_));
  NAND2_X1   g15540(.A1(new_n15640_), .A2(new_n15630_), .ZN(new_n15641_));
  NAND2_X1   g15541(.A1(new_n15631_), .A2(new_n15632_), .ZN(new_n15642_));
  NAND2_X1   g15542(.A1(new_n15642_), .A2(new_n15556_), .ZN(new_n15643_));
  AOI21_X1   g15543(.A1(new_n15643_), .A2(new_n15641_), .B(new_n15636_), .ZN(new_n15644_));
  NOR2_X1    g15544(.A1(new_n15458_), .A2(new_n15644_), .ZN(new_n15645_));
  OAI21_X1   g15545(.A1(new_n15645_), .A2(new_n15639_), .B(new_n15433_), .ZN(new_n15646_));
  NAND2_X1   g15546(.A1(new_n15458_), .A2(new_n15644_), .ZN(new_n15647_));
  NAND4_X1   g15547(.A1(new_n15638_), .A2(new_n15436_), .A3(new_n15430_), .A4(new_n15433_), .ZN(new_n15648_));
  NAND3_X1   g15548(.A1(new_n15647_), .A2(new_n15648_), .A3(new_n15439_), .ZN(new_n15649_));
  AOI22_X1   g15549(.A1(new_n15072_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n10962_), .ZN(new_n15650_));
  OAI21_X1   g15550(.A1(new_n15650_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n15651_));
  NOR2_X1    g15551(.A1(new_n15071_), .A2(new_n15651_), .ZN(new_n15652_));
  INV_X1     g15552(.I(new_n15651_), .ZN(new_n15653_));
  NOR2_X1    g15553(.A1(new_n14053_), .A2(new_n15653_), .ZN(new_n15654_));
  NOR2_X1    g15554(.A1(new_n15652_), .A2(new_n15654_), .ZN(new_n15655_));
  NAND3_X1   g15555(.A1(new_n15646_), .A2(new_n15649_), .A3(new_n15655_), .ZN(new_n15656_));
  AOI21_X1   g15556(.A1(new_n15647_), .A2(new_n15648_), .B(new_n15439_), .ZN(new_n15657_));
  NOR3_X1    g15557(.A1(new_n15645_), .A2(new_n15639_), .A3(new_n15433_), .ZN(new_n15658_));
  INV_X1     g15558(.I(new_n15655_), .ZN(new_n15659_));
  OAI21_X1   g15559(.A1(new_n15658_), .A2(new_n15657_), .B(new_n15659_), .ZN(new_n15660_));
  AOI22_X1   g15560(.A1(new_n15554_), .A2(new_n15552_), .B1(new_n15660_), .B2(new_n15656_), .ZN(new_n15661_));
  OAI21_X1   g15561(.A1(new_n15459_), .A2(new_n15330_), .B(new_n15460_), .ZN(new_n15662_));
  OAI21_X1   g15562(.A1(new_n15332_), .A2(new_n15662_), .B(new_n15552_), .ZN(new_n15663_));
  OAI21_X1   g15563(.A1(new_n15658_), .A2(new_n15657_), .B(new_n15655_), .ZN(new_n15664_));
  NAND3_X1   g15564(.A1(new_n15646_), .A2(new_n15649_), .A3(new_n15659_), .ZN(new_n15665_));
  AOI21_X1   g15565(.A1(new_n15664_), .A2(new_n15665_), .B(new_n15663_), .ZN(new_n15666_));
  NOR2_X1    g15566(.A1(new_n15666_), .A2(new_n15661_), .ZN(new_n15667_));
  INV_X1     g15567(.I(new_n15667_), .ZN(new_n15668_));
  AOI22_X1   g15568(.A1(new_n14281_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n14274_), .ZN(new_n15669_));
  OAI21_X1   g15569(.A1(new_n15669_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n15670_));
  XNOR2_X1   g15570(.A1(new_n14280_), .A2(new_n15670_), .ZN(new_n15671_));
  NAND2_X1   g15571(.A1(new_n15668_), .A2(new_n15671_), .ZN(new_n15672_));
  XOR2_X1    g15572(.A1(new_n15672_), .A2(new_n15487_), .Z(new_n15673_));
  XOR2_X1    g15573(.A1(new_n15673_), .A2(new_n15485_), .Z(new_n15674_));
  INV_X1     g15574(.I(new_n15305_), .ZN(new_n15675_));
  NOR3_X1    g15575(.A1(new_n15300_), .A2(new_n15675_), .A3(new_n15515_), .ZN(new_n15676_));
  NAND2_X1   g15576(.A1(new_n15675_), .A2(new_n15515_), .ZN(new_n15677_));
  OAI22_X1   g15577(.A1(new_n15676_), .A2(new_n15114_), .B1(new_n15309_), .B2(new_n15677_), .ZN(new_n15678_));
  NAND2_X1   g15578(.A1(new_n15515_), .A2(new_n9404_), .ZN(new_n15679_));
  NOR2_X1    g15579(.A1(new_n3455_), .A2(new_n9407_), .ZN(new_n15680_));
  AOI21_X1   g15580(.A1(new_n15675_), .A2(new_n15680_), .B(\a[2] ), .ZN(new_n15681_));
  AOI21_X1   g15581(.A1(new_n15681_), .A2(new_n15679_), .B(new_n3414_), .ZN(new_n15682_));
  XNOR2_X1   g15582(.A1(new_n15678_), .A2(new_n15682_), .ZN(new_n15683_));
  AOI22_X1   g15583(.A1(new_n15127_), .A2(new_n8832_), .B1(new_n2898_), .B2(new_n15115_), .ZN(new_n15684_));
  OAI21_X1   g15584(.A1(new_n15684_), .A2(\a[5] ), .B(new_n2898_), .ZN(new_n15685_));
  XOR2_X1    g15585(.A1(new_n15125_), .A2(new_n15685_), .Z(new_n15686_));
  XOR2_X1    g15586(.A1(new_n15683_), .A2(new_n15686_), .Z(new_n15687_));
  INV_X1     g15587(.I(new_n15686_), .ZN(new_n15688_));
  NAND2_X1   g15588(.A1(new_n15683_), .A2(new_n15688_), .ZN(new_n15689_));
  NOR2_X1    g15589(.A1(new_n15683_), .A2(new_n15688_), .ZN(new_n15690_));
  INV_X1     g15590(.I(new_n15690_), .ZN(new_n15691_));
  NAND2_X1   g15591(.A1(new_n15691_), .A2(new_n15689_), .ZN(new_n15692_));
  NAND2_X1   g15592(.A1(new_n15674_), .A2(new_n15692_), .ZN(new_n15693_));
  OAI21_X1   g15593(.A1(new_n15674_), .A2(new_n15687_), .B(new_n15693_), .ZN(new_n15694_));
  NAND2_X1   g15594(.A1(new_n15694_), .A2(new_n15551_), .ZN(new_n15695_));
  AOI21_X1   g15595(.A1(new_n15539_), .A2(new_n15545_), .B(new_n15695_), .ZN(new_n15696_));
  NAND3_X1   g15596(.A1(new_n15525_), .A2(new_n15526_), .A3(new_n15522_), .ZN(new_n15697_));
  OAI21_X1   g15597(.A1(new_n15501_), .A2(new_n15497_), .B(new_n15523_), .ZN(new_n15698_));
  NAND3_X1   g15598(.A1(new_n15698_), .A2(new_n15697_), .A3(new_n15298_), .ZN(new_n15699_));
  AOI21_X1   g15599(.A1(new_n15698_), .A2(new_n15697_), .B(new_n15298_), .ZN(new_n15700_));
  OAI21_X1   g15600(.A1(new_n15321_), .A2(new_n15700_), .B(new_n15699_), .ZN(new_n15701_));
  INV_X1     g15601(.I(new_n15551_), .ZN(new_n15702_));
  NOR2_X1    g15602(.A1(new_n15674_), .A2(new_n15687_), .ZN(new_n15703_));
  AOI21_X1   g15603(.A1(new_n15674_), .A2(new_n15692_), .B(new_n15703_), .ZN(new_n15704_));
  NOR2_X1    g15604(.A1(new_n15704_), .A2(new_n15702_), .ZN(new_n15705_));
  NOR3_X1    g15605(.A1(new_n15152_), .A2(new_n15705_), .A3(new_n15701_), .ZN(new_n15706_));
  OAI21_X1   g15606(.A1(new_n15696_), .A2(new_n15706_), .B(new_n15542_), .ZN(new_n15707_));
  OAI21_X1   g15607(.A1(new_n15152_), .A2(new_n15701_), .B(new_n15705_), .ZN(new_n15708_));
  NAND3_X1   g15608(.A1(new_n15539_), .A2(new_n15545_), .A3(new_n15695_), .ZN(new_n15709_));
  NAND3_X1   g15609(.A1(new_n15709_), .A2(new_n15708_), .A3(new_n15541_), .ZN(new_n15710_));
  NAND2_X1   g15610(.A1(new_n15707_), .A2(new_n15710_), .ZN(new_n15711_));
  OAI21_X1   g15611(.A1(new_n15536_), .A2(new_n15540_), .B(new_n15711_), .ZN(new_n15712_));
  AOI21_X1   g15612(.A1(new_n15709_), .A2(new_n15708_), .B(new_n15541_), .ZN(new_n15713_));
  NOR3_X1    g15613(.A1(new_n15696_), .A2(new_n15706_), .A3(new_n15542_), .ZN(new_n15714_));
  NOR2_X1    g15614(.A1(new_n15713_), .A2(new_n15714_), .ZN(new_n15715_));
  NAND4_X1   g15615(.A1(\result[3] ), .A2(new_n15323_), .A3(new_n15715_), .A4(new_n15532_), .ZN(new_n15716_));
  NAND2_X1   g15616(.A1(new_n15712_), .A2(new_n15716_), .ZN(\result[6] ));
  NAND2_X1   g15617(.A1(new_n15327_), .A2(new_n15532_), .ZN(new_n15718_));
  AOI22_X1   g15618(.A1(new_n14602_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n14603_), .ZN(new_n15719_));
  OAI21_X1   g15619(.A1(new_n15719_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n15720_));
  XNOR2_X1   g15620(.A1(new_n14601_), .A2(new_n15720_), .ZN(new_n15721_));
  NAND2_X1   g15621(.A1(new_n15668_), .A2(new_n15480_), .ZN(new_n15722_));
  NOR3_X1    g15622(.A1(new_n15475_), .A2(new_n15480_), .A3(new_n15482_), .ZN(new_n15723_));
  NAND2_X1   g15623(.A1(new_n15667_), .A2(new_n15485_), .ZN(new_n15724_));
  NAND3_X1   g15624(.A1(new_n15723_), .A2(new_n15724_), .A3(new_n15671_), .ZN(new_n15725_));
  NAND2_X1   g15625(.A1(new_n15725_), .A2(new_n15722_), .ZN(new_n15726_));
  OAI22_X1   g15626(.A1(new_n10965_), .A2(new_n6757_), .B1(new_n1078_), .B2(new_n10570_), .ZN(new_n15727_));
  AOI21_X1   g15627(.A1(new_n15727_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n15728_));
  XNOR2_X1   g15628(.A1(new_n14077_), .A2(new_n15728_), .ZN(new_n15729_));
  NAND2_X1   g15629(.A1(new_n15663_), .A2(new_n15664_), .ZN(new_n15730_));
  NAND2_X1   g15630(.A1(new_n15730_), .A2(new_n15665_), .ZN(new_n15731_));
  AOI22_X1   g15631(.A1(new_n12891_), .A2(new_n5421_), .B1(new_n10924_), .B2(new_n4660_), .ZN(new_n15732_));
  OAI21_X1   g15632(.A1(new_n15732_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n15733_));
  XNOR2_X1   g15633(.A1(new_n12889_), .A2(new_n15733_), .ZN(new_n15734_));
  INV_X1     g15634(.I(new_n15631_), .ZN(new_n15735_));
  OAI21_X1   g15635(.A1(new_n15735_), .A2(new_n15556_), .B(new_n15632_), .ZN(new_n15736_));
  OAI22_X1   g15636(.A1(new_n12601_), .A2(new_n5336_), .B1(new_n5398_), .B2(new_n10595_), .ZN(new_n15737_));
  AOI21_X1   g15637(.A1(new_n15737_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n15738_));
  XOR2_X1    g15638(.A1(new_n12600_), .A2(new_n15738_), .Z(new_n15739_));
  NAND2_X1   g15639(.A1(new_n15611_), .A2(new_n15612_), .ZN(new_n15740_));
  NOR2_X1    g15640(.A1(new_n15740_), .A2(new_n15399_), .ZN(new_n15741_));
  NOR2_X1    g15641(.A1(new_n15741_), .A2(new_n15613_), .ZN(new_n15742_));
  AOI22_X1   g15642(.A1(new_n15742_), .A2(new_n15416_), .B1(new_n15399_), .B2(new_n15740_), .ZN(new_n15743_));
  INV_X1     g15643(.I(new_n15743_), .ZN(new_n15744_));
  OAI22_X1   g15644(.A1(new_n10870_), .A2(new_n4612_), .B1(new_n4781_), .B2(new_n10868_), .ZN(new_n15745_));
  OAI21_X1   g15645(.A1(new_n1128_), .A2(new_n10881_), .B(new_n15745_), .ZN(new_n15746_));
  AOI21_X1   g15646(.A1(new_n15746_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n15747_));
  XNOR2_X1   g15647(.A1(new_n11802_), .A2(new_n15747_), .ZN(new_n15748_));
  OAI21_X1   g15648(.A1(new_n15574_), .A2(new_n15572_), .B(new_n15360_), .ZN(new_n15749_));
  NAND3_X1   g15649(.A1(new_n15582_), .A2(new_n15359_), .A3(new_n15573_), .ZN(new_n15750_));
  NAND3_X1   g15650(.A1(new_n15373_), .A2(new_n15750_), .A3(new_n15579_), .ZN(new_n15751_));
  NAND2_X1   g15651(.A1(new_n15751_), .A2(new_n15749_), .ZN(new_n15752_));
  NOR2_X1    g15652(.A1(new_n3416_), .A2(\a[2] ), .ZN(new_n15753_));
  INV_X1     g15653(.I(new_n15753_), .ZN(new_n15754_));
  NAND3_X1   g15654(.A1(new_n15511_), .A2(\a[2] ), .A3(new_n15754_), .ZN(new_n15755_));
  OAI21_X1   g15655(.A1(new_n15515_), .A2(new_n3415_), .B(new_n451_), .ZN(new_n15756_));
  NOR2_X1    g15656(.A1(new_n10633_), .A2(new_n511_), .ZN(new_n15757_));
  INV_X1     g15657(.I(new_n15757_), .ZN(new_n15758_));
  AOI22_X1   g15658(.A1(new_n10638_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n10828_), .ZN(new_n15759_));
  AOI21_X1   g15659(.A1(new_n15758_), .A2(new_n15759_), .B(new_n82_), .ZN(new_n15760_));
  NAND2_X1   g15660(.A1(new_n11987_), .A2(new_n15760_), .ZN(new_n15761_));
  INV_X1     g15661(.I(new_n15761_), .ZN(new_n15762_));
  AOI21_X1   g15662(.A1(new_n15755_), .A2(new_n15756_), .B(new_n15762_), .ZN(new_n15763_));
  NOR3_X1    g15663(.A1(new_n15515_), .A2(new_n451_), .A3(new_n15753_), .ZN(new_n15764_));
  AOI21_X1   g15664(.A1(new_n15511_), .A2(new_n15754_), .B(\a[2] ), .ZN(new_n15765_));
  NOR3_X1    g15665(.A1(new_n15765_), .A2(new_n15764_), .A3(new_n15761_), .ZN(new_n15766_));
  OAI22_X1   g15666(.A1(new_n10844_), .A2(new_n4527_), .B1(new_n10631_), .B2(new_n4529_), .ZN(new_n15767_));
  OAI21_X1   g15667(.A1(new_n79_), .A2(new_n10856_), .B(new_n15767_), .ZN(new_n15768_));
  AOI21_X1   g15668(.A1(new_n15768_), .A2(new_n72_), .B(new_n79_), .ZN(new_n15769_));
  XOR2_X1    g15669(.A1(new_n11631_), .A2(new_n15769_), .Z(new_n15770_));
  NAND2_X1   g15670(.A1(new_n10638_), .A2(new_n962_), .ZN(new_n15771_));
  AOI22_X1   g15671(.A1(new_n10828_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n10652_), .ZN(new_n15772_));
  AOI21_X1   g15672(.A1(new_n15771_), .A2(new_n15772_), .B(new_n82_), .ZN(new_n15773_));
  NAND3_X1   g15673(.A1(new_n11268_), .A2(new_n15340_), .A3(new_n15773_), .ZN(new_n15774_));
  INV_X1     g15674(.I(new_n15774_), .ZN(new_n15775_));
  XOR2_X1    g15675(.A1(new_n15770_), .A2(new_n15775_), .Z(new_n15776_));
  INV_X1     g15676(.I(new_n15776_), .ZN(new_n15777_));
  OAI21_X1   g15677(.A1(new_n15763_), .A2(new_n15766_), .B(new_n15777_), .ZN(new_n15778_));
  OAI21_X1   g15678(.A1(new_n15765_), .A2(new_n15764_), .B(new_n15761_), .ZN(new_n15779_));
  NAND3_X1   g15679(.A1(new_n15755_), .A2(new_n15756_), .A3(new_n15762_), .ZN(new_n15780_));
  AND2_X2    g15680(.A1(new_n15770_), .A2(new_n15774_), .Z(new_n15781_));
  NOR2_X1    g15681(.A1(new_n15770_), .A2(new_n15774_), .ZN(new_n15782_));
  NOR2_X1    g15682(.A1(new_n15781_), .A2(new_n15782_), .ZN(new_n15783_));
  INV_X1     g15683(.I(new_n15783_), .ZN(new_n15784_));
  NAND3_X1   g15684(.A1(new_n15779_), .A2(new_n15780_), .A3(new_n15784_), .ZN(new_n15785_));
  AOI21_X1   g15685(.A1(new_n15558_), .A2(new_n15563_), .B(new_n15567_), .ZN(new_n15786_));
  NAND2_X1   g15686(.A1(new_n15561_), .A2(new_n15786_), .ZN(new_n15787_));
  OAI21_X1   g15687(.A1(new_n15558_), .A2(new_n15563_), .B(new_n15787_), .ZN(new_n15788_));
  INV_X1     g15688(.I(new_n15788_), .ZN(new_n15789_));
  NAND3_X1   g15689(.A1(new_n15778_), .A2(new_n15785_), .A3(new_n15789_), .ZN(new_n15790_));
  AOI21_X1   g15690(.A1(new_n15779_), .A2(new_n15780_), .B(new_n15776_), .ZN(new_n15791_));
  NOR3_X1    g15691(.A1(new_n15763_), .A2(new_n15766_), .A3(new_n15783_), .ZN(new_n15792_));
  OAI21_X1   g15692(.A1(new_n15792_), .A2(new_n15791_), .B(new_n15788_), .ZN(new_n15793_));
  OAI22_X1   g15693(.A1(new_n10985_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n10896_), .ZN(new_n15794_));
  AOI21_X1   g15694(.A1(new_n15794_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n15795_));
  XNOR2_X1   g15695(.A1(new_n10984_), .A2(new_n15795_), .ZN(new_n15796_));
  INV_X1     g15696(.I(new_n15796_), .ZN(new_n15797_));
  NAND3_X1   g15697(.A1(new_n15793_), .A2(new_n15790_), .A3(new_n15797_), .ZN(new_n15798_));
  NOR3_X1    g15698(.A1(new_n15792_), .A2(new_n15791_), .A3(new_n15788_), .ZN(new_n15799_));
  AOI21_X1   g15699(.A1(new_n15778_), .A2(new_n15785_), .B(new_n15789_), .ZN(new_n15800_));
  OAI21_X1   g15700(.A1(new_n15799_), .A2(new_n15800_), .B(new_n15796_), .ZN(new_n15801_));
  AOI21_X1   g15701(.A1(new_n15801_), .A2(new_n15798_), .B(new_n15752_), .ZN(new_n15802_));
  INV_X1     g15702(.I(new_n15752_), .ZN(new_n15803_));
  NOR3_X1    g15703(.A1(new_n15799_), .A2(new_n15800_), .A3(new_n15796_), .ZN(new_n15804_));
  AOI21_X1   g15704(.A1(new_n15793_), .A2(new_n15790_), .B(new_n15797_), .ZN(new_n15805_));
  NOR3_X1    g15705(.A1(new_n15804_), .A2(new_n15805_), .A3(new_n15803_), .ZN(new_n15806_));
  OAI21_X1   g15706(.A1(new_n15806_), .A2(new_n15802_), .B(new_n15748_), .ZN(new_n15807_));
  INV_X1     g15707(.I(new_n15748_), .ZN(new_n15808_));
  OAI21_X1   g15708(.A1(new_n15804_), .A2(new_n15805_), .B(new_n15803_), .ZN(new_n15809_));
  NAND3_X1   g15709(.A1(new_n15801_), .A2(new_n15798_), .A3(new_n15752_), .ZN(new_n15810_));
  NAND3_X1   g15710(.A1(new_n15809_), .A2(new_n15810_), .A3(new_n15808_), .ZN(new_n15811_));
  NAND2_X1   g15711(.A1(new_n15585_), .A2(new_n15588_), .ZN(new_n15812_));
  INV_X1     g15712(.I(new_n15812_), .ZN(new_n15813_));
  OAI21_X1   g15713(.A1(new_n15812_), .A2(new_n15392_), .B(new_n15597_), .ZN(new_n15814_));
  OAI22_X1   g15714(.A1(new_n15814_), .A2(new_n15557_), .B1(new_n15371_), .B2(new_n15813_), .ZN(new_n15815_));
  NAND3_X1   g15715(.A1(new_n15807_), .A2(new_n15811_), .A3(new_n15815_), .ZN(new_n15816_));
  AOI21_X1   g15716(.A1(new_n15809_), .A2(new_n15810_), .B(new_n15808_), .ZN(new_n15817_));
  NOR3_X1    g15717(.A1(new_n15806_), .A2(new_n15802_), .A3(new_n15748_), .ZN(new_n15818_));
  INV_X1     g15718(.I(new_n15815_), .ZN(new_n15819_));
  OAI21_X1   g15719(.A1(new_n15818_), .A2(new_n15817_), .B(new_n15819_), .ZN(new_n15820_));
  AOI21_X1   g15720(.A1(new_n15820_), .A2(new_n15816_), .B(new_n15744_), .ZN(new_n15821_));
  NOR3_X1    g15721(.A1(new_n15818_), .A2(new_n15817_), .A3(new_n15819_), .ZN(new_n15822_));
  AOI21_X1   g15722(.A1(new_n15807_), .A2(new_n15811_), .B(new_n15815_), .ZN(new_n15823_));
  NOR3_X1    g15723(.A1(new_n15822_), .A2(new_n15823_), .A3(new_n15743_), .ZN(new_n15824_));
  OAI21_X1   g15724(.A1(new_n15824_), .A2(new_n15821_), .B(new_n15739_), .ZN(new_n15825_));
  INV_X1     g15725(.I(new_n15739_), .ZN(new_n15826_));
  OAI21_X1   g15726(.A1(new_n15822_), .A2(new_n15823_), .B(new_n15743_), .ZN(new_n15827_));
  NAND3_X1   g15727(.A1(new_n15820_), .A2(new_n15816_), .A3(new_n15744_), .ZN(new_n15828_));
  NAND3_X1   g15728(.A1(new_n15827_), .A2(new_n15828_), .A3(new_n15826_), .ZN(new_n15829_));
  AOI22_X1   g15729(.A1(new_n12909_), .A2(new_n5968_), .B1(new_n10949_), .B2(new_n785_), .ZN(new_n15830_));
  OAI21_X1   g15730(.A1(new_n15830_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n15831_));
  XOR2_X1    g15731(.A1(new_n12907_), .A2(new_n15831_), .Z(new_n15832_));
  INV_X1     g15732(.I(new_n15832_), .ZN(new_n15833_));
  NAND3_X1   g15733(.A1(new_n15825_), .A2(new_n15829_), .A3(new_n15833_), .ZN(new_n15834_));
  AOI21_X1   g15734(.A1(new_n15827_), .A2(new_n15828_), .B(new_n15826_), .ZN(new_n15835_));
  NOR3_X1    g15735(.A1(new_n15824_), .A2(new_n15821_), .A3(new_n15739_), .ZN(new_n15836_));
  OAI21_X1   g15736(.A1(new_n15836_), .A2(new_n15835_), .B(new_n15832_), .ZN(new_n15837_));
  AOI21_X1   g15737(.A1(new_n15837_), .A2(new_n15834_), .B(new_n15736_), .ZN(new_n15838_));
  INV_X1     g15738(.I(new_n15736_), .ZN(new_n15839_));
  NOR3_X1    g15739(.A1(new_n15836_), .A2(new_n15835_), .A3(new_n15832_), .ZN(new_n15840_));
  AOI21_X1   g15740(.A1(new_n15825_), .A2(new_n15829_), .B(new_n15833_), .ZN(new_n15841_));
  NOR3_X1    g15741(.A1(new_n15840_), .A2(new_n15841_), .A3(new_n15839_), .ZN(new_n15842_));
  OAI21_X1   g15742(.A1(new_n15842_), .A2(new_n15838_), .B(new_n15734_), .ZN(new_n15843_));
  INV_X1     g15743(.I(new_n15734_), .ZN(new_n15844_));
  OAI21_X1   g15744(.A1(new_n15840_), .A2(new_n15841_), .B(new_n15839_), .ZN(new_n15845_));
  NAND3_X1   g15745(.A1(new_n15837_), .A2(new_n15834_), .A3(new_n15736_), .ZN(new_n15846_));
  NAND3_X1   g15746(.A1(new_n15845_), .A2(new_n15846_), .A3(new_n15844_), .ZN(new_n15847_));
  NOR2_X1    g15747(.A1(new_n15628_), .A2(new_n15633_), .ZN(new_n15848_));
  INV_X1     g15748(.I(new_n15848_), .ZN(new_n15849_));
  AOI21_X1   g15749(.A1(new_n15848_), .A2(new_n15433_), .B(new_n15636_), .ZN(new_n15850_));
  AOI22_X1   g15750(.A1(new_n15850_), .A2(new_n15442_), .B1(new_n15439_), .B2(new_n15849_), .ZN(new_n15851_));
  INV_X1     g15751(.I(new_n15851_), .ZN(new_n15852_));
  NAND3_X1   g15752(.A1(new_n15843_), .A2(new_n15847_), .A3(new_n15852_), .ZN(new_n15853_));
  AOI21_X1   g15753(.A1(new_n15845_), .A2(new_n15846_), .B(new_n15844_), .ZN(new_n15854_));
  NOR3_X1    g15754(.A1(new_n15842_), .A2(new_n15838_), .A3(new_n15734_), .ZN(new_n15855_));
  OAI21_X1   g15755(.A1(new_n15855_), .A2(new_n15854_), .B(new_n15851_), .ZN(new_n15856_));
  AOI21_X1   g15756(.A1(new_n15856_), .A2(new_n15853_), .B(new_n15731_), .ZN(new_n15857_));
  INV_X1     g15757(.I(new_n15665_), .ZN(new_n15858_));
  AOI21_X1   g15758(.A1(new_n15663_), .A2(new_n15664_), .B(new_n15858_), .ZN(new_n15859_));
  NOR3_X1    g15759(.A1(new_n15855_), .A2(new_n15854_), .A3(new_n15851_), .ZN(new_n15860_));
  AOI21_X1   g15760(.A1(new_n15843_), .A2(new_n15847_), .B(new_n15852_), .ZN(new_n15861_));
  NOR3_X1    g15761(.A1(new_n15860_), .A2(new_n15861_), .A3(new_n15859_), .ZN(new_n15862_));
  OAI21_X1   g15762(.A1(new_n15857_), .A2(new_n15862_), .B(new_n15729_), .ZN(new_n15863_));
  INV_X1     g15763(.I(new_n15729_), .ZN(new_n15864_));
  OAI21_X1   g15764(.A1(new_n15860_), .A2(new_n15861_), .B(new_n15859_), .ZN(new_n15865_));
  NAND3_X1   g15765(.A1(new_n15856_), .A2(new_n15853_), .A3(new_n15731_), .ZN(new_n15866_));
  NAND3_X1   g15766(.A1(new_n15866_), .A2(new_n15865_), .A3(new_n15864_), .ZN(new_n15867_));
  OAI22_X1   g15767(.A1(new_n15313_), .A2(new_n8831_), .B1(new_n3040_), .B2(new_n15305_), .ZN(new_n15868_));
  AOI21_X1   g15768(.A1(new_n15868_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n15869_));
  INV_X1     g15769(.I(new_n15869_), .ZN(new_n15870_));
  NOR2_X1    g15770(.A1(new_n15312_), .A2(new_n15870_), .ZN(new_n15871_));
  AOI21_X1   g15771(.A1(new_n15311_), .A2(new_n15308_), .B(new_n15869_), .ZN(new_n15872_));
  NOR2_X1    g15772(.A1(new_n15871_), .A2(new_n15872_), .ZN(new_n15873_));
  INV_X1     g15773(.I(new_n15873_), .ZN(new_n15874_));
  NAND3_X1   g15774(.A1(new_n15874_), .A2(new_n15863_), .A3(new_n15867_), .ZN(new_n15875_));
  AOI21_X1   g15775(.A1(new_n15866_), .A2(new_n15865_), .B(new_n15864_), .ZN(new_n15876_));
  NOR3_X1    g15776(.A1(new_n15857_), .A2(new_n15862_), .A3(new_n15729_), .ZN(new_n15877_));
  OAI21_X1   g15777(.A1(new_n15876_), .A2(new_n15877_), .B(new_n15873_), .ZN(new_n15878_));
  AOI21_X1   g15778(.A1(new_n15875_), .A2(new_n15878_), .B(new_n15726_), .ZN(new_n15879_));
  AND3_X2    g15779(.A1(new_n15875_), .A2(new_n15726_), .A3(new_n15878_), .Z(new_n15880_));
  OAI21_X1   g15780(.A1(new_n15880_), .A2(new_n15879_), .B(new_n15721_), .ZN(new_n15881_));
  OR3_X2     g15781(.A1(new_n15880_), .A2(new_n15721_), .A3(new_n15879_), .Z(new_n15882_));
  AOI21_X1   g15782(.A1(new_n15674_), .A2(new_n15689_), .B(new_n15690_), .ZN(new_n15883_));
  INV_X1     g15783(.I(new_n15883_), .ZN(new_n15884_));
  NAND3_X1   g15784(.A1(new_n15884_), .A2(new_n15881_), .A3(new_n15882_), .ZN(new_n15885_));
  NAND2_X1   g15785(.A1(new_n15882_), .A2(new_n15881_), .ZN(new_n15886_));
  NAND2_X1   g15786(.A1(new_n15886_), .A2(new_n15883_), .ZN(new_n15887_));
  NAND2_X1   g15787(.A1(new_n15885_), .A2(new_n15887_), .ZN(new_n15888_));
  AND3_X2    g15788(.A1(new_n14429_), .A2(new_n14921_), .A3(new_n15151_), .Z(new_n15889_));
  OAI21_X1   g15789(.A1(new_n15889_), .A2(new_n15150_), .B(new_n15545_), .ZN(new_n15890_));
  NOR2_X1    g15790(.A1(new_n15542_), .A2(new_n15702_), .ZN(new_n15891_));
  INV_X1     g15791(.I(new_n15891_), .ZN(new_n15892_));
  OAI21_X1   g15792(.A1(new_n15541_), .A2(new_n15551_), .B(new_n15694_), .ZN(new_n15893_));
  OAI21_X1   g15793(.A1(new_n15890_), .A2(new_n15893_), .B(new_n15892_), .ZN(new_n15894_));
  NAND2_X1   g15794(.A1(new_n15894_), .A2(new_n15888_), .ZN(new_n15895_));
  XOR2_X1    g15795(.A1(new_n15718_), .A2(new_n15895_), .Z(new_n15896_));
  XOR2_X1    g15796(.A1(new_n15896_), .A2(new_n15711_), .Z(\result[7] ));
  AOI21_X1   g15797(.A1(new_n15712_), .A2(new_n15716_), .B(new_n15895_), .ZN(new_n15898_));
  NOR2_X1    g15798(.A1(new_n15152_), .A2(new_n15701_), .ZN(new_n15899_));
  AOI21_X1   g15799(.A1(new_n15542_), .A2(new_n15702_), .B(new_n15704_), .ZN(new_n15900_));
  AOI21_X1   g15800(.A1(new_n15899_), .A2(new_n15900_), .B(new_n15891_), .ZN(new_n15901_));
  NAND2_X1   g15801(.A1(new_n15884_), .A2(new_n15886_), .ZN(new_n15902_));
  OAI22_X1   g15802(.A1(new_n15305_), .A2(new_n8830_), .B1(new_n15114_), .B2(new_n3042_), .ZN(new_n15903_));
  OAI21_X1   g15803(.A1(new_n3040_), .A2(new_n15515_), .B(new_n15903_), .ZN(new_n15904_));
  AOI21_X1   g15804(.A1(new_n15904_), .A2(new_n452_), .B(new_n3040_), .ZN(new_n15905_));
  XOR2_X1    g15805(.A1(new_n15518_), .A2(new_n15905_), .Z(new_n15906_));
  INV_X1     g15806(.I(new_n15721_), .ZN(new_n15907_));
  NAND2_X1   g15807(.A1(new_n15851_), .A2(new_n15729_), .ZN(new_n15908_));
  NAND2_X1   g15808(.A1(new_n15852_), .A2(new_n15864_), .ZN(new_n15909_));
  AOI22_X1   g15809(.A1(new_n15843_), .A2(new_n15847_), .B1(new_n15908_), .B2(new_n15909_), .ZN(new_n15910_));
  NAND2_X1   g15810(.A1(new_n15843_), .A2(new_n15847_), .ZN(new_n15911_));
  XOR2_X1    g15811(.A1(new_n15851_), .A2(new_n15864_), .Z(new_n15912_));
  NOR2_X1    g15812(.A1(new_n15911_), .A2(new_n15912_), .ZN(new_n15913_));
  OAI22_X1   g15813(.A1(new_n15913_), .A2(new_n15910_), .B1(new_n15907_), .B2(new_n15731_), .ZN(new_n15914_));
  NAND2_X1   g15814(.A1(new_n15731_), .A2(new_n15907_), .ZN(new_n15915_));
  NAND2_X1   g15815(.A1(new_n15914_), .A2(new_n15915_), .ZN(new_n15916_));
  OAI22_X1   g15816(.A1(new_n10570_), .A2(new_n6756_), .B1(new_n2258_), .B2(new_n10961_), .ZN(new_n15917_));
  OAI21_X1   g15817(.A1(new_n10564_), .A2(new_n1078_), .B(new_n15917_), .ZN(new_n15918_));
  AOI21_X1   g15818(.A1(new_n15918_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n15919_));
  XNOR2_X1   g15819(.A1(new_n10976_), .A2(new_n15919_), .ZN(new_n15920_));
  INV_X1     g15820(.I(new_n15920_), .ZN(new_n15921_));
  NAND2_X1   g15821(.A1(new_n15911_), .A2(new_n15908_), .ZN(new_n15922_));
  NAND2_X1   g15822(.A1(new_n15922_), .A2(new_n15909_), .ZN(new_n15923_));
  OAI22_X1   g15823(.A1(new_n1851_), .A2(new_n10938_), .B1(new_n10952_), .B2(new_n5966_), .ZN(new_n15924_));
  OAI21_X1   g15824(.A1(new_n10577_), .A2(new_n643_), .B(new_n15924_), .ZN(new_n15925_));
  AOI21_X1   g15825(.A1(new_n15925_), .A2(new_n279_), .B(new_n643_), .ZN(new_n15926_));
  XOR2_X1    g15826(.A1(new_n13544_), .A2(new_n15926_), .Z(new_n15927_));
  NAND2_X1   g15827(.A1(new_n15819_), .A2(new_n15739_), .ZN(new_n15928_));
  NAND2_X1   g15828(.A1(new_n15826_), .A2(new_n15815_), .ZN(new_n15929_));
  AOI22_X1   g15829(.A1(new_n15807_), .A2(new_n15811_), .B1(new_n15928_), .B2(new_n15929_), .ZN(new_n15930_));
  NAND2_X1   g15830(.A1(new_n15807_), .A2(new_n15811_), .ZN(new_n15931_));
  XOR2_X1    g15831(.A1(new_n15815_), .A2(new_n15739_), .Z(new_n15932_));
  NOR2_X1    g15832(.A1(new_n15931_), .A2(new_n15932_), .ZN(new_n15933_));
  OAI22_X1   g15833(.A1(new_n15933_), .A2(new_n15930_), .B1(new_n15844_), .B2(new_n15744_), .ZN(new_n15934_));
  NAND2_X1   g15834(.A1(new_n15744_), .A2(new_n15844_), .ZN(new_n15935_));
  NAND2_X1   g15835(.A1(new_n15934_), .A2(new_n15935_), .ZN(new_n15936_));
  OAI22_X1   g15836(.A1(new_n10589_), .A2(new_n5398_), .B1(new_n12623_), .B2(new_n5336_), .ZN(new_n15937_));
  AOI21_X1   g15837(.A1(new_n15937_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n15938_));
  XOR2_X1    g15838(.A1(new_n12622_), .A2(new_n15938_), .Z(new_n15939_));
  INV_X1     g15839(.I(new_n15939_), .ZN(new_n15940_));
  NAND2_X1   g15840(.A1(new_n15931_), .A2(new_n15928_), .ZN(new_n15941_));
  NAND2_X1   g15841(.A1(new_n15941_), .A2(new_n15929_), .ZN(new_n15942_));
  INV_X1     g15842(.I(new_n15942_), .ZN(new_n15943_));
  OAI22_X1   g15843(.A1(new_n10606_), .A2(new_n1239_), .B1(new_n4981_), .B2(new_n10901_), .ZN(new_n15944_));
  AOI21_X1   g15844(.A1(new_n15944_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n15945_));
  XOR2_X1    g15845(.A1(new_n12211_), .A2(new_n15945_), .Z(new_n15946_));
  INV_X1     g15846(.I(new_n15946_), .ZN(new_n15947_));
  NOR2_X1    g15847(.A1(new_n15803_), .A2(new_n15796_), .ZN(new_n15948_));
  NAND2_X1   g15848(.A1(new_n15803_), .A2(new_n15796_), .ZN(new_n15949_));
  NAND3_X1   g15849(.A1(new_n15793_), .A2(new_n15790_), .A3(new_n15808_), .ZN(new_n15950_));
  OAI21_X1   g15850(.A1(new_n15799_), .A2(new_n15800_), .B(new_n15748_), .ZN(new_n15951_));
  NAND2_X1   g15851(.A1(new_n15951_), .A2(new_n15950_), .ZN(new_n15952_));
  AOI21_X1   g15852(.A1(new_n15952_), .A2(new_n15949_), .B(new_n15948_), .ZN(new_n15953_));
  OAI22_X1   g15853(.A1(new_n10844_), .A2(new_n4529_), .B1(new_n4527_), .B2(new_n10856_), .ZN(new_n15954_));
  OAI21_X1   g15854(.A1(new_n10870_), .A2(new_n79_), .B(new_n15954_), .ZN(new_n15955_));
  AOI21_X1   g15855(.A1(new_n15955_), .A2(new_n72_), .B(new_n79_), .ZN(new_n15956_));
  XOR2_X1    g15856(.A1(new_n11648_), .A2(new_n15956_), .Z(new_n15957_));
  INV_X1     g15857(.I(new_n15957_), .ZN(new_n15958_));
  AOI21_X1   g15858(.A1(new_n15779_), .A2(new_n15780_), .B(new_n15781_), .ZN(new_n15959_));
  NOR2_X1    g15859(.A1(new_n15959_), .A2(new_n15782_), .ZN(new_n15960_));
  NAND2_X1   g15860(.A1(new_n15755_), .A2(new_n15756_), .ZN(new_n15961_));
  NOR2_X1    g15861(.A1(new_n10631_), .A2(new_n511_), .ZN(new_n15962_));
  OAI22_X1   g15862(.A1(new_n10633_), .A2(new_n88_), .B1(new_n92_), .B2(new_n11264_), .ZN(new_n15963_));
  OAI21_X1   g15863(.A1(new_n15962_), .A2(new_n15963_), .B(new_n961_), .ZN(new_n15964_));
  NOR2_X1    g15864(.A1(new_n11445_), .A2(new_n15964_), .ZN(new_n15965_));
  AOI21_X1   g15865(.A1(new_n15961_), .A2(new_n15761_), .B(new_n15965_), .ZN(new_n15966_));
  NOR2_X1    g15866(.A1(new_n15765_), .A2(new_n15764_), .ZN(new_n15967_));
  INV_X1     g15867(.I(new_n15965_), .ZN(new_n15968_));
  NOR3_X1    g15868(.A1(new_n15967_), .A2(new_n15762_), .A3(new_n15968_), .ZN(new_n15969_));
  OAI22_X1   g15869(.A1(new_n10881_), .A2(new_n4781_), .B1(new_n10868_), .B2(new_n4612_), .ZN(new_n15970_));
  OAI21_X1   g15870(.A1(new_n10619_), .A2(new_n1128_), .B(new_n15970_), .ZN(new_n15971_));
  AOI21_X1   g15871(.A1(new_n15971_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n15972_));
  XOR2_X1    g15872(.A1(new_n12074_), .A2(new_n15972_), .Z(new_n15973_));
  NOR3_X1    g15873(.A1(new_n15969_), .A2(new_n15966_), .A3(new_n15973_), .ZN(new_n15974_));
  OAI21_X1   g15874(.A1(new_n15967_), .A2(new_n15762_), .B(new_n15968_), .ZN(new_n15975_));
  NAND3_X1   g15875(.A1(new_n15961_), .A2(new_n15761_), .A3(new_n15965_), .ZN(new_n15976_));
  INV_X1     g15876(.I(new_n15973_), .ZN(new_n15977_));
  AOI21_X1   g15877(.A1(new_n15975_), .A2(new_n15976_), .B(new_n15977_), .ZN(new_n15978_));
  OAI21_X1   g15878(.A1(new_n15974_), .A2(new_n15978_), .B(new_n15960_), .ZN(new_n15979_));
  NOR2_X1    g15879(.A1(new_n15763_), .A2(new_n15766_), .ZN(new_n15980_));
  INV_X1     g15880(.I(new_n15782_), .ZN(new_n15981_));
  OAI21_X1   g15881(.A1(new_n15980_), .A2(new_n15781_), .B(new_n15981_), .ZN(new_n15982_));
  NAND3_X1   g15882(.A1(new_n15975_), .A2(new_n15976_), .A3(new_n15977_), .ZN(new_n15983_));
  OAI21_X1   g15883(.A1(new_n15969_), .A2(new_n15966_), .B(new_n15973_), .ZN(new_n15984_));
  NAND3_X1   g15884(.A1(new_n15982_), .A2(new_n15984_), .A3(new_n15983_), .ZN(new_n15985_));
  AOI21_X1   g15885(.A1(new_n15979_), .A2(new_n15985_), .B(new_n15958_), .ZN(new_n15986_));
  AOI21_X1   g15886(.A1(new_n15983_), .A2(new_n15984_), .B(new_n15982_), .ZN(new_n15987_));
  NOR3_X1    g15887(.A1(new_n15974_), .A2(new_n15978_), .A3(new_n15960_), .ZN(new_n15988_));
  NOR3_X1    g15888(.A1(new_n15987_), .A2(new_n15988_), .A3(new_n15957_), .ZN(new_n15989_));
  NOR2_X1    g15889(.A1(new_n15789_), .A2(new_n15748_), .ZN(new_n15990_));
  NOR2_X1    g15890(.A1(new_n15788_), .A2(new_n15808_), .ZN(new_n15991_));
  NOR3_X1    g15891(.A1(new_n15792_), .A2(new_n15791_), .A3(new_n15991_), .ZN(new_n15992_));
  NOR2_X1    g15892(.A1(new_n15992_), .A2(new_n15990_), .ZN(new_n15993_));
  NOR3_X1    g15893(.A1(new_n15989_), .A2(new_n15986_), .A3(new_n15993_), .ZN(new_n15994_));
  OAI21_X1   g15894(.A1(new_n15987_), .A2(new_n15988_), .B(new_n15957_), .ZN(new_n15995_));
  NAND3_X1   g15895(.A1(new_n15979_), .A2(new_n15985_), .A3(new_n15958_), .ZN(new_n15996_));
  INV_X1     g15896(.I(new_n15993_), .ZN(new_n15997_));
  AOI21_X1   g15897(.A1(new_n15995_), .A2(new_n15996_), .B(new_n15997_), .ZN(new_n15998_));
  OAI21_X1   g15898(.A1(new_n15994_), .A2(new_n15998_), .B(new_n15953_), .ZN(new_n15999_));
  INV_X1     g15899(.I(new_n15948_), .ZN(new_n16000_));
  NOR3_X1    g15900(.A1(new_n15799_), .A2(new_n15800_), .A3(new_n15748_), .ZN(new_n16001_));
  AOI21_X1   g15901(.A1(new_n15793_), .A2(new_n15790_), .B(new_n15808_), .ZN(new_n16002_));
  OAI21_X1   g15902(.A1(new_n16001_), .A2(new_n16002_), .B(new_n15949_), .ZN(new_n16003_));
  NAND2_X1   g15903(.A1(new_n16003_), .A2(new_n16000_), .ZN(new_n16004_));
  NAND3_X1   g15904(.A1(new_n15995_), .A2(new_n15996_), .A3(new_n15997_), .ZN(new_n16005_));
  OAI21_X1   g15905(.A1(new_n15989_), .A2(new_n15986_), .B(new_n15993_), .ZN(new_n16006_));
  NAND3_X1   g15906(.A1(new_n16006_), .A2(new_n16005_), .A3(new_n16004_), .ZN(new_n16007_));
  AOI21_X1   g15907(.A1(new_n15999_), .A2(new_n16007_), .B(new_n15947_), .ZN(new_n16008_));
  AOI21_X1   g15908(.A1(new_n16006_), .A2(new_n16005_), .B(new_n16004_), .ZN(new_n16009_));
  NOR3_X1    g15909(.A1(new_n15994_), .A2(new_n15998_), .A3(new_n15953_), .ZN(new_n16010_));
  NOR3_X1    g15910(.A1(new_n16010_), .A2(new_n16009_), .A3(new_n15946_), .ZN(new_n16011_));
  OAI22_X1   g15911(.A1(new_n10583_), .A2(new_n1620_), .B1(new_n5420_), .B2(new_n10928_), .ZN(new_n16012_));
  AOI21_X1   g15912(.A1(new_n16012_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n16013_));
  XNOR2_X1   g15913(.A1(new_n13378_), .A2(new_n16013_), .ZN(new_n16014_));
  NOR3_X1    g15914(.A1(new_n16008_), .A2(new_n16011_), .A3(new_n16014_), .ZN(new_n16015_));
  OAI21_X1   g15915(.A1(new_n16010_), .A2(new_n16009_), .B(new_n15946_), .ZN(new_n16016_));
  NAND3_X1   g15916(.A1(new_n15999_), .A2(new_n16007_), .A3(new_n15947_), .ZN(new_n16017_));
  INV_X1     g15917(.I(new_n16014_), .ZN(new_n16018_));
  AOI21_X1   g15918(.A1(new_n16016_), .A2(new_n16017_), .B(new_n16018_), .ZN(new_n16019_));
  OAI21_X1   g15919(.A1(new_n16015_), .A2(new_n16019_), .B(new_n15943_), .ZN(new_n16020_));
  NAND3_X1   g15920(.A1(new_n16016_), .A2(new_n16017_), .A3(new_n16018_), .ZN(new_n16021_));
  OAI21_X1   g15921(.A1(new_n16008_), .A2(new_n16011_), .B(new_n16014_), .ZN(new_n16022_));
  NAND3_X1   g15922(.A1(new_n16022_), .A2(new_n16021_), .A3(new_n15942_), .ZN(new_n16023_));
  AOI21_X1   g15923(.A1(new_n16020_), .A2(new_n16023_), .B(new_n15940_), .ZN(new_n16024_));
  AOI21_X1   g15924(.A1(new_n16022_), .A2(new_n16021_), .B(new_n15942_), .ZN(new_n16025_));
  NOR3_X1    g15925(.A1(new_n16015_), .A2(new_n16019_), .A3(new_n15943_), .ZN(new_n16026_));
  NOR3_X1    g15926(.A1(new_n16026_), .A2(new_n16025_), .A3(new_n15939_), .ZN(new_n16027_));
  NOR2_X1    g15927(.A1(new_n16027_), .A2(new_n16024_), .ZN(new_n16028_));
  NOR2_X1    g15928(.A1(new_n15839_), .A2(new_n15832_), .ZN(new_n16029_));
  INV_X1     g15929(.I(new_n16029_), .ZN(new_n16030_));
  NAND2_X1   g15930(.A1(new_n15839_), .A2(new_n15832_), .ZN(new_n16031_));
  NOR3_X1    g15931(.A1(new_n15836_), .A2(new_n15835_), .A3(new_n15734_), .ZN(new_n16032_));
  AOI21_X1   g15932(.A1(new_n15825_), .A2(new_n15829_), .B(new_n15844_), .ZN(new_n16033_));
  OAI21_X1   g15933(.A1(new_n16032_), .A2(new_n16033_), .B(new_n16031_), .ZN(new_n16034_));
  NAND2_X1   g15934(.A1(new_n16034_), .A2(new_n16030_), .ZN(new_n16035_));
  NAND2_X1   g15935(.A1(new_n16028_), .A2(new_n16035_), .ZN(new_n16036_));
  OAI21_X1   g15936(.A1(new_n16026_), .A2(new_n16025_), .B(new_n15939_), .ZN(new_n16037_));
  NAND3_X1   g15937(.A1(new_n16020_), .A2(new_n16023_), .A3(new_n15940_), .ZN(new_n16038_));
  NAND2_X1   g15938(.A1(new_n16037_), .A2(new_n16038_), .ZN(new_n16039_));
  NAND3_X1   g15939(.A1(new_n15825_), .A2(new_n15829_), .A3(new_n15844_), .ZN(new_n16040_));
  OAI21_X1   g15940(.A1(new_n15836_), .A2(new_n15835_), .B(new_n15734_), .ZN(new_n16041_));
  NAND2_X1   g15941(.A1(new_n16041_), .A2(new_n16040_), .ZN(new_n16042_));
  AOI21_X1   g15942(.A1(new_n16042_), .A2(new_n16031_), .B(new_n16029_), .ZN(new_n16043_));
  NAND2_X1   g15943(.A1(new_n16039_), .A2(new_n16043_), .ZN(new_n16044_));
  AOI21_X1   g15944(.A1(new_n16036_), .A2(new_n16044_), .B(new_n15936_), .ZN(new_n16045_));
  INV_X1     g15945(.I(new_n15936_), .ZN(new_n16046_));
  NOR2_X1    g15946(.A1(new_n16039_), .A2(new_n16043_), .ZN(new_n16047_));
  NOR2_X1    g15947(.A1(new_n16028_), .A2(new_n16035_), .ZN(new_n16048_));
  NOR3_X1    g15948(.A1(new_n16048_), .A2(new_n16047_), .A3(new_n16046_), .ZN(new_n16049_));
  OAI21_X1   g15949(.A1(new_n16045_), .A2(new_n16049_), .B(new_n15927_), .ZN(new_n16050_));
  INV_X1     g15950(.I(new_n15927_), .ZN(new_n16051_));
  OAI21_X1   g15951(.A1(new_n16048_), .A2(new_n16047_), .B(new_n16046_), .ZN(new_n16052_));
  NAND3_X1   g15952(.A1(new_n16036_), .A2(new_n16044_), .A3(new_n15936_), .ZN(new_n16053_));
  NAND3_X1   g15953(.A1(new_n16052_), .A2(new_n16053_), .A3(new_n16051_), .ZN(new_n16054_));
  OAI22_X1   g15954(.A1(new_n14276_), .A2(new_n2718_), .B1(new_n7836_), .B2(new_n14594_), .ZN(new_n16055_));
  OAI21_X1   g15955(.A1(new_n14886_), .A2(new_n2495_), .B(new_n16055_), .ZN(new_n16056_));
  AOI21_X1   g15956(.A1(new_n16056_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n16057_));
  XOR2_X1    g15957(.A1(new_n14891_), .A2(new_n16057_), .Z(new_n16058_));
  INV_X1     g15958(.I(new_n16058_), .ZN(new_n16059_));
  NAND3_X1   g15959(.A1(new_n16050_), .A2(new_n16054_), .A3(new_n16059_), .ZN(new_n16060_));
  AOI21_X1   g15960(.A1(new_n16052_), .A2(new_n16053_), .B(new_n16051_), .ZN(new_n16061_));
  NOR3_X1    g15961(.A1(new_n16045_), .A2(new_n16049_), .A3(new_n15927_), .ZN(new_n16062_));
  OAI21_X1   g15962(.A1(new_n16062_), .A2(new_n16061_), .B(new_n16058_), .ZN(new_n16063_));
  AOI21_X1   g15963(.A1(new_n16063_), .A2(new_n16060_), .B(new_n15923_), .ZN(new_n16064_));
  INV_X1     g15964(.I(new_n15923_), .ZN(new_n16065_));
  NOR3_X1    g15965(.A1(new_n16062_), .A2(new_n16061_), .A3(new_n16058_), .ZN(new_n16066_));
  AOI21_X1   g15966(.A1(new_n16050_), .A2(new_n16054_), .B(new_n16059_), .ZN(new_n16067_));
  NOR3_X1    g15967(.A1(new_n16066_), .A2(new_n16067_), .A3(new_n16065_), .ZN(new_n16068_));
  OAI21_X1   g15968(.A1(new_n16068_), .A2(new_n16064_), .B(new_n15921_), .ZN(new_n16069_));
  OAI21_X1   g15969(.A1(new_n16066_), .A2(new_n16067_), .B(new_n16065_), .ZN(new_n16070_));
  NAND3_X1   g15970(.A1(new_n16063_), .A2(new_n16060_), .A3(new_n15923_), .ZN(new_n16071_));
  NAND3_X1   g15971(.A1(new_n16070_), .A2(new_n16071_), .A3(new_n15920_), .ZN(new_n16072_));
  AOI21_X1   g15972(.A1(new_n15725_), .A2(new_n15722_), .B(new_n15873_), .ZN(new_n16073_));
  INV_X1     g15973(.I(new_n16073_), .ZN(new_n16074_));
  NAND3_X1   g15974(.A1(new_n15725_), .A2(new_n15722_), .A3(new_n15873_), .ZN(new_n16075_));
  NOR3_X1    g15975(.A1(new_n15876_), .A2(new_n15877_), .A3(new_n15721_), .ZN(new_n16076_));
  AOI21_X1   g15976(.A1(new_n15863_), .A2(new_n15867_), .B(new_n15907_), .ZN(new_n16077_));
  OAI21_X1   g15977(.A1(new_n16076_), .A2(new_n16077_), .B(new_n16075_), .ZN(new_n16078_));
  NAND2_X1   g15978(.A1(new_n16078_), .A2(new_n16074_), .ZN(new_n16079_));
  NAND3_X1   g15979(.A1(new_n16079_), .A2(new_n16069_), .A3(new_n16072_), .ZN(new_n16080_));
  AOI21_X1   g15980(.A1(new_n16070_), .A2(new_n16071_), .B(new_n15920_), .ZN(new_n16081_));
  NOR3_X1    g15981(.A1(new_n16068_), .A2(new_n16064_), .A3(new_n15921_), .ZN(new_n16082_));
  NAND3_X1   g15982(.A1(new_n15863_), .A2(new_n15867_), .A3(new_n15907_), .ZN(new_n16083_));
  OAI21_X1   g15983(.A1(new_n15876_), .A2(new_n15877_), .B(new_n15721_), .ZN(new_n16084_));
  NAND2_X1   g15984(.A1(new_n16084_), .A2(new_n16083_), .ZN(new_n16085_));
  AOI21_X1   g15985(.A1(new_n16085_), .A2(new_n16075_), .B(new_n16073_), .ZN(new_n16086_));
  OAI21_X1   g15986(.A1(new_n16081_), .A2(new_n16082_), .B(new_n16086_), .ZN(new_n16087_));
  AOI21_X1   g15987(.A1(new_n16087_), .A2(new_n16080_), .B(new_n15916_), .ZN(new_n16088_));
  INV_X1     g15988(.I(new_n15916_), .ZN(new_n16089_));
  NOR3_X1    g15989(.A1(new_n16086_), .A2(new_n16082_), .A3(new_n16081_), .ZN(new_n16090_));
  AOI21_X1   g15990(.A1(new_n16069_), .A2(new_n16072_), .B(new_n16079_), .ZN(new_n16091_));
  NOR3_X1    g15991(.A1(new_n16091_), .A2(new_n16089_), .A3(new_n16090_), .ZN(new_n16092_));
  OAI21_X1   g15992(.A1(new_n16092_), .A2(new_n16088_), .B(new_n15906_), .ZN(new_n16093_));
  INV_X1     g15993(.I(new_n15906_), .ZN(new_n16094_));
  OAI21_X1   g15994(.A1(new_n16091_), .A2(new_n16090_), .B(new_n16089_), .ZN(new_n16095_));
  NAND3_X1   g15995(.A1(new_n16087_), .A2(new_n16080_), .A3(new_n15916_), .ZN(new_n16096_));
  NAND3_X1   g15996(.A1(new_n16095_), .A2(new_n16096_), .A3(new_n16094_), .ZN(new_n16097_));
  AOI22_X1   g15997(.A1(new_n16093_), .A2(new_n16097_), .B1(new_n15885_), .B2(new_n15887_), .ZN(new_n16098_));
  XOR2_X1    g15998(.A1(new_n16098_), .A2(new_n15902_), .Z(new_n16099_));
  XOR2_X1    g15999(.A1(new_n16099_), .A2(new_n15901_), .Z(new_n16100_));
  XOR2_X1    g16000(.A1(new_n15898_), .A2(new_n16100_), .Z(\result[8] ));
  AOI21_X1   g16001(.A1(new_n15327_), .A2(new_n15532_), .B(new_n15715_), .ZN(new_n16102_));
  NOR3_X1    g16002(.A1(new_n15536_), .A2(new_n15540_), .A3(new_n15711_), .ZN(new_n16103_));
  INV_X1     g16003(.I(new_n15895_), .ZN(new_n16104_));
  OAI21_X1   g16004(.A1(new_n16103_), .A2(new_n16102_), .B(new_n16104_), .ZN(new_n16105_));
  XOR2_X1    g16005(.A1(new_n16099_), .A2(new_n15894_), .Z(new_n16106_));
  INV_X1     g16006(.I(new_n15886_), .ZN(new_n16107_));
  AOI21_X1   g16007(.A1(new_n16095_), .A2(new_n16096_), .B(new_n16094_), .ZN(new_n16108_));
  NOR3_X1    g16008(.A1(new_n16092_), .A2(new_n16088_), .A3(new_n15906_), .ZN(new_n16109_));
  NOR3_X1    g16009(.A1(new_n16109_), .A2(new_n16108_), .A3(new_n15884_), .ZN(new_n16110_));
  OAI21_X1   g16010(.A1(new_n16109_), .A2(new_n16108_), .B(new_n15884_), .ZN(new_n16111_));
  AOI21_X1   g16011(.A1(new_n16107_), .A2(new_n16111_), .B(new_n16110_), .ZN(new_n16112_));
  NAND2_X1   g16012(.A1(new_n15894_), .A2(new_n16112_), .ZN(new_n16113_));
  AOI22_X1   g16013(.A1(new_n14281_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n14274_), .ZN(new_n16114_));
  OAI21_X1   g16014(.A1(new_n16114_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n16115_));
  XOR2_X1    g16015(.A1(new_n14280_), .A2(new_n16115_), .Z(new_n16116_));
  NAND2_X1   g16016(.A1(new_n16046_), .A2(new_n15927_), .ZN(new_n16117_));
  NAND2_X1   g16017(.A1(new_n15936_), .A2(new_n16051_), .ZN(new_n16118_));
  NAND2_X1   g16018(.A1(new_n16117_), .A2(new_n16118_), .ZN(new_n16119_));
  XOR2_X1    g16019(.A1(new_n15936_), .A2(new_n15927_), .Z(new_n16120_));
  NOR2_X1    g16020(.A1(new_n16039_), .A2(new_n16120_), .ZN(new_n16121_));
  AOI21_X1   g16021(.A1(new_n16039_), .A2(new_n16119_), .B(new_n16121_), .ZN(new_n16122_));
  AOI21_X1   g16022(.A1(new_n15921_), .A2(new_n16043_), .B(new_n16122_), .ZN(new_n16123_));
  NOR2_X1    g16023(.A1(new_n15921_), .A2(new_n16043_), .ZN(new_n16124_));
  NOR2_X1    g16024(.A1(new_n16123_), .A2(new_n16124_), .ZN(new_n16125_));
  INV_X1     g16025(.I(new_n16125_), .ZN(new_n16126_));
  AOI22_X1   g16026(.A1(new_n15072_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n10962_), .ZN(new_n16127_));
  OAI21_X1   g16027(.A1(new_n16127_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n16128_));
  NOR2_X1    g16028(.A1(new_n15071_), .A2(new_n16128_), .ZN(new_n16129_));
  INV_X1     g16029(.I(new_n16128_), .ZN(new_n16130_));
  NOR2_X1    g16030(.A1(new_n14053_), .A2(new_n16130_), .ZN(new_n16131_));
  NOR2_X1    g16031(.A1(new_n16129_), .A2(new_n16131_), .ZN(new_n16132_));
  INV_X1     g16032(.I(new_n16132_), .ZN(new_n16133_));
  INV_X1     g16033(.I(new_n16118_), .ZN(new_n16134_));
  AOI21_X1   g16034(.A1(new_n16039_), .A2(new_n16117_), .B(new_n16134_), .ZN(new_n16135_));
  OAI22_X1   g16035(.A1(new_n10913_), .A2(new_n5398_), .B1(new_n12768_), .B2(new_n5336_), .ZN(new_n16136_));
  AOI21_X1   g16036(.A1(new_n16136_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n16137_));
  XOR2_X1    g16037(.A1(new_n12767_), .A2(new_n16137_), .Z(new_n16138_));
  NAND2_X1   g16038(.A1(new_n15995_), .A2(new_n15996_), .ZN(new_n16139_));
  NAND2_X1   g16039(.A1(new_n15993_), .A2(new_n15946_), .ZN(new_n16140_));
  NAND2_X1   g16040(.A1(new_n15997_), .A2(new_n15947_), .ZN(new_n16141_));
  NAND2_X1   g16041(.A1(new_n16141_), .A2(new_n16140_), .ZN(new_n16142_));
  XOR2_X1    g16042(.A1(new_n15993_), .A2(new_n15947_), .Z(new_n16143_));
  NOR2_X1    g16043(.A1(new_n16143_), .A2(new_n16139_), .ZN(new_n16144_));
  AOI21_X1   g16044(.A1(new_n16139_), .A2(new_n16142_), .B(new_n16144_), .ZN(new_n16145_));
  NOR2_X1    g16045(.A1(new_n16004_), .A2(new_n15940_), .ZN(new_n16146_));
  NOR2_X1    g16046(.A1(new_n16145_), .A2(new_n16146_), .ZN(new_n16147_));
  NOR2_X1    g16047(.A1(new_n15953_), .A2(new_n15939_), .ZN(new_n16148_));
  OR2_X2     g16048(.A1(new_n16147_), .A2(new_n16148_), .Z(new_n16149_));
  AOI22_X1   g16049(.A1(new_n10625_), .A2(new_n4526_), .B1(new_n4570_), .B2(new_n10857_), .ZN(new_n16150_));
  AOI21_X1   g16050(.A1(new_n101_), .A2(new_n10875_), .B(new_n16150_), .ZN(new_n16151_));
  OAI21_X1   g16051(.A1(new_n16151_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n16152_));
  XNOR2_X1   g16052(.A1(new_n11722_), .A2(new_n16152_), .ZN(new_n16153_));
  INV_X1     g16053(.I(new_n16153_), .ZN(new_n16154_));
  NAND2_X1   g16054(.A1(new_n15961_), .A2(new_n15761_), .ZN(new_n16155_));
  INV_X1     g16055(.I(new_n16155_), .ZN(new_n16156_));
  OAI21_X1   g16056(.A1(new_n15982_), .A2(new_n15965_), .B(new_n16156_), .ZN(new_n16157_));
  NAND2_X1   g16057(.A1(new_n15982_), .A2(new_n15965_), .ZN(new_n16158_));
  NAND2_X1   g16058(.A1(new_n16157_), .A2(new_n16158_), .ZN(new_n16159_));
  INV_X1     g16059(.I(new_n16159_), .ZN(new_n16160_));
  NOR2_X1    g16060(.A1(new_n10631_), .A2(new_n88_), .ZN(new_n16161_));
  INV_X1     g16061(.I(new_n16161_), .ZN(new_n16162_));
  AOI22_X1   g16062(.A1(new_n10843_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n10833_), .ZN(new_n16163_));
  AOI21_X1   g16063(.A1(new_n16162_), .A2(new_n16163_), .B(new_n82_), .ZN(new_n16164_));
  NAND2_X1   g16064(.A1(new_n11607_), .A2(new_n16164_), .ZN(new_n16165_));
  INV_X1     g16065(.I(new_n16165_), .ZN(new_n16166_));
  OAI21_X1   g16066(.A1(new_n15967_), .A2(new_n15761_), .B(new_n16166_), .ZN(new_n16167_));
  NAND3_X1   g16067(.A1(new_n15961_), .A2(new_n15762_), .A3(new_n16165_), .ZN(new_n16168_));
  AOI21_X1   g16068(.A1(new_n16167_), .A2(new_n16168_), .B(new_n15961_), .ZN(new_n16169_));
  AOI21_X1   g16069(.A1(new_n15961_), .A2(new_n15762_), .B(new_n16165_), .ZN(new_n16170_));
  NOR3_X1    g16070(.A1(new_n15967_), .A2(new_n15761_), .A3(new_n16166_), .ZN(new_n16171_));
  NOR3_X1    g16071(.A1(new_n16171_), .A2(new_n16170_), .A3(new_n15967_), .ZN(new_n16172_));
  NOR2_X1    g16072(.A1(new_n16172_), .A2(new_n16169_), .ZN(new_n16173_));
  OAI22_X1   g16073(.A1(new_n10619_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10881_), .ZN(new_n16174_));
  OAI21_X1   g16074(.A1(new_n1128_), .A2(new_n10611_), .B(new_n16174_), .ZN(new_n16175_));
  AOI21_X1   g16075(.A1(new_n16175_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n16176_));
  XOR2_X1    g16076(.A1(new_n12090_), .A2(new_n16176_), .Z(new_n16177_));
  INV_X1     g16077(.I(new_n16177_), .ZN(new_n16178_));
  NAND2_X1   g16078(.A1(new_n16173_), .A2(new_n16178_), .ZN(new_n16179_));
  OAI21_X1   g16079(.A1(new_n16171_), .A2(new_n16170_), .B(new_n15967_), .ZN(new_n16180_));
  NAND3_X1   g16080(.A1(new_n16167_), .A2(new_n16168_), .A3(new_n15961_), .ZN(new_n16181_));
  NAND2_X1   g16081(.A1(new_n16180_), .A2(new_n16181_), .ZN(new_n16182_));
  NAND2_X1   g16082(.A1(new_n16182_), .A2(new_n16177_), .ZN(new_n16183_));
  NAND2_X1   g16083(.A1(new_n16179_), .A2(new_n16183_), .ZN(new_n16184_));
  NAND2_X1   g16084(.A1(new_n16184_), .A2(new_n16160_), .ZN(new_n16185_));
  NAND3_X1   g16085(.A1(new_n16159_), .A2(new_n16179_), .A3(new_n16183_), .ZN(new_n16186_));
  AOI21_X1   g16086(.A1(new_n16185_), .A2(new_n16186_), .B(new_n16154_), .ZN(new_n16187_));
  AOI21_X1   g16087(.A1(new_n16179_), .A2(new_n16183_), .B(new_n16159_), .ZN(new_n16188_));
  INV_X1     g16088(.I(new_n16186_), .ZN(new_n16189_));
  NOR3_X1    g16089(.A1(new_n16189_), .A2(new_n16153_), .A3(new_n16188_), .ZN(new_n16190_));
  NOR2_X1    g16090(.A1(new_n15973_), .A2(new_n15957_), .ZN(new_n16191_));
  INV_X1     g16091(.I(new_n16191_), .ZN(new_n16192_));
  NAND2_X1   g16092(.A1(new_n15975_), .A2(new_n15976_), .ZN(new_n16193_));
  NOR2_X1    g16093(.A1(new_n15960_), .A2(new_n16193_), .ZN(new_n16194_));
  NOR2_X1    g16094(.A1(new_n15969_), .A2(new_n15966_), .ZN(new_n16195_));
  NOR2_X1    g16095(.A1(new_n15982_), .A2(new_n16195_), .ZN(new_n16196_));
  OAI22_X1   g16096(.A1(new_n16196_), .A2(new_n16194_), .B1(new_n15958_), .B2(new_n15977_), .ZN(new_n16197_));
  NAND2_X1   g16097(.A1(new_n16197_), .A2(new_n16192_), .ZN(new_n16198_));
  AOI22_X1   g16098(.A1(new_n12578_), .A2(new_n5783_), .B1(new_n247_), .B2(new_n10600_), .ZN(new_n16199_));
  OAI21_X1   g16099(.A1(new_n16199_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n16200_));
  XNOR2_X1   g16100(.A1(new_n12576_), .A2(new_n16200_), .ZN(new_n16201_));
  INV_X1     g16101(.I(new_n16201_), .ZN(new_n16202_));
  NOR2_X1    g16102(.A1(new_n16198_), .A2(new_n16202_), .ZN(new_n16203_));
  AOI21_X1   g16103(.A1(new_n16197_), .A2(new_n16192_), .B(new_n16201_), .ZN(new_n16204_));
  OAI22_X1   g16104(.A1(new_n16190_), .A2(new_n16187_), .B1(new_n16204_), .B2(new_n16203_), .ZN(new_n16205_));
  OAI21_X1   g16105(.A1(new_n16189_), .A2(new_n16188_), .B(new_n16153_), .ZN(new_n16206_));
  NAND3_X1   g16106(.A1(new_n16185_), .A2(new_n16154_), .A3(new_n16186_), .ZN(new_n16207_));
  AOI21_X1   g16107(.A1(new_n16197_), .A2(new_n16192_), .B(new_n16202_), .ZN(new_n16208_));
  INV_X1     g16108(.I(new_n16208_), .ZN(new_n16209_));
  NAND3_X1   g16109(.A1(new_n16197_), .A2(new_n16192_), .A3(new_n16202_), .ZN(new_n16210_));
  NAND2_X1   g16110(.A1(new_n16209_), .A2(new_n16210_), .ZN(new_n16211_));
  NAND3_X1   g16111(.A1(new_n16211_), .A2(new_n16206_), .A3(new_n16207_), .ZN(new_n16212_));
  NAND2_X1   g16112(.A1(new_n16139_), .A2(new_n16140_), .ZN(new_n16213_));
  NAND2_X1   g16113(.A1(new_n16213_), .A2(new_n16141_), .ZN(new_n16214_));
  NAND3_X1   g16114(.A1(new_n16205_), .A2(new_n16212_), .A3(new_n16214_), .ZN(new_n16215_));
  INV_X1     g16115(.I(new_n16203_), .ZN(new_n16216_));
  INV_X1     g16116(.I(new_n16204_), .ZN(new_n16217_));
  AOI22_X1   g16117(.A1(new_n16206_), .A2(new_n16207_), .B1(new_n16216_), .B2(new_n16217_), .ZN(new_n16218_));
  INV_X1     g16118(.I(new_n16210_), .ZN(new_n16219_));
  NOR2_X1    g16119(.A1(new_n16219_), .A2(new_n16208_), .ZN(new_n16220_));
  NOR3_X1    g16120(.A1(new_n16220_), .A2(new_n16190_), .A3(new_n16187_), .ZN(new_n16221_));
  INV_X1     g16121(.I(new_n16214_), .ZN(new_n16222_));
  OAI21_X1   g16122(.A1(new_n16218_), .A2(new_n16221_), .B(new_n16222_), .ZN(new_n16223_));
  OAI22_X1   g16123(.A1(new_n13395_), .A2(new_n5420_), .B1(new_n1620_), .B2(new_n10938_), .ZN(new_n16224_));
  AOI21_X1   g16124(.A1(new_n16224_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n16225_));
  XOR2_X1    g16125(.A1(new_n13394_), .A2(new_n16225_), .Z(new_n16226_));
  INV_X1     g16126(.I(new_n16226_), .ZN(new_n16227_));
  NAND3_X1   g16127(.A1(new_n16223_), .A2(new_n16215_), .A3(new_n16227_), .ZN(new_n16228_));
  NOR3_X1    g16128(.A1(new_n16218_), .A2(new_n16221_), .A3(new_n16222_), .ZN(new_n16229_));
  AOI21_X1   g16129(.A1(new_n16205_), .A2(new_n16212_), .B(new_n16214_), .ZN(new_n16230_));
  OAI21_X1   g16130(.A1(new_n16229_), .A2(new_n16230_), .B(new_n16226_), .ZN(new_n16231_));
  AOI21_X1   g16131(.A1(new_n16231_), .A2(new_n16228_), .B(new_n16149_), .ZN(new_n16232_));
  NOR2_X1    g16132(.A1(new_n16147_), .A2(new_n16148_), .ZN(new_n16233_));
  NOR3_X1    g16133(.A1(new_n16229_), .A2(new_n16230_), .A3(new_n16226_), .ZN(new_n16234_));
  AOI21_X1   g16134(.A1(new_n16223_), .A2(new_n16215_), .B(new_n16227_), .ZN(new_n16235_));
  NOR3_X1    g16135(.A1(new_n16234_), .A2(new_n16235_), .A3(new_n16233_), .ZN(new_n16236_));
  OAI21_X1   g16136(.A1(new_n16236_), .A2(new_n16232_), .B(new_n16138_), .ZN(new_n16237_));
  INV_X1     g16137(.I(new_n16138_), .ZN(new_n16238_));
  OAI21_X1   g16138(.A1(new_n16234_), .A2(new_n16235_), .B(new_n16233_), .ZN(new_n16239_));
  NAND3_X1   g16139(.A1(new_n16231_), .A2(new_n16228_), .A3(new_n16149_), .ZN(new_n16240_));
  NAND3_X1   g16140(.A1(new_n16239_), .A2(new_n16240_), .A3(new_n16238_), .ZN(new_n16241_));
  NOR2_X1    g16141(.A1(new_n15943_), .A2(new_n16014_), .ZN(new_n16242_));
  INV_X1     g16142(.I(new_n16242_), .ZN(new_n16243_));
  NAND2_X1   g16143(.A1(new_n15943_), .A2(new_n16014_), .ZN(new_n16244_));
  NAND3_X1   g16144(.A1(new_n16016_), .A2(new_n16017_), .A3(new_n15940_), .ZN(new_n16245_));
  OAI21_X1   g16145(.A1(new_n16008_), .A2(new_n16011_), .B(new_n15939_), .ZN(new_n16246_));
  NAND2_X1   g16146(.A1(new_n16246_), .A2(new_n16245_), .ZN(new_n16247_));
  NAND2_X1   g16147(.A1(new_n16247_), .A2(new_n16244_), .ZN(new_n16248_));
  NAND2_X1   g16148(.A1(new_n16248_), .A2(new_n16243_), .ZN(new_n16249_));
  NAND3_X1   g16149(.A1(new_n16237_), .A2(new_n16241_), .A3(new_n16249_), .ZN(new_n16250_));
  AOI21_X1   g16150(.A1(new_n16239_), .A2(new_n16240_), .B(new_n16238_), .ZN(new_n16251_));
  NOR3_X1    g16151(.A1(new_n16236_), .A2(new_n16232_), .A3(new_n16138_), .ZN(new_n16252_));
  AOI22_X1   g16152(.A1(new_n16246_), .A2(new_n16245_), .B1(new_n15943_), .B2(new_n16014_), .ZN(new_n16253_));
  NOR2_X1    g16153(.A1(new_n16253_), .A2(new_n16242_), .ZN(new_n16254_));
  OAI21_X1   g16154(.A1(new_n16252_), .A2(new_n16251_), .B(new_n16254_), .ZN(new_n16255_));
  NAND2_X1   g16155(.A1(new_n16255_), .A2(new_n16250_), .ZN(new_n16256_));
  NAND2_X1   g16156(.A1(new_n16256_), .A2(new_n16135_), .ZN(new_n16257_));
  INV_X1     g16157(.I(new_n16135_), .ZN(new_n16258_));
  NAND3_X1   g16158(.A1(new_n16258_), .A2(new_n16255_), .A3(new_n16250_), .ZN(new_n16259_));
  AOI21_X1   g16159(.A1(new_n16257_), .A2(new_n16259_), .B(new_n16133_), .ZN(new_n16260_));
  AOI21_X1   g16160(.A1(new_n16250_), .A2(new_n16255_), .B(new_n16258_), .ZN(new_n16261_));
  NOR2_X1    g16161(.A1(new_n16256_), .A2(new_n16135_), .ZN(new_n16262_));
  NOR3_X1    g16162(.A1(new_n16262_), .A2(new_n16261_), .A3(new_n16132_), .ZN(new_n16263_));
  AOI22_X1   g16163(.A1(new_n15127_), .A2(new_n7838_), .B1(new_n2469_), .B2(new_n15115_), .ZN(new_n16264_));
  OAI21_X1   g16164(.A1(new_n16264_), .A2(\a[8] ), .B(new_n2469_), .ZN(new_n16265_));
  XNOR2_X1   g16165(.A1(new_n15125_), .A2(new_n16265_), .ZN(new_n16266_));
  NOR3_X1    g16166(.A1(new_n16263_), .A2(new_n16260_), .A3(new_n16266_), .ZN(new_n16267_));
  OAI21_X1   g16167(.A1(new_n16262_), .A2(new_n16261_), .B(new_n16132_), .ZN(new_n16268_));
  NAND3_X1   g16168(.A1(new_n16257_), .A2(new_n16133_), .A3(new_n16259_), .ZN(new_n16269_));
  INV_X1     g16169(.I(new_n16266_), .ZN(new_n16270_));
  AOI21_X1   g16170(.A1(new_n16268_), .A2(new_n16269_), .B(new_n16270_), .ZN(new_n16271_));
  NOR2_X1    g16171(.A1(new_n16267_), .A2(new_n16271_), .ZN(new_n16272_));
  NOR2_X1    g16172(.A1(new_n16272_), .A2(new_n16126_), .ZN(new_n16273_));
  NOR3_X1    g16173(.A1(new_n16267_), .A2(new_n16271_), .A3(new_n16125_), .ZN(new_n16274_));
  OAI21_X1   g16174(.A1(new_n16273_), .A2(new_n16274_), .B(new_n16116_), .ZN(new_n16275_));
  OR3_X2     g16175(.A1(new_n16273_), .A2(new_n16116_), .A3(new_n16274_), .Z(new_n16276_));
  NAND2_X1   g16176(.A1(new_n16276_), .A2(new_n16275_), .ZN(new_n16277_));
  NAND3_X1   g16177(.A1(new_n16050_), .A2(new_n16054_), .A3(new_n15920_), .ZN(new_n16278_));
  OAI21_X1   g16178(.A1(new_n16062_), .A2(new_n16061_), .B(new_n15921_), .ZN(new_n16279_));
  AOI22_X1   g16179(.A1(new_n16279_), .A2(new_n16278_), .B1(new_n16065_), .B2(new_n16058_), .ZN(new_n16280_));
  AOI21_X1   g16180(.A1(new_n15923_), .A2(new_n16059_), .B(new_n16280_), .ZN(new_n16281_));
  NAND2_X1   g16181(.A1(new_n15515_), .A2(new_n5033_), .ZN(new_n16282_));
  NOR2_X1    g16182(.A1(new_n5031_), .A2(new_n2898_), .ZN(new_n16283_));
  AOI21_X1   g16183(.A1(new_n15675_), .A2(new_n16283_), .B(\a[5] ), .ZN(new_n16284_));
  AOI21_X1   g16184(.A1(new_n16284_), .A2(new_n16282_), .B(new_n3040_), .ZN(new_n16285_));
  XNOR2_X1   g16185(.A1(new_n15678_), .A2(new_n16285_), .ZN(new_n16286_));
  XOR2_X1    g16186(.A1(new_n16281_), .A2(new_n16286_), .Z(new_n16287_));
  NAND2_X1   g16187(.A1(new_n16069_), .A2(new_n16072_), .ZN(new_n16288_));
  OAI21_X1   g16188(.A1(new_n16094_), .A2(new_n15916_), .B(new_n16288_), .ZN(new_n16289_));
  NAND2_X1   g16189(.A1(new_n16094_), .A2(new_n15916_), .ZN(new_n16290_));
  NAND2_X1   g16190(.A1(new_n16289_), .A2(new_n16290_), .ZN(new_n16291_));
  XNOR2_X1   g16191(.A1(new_n16291_), .A2(new_n16287_), .ZN(new_n16292_));
  NAND2_X1   g16192(.A1(new_n16292_), .A2(new_n16277_), .ZN(new_n16293_));
  XOR2_X1    g16193(.A1(new_n16291_), .A2(new_n16287_), .Z(new_n16294_));
  NAND3_X1   g16194(.A1(new_n16294_), .A2(new_n16275_), .A3(new_n16276_), .ZN(new_n16295_));
  AND2_X2    g16195(.A1(new_n16295_), .A2(new_n16293_), .Z(new_n16296_));
  XOR2_X1    g16196(.A1(new_n16288_), .A2(new_n15916_), .Z(new_n16297_));
  XOR2_X1    g16197(.A1(new_n16297_), .A2(new_n15906_), .Z(new_n16298_));
  NOR2_X1    g16198(.A1(new_n16298_), .A2(new_n16086_), .ZN(new_n16299_));
  AOI21_X1   g16199(.A1(new_n16293_), .A2(new_n16295_), .B(new_n16299_), .ZN(new_n16300_));
  XOR2_X1    g16200(.A1(new_n16297_), .A2(new_n16094_), .Z(new_n16301_));
  NAND2_X1   g16201(.A1(new_n16301_), .A2(new_n16079_), .ZN(new_n16302_));
  NAND2_X1   g16202(.A1(new_n16113_), .A2(new_n16302_), .ZN(new_n16303_));
  AOI22_X1   g16203(.A1(new_n16303_), .A2(new_n16296_), .B1(new_n16113_), .B2(new_n16300_), .ZN(new_n16304_));
  INV_X1     g16204(.I(new_n16304_), .ZN(new_n16305_));
  OAI21_X1   g16205(.A1(new_n16105_), .A2(new_n16106_), .B(new_n16305_), .ZN(new_n16306_));
  NAND4_X1   g16206(.A1(\result[6] ), .A2(new_n16104_), .A3(new_n16100_), .A4(new_n16304_), .ZN(new_n16307_));
  NAND2_X1   g16207(.A1(new_n16306_), .A2(new_n16307_), .ZN(\result[9] ));
  NAND2_X1   g16208(.A1(new_n15898_), .A2(new_n16100_), .ZN(new_n16309_));
  XOR2_X1    g16209(.A1(new_n16277_), .A2(new_n16287_), .Z(new_n16310_));
  NAND3_X1   g16210(.A1(new_n15894_), .A2(new_n16112_), .A3(new_n16310_), .ZN(new_n16311_));
  AOI21_X1   g16211(.A1(new_n15894_), .A2(new_n16112_), .B(new_n16310_), .ZN(new_n16312_));
  NAND2_X1   g16212(.A1(new_n16299_), .A2(new_n16291_), .ZN(new_n16313_));
  OAI21_X1   g16213(.A1(new_n16312_), .A2(new_n16313_), .B(new_n16311_), .ZN(new_n16314_));
  NAND2_X1   g16214(.A1(new_n16281_), .A2(new_n16286_), .ZN(new_n16315_));
  NOR2_X1    g16215(.A1(new_n16281_), .A2(new_n16286_), .ZN(new_n16316_));
  AOI21_X1   g16216(.A1(new_n16277_), .A2(new_n16315_), .B(new_n16316_), .ZN(new_n16317_));
  INV_X1     g16217(.I(new_n16317_), .ZN(new_n16318_));
  OAI22_X1   g16218(.A1(new_n15313_), .A2(new_n7837_), .B1(new_n2495_), .B2(new_n15305_), .ZN(new_n16319_));
  AOI21_X1   g16219(.A1(new_n16319_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n16320_));
  XNOR2_X1   g16220(.A1(new_n15312_), .A2(new_n16320_), .ZN(new_n16321_));
  NAND2_X1   g16221(.A1(new_n16237_), .A2(new_n16241_), .ZN(new_n16322_));
  NOR2_X1    g16222(.A1(new_n16249_), .A2(new_n16133_), .ZN(new_n16323_));
  NOR2_X1    g16223(.A1(new_n16254_), .A2(new_n16132_), .ZN(new_n16324_));
  OAI21_X1   g16224(.A1(new_n16323_), .A2(new_n16324_), .B(new_n16322_), .ZN(new_n16325_));
  NOR2_X1    g16225(.A1(new_n16252_), .A2(new_n16251_), .ZN(new_n16326_));
  OAI21_X1   g16226(.A1(new_n16253_), .A2(new_n16242_), .B(new_n16132_), .ZN(new_n16327_));
  NAND3_X1   g16227(.A1(new_n16248_), .A2(new_n16133_), .A3(new_n16243_), .ZN(new_n16328_));
  NAND2_X1   g16228(.A1(new_n16328_), .A2(new_n16327_), .ZN(new_n16329_));
  NAND2_X1   g16229(.A1(new_n16326_), .A2(new_n16329_), .ZN(new_n16330_));
  NAND2_X1   g16230(.A1(new_n16325_), .A2(new_n16330_), .ZN(new_n16331_));
  NAND2_X1   g16231(.A1(new_n16135_), .A2(new_n16116_), .ZN(new_n16332_));
  NOR2_X1    g16232(.A1(new_n16135_), .A2(new_n16116_), .ZN(new_n16333_));
  AOI21_X1   g16233(.A1(new_n16331_), .A2(new_n16332_), .B(new_n16333_), .ZN(new_n16334_));
  INV_X1     g16234(.I(new_n16334_), .ZN(new_n16335_));
  AOI22_X1   g16235(.A1(new_n12909_), .A2(new_n5421_), .B1(new_n10949_), .B2(new_n4660_), .ZN(new_n16336_));
  OAI21_X1   g16236(.A1(new_n16336_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n16337_));
  XOR2_X1    g16237(.A1(new_n12907_), .A2(new_n16337_), .Z(new_n16338_));
  NOR2_X1    g16238(.A1(new_n16233_), .A2(new_n16226_), .ZN(new_n16339_));
  NAND3_X1   g16239(.A1(new_n16223_), .A2(new_n16215_), .A3(new_n16238_), .ZN(new_n16340_));
  OAI21_X1   g16240(.A1(new_n16229_), .A2(new_n16230_), .B(new_n16138_), .ZN(new_n16341_));
  AOI22_X1   g16241(.A1(new_n16341_), .A2(new_n16340_), .B1(new_n16233_), .B2(new_n16226_), .ZN(new_n16342_));
  NOR2_X1    g16242(.A1(new_n16342_), .A2(new_n16339_), .ZN(new_n16343_));
  INV_X1     g16243(.I(new_n16343_), .ZN(new_n16344_));
  OAI22_X1   g16244(.A1(new_n12601_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n10595_), .ZN(new_n16345_));
  AOI21_X1   g16245(.A1(new_n16345_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n16346_));
  XOR2_X1    g16246(.A1(new_n12600_), .A2(new_n16346_), .Z(new_n16347_));
  OAI21_X1   g16247(.A1(new_n16190_), .A2(new_n16187_), .B(new_n16216_), .ZN(new_n16348_));
  NAND2_X1   g16248(.A1(new_n16348_), .A2(new_n16217_), .ZN(new_n16349_));
  OAI22_X1   g16249(.A1(new_n10870_), .A2(new_n4529_), .B1(new_n4527_), .B2(new_n10868_), .ZN(new_n16350_));
  OAI21_X1   g16250(.A1(new_n79_), .A2(new_n10881_), .B(new_n16350_), .ZN(new_n16351_));
  AOI21_X1   g16251(.A1(new_n16351_), .A2(new_n72_), .B(new_n79_), .ZN(new_n16352_));
  XNOR2_X1   g16252(.A1(new_n11802_), .A2(new_n16352_), .ZN(new_n16353_));
  NOR2_X1    g16253(.A1(new_n16177_), .A2(new_n16153_), .ZN(new_n16354_));
  INV_X1     g16254(.I(new_n16354_), .ZN(new_n16355_));
  NAND2_X1   g16255(.A1(new_n16177_), .A2(new_n16153_), .ZN(new_n16356_));
  AOI21_X1   g16256(.A1(new_n16157_), .A2(new_n16158_), .B(new_n16182_), .ZN(new_n16357_));
  AOI21_X1   g16257(.A1(new_n15960_), .A2(new_n15968_), .B(new_n16155_), .ZN(new_n16358_));
  NOR2_X1    g16258(.A1(new_n15960_), .A2(new_n15968_), .ZN(new_n16359_));
  NOR3_X1    g16259(.A1(new_n16173_), .A2(new_n16358_), .A3(new_n16359_), .ZN(new_n16360_));
  OAI21_X1   g16260(.A1(new_n16357_), .A2(new_n16360_), .B(new_n16356_), .ZN(new_n16361_));
  NAND2_X1   g16261(.A1(new_n16361_), .A2(new_n16355_), .ZN(new_n16362_));
  NOR3_X1    g16262(.A1(new_n15967_), .A2(new_n15762_), .A3(new_n16165_), .ZN(new_n16363_));
  NOR3_X1    g16263(.A1(new_n16358_), .A2(new_n16182_), .A3(new_n16359_), .ZN(new_n16364_));
  NOR2_X1    g16264(.A1(new_n15967_), .A2(new_n15761_), .ZN(new_n16365_));
  INV_X1     g16265(.I(new_n16365_), .ZN(new_n16366_));
  INV_X1     g16266(.I(new_n5035_), .ZN(new_n16367_));
  NOR2_X1    g16267(.A1(new_n15515_), .A2(new_n5034_), .ZN(new_n16368_));
  OAI22_X1   g16268(.A1(new_n16368_), .A2(\a[5] ), .B1(new_n16367_), .B2(new_n15515_), .ZN(new_n16369_));
  NOR2_X1    g16269(.A1(new_n16369_), .A2(new_n15967_), .ZN(new_n16370_));
  NAND2_X1   g16270(.A1(new_n15511_), .A2(new_n5036_), .ZN(new_n16371_));
  AOI22_X1   g16271(.A1(new_n16371_), .A2(new_n452_), .B1(new_n5035_), .B2(new_n15511_), .ZN(new_n16372_));
  NOR2_X1    g16272(.A1(new_n16372_), .A2(new_n15961_), .ZN(new_n16373_));
  AOI22_X1   g16273(.A1(new_n10857_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n10630_), .ZN(new_n16374_));
  OAI21_X1   g16274(.A1(new_n88_), .A2(new_n10844_), .B(new_n16374_), .ZN(new_n16375_));
  NAND3_X1   g16275(.A1(new_n13210_), .A2(new_n961_), .A3(new_n16375_), .ZN(new_n16376_));
  OAI21_X1   g16276(.A1(new_n16370_), .A2(new_n16373_), .B(new_n16376_), .ZN(new_n16377_));
  NAND2_X1   g16277(.A1(new_n16372_), .A2(new_n15961_), .ZN(new_n16378_));
  NAND2_X1   g16278(.A1(new_n16369_), .A2(new_n15967_), .ZN(new_n16379_));
  INV_X1     g16279(.I(new_n16376_), .ZN(new_n16380_));
  NAND3_X1   g16280(.A1(new_n16379_), .A2(new_n16378_), .A3(new_n16380_), .ZN(new_n16381_));
  AOI21_X1   g16281(.A1(new_n16377_), .A2(new_n16381_), .B(new_n16366_), .ZN(new_n16382_));
  NAND3_X1   g16282(.A1(new_n16379_), .A2(new_n16378_), .A3(new_n16376_), .ZN(new_n16383_));
  OAI21_X1   g16283(.A1(new_n16370_), .A2(new_n16373_), .B(new_n16380_), .ZN(new_n16384_));
  AOI21_X1   g16284(.A1(new_n16384_), .A2(new_n16383_), .B(new_n16365_), .ZN(new_n16385_));
  NOR2_X1    g16285(.A1(new_n16382_), .A2(new_n16385_), .ZN(new_n16386_));
  OAI21_X1   g16286(.A1(new_n16363_), .A2(new_n16364_), .B(new_n16386_), .ZN(new_n16387_));
  INV_X1     g16287(.I(new_n16363_), .ZN(new_n16388_));
  NAND3_X1   g16288(.A1(new_n16157_), .A2(new_n16173_), .A3(new_n16158_), .ZN(new_n16389_));
  AOI21_X1   g16289(.A1(new_n16379_), .A2(new_n16378_), .B(new_n16380_), .ZN(new_n16390_));
  NOR3_X1    g16290(.A1(new_n16370_), .A2(new_n16373_), .A3(new_n16376_), .ZN(new_n16391_));
  OAI21_X1   g16291(.A1(new_n16390_), .A2(new_n16391_), .B(new_n16365_), .ZN(new_n16392_));
  NOR3_X1    g16292(.A1(new_n16370_), .A2(new_n16373_), .A3(new_n16380_), .ZN(new_n16393_));
  AOI21_X1   g16293(.A1(new_n16379_), .A2(new_n16378_), .B(new_n16376_), .ZN(new_n16394_));
  OAI21_X1   g16294(.A1(new_n16394_), .A2(new_n16393_), .B(new_n16366_), .ZN(new_n16395_));
  NAND2_X1   g16295(.A1(new_n16392_), .A2(new_n16395_), .ZN(new_n16396_));
  NAND3_X1   g16296(.A1(new_n16396_), .A2(new_n16389_), .A3(new_n16388_), .ZN(new_n16397_));
  OAI22_X1   g16297(.A1(new_n10619_), .A2(new_n4612_), .B1(new_n4781_), .B2(new_n10611_), .ZN(new_n16398_));
  OAI21_X1   g16298(.A1(new_n1128_), .A2(new_n10896_), .B(new_n16398_), .ZN(new_n16399_));
  AOI21_X1   g16299(.A1(new_n16399_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n16400_));
  XNOR2_X1   g16300(.A1(new_n10984_), .A2(new_n16400_), .ZN(new_n16401_));
  INV_X1     g16301(.I(new_n16401_), .ZN(new_n16402_));
  NAND3_X1   g16302(.A1(new_n16387_), .A2(new_n16397_), .A3(new_n16402_), .ZN(new_n16403_));
  AOI21_X1   g16303(.A1(new_n16388_), .A2(new_n16389_), .B(new_n16396_), .ZN(new_n16404_));
  NOR3_X1    g16304(.A1(new_n16386_), .A2(new_n16364_), .A3(new_n16363_), .ZN(new_n16405_));
  OAI21_X1   g16305(.A1(new_n16404_), .A2(new_n16405_), .B(new_n16401_), .ZN(new_n16406_));
  AOI21_X1   g16306(.A1(new_n16406_), .A2(new_n16403_), .B(new_n16362_), .ZN(new_n16407_));
  OR2_X2     g16307(.A1(new_n16357_), .A2(new_n16360_), .Z(new_n16408_));
  AOI21_X1   g16308(.A1(new_n16408_), .A2(new_n16356_), .B(new_n16354_), .ZN(new_n16409_));
  NOR3_X1    g16309(.A1(new_n16404_), .A2(new_n16405_), .A3(new_n16401_), .ZN(new_n16410_));
  AOI21_X1   g16310(.A1(new_n16387_), .A2(new_n16397_), .B(new_n16402_), .ZN(new_n16411_));
  NOR3_X1    g16311(.A1(new_n16409_), .A2(new_n16410_), .A3(new_n16411_), .ZN(new_n16412_));
  OAI21_X1   g16312(.A1(new_n16412_), .A2(new_n16407_), .B(new_n16353_), .ZN(new_n16413_));
  INV_X1     g16313(.I(new_n16353_), .ZN(new_n16414_));
  OAI21_X1   g16314(.A1(new_n16410_), .A2(new_n16411_), .B(new_n16409_), .ZN(new_n16415_));
  NAND3_X1   g16315(.A1(new_n16406_), .A2(new_n16403_), .A3(new_n16362_), .ZN(new_n16416_));
  NAND3_X1   g16316(.A1(new_n16415_), .A2(new_n16414_), .A3(new_n16416_), .ZN(new_n16417_));
  AOI22_X1   g16317(.A1(new_n12891_), .A2(new_n5337_), .B1(new_n10924_), .B2(new_n4717_), .ZN(new_n16418_));
  OAI21_X1   g16318(.A1(new_n16418_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n16419_));
  XNOR2_X1   g16319(.A1(new_n12889_), .A2(new_n16419_), .ZN(new_n16420_));
  INV_X1     g16320(.I(new_n16420_), .ZN(new_n16421_));
  NAND3_X1   g16321(.A1(new_n16417_), .A2(new_n16413_), .A3(new_n16421_), .ZN(new_n16422_));
  AOI21_X1   g16322(.A1(new_n16415_), .A2(new_n16416_), .B(new_n16414_), .ZN(new_n16423_));
  NOR3_X1    g16323(.A1(new_n16412_), .A2(new_n16407_), .A3(new_n16353_), .ZN(new_n16424_));
  OAI21_X1   g16324(.A1(new_n16423_), .A2(new_n16424_), .B(new_n16420_), .ZN(new_n16425_));
  AOI21_X1   g16325(.A1(new_n16425_), .A2(new_n16422_), .B(new_n16349_), .ZN(new_n16426_));
  NAND2_X1   g16326(.A1(new_n16206_), .A2(new_n16207_), .ZN(new_n16427_));
  AOI21_X1   g16327(.A1(new_n16427_), .A2(new_n16216_), .B(new_n16204_), .ZN(new_n16428_));
  NOR3_X1    g16328(.A1(new_n16423_), .A2(new_n16424_), .A3(new_n16420_), .ZN(new_n16429_));
  AOI21_X1   g16329(.A1(new_n16417_), .A2(new_n16413_), .B(new_n16421_), .ZN(new_n16430_));
  NOR3_X1    g16330(.A1(new_n16429_), .A2(new_n16430_), .A3(new_n16428_), .ZN(new_n16431_));
  OAI21_X1   g16331(.A1(new_n16431_), .A2(new_n16426_), .B(new_n16347_), .ZN(new_n16432_));
  INV_X1     g16332(.I(new_n16347_), .ZN(new_n16433_));
  OAI21_X1   g16333(.A1(new_n16429_), .A2(new_n16430_), .B(new_n16428_), .ZN(new_n16434_));
  NAND3_X1   g16334(.A1(new_n16425_), .A2(new_n16422_), .A3(new_n16349_), .ZN(new_n16435_));
  NAND3_X1   g16335(.A1(new_n16434_), .A2(new_n16435_), .A3(new_n16433_), .ZN(new_n16436_));
  OAI22_X1   g16336(.A1(new_n16218_), .A2(new_n16221_), .B1(new_n16238_), .B2(new_n16214_), .ZN(new_n16437_));
  NAND2_X1   g16337(.A1(new_n16214_), .A2(new_n16238_), .ZN(new_n16438_));
  NAND2_X1   g16338(.A1(new_n16437_), .A2(new_n16438_), .ZN(new_n16439_));
  NAND3_X1   g16339(.A1(new_n16432_), .A2(new_n16436_), .A3(new_n16439_), .ZN(new_n16440_));
  AOI21_X1   g16340(.A1(new_n16434_), .A2(new_n16435_), .B(new_n16433_), .ZN(new_n16441_));
  NOR3_X1    g16341(.A1(new_n16431_), .A2(new_n16426_), .A3(new_n16347_), .ZN(new_n16442_));
  INV_X1     g16342(.I(new_n16439_), .ZN(new_n16443_));
  OAI21_X1   g16343(.A1(new_n16442_), .A2(new_n16441_), .B(new_n16443_), .ZN(new_n16444_));
  AOI21_X1   g16344(.A1(new_n16444_), .A2(new_n16440_), .B(new_n16344_), .ZN(new_n16445_));
  NOR3_X1    g16345(.A1(new_n16442_), .A2(new_n16441_), .A3(new_n16443_), .ZN(new_n16446_));
  AOI21_X1   g16346(.A1(new_n16432_), .A2(new_n16436_), .B(new_n16439_), .ZN(new_n16447_));
  NOR3_X1    g16347(.A1(new_n16446_), .A2(new_n16447_), .A3(new_n16343_), .ZN(new_n16448_));
  OAI21_X1   g16348(.A1(new_n16448_), .A2(new_n16445_), .B(new_n16338_), .ZN(new_n16449_));
  INV_X1     g16349(.I(new_n16338_), .ZN(new_n16450_));
  OAI21_X1   g16350(.A1(new_n16446_), .A2(new_n16447_), .B(new_n16343_), .ZN(new_n16451_));
  NAND3_X1   g16351(.A1(new_n16444_), .A2(new_n16440_), .A3(new_n16344_), .ZN(new_n16452_));
  NAND3_X1   g16352(.A1(new_n16451_), .A2(new_n16452_), .A3(new_n16450_), .ZN(new_n16453_));
  INV_X1     g16353(.I(new_n16327_), .ZN(new_n16454_));
  NOR3_X1    g16354(.A1(new_n16253_), .A2(new_n16132_), .A3(new_n16242_), .ZN(new_n16455_));
  OAI22_X1   g16355(.A1(new_n10965_), .A2(new_n5967_), .B1(new_n643_), .B2(new_n10570_), .ZN(new_n16456_));
  AOI21_X1   g16356(.A1(new_n16456_), .A2(new_n279_), .B(new_n643_), .ZN(new_n16457_));
  XNOR2_X1   g16357(.A1(new_n14077_), .A2(new_n16457_), .ZN(new_n16458_));
  INV_X1     g16358(.I(new_n16458_), .ZN(new_n16459_));
  OAI21_X1   g16359(.A1(new_n16454_), .A2(new_n16455_), .B(new_n16459_), .ZN(new_n16460_));
  NOR2_X1    g16360(.A1(new_n16460_), .A2(new_n16324_), .ZN(new_n16461_));
  NOR2_X1    g16361(.A1(new_n16254_), .A2(new_n16132_), .ZN(new_n16462_));
  OAI21_X1   g16362(.A1(new_n16461_), .A2(new_n16462_), .B(new_n16326_), .ZN(new_n16463_));
  NAND2_X1   g16363(.A1(new_n16249_), .A2(new_n16133_), .ZN(new_n16464_));
  NAND3_X1   g16364(.A1(new_n16329_), .A2(new_n16464_), .A3(new_n16459_), .ZN(new_n16465_));
  INV_X1     g16365(.I(new_n16462_), .ZN(new_n16466_));
  NAND3_X1   g16366(.A1(new_n16465_), .A2(new_n16322_), .A3(new_n16466_), .ZN(new_n16467_));
  NAND2_X1   g16367(.A1(new_n16463_), .A2(new_n16467_), .ZN(new_n16468_));
  AOI22_X1   g16368(.A1(new_n14602_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n14603_), .ZN(new_n16469_));
  OAI21_X1   g16369(.A1(new_n16469_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n16470_));
  XNOR2_X1   g16370(.A1(new_n14601_), .A2(new_n16470_), .ZN(new_n16471_));
  NAND2_X1   g16371(.A1(new_n16468_), .A2(new_n16471_), .ZN(new_n16472_));
  INV_X1     g16372(.I(new_n16471_), .ZN(new_n16473_));
  NAND3_X1   g16373(.A1(new_n16463_), .A2(new_n16467_), .A3(new_n16473_), .ZN(new_n16474_));
  AOI22_X1   g16374(.A1(new_n16472_), .A2(new_n16474_), .B1(new_n16449_), .B2(new_n16453_), .ZN(new_n16475_));
  NAND2_X1   g16375(.A1(new_n16449_), .A2(new_n16453_), .ZN(new_n16476_));
  NAND3_X1   g16376(.A1(new_n16463_), .A2(new_n16467_), .A3(new_n16471_), .ZN(new_n16477_));
  AOI21_X1   g16377(.A1(new_n16465_), .A2(new_n16466_), .B(new_n16322_), .ZN(new_n16478_));
  NOR3_X1    g16378(.A1(new_n16461_), .A2(new_n16326_), .A3(new_n16462_), .ZN(new_n16479_));
  OAI21_X1   g16379(.A1(new_n16479_), .A2(new_n16478_), .B(new_n16473_), .ZN(new_n16480_));
  AOI21_X1   g16380(.A1(new_n16477_), .A2(new_n16480_), .B(new_n16476_), .ZN(new_n16481_));
  NOR2_X1    g16381(.A1(new_n16481_), .A2(new_n16475_), .ZN(new_n16482_));
  NOR2_X1    g16382(.A1(new_n16125_), .A2(new_n16266_), .ZN(new_n16483_));
  INV_X1     g16383(.I(new_n16483_), .ZN(new_n16484_));
  NOR3_X1    g16384(.A1(new_n16263_), .A2(new_n16260_), .A3(new_n16116_), .ZN(new_n16485_));
  INV_X1     g16385(.I(new_n16116_), .ZN(new_n16486_));
  AOI21_X1   g16386(.A1(new_n16268_), .A2(new_n16269_), .B(new_n16486_), .ZN(new_n16487_));
  OAI22_X1   g16387(.A1(new_n16485_), .A2(new_n16487_), .B1(new_n16126_), .B2(new_n16270_), .ZN(new_n16488_));
  NAND2_X1   g16388(.A1(new_n16488_), .A2(new_n16484_), .ZN(new_n16489_));
  NAND2_X1   g16389(.A1(new_n16489_), .A2(new_n16482_), .ZN(new_n16490_));
  NOR2_X1    g16390(.A1(new_n16489_), .A2(new_n16482_), .ZN(new_n16491_));
  INV_X1     g16391(.I(new_n16491_), .ZN(new_n16492_));
  AOI21_X1   g16392(.A1(new_n16492_), .A2(new_n16490_), .B(new_n16335_), .ZN(new_n16493_));
  INV_X1     g16393(.I(new_n16490_), .ZN(new_n16494_));
  NOR3_X1    g16394(.A1(new_n16494_), .A2(new_n16334_), .A3(new_n16491_), .ZN(new_n16495_));
  OAI21_X1   g16395(.A1(new_n16493_), .A2(new_n16495_), .B(new_n16321_), .ZN(new_n16496_));
  INV_X1     g16396(.I(new_n16321_), .ZN(new_n16497_));
  OAI21_X1   g16397(.A1(new_n16494_), .A2(new_n16491_), .B(new_n16334_), .ZN(new_n16498_));
  NAND3_X1   g16398(.A1(new_n16492_), .A2(new_n16335_), .A3(new_n16490_), .ZN(new_n16499_));
  NAND3_X1   g16399(.A1(new_n16498_), .A2(new_n16499_), .A3(new_n16497_), .ZN(new_n16500_));
  NAND2_X1   g16400(.A1(new_n16496_), .A2(new_n16500_), .ZN(new_n16501_));
  NOR2_X1    g16401(.A1(new_n16501_), .A2(new_n16318_), .ZN(new_n16502_));
  AOI21_X1   g16402(.A1(new_n16498_), .A2(new_n16499_), .B(new_n16497_), .ZN(new_n16503_));
  NOR3_X1    g16403(.A1(new_n16493_), .A2(new_n16495_), .A3(new_n16321_), .ZN(new_n16504_));
  NOR2_X1    g16404(.A1(new_n16503_), .A2(new_n16504_), .ZN(new_n16505_));
  NOR2_X1    g16405(.A1(new_n16505_), .A2(new_n16317_), .ZN(new_n16506_));
  OAI21_X1   g16406(.A1(new_n16502_), .A2(new_n16506_), .B(new_n16314_), .ZN(new_n16507_));
  XOR2_X1    g16407(.A1(new_n16309_), .A2(new_n16507_), .Z(new_n16508_));
  XOR2_X1    g16408(.A1(new_n16508_), .A2(new_n16305_), .Z(\result[10] ));
  AOI21_X1   g16409(.A1(new_n16306_), .A2(new_n16307_), .B(new_n16507_), .ZN(new_n16510_));
  NAND3_X1   g16410(.A1(new_n16093_), .A2(new_n16097_), .A3(new_n15883_), .ZN(new_n16511_));
  AOI21_X1   g16411(.A1(new_n16093_), .A2(new_n16097_), .B(new_n15883_), .ZN(new_n16512_));
  OAI21_X1   g16412(.A1(new_n15886_), .A2(new_n16512_), .B(new_n16511_), .ZN(new_n16513_));
  XNOR2_X1   g16413(.A1(new_n16277_), .A2(new_n16287_), .ZN(new_n16514_));
  NOR3_X1    g16414(.A1(new_n15901_), .A2(new_n16513_), .A3(new_n16514_), .ZN(new_n16515_));
  OAI21_X1   g16415(.A1(new_n15901_), .A2(new_n16513_), .B(new_n16514_), .ZN(new_n16516_));
  AOI21_X1   g16416(.A1(new_n16289_), .A2(new_n16290_), .B(new_n16302_), .ZN(new_n16517_));
  AOI21_X1   g16417(.A1(new_n16516_), .A2(new_n16517_), .B(new_n16515_), .ZN(new_n16518_));
  OAI22_X1   g16418(.A1(new_n15305_), .A2(new_n7836_), .B1(new_n15114_), .B2(new_n2718_), .ZN(new_n16519_));
  OAI21_X1   g16419(.A1(new_n2495_), .A2(new_n15515_), .B(new_n16519_), .ZN(new_n16520_));
  AOI21_X1   g16420(.A1(new_n16520_), .A2(new_n498_), .B(new_n2495_), .ZN(new_n16521_));
  XOR2_X1    g16421(.A1(new_n15518_), .A2(new_n16521_), .Z(new_n16522_));
  INV_X1     g16422(.I(new_n16522_), .ZN(new_n16523_));
  NAND2_X1   g16423(.A1(new_n16335_), .A2(new_n16473_), .ZN(new_n16524_));
  XOR2_X1    g16424(.A1(new_n16476_), .A2(new_n16468_), .Z(new_n16525_));
  OAI21_X1   g16425(.A1(new_n16335_), .A2(new_n16473_), .B(new_n16525_), .ZN(new_n16526_));
  NAND2_X1   g16426(.A1(new_n16526_), .A2(new_n16524_), .ZN(new_n16527_));
  INV_X1     g16427(.I(new_n16527_), .ZN(new_n16528_));
  OAI22_X1   g16428(.A1(new_n10570_), .A2(new_n5966_), .B1(new_n1851_), .B2(new_n10961_), .ZN(new_n16529_));
  OAI21_X1   g16429(.A1(new_n10564_), .A2(new_n643_), .B(new_n16529_), .ZN(new_n16530_));
  AOI21_X1   g16430(.A1(new_n16530_), .A2(new_n279_), .B(new_n643_), .ZN(new_n16531_));
  XOR2_X1    g16431(.A1(new_n10976_), .A2(new_n16531_), .Z(new_n16532_));
  INV_X1     g16432(.I(new_n16532_), .ZN(new_n16533_));
  OAI21_X1   g16433(.A1(new_n16326_), .A2(new_n16323_), .B(new_n16464_), .ZN(new_n16534_));
  NAND2_X1   g16434(.A1(new_n16534_), .A2(new_n16459_), .ZN(new_n16535_));
  NOR2_X1    g16435(.A1(new_n16534_), .A2(new_n16459_), .ZN(new_n16536_));
  OAI21_X1   g16436(.A1(new_n16476_), .A2(new_n16536_), .B(new_n16535_), .ZN(new_n16537_));
  INV_X1     g16437(.I(new_n16537_), .ZN(new_n16538_));
  OAI22_X1   g16438(.A1(new_n1622_), .A2(new_n10938_), .B1(new_n10952_), .B2(new_n5419_), .ZN(new_n16539_));
  OAI21_X1   g16439(.A1(new_n10577_), .A2(new_n1620_), .B(new_n16539_), .ZN(new_n16540_));
  AOI21_X1   g16440(.A1(new_n16540_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n16541_));
  XOR2_X1    g16441(.A1(new_n13544_), .A2(new_n16541_), .Z(new_n16542_));
  INV_X1     g16442(.I(new_n16542_), .ZN(new_n16543_));
  NOR2_X1    g16443(.A1(new_n16423_), .A2(new_n16424_), .ZN(new_n16544_));
  XOR2_X1    g16444(.A1(new_n16428_), .A2(new_n16347_), .Z(new_n16545_));
  NAND2_X1   g16445(.A1(new_n16545_), .A2(new_n16544_), .ZN(new_n16546_));
  NAND2_X1   g16446(.A1(new_n16417_), .A2(new_n16413_), .ZN(new_n16547_));
  NAND2_X1   g16447(.A1(new_n16428_), .A2(new_n16347_), .ZN(new_n16548_));
  NAND2_X1   g16448(.A1(new_n16349_), .A2(new_n16433_), .ZN(new_n16549_));
  NAND2_X1   g16449(.A1(new_n16549_), .A2(new_n16548_), .ZN(new_n16550_));
  AOI22_X1   g16450(.A1(new_n16443_), .A2(new_n16420_), .B1(new_n16550_), .B2(new_n16547_), .ZN(new_n16551_));
  AOI22_X1   g16451(.A1(new_n16551_), .A2(new_n16546_), .B1(new_n16421_), .B2(new_n16439_), .ZN(new_n16552_));
  OAI22_X1   g16452(.A1(new_n10896_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10611_), .ZN(new_n16553_));
  OAI21_X1   g16453(.A1(new_n10606_), .A2(new_n1128_), .B(new_n16553_), .ZN(new_n16554_));
  AOI21_X1   g16454(.A1(new_n16554_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n16555_));
  XOR2_X1    g16455(.A1(new_n12211_), .A2(new_n16555_), .Z(new_n16556_));
  INV_X1     g16456(.I(new_n16556_), .ZN(new_n16557_));
  NOR2_X1    g16457(.A1(new_n16409_), .A2(new_n16401_), .ZN(new_n16558_));
  NAND2_X1   g16458(.A1(new_n16409_), .A2(new_n16401_), .ZN(new_n16559_));
  NAND3_X1   g16459(.A1(new_n16387_), .A2(new_n16397_), .A3(new_n16414_), .ZN(new_n16560_));
  OAI21_X1   g16460(.A1(new_n16404_), .A2(new_n16405_), .B(new_n16353_), .ZN(new_n16561_));
  NAND2_X1   g16461(.A1(new_n16561_), .A2(new_n16560_), .ZN(new_n16562_));
  AOI21_X1   g16462(.A1(new_n16562_), .A2(new_n16559_), .B(new_n16558_), .ZN(new_n16563_));
  NAND2_X1   g16463(.A1(new_n16396_), .A2(new_n16353_), .ZN(new_n16564_));
  NAND3_X1   g16464(.A1(new_n16564_), .A2(new_n16388_), .A3(new_n16389_), .ZN(new_n16565_));
  NOR2_X1    g16465(.A1(new_n16396_), .A2(new_n16353_), .ZN(new_n16566_));
  INV_X1     g16466(.I(new_n16566_), .ZN(new_n16567_));
  AOI21_X1   g16467(.A1(new_n16365_), .A2(new_n16383_), .B(new_n16394_), .ZN(new_n16568_));
  NOR2_X1    g16468(.A1(new_n16369_), .A2(new_n15961_), .ZN(new_n16569_));
  NOR2_X1    g16469(.A1(new_n10870_), .A2(new_n511_), .ZN(new_n16570_));
  INV_X1     g16470(.I(new_n16570_), .ZN(new_n16571_));
  AOI22_X1   g16471(.A1(new_n10857_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n10843_), .ZN(new_n16572_));
  AOI21_X1   g16472(.A1(new_n16571_), .A2(new_n16572_), .B(new_n82_), .ZN(new_n16573_));
  NAND2_X1   g16473(.A1(new_n13225_), .A2(new_n16573_), .ZN(new_n16574_));
  INV_X1     g16474(.I(new_n16574_), .ZN(new_n16575_));
  NAND2_X1   g16475(.A1(new_n16569_), .A2(new_n16575_), .ZN(new_n16576_));
  INV_X1     g16476(.I(new_n16576_), .ZN(new_n16577_));
  OAI21_X1   g16477(.A1(new_n16369_), .A2(new_n15961_), .B(new_n16574_), .ZN(new_n16578_));
  INV_X1     g16478(.I(new_n16578_), .ZN(new_n16579_));
  OAI22_X1   g16479(.A1(new_n10881_), .A2(new_n4527_), .B1(new_n10868_), .B2(new_n4529_), .ZN(new_n16580_));
  OAI21_X1   g16480(.A1(new_n10619_), .A2(new_n79_), .B(new_n16580_), .ZN(new_n16581_));
  AOI21_X1   g16481(.A1(new_n16581_), .A2(new_n72_), .B(new_n79_), .ZN(new_n16582_));
  XOR2_X1    g16482(.A1(new_n12074_), .A2(new_n16582_), .Z(new_n16583_));
  OAI21_X1   g16483(.A1(new_n16577_), .A2(new_n16579_), .B(new_n16583_), .ZN(new_n16584_));
  INV_X1     g16484(.I(new_n16583_), .ZN(new_n16585_));
  NAND3_X1   g16485(.A1(new_n16576_), .A2(new_n16578_), .A3(new_n16585_), .ZN(new_n16586_));
  AOI21_X1   g16486(.A1(new_n16584_), .A2(new_n16586_), .B(new_n16568_), .ZN(new_n16587_));
  OAI21_X1   g16487(.A1(new_n16366_), .A2(new_n16393_), .B(new_n16384_), .ZN(new_n16588_));
  NAND3_X1   g16488(.A1(new_n16576_), .A2(new_n16578_), .A3(new_n16583_), .ZN(new_n16589_));
  OAI21_X1   g16489(.A1(new_n16577_), .A2(new_n16579_), .B(new_n16585_), .ZN(new_n16590_));
  AOI21_X1   g16490(.A1(new_n16590_), .A2(new_n16589_), .B(new_n16588_), .ZN(new_n16591_));
  NOR2_X1    g16491(.A1(new_n16587_), .A2(new_n16591_), .ZN(new_n16592_));
  NAND3_X1   g16492(.A1(new_n16565_), .A2(new_n16592_), .A3(new_n16567_), .ZN(new_n16593_));
  NOR2_X1    g16493(.A1(new_n16386_), .A2(new_n16414_), .ZN(new_n16594_));
  NOR3_X1    g16494(.A1(new_n16594_), .A2(new_n16363_), .A3(new_n16364_), .ZN(new_n16595_));
  INV_X1     g16495(.I(new_n16592_), .ZN(new_n16596_));
  OAI21_X1   g16496(.A1(new_n16595_), .A2(new_n16566_), .B(new_n16596_), .ZN(new_n16597_));
  OAI22_X1   g16497(.A1(new_n10589_), .A2(new_n1239_), .B1(new_n12623_), .B2(new_n4981_), .ZN(new_n16598_));
  AOI21_X1   g16498(.A1(new_n16598_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n16599_));
  XOR2_X1    g16499(.A1(new_n12622_), .A2(new_n16599_), .Z(new_n16600_));
  INV_X1     g16500(.I(new_n16600_), .ZN(new_n16601_));
  NAND3_X1   g16501(.A1(new_n16597_), .A2(new_n16593_), .A3(new_n16601_), .ZN(new_n16602_));
  NOR3_X1    g16502(.A1(new_n16596_), .A2(new_n16595_), .A3(new_n16566_), .ZN(new_n16603_));
  AOI21_X1   g16503(.A1(new_n16565_), .A2(new_n16567_), .B(new_n16592_), .ZN(new_n16604_));
  OAI21_X1   g16504(.A1(new_n16603_), .A2(new_n16604_), .B(new_n16600_), .ZN(new_n16605_));
  NAND2_X1   g16505(.A1(new_n16602_), .A2(new_n16605_), .ZN(new_n16606_));
  NAND2_X1   g16506(.A1(new_n16606_), .A2(new_n16563_), .ZN(new_n16607_));
  INV_X1     g16507(.I(new_n16563_), .ZN(new_n16608_));
  NOR3_X1    g16508(.A1(new_n16603_), .A2(new_n16604_), .A3(new_n16600_), .ZN(new_n16609_));
  AOI21_X1   g16509(.A1(new_n16597_), .A2(new_n16593_), .B(new_n16601_), .ZN(new_n16610_));
  NOR2_X1    g16510(.A1(new_n16610_), .A2(new_n16609_), .ZN(new_n16611_));
  NAND2_X1   g16511(.A1(new_n16608_), .A2(new_n16611_), .ZN(new_n16612_));
  AOI21_X1   g16512(.A1(new_n16612_), .A2(new_n16607_), .B(new_n16557_), .ZN(new_n16613_));
  NOR2_X1    g16513(.A1(new_n16608_), .A2(new_n16611_), .ZN(new_n16614_));
  NOR2_X1    g16514(.A1(new_n16606_), .A2(new_n16563_), .ZN(new_n16615_));
  NOR3_X1    g16515(.A1(new_n16614_), .A2(new_n16615_), .A3(new_n16556_), .ZN(new_n16616_));
  INV_X1     g16516(.I(new_n16549_), .ZN(new_n16617_));
  NOR2_X1    g16517(.A1(new_n16349_), .A2(new_n16433_), .ZN(new_n16618_));
  NOR2_X1    g16518(.A1(new_n16547_), .A2(new_n16618_), .ZN(new_n16619_));
  OAI22_X1   g16519(.A1(new_n10583_), .A2(new_n5398_), .B1(new_n5336_), .B2(new_n10928_), .ZN(new_n16620_));
  AOI21_X1   g16520(.A1(new_n16620_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n16621_));
  XNOR2_X1   g16521(.A1(new_n13378_), .A2(new_n16621_), .ZN(new_n16622_));
  INV_X1     g16522(.I(new_n16622_), .ZN(new_n16623_));
  NOR3_X1    g16523(.A1(new_n16619_), .A2(new_n16617_), .A3(new_n16623_), .ZN(new_n16624_));
  NAND2_X1   g16524(.A1(new_n16544_), .A2(new_n16548_), .ZN(new_n16625_));
  AOI21_X1   g16525(.A1(new_n16625_), .A2(new_n16549_), .B(new_n16622_), .ZN(new_n16626_));
  OAI22_X1   g16526(.A1(new_n16626_), .A2(new_n16624_), .B1(new_n16613_), .B2(new_n16616_), .ZN(new_n16627_));
  NOR2_X1    g16527(.A1(new_n16616_), .A2(new_n16613_), .ZN(new_n16628_));
  OAI21_X1   g16528(.A1(new_n16619_), .A2(new_n16617_), .B(new_n16622_), .ZN(new_n16629_));
  NAND3_X1   g16529(.A1(new_n16625_), .A2(new_n16549_), .A3(new_n16623_), .ZN(new_n16630_));
  NAND2_X1   g16530(.A1(new_n16630_), .A2(new_n16629_), .ZN(new_n16631_));
  NAND2_X1   g16531(.A1(new_n16631_), .A2(new_n16628_), .ZN(new_n16632_));
  NAND2_X1   g16532(.A1(new_n16632_), .A2(new_n16627_), .ZN(new_n16633_));
  NOR2_X1    g16533(.A1(new_n16343_), .A2(new_n16338_), .ZN(new_n16634_));
  INV_X1     g16534(.I(new_n16634_), .ZN(new_n16635_));
  NOR3_X1    g16535(.A1(new_n16342_), .A2(new_n16450_), .A3(new_n16339_), .ZN(new_n16636_));
  INV_X1     g16536(.I(new_n16636_), .ZN(new_n16637_));
  OAI21_X1   g16537(.A1(new_n16446_), .A2(new_n16447_), .B(new_n16637_), .ZN(new_n16638_));
  AOI21_X1   g16538(.A1(new_n16638_), .A2(new_n16635_), .B(new_n16633_), .ZN(new_n16639_));
  OAI21_X1   g16539(.A1(new_n16614_), .A2(new_n16615_), .B(new_n16556_), .ZN(new_n16640_));
  NAND3_X1   g16540(.A1(new_n16612_), .A2(new_n16607_), .A3(new_n16557_), .ZN(new_n16641_));
  NAND3_X1   g16541(.A1(new_n16625_), .A2(new_n16549_), .A3(new_n16622_), .ZN(new_n16642_));
  OAI21_X1   g16542(.A1(new_n16619_), .A2(new_n16617_), .B(new_n16623_), .ZN(new_n16643_));
  AOI22_X1   g16543(.A1(new_n16642_), .A2(new_n16643_), .B1(new_n16640_), .B2(new_n16641_), .ZN(new_n16644_));
  AOI21_X1   g16544(.A1(new_n16628_), .A2(new_n16631_), .B(new_n16644_), .ZN(new_n16645_));
  AOI21_X1   g16545(.A1(new_n16444_), .A2(new_n16440_), .B(new_n16636_), .ZN(new_n16646_));
  NOR3_X1    g16546(.A1(new_n16646_), .A2(new_n16645_), .A3(new_n16634_), .ZN(new_n16647_));
  OAI21_X1   g16547(.A1(new_n16639_), .A2(new_n16647_), .B(new_n16552_), .ZN(new_n16648_));
  INV_X1     g16548(.I(new_n16552_), .ZN(new_n16649_));
  OAI21_X1   g16549(.A1(new_n16646_), .A2(new_n16634_), .B(new_n16645_), .ZN(new_n16650_));
  NAND3_X1   g16550(.A1(new_n16638_), .A2(new_n16633_), .A3(new_n16635_), .ZN(new_n16651_));
  NAND3_X1   g16551(.A1(new_n16650_), .A2(new_n16651_), .A3(new_n16649_), .ZN(new_n16652_));
  AOI21_X1   g16552(.A1(new_n16648_), .A2(new_n16652_), .B(new_n16543_), .ZN(new_n16653_));
  AOI21_X1   g16553(.A1(new_n16650_), .A2(new_n16651_), .B(new_n16649_), .ZN(new_n16654_));
  NOR3_X1    g16554(.A1(new_n16639_), .A2(new_n16647_), .A3(new_n16552_), .ZN(new_n16655_));
  NOR3_X1    g16555(.A1(new_n16654_), .A2(new_n16655_), .A3(new_n16542_), .ZN(new_n16656_));
  OAI22_X1   g16556(.A1(new_n14276_), .A2(new_n2258_), .B1(new_n6756_), .B2(new_n14594_), .ZN(new_n16657_));
  OAI21_X1   g16557(.A1(new_n14886_), .A2(new_n1078_), .B(new_n16657_), .ZN(new_n16658_));
  AOI21_X1   g16558(.A1(new_n16658_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n16659_));
  XOR2_X1    g16559(.A1(new_n14891_), .A2(new_n16659_), .Z(new_n16660_));
  NOR3_X1    g16560(.A1(new_n16656_), .A2(new_n16653_), .A3(new_n16660_), .ZN(new_n16661_));
  OAI21_X1   g16561(.A1(new_n16654_), .A2(new_n16655_), .B(new_n16542_), .ZN(new_n16662_));
  NAND3_X1   g16562(.A1(new_n16648_), .A2(new_n16652_), .A3(new_n16543_), .ZN(new_n16663_));
  INV_X1     g16563(.I(new_n16660_), .ZN(new_n16664_));
  AOI21_X1   g16564(.A1(new_n16662_), .A2(new_n16663_), .B(new_n16664_), .ZN(new_n16665_));
  OAI21_X1   g16565(.A1(new_n16661_), .A2(new_n16665_), .B(new_n16538_), .ZN(new_n16666_));
  NAND3_X1   g16566(.A1(new_n16662_), .A2(new_n16663_), .A3(new_n16664_), .ZN(new_n16667_));
  OAI21_X1   g16567(.A1(new_n16656_), .A2(new_n16653_), .B(new_n16660_), .ZN(new_n16668_));
  NAND3_X1   g16568(.A1(new_n16668_), .A2(new_n16667_), .A3(new_n16537_), .ZN(new_n16669_));
  AOI21_X1   g16569(.A1(new_n16666_), .A2(new_n16669_), .B(new_n16533_), .ZN(new_n16670_));
  AOI21_X1   g16570(.A1(new_n16668_), .A2(new_n16667_), .B(new_n16537_), .ZN(new_n16671_));
  NOR3_X1    g16571(.A1(new_n16661_), .A2(new_n16665_), .A3(new_n16538_), .ZN(new_n16672_));
  NOR3_X1    g16572(.A1(new_n16672_), .A2(new_n16671_), .A3(new_n16532_), .ZN(new_n16673_));
  AOI21_X1   g16573(.A1(new_n16488_), .A2(new_n16484_), .B(new_n16321_), .ZN(new_n16674_));
  NAND3_X1   g16574(.A1(new_n16488_), .A2(new_n16321_), .A3(new_n16484_), .ZN(new_n16675_));
  AOI21_X1   g16575(.A1(new_n16463_), .A2(new_n16467_), .B(new_n16473_), .ZN(new_n16676_));
  INV_X1     g16576(.I(new_n16474_), .ZN(new_n16677_));
  OAI21_X1   g16577(.A1(new_n16676_), .A2(new_n16677_), .B(new_n16476_), .ZN(new_n16678_));
  NAND2_X1   g16578(.A1(new_n16480_), .A2(new_n16477_), .ZN(new_n16679_));
  NAND3_X1   g16579(.A1(new_n16679_), .A2(new_n16449_), .A3(new_n16453_), .ZN(new_n16680_));
  NAND3_X1   g16580(.A1(new_n16680_), .A2(new_n16678_), .A3(new_n16335_), .ZN(new_n16681_));
  OAI21_X1   g16581(.A1(new_n16481_), .A2(new_n16475_), .B(new_n16334_), .ZN(new_n16682_));
  NAND2_X1   g16582(.A1(new_n16682_), .A2(new_n16681_), .ZN(new_n16683_));
  AOI21_X1   g16583(.A1(new_n16683_), .A2(new_n16675_), .B(new_n16674_), .ZN(new_n16684_));
  NOR3_X1    g16584(.A1(new_n16673_), .A2(new_n16670_), .A3(new_n16684_), .ZN(new_n16685_));
  OAI21_X1   g16585(.A1(new_n16672_), .A2(new_n16671_), .B(new_n16532_), .ZN(new_n16686_));
  NAND3_X1   g16586(.A1(new_n16666_), .A2(new_n16669_), .A3(new_n16533_), .ZN(new_n16687_));
  NAND3_X1   g16587(.A1(new_n16268_), .A2(new_n16269_), .A3(new_n16486_), .ZN(new_n16688_));
  OAI21_X1   g16588(.A1(new_n16263_), .A2(new_n16260_), .B(new_n16116_), .ZN(new_n16689_));
  AOI22_X1   g16589(.A1(new_n16689_), .A2(new_n16688_), .B1(new_n16125_), .B2(new_n16266_), .ZN(new_n16690_));
  OAI21_X1   g16590(.A1(new_n16690_), .A2(new_n16483_), .B(new_n16497_), .ZN(new_n16691_));
  NOR3_X1    g16591(.A1(new_n16690_), .A2(new_n16497_), .A3(new_n16483_), .ZN(new_n16692_));
  NOR3_X1    g16592(.A1(new_n16481_), .A2(new_n16475_), .A3(new_n16334_), .ZN(new_n16693_));
  AOI21_X1   g16593(.A1(new_n16680_), .A2(new_n16678_), .B(new_n16335_), .ZN(new_n16694_));
  NOR2_X1    g16594(.A1(new_n16694_), .A2(new_n16693_), .ZN(new_n16695_));
  OAI21_X1   g16595(.A1(new_n16695_), .A2(new_n16692_), .B(new_n16691_), .ZN(new_n16696_));
  AOI21_X1   g16596(.A1(new_n16686_), .A2(new_n16687_), .B(new_n16696_), .ZN(new_n16697_));
  OAI21_X1   g16597(.A1(new_n16685_), .A2(new_n16697_), .B(new_n16528_), .ZN(new_n16698_));
  NAND3_X1   g16598(.A1(new_n16686_), .A2(new_n16687_), .A3(new_n16696_), .ZN(new_n16699_));
  OAI21_X1   g16599(.A1(new_n16673_), .A2(new_n16670_), .B(new_n16684_), .ZN(new_n16700_));
  NAND3_X1   g16600(.A1(new_n16700_), .A2(new_n16699_), .A3(new_n16527_), .ZN(new_n16701_));
  AOI21_X1   g16601(.A1(new_n16698_), .A2(new_n16701_), .B(new_n16523_), .ZN(new_n16702_));
  AOI21_X1   g16602(.A1(new_n16700_), .A2(new_n16699_), .B(new_n16527_), .ZN(new_n16703_));
  NOR3_X1    g16603(.A1(new_n16685_), .A2(new_n16697_), .A3(new_n16528_), .ZN(new_n16704_));
  NOR3_X1    g16604(.A1(new_n16704_), .A2(new_n16703_), .A3(new_n16522_), .ZN(new_n16705_));
  NOR2_X1    g16605(.A1(new_n16501_), .A2(new_n16317_), .ZN(new_n16706_));
  NOR2_X1    g16606(.A1(new_n16505_), .A2(new_n16318_), .ZN(new_n16707_));
  OAI22_X1   g16607(.A1(new_n16707_), .A2(new_n16706_), .B1(new_n16702_), .B2(new_n16705_), .ZN(new_n16708_));
  NOR2_X1    g16608(.A1(new_n16708_), .A2(new_n16506_), .ZN(new_n16709_));
  NOR2_X1    g16609(.A1(new_n16505_), .A2(new_n16317_), .ZN(new_n16710_));
  NOR2_X1    g16610(.A1(new_n16709_), .A2(new_n16710_), .ZN(new_n16711_));
  XOR2_X1    g16611(.A1(new_n16711_), .A2(new_n16518_), .Z(new_n16712_));
  XOR2_X1    g16612(.A1(new_n16510_), .A2(new_n16712_), .Z(\result[11] ));
  AOI21_X1   g16613(.A1(new_n15898_), .A2(new_n16100_), .B(new_n16304_), .ZN(new_n16714_));
  NOR3_X1    g16614(.A1(new_n16105_), .A2(new_n16106_), .A3(new_n16305_), .ZN(new_n16715_));
  INV_X1     g16615(.I(new_n16507_), .ZN(new_n16716_));
  OAI21_X1   g16616(.A1(new_n16715_), .A2(new_n16714_), .B(new_n16716_), .ZN(new_n16717_));
  XOR2_X1    g16617(.A1(new_n16711_), .A2(new_n16314_), .Z(new_n16718_));
  NOR3_X1    g16618(.A1(new_n16705_), .A2(new_n16702_), .A3(new_n16501_), .ZN(new_n16719_));
  OAI21_X1   g16619(.A1(new_n16705_), .A2(new_n16702_), .B(new_n16501_), .ZN(new_n16720_));
  AOI21_X1   g16620(.A1(new_n16317_), .A2(new_n16720_), .B(new_n16719_), .ZN(new_n16721_));
  NAND2_X1   g16621(.A1(new_n16314_), .A2(new_n16721_), .ZN(new_n16722_));
  NAND2_X1   g16622(.A1(new_n16686_), .A2(new_n16687_), .ZN(new_n16723_));
  XOR2_X1    g16623(.A1(new_n16723_), .A2(new_n16527_), .Z(new_n16724_));
  XOR2_X1    g16624(.A1(new_n16724_), .A2(new_n16522_), .Z(new_n16725_));
  NOR2_X1    g16625(.A1(new_n16725_), .A2(new_n16684_), .ZN(new_n16726_));
  OAI22_X1   g16626(.A1(new_n10913_), .A2(new_n1239_), .B1(new_n12768_), .B2(new_n4981_), .ZN(new_n16727_));
  AOI21_X1   g16627(.A1(new_n16727_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n16728_));
  XOR2_X1    g16628(.A1(new_n12767_), .A2(new_n16728_), .Z(new_n16729_));
  NOR2_X1    g16629(.A1(new_n16563_), .A2(new_n16600_), .ZN(new_n16730_));
  NAND2_X1   g16630(.A1(new_n16563_), .A2(new_n16600_), .ZN(new_n16731_));
  NOR2_X1    g16631(.A1(new_n16603_), .A2(new_n16604_), .ZN(new_n16732_));
  XOR2_X1    g16632(.A1(new_n16732_), .A2(new_n16556_), .Z(new_n16733_));
  AOI21_X1   g16633(.A1(new_n16733_), .A2(new_n16731_), .B(new_n16730_), .ZN(new_n16734_));
  INV_X1     g16634(.I(new_n16734_), .ZN(new_n16735_));
  OAI22_X1   g16635(.A1(new_n10619_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10881_), .ZN(new_n16736_));
  OAI21_X1   g16636(.A1(new_n79_), .A2(new_n10611_), .B(new_n16736_), .ZN(new_n16737_));
  AOI21_X1   g16637(.A1(new_n16737_), .A2(new_n72_), .B(new_n79_), .ZN(new_n16738_));
  XOR2_X1    g16638(.A1(new_n12090_), .A2(new_n16738_), .Z(new_n16739_));
  XOR2_X1    g16639(.A1(new_n16569_), .A2(new_n16574_), .Z(new_n16740_));
  INV_X1     g16640(.I(new_n16740_), .ZN(new_n16741_));
  NOR2_X1    g16641(.A1(new_n10870_), .A2(new_n88_), .ZN(new_n16742_));
  OAI22_X1   g16642(.A1(new_n10868_), .A2(new_n511_), .B1(new_n92_), .B2(new_n10856_), .ZN(new_n16743_));
  OAI21_X1   g16643(.A1(new_n16742_), .A2(new_n16743_), .B(new_n961_), .ZN(new_n16744_));
  NOR2_X1    g16644(.A1(new_n11722_), .A2(new_n16744_), .ZN(new_n16745_));
  NOR2_X1    g16645(.A1(new_n16741_), .A2(new_n16745_), .ZN(new_n16746_));
  INV_X1     g16646(.I(new_n16746_), .ZN(new_n16747_));
  NAND2_X1   g16647(.A1(new_n16741_), .A2(new_n16745_), .ZN(new_n16748_));
  NAND2_X1   g16648(.A1(new_n16747_), .A2(new_n16748_), .ZN(new_n16749_));
  NAND2_X1   g16649(.A1(new_n16588_), .A2(new_n16589_), .ZN(new_n16750_));
  NAND2_X1   g16650(.A1(new_n16750_), .A2(new_n16590_), .ZN(new_n16751_));
  AOI22_X1   g16651(.A1(new_n12204_), .A2(new_n4767_), .B1(new_n4613_), .B2(new_n10897_), .ZN(new_n16752_));
  AOI21_X1   g16652(.A1(new_n117_), .A2(new_n10600_), .B(new_n16752_), .ZN(new_n16753_));
  OAI21_X1   g16653(.A1(new_n16753_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n16754_));
  XNOR2_X1   g16654(.A1(new_n12576_), .A2(new_n16754_), .ZN(new_n16755_));
  XOR2_X1    g16655(.A1(new_n16751_), .A2(new_n16755_), .Z(new_n16756_));
  XOR2_X1    g16656(.A1(new_n16756_), .A2(new_n16749_), .Z(new_n16757_));
  XNOR2_X1   g16657(.A1(new_n16757_), .A2(new_n16739_), .ZN(new_n16758_));
  AOI22_X1   g16658(.A1(new_n16596_), .A2(new_n16556_), .B1(new_n16565_), .B2(new_n16567_), .ZN(new_n16759_));
  NOR2_X1    g16659(.A1(new_n16596_), .A2(new_n16556_), .ZN(new_n16760_));
  NOR2_X1    g16660(.A1(new_n16759_), .A2(new_n16760_), .ZN(new_n16761_));
  INV_X1     g16661(.I(new_n16761_), .ZN(new_n16762_));
  NAND2_X1   g16662(.A1(new_n16758_), .A2(new_n16762_), .ZN(new_n16763_));
  XOR2_X1    g16663(.A1(new_n16757_), .A2(new_n16739_), .Z(new_n16764_));
  NAND2_X1   g16664(.A1(new_n16764_), .A2(new_n16761_), .ZN(new_n16765_));
  OAI22_X1   g16665(.A1(new_n13395_), .A2(new_n5336_), .B1(new_n5398_), .B2(new_n10938_), .ZN(new_n16766_));
  AOI21_X1   g16666(.A1(new_n16766_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n16767_));
  XOR2_X1    g16667(.A1(new_n13394_), .A2(new_n16767_), .Z(new_n16768_));
  INV_X1     g16668(.I(new_n16768_), .ZN(new_n16769_));
  NAND3_X1   g16669(.A1(new_n16763_), .A2(new_n16765_), .A3(new_n16769_), .ZN(new_n16770_));
  INV_X1     g16670(.I(new_n16770_), .ZN(new_n16771_));
  AOI21_X1   g16671(.A1(new_n16763_), .A2(new_n16765_), .B(new_n16769_), .ZN(new_n16772_));
  NOR2_X1    g16672(.A1(new_n16771_), .A2(new_n16772_), .ZN(new_n16773_));
  NOR2_X1    g16673(.A1(new_n16773_), .A2(new_n16735_), .ZN(new_n16774_));
  INV_X1     g16674(.I(new_n16772_), .ZN(new_n16775_));
  NAND2_X1   g16675(.A1(new_n16775_), .A2(new_n16770_), .ZN(new_n16776_));
  NOR2_X1    g16676(.A1(new_n16776_), .A2(new_n16734_), .ZN(new_n16777_));
  OAI21_X1   g16677(.A1(new_n16777_), .A2(new_n16774_), .B(new_n16729_), .ZN(new_n16778_));
  INV_X1     g16678(.I(new_n16729_), .ZN(new_n16779_));
  NAND2_X1   g16679(.A1(new_n16776_), .A2(new_n16734_), .ZN(new_n16780_));
  NAND2_X1   g16680(.A1(new_n16773_), .A2(new_n16735_), .ZN(new_n16781_));
  NAND3_X1   g16681(.A1(new_n16780_), .A2(new_n16781_), .A3(new_n16779_), .ZN(new_n16782_));
  NAND2_X1   g16682(.A1(new_n16778_), .A2(new_n16782_), .ZN(new_n16783_));
  OAI21_X1   g16683(.A1(new_n16628_), .A2(new_n16624_), .B(new_n16643_), .ZN(new_n16784_));
  OAI22_X1   g16684(.A1(new_n14054_), .A2(new_n5420_), .B1(new_n1620_), .B2(new_n10961_), .ZN(new_n16785_));
  AOI21_X1   g16685(.A1(new_n16785_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n16786_));
  XOR2_X1    g16686(.A1(new_n14053_), .A2(new_n16786_), .Z(new_n16787_));
  INV_X1     g16687(.I(new_n16787_), .ZN(new_n16788_));
  NOR2_X1    g16688(.A1(new_n16784_), .A2(new_n16788_), .ZN(new_n16789_));
  INV_X1     g16689(.I(new_n16789_), .ZN(new_n16790_));
  NAND2_X1   g16690(.A1(new_n16784_), .A2(new_n16788_), .ZN(new_n16791_));
  NAND2_X1   g16691(.A1(new_n16790_), .A2(new_n16791_), .ZN(new_n16792_));
  XOR2_X1    g16692(.A1(new_n16784_), .A2(new_n16787_), .Z(new_n16793_));
  NOR2_X1    g16693(.A1(new_n16783_), .A2(new_n16793_), .ZN(new_n16794_));
  AOI21_X1   g16694(.A1(new_n16783_), .A2(new_n16792_), .B(new_n16794_), .ZN(new_n16795_));
  NAND2_X1   g16695(.A1(new_n16552_), .A2(new_n16542_), .ZN(new_n16796_));
  NAND2_X1   g16696(.A1(new_n16633_), .A2(new_n16796_), .ZN(new_n16797_));
  NAND2_X1   g16697(.A1(new_n16649_), .A2(new_n16543_), .ZN(new_n16798_));
  NAND2_X1   g16698(.A1(new_n16797_), .A2(new_n16798_), .ZN(new_n16799_));
  AOI22_X1   g16699(.A1(new_n14281_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n14274_), .ZN(new_n16800_));
  OAI21_X1   g16700(.A1(new_n16800_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n16801_));
  XOR2_X1    g16701(.A1(new_n14280_), .A2(new_n16801_), .Z(new_n16802_));
  INV_X1     g16702(.I(new_n16802_), .ZN(new_n16803_));
  NOR2_X1    g16703(.A1(new_n16799_), .A2(new_n16803_), .ZN(new_n16804_));
  NAND2_X1   g16704(.A1(new_n16799_), .A2(new_n16803_), .ZN(new_n16805_));
  INV_X1     g16705(.I(new_n16805_), .ZN(new_n16806_));
  NOR2_X1    g16706(.A1(new_n16806_), .A2(new_n16804_), .ZN(new_n16807_));
  NOR2_X1    g16707(.A1(new_n16795_), .A2(new_n16807_), .ZN(new_n16808_));
  XOR2_X1    g16708(.A1(new_n16799_), .A2(new_n16803_), .Z(new_n16809_));
  AOI21_X1   g16709(.A1(new_n16795_), .A2(new_n16809_), .B(new_n16808_), .ZN(new_n16810_));
  NOR2_X1    g16710(.A1(new_n16646_), .A2(new_n16634_), .ZN(new_n16811_));
  AOI21_X1   g16711(.A1(new_n16798_), .A2(new_n16796_), .B(new_n16645_), .ZN(new_n16812_));
  XOR2_X1    g16712(.A1(new_n16552_), .A2(new_n16542_), .Z(new_n16813_));
  AOI21_X1   g16713(.A1(new_n16645_), .A2(new_n16813_), .B(new_n16812_), .ZN(new_n16814_));
  AOI21_X1   g16714(.A1(new_n16811_), .A2(new_n16532_), .B(new_n16814_), .ZN(new_n16815_));
  NOR2_X1    g16715(.A1(new_n16811_), .A2(new_n16532_), .ZN(new_n16816_));
  NOR2_X1    g16716(.A1(new_n16815_), .A2(new_n16816_), .ZN(new_n16817_));
  AOI22_X1   g16717(.A1(new_n15127_), .A2(new_n6758_), .B1(new_n805_), .B2(new_n15115_), .ZN(new_n16818_));
  OAI21_X1   g16718(.A1(new_n16818_), .A2(\a[11] ), .B(new_n805_), .ZN(new_n16819_));
  XNOR2_X1   g16719(.A1(new_n15125_), .A2(new_n16819_), .ZN(new_n16820_));
  NAND2_X1   g16720(.A1(new_n16817_), .A2(new_n16820_), .ZN(new_n16821_));
  NOR2_X1    g16721(.A1(new_n16817_), .A2(new_n16820_), .ZN(new_n16822_));
  INV_X1     g16722(.I(new_n16822_), .ZN(new_n16823_));
  AND2_X2    g16723(.A1(new_n16823_), .A2(new_n16821_), .Z(new_n16824_));
  XOR2_X1    g16724(.A1(new_n16817_), .A2(new_n16820_), .Z(new_n16825_));
  NAND2_X1   g16725(.A1(new_n16810_), .A2(new_n16825_), .ZN(new_n16826_));
  OAI21_X1   g16726(.A1(new_n16824_), .A2(new_n16810_), .B(new_n16826_), .ZN(new_n16827_));
  NAND3_X1   g16727(.A1(new_n16662_), .A2(new_n16663_), .A3(new_n16533_), .ZN(new_n16828_));
  OAI21_X1   g16728(.A1(new_n16656_), .A2(new_n16653_), .B(new_n16532_), .ZN(new_n16829_));
  AOI22_X1   g16729(.A1(new_n16829_), .A2(new_n16828_), .B1(new_n16538_), .B2(new_n16660_), .ZN(new_n16830_));
  AOI21_X1   g16730(.A1(new_n16537_), .A2(new_n16664_), .B(new_n16830_), .ZN(new_n16831_));
  NAND2_X1   g16731(.A1(new_n15515_), .A2(new_n5110_), .ZN(new_n16832_));
  NOR2_X1    g16732(.A1(new_n5108_), .A2(new_n2469_), .ZN(new_n16833_));
  AOI21_X1   g16733(.A1(new_n15675_), .A2(new_n16833_), .B(\a[8] ), .ZN(new_n16834_));
  AOI21_X1   g16734(.A1(new_n16834_), .A2(new_n16832_), .B(new_n2495_), .ZN(new_n16835_));
  XNOR2_X1   g16735(.A1(new_n15678_), .A2(new_n16835_), .ZN(new_n16836_));
  XNOR2_X1   g16736(.A1(new_n16831_), .A2(new_n16836_), .ZN(new_n16837_));
  OAI21_X1   g16737(.A1(new_n16523_), .A2(new_n16527_), .B(new_n16723_), .ZN(new_n16838_));
  OAI21_X1   g16738(.A1(new_n16522_), .A2(new_n16528_), .B(new_n16838_), .ZN(new_n16839_));
  XOR2_X1    g16739(.A1(new_n16839_), .A2(new_n16837_), .Z(new_n16840_));
  NAND2_X1   g16740(.A1(new_n16840_), .A2(new_n16827_), .ZN(new_n16841_));
  INV_X1     g16741(.I(new_n16827_), .ZN(new_n16842_));
  INV_X1     g16742(.I(new_n16837_), .ZN(new_n16843_));
  XOR2_X1    g16743(.A1(new_n16839_), .A2(new_n16843_), .Z(new_n16844_));
  NAND2_X1   g16744(.A1(new_n16844_), .A2(new_n16842_), .ZN(new_n16845_));
  AOI21_X1   g16745(.A1(new_n16845_), .A2(new_n16841_), .B(new_n16726_), .ZN(new_n16846_));
  NAND2_X1   g16746(.A1(new_n16846_), .A2(new_n16722_), .ZN(new_n16847_));
  XOR2_X1    g16747(.A1(new_n16839_), .A2(new_n16843_), .Z(new_n16848_));
  NOR2_X1    g16748(.A1(new_n16848_), .A2(new_n16842_), .ZN(new_n16849_));
  AOI21_X1   g16749(.A1(new_n16842_), .A2(new_n16844_), .B(new_n16849_), .ZN(new_n16850_));
  OAI21_X1   g16750(.A1(new_n16704_), .A2(new_n16703_), .B(new_n16522_), .ZN(new_n16851_));
  NAND3_X1   g16751(.A1(new_n16698_), .A2(new_n16701_), .A3(new_n16523_), .ZN(new_n16852_));
  NAND3_X1   g16752(.A1(new_n16851_), .A2(new_n16852_), .A3(new_n16505_), .ZN(new_n16853_));
  AOI21_X1   g16753(.A1(new_n16851_), .A2(new_n16852_), .B(new_n16505_), .ZN(new_n16854_));
  OAI21_X1   g16754(.A1(new_n16318_), .A2(new_n16854_), .B(new_n16853_), .ZN(new_n16855_));
  OAI22_X1   g16755(.A1(new_n16518_), .A2(new_n16855_), .B1(new_n16684_), .B2(new_n16725_), .ZN(new_n16856_));
  NAND2_X1   g16756(.A1(new_n16850_), .A2(new_n16856_), .ZN(new_n16857_));
  NAND2_X1   g16757(.A1(new_n16857_), .A2(new_n16847_), .ZN(new_n16858_));
  OAI21_X1   g16758(.A1(new_n16717_), .A2(new_n16718_), .B(new_n16858_), .ZN(new_n16859_));
  AOI22_X1   g16759(.A1(new_n16850_), .A2(new_n16856_), .B1(new_n16846_), .B2(new_n16722_), .ZN(new_n16860_));
  NAND4_X1   g16760(.A1(\result[9] ), .A2(new_n16716_), .A3(new_n16712_), .A4(new_n16860_), .ZN(new_n16861_));
  NAND2_X1   g16761(.A1(new_n16859_), .A2(new_n16861_), .ZN(\result[12] ));
  NAND2_X1   g16762(.A1(new_n16510_), .A2(new_n16712_), .ZN(new_n16863_));
  XNOR2_X1   g16763(.A1(new_n16827_), .A2(new_n16837_), .ZN(new_n16864_));
  NAND3_X1   g16764(.A1(new_n16314_), .A2(new_n16721_), .A3(new_n16864_), .ZN(new_n16865_));
  AOI21_X1   g16765(.A1(new_n16314_), .A2(new_n16721_), .B(new_n16864_), .ZN(new_n16866_));
  AND4_X2    g16766(.A1(new_n16523_), .A2(new_n16723_), .A3(new_n16527_), .A4(new_n16696_), .Z(new_n16867_));
  INV_X1     g16767(.I(new_n16867_), .ZN(new_n16868_));
  OAI21_X1   g16768(.A1(new_n16866_), .A2(new_n16868_), .B(new_n16865_), .ZN(new_n16869_));
  NAND2_X1   g16769(.A1(new_n16831_), .A2(new_n16836_), .ZN(new_n16870_));
  NOR2_X1    g16770(.A1(new_n16831_), .A2(new_n16836_), .ZN(new_n16871_));
  AOI21_X1   g16771(.A1(new_n16827_), .A2(new_n16870_), .B(new_n16871_), .ZN(new_n16872_));
  INV_X1     g16772(.I(new_n16872_), .ZN(new_n16873_));
  AOI22_X1   g16773(.A1(new_n14602_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n14603_), .ZN(new_n16874_));
  OAI21_X1   g16774(.A1(new_n16874_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n16875_));
  XNOR2_X1   g16775(.A1(new_n14601_), .A2(new_n16875_), .ZN(new_n16876_));
  INV_X1     g16776(.I(new_n16876_), .ZN(new_n16877_));
  INV_X1     g16777(.I(new_n16791_), .ZN(new_n16878_));
  OAI21_X1   g16778(.A1(new_n16789_), .A2(new_n16878_), .B(new_n16783_), .ZN(new_n16879_));
  OAI21_X1   g16779(.A1(new_n16783_), .A2(new_n16793_), .B(new_n16879_), .ZN(new_n16880_));
  INV_X1     g16780(.I(new_n16804_), .ZN(new_n16881_));
  AOI21_X1   g16781(.A1(new_n16880_), .A2(new_n16881_), .B(new_n16806_), .ZN(new_n16882_));
  AOI21_X1   g16782(.A1(new_n16778_), .A2(new_n16782_), .B(new_n16789_), .ZN(new_n16883_));
  OAI22_X1   g16783(.A1(new_n10965_), .A2(new_n5420_), .B1(new_n1620_), .B2(new_n10570_), .ZN(new_n16884_));
  AOI21_X1   g16784(.A1(new_n16884_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n16885_));
  XNOR2_X1   g16785(.A1(new_n14077_), .A2(new_n16885_), .ZN(new_n16886_));
  INV_X1     g16786(.I(new_n16886_), .ZN(new_n16887_));
  NOR3_X1    g16787(.A1(new_n16883_), .A2(new_n16878_), .A3(new_n16887_), .ZN(new_n16888_));
  OAI21_X1   g16788(.A1(new_n16883_), .A2(new_n16878_), .B(new_n16887_), .ZN(new_n16889_));
  INV_X1     g16789(.I(new_n16889_), .ZN(new_n16890_));
  NOR2_X1    g16790(.A1(new_n16761_), .A2(new_n16729_), .ZN(new_n16891_));
  INV_X1     g16791(.I(new_n16891_), .ZN(new_n16892_));
  OAI22_X1   g16792(.A1(new_n10606_), .A2(new_n4612_), .B1(new_n4781_), .B2(new_n10599_), .ZN(new_n16893_));
  OAI21_X1   g16793(.A1(new_n10595_), .A2(new_n1128_), .B(new_n16893_), .ZN(new_n16894_));
  AOI21_X1   g16794(.A1(new_n16894_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n16895_));
  XOR2_X1    g16795(.A1(new_n12600_), .A2(new_n16895_), .Z(new_n16896_));
  OR2_X2     g16796(.A1(new_n16755_), .A2(new_n16739_), .Z(new_n16897_));
  NAND2_X1   g16797(.A1(new_n16755_), .A2(new_n16739_), .ZN(new_n16898_));
  XOR2_X1    g16798(.A1(new_n16749_), .A2(new_n16751_), .Z(new_n16899_));
  NAND2_X1   g16799(.A1(new_n16899_), .A2(new_n16898_), .ZN(new_n16900_));
  NAND2_X1   g16800(.A1(new_n16900_), .A2(new_n16897_), .ZN(new_n16901_));
  INV_X1     g16801(.I(new_n16751_), .ZN(new_n16902_));
  NAND2_X1   g16802(.A1(new_n10875_), .A2(new_n87_), .ZN(new_n16903_));
  AOI22_X1   g16803(.A1(new_n10882_), .A2(new_n962_), .B1(new_n10625_), .B2(new_n4406_), .ZN(new_n16904_));
  AOI21_X1   g16804(.A1(new_n16904_), .A2(new_n16903_), .B(new_n82_), .ZN(new_n16905_));
  NAND2_X1   g16805(.A1(new_n11802_), .A2(new_n16905_), .ZN(new_n16906_));
  NOR2_X1    g16806(.A1(new_n15515_), .A2(new_n5111_), .ZN(new_n16907_));
  OAI22_X1   g16807(.A1(new_n16907_), .A2(\a[8] ), .B1(new_n5113_), .B2(new_n15515_), .ZN(new_n16908_));
  INV_X1     g16808(.I(new_n16908_), .ZN(new_n16909_));
  OAI22_X1   g16809(.A1(new_n10619_), .A2(new_n4529_), .B1(new_n4527_), .B2(new_n10611_), .ZN(new_n16910_));
  OAI21_X1   g16810(.A1(new_n79_), .A2(new_n10896_), .B(new_n16910_), .ZN(new_n16911_));
  AOI21_X1   g16811(.A1(new_n16911_), .A2(new_n72_), .B(new_n79_), .ZN(new_n16912_));
  XOR2_X1    g16812(.A1(new_n10984_), .A2(new_n16912_), .Z(new_n16913_));
  XOR2_X1    g16813(.A1(new_n16576_), .A2(new_n16913_), .Z(new_n16914_));
  XOR2_X1    g16814(.A1(new_n16914_), .A2(new_n16909_), .Z(new_n16915_));
  XOR2_X1    g16815(.A1(new_n16915_), .A2(new_n16906_), .Z(new_n16916_));
  OAI21_X1   g16816(.A1(new_n16916_), .A2(new_n16748_), .B(new_n16747_), .ZN(new_n16917_));
  NAND2_X1   g16817(.A1(new_n16917_), .A2(new_n16902_), .ZN(new_n16918_));
  OR2_X2     g16818(.A1(new_n16917_), .A2(new_n16902_), .Z(new_n16919_));
  OAI22_X1   g16819(.A1(new_n12890_), .A2(new_n4981_), .B1(new_n10923_), .B2(new_n1239_), .ZN(new_n16920_));
  AOI21_X1   g16820(.A1(new_n16920_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n16921_));
  XOR2_X1    g16821(.A1(new_n12889_), .A2(new_n16921_), .Z(new_n16922_));
  INV_X1     g16822(.I(new_n16922_), .ZN(new_n16923_));
  NAND3_X1   g16823(.A1(new_n16919_), .A2(new_n16918_), .A3(new_n16923_), .ZN(new_n16924_));
  INV_X1     g16824(.I(new_n16918_), .ZN(new_n16925_));
  NOR2_X1    g16825(.A1(new_n16917_), .A2(new_n16902_), .ZN(new_n16926_));
  OAI21_X1   g16826(.A1(new_n16925_), .A2(new_n16926_), .B(new_n16922_), .ZN(new_n16927_));
  AOI21_X1   g16827(.A1(new_n16927_), .A2(new_n16924_), .B(new_n16901_), .ZN(new_n16928_));
  INV_X1     g16828(.I(new_n16901_), .ZN(new_n16929_));
  NOR3_X1    g16829(.A1(new_n16925_), .A2(new_n16926_), .A3(new_n16922_), .ZN(new_n16930_));
  AOI21_X1   g16830(.A1(new_n16919_), .A2(new_n16918_), .B(new_n16923_), .ZN(new_n16931_));
  NOR3_X1    g16831(.A1(new_n16930_), .A2(new_n16931_), .A3(new_n16929_), .ZN(new_n16932_));
  OAI21_X1   g16832(.A1(new_n16932_), .A2(new_n16928_), .B(new_n16896_), .ZN(new_n16933_));
  INV_X1     g16833(.I(new_n16896_), .ZN(new_n16934_));
  OAI21_X1   g16834(.A1(new_n16930_), .A2(new_n16931_), .B(new_n16929_), .ZN(new_n16935_));
  NAND3_X1   g16835(.A1(new_n16927_), .A2(new_n16924_), .A3(new_n16901_), .ZN(new_n16936_));
  NAND3_X1   g16836(.A1(new_n16935_), .A2(new_n16936_), .A3(new_n16934_), .ZN(new_n16937_));
  NAND2_X1   g16837(.A1(new_n16933_), .A2(new_n16937_), .ZN(new_n16938_));
  XOR2_X1    g16838(.A1(new_n16761_), .A2(new_n16729_), .Z(new_n16939_));
  NAND3_X1   g16839(.A1(new_n16938_), .A2(new_n16892_), .A3(new_n16939_), .ZN(new_n16940_));
  NOR2_X1    g16840(.A1(new_n16761_), .A2(new_n16729_), .ZN(new_n16942_));
  INV_X1     g16841(.I(new_n16942_), .ZN(new_n16943_));
  AOI21_X1   g16842(.A1(new_n16940_), .A2(new_n16943_), .B(new_n16764_), .ZN(new_n16944_));
  AOI21_X1   g16843(.A1(new_n16935_), .A2(new_n16936_), .B(new_n16934_), .ZN(new_n16945_));
  NOR3_X1    g16844(.A1(new_n16932_), .A2(new_n16928_), .A3(new_n16896_), .ZN(new_n16946_));
  OAI21_X1   g16845(.A1(new_n16946_), .A2(new_n16945_), .B(new_n16939_), .ZN(new_n16947_));
  NOR2_X1    g16846(.A1(new_n16947_), .A2(new_n16891_), .ZN(new_n16948_));
  NOR3_X1    g16847(.A1(new_n16948_), .A2(new_n16758_), .A3(new_n16942_), .ZN(new_n16949_));
  NOR2_X1    g16848(.A1(new_n16949_), .A2(new_n16944_), .ZN(new_n16950_));
  OAI21_X1   g16849(.A1(new_n16948_), .A2(new_n16942_), .B(new_n16758_), .ZN(new_n16951_));
  NAND3_X1   g16850(.A1(new_n16940_), .A2(new_n16764_), .A3(new_n16943_), .ZN(new_n16952_));
  NOR2_X1    g16851(.A1(new_n16734_), .A2(new_n16768_), .ZN(new_n16953_));
  NAND3_X1   g16852(.A1(new_n16763_), .A2(new_n16765_), .A3(new_n16779_), .ZN(new_n16954_));
  NOR2_X1    g16853(.A1(new_n16764_), .A2(new_n16761_), .ZN(new_n16955_));
  NOR2_X1    g16854(.A1(new_n16758_), .A2(new_n16762_), .ZN(new_n16956_));
  OAI21_X1   g16855(.A1(new_n16956_), .A2(new_n16955_), .B(new_n16729_), .ZN(new_n16957_));
  AOI22_X1   g16856(.A1(new_n16957_), .A2(new_n16954_), .B1(new_n16734_), .B2(new_n16768_), .ZN(new_n16958_));
  NOR2_X1    g16857(.A1(new_n16958_), .A2(new_n16953_), .ZN(new_n16959_));
  AOI22_X1   g16858(.A1(new_n12909_), .A2(new_n5337_), .B1(new_n10949_), .B2(new_n4717_), .ZN(new_n16960_));
  OAI21_X1   g16859(.A1(new_n16960_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n16961_));
  XOR2_X1    g16860(.A1(new_n12907_), .A2(new_n16961_), .Z(new_n16962_));
  NAND2_X1   g16861(.A1(new_n16959_), .A2(new_n16962_), .ZN(new_n16963_));
  NOR2_X1    g16862(.A1(new_n16959_), .A2(new_n16962_), .ZN(new_n16964_));
  INV_X1     g16863(.I(new_n16964_), .ZN(new_n16965_));
  AOI22_X1   g16864(.A1(new_n16965_), .A2(new_n16963_), .B1(new_n16951_), .B2(new_n16952_), .ZN(new_n16966_));
  XOR2_X1    g16865(.A1(new_n16959_), .A2(new_n16962_), .Z(new_n16967_));
  AOI21_X1   g16866(.A1(new_n16950_), .A2(new_n16967_), .B(new_n16966_), .ZN(new_n16968_));
  NOR3_X1    g16867(.A1(new_n16890_), .A2(new_n16968_), .A3(new_n16888_), .ZN(new_n16969_));
  INV_X1     g16868(.I(new_n16888_), .ZN(new_n16970_));
  INV_X1     g16869(.I(new_n16963_), .ZN(new_n16971_));
  NOR2_X1    g16870(.A1(new_n16971_), .A2(new_n16964_), .ZN(new_n16972_));
  NAND2_X1   g16871(.A1(new_n16950_), .A2(new_n16967_), .ZN(new_n16973_));
  OAI21_X1   g16872(.A1(new_n16950_), .A2(new_n16972_), .B(new_n16973_), .ZN(new_n16974_));
  AOI21_X1   g16873(.A1(new_n16970_), .A2(new_n16889_), .B(new_n16974_), .ZN(new_n16975_));
  OAI21_X1   g16874(.A1(new_n16969_), .A2(new_n16975_), .B(new_n16882_), .ZN(new_n16976_));
  OAI21_X1   g16875(.A1(new_n16795_), .A2(new_n16804_), .B(new_n16805_), .ZN(new_n16977_));
  NAND3_X1   g16876(.A1(new_n16974_), .A2(new_n16970_), .A3(new_n16889_), .ZN(new_n16978_));
  OAI21_X1   g16877(.A1(new_n16888_), .A2(new_n16890_), .B(new_n16968_), .ZN(new_n16979_));
  NAND3_X1   g16878(.A1(new_n16978_), .A2(new_n16977_), .A3(new_n16979_), .ZN(new_n16980_));
  AOI21_X1   g16879(.A1(new_n16976_), .A2(new_n16980_), .B(new_n16877_), .ZN(new_n16981_));
  AOI21_X1   g16880(.A1(new_n16978_), .A2(new_n16979_), .B(new_n16977_), .ZN(new_n16982_));
  NOR3_X1    g16881(.A1(new_n16882_), .A2(new_n16975_), .A3(new_n16969_), .ZN(new_n16983_));
  NOR3_X1    g16882(.A1(new_n16983_), .A2(new_n16982_), .A3(new_n16876_), .ZN(new_n16984_));
  NOR2_X1    g16883(.A1(new_n16981_), .A2(new_n16984_), .ZN(new_n16985_));
  INV_X1     g16884(.I(new_n16810_), .ZN(new_n16986_));
  OAI22_X1   g16885(.A1(new_n15313_), .A2(new_n6757_), .B1(new_n1078_), .B2(new_n15305_), .ZN(new_n16987_));
  AOI21_X1   g16886(.A1(new_n16987_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n16988_));
  XNOR2_X1   g16887(.A1(new_n15312_), .A2(new_n16988_), .ZN(new_n16989_));
  INV_X1     g16888(.I(new_n16989_), .ZN(new_n16990_));
  NAND3_X1   g16889(.A1(new_n16825_), .A2(new_n16823_), .A3(new_n16990_), .ZN(new_n16991_));
  NOR2_X1    g16890(.A1(new_n16817_), .A2(new_n16820_), .ZN(new_n16992_));
  INV_X1     g16891(.I(new_n16992_), .ZN(new_n16993_));
  AOI21_X1   g16892(.A1(new_n16991_), .A2(new_n16993_), .B(new_n16986_), .ZN(new_n16994_));
  INV_X1     g16893(.I(new_n16994_), .ZN(new_n16995_));
  NAND3_X1   g16894(.A1(new_n16986_), .A2(new_n16991_), .A3(new_n16993_), .ZN(new_n16996_));
  NAND3_X1   g16895(.A1(new_n16995_), .A2(new_n16985_), .A3(new_n16996_), .ZN(new_n16997_));
  OAI21_X1   g16896(.A1(new_n16983_), .A2(new_n16982_), .B(new_n16876_), .ZN(new_n16998_));
  NAND3_X1   g16897(.A1(new_n16976_), .A2(new_n16877_), .A3(new_n16980_), .ZN(new_n16999_));
  NAND2_X1   g16898(.A1(new_n16999_), .A2(new_n16998_), .ZN(new_n17000_));
  INV_X1     g16899(.I(new_n16996_), .ZN(new_n17001_));
  OAI21_X1   g16900(.A1(new_n17001_), .A2(new_n16994_), .B(new_n17000_), .ZN(new_n17002_));
  NAND2_X1   g16901(.A1(new_n16997_), .A2(new_n17002_), .ZN(new_n17003_));
  NOR2_X1    g16902(.A1(new_n17003_), .A2(new_n16873_), .ZN(new_n17004_));
  NOR3_X1    g16903(.A1(new_n17001_), .A2(new_n17000_), .A3(new_n16994_), .ZN(new_n17005_));
  AOI21_X1   g16904(.A1(new_n16995_), .A2(new_n16996_), .B(new_n16985_), .ZN(new_n17006_));
  NOR2_X1    g16905(.A1(new_n17006_), .A2(new_n17005_), .ZN(new_n17007_));
  NOR2_X1    g16906(.A1(new_n17007_), .A2(new_n16872_), .ZN(new_n17008_));
  OAI21_X1   g16907(.A1(new_n17004_), .A2(new_n17008_), .B(new_n16869_), .ZN(new_n17009_));
  XOR2_X1    g16908(.A1(new_n16863_), .A2(new_n17009_), .Z(new_n17010_));
  XOR2_X1    g16909(.A1(new_n17010_), .A2(new_n16858_), .Z(\result[13] ));
  AOI21_X1   g16910(.A1(new_n16859_), .A2(new_n16861_), .B(new_n17009_), .ZN(new_n17012_));
  XOR2_X1    g16911(.A1(new_n16827_), .A2(new_n16837_), .Z(new_n17013_));
  NOR3_X1    g16912(.A1(new_n16518_), .A2(new_n16855_), .A3(new_n17013_), .ZN(new_n17014_));
  OAI21_X1   g16913(.A1(new_n16518_), .A2(new_n16855_), .B(new_n17013_), .ZN(new_n17015_));
  AOI21_X1   g16914(.A1(new_n17015_), .A2(new_n16867_), .B(new_n17014_), .ZN(new_n17016_));
  NAND2_X1   g16915(.A1(new_n16919_), .A2(new_n16918_), .ZN(new_n17017_));
  XOR2_X1    g16916(.A1(new_n17017_), .A2(new_n16929_), .Z(new_n17018_));
  OR2_X2     g16917(.A1(new_n17018_), .A2(new_n16934_), .Z(new_n17019_));
  NAND2_X1   g16918(.A1(new_n17018_), .A2(new_n16934_), .ZN(new_n17020_));
  AOI21_X1   g16919(.A1(new_n17019_), .A2(new_n17020_), .B(new_n16922_), .ZN(new_n17021_));
  INV_X1     g16920(.I(new_n17021_), .ZN(new_n17022_));
  OAI21_X1   g16921(.A1(new_n16946_), .A2(new_n16945_), .B(new_n16779_), .ZN(new_n17023_));
  NAND2_X1   g16922(.A1(new_n17023_), .A2(new_n16761_), .ZN(new_n17024_));
  NOR3_X1    g16923(.A1(new_n16946_), .A2(new_n16945_), .A3(new_n16779_), .ZN(new_n17025_));
  NOR2_X1    g16924(.A1(new_n17025_), .A2(new_n16758_), .ZN(new_n17026_));
  NOR2_X1    g16925(.A1(new_n16577_), .A2(new_n16909_), .ZN(new_n17027_));
  INV_X1     g16926(.I(new_n17027_), .ZN(new_n17028_));
  NAND2_X1   g16927(.A1(new_n16577_), .A2(new_n16909_), .ZN(new_n17029_));
  NAND2_X1   g16928(.A1(new_n17028_), .A2(new_n17029_), .ZN(new_n17030_));
  XNOR2_X1   g16929(.A1(new_n17030_), .A2(new_n16906_), .ZN(new_n17031_));
  NAND2_X1   g16930(.A1(new_n16747_), .A2(new_n16748_), .ZN(new_n17032_));
  NAND2_X1   g16931(.A1(new_n17032_), .A2(new_n16751_), .ZN(new_n17033_));
  XOR2_X1    g16932(.A1(new_n16576_), .A2(new_n16908_), .Z(new_n17034_));
  NAND2_X1   g16933(.A1(new_n17034_), .A2(new_n16906_), .ZN(new_n17035_));
  NOR2_X1    g16934(.A1(new_n10619_), .A2(new_n511_), .ZN(new_n17036_));
  INV_X1     g16935(.I(new_n17036_), .ZN(new_n17037_));
  AOI22_X1   g16936(.A1(new_n10882_), .A2(new_n87_), .B1(new_n10875_), .B2(new_n4406_), .ZN(new_n17038_));
  AOI21_X1   g16937(.A1(new_n17037_), .A2(new_n17038_), .B(new_n82_), .ZN(new_n17039_));
  NAND2_X1   g16938(.A1(new_n13877_), .A2(new_n17039_), .ZN(new_n17040_));
  INV_X1     g16939(.I(new_n17040_), .ZN(new_n17041_));
  OAI22_X1   g16940(.A1(new_n10896_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10611_), .ZN(new_n17042_));
  OAI21_X1   g16941(.A1(new_n10606_), .A2(new_n79_), .B(new_n17042_), .ZN(new_n17043_));
  AOI21_X1   g16942(.A1(new_n17043_), .A2(new_n72_), .B(new_n79_), .ZN(new_n17044_));
  XOR2_X1    g16943(.A1(new_n12211_), .A2(new_n17044_), .Z(new_n17045_));
  NOR2_X1    g16944(.A1(new_n17045_), .A2(new_n17041_), .ZN(new_n17046_));
  XOR2_X1    g16945(.A1(new_n17027_), .A2(new_n17046_), .Z(new_n17047_));
  XOR2_X1    g16946(.A1(new_n17047_), .A2(new_n17035_), .Z(new_n17048_));
  OAI22_X1   g16947(.A1(new_n10595_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10599_), .ZN(new_n17049_));
  OAI21_X1   g16948(.A1(new_n10589_), .A2(new_n1128_), .B(new_n17049_), .ZN(new_n17050_));
  AOI21_X1   g16949(.A1(new_n17050_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n17051_));
  XOR2_X1    g16950(.A1(new_n12622_), .A2(new_n17051_), .Z(new_n17052_));
  NOR2_X1    g16951(.A1(new_n17048_), .A2(new_n17052_), .ZN(new_n17053_));
  NAND2_X1   g16952(.A1(new_n17053_), .A2(new_n17033_), .ZN(new_n17054_));
  NOR2_X1    g16953(.A1(new_n17053_), .A2(new_n17033_), .ZN(new_n17055_));
  INV_X1     g16954(.I(new_n17055_), .ZN(new_n17056_));
  AOI22_X1   g16955(.A1(new_n17056_), .A2(new_n17054_), .B1(new_n16913_), .B2(new_n17031_), .ZN(new_n17057_));
  NAND2_X1   g16956(.A1(new_n17031_), .A2(new_n16913_), .ZN(new_n17058_));
  INV_X1     g16957(.I(new_n17054_), .ZN(new_n17059_));
  NOR3_X1    g16958(.A1(new_n17059_), .A2(new_n17055_), .A3(new_n17058_), .ZN(new_n17060_));
  NOR2_X1    g16959(.A1(new_n17057_), .A2(new_n17060_), .ZN(new_n17061_));
  NOR2_X1    g16960(.A1(new_n16929_), .A2(new_n16896_), .ZN(new_n17062_));
  INV_X1     g16961(.I(new_n17062_), .ZN(new_n17063_));
  NOR2_X1    g16962(.A1(new_n16901_), .A2(new_n16934_), .ZN(new_n17064_));
  OR3_X2     g16963(.A1(new_n17064_), .A2(new_n16925_), .A3(new_n16926_), .Z(new_n17065_));
  OAI22_X1   g16964(.A1(new_n10583_), .A2(new_n1239_), .B1(new_n4981_), .B2(new_n10928_), .ZN(new_n17066_));
  AOI21_X1   g16965(.A1(new_n17066_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n17067_));
  XNOR2_X1   g16966(.A1(new_n13378_), .A2(new_n17067_), .ZN(new_n17068_));
  NAND3_X1   g16967(.A1(new_n17065_), .A2(new_n17063_), .A3(new_n17068_), .ZN(new_n17069_));
  AOI21_X1   g16968(.A1(new_n17065_), .A2(new_n17063_), .B(new_n17068_), .ZN(new_n17070_));
  INV_X1     g16969(.I(new_n17070_), .ZN(new_n17071_));
  AOI21_X1   g16970(.A1(new_n17071_), .A2(new_n17069_), .B(new_n17061_), .ZN(new_n17072_));
  INV_X1     g16971(.I(new_n17061_), .ZN(new_n17073_));
  INV_X1     g16972(.I(new_n17068_), .ZN(new_n17074_));
  AOI21_X1   g16973(.A1(new_n17065_), .A2(new_n17063_), .B(new_n17074_), .ZN(new_n17075_));
  INV_X1     g16974(.I(new_n17075_), .ZN(new_n17076_));
  NAND3_X1   g16975(.A1(new_n17065_), .A2(new_n17063_), .A3(new_n17074_), .ZN(new_n17077_));
  AOI21_X1   g16976(.A1(new_n17076_), .A2(new_n17077_), .B(new_n17073_), .ZN(new_n17078_));
  OAI22_X1   g16977(.A1(new_n4719_), .A2(new_n10938_), .B1(new_n10952_), .B2(new_n5335_), .ZN(new_n17079_));
  OAI21_X1   g16978(.A1(new_n10577_), .A2(new_n5398_), .B(new_n17079_), .ZN(new_n17080_));
  AOI21_X1   g16979(.A1(new_n17080_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n17081_));
  XOR2_X1    g16980(.A1(new_n13544_), .A2(new_n17081_), .Z(new_n17082_));
  INV_X1     g16981(.I(new_n17082_), .ZN(new_n17083_));
  OAI21_X1   g16982(.A1(new_n17078_), .A2(new_n17072_), .B(new_n17083_), .ZN(new_n17084_));
  AOI21_X1   g16983(.A1(new_n17026_), .A2(new_n17024_), .B(new_n17084_), .ZN(new_n17085_));
  AOI21_X1   g16984(.A1(new_n16938_), .A2(new_n16779_), .B(new_n16762_), .ZN(new_n17086_));
  OAI21_X1   g16985(.A1(new_n16938_), .A2(new_n16779_), .B(new_n16764_), .ZN(new_n17087_));
  INV_X1     g16986(.I(new_n17069_), .ZN(new_n17088_));
  OAI21_X1   g16987(.A1(new_n17088_), .A2(new_n17070_), .B(new_n17073_), .ZN(new_n17089_));
  AND3_X2    g16988(.A1(new_n17065_), .A2(new_n17063_), .A3(new_n17074_), .Z(new_n17090_));
  OAI21_X1   g16989(.A1(new_n17090_), .A2(new_n17075_), .B(new_n17061_), .ZN(new_n17091_));
  AOI21_X1   g16990(.A1(new_n17089_), .A2(new_n17091_), .B(new_n17082_), .ZN(new_n17092_));
  NOR3_X1    g16991(.A1(new_n17092_), .A2(new_n17086_), .A3(new_n17087_), .ZN(new_n17093_));
  OAI21_X1   g16992(.A1(new_n17085_), .A2(new_n17093_), .B(new_n17022_), .ZN(new_n17094_));
  OAI21_X1   g16993(.A1(new_n17086_), .A2(new_n17087_), .B(new_n17092_), .ZN(new_n17095_));
  NAND3_X1   g16994(.A1(new_n17084_), .A2(new_n17026_), .A3(new_n17024_), .ZN(new_n17096_));
  NAND3_X1   g16995(.A1(new_n17095_), .A2(new_n17096_), .A3(new_n17021_), .ZN(new_n17097_));
  NAND2_X1   g16996(.A1(new_n17094_), .A2(new_n17097_), .ZN(new_n17098_));
  NAND3_X1   g16997(.A1(new_n16951_), .A2(new_n16952_), .A3(new_n16963_), .ZN(new_n17099_));
  OAI22_X1   g16998(.A1(new_n10570_), .A2(new_n5419_), .B1(new_n1622_), .B2(new_n10961_), .ZN(new_n17100_));
  OAI21_X1   g16999(.A1(new_n10564_), .A2(new_n1620_), .B(new_n17100_), .ZN(new_n17101_));
  AOI21_X1   g17000(.A1(new_n17101_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n17102_));
  XOR2_X1    g17001(.A1(new_n10976_), .A2(new_n17102_), .Z(new_n17103_));
  NAND3_X1   g17002(.A1(new_n17099_), .A2(new_n16965_), .A3(new_n17103_), .ZN(new_n17104_));
  INV_X1     g17003(.I(new_n17104_), .ZN(new_n17105_));
  AOI21_X1   g17004(.A1(new_n17099_), .A2(new_n16965_), .B(new_n17103_), .ZN(new_n17106_));
  OAI21_X1   g17005(.A1(new_n17105_), .A2(new_n17106_), .B(new_n17098_), .ZN(new_n17107_));
  AOI21_X1   g17006(.A1(new_n17095_), .A2(new_n17096_), .B(new_n17021_), .ZN(new_n17108_));
  NOR3_X1    g17007(.A1(new_n17085_), .A2(new_n17093_), .A3(new_n17022_), .ZN(new_n17109_));
  NOR2_X1    g17008(.A1(new_n17109_), .A2(new_n17108_), .ZN(new_n17110_));
  INV_X1     g17009(.I(new_n17103_), .ZN(new_n17111_));
  AOI21_X1   g17010(.A1(new_n17099_), .A2(new_n16965_), .B(new_n17111_), .ZN(new_n17112_));
  NAND3_X1   g17011(.A1(new_n17099_), .A2(new_n16965_), .A3(new_n17111_), .ZN(new_n17113_));
  INV_X1     g17012(.I(new_n17113_), .ZN(new_n17114_));
  OAI21_X1   g17013(.A1(new_n17114_), .A2(new_n17112_), .B(new_n17110_), .ZN(new_n17115_));
  NAND2_X1   g17014(.A1(new_n17115_), .A2(new_n17107_), .ZN(new_n17116_));
  NOR2_X1    g17015(.A1(new_n16974_), .A2(new_n16888_), .ZN(new_n17117_));
  OAI22_X1   g17016(.A1(new_n14276_), .A2(new_n1851_), .B1(new_n5966_), .B2(new_n14594_), .ZN(new_n17118_));
  OAI21_X1   g17017(.A1(new_n14886_), .A2(new_n643_), .B(new_n17118_), .ZN(new_n17119_));
  AOI21_X1   g17018(.A1(new_n17119_), .A2(new_n279_), .B(new_n643_), .ZN(new_n17120_));
  XOR2_X1    g17019(.A1(new_n14891_), .A2(new_n17120_), .Z(new_n17121_));
  INV_X1     g17020(.I(new_n17121_), .ZN(new_n17122_));
  NOR3_X1    g17021(.A1(new_n17117_), .A2(new_n16890_), .A3(new_n17122_), .ZN(new_n17123_));
  NAND2_X1   g17022(.A1(new_n16970_), .A2(new_n16968_), .ZN(new_n17124_));
  AOI21_X1   g17023(.A1(new_n17124_), .A2(new_n16889_), .B(new_n17121_), .ZN(new_n17125_));
  OAI21_X1   g17024(.A1(new_n17123_), .A2(new_n17125_), .B(new_n17116_), .ZN(new_n17126_));
  INV_X1     g17025(.I(new_n17106_), .ZN(new_n17127_));
  AOI21_X1   g17026(.A1(new_n17127_), .A2(new_n17104_), .B(new_n17110_), .ZN(new_n17128_));
  INV_X1     g17027(.I(new_n17112_), .ZN(new_n17129_));
  AOI21_X1   g17028(.A1(new_n17129_), .A2(new_n17113_), .B(new_n17098_), .ZN(new_n17130_));
  NOR2_X1    g17029(.A1(new_n17128_), .A2(new_n17130_), .ZN(new_n17131_));
  AOI21_X1   g17030(.A1(new_n17124_), .A2(new_n16889_), .B(new_n17122_), .ZN(new_n17132_));
  NOR3_X1    g17031(.A1(new_n17117_), .A2(new_n16890_), .A3(new_n17121_), .ZN(new_n17133_));
  OAI21_X1   g17032(.A1(new_n17133_), .A2(new_n17132_), .B(new_n17131_), .ZN(new_n17134_));
  NAND2_X1   g17033(.A1(new_n17134_), .A2(new_n17126_), .ZN(new_n17135_));
  NAND2_X1   g17034(.A1(new_n16977_), .A2(new_n16877_), .ZN(new_n17136_));
  OAI22_X1   g17035(.A1(new_n16975_), .A2(new_n16969_), .B1(new_n16977_), .B2(new_n16877_), .ZN(new_n17137_));
  OAI22_X1   g17036(.A1(new_n15305_), .A2(new_n6756_), .B1(new_n15114_), .B2(new_n2258_), .ZN(new_n17138_));
  OAI21_X1   g17037(.A1(new_n1078_), .A2(new_n15515_), .B(new_n17138_), .ZN(new_n17139_));
  AOI21_X1   g17038(.A1(new_n17139_), .A2(new_n294_), .B(new_n1078_), .ZN(new_n17140_));
  XOR2_X1    g17039(.A1(new_n15518_), .A2(new_n17140_), .Z(new_n17141_));
  NAND3_X1   g17040(.A1(new_n17137_), .A2(new_n17136_), .A3(new_n17141_), .ZN(new_n17142_));
  INV_X1     g17041(.I(new_n17136_), .ZN(new_n17143_));
  AOI22_X1   g17042(.A1(new_n16882_), .A2(new_n16876_), .B1(new_n16978_), .B2(new_n16979_), .ZN(new_n17144_));
  INV_X1     g17043(.I(new_n17141_), .ZN(new_n17145_));
  OAI21_X1   g17044(.A1(new_n17144_), .A2(new_n17143_), .B(new_n17145_), .ZN(new_n17146_));
  NAND2_X1   g17045(.A1(new_n17146_), .A2(new_n17142_), .ZN(new_n17147_));
  NAND2_X1   g17046(.A1(new_n17147_), .A2(new_n17135_), .ZN(new_n17148_));
  NAND3_X1   g17047(.A1(new_n17124_), .A2(new_n16889_), .A3(new_n17121_), .ZN(new_n17149_));
  OAI21_X1   g17048(.A1(new_n17117_), .A2(new_n16890_), .B(new_n17122_), .ZN(new_n17150_));
  AOI21_X1   g17049(.A1(new_n17150_), .A2(new_n17149_), .B(new_n17131_), .ZN(new_n17151_));
  INV_X1     g17050(.I(new_n17132_), .ZN(new_n17152_));
  NAND3_X1   g17051(.A1(new_n17124_), .A2(new_n16889_), .A3(new_n17122_), .ZN(new_n17153_));
  NAND2_X1   g17052(.A1(new_n17152_), .A2(new_n17153_), .ZN(new_n17154_));
  AOI21_X1   g17053(.A1(new_n17154_), .A2(new_n17131_), .B(new_n17151_), .ZN(new_n17155_));
  AOI21_X1   g17054(.A1(new_n17137_), .A2(new_n17136_), .B(new_n17145_), .ZN(new_n17156_));
  NAND3_X1   g17055(.A1(new_n17137_), .A2(new_n17136_), .A3(new_n17145_), .ZN(new_n17157_));
  INV_X1     g17056(.I(new_n17157_), .ZN(new_n17158_));
  OAI21_X1   g17057(.A1(new_n17158_), .A2(new_n17156_), .B(new_n17155_), .ZN(new_n17159_));
  INV_X1     g17058(.I(new_n16807_), .ZN(new_n17160_));
  NAND2_X1   g17059(.A1(new_n16880_), .A2(new_n17160_), .ZN(new_n17161_));
  NAND2_X1   g17060(.A1(new_n16795_), .A2(new_n16809_), .ZN(new_n17162_));
  AOI22_X1   g17061(.A1(new_n17161_), .A2(new_n17162_), .B1(new_n16817_), .B2(new_n16820_), .ZN(new_n17163_));
  OAI21_X1   g17062(.A1(new_n17163_), .A2(new_n16822_), .B(new_n16990_), .ZN(new_n17164_));
  NOR3_X1    g17063(.A1(new_n17163_), .A2(new_n16822_), .A3(new_n16990_), .ZN(new_n17165_));
  OR3_X2     g17064(.A1(new_n16981_), .A2(new_n16984_), .A3(new_n17165_), .Z(new_n17166_));
  NAND4_X1   g17065(.A1(new_n17159_), .A2(new_n17148_), .A3(new_n17166_), .A4(new_n17164_), .ZN(new_n17167_));
  AOI22_X1   g17066(.A1(new_n17146_), .A2(new_n17142_), .B1(new_n17126_), .B2(new_n17134_), .ZN(new_n17168_));
  INV_X1     g17067(.I(new_n17156_), .ZN(new_n17169_));
  AOI21_X1   g17068(.A1(new_n17169_), .A2(new_n17157_), .B(new_n17135_), .ZN(new_n17170_));
  INV_X1     g17069(.I(new_n17164_), .ZN(new_n17171_));
  NOR3_X1    g17070(.A1(new_n16981_), .A2(new_n16984_), .A3(new_n17165_), .ZN(new_n17172_));
  OAI22_X1   g17071(.A1(new_n17170_), .A2(new_n17168_), .B1(new_n17171_), .B2(new_n17172_), .ZN(new_n17173_));
  NAND2_X1   g17072(.A1(new_n17167_), .A2(new_n17173_), .ZN(new_n17174_));
  INV_X1     g17073(.I(new_n17174_), .ZN(new_n17175_));
  NOR2_X1    g17074(.A1(new_n17003_), .A2(new_n16872_), .ZN(new_n17176_));
  NOR2_X1    g17075(.A1(new_n17007_), .A2(new_n16873_), .ZN(new_n17177_));
  NOR2_X1    g17076(.A1(new_n17176_), .A2(new_n17177_), .ZN(new_n17178_));
  NOR3_X1    g17077(.A1(new_n17178_), .A2(new_n17008_), .A3(new_n17175_), .ZN(new_n17179_));
  NOR2_X1    g17078(.A1(new_n17007_), .A2(new_n16872_), .ZN(new_n17180_));
  NOR2_X1    g17079(.A1(new_n17179_), .A2(new_n17180_), .ZN(new_n17181_));
  XOR2_X1    g17080(.A1(new_n17181_), .A2(new_n17016_), .Z(new_n17182_));
  XOR2_X1    g17081(.A1(new_n17012_), .A2(new_n17182_), .Z(\result[14] ));
  INV_X1     g17082(.I(new_n17009_), .ZN(new_n17184_));
  NOR4_X1    g17083(.A1(new_n17170_), .A2(new_n17168_), .A3(new_n17171_), .A4(new_n17172_), .ZN(new_n17185_));
  NAND3_X1   g17084(.A1(new_n17167_), .A2(new_n17007_), .A3(new_n17173_), .ZN(new_n17186_));
  AOI21_X1   g17085(.A1(new_n17167_), .A2(new_n17173_), .B(new_n17007_), .ZN(new_n17187_));
  OAI21_X1   g17086(.A1(new_n17187_), .A2(new_n16873_), .B(new_n17186_), .ZN(new_n17188_));
  NOR2_X1    g17087(.A1(new_n17048_), .A2(new_n17033_), .ZN(new_n17189_));
  NAND2_X1   g17088(.A1(new_n17048_), .A2(new_n17033_), .ZN(new_n17190_));
  NOR2_X1    g17089(.A1(new_n17058_), .A2(new_n17052_), .ZN(new_n17191_));
  AOI21_X1   g17090(.A1(new_n17191_), .A2(new_n17190_), .B(new_n17189_), .ZN(new_n17192_));
  NOR2_X1    g17091(.A1(new_n17035_), .A2(new_n17041_), .ZN(new_n17193_));
  AOI21_X1   g17092(.A1(new_n17034_), .A2(new_n16906_), .B(new_n17040_), .ZN(new_n17194_));
  NOR4_X1    g17093(.A1(new_n17194_), .A2(new_n16577_), .A3(new_n16909_), .A4(new_n17045_), .ZN(new_n17195_));
  NOR2_X1    g17094(.A1(new_n17195_), .A2(new_n17193_), .ZN(new_n17196_));
  AOI22_X1   g17095(.A1(new_n12204_), .A2(new_n4526_), .B1(new_n4570_), .B2(new_n10897_), .ZN(new_n17197_));
  AOI21_X1   g17096(.A1(new_n101_), .A2(new_n10600_), .B(new_n17197_), .ZN(new_n17198_));
  OAI21_X1   g17097(.A1(new_n17198_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n17199_));
  XNOR2_X1   g17098(.A1(new_n12576_), .A2(new_n17199_), .ZN(new_n17200_));
  NOR2_X1    g17099(.A1(new_n10619_), .A2(new_n88_), .ZN(new_n17201_));
  INV_X1     g17100(.I(new_n17201_), .ZN(new_n17202_));
  AOI22_X1   g17101(.A1(new_n10612_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n10882_), .ZN(new_n17203_));
  AOI21_X1   g17102(.A1(new_n17202_), .A2(new_n17203_), .B(new_n82_), .ZN(new_n17204_));
  NAND2_X1   g17103(.A1(new_n13894_), .A2(new_n17204_), .ZN(new_n17205_));
  XNOR2_X1   g17104(.A1(new_n17200_), .A2(new_n17205_), .ZN(new_n17206_));
  NOR2_X1    g17105(.A1(new_n17206_), .A2(new_n17040_), .ZN(new_n17207_));
  NAND2_X1   g17106(.A1(new_n17200_), .A2(new_n17205_), .ZN(new_n17208_));
  NOR2_X1    g17107(.A1(new_n17200_), .A2(new_n17205_), .ZN(new_n17209_));
  INV_X1     g17108(.I(new_n17209_), .ZN(new_n17210_));
  AOI21_X1   g17109(.A1(new_n17210_), .A2(new_n17208_), .B(new_n17041_), .ZN(new_n17211_));
  NOR2_X1    g17110(.A1(new_n17207_), .A2(new_n17211_), .ZN(new_n17212_));
  OAI22_X1   g17111(.A1(new_n10589_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10595_), .ZN(new_n17213_));
  OAI21_X1   g17112(.A1(new_n10913_), .A2(new_n1128_), .B(new_n17213_), .ZN(new_n17214_));
  AOI21_X1   g17113(.A1(new_n17214_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n17215_));
  XOR2_X1    g17114(.A1(new_n12767_), .A2(new_n17215_), .Z(new_n17216_));
  XNOR2_X1   g17115(.A1(new_n17212_), .A2(new_n17216_), .ZN(new_n17217_));
  INV_X1     g17116(.I(new_n17212_), .ZN(new_n17218_));
  INV_X1     g17117(.I(new_n17216_), .ZN(new_n17219_));
  NOR2_X1    g17118(.A1(new_n17218_), .A2(new_n17219_), .ZN(new_n17220_));
  NOR2_X1    g17119(.A1(new_n17212_), .A2(new_n17216_), .ZN(new_n17221_));
  OAI21_X1   g17120(.A1(new_n17220_), .A2(new_n17221_), .B(new_n17196_), .ZN(new_n17222_));
  OAI21_X1   g17121(.A1(new_n17196_), .A2(new_n17217_), .B(new_n17222_), .ZN(new_n17223_));
  OAI22_X1   g17122(.A1(new_n13395_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n10938_), .ZN(new_n17224_));
  AOI21_X1   g17123(.A1(new_n17224_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n17225_));
  XOR2_X1    g17124(.A1(new_n13394_), .A2(new_n17225_), .Z(new_n17226_));
  INV_X1     g17125(.I(new_n17226_), .ZN(new_n17227_));
  NOR2_X1    g17126(.A1(new_n17223_), .A2(new_n17227_), .ZN(new_n17228_));
  NAND2_X1   g17127(.A1(new_n17223_), .A2(new_n17227_), .ZN(new_n17229_));
  INV_X1     g17128(.I(new_n17229_), .ZN(new_n17230_));
  NOR2_X1    g17129(.A1(new_n17230_), .A2(new_n17228_), .ZN(new_n17231_));
  XOR2_X1    g17130(.A1(new_n17223_), .A2(new_n17227_), .Z(new_n17232_));
  NAND2_X1   g17131(.A1(new_n17232_), .A2(new_n17192_), .ZN(new_n17233_));
  OAI21_X1   g17132(.A1(new_n17192_), .A2(new_n17231_), .B(new_n17233_), .ZN(new_n17234_));
  AOI21_X1   g17133(.A1(new_n17073_), .A2(new_n17069_), .B(new_n17070_), .ZN(new_n17235_));
  OAI22_X1   g17134(.A1(new_n14054_), .A2(new_n5336_), .B1(new_n5398_), .B2(new_n10961_), .ZN(new_n17236_));
  AOI21_X1   g17135(.A1(new_n17236_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n17237_));
  XOR2_X1    g17136(.A1(new_n14053_), .A2(new_n17237_), .Z(new_n17238_));
  NAND2_X1   g17137(.A1(new_n17235_), .A2(new_n17238_), .ZN(new_n17239_));
  NOR2_X1    g17138(.A1(new_n17235_), .A2(new_n17238_), .ZN(new_n17240_));
  INV_X1     g17139(.I(new_n17240_), .ZN(new_n17241_));
  NAND2_X1   g17140(.A1(new_n17241_), .A2(new_n17239_), .ZN(new_n17242_));
  XNOR2_X1   g17141(.A1(new_n17235_), .A2(new_n17238_), .ZN(new_n17243_));
  NOR2_X1    g17142(.A1(new_n17243_), .A2(new_n17234_), .ZN(new_n17244_));
  AOI21_X1   g17143(.A1(new_n17234_), .A2(new_n17242_), .B(new_n17244_), .ZN(new_n17245_));
  NAND2_X1   g17144(.A1(new_n17026_), .A2(new_n17024_), .ZN(new_n17246_));
  NOR2_X1    g17145(.A1(new_n17078_), .A2(new_n17072_), .ZN(new_n17247_));
  NOR2_X1    g17146(.A1(new_n17246_), .A2(new_n17247_), .ZN(new_n17248_));
  NAND2_X1   g17147(.A1(new_n17246_), .A2(new_n17247_), .ZN(new_n17249_));
  NOR2_X1    g17148(.A1(new_n17022_), .A2(new_n17082_), .ZN(new_n17250_));
  AOI21_X1   g17149(.A1(new_n17249_), .A2(new_n17250_), .B(new_n17248_), .ZN(new_n17251_));
  AOI22_X1   g17150(.A1(new_n14281_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n14274_), .ZN(new_n17252_));
  OAI21_X1   g17151(.A1(new_n17252_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n17253_));
  XOR2_X1    g17152(.A1(new_n14280_), .A2(new_n17253_), .Z(new_n17254_));
  NAND2_X1   g17153(.A1(new_n17251_), .A2(new_n17254_), .ZN(new_n17255_));
  OR2_X2     g17154(.A1(new_n17251_), .A2(new_n17254_), .Z(new_n17256_));
  AOI21_X1   g17155(.A1(new_n17256_), .A2(new_n17255_), .B(new_n17245_), .ZN(new_n17257_));
  INV_X1     g17156(.I(new_n17245_), .ZN(new_n17258_));
  INV_X1     g17157(.I(new_n17254_), .ZN(new_n17259_));
  XOR2_X1    g17158(.A1(new_n17251_), .A2(new_n17259_), .Z(new_n17260_));
  NOR2_X1    g17159(.A1(new_n17260_), .A2(new_n17258_), .ZN(new_n17261_));
  NOR2_X1    g17160(.A1(new_n17261_), .A2(new_n17257_), .ZN(new_n17262_));
  AOI21_X1   g17161(.A1(new_n17098_), .A2(new_n17104_), .B(new_n17106_), .ZN(new_n17263_));
  AOI22_X1   g17162(.A1(new_n15127_), .A2(new_n5968_), .B1(new_n785_), .B2(new_n15115_), .ZN(new_n17264_));
  OAI21_X1   g17163(.A1(new_n17264_), .A2(\a[14] ), .B(new_n785_), .ZN(new_n17265_));
  XNOR2_X1   g17164(.A1(new_n15125_), .A2(new_n17265_), .ZN(new_n17266_));
  NAND2_X1   g17165(.A1(new_n17263_), .A2(new_n17266_), .ZN(new_n17267_));
  NOR2_X1    g17166(.A1(new_n17263_), .A2(new_n17266_), .ZN(new_n17268_));
  INV_X1     g17167(.I(new_n17268_), .ZN(new_n17269_));
  AOI21_X1   g17168(.A1(new_n17267_), .A2(new_n17269_), .B(new_n17262_), .ZN(new_n17270_));
  XNOR2_X1   g17169(.A1(new_n17263_), .A2(new_n17266_), .ZN(new_n17271_));
  NOR3_X1    g17170(.A1(new_n17271_), .A2(new_n17257_), .A3(new_n17261_), .ZN(new_n17272_));
  NOR2_X1    g17171(.A1(new_n17270_), .A2(new_n17272_), .ZN(new_n17273_));
  AOI21_X1   g17172(.A1(new_n17116_), .A2(new_n17149_), .B(new_n17125_), .ZN(new_n17274_));
  NAND2_X1   g17173(.A1(new_n15515_), .A2(new_n5249_), .ZN(new_n17275_));
  NOR2_X1    g17174(.A1(new_n5247_), .A2(new_n805_), .ZN(new_n17276_));
  AOI21_X1   g17175(.A1(new_n15675_), .A2(new_n17276_), .B(\a[11] ), .ZN(new_n17277_));
  AOI21_X1   g17176(.A1(new_n17277_), .A2(new_n17275_), .B(new_n1078_), .ZN(new_n17278_));
  XNOR2_X1   g17177(.A1(new_n15678_), .A2(new_n17278_), .ZN(new_n17279_));
  NAND2_X1   g17178(.A1(new_n17274_), .A2(new_n17279_), .ZN(new_n17280_));
  INV_X1     g17179(.I(new_n17280_), .ZN(new_n17281_));
  NOR2_X1    g17180(.A1(new_n17274_), .A2(new_n17279_), .ZN(new_n17282_));
  NOR2_X1    g17181(.A1(new_n17281_), .A2(new_n17282_), .ZN(new_n17283_));
  NOR2_X1    g17182(.A1(new_n17283_), .A2(new_n17273_), .ZN(new_n17284_));
  XOR2_X1    g17183(.A1(new_n17274_), .A2(new_n17279_), .Z(new_n17285_));
  AOI21_X1   g17184(.A1(new_n17273_), .A2(new_n17285_), .B(new_n17284_), .ZN(new_n17286_));
  AOI21_X1   g17185(.A1(new_n17137_), .A2(new_n17136_), .B(new_n17141_), .ZN(new_n17287_));
  AOI21_X1   g17186(.A1(new_n17135_), .A2(new_n17142_), .B(new_n17287_), .ZN(new_n17288_));
  NOR2_X1    g17187(.A1(new_n17286_), .A2(new_n17288_), .ZN(new_n17289_));
  OAI21_X1   g17188(.A1(new_n17016_), .A2(new_n17188_), .B(new_n17289_), .ZN(new_n17290_));
  AOI22_X1   g17189(.A1(new_n17159_), .A2(new_n17148_), .B1(new_n17166_), .B2(new_n17164_), .ZN(new_n17291_));
  NOR3_X1    g17190(.A1(new_n17291_), .A2(new_n17003_), .A3(new_n17185_), .ZN(new_n17292_));
  OAI21_X1   g17191(.A1(new_n17291_), .A2(new_n17185_), .B(new_n17003_), .ZN(new_n17293_));
  AOI21_X1   g17192(.A1(new_n17293_), .A2(new_n16872_), .B(new_n17292_), .ZN(new_n17294_));
  INV_X1     g17193(.I(new_n17289_), .ZN(new_n17295_));
  NAND3_X1   g17194(.A1(new_n16869_), .A2(new_n17294_), .A3(new_n17295_), .ZN(new_n17296_));
  AOI21_X1   g17195(.A1(new_n17290_), .A2(new_n17296_), .B(new_n17185_), .ZN(new_n17297_));
  AOI21_X1   g17196(.A1(new_n16869_), .A2(new_n17294_), .B(new_n17295_), .ZN(new_n17298_));
  NOR3_X1    g17197(.A1(new_n17016_), .A2(new_n17289_), .A3(new_n17188_), .ZN(new_n17299_));
  NOR3_X1    g17198(.A1(new_n17299_), .A2(new_n17298_), .A3(new_n17167_), .ZN(new_n17300_));
  NOR2_X1    g17199(.A1(new_n17300_), .A2(new_n17297_), .ZN(new_n17301_));
  NAND4_X1   g17200(.A1(\result[12] ), .A2(new_n17184_), .A3(new_n17182_), .A4(new_n17301_), .ZN(new_n17302_));
  AOI21_X1   g17201(.A1(new_n16510_), .A2(new_n16712_), .B(new_n16860_), .ZN(new_n17303_));
  NOR3_X1    g17202(.A1(new_n16717_), .A2(new_n16718_), .A3(new_n16858_), .ZN(new_n17304_));
  OAI21_X1   g17203(.A1(new_n17304_), .A2(new_n17303_), .B(new_n17184_), .ZN(new_n17305_));
  XOR2_X1    g17204(.A1(new_n17181_), .A2(new_n16869_), .Z(new_n17306_));
  OAI21_X1   g17205(.A1(new_n17299_), .A2(new_n17298_), .B(new_n17167_), .ZN(new_n17307_));
  NAND3_X1   g17206(.A1(new_n17290_), .A2(new_n17296_), .A3(new_n17185_), .ZN(new_n17308_));
  NAND2_X1   g17207(.A1(new_n17307_), .A2(new_n17308_), .ZN(new_n17309_));
  OAI21_X1   g17208(.A1(new_n17305_), .A2(new_n17306_), .B(new_n17309_), .ZN(new_n17310_));
  NAND2_X1   g17209(.A1(new_n17310_), .A2(new_n17302_), .ZN(\result[15] ));
  NAND2_X1   g17210(.A1(new_n17012_), .A2(new_n17182_), .ZN(new_n17312_));
  NAND2_X1   g17211(.A1(new_n16869_), .A2(new_n17294_), .ZN(new_n17313_));
  AOI21_X1   g17212(.A1(new_n17286_), .A2(new_n17167_), .B(new_n17288_), .ZN(new_n17314_));
  INV_X1     g17213(.I(new_n17314_), .ZN(new_n17315_));
  OAI22_X1   g17214(.A1(new_n17313_), .A2(new_n17315_), .B1(new_n17167_), .B2(new_n17286_), .ZN(new_n17316_));
  NOR2_X1    g17215(.A1(new_n17273_), .A2(new_n17281_), .ZN(new_n17317_));
  NOR2_X1    g17216(.A1(new_n17317_), .A2(new_n17282_), .ZN(new_n17318_));
  INV_X1     g17217(.I(new_n17318_), .ZN(new_n17319_));
  AOI22_X1   g17218(.A1(new_n14602_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n14603_), .ZN(new_n17320_));
  OAI21_X1   g17219(.A1(new_n17320_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n17321_));
  XNOR2_X1   g17220(.A1(new_n14601_), .A2(new_n17321_), .ZN(new_n17322_));
  INV_X1     g17221(.I(new_n17322_), .ZN(new_n17323_));
  NAND2_X1   g17222(.A1(new_n17255_), .A2(new_n17258_), .ZN(new_n17324_));
  NAND2_X1   g17223(.A1(new_n17324_), .A2(new_n17256_), .ZN(new_n17325_));
  AOI21_X1   g17224(.A1(new_n17234_), .A2(new_n17239_), .B(new_n17240_), .ZN(new_n17326_));
  OAI22_X1   g17225(.A1(new_n10965_), .A2(new_n5336_), .B1(new_n5398_), .B2(new_n10570_), .ZN(new_n17327_));
  AOI21_X1   g17226(.A1(new_n17327_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n17328_));
  XNOR2_X1   g17227(.A1(new_n14077_), .A2(new_n17328_), .ZN(new_n17329_));
  NAND2_X1   g17228(.A1(new_n17326_), .A2(new_n17329_), .ZN(new_n17330_));
  NOR2_X1    g17229(.A1(new_n17326_), .A2(new_n17329_), .ZN(new_n17331_));
  INV_X1     g17230(.I(new_n17331_), .ZN(new_n17332_));
  NAND2_X1   g17231(.A1(new_n17332_), .A2(new_n17330_), .ZN(new_n17333_));
  OAI21_X1   g17232(.A1(new_n17192_), .A2(new_n17228_), .B(new_n17229_), .ZN(new_n17334_));
  INV_X1     g17233(.I(new_n17334_), .ZN(new_n17335_));
  INV_X1     g17234(.I(new_n17217_), .ZN(new_n17336_));
  OAI22_X1   g17235(.A1(new_n10606_), .A2(new_n4529_), .B1(new_n4527_), .B2(new_n10599_), .ZN(new_n17337_));
  OAI21_X1   g17236(.A1(new_n10595_), .A2(new_n79_), .B(new_n17337_), .ZN(new_n17338_));
  AOI21_X1   g17237(.A1(new_n17338_), .A2(new_n72_), .B(new_n79_), .ZN(new_n17339_));
  XOR2_X1    g17238(.A1(new_n12600_), .A2(new_n17339_), .Z(new_n17340_));
  INV_X1     g17239(.I(new_n17340_), .ZN(new_n17341_));
  OAI21_X1   g17240(.A1(new_n15515_), .A2(new_n5250_), .B(new_n294_), .ZN(new_n17342_));
  OAI21_X1   g17241(.A1(new_n5252_), .A2(new_n15515_), .B(new_n17342_), .ZN(new_n17343_));
  NOR2_X1    g17242(.A1(new_n10611_), .A2(new_n88_), .ZN(new_n17344_));
  INV_X1     g17243(.I(new_n17344_), .ZN(new_n17345_));
  AOI22_X1   g17244(.A1(new_n10620_), .A2(new_n4406_), .B1(new_n962_), .B2(new_n10897_), .ZN(new_n17346_));
  AOI21_X1   g17245(.A1(new_n17346_), .A2(new_n17345_), .B(new_n82_), .ZN(new_n17347_));
  AOI21_X1   g17246(.A1(new_n10984_), .A2(new_n17347_), .B(new_n17343_), .ZN(new_n17348_));
  INV_X1     g17247(.I(new_n17343_), .ZN(new_n17349_));
  NAND2_X1   g17248(.A1(new_n10984_), .A2(new_n17347_), .ZN(new_n17350_));
  NOR2_X1    g17249(.A1(new_n17349_), .A2(new_n17350_), .ZN(new_n17351_));
  NOR2_X1    g17250(.A1(new_n17351_), .A2(new_n17348_), .ZN(new_n17352_));
  AOI21_X1   g17251(.A1(new_n17041_), .A2(new_n17208_), .B(new_n17209_), .ZN(new_n17353_));
  AOI22_X1   g17252(.A1(new_n10914_), .A2(new_n4767_), .B1(new_n4613_), .B2(new_n12616_), .ZN(new_n17354_));
  AOI21_X1   g17253(.A1(new_n117_), .A2(new_n10924_), .B(new_n17354_), .ZN(new_n17355_));
  OAI21_X1   g17254(.A1(new_n17355_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n17356_));
  XOR2_X1    g17255(.A1(new_n12889_), .A2(new_n17356_), .Z(new_n17357_));
  XOR2_X1    g17256(.A1(new_n17357_), .A2(new_n17353_), .Z(new_n17358_));
  XOR2_X1    g17257(.A1(new_n17358_), .A2(new_n17352_), .Z(new_n17359_));
  XOR2_X1    g17258(.A1(new_n17359_), .A2(new_n17341_), .Z(new_n17360_));
  NAND2_X1   g17259(.A1(new_n17360_), .A2(new_n17336_), .ZN(new_n17361_));
  XNOR2_X1   g17260(.A1(new_n17361_), .A2(new_n17221_), .ZN(new_n17362_));
  XOR2_X1    g17261(.A1(new_n17362_), .A2(new_n17196_), .Z(new_n17363_));
  OAI22_X1   g17262(.A1(new_n12908_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n10952_), .ZN(new_n17364_));
  AOI21_X1   g17263(.A1(new_n17364_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n17365_));
  XNOR2_X1   g17264(.A1(new_n12907_), .A2(new_n17365_), .ZN(new_n17366_));
  XOR2_X1    g17265(.A1(new_n17363_), .A2(new_n17366_), .Z(new_n17367_));
  INV_X1     g17266(.I(new_n17366_), .ZN(new_n17368_));
  NOR2_X1    g17267(.A1(new_n17363_), .A2(new_n17368_), .ZN(new_n17369_));
  AND2_X2    g17268(.A1(new_n17363_), .A2(new_n17368_), .Z(new_n17370_));
  NOR2_X1    g17269(.A1(new_n17370_), .A2(new_n17369_), .ZN(new_n17371_));
  MUX2_X1    g17270(.I0(new_n17367_), .I1(new_n17371_), .S(new_n17335_), .Z(new_n17372_));
  XOR2_X1    g17271(.A1(new_n17372_), .A2(new_n17333_), .Z(new_n17373_));
  NOR2_X1    g17272(.A1(new_n17373_), .A2(new_n17325_), .ZN(new_n17374_));
  INV_X1     g17273(.I(new_n17374_), .ZN(new_n17375_));
  NAND2_X1   g17274(.A1(new_n17373_), .A2(new_n17325_), .ZN(new_n17376_));
  AOI21_X1   g17275(.A1(new_n17375_), .A2(new_n17376_), .B(new_n17323_), .ZN(new_n17377_));
  INV_X1     g17276(.I(new_n17376_), .ZN(new_n17378_));
  NOR3_X1    g17277(.A1(new_n17378_), .A2(new_n17322_), .A3(new_n17374_), .ZN(new_n17379_));
  NOR2_X1    g17278(.A1(new_n17377_), .A2(new_n17379_), .ZN(new_n17380_));
  INV_X1     g17279(.I(new_n17380_), .ZN(new_n17381_));
  AOI21_X1   g17280(.A1(new_n17263_), .A2(new_n17266_), .B(new_n17262_), .ZN(new_n17382_));
  NOR2_X1    g17281(.A1(new_n17382_), .A2(new_n17268_), .ZN(new_n17383_));
  OAI22_X1   g17282(.A1(new_n15313_), .A2(new_n5967_), .B1(new_n643_), .B2(new_n15305_), .ZN(new_n17384_));
  AOI21_X1   g17283(.A1(new_n17384_), .A2(new_n279_), .B(new_n643_), .ZN(new_n17385_));
  XNOR2_X1   g17284(.A1(new_n15312_), .A2(new_n17385_), .ZN(new_n17386_));
  NAND2_X1   g17285(.A1(new_n17383_), .A2(new_n17386_), .ZN(new_n17387_));
  INV_X1     g17286(.I(new_n17387_), .ZN(new_n17388_));
  NOR2_X1    g17287(.A1(new_n17383_), .A2(new_n17386_), .ZN(new_n17389_));
  OAI21_X1   g17288(.A1(new_n17388_), .A2(new_n17389_), .B(new_n17381_), .ZN(new_n17390_));
  INV_X1     g17289(.I(new_n17386_), .ZN(new_n17391_));
  NOR2_X1    g17290(.A1(new_n17383_), .A2(new_n17391_), .ZN(new_n17392_));
  NAND2_X1   g17291(.A1(new_n17383_), .A2(new_n17391_), .ZN(new_n17393_));
  INV_X1     g17292(.I(new_n17393_), .ZN(new_n17394_));
  OAI21_X1   g17293(.A1(new_n17394_), .A2(new_n17392_), .B(new_n17380_), .ZN(new_n17395_));
  NAND2_X1   g17294(.A1(new_n17390_), .A2(new_n17395_), .ZN(new_n17396_));
  NOR2_X1    g17295(.A1(new_n17396_), .A2(new_n17319_), .ZN(new_n17397_));
  INV_X1     g17296(.I(new_n17389_), .ZN(new_n17398_));
  AOI21_X1   g17297(.A1(new_n17398_), .A2(new_n17387_), .B(new_n17380_), .ZN(new_n17399_));
  OR2_X2     g17298(.A1(new_n17382_), .A2(new_n17268_), .Z(new_n17400_));
  NAND2_X1   g17299(.A1(new_n17400_), .A2(new_n17386_), .ZN(new_n17401_));
  AOI21_X1   g17300(.A1(new_n17401_), .A2(new_n17393_), .B(new_n17381_), .ZN(new_n17402_));
  NOR2_X1    g17301(.A1(new_n17399_), .A2(new_n17402_), .ZN(new_n17403_));
  NOR2_X1    g17302(.A1(new_n17403_), .A2(new_n17318_), .ZN(new_n17404_));
  OAI21_X1   g17303(.A1(new_n17397_), .A2(new_n17404_), .B(new_n17316_), .ZN(new_n17405_));
  XOR2_X1    g17304(.A1(new_n17405_), .A2(new_n17309_), .Z(new_n17406_));
  XOR2_X1    g17305(.A1(new_n17406_), .A2(new_n17312_), .Z(\result[16] ));
  AOI21_X1   g17306(.A1(new_n17310_), .A2(new_n17302_), .B(new_n17405_), .ZN(new_n17408_));
  NOR2_X1    g17307(.A1(new_n17016_), .A2(new_n17188_), .ZN(new_n17409_));
  NOR2_X1    g17308(.A1(new_n17286_), .A2(new_n17167_), .ZN(new_n17410_));
  AOI21_X1   g17309(.A1(new_n17409_), .A2(new_n17314_), .B(new_n17410_), .ZN(new_n17411_));
  INV_X1     g17310(.I(new_n17369_), .ZN(new_n17412_));
  AOI21_X1   g17311(.A1(new_n17334_), .A2(new_n17412_), .B(new_n17370_), .ZN(new_n17413_));
  INV_X1     g17312(.I(new_n17357_), .ZN(new_n17414_));
  XNOR2_X1   g17313(.A1(new_n17352_), .A2(new_n17353_), .ZN(new_n17415_));
  OR2_X2     g17314(.A1(new_n17415_), .A2(new_n17341_), .Z(new_n17416_));
  NAND2_X1   g17315(.A1(new_n17415_), .A2(new_n17341_), .ZN(new_n17417_));
  AOI21_X1   g17316(.A1(new_n17416_), .A2(new_n17417_), .B(new_n17414_), .ZN(new_n17418_));
  AOI21_X1   g17317(.A1(new_n17360_), .A2(new_n17218_), .B(new_n17219_), .ZN(new_n17419_));
  NOR2_X1    g17318(.A1(new_n17360_), .A2(new_n17218_), .ZN(new_n17420_));
  NOR3_X1    g17319(.A1(new_n17419_), .A2(new_n17420_), .A3(new_n17196_), .ZN(new_n17421_));
  NAND2_X1   g17320(.A1(new_n17352_), .A2(new_n17353_), .ZN(new_n17422_));
  INV_X1     g17321(.I(new_n17422_), .ZN(new_n17423_));
  NOR2_X1    g17322(.A1(new_n17343_), .A2(new_n17350_), .ZN(new_n17424_));
  INV_X1     g17323(.I(new_n17424_), .ZN(new_n17425_));
  NOR2_X1    g17324(.A1(new_n10606_), .A2(new_n511_), .ZN(new_n17426_));
  INV_X1     g17325(.I(new_n17426_), .ZN(new_n17427_));
  AOI22_X1   g17326(.A1(new_n10897_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n10612_), .ZN(new_n17428_));
  AOI21_X1   g17327(.A1(new_n17427_), .A2(new_n17428_), .B(new_n82_), .ZN(new_n17429_));
  OAI21_X1   g17328(.A1(new_n12209_), .A2(new_n12210_), .B(new_n17429_), .ZN(new_n17430_));
  OAI22_X1   g17329(.A1(new_n10595_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10599_), .ZN(new_n17431_));
  OAI21_X1   g17330(.A1(new_n10589_), .A2(new_n79_), .B(new_n17431_), .ZN(new_n17432_));
  AOI21_X1   g17331(.A1(new_n17432_), .A2(new_n72_), .B(new_n79_), .ZN(new_n17433_));
  XOR2_X1    g17332(.A1(new_n12622_), .A2(new_n17433_), .Z(new_n17434_));
  XOR2_X1    g17333(.A1(new_n17434_), .A2(new_n17430_), .Z(new_n17435_));
  NOR2_X1    g17334(.A1(new_n17435_), .A2(new_n17425_), .ZN(new_n17436_));
  INV_X1     g17335(.I(new_n17430_), .ZN(new_n17437_));
  NAND2_X1   g17336(.A1(new_n17434_), .A2(new_n17437_), .ZN(new_n17438_));
  NOR2_X1    g17337(.A1(new_n17434_), .A2(new_n17437_), .ZN(new_n17439_));
  INV_X1     g17338(.I(new_n17439_), .ZN(new_n17440_));
  AOI21_X1   g17339(.A1(new_n17440_), .A2(new_n17438_), .B(new_n17424_), .ZN(new_n17441_));
  OAI22_X1   g17340(.A1(new_n10923_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10913_), .ZN(new_n17442_));
  OAI21_X1   g17341(.A1(new_n10583_), .A2(new_n1128_), .B(new_n17442_), .ZN(new_n17443_));
  AOI21_X1   g17342(.A1(new_n17443_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n17444_));
  XOR2_X1    g17343(.A1(new_n13378_), .A2(new_n17444_), .Z(new_n17445_));
  OAI21_X1   g17344(.A1(new_n17436_), .A2(new_n17441_), .B(new_n17445_), .ZN(new_n17446_));
  XOR2_X1    g17345(.A1(new_n17446_), .A2(new_n17423_), .Z(new_n17447_));
  XNOR2_X1   g17346(.A1(new_n17447_), .A2(new_n17416_), .ZN(new_n17448_));
  OAI22_X1   g17347(.A1(new_n1973_), .A2(new_n10938_), .B1(new_n10952_), .B2(new_n4902_), .ZN(new_n17449_));
  OAI21_X1   g17348(.A1(new_n10577_), .A2(new_n1239_), .B(new_n17449_), .ZN(new_n17450_));
  AOI21_X1   g17349(.A1(new_n17450_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n17451_));
  XOR2_X1    g17350(.A1(new_n13544_), .A2(new_n17451_), .Z(new_n17452_));
  NOR2_X1    g17351(.A1(new_n17448_), .A2(new_n17452_), .ZN(new_n17453_));
  XNOR2_X1   g17352(.A1(new_n17421_), .A2(new_n17453_), .ZN(new_n17454_));
  XOR2_X1    g17353(.A1(new_n17454_), .A2(new_n17418_), .Z(new_n17455_));
  OAI22_X1   g17354(.A1(new_n10570_), .A2(new_n5335_), .B1(new_n4719_), .B2(new_n10961_), .ZN(new_n17456_));
  OAI21_X1   g17355(.A1(new_n10564_), .A2(new_n5398_), .B(new_n17456_), .ZN(new_n17457_));
  AOI21_X1   g17356(.A1(new_n17457_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n17458_));
  XOR2_X1    g17357(.A1(new_n10976_), .A2(new_n17458_), .Z(new_n17459_));
  AND2_X2    g17358(.A1(new_n17455_), .A2(new_n17459_), .Z(new_n17460_));
  NOR2_X1    g17359(.A1(new_n17455_), .A2(new_n17459_), .ZN(new_n17461_));
  NOR2_X1    g17360(.A1(new_n17460_), .A2(new_n17461_), .ZN(new_n17462_));
  NOR2_X1    g17361(.A1(new_n17462_), .A2(new_n17413_), .ZN(new_n17463_));
  INV_X1     g17362(.I(new_n17413_), .ZN(new_n17464_));
  XNOR2_X1   g17363(.A1(new_n17455_), .A2(new_n17459_), .ZN(new_n17465_));
  NOR2_X1    g17364(.A1(new_n17465_), .A2(new_n17464_), .ZN(new_n17466_));
  NOR2_X1    g17365(.A1(new_n17466_), .A2(new_n17463_), .ZN(new_n17467_));
  AND2_X2    g17366(.A1(new_n17372_), .A2(new_n17330_), .Z(new_n17468_));
  NOR2_X1    g17367(.A1(new_n17468_), .A2(new_n17331_), .ZN(new_n17469_));
  OAI22_X1   g17368(.A1(new_n14276_), .A2(new_n1622_), .B1(new_n5419_), .B2(new_n14594_), .ZN(new_n17470_));
  OAI21_X1   g17369(.A1(new_n14886_), .A2(new_n1620_), .B(new_n17470_), .ZN(new_n17471_));
  AOI21_X1   g17370(.A1(new_n17471_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n17472_));
  XOR2_X1    g17371(.A1(new_n14891_), .A2(new_n17472_), .Z(new_n17473_));
  NAND2_X1   g17372(.A1(new_n17469_), .A2(new_n17473_), .ZN(new_n17474_));
  NOR2_X1    g17373(.A1(new_n17469_), .A2(new_n17473_), .ZN(new_n17475_));
  INV_X1     g17374(.I(new_n17475_), .ZN(new_n17476_));
  AOI21_X1   g17375(.A1(new_n17476_), .A2(new_n17474_), .B(new_n17467_), .ZN(new_n17477_));
  XOR2_X1    g17376(.A1(new_n17469_), .A2(new_n17473_), .Z(new_n17478_));
  AOI21_X1   g17377(.A1(new_n17478_), .A2(new_n17467_), .B(new_n17477_), .ZN(new_n17479_));
  NAND2_X1   g17378(.A1(new_n17325_), .A2(new_n17323_), .ZN(new_n17480_));
  INV_X1     g17379(.I(new_n17373_), .ZN(new_n17481_));
  OAI21_X1   g17380(.A1(new_n17325_), .A2(new_n17323_), .B(new_n17481_), .ZN(new_n17482_));
  OAI22_X1   g17381(.A1(new_n15305_), .A2(new_n5966_), .B1(new_n15114_), .B2(new_n1851_), .ZN(new_n17483_));
  OAI21_X1   g17382(.A1(new_n643_), .A2(new_n15515_), .B(new_n17483_), .ZN(new_n17484_));
  AOI21_X1   g17383(.A1(new_n17484_), .A2(new_n279_), .B(new_n643_), .ZN(new_n17485_));
  XOR2_X1    g17384(.A1(new_n15518_), .A2(new_n17485_), .Z(new_n17486_));
  NAND3_X1   g17385(.A1(new_n17482_), .A2(new_n17480_), .A3(new_n17486_), .ZN(new_n17487_));
  NAND2_X1   g17386(.A1(new_n17482_), .A2(new_n17480_), .ZN(new_n17488_));
  INV_X1     g17387(.I(new_n17486_), .ZN(new_n17489_));
  NAND2_X1   g17388(.A1(new_n17488_), .A2(new_n17489_), .ZN(new_n17490_));
  AOI21_X1   g17389(.A1(new_n17490_), .A2(new_n17487_), .B(new_n17479_), .ZN(new_n17491_));
  NAND2_X1   g17390(.A1(new_n17488_), .A2(new_n17486_), .ZN(new_n17492_));
  NAND3_X1   g17391(.A1(new_n17482_), .A2(new_n17480_), .A3(new_n17489_), .ZN(new_n17493_));
  NAND2_X1   g17392(.A1(new_n17492_), .A2(new_n17493_), .ZN(new_n17494_));
  NAND2_X1   g17393(.A1(new_n17494_), .A2(new_n17479_), .ZN(new_n17495_));
  INV_X1     g17394(.I(new_n17495_), .ZN(new_n17496_));
  NAND2_X1   g17395(.A1(new_n17387_), .A2(new_n17380_), .ZN(new_n17497_));
  INV_X1     g17396(.I(new_n17497_), .ZN(new_n17498_));
  NOR4_X1    g17397(.A1(new_n17496_), .A2(new_n17498_), .A3(new_n17389_), .A4(new_n17491_), .ZN(new_n17499_));
  INV_X1     g17398(.I(new_n17479_), .ZN(new_n17500_));
  NAND2_X1   g17399(.A1(new_n17490_), .A2(new_n17487_), .ZN(new_n17501_));
  NAND2_X1   g17400(.A1(new_n17500_), .A2(new_n17501_), .ZN(new_n17502_));
  AOI22_X1   g17401(.A1(new_n17502_), .A2(new_n17495_), .B1(new_n17398_), .B2(new_n17497_), .ZN(new_n17503_));
  NOR2_X1    g17402(.A1(new_n17499_), .A2(new_n17503_), .ZN(new_n17504_));
  XOR2_X1    g17403(.A1(new_n17403_), .A2(new_n17319_), .Z(new_n17505_));
  NOR3_X1    g17404(.A1(new_n17505_), .A2(new_n17404_), .A3(new_n17504_), .ZN(new_n17506_));
  NOR2_X1    g17405(.A1(new_n17403_), .A2(new_n17318_), .ZN(new_n17507_));
  NOR2_X1    g17406(.A1(new_n17506_), .A2(new_n17507_), .ZN(new_n17508_));
  XOR2_X1    g17407(.A1(new_n17508_), .A2(new_n17411_), .Z(new_n17509_));
  XOR2_X1    g17408(.A1(new_n17408_), .A2(new_n17509_), .Z(\result[17] ));
  NOR3_X1    g17409(.A1(new_n17305_), .A2(new_n17306_), .A3(new_n17309_), .ZN(new_n17511_));
  AOI21_X1   g17410(.A1(new_n17012_), .A2(new_n17182_), .B(new_n17301_), .ZN(new_n17512_));
  INV_X1     g17411(.I(new_n17405_), .ZN(new_n17513_));
  OAI21_X1   g17412(.A1(new_n17511_), .A2(new_n17512_), .B(new_n17513_), .ZN(new_n17514_));
  XOR2_X1    g17413(.A1(new_n17508_), .A2(new_n17316_), .Z(new_n17515_));
  NAND4_X1   g17414(.A1(new_n17502_), .A2(new_n17495_), .A3(new_n17398_), .A4(new_n17497_), .ZN(new_n17516_));
  OAI22_X1   g17415(.A1(new_n17496_), .A2(new_n17491_), .B1(new_n17498_), .B2(new_n17389_), .ZN(new_n17517_));
  NAND3_X1   g17416(.A1(new_n17517_), .A2(new_n17403_), .A3(new_n17516_), .ZN(new_n17518_));
  AOI21_X1   g17417(.A1(new_n17517_), .A2(new_n17516_), .B(new_n17403_), .ZN(new_n17519_));
  OAI21_X1   g17418(.A1(new_n17519_), .A2(new_n17319_), .B(new_n17518_), .ZN(new_n17520_));
  INV_X1     g17419(.I(new_n17460_), .ZN(new_n17521_));
  AOI21_X1   g17420(.A1(new_n17464_), .A2(new_n17521_), .B(new_n17461_), .ZN(new_n17522_));
  INV_X1     g17421(.I(new_n17522_), .ZN(new_n17523_));
  AOI21_X1   g17422(.A1(new_n17434_), .A2(new_n17437_), .B(new_n17425_), .ZN(new_n17524_));
  NOR2_X1    g17423(.A1(new_n17524_), .A2(new_n17439_), .ZN(new_n17525_));
  NOR2_X1    g17424(.A1(new_n10606_), .A2(new_n88_), .ZN(new_n17526_));
  INV_X1     g17425(.I(new_n17526_), .ZN(new_n17527_));
  AOI22_X1   g17426(.A1(new_n10600_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n10897_), .ZN(new_n17528_));
  AOI21_X1   g17427(.A1(new_n17527_), .A2(new_n17528_), .B(new_n82_), .ZN(new_n17529_));
  NAND2_X1   g17428(.A1(new_n14188_), .A2(new_n17529_), .ZN(new_n17530_));
  XOR2_X1    g17429(.A1(new_n17530_), .A2(new_n17430_), .Z(new_n17531_));
  NOR2_X1    g17430(.A1(new_n17530_), .A2(new_n17437_), .ZN(new_n17532_));
  INV_X1     g17431(.I(new_n17530_), .ZN(new_n17533_));
  NOR2_X1    g17432(.A1(new_n17533_), .A2(new_n17430_), .ZN(new_n17534_));
  OAI21_X1   g17433(.A1(new_n17532_), .A2(new_n17534_), .B(new_n17525_), .ZN(new_n17535_));
  OAI21_X1   g17434(.A1(new_n17525_), .A2(new_n17531_), .B(new_n17535_), .ZN(new_n17536_));
  OAI22_X1   g17435(.A1(new_n10583_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10923_), .ZN(new_n17537_));
  OAI21_X1   g17436(.A1(new_n1128_), .A2(new_n10938_), .B(new_n17537_), .ZN(new_n17538_));
  AOI21_X1   g17437(.A1(new_n17538_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n17539_));
  XOR2_X1    g17438(.A1(new_n13394_), .A2(new_n17539_), .Z(new_n17540_));
  OAI22_X1   g17439(.A1(new_n10589_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10595_), .ZN(new_n17541_));
  OAI21_X1   g17440(.A1(new_n10913_), .A2(new_n79_), .B(new_n17541_), .ZN(new_n17542_));
  AOI21_X1   g17441(.A1(new_n17542_), .A2(new_n72_), .B(new_n79_), .ZN(new_n17543_));
  XOR2_X1    g17442(.A1(new_n12767_), .A2(new_n17543_), .Z(new_n17544_));
  XNOR2_X1   g17443(.A1(new_n17540_), .A2(new_n17544_), .ZN(new_n17545_));
  INV_X1     g17444(.I(new_n17545_), .ZN(new_n17546_));
  NAND2_X1   g17445(.A1(new_n17540_), .A2(new_n17544_), .ZN(new_n17547_));
  INV_X1     g17446(.I(new_n17547_), .ZN(new_n17548_));
  NOR2_X1    g17447(.A1(new_n17540_), .A2(new_n17544_), .ZN(new_n17549_));
  NOR2_X1    g17448(.A1(new_n17548_), .A2(new_n17549_), .ZN(new_n17550_));
  NOR2_X1    g17449(.A1(new_n17550_), .A2(new_n17536_), .ZN(new_n17551_));
  AOI21_X1   g17450(.A1(new_n17536_), .A2(new_n17546_), .B(new_n17551_), .ZN(new_n17552_));
  NOR2_X1    g17451(.A1(new_n17436_), .A2(new_n17441_), .ZN(new_n17553_));
  NOR2_X1    g17452(.A1(new_n17416_), .A2(new_n17553_), .ZN(new_n17554_));
  NAND2_X1   g17453(.A1(new_n17423_), .A2(new_n17445_), .ZN(new_n17555_));
  AOI21_X1   g17454(.A1(new_n17416_), .A2(new_n17553_), .B(new_n17555_), .ZN(new_n17556_));
  NOR2_X1    g17455(.A1(new_n17556_), .A2(new_n17554_), .ZN(new_n17557_));
  OAI22_X1   g17456(.A1(new_n14054_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n10961_), .ZN(new_n17558_));
  AOI21_X1   g17457(.A1(new_n17558_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n17559_));
  XOR2_X1    g17458(.A1(new_n14053_), .A2(new_n17559_), .Z(new_n17560_));
  AND2_X2    g17459(.A1(new_n17560_), .A2(new_n17557_), .Z(new_n17561_));
  NOR2_X1    g17460(.A1(new_n17560_), .A2(new_n17557_), .ZN(new_n17562_));
  NOR2_X1    g17461(.A1(new_n17561_), .A2(new_n17562_), .ZN(new_n17563_));
  NOR2_X1    g17462(.A1(new_n17563_), .A2(new_n17552_), .ZN(new_n17564_));
  XNOR2_X1   g17463(.A1(new_n17560_), .A2(new_n17557_), .ZN(new_n17565_));
  INV_X1     g17464(.I(new_n17565_), .ZN(new_n17566_));
  AOI21_X1   g17465(.A1(new_n17552_), .A2(new_n17566_), .B(new_n17564_), .ZN(new_n17567_));
  INV_X1     g17466(.I(new_n17448_), .ZN(new_n17568_));
  NAND2_X1   g17467(.A1(new_n17421_), .A2(new_n17568_), .ZN(new_n17569_));
  INV_X1     g17468(.I(new_n17418_), .ZN(new_n17570_));
  NOR2_X1    g17469(.A1(new_n17570_), .A2(new_n17452_), .ZN(new_n17571_));
  OAI21_X1   g17470(.A1(new_n17421_), .A2(new_n17568_), .B(new_n17571_), .ZN(new_n17572_));
  NAND2_X1   g17471(.A1(new_n17572_), .A2(new_n17569_), .ZN(new_n17573_));
  AOI22_X1   g17472(.A1(new_n14281_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n14274_), .ZN(new_n17574_));
  OAI21_X1   g17473(.A1(new_n17574_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n17575_));
  XOR2_X1    g17474(.A1(new_n14280_), .A2(new_n17575_), .Z(new_n17576_));
  INV_X1     g17475(.I(new_n17576_), .ZN(new_n17577_));
  NOR2_X1    g17476(.A1(new_n17573_), .A2(new_n17577_), .ZN(new_n17578_));
  INV_X1     g17477(.I(new_n17578_), .ZN(new_n17579_));
  NAND2_X1   g17478(.A1(new_n17573_), .A2(new_n17577_), .ZN(new_n17580_));
  AOI21_X1   g17479(.A1(new_n17579_), .A2(new_n17580_), .B(new_n17567_), .ZN(new_n17581_));
  INV_X1     g17480(.I(new_n17567_), .ZN(new_n17582_));
  XOR2_X1    g17481(.A1(new_n17573_), .A2(new_n17576_), .Z(new_n17583_));
  NOR2_X1    g17482(.A1(new_n17583_), .A2(new_n17582_), .ZN(new_n17584_));
  AOI22_X1   g17483(.A1(new_n15127_), .A2(new_n5421_), .B1(new_n4660_), .B2(new_n15115_), .ZN(new_n17585_));
  OAI21_X1   g17484(.A1(new_n17585_), .A2(\a[17] ), .B(new_n4660_), .ZN(new_n17586_));
  XNOR2_X1   g17485(.A1(new_n15125_), .A2(new_n17586_), .ZN(new_n17587_));
  INV_X1     g17486(.I(new_n17587_), .ZN(new_n17588_));
  NOR3_X1    g17487(.A1(new_n17584_), .A2(new_n17581_), .A3(new_n17588_), .ZN(new_n17589_));
  NOR2_X1    g17488(.A1(new_n17584_), .A2(new_n17581_), .ZN(new_n17590_));
  NOR2_X1    g17489(.A1(new_n17590_), .A2(new_n17587_), .ZN(new_n17591_));
  OAI21_X1   g17490(.A1(new_n17589_), .A2(new_n17591_), .B(new_n17523_), .ZN(new_n17592_));
  XOR2_X1    g17491(.A1(new_n17590_), .A2(new_n17588_), .Z(new_n17593_));
  OAI21_X1   g17492(.A1(new_n17593_), .A2(new_n17523_), .B(new_n17592_), .ZN(new_n17594_));
  INV_X1     g17493(.I(new_n17474_), .ZN(new_n17595_));
  OAI21_X1   g17494(.A1(new_n17467_), .A2(new_n17595_), .B(new_n17476_), .ZN(new_n17596_));
  NAND2_X1   g17495(.A1(new_n15515_), .A2(new_n4943_), .ZN(new_n17597_));
  NOR2_X1    g17496(.A1(new_n4941_), .A2(new_n785_), .ZN(new_n17598_));
  AOI21_X1   g17497(.A1(new_n15675_), .A2(new_n17598_), .B(\a[14] ), .ZN(new_n17599_));
  AOI21_X1   g17498(.A1(new_n17599_), .A2(new_n17597_), .B(new_n643_), .ZN(new_n17600_));
  XNOR2_X1   g17499(.A1(new_n15678_), .A2(new_n17600_), .ZN(new_n17601_));
  INV_X1     g17500(.I(new_n17601_), .ZN(new_n17602_));
  OR2_X2     g17501(.A1(new_n17596_), .A2(new_n17602_), .Z(new_n17603_));
  NAND2_X1   g17502(.A1(new_n17596_), .A2(new_n17602_), .ZN(new_n17604_));
  NAND2_X1   g17503(.A1(new_n17603_), .A2(new_n17604_), .ZN(new_n17605_));
  XOR2_X1    g17504(.A1(new_n17596_), .A2(new_n17601_), .Z(new_n17606_));
  NOR2_X1    g17505(.A1(new_n17606_), .A2(new_n17594_), .ZN(new_n17607_));
  AOI21_X1   g17506(.A1(new_n17594_), .A2(new_n17605_), .B(new_n17607_), .ZN(new_n17608_));
  NAND2_X1   g17507(.A1(new_n17500_), .A2(new_n17487_), .ZN(new_n17609_));
  NAND2_X1   g17508(.A1(new_n17609_), .A2(new_n17490_), .ZN(new_n17610_));
  INV_X1     g17509(.I(new_n17610_), .ZN(new_n17611_));
  NOR2_X1    g17510(.A1(new_n17608_), .A2(new_n17611_), .ZN(new_n17612_));
  OAI21_X1   g17511(.A1(new_n17411_), .A2(new_n17520_), .B(new_n17612_), .ZN(new_n17613_));
  NOR3_X1    g17512(.A1(new_n17499_), .A2(new_n17396_), .A3(new_n17503_), .ZN(new_n17614_));
  OAI21_X1   g17513(.A1(new_n17499_), .A2(new_n17503_), .B(new_n17396_), .ZN(new_n17615_));
  AOI21_X1   g17514(.A1(new_n17318_), .A2(new_n17615_), .B(new_n17614_), .ZN(new_n17616_));
  INV_X1     g17515(.I(new_n17612_), .ZN(new_n17617_));
  NAND3_X1   g17516(.A1(new_n17316_), .A2(new_n17616_), .A3(new_n17617_), .ZN(new_n17618_));
  AOI21_X1   g17517(.A1(new_n17618_), .A2(new_n17613_), .B(new_n17499_), .ZN(new_n17619_));
  AOI21_X1   g17518(.A1(new_n17316_), .A2(new_n17616_), .B(new_n17617_), .ZN(new_n17620_));
  NOR3_X1    g17519(.A1(new_n17411_), .A2(new_n17520_), .A3(new_n17612_), .ZN(new_n17621_));
  NOR3_X1    g17520(.A1(new_n17620_), .A2(new_n17621_), .A3(new_n17516_), .ZN(new_n17622_));
  OR2_X2     g17521(.A1(new_n17619_), .A2(new_n17622_), .Z(new_n17623_));
  OAI21_X1   g17522(.A1(new_n17514_), .A2(new_n17515_), .B(new_n17623_), .ZN(new_n17624_));
  NOR2_X1    g17523(.A1(new_n17619_), .A2(new_n17622_), .ZN(new_n17625_));
  NAND4_X1   g17524(.A1(\result[15] ), .A2(new_n17513_), .A3(new_n17509_), .A4(new_n17625_), .ZN(new_n17626_));
  NAND2_X1   g17525(.A1(new_n17624_), .A2(new_n17626_), .ZN(\result[18] ));
  NOR2_X1    g17526(.A1(new_n17514_), .A2(new_n17515_), .ZN(new_n17628_));
  NAND2_X1   g17527(.A1(new_n17316_), .A2(new_n17616_), .ZN(new_n17629_));
  AOI21_X1   g17528(.A1(new_n17608_), .A2(new_n17516_), .B(new_n17611_), .ZN(new_n17630_));
  INV_X1     g17529(.I(new_n17630_), .ZN(new_n17631_));
  OAI22_X1   g17530(.A1(new_n17629_), .A2(new_n17631_), .B1(new_n17516_), .B2(new_n17608_), .ZN(new_n17632_));
  INV_X1     g17531(.I(new_n17604_), .ZN(new_n17633_));
  AND2_X2    g17532(.A1(new_n17603_), .A2(new_n17594_), .Z(new_n17634_));
  INV_X1     g17533(.I(new_n17591_), .ZN(new_n17635_));
  OAI21_X1   g17534(.A1(new_n17522_), .A2(new_n17589_), .B(new_n17635_), .ZN(new_n17636_));
  NOR2_X1    g17535(.A1(new_n17552_), .A2(new_n17561_), .ZN(new_n17637_));
  NOR2_X1    g17536(.A1(new_n17637_), .A2(new_n17562_), .ZN(new_n17638_));
  OAI22_X1   g17537(.A1(new_n10965_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n10570_), .ZN(new_n17639_));
  AOI21_X1   g17538(.A1(new_n17639_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n17640_));
  XNOR2_X1   g17539(.A1(new_n14077_), .A2(new_n17640_), .ZN(new_n17641_));
  NAND2_X1   g17540(.A1(new_n17638_), .A2(new_n17641_), .ZN(new_n17642_));
  OR2_X2     g17541(.A1(new_n17638_), .A2(new_n17641_), .Z(new_n17643_));
  NAND2_X1   g17542(.A1(new_n17643_), .A2(new_n17642_), .ZN(new_n17644_));
  INV_X1     g17543(.I(new_n17525_), .ZN(new_n17645_));
  INV_X1     g17544(.I(new_n17532_), .ZN(new_n17646_));
  AOI21_X1   g17545(.A1(new_n17645_), .A2(new_n17646_), .B(new_n17534_), .ZN(new_n17647_));
  INV_X1     g17546(.I(new_n17647_), .ZN(new_n17648_));
  OAI21_X1   g17547(.A1(new_n15515_), .A2(new_n4944_), .B(new_n279_), .ZN(new_n17649_));
  OAI21_X1   g17548(.A1(new_n4946_), .A2(new_n15515_), .B(new_n17649_), .ZN(new_n17650_));
  INV_X1     g17549(.I(new_n17650_), .ZN(new_n17651_));
  NAND2_X1   g17550(.A1(new_n12614_), .A2(new_n962_), .ZN(new_n17652_));
  AOI22_X1   g17551(.A1(new_n12204_), .A2(new_n4406_), .B1(new_n87_), .B2(new_n10600_), .ZN(new_n17653_));
  AOI21_X1   g17552(.A1(new_n17653_), .A2(new_n17652_), .B(new_n82_), .ZN(new_n17654_));
  NAND2_X1   g17553(.A1(new_n13949_), .A2(new_n17654_), .ZN(new_n17655_));
  XOR2_X1    g17554(.A1(new_n17655_), .A2(new_n17533_), .Z(new_n17656_));
  NOR2_X1    g17555(.A1(new_n17656_), .A2(new_n17651_), .ZN(new_n17657_));
  AOI21_X1   g17556(.A1(new_n13949_), .A2(new_n17654_), .B(new_n17533_), .ZN(new_n17658_));
  NOR2_X1    g17557(.A1(new_n17655_), .A2(new_n17530_), .ZN(new_n17659_));
  NOR2_X1    g17558(.A1(new_n17658_), .A2(new_n17659_), .ZN(new_n17660_));
  NOR2_X1    g17559(.A1(new_n17660_), .A2(new_n17650_), .ZN(new_n17661_));
  NOR2_X1    g17560(.A1(new_n17657_), .A2(new_n17661_), .ZN(new_n17662_));
  AOI22_X1   g17561(.A1(new_n10914_), .A2(new_n4526_), .B1(new_n4570_), .B2(new_n12616_), .ZN(new_n17663_));
  AOI21_X1   g17562(.A1(new_n101_), .A2(new_n10924_), .B(new_n17663_), .ZN(new_n17664_));
  OAI21_X1   g17563(.A1(new_n17664_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n17665_));
  XNOR2_X1   g17564(.A1(new_n12889_), .A2(new_n17665_), .ZN(new_n17666_));
  XOR2_X1    g17565(.A1(new_n17666_), .A2(new_n17662_), .Z(new_n17667_));
  NAND2_X1   g17566(.A1(new_n17648_), .A2(new_n17667_), .ZN(new_n17668_));
  AND2_X2    g17567(.A1(new_n17666_), .A2(new_n17662_), .Z(new_n17669_));
  NOR2_X1    g17568(.A1(new_n17666_), .A2(new_n17662_), .ZN(new_n17670_));
  OAI21_X1   g17569(.A1(new_n17669_), .A2(new_n17670_), .B(new_n17647_), .ZN(new_n17671_));
  NAND2_X1   g17570(.A1(new_n17668_), .A2(new_n17671_), .ZN(new_n17672_));
  NOR2_X1    g17571(.A1(new_n17548_), .A2(new_n17536_), .ZN(new_n17673_));
  NOR2_X1    g17572(.A1(new_n17673_), .A2(new_n17549_), .ZN(new_n17674_));
  OAI22_X1   g17573(.A1(new_n10583_), .A2(new_n4612_), .B1(new_n4781_), .B2(new_n10938_), .ZN(new_n17675_));
  OAI21_X1   g17574(.A1(new_n1128_), .A2(new_n10952_), .B(new_n17675_), .ZN(new_n17676_));
  AOI21_X1   g17575(.A1(new_n17676_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n17677_));
  XNOR2_X1   g17576(.A1(new_n12907_), .A2(new_n17677_), .ZN(new_n17678_));
  AND2_X2    g17577(.A1(new_n17674_), .A2(new_n17678_), .Z(new_n17679_));
  NOR2_X1    g17578(.A1(new_n17674_), .A2(new_n17678_), .ZN(new_n17680_));
  OAI21_X1   g17579(.A1(new_n17679_), .A2(new_n17680_), .B(new_n17672_), .ZN(new_n17681_));
  XOR2_X1    g17580(.A1(new_n17674_), .A2(new_n17678_), .Z(new_n17682_));
  NAND3_X1   g17581(.A1(new_n17682_), .A2(new_n17668_), .A3(new_n17671_), .ZN(new_n17683_));
  NAND2_X1   g17582(.A1(new_n17683_), .A2(new_n17681_), .ZN(new_n17684_));
  AOI22_X1   g17583(.A1(new_n14602_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n14603_), .ZN(new_n17685_));
  OAI21_X1   g17584(.A1(new_n17685_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n17686_));
  XNOR2_X1   g17585(.A1(new_n14601_), .A2(new_n17686_), .ZN(new_n17687_));
  XOR2_X1    g17586(.A1(new_n17684_), .A2(new_n17687_), .Z(new_n17688_));
  XNOR2_X1   g17587(.A1(new_n17684_), .A2(new_n17687_), .ZN(new_n17689_));
  MUX2_X1    g17588(.I0(new_n17689_), .I1(new_n17688_), .S(new_n17644_), .Z(new_n17690_));
  NOR2_X1    g17589(.A1(new_n17690_), .A2(new_n17583_), .ZN(new_n17691_));
  XNOR2_X1   g17590(.A1(new_n17691_), .A2(new_n17580_), .ZN(new_n17692_));
  NAND2_X1   g17591(.A1(new_n17692_), .A2(new_n17567_), .ZN(new_n17693_));
  OR2_X2     g17592(.A1(new_n17692_), .A2(new_n17567_), .Z(new_n17694_));
  NAND2_X1   g17593(.A1(new_n17694_), .A2(new_n17693_), .ZN(new_n17695_));
  OAI22_X1   g17594(.A1(new_n15313_), .A2(new_n5420_), .B1(new_n1620_), .B2(new_n15305_), .ZN(new_n17696_));
  AOI21_X1   g17595(.A1(new_n17696_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n17697_));
  XNOR2_X1   g17596(.A1(new_n15312_), .A2(new_n17697_), .ZN(new_n17698_));
  XOR2_X1    g17597(.A1(new_n17695_), .A2(new_n17698_), .Z(new_n17699_));
  NAND2_X1   g17598(.A1(new_n17699_), .A2(new_n17636_), .ZN(new_n17700_));
  INV_X1     g17599(.I(new_n17698_), .ZN(new_n17701_));
  XOR2_X1    g17600(.A1(new_n17695_), .A2(new_n17701_), .Z(new_n17702_));
  INV_X1     g17601(.I(new_n17702_), .ZN(new_n17703_));
  OAI21_X1   g17602(.A1(new_n17636_), .A2(new_n17703_), .B(new_n17700_), .ZN(new_n17704_));
  NOR3_X1    g17603(.A1(new_n17634_), .A2(new_n17633_), .A3(new_n17704_), .ZN(new_n17705_));
  NOR2_X1    g17604(.A1(new_n17634_), .A2(new_n17633_), .ZN(new_n17706_));
  INV_X1     g17605(.I(new_n17704_), .ZN(new_n17707_));
  NOR2_X1    g17606(.A1(new_n17706_), .A2(new_n17707_), .ZN(new_n17708_));
  OAI21_X1   g17607(.A1(new_n17705_), .A2(new_n17708_), .B(new_n17632_), .ZN(new_n17709_));
  XOR2_X1    g17608(.A1(new_n17628_), .A2(new_n17709_), .Z(new_n17710_));
  XOR2_X1    g17609(.A1(new_n17710_), .A2(new_n17625_), .Z(\result[19] ));
  AOI21_X1   g17610(.A1(new_n17624_), .A2(new_n17626_), .B(new_n17709_), .ZN(new_n17712_));
  NOR2_X1    g17611(.A1(new_n17411_), .A2(new_n17520_), .ZN(new_n17713_));
  INV_X1     g17612(.I(new_n17608_), .ZN(new_n17714_));
  AOI22_X1   g17613(.A1(new_n17713_), .A2(new_n17630_), .B1(new_n17499_), .B2(new_n17714_), .ZN(new_n17715_));
  NAND2_X1   g17614(.A1(new_n17695_), .A2(new_n17701_), .ZN(new_n17716_));
  INV_X1     g17615(.I(new_n17687_), .ZN(new_n17717_));
  XOR2_X1    g17616(.A1(new_n17644_), .A2(new_n17684_), .Z(new_n17718_));
  NOR2_X1    g17617(.A1(new_n17718_), .A2(new_n17717_), .ZN(new_n17719_));
  NOR2_X1    g17618(.A1(new_n17690_), .A2(new_n17576_), .ZN(new_n17720_));
  NOR2_X1    g17619(.A1(new_n17720_), .A2(new_n17573_), .ZN(new_n17721_));
  NAND2_X1   g17620(.A1(new_n17690_), .A2(new_n17576_), .ZN(new_n17722_));
  NAND2_X1   g17621(.A1(new_n17722_), .A2(new_n17582_), .ZN(new_n17723_));
  NOR2_X1    g17622(.A1(new_n17721_), .A2(new_n17723_), .ZN(new_n17724_));
  NOR2_X1    g17623(.A1(new_n17647_), .A2(new_n17669_), .ZN(new_n17725_));
  NOR2_X1    g17624(.A1(new_n17725_), .A2(new_n17670_), .ZN(new_n17726_));
  NOR2_X1    g17625(.A1(new_n10589_), .A2(new_n511_), .ZN(new_n17727_));
  INV_X1     g17626(.I(new_n17727_), .ZN(new_n17728_));
  AOI22_X1   g17627(.A1(new_n12614_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n10600_), .ZN(new_n17729_));
  AOI21_X1   g17628(.A1(new_n17728_), .A2(new_n17729_), .B(new_n82_), .ZN(new_n17730_));
  NAND2_X1   g17629(.A1(new_n13972_), .A2(new_n17730_), .ZN(new_n17731_));
  INV_X1     g17630(.I(new_n17731_), .ZN(new_n17732_));
  INV_X1     g17631(.I(new_n17658_), .ZN(new_n17733_));
  AOI21_X1   g17632(.A1(new_n17733_), .A2(new_n17651_), .B(new_n17659_), .ZN(new_n17734_));
  INV_X1     g17633(.I(new_n17734_), .ZN(new_n17735_));
  OAI22_X1   g17634(.A1(new_n10923_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10913_), .ZN(new_n17736_));
  OAI21_X1   g17635(.A1(new_n10583_), .A2(new_n79_), .B(new_n17736_), .ZN(new_n17737_));
  AOI21_X1   g17636(.A1(new_n17737_), .A2(new_n72_), .B(new_n79_), .ZN(new_n17738_));
  XNOR2_X1   g17637(.A1(new_n13378_), .A2(new_n17738_), .ZN(new_n17739_));
  XOR2_X1    g17638(.A1(new_n17739_), .A2(new_n17735_), .Z(new_n17740_));
  NOR2_X1    g17639(.A1(new_n17740_), .A2(new_n17732_), .ZN(new_n17741_));
  AND2_X2    g17640(.A1(new_n17739_), .A2(new_n17734_), .Z(new_n17742_));
  NOR2_X1    g17641(.A1(new_n17739_), .A2(new_n17734_), .ZN(new_n17743_));
  NOR2_X1    g17642(.A1(new_n17742_), .A2(new_n17743_), .ZN(new_n17744_));
  NOR2_X1    g17643(.A1(new_n17744_), .A2(new_n17731_), .ZN(new_n17745_));
  NOR2_X1    g17644(.A1(new_n17745_), .A2(new_n17741_), .ZN(new_n17746_));
  OAI22_X1   g17645(.A1(new_n10577_), .A2(new_n1128_), .B1(new_n4782_), .B2(new_n10953_), .ZN(new_n17747_));
  AOI21_X1   g17646(.A1(new_n17747_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n17748_));
  XOR2_X1    g17647(.A1(new_n13544_), .A2(new_n17748_), .Z(new_n17749_));
  INV_X1     g17648(.I(new_n17749_), .ZN(new_n17750_));
  NOR2_X1    g17649(.A1(new_n17750_), .A2(new_n17746_), .ZN(new_n17751_));
  INV_X1     g17650(.I(new_n17751_), .ZN(new_n17752_));
  NAND2_X1   g17651(.A1(new_n17750_), .A2(new_n17746_), .ZN(new_n17753_));
  AOI21_X1   g17652(.A1(new_n17752_), .A2(new_n17753_), .B(new_n17726_), .ZN(new_n17754_));
  XOR2_X1    g17653(.A1(new_n17746_), .A2(new_n17749_), .Z(new_n17755_));
  NOR3_X1    g17654(.A1(new_n17755_), .A2(new_n17670_), .A3(new_n17725_), .ZN(new_n17756_));
  NOR2_X1    g17655(.A1(new_n17756_), .A2(new_n17754_), .ZN(new_n17757_));
  NOR2_X1    g17656(.A1(new_n17679_), .A2(new_n17672_), .ZN(new_n17758_));
  NOR2_X1    g17657(.A1(new_n17758_), .A2(new_n17680_), .ZN(new_n17759_));
  OAI22_X1   g17658(.A1(new_n10570_), .A2(new_n4902_), .B1(new_n1973_), .B2(new_n10961_), .ZN(new_n17760_));
  OAI21_X1   g17659(.A1(new_n10564_), .A2(new_n1239_), .B(new_n17760_), .ZN(new_n17761_));
  AOI21_X1   g17660(.A1(new_n17761_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n17762_));
  XOR2_X1    g17661(.A1(new_n10976_), .A2(new_n17762_), .Z(new_n17763_));
  NAND2_X1   g17662(.A1(new_n17759_), .A2(new_n17763_), .ZN(new_n17764_));
  NOR2_X1    g17663(.A1(new_n17759_), .A2(new_n17763_), .ZN(new_n17765_));
  INV_X1     g17664(.I(new_n17765_), .ZN(new_n17766_));
  AOI21_X1   g17665(.A1(new_n17766_), .A2(new_n17764_), .B(new_n17757_), .ZN(new_n17767_));
  INV_X1     g17666(.I(new_n17757_), .ZN(new_n17768_));
  XNOR2_X1   g17667(.A1(new_n17759_), .A2(new_n17763_), .ZN(new_n17769_));
  NOR2_X1    g17668(.A1(new_n17769_), .A2(new_n17768_), .ZN(new_n17770_));
  INV_X1     g17669(.I(new_n17642_), .ZN(new_n17771_));
  OAI21_X1   g17670(.A1(new_n17771_), .A2(new_n17684_), .B(new_n17643_), .ZN(new_n17772_));
  OAI22_X1   g17671(.A1(new_n14276_), .A2(new_n4719_), .B1(new_n5335_), .B2(new_n14594_), .ZN(new_n17773_));
  OAI21_X1   g17672(.A1(new_n14886_), .A2(new_n5398_), .B(new_n17773_), .ZN(new_n17774_));
  AOI21_X1   g17673(.A1(new_n17774_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n17775_));
  XOR2_X1    g17674(.A1(new_n14891_), .A2(new_n17775_), .Z(new_n17776_));
  INV_X1     g17675(.I(new_n17776_), .ZN(new_n17777_));
  NOR2_X1    g17676(.A1(new_n17772_), .A2(new_n17777_), .ZN(new_n17778_));
  NAND2_X1   g17677(.A1(new_n17772_), .A2(new_n17777_), .ZN(new_n17779_));
  INV_X1     g17678(.I(new_n17779_), .ZN(new_n17780_));
  OAI22_X1   g17679(.A1(new_n17780_), .A2(new_n17778_), .B1(new_n17767_), .B2(new_n17770_), .ZN(new_n17781_));
  NOR2_X1    g17680(.A1(new_n17770_), .A2(new_n17767_), .ZN(new_n17782_));
  XOR2_X1    g17681(.A1(new_n17772_), .A2(new_n17777_), .Z(new_n17783_));
  NAND2_X1   g17682(.A1(new_n17783_), .A2(new_n17782_), .ZN(new_n17784_));
  NAND2_X1   g17683(.A1(new_n17784_), .A2(new_n17781_), .ZN(new_n17785_));
  INV_X1     g17684(.I(new_n17785_), .ZN(new_n17786_));
  OAI22_X1   g17685(.A1(new_n15305_), .A2(new_n5419_), .B1(new_n15114_), .B2(new_n1622_), .ZN(new_n17787_));
  OAI21_X1   g17686(.A1(new_n1620_), .A2(new_n15515_), .B(new_n17787_), .ZN(new_n17788_));
  AOI21_X1   g17687(.A1(new_n17788_), .A2(new_n126_), .B(new_n1620_), .ZN(new_n17789_));
  XOR2_X1    g17688(.A1(new_n15518_), .A2(new_n17789_), .Z(new_n17790_));
  NOR2_X1    g17689(.A1(new_n17786_), .A2(new_n17790_), .ZN(new_n17791_));
  XOR2_X1    g17690(.A1(new_n17791_), .A2(new_n17724_), .Z(new_n17792_));
  XOR2_X1    g17691(.A1(new_n17792_), .A2(new_n17719_), .Z(new_n17793_));
  NAND2_X1   g17692(.A1(new_n17702_), .A2(new_n17793_), .ZN(new_n17794_));
  XNOR2_X1   g17693(.A1(new_n17794_), .A2(new_n17716_), .ZN(new_n17795_));
  XOR2_X1    g17694(.A1(new_n17795_), .A2(new_n17636_), .Z(new_n17796_));
  XOR2_X1    g17695(.A1(new_n17706_), .A2(new_n17704_), .Z(new_n17797_));
  NOR2_X1    g17696(.A1(new_n17797_), .A2(new_n17796_), .ZN(new_n17798_));
  XOR2_X1    g17697(.A1(new_n17798_), .A2(new_n17708_), .Z(new_n17799_));
  XOR2_X1    g17698(.A1(new_n17799_), .A2(new_n17715_), .Z(new_n17800_));
  INV_X1     g17699(.I(new_n17800_), .ZN(new_n17801_));
  XOR2_X1    g17700(.A1(new_n17712_), .A2(new_n17801_), .Z(\result[20] ));
  INV_X1     g17701(.I(new_n17709_), .ZN(new_n17803_));
  AOI21_X1   g17702(.A1(new_n17793_), .A2(new_n17695_), .B(new_n17701_), .ZN(new_n17804_));
  OAI21_X1   g17703(.A1(new_n17793_), .A2(new_n17695_), .B(new_n17636_), .ZN(new_n17805_));
  NOR2_X1    g17704(.A1(new_n17804_), .A2(new_n17805_), .ZN(new_n17806_));
  INV_X1     g17705(.I(new_n17796_), .ZN(new_n17807_));
  NOR2_X1    g17706(.A1(new_n17807_), .A2(new_n17704_), .ZN(new_n17808_));
  NAND2_X1   g17707(.A1(new_n17807_), .A2(new_n17704_), .ZN(new_n17809_));
  AOI21_X1   g17708(.A1(new_n17706_), .A2(new_n17809_), .B(new_n17808_), .ZN(new_n17810_));
  INV_X1     g17709(.I(new_n17810_), .ZN(new_n17811_));
  NOR2_X1    g17710(.A1(new_n17785_), .A2(new_n17719_), .ZN(new_n17812_));
  NOR2_X1    g17711(.A1(new_n17812_), .A2(new_n17790_), .ZN(new_n17813_));
  AOI22_X1   g17712(.A1(new_n17813_), .A2(new_n17724_), .B1(new_n17719_), .B2(new_n17785_), .ZN(new_n17814_));
  OAI21_X1   g17713(.A1(new_n17726_), .A2(new_n17751_), .B(new_n17753_), .ZN(new_n17815_));
  INV_X1     g17714(.I(new_n17815_), .ZN(new_n17816_));
  OAI22_X1   g17715(.A1(new_n10583_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10923_), .ZN(new_n17817_));
  OAI21_X1   g17716(.A1(new_n79_), .A2(new_n10938_), .B(new_n17817_), .ZN(new_n17818_));
  AOI21_X1   g17717(.A1(new_n17818_), .A2(new_n72_), .B(new_n79_), .ZN(new_n17819_));
  XOR2_X1    g17718(.A1(new_n13394_), .A2(new_n17819_), .Z(new_n17820_));
  NOR2_X1    g17719(.A1(new_n10913_), .A2(new_n511_), .ZN(new_n17821_));
  INV_X1     g17720(.I(new_n17821_), .ZN(new_n17822_));
  AOI22_X1   g17721(.A1(new_n12616_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n12614_), .ZN(new_n17823_));
  AOI21_X1   g17722(.A1(new_n17822_), .A2(new_n17823_), .B(new_n82_), .ZN(new_n17824_));
  OAI21_X1   g17723(.A1(new_n12766_), .A2(new_n12764_), .B(new_n17824_), .ZN(new_n17825_));
  INV_X1     g17724(.I(new_n17825_), .ZN(new_n17826_));
  XOR2_X1    g17725(.A1(new_n17820_), .A2(new_n17826_), .Z(new_n17827_));
  NOR2_X1    g17726(.A1(new_n17827_), .A2(new_n17732_), .ZN(new_n17828_));
  INV_X1     g17727(.I(new_n17820_), .ZN(new_n17829_));
  NOR2_X1    g17728(.A1(new_n17829_), .A2(new_n17826_), .ZN(new_n17830_));
  NOR2_X1    g17729(.A1(new_n17820_), .A2(new_n17825_), .ZN(new_n17831_));
  NOR2_X1    g17730(.A1(new_n17830_), .A2(new_n17831_), .ZN(new_n17832_));
  NOR2_X1    g17731(.A1(new_n17832_), .A2(new_n17731_), .ZN(new_n17833_));
  NOR2_X1    g17732(.A1(new_n17833_), .A2(new_n17828_), .ZN(new_n17834_));
  INV_X1     g17733(.I(new_n17742_), .ZN(new_n17835_));
  AOI21_X1   g17734(.A1(new_n17835_), .A2(new_n17731_), .B(new_n17743_), .ZN(new_n17836_));
  INV_X1     g17735(.I(new_n17836_), .ZN(new_n17837_));
  OAI22_X1   g17736(.A1(new_n10577_), .A2(new_n4781_), .B1(new_n4612_), .B2(new_n10952_), .ZN(new_n17838_));
  OAI21_X1   g17737(.A1(new_n1128_), .A2(new_n10961_), .B(new_n17838_), .ZN(new_n17839_));
  AOI21_X1   g17738(.A1(new_n17839_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n17840_));
  XOR2_X1    g17739(.A1(new_n14053_), .A2(new_n17840_), .Z(new_n17841_));
  XOR2_X1    g17740(.A1(new_n17841_), .A2(new_n17837_), .Z(new_n17842_));
  NOR2_X1    g17741(.A1(new_n17842_), .A2(new_n17834_), .ZN(new_n17843_));
  AND2_X2    g17742(.A1(new_n17841_), .A2(new_n17836_), .Z(new_n17844_));
  NOR2_X1    g17743(.A1(new_n17841_), .A2(new_n17836_), .ZN(new_n17845_));
  NOR2_X1    g17744(.A1(new_n17844_), .A2(new_n17845_), .ZN(new_n17846_));
  NOR3_X1    g17745(.A1(new_n17846_), .A2(new_n17828_), .A3(new_n17833_), .ZN(new_n17847_));
  NOR2_X1    g17746(.A1(new_n17847_), .A2(new_n17843_), .ZN(new_n17848_));
  AOI22_X1   g17747(.A1(new_n14281_), .A2(new_n5783_), .B1(new_n247_), .B2(new_n14274_), .ZN(new_n17849_));
  OAI21_X1   g17748(.A1(new_n17849_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n17850_));
  XOR2_X1    g17749(.A1(new_n14280_), .A2(new_n17850_), .Z(new_n17851_));
  NAND2_X1   g17750(.A1(new_n17848_), .A2(new_n17851_), .ZN(new_n17852_));
  INV_X1     g17751(.I(new_n17848_), .ZN(new_n17853_));
  INV_X1     g17752(.I(new_n17851_), .ZN(new_n17854_));
  NAND2_X1   g17753(.A1(new_n17853_), .A2(new_n17854_), .ZN(new_n17855_));
  AOI21_X1   g17754(.A1(new_n17855_), .A2(new_n17852_), .B(new_n17816_), .ZN(new_n17856_));
  XOR2_X1    g17755(.A1(new_n17848_), .A2(new_n17851_), .Z(new_n17857_));
  AOI21_X1   g17756(.A1(new_n17857_), .A2(new_n17816_), .B(new_n17856_), .ZN(new_n17858_));
  NAND2_X1   g17757(.A1(new_n17764_), .A2(new_n17768_), .ZN(new_n17859_));
  NAND2_X1   g17758(.A1(new_n17859_), .A2(new_n17766_), .ZN(new_n17860_));
  INV_X1     g17759(.I(new_n17860_), .ZN(new_n17861_));
  AOI22_X1   g17760(.A1(new_n15127_), .A2(new_n5337_), .B1(new_n4717_), .B2(new_n15115_), .ZN(new_n17862_));
  OAI21_X1   g17761(.A1(new_n17862_), .A2(\a[20] ), .B(new_n4717_), .ZN(new_n17863_));
  XNOR2_X1   g17762(.A1(new_n15125_), .A2(new_n17863_), .ZN(new_n17864_));
  AND2_X2    g17763(.A1(new_n17864_), .A2(new_n17861_), .Z(new_n17865_));
  NOR2_X1    g17764(.A1(new_n17864_), .A2(new_n17861_), .ZN(new_n17866_));
  NOR2_X1    g17765(.A1(new_n17865_), .A2(new_n17866_), .ZN(new_n17867_));
  NOR2_X1    g17766(.A1(new_n17867_), .A2(new_n17858_), .ZN(new_n17868_));
  XOR2_X1    g17767(.A1(new_n17864_), .A2(new_n17860_), .Z(new_n17869_));
  INV_X1     g17768(.I(new_n17869_), .ZN(new_n17870_));
  AOI21_X1   g17769(.A1(new_n17858_), .A2(new_n17870_), .B(new_n17868_), .ZN(new_n17871_));
  OAI21_X1   g17770(.A1(new_n17782_), .A2(new_n17778_), .B(new_n17779_), .ZN(new_n17872_));
  NAND2_X1   g17771(.A1(new_n15515_), .A2(new_n4663_), .ZN(new_n17873_));
  NOR2_X1    g17772(.A1(new_n4661_), .A2(new_n4660_), .ZN(new_n17874_));
  AOI21_X1   g17773(.A1(new_n15675_), .A2(new_n17874_), .B(\a[17] ), .ZN(new_n17875_));
  AOI21_X1   g17774(.A1(new_n17875_), .A2(new_n17873_), .B(new_n1620_), .ZN(new_n17876_));
  XNOR2_X1   g17775(.A1(new_n15678_), .A2(new_n17876_), .ZN(new_n17877_));
  INV_X1     g17776(.I(new_n17877_), .ZN(new_n17878_));
  NOR2_X1    g17777(.A1(new_n17872_), .A2(new_n17878_), .ZN(new_n17879_));
  INV_X1     g17778(.I(new_n17879_), .ZN(new_n17880_));
  NAND2_X1   g17779(.A1(new_n17872_), .A2(new_n17878_), .ZN(new_n17881_));
  AOI21_X1   g17780(.A1(new_n17880_), .A2(new_n17881_), .B(new_n17871_), .ZN(new_n17882_));
  XOR2_X1    g17781(.A1(new_n17872_), .A2(new_n17877_), .Z(new_n17883_));
  INV_X1     g17782(.I(new_n17883_), .ZN(new_n17884_));
  AOI21_X1   g17783(.A1(new_n17871_), .A2(new_n17884_), .B(new_n17882_), .ZN(new_n17885_));
  NOR2_X1    g17784(.A1(new_n17885_), .A2(new_n17814_), .ZN(new_n17886_));
  OAI21_X1   g17785(.A1(new_n17811_), .A2(new_n17715_), .B(new_n17886_), .ZN(new_n17887_));
  INV_X1     g17786(.I(new_n17886_), .ZN(new_n17888_));
  NAND3_X1   g17787(.A1(new_n17632_), .A2(new_n17810_), .A3(new_n17888_), .ZN(new_n17889_));
  AOI21_X1   g17788(.A1(new_n17887_), .A2(new_n17889_), .B(new_n17806_), .ZN(new_n17890_));
  INV_X1     g17789(.I(new_n17806_), .ZN(new_n17891_));
  AOI21_X1   g17790(.A1(new_n17632_), .A2(new_n17810_), .B(new_n17888_), .ZN(new_n17892_));
  NOR3_X1    g17791(.A1(new_n17811_), .A2(new_n17715_), .A3(new_n17886_), .ZN(new_n17893_));
  NOR3_X1    g17792(.A1(new_n17893_), .A2(new_n17892_), .A3(new_n17891_), .ZN(new_n17894_));
  NOR2_X1    g17793(.A1(new_n17890_), .A2(new_n17894_), .ZN(new_n17895_));
  NAND4_X1   g17794(.A1(\result[18] ), .A2(new_n17803_), .A3(new_n17801_), .A4(new_n17895_), .ZN(new_n17896_));
  AOI21_X1   g17795(.A1(new_n17408_), .A2(new_n17509_), .B(new_n17625_), .ZN(new_n17897_));
  NOR3_X1    g17796(.A1(new_n17514_), .A2(new_n17623_), .A3(new_n17515_), .ZN(new_n17898_));
  OAI21_X1   g17797(.A1(new_n17898_), .A2(new_n17897_), .B(new_n17803_), .ZN(new_n17899_));
  OR2_X2     g17798(.A1(new_n17890_), .A2(new_n17894_), .Z(new_n17900_));
  OAI21_X1   g17799(.A1(new_n17899_), .A2(new_n17800_), .B(new_n17900_), .ZN(new_n17901_));
  NAND2_X1   g17800(.A1(new_n17901_), .A2(new_n17896_), .ZN(\result[21] ));
  NAND2_X1   g17801(.A1(new_n17712_), .A2(new_n17801_), .ZN(new_n17903_));
  NOR2_X1    g17802(.A1(new_n17811_), .A2(new_n17715_), .ZN(new_n17904_));
  NOR2_X1    g17803(.A1(new_n17891_), .A2(new_n17814_), .ZN(new_n17905_));
  AOI21_X1   g17804(.A1(new_n17891_), .A2(new_n17814_), .B(new_n17885_), .ZN(new_n17906_));
  AOI21_X1   g17805(.A1(new_n17904_), .A2(new_n17906_), .B(new_n17905_), .ZN(new_n17907_));
  OAI21_X1   g17806(.A1(new_n17871_), .A2(new_n17879_), .B(new_n17881_), .ZN(new_n17908_));
  NOR2_X1    g17807(.A1(new_n17865_), .A2(new_n17858_), .ZN(new_n17909_));
  NOR2_X1    g17808(.A1(new_n17909_), .A2(new_n17866_), .ZN(new_n17910_));
  INV_X1     g17809(.I(new_n17910_), .ZN(new_n17911_));
  INV_X1     g17810(.I(new_n17844_), .ZN(new_n17912_));
  AOI21_X1   g17811(.A1(new_n17912_), .A2(new_n17834_), .B(new_n17845_), .ZN(new_n17913_));
  OAI22_X1   g17812(.A1(new_n10577_), .A2(new_n4612_), .B1(new_n4781_), .B2(new_n10961_), .ZN(new_n17914_));
  OAI21_X1   g17813(.A1(new_n1128_), .A2(new_n10570_), .B(new_n17914_), .ZN(new_n17915_));
  AOI21_X1   g17814(.A1(new_n17915_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n17916_));
  XNOR2_X1   g17815(.A1(new_n14077_), .A2(new_n17916_), .ZN(new_n17917_));
  AND2_X2    g17816(.A1(new_n17913_), .A2(new_n17917_), .Z(new_n17918_));
  NOR2_X1    g17817(.A1(new_n17913_), .A2(new_n17917_), .ZN(new_n17919_));
  NOR2_X1    g17818(.A1(new_n17918_), .A2(new_n17919_), .ZN(new_n17920_));
  INV_X1     g17819(.I(new_n17831_), .ZN(new_n17921_));
  OAI21_X1   g17820(.A1(new_n17732_), .A2(new_n17830_), .B(new_n17921_), .ZN(new_n17922_));
  OAI21_X1   g17821(.A1(new_n15515_), .A2(new_n4664_), .B(new_n126_), .ZN(new_n17923_));
  OAI21_X1   g17822(.A1(new_n4666_), .A2(new_n15515_), .B(new_n17923_), .ZN(new_n17924_));
  INV_X1     g17823(.I(new_n17924_), .ZN(new_n17925_));
  NOR2_X1    g17824(.A1(new_n10913_), .A2(new_n88_), .ZN(new_n17926_));
  INV_X1     g17825(.I(new_n17926_), .ZN(new_n17927_));
  AOI22_X1   g17826(.A1(new_n10924_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n12616_), .ZN(new_n17928_));
  AOI21_X1   g17827(.A1(new_n17928_), .A2(new_n17927_), .B(new_n82_), .ZN(new_n17929_));
  AOI21_X1   g17828(.A1(new_n14531_), .A2(new_n17929_), .B(new_n17925_), .ZN(new_n17930_));
  NAND2_X1   g17829(.A1(new_n14531_), .A2(new_n17929_), .ZN(new_n17931_));
  NOR2_X1    g17830(.A1(new_n17931_), .A2(new_n17924_), .ZN(new_n17932_));
  NOR2_X1    g17831(.A1(new_n17932_), .A2(new_n17930_), .ZN(new_n17933_));
  NOR2_X1    g17832(.A1(new_n17933_), .A2(new_n17731_), .ZN(new_n17934_));
  XOR2_X1    g17833(.A1(new_n17931_), .A2(new_n17925_), .Z(new_n17935_));
  NOR2_X1    g17834(.A1(new_n17935_), .A2(new_n17732_), .ZN(new_n17936_));
  NOR2_X1    g17835(.A1(new_n17936_), .A2(new_n17934_), .ZN(new_n17937_));
  XOR2_X1    g17836(.A1(new_n17922_), .A2(new_n17937_), .Z(new_n17938_));
  OAI22_X1   g17837(.A1(new_n10583_), .A2(new_n4529_), .B1(new_n4527_), .B2(new_n10938_), .ZN(new_n17939_));
  OAI21_X1   g17838(.A1(new_n79_), .A2(new_n10952_), .B(new_n17939_), .ZN(new_n17940_));
  AOI21_X1   g17839(.A1(new_n17940_), .A2(new_n72_), .B(new_n79_), .ZN(new_n17941_));
  XNOR2_X1   g17840(.A1(new_n12907_), .A2(new_n17941_), .ZN(new_n17942_));
  INV_X1     g17841(.I(new_n17942_), .ZN(new_n17943_));
  NOR2_X1    g17842(.A1(new_n17938_), .A2(new_n17943_), .ZN(new_n17944_));
  NAND2_X1   g17843(.A1(new_n17938_), .A2(new_n17943_), .ZN(new_n17945_));
  INV_X1     g17844(.I(new_n17945_), .ZN(new_n17946_));
  NOR2_X1    g17845(.A1(new_n17946_), .A2(new_n17944_), .ZN(new_n17947_));
  AOI22_X1   g17846(.A1(new_n14602_), .A2(new_n5783_), .B1(new_n247_), .B2(new_n14603_), .ZN(new_n17948_));
  OAI21_X1   g17847(.A1(new_n17948_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n17949_));
  XOR2_X1    g17848(.A1(new_n14601_), .A2(new_n17949_), .Z(new_n17950_));
  XOR2_X1    g17849(.A1(new_n17947_), .A2(new_n17950_), .Z(new_n17951_));
  NOR2_X1    g17850(.A1(new_n17951_), .A2(new_n17920_), .ZN(new_n17952_));
  XOR2_X1    g17851(.A1(new_n17947_), .A2(new_n17950_), .Z(new_n17953_));
  AOI21_X1   g17852(.A1(new_n17920_), .A2(new_n17953_), .B(new_n17952_), .ZN(new_n17954_));
  INV_X1     g17853(.I(new_n17954_), .ZN(new_n17955_));
  NAND2_X1   g17854(.A1(new_n17955_), .A2(new_n17857_), .ZN(new_n17956_));
  XOR2_X1    g17855(.A1(new_n17956_), .A2(new_n17855_), .Z(new_n17957_));
  NAND2_X1   g17856(.A1(new_n17957_), .A2(new_n17816_), .ZN(new_n17958_));
  OR2_X2     g17857(.A1(new_n17957_), .A2(new_n17816_), .Z(new_n17959_));
  NAND2_X1   g17858(.A1(new_n17959_), .A2(new_n17958_), .ZN(new_n17960_));
  OAI22_X1   g17859(.A1(new_n15313_), .A2(new_n5336_), .B1(new_n5398_), .B2(new_n15305_), .ZN(new_n17961_));
  AOI21_X1   g17860(.A1(new_n17961_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n17962_));
  XNOR2_X1   g17861(.A1(new_n15312_), .A2(new_n17962_), .ZN(new_n17963_));
  INV_X1     g17862(.I(new_n17963_), .ZN(new_n17964_));
  NOR2_X1    g17863(.A1(new_n17960_), .A2(new_n17964_), .ZN(new_n17965_));
  AOI21_X1   g17864(.A1(new_n17959_), .A2(new_n17958_), .B(new_n17963_), .ZN(new_n17966_));
  OAI21_X1   g17865(.A1(new_n17965_), .A2(new_n17966_), .B(new_n17911_), .ZN(new_n17967_));
  XOR2_X1    g17866(.A1(new_n17960_), .A2(new_n17964_), .Z(new_n17968_));
  NAND2_X1   g17867(.A1(new_n17968_), .A2(new_n17910_), .ZN(new_n17969_));
  NAND2_X1   g17868(.A1(new_n17969_), .A2(new_n17967_), .ZN(new_n17970_));
  XOR2_X1    g17869(.A1(new_n17970_), .A2(new_n17908_), .Z(new_n17971_));
  NOR2_X1    g17870(.A1(new_n17907_), .A2(new_n17971_), .ZN(new_n17972_));
  XOR2_X1    g17871(.A1(new_n17895_), .A2(new_n17972_), .Z(new_n17973_));
  XOR2_X1    g17872(.A1(new_n17973_), .A2(new_n17903_), .Z(\result[22] ));
  INV_X1     g17873(.I(new_n17972_), .ZN(new_n17975_));
  AOI21_X1   g17874(.A1(new_n17901_), .A2(new_n17896_), .B(new_n17975_), .ZN(new_n17976_));
  NAND2_X1   g17875(.A1(new_n17632_), .A2(new_n17810_), .ZN(new_n17977_));
  INV_X1     g17876(.I(new_n17906_), .ZN(new_n17978_));
  OAI22_X1   g17877(.A1(new_n17977_), .A2(new_n17978_), .B1(new_n17891_), .B2(new_n17814_), .ZN(new_n17979_));
  NAND2_X1   g17878(.A1(new_n17970_), .A2(new_n17908_), .ZN(new_n17980_));
  XNOR2_X1   g17879(.A1(new_n17920_), .A2(new_n17947_), .ZN(new_n17981_));
  NOR2_X1    g17880(.A1(new_n17981_), .A2(new_n17950_), .ZN(new_n17982_));
  AOI21_X1   g17881(.A1(new_n17955_), .A2(new_n17854_), .B(new_n17853_), .ZN(new_n17983_));
  OAI21_X1   g17882(.A1(new_n17955_), .A2(new_n17854_), .B(new_n17815_), .ZN(new_n17984_));
  NOR2_X1    g17883(.A1(new_n17983_), .A2(new_n17984_), .ZN(new_n17985_));
  INV_X1     g17884(.I(new_n17937_), .ZN(new_n17986_));
  NOR2_X1    g17885(.A1(new_n17922_), .A2(new_n17986_), .ZN(new_n17987_));
  INV_X1     g17886(.I(new_n17930_), .ZN(new_n17988_));
  AOI21_X1   g17887(.A1(new_n17988_), .A2(new_n17732_), .B(new_n17932_), .ZN(new_n17989_));
  NOR2_X1    g17888(.A1(new_n10583_), .A2(new_n511_), .ZN(new_n17990_));
  INV_X1     g17889(.I(new_n17990_), .ZN(new_n17991_));
  AOI22_X1   g17890(.A1(new_n10924_), .A2(new_n87_), .B1(new_n4406_), .B2(new_n10914_), .ZN(new_n17992_));
  AOI21_X1   g17891(.A1(new_n17991_), .A2(new_n17992_), .B(new_n82_), .ZN(new_n17993_));
  NAND2_X1   g17892(.A1(new_n13378_), .A2(new_n17993_), .ZN(new_n17994_));
  OAI22_X1   g17893(.A1(new_n10577_), .A2(new_n79_), .B1(new_n4530_), .B2(new_n10953_), .ZN(new_n17995_));
  AOI21_X1   g17894(.A1(new_n17995_), .A2(new_n72_), .B(new_n79_), .ZN(new_n17996_));
  XOR2_X1    g17895(.A1(new_n13544_), .A2(new_n17996_), .Z(new_n17997_));
  XOR2_X1    g17896(.A1(new_n17997_), .A2(new_n17994_), .Z(new_n17998_));
  NOR2_X1    g17897(.A1(new_n17998_), .A2(new_n17989_), .ZN(new_n17999_));
  INV_X1     g17898(.I(new_n17989_), .ZN(new_n18000_));
  INV_X1     g17899(.I(new_n17994_), .ZN(new_n18001_));
  AND2_X2    g17900(.A1(new_n17997_), .A2(new_n18001_), .Z(new_n18002_));
  NOR2_X1    g17901(.A1(new_n17997_), .A2(new_n18001_), .ZN(new_n18003_));
  NOR2_X1    g17902(.A1(new_n18002_), .A2(new_n18003_), .ZN(new_n18004_));
  NOR2_X1    g17903(.A1(new_n18004_), .A2(new_n18000_), .ZN(new_n18005_));
  NOR2_X1    g17904(.A1(new_n18005_), .A2(new_n17999_), .ZN(new_n18006_));
  INV_X1     g17905(.I(new_n18006_), .ZN(new_n18007_));
  NOR2_X1    g17906(.A1(new_n10570_), .A2(new_n10961_), .ZN(new_n18008_));
  OAI22_X1   g17907(.A1(new_n10564_), .A2(new_n1128_), .B1(new_n4782_), .B2(new_n18008_), .ZN(new_n18009_));
  AOI21_X1   g17908(.A1(new_n18009_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n18010_));
  XNOR2_X1   g17909(.A1(new_n10976_), .A2(new_n18010_), .ZN(new_n18011_));
  NAND2_X1   g17910(.A1(new_n18007_), .A2(new_n18011_), .ZN(new_n18012_));
  XOR2_X1    g17911(.A1(new_n18012_), .A2(new_n17944_), .Z(new_n18013_));
  XOR2_X1    g17912(.A1(new_n18013_), .A2(new_n17987_), .Z(new_n18014_));
  NOR2_X1    g17913(.A1(new_n17918_), .A2(new_n17947_), .ZN(new_n18015_));
  NOR2_X1    g17914(.A1(new_n18015_), .A2(new_n17919_), .ZN(new_n18016_));
  INV_X1     g17915(.I(new_n18016_), .ZN(new_n18017_));
  OAI22_X1   g17916(.A1(new_n14276_), .A2(new_n1973_), .B1(new_n4902_), .B2(new_n14594_), .ZN(new_n18018_));
  OAI21_X1   g17917(.A1(new_n14886_), .A2(new_n1239_), .B(new_n18018_), .ZN(new_n18019_));
  AOI21_X1   g17918(.A1(new_n18019_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n18020_));
  XOR2_X1    g17919(.A1(new_n14891_), .A2(new_n18020_), .Z(new_n18021_));
  INV_X1     g17920(.I(new_n18021_), .ZN(new_n18022_));
  NOR2_X1    g17921(.A1(new_n18017_), .A2(new_n18022_), .ZN(new_n18023_));
  NOR2_X1    g17922(.A1(new_n18016_), .A2(new_n18021_), .ZN(new_n18024_));
  NOR2_X1    g17923(.A1(new_n18023_), .A2(new_n18024_), .ZN(new_n18025_));
  NOR2_X1    g17924(.A1(new_n18025_), .A2(new_n18014_), .ZN(new_n18026_));
  XOR2_X1    g17925(.A1(new_n18016_), .A2(new_n18021_), .Z(new_n18027_));
  AOI21_X1   g17926(.A1(new_n18014_), .A2(new_n18027_), .B(new_n18026_), .ZN(new_n18028_));
  OAI22_X1   g17927(.A1(new_n15305_), .A2(new_n5335_), .B1(new_n15114_), .B2(new_n4719_), .ZN(new_n18029_));
  OAI21_X1   g17928(.A1(new_n5398_), .A2(new_n15515_), .B(new_n18029_), .ZN(new_n18030_));
  AOI21_X1   g17929(.A1(new_n18030_), .A2(new_n90_), .B(new_n5398_), .ZN(new_n18031_));
  XOR2_X1    g17930(.A1(new_n15518_), .A2(new_n18031_), .Z(new_n18032_));
  NOR2_X1    g17931(.A1(new_n18028_), .A2(new_n18032_), .ZN(new_n18033_));
  XOR2_X1    g17932(.A1(new_n18033_), .A2(new_n17985_), .Z(new_n18034_));
  XOR2_X1    g17933(.A1(new_n18034_), .A2(new_n17982_), .Z(new_n18035_));
  NAND2_X1   g17934(.A1(new_n17968_), .A2(new_n18035_), .ZN(new_n18036_));
  XOR2_X1    g17935(.A1(new_n18036_), .A2(new_n17966_), .Z(new_n18037_));
  XOR2_X1    g17936(.A1(new_n18037_), .A2(new_n17910_), .Z(new_n18038_));
  XOR2_X1    g17937(.A1(new_n17970_), .A2(new_n17908_), .Z(new_n18039_));
  NAND2_X1   g17938(.A1(new_n18038_), .A2(new_n18039_), .ZN(new_n18040_));
  XNOR2_X1   g17939(.A1(new_n18040_), .A2(new_n17980_), .ZN(new_n18041_));
  XOR2_X1    g17940(.A1(new_n17979_), .A2(new_n18041_), .Z(new_n18042_));
  INV_X1     g17941(.I(new_n18042_), .ZN(new_n18043_));
  XOR2_X1    g17942(.A1(new_n17976_), .A2(new_n18043_), .Z(\result[23] ));
  NOR3_X1    g17943(.A1(new_n17899_), .A2(new_n17900_), .A3(new_n17800_), .ZN(new_n18045_));
  AOI21_X1   g17944(.A1(new_n17712_), .A2(new_n17801_), .B(new_n17895_), .ZN(new_n18046_));
  OAI21_X1   g17945(.A1(new_n18045_), .A2(new_n18046_), .B(new_n17972_), .ZN(new_n18047_));
  AOI21_X1   g17946(.A1(new_n18035_), .A2(new_n17960_), .B(new_n17964_), .ZN(new_n18048_));
  OAI21_X1   g17947(.A1(new_n18035_), .A2(new_n17960_), .B(new_n17911_), .ZN(new_n18049_));
  NOR2_X1    g17948(.A1(new_n18048_), .A2(new_n18049_), .ZN(new_n18050_));
  INV_X1     g17949(.I(new_n17908_), .ZN(new_n18051_));
  NOR2_X1    g17950(.A1(new_n18038_), .A2(new_n17970_), .ZN(new_n18052_));
  NAND2_X1   g17951(.A1(new_n18038_), .A2(new_n17970_), .ZN(new_n18053_));
  AOI21_X1   g17952(.A1(new_n18051_), .A2(new_n18053_), .B(new_n18052_), .ZN(new_n18054_));
  INV_X1     g17953(.I(new_n18054_), .ZN(new_n18055_));
  INV_X1     g17954(.I(new_n18002_), .ZN(new_n18056_));
  AOI21_X1   g17955(.A1(new_n18056_), .A2(new_n18000_), .B(new_n18003_), .ZN(new_n18057_));
  NOR2_X1    g17956(.A1(new_n10583_), .A2(new_n88_), .ZN(new_n18058_));
  INV_X1     g17957(.I(new_n18058_), .ZN(new_n18059_));
  AOI22_X1   g17958(.A1(new_n10937_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n10924_), .ZN(new_n18060_));
  AOI21_X1   g17959(.A1(new_n18059_), .A2(new_n18060_), .B(new_n82_), .ZN(new_n18061_));
  NAND2_X1   g17960(.A1(new_n14014_), .A2(new_n18061_), .ZN(new_n18062_));
  XOR2_X1    g17961(.A1(new_n18062_), .A2(new_n17994_), .Z(new_n18063_));
  NOR2_X1    g17962(.A1(new_n18057_), .A2(new_n18063_), .ZN(new_n18064_));
  INV_X1     g17963(.I(new_n18057_), .ZN(new_n18065_));
  NOR2_X1    g17964(.A1(new_n18062_), .A2(new_n18001_), .ZN(new_n18066_));
  INV_X1     g17965(.I(new_n18062_), .ZN(new_n18067_));
  NOR2_X1    g17966(.A1(new_n18067_), .A2(new_n17994_), .ZN(new_n18068_));
  NOR2_X1    g17967(.A1(new_n18068_), .A2(new_n18066_), .ZN(new_n18069_));
  NOR2_X1    g17968(.A1(new_n18065_), .A2(new_n18069_), .ZN(new_n18070_));
  NOR2_X1    g17969(.A1(new_n18070_), .A2(new_n18064_), .ZN(new_n18071_));
  INV_X1     g17970(.I(new_n18071_), .ZN(new_n18072_));
  AOI22_X1   g17971(.A1(new_n10971_), .A2(new_n4767_), .B1(new_n4613_), .B2(new_n10571_), .ZN(new_n18073_));
  AOI21_X1   g17972(.A1(new_n117_), .A2(new_n14274_), .B(new_n18073_), .ZN(new_n18074_));
  OAI21_X1   g17973(.A1(new_n18074_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n18075_));
  XOR2_X1    g17974(.A1(new_n14280_), .A2(new_n18075_), .Z(new_n18076_));
  OAI22_X1   g17975(.A1(new_n10577_), .A2(new_n4527_), .B1(new_n4529_), .B2(new_n10952_), .ZN(new_n18077_));
  OAI21_X1   g17976(.A1(new_n79_), .A2(new_n10961_), .B(new_n18077_), .ZN(new_n18078_));
  AOI21_X1   g17977(.A1(new_n18078_), .A2(new_n72_), .B(new_n79_), .ZN(new_n18079_));
  XOR2_X1    g17978(.A1(new_n14053_), .A2(new_n18079_), .Z(new_n18080_));
  INV_X1     g17979(.I(new_n18080_), .ZN(new_n18081_));
  XOR2_X1    g17980(.A1(new_n18076_), .A2(new_n18081_), .Z(new_n18082_));
  INV_X1     g17981(.I(new_n18082_), .ZN(new_n18083_));
  AND2_X2    g17982(.A1(new_n18076_), .A2(new_n18080_), .Z(new_n18084_));
  NOR2_X1    g17983(.A1(new_n18076_), .A2(new_n18080_), .ZN(new_n18085_));
  NOR2_X1    g17984(.A1(new_n18084_), .A2(new_n18085_), .ZN(new_n18086_));
  NOR2_X1    g17985(.A1(new_n18086_), .A2(new_n18072_), .ZN(new_n18087_));
  AOI21_X1   g17986(.A1(new_n18072_), .A2(new_n18083_), .B(new_n18087_), .ZN(new_n18088_));
  OAI21_X1   g17987(.A1(new_n18007_), .A2(new_n17987_), .B(new_n17944_), .ZN(new_n18089_));
  INV_X1     g17988(.I(new_n18089_), .ZN(new_n18090_));
  AOI22_X1   g17989(.A1(new_n18090_), .A2(new_n18011_), .B1(new_n17987_), .B2(new_n18007_), .ZN(new_n18091_));
  AOI22_X1   g17990(.A1(new_n15127_), .A2(new_n5783_), .B1(new_n247_), .B2(new_n15115_), .ZN(new_n18092_));
  OAI21_X1   g17991(.A1(new_n18092_), .A2(\a[23] ), .B(new_n247_), .ZN(new_n18093_));
  XNOR2_X1   g17992(.A1(new_n15125_), .A2(new_n18093_), .ZN(new_n18094_));
  AND2_X2    g17993(.A1(new_n18094_), .A2(new_n18091_), .Z(new_n18095_));
  NOR2_X1    g17994(.A1(new_n18094_), .A2(new_n18091_), .ZN(new_n18096_));
  NOR2_X1    g17995(.A1(new_n18095_), .A2(new_n18096_), .ZN(new_n18097_));
  NOR2_X1    g17996(.A1(new_n18097_), .A2(new_n18088_), .ZN(new_n18098_));
  INV_X1     g17997(.I(new_n18088_), .ZN(new_n18099_));
  XNOR2_X1   g17998(.A1(new_n18094_), .A2(new_n18091_), .ZN(new_n18100_));
  NOR2_X1    g17999(.A1(new_n18100_), .A2(new_n18099_), .ZN(new_n18101_));
  NOR2_X1    g18000(.A1(new_n18098_), .A2(new_n18101_), .ZN(new_n18102_));
  INV_X1     g18001(.I(new_n18024_), .ZN(new_n18103_));
  OAI21_X1   g18002(.A1(new_n18014_), .A2(new_n18023_), .B(new_n18103_), .ZN(new_n18104_));
  NAND2_X1   g18003(.A1(new_n15515_), .A2(new_n4722_), .ZN(new_n18105_));
  NOR2_X1    g18004(.A1(new_n4720_), .A2(new_n4717_), .ZN(new_n18106_));
  AOI21_X1   g18005(.A1(new_n15675_), .A2(new_n18106_), .B(\a[20] ), .ZN(new_n18107_));
  AOI21_X1   g18006(.A1(new_n18107_), .A2(new_n18105_), .B(new_n5398_), .ZN(new_n18108_));
  XNOR2_X1   g18007(.A1(new_n15678_), .A2(new_n18108_), .ZN(new_n18109_));
  INV_X1     g18008(.I(new_n18109_), .ZN(new_n18110_));
  NOR2_X1    g18009(.A1(new_n18104_), .A2(new_n18110_), .ZN(new_n18111_));
  AND2_X2    g18010(.A1(new_n18104_), .A2(new_n18110_), .Z(new_n18112_));
  NOR2_X1    g18011(.A1(new_n18112_), .A2(new_n18111_), .ZN(new_n18113_));
  NOR2_X1    g18012(.A1(new_n18113_), .A2(new_n18102_), .ZN(new_n18114_));
  XOR2_X1    g18013(.A1(new_n18104_), .A2(new_n18109_), .Z(new_n18115_));
  INV_X1     g18014(.I(new_n18115_), .ZN(new_n18116_));
  AOI21_X1   g18015(.A1(new_n18102_), .A2(new_n18116_), .B(new_n18114_), .ZN(new_n18117_));
  INV_X1     g18016(.I(new_n18028_), .ZN(new_n18118_));
  NOR2_X1    g18017(.A1(new_n18118_), .A2(new_n17985_), .ZN(new_n18119_));
  NOR4_X1    g18018(.A1(new_n18119_), .A2(new_n17950_), .A3(new_n17981_), .A4(new_n18032_), .ZN(new_n18120_));
  AOI21_X1   g18019(.A1(new_n17985_), .A2(new_n18118_), .B(new_n18120_), .ZN(new_n18121_));
  NOR2_X1    g18020(.A1(new_n18121_), .A2(new_n18117_), .ZN(new_n18122_));
  OAI21_X1   g18021(.A1(new_n17907_), .A2(new_n18055_), .B(new_n18122_), .ZN(new_n18123_));
  INV_X1     g18022(.I(new_n18122_), .ZN(new_n18124_));
  NAND3_X1   g18023(.A1(new_n17979_), .A2(new_n18054_), .A3(new_n18124_), .ZN(new_n18125_));
  AOI21_X1   g18024(.A1(new_n18123_), .A2(new_n18125_), .B(new_n18050_), .ZN(new_n18126_));
  INV_X1     g18025(.I(new_n18050_), .ZN(new_n18127_));
  AOI21_X1   g18026(.A1(new_n17979_), .A2(new_n18054_), .B(new_n18124_), .ZN(new_n18128_));
  NOR3_X1    g18027(.A1(new_n17907_), .A2(new_n18055_), .A3(new_n18122_), .ZN(new_n18129_));
  NOR3_X1    g18028(.A1(new_n18129_), .A2(new_n18128_), .A3(new_n18127_), .ZN(new_n18130_));
  NOR2_X1    g18029(.A1(new_n18130_), .A2(new_n18126_), .ZN(new_n18131_));
  INV_X1     g18030(.I(new_n18131_), .ZN(new_n18132_));
  OAI21_X1   g18031(.A1(new_n18047_), .A2(new_n18042_), .B(new_n18132_), .ZN(new_n18133_));
  NAND4_X1   g18032(.A1(\result[21] ), .A2(new_n17972_), .A3(new_n18043_), .A4(new_n18131_), .ZN(new_n18134_));
  NAND2_X1   g18033(.A1(new_n18133_), .A2(new_n18134_), .ZN(\result[24] ));
  NAND2_X1   g18034(.A1(new_n17976_), .A2(new_n18043_), .ZN(new_n18136_));
  NOR2_X1    g18035(.A1(new_n17907_), .A2(new_n18055_), .ZN(new_n18137_));
  NOR2_X1    g18036(.A1(new_n18127_), .A2(new_n18117_), .ZN(new_n18138_));
  AOI21_X1   g18037(.A1(new_n18127_), .A2(new_n18117_), .B(new_n18121_), .ZN(new_n18139_));
  AOI21_X1   g18038(.A1(new_n18137_), .A2(new_n18139_), .B(new_n18138_), .ZN(new_n18140_));
  NOR2_X1    g18039(.A1(new_n18102_), .A2(new_n18111_), .ZN(new_n18141_));
  NOR2_X1    g18040(.A1(new_n18141_), .A2(new_n18112_), .ZN(new_n18142_));
  INV_X1     g18041(.I(new_n18066_), .ZN(new_n18143_));
  AOI21_X1   g18042(.A1(new_n18065_), .A2(new_n18143_), .B(new_n18068_), .ZN(new_n18144_));
  NOR2_X1    g18043(.A1(new_n15515_), .A2(new_n4723_), .ZN(new_n18145_));
  OAI22_X1   g18044(.A1(new_n18145_), .A2(\a[20] ), .B1(new_n4725_), .B2(new_n15515_), .ZN(new_n18146_));
  INV_X1     g18045(.I(new_n18146_), .ZN(new_n18147_));
  NOR2_X1    g18046(.A1(new_n10938_), .A2(new_n88_), .ZN(new_n18148_));
  INV_X1     g18047(.I(new_n18148_), .ZN(new_n18149_));
  AOI22_X1   g18048(.A1(new_n10584_), .A2(new_n4406_), .B1(new_n962_), .B2(new_n10949_), .ZN(new_n18150_));
  AOI21_X1   g18049(.A1(new_n18150_), .A2(new_n18149_), .B(new_n82_), .ZN(new_n18151_));
  NAND2_X1   g18050(.A1(new_n12907_), .A2(new_n18151_), .ZN(new_n18152_));
  XNOR2_X1   g18051(.A1(new_n18152_), .A2(new_n18062_), .ZN(new_n18153_));
  NOR2_X1    g18052(.A1(new_n18153_), .A2(new_n18147_), .ZN(new_n18154_));
  AOI21_X1   g18053(.A1(new_n12907_), .A2(new_n18151_), .B(new_n18067_), .ZN(new_n18155_));
  NOR2_X1    g18054(.A1(new_n18152_), .A2(new_n18062_), .ZN(new_n18156_));
  NOR2_X1    g18055(.A1(new_n18155_), .A2(new_n18156_), .ZN(new_n18157_));
  NOR2_X1    g18056(.A1(new_n18157_), .A2(new_n18146_), .ZN(new_n18158_));
  NOR2_X1    g18057(.A1(new_n18158_), .A2(new_n18154_), .ZN(new_n18159_));
  OAI22_X1   g18058(.A1(new_n10577_), .A2(new_n4529_), .B1(new_n4527_), .B2(new_n10961_), .ZN(new_n18160_));
  OAI21_X1   g18059(.A1(new_n79_), .A2(new_n10570_), .B(new_n18160_), .ZN(new_n18161_));
  AOI21_X1   g18060(.A1(new_n18161_), .A2(new_n72_), .B(new_n79_), .ZN(new_n18162_));
  XNOR2_X1   g18061(.A1(new_n14077_), .A2(new_n18162_), .ZN(new_n18163_));
  AND2_X2    g18062(.A1(new_n18159_), .A2(new_n18163_), .Z(new_n18164_));
  NOR2_X1    g18063(.A1(new_n18159_), .A2(new_n18163_), .ZN(new_n18165_));
  NOR2_X1    g18064(.A1(new_n18164_), .A2(new_n18165_), .ZN(new_n18166_));
  NOR2_X1    g18065(.A1(new_n18144_), .A2(new_n18166_), .ZN(new_n18167_));
  INV_X1     g18066(.I(new_n18144_), .ZN(new_n18168_));
  XNOR2_X1   g18067(.A1(new_n18159_), .A2(new_n18163_), .ZN(new_n18169_));
  NOR2_X1    g18068(.A1(new_n18168_), .A2(new_n18169_), .ZN(new_n18170_));
  NOR2_X1    g18069(.A1(new_n18170_), .A2(new_n18167_), .ZN(new_n18171_));
  INV_X1     g18070(.I(new_n18171_), .ZN(new_n18172_));
  NOR2_X1    g18071(.A1(new_n18072_), .A2(new_n18084_), .ZN(new_n18173_));
  NOR2_X1    g18072(.A1(new_n18173_), .A2(new_n18085_), .ZN(new_n18174_));
  AOI22_X1   g18073(.A1(new_n10971_), .A2(new_n4613_), .B1(new_n4767_), .B2(new_n14274_), .ZN(new_n18175_));
  AOI21_X1   g18074(.A1(new_n117_), .A2(new_n14603_), .B(new_n18175_), .ZN(new_n18176_));
  OAI21_X1   g18075(.A1(new_n18176_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n18177_));
  XNOR2_X1   g18076(.A1(new_n14601_), .A2(new_n18177_), .ZN(new_n18178_));
  INV_X1     g18077(.I(new_n18178_), .ZN(new_n18179_));
  XOR2_X1    g18078(.A1(new_n18174_), .A2(new_n18179_), .Z(new_n18180_));
  INV_X1     g18079(.I(new_n18180_), .ZN(new_n18181_));
  NOR3_X1    g18080(.A1(new_n18173_), .A2(new_n18085_), .A3(new_n18179_), .ZN(new_n18182_));
  NOR2_X1    g18081(.A1(new_n18174_), .A2(new_n18178_), .ZN(new_n18183_));
  NOR2_X1    g18082(.A1(new_n18183_), .A2(new_n18182_), .ZN(new_n18184_));
  NOR2_X1    g18083(.A1(new_n18184_), .A2(new_n18172_), .ZN(new_n18185_));
  AOI21_X1   g18084(.A1(new_n18181_), .A2(new_n18172_), .B(new_n18185_), .ZN(new_n18186_));
  INV_X1     g18085(.I(new_n18095_), .ZN(new_n18187_));
  AOI21_X1   g18086(.A1(new_n18187_), .A2(new_n18099_), .B(new_n18096_), .ZN(new_n18188_));
  OAI22_X1   g18087(.A1(new_n15313_), .A2(new_n4981_), .B1(new_n1239_), .B2(new_n15305_), .ZN(new_n18189_));
  AOI21_X1   g18088(.A1(new_n18189_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n18190_));
  XNOR2_X1   g18089(.A1(new_n15312_), .A2(new_n18190_), .ZN(new_n18191_));
  AND2_X2    g18090(.A1(new_n18188_), .A2(new_n18191_), .Z(new_n18192_));
  NOR2_X1    g18091(.A1(new_n18188_), .A2(new_n18191_), .ZN(new_n18193_));
  NOR2_X1    g18092(.A1(new_n18192_), .A2(new_n18193_), .ZN(new_n18194_));
  NOR2_X1    g18093(.A1(new_n18194_), .A2(new_n18186_), .ZN(new_n18195_));
  INV_X1     g18094(.I(new_n18186_), .ZN(new_n18196_));
  XNOR2_X1   g18095(.A1(new_n18188_), .A2(new_n18191_), .ZN(new_n18197_));
  NOR2_X1    g18096(.A1(new_n18197_), .A2(new_n18196_), .ZN(new_n18198_));
  NOR2_X1    g18097(.A1(new_n18195_), .A2(new_n18198_), .ZN(new_n18199_));
  NAND2_X1   g18098(.A1(new_n18199_), .A2(new_n18142_), .ZN(new_n18200_));
  INV_X1     g18099(.I(new_n18142_), .ZN(new_n18201_));
  OAI21_X1   g18100(.A1(new_n18195_), .A2(new_n18198_), .B(new_n18201_), .ZN(new_n18202_));
  AOI21_X1   g18101(.A1(new_n18200_), .A2(new_n18202_), .B(new_n18140_), .ZN(new_n18203_));
  XOR2_X1    g18102(.A1(new_n18136_), .A2(new_n18203_), .Z(new_n18204_));
  XOR2_X1    g18103(.A1(new_n18204_), .A2(new_n18131_), .Z(\result[25] ));
  INV_X1     g18104(.I(new_n18203_), .ZN(new_n18206_));
  AOI21_X1   g18105(.A1(new_n18133_), .A2(new_n18134_), .B(new_n18206_), .ZN(new_n18207_));
  INV_X1     g18106(.I(new_n18164_), .ZN(new_n18208_));
  AOI21_X1   g18107(.A1(new_n18168_), .A2(new_n18208_), .B(new_n18165_), .ZN(new_n18209_));
  NOR2_X1    g18108(.A1(new_n10577_), .A2(new_n511_), .ZN(new_n18210_));
  INV_X1     g18109(.I(new_n18210_), .ZN(new_n18211_));
  NOR2_X1    g18110(.A1(new_n10953_), .A2(new_n4545_), .ZN(new_n18212_));
  AOI21_X1   g18111(.A1(new_n18211_), .A2(new_n18212_), .B(new_n82_), .ZN(new_n18213_));
  NAND2_X1   g18112(.A1(new_n15444_), .A2(new_n18213_), .ZN(new_n18214_));
  INV_X1     g18113(.I(new_n18214_), .ZN(new_n18215_));
  INV_X1     g18114(.I(new_n18155_), .ZN(new_n18216_));
  AOI21_X1   g18115(.A1(new_n18216_), .A2(new_n18147_), .B(new_n18156_), .ZN(new_n18217_));
  INV_X1     g18116(.I(new_n18217_), .ZN(new_n18218_));
  OAI22_X1   g18117(.A1(new_n10564_), .A2(new_n79_), .B1(new_n4530_), .B2(new_n18008_), .ZN(new_n18219_));
  AOI21_X1   g18118(.A1(new_n18219_), .A2(new_n72_), .B(new_n79_), .ZN(new_n18220_));
  AND2_X2    g18119(.A1(new_n10976_), .A2(new_n18220_), .Z(new_n18221_));
  NOR2_X1    g18120(.A1(new_n10976_), .A2(new_n18220_), .ZN(new_n18222_));
  NOR2_X1    g18121(.A1(new_n18221_), .A2(new_n18222_), .ZN(new_n18223_));
  XOR2_X1    g18122(.A1(new_n18223_), .A2(new_n18218_), .Z(new_n18224_));
  NOR2_X1    g18123(.A1(new_n18224_), .A2(new_n18215_), .ZN(new_n18225_));
  NOR3_X1    g18124(.A1(new_n18221_), .A2(new_n18218_), .A3(new_n18222_), .ZN(new_n18226_));
  NOR2_X1    g18125(.A1(new_n18223_), .A2(new_n18217_), .ZN(new_n18227_));
  NOR2_X1    g18126(.A1(new_n18227_), .A2(new_n18226_), .ZN(new_n18228_));
  NOR2_X1    g18127(.A1(new_n18228_), .A2(new_n18214_), .ZN(new_n18229_));
  NOR2_X1    g18128(.A1(new_n18225_), .A2(new_n18229_), .ZN(new_n18230_));
  OAI22_X1   g18129(.A1(new_n14886_), .A2(new_n1128_), .B1(new_n4782_), .B2(new_n14598_), .ZN(new_n18231_));
  AOI21_X1   g18130(.A1(new_n18231_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n18232_));
  XOR2_X1    g18131(.A1(new_n14891_), .A2(new_n18232_), .Z(new_n18233_));
  INV_X1     g18132(.I(new_n18233_), .ZN(new_n18234_));
  NOR2_X1    g18133(.A1(new_n18230_), .A2(new_n18234_), .ZN(new_n18235_));
  INV_X1     g18134(.I(new_n18235_), .ZN(new_n18236_));
  NAND2_X1   g18135(.A1(new_n18230_), .A2(new_n18234_), .ZN(new_n18237_));
  AOI21_X1   g18136(.A1(new_n18236_), .A2(new_n18237_), .B(new_n18209_), .ZN(new_n18238_));
  INV_X1     g18137(.I(new_n18209_), .ZN(new_n18239_));
  XOR2_X1    g18138(.A1(new_n18230_), .A2(new_n18233_), .Z(new_n18240_));
  NOR2_X1    g18139(.A1(new_n18240_), .A2(new_n18239_), .ZN(new_n18241_));
  NOR2_X1    g18140(.A1(new_n18241_), .A2(new_n18238_), .ZN(new_n18242_));
  NOR2_X1    g18141(.A1(new_n18182_), .A2(new_n18171_), .ZN(new_n18243_));
  OAI22_X1   g18142(.A1(new_n15305_), .A2(new_n4902_), .B1(new_n15114_), .B2(new_n1973_), .ZN(new_n18244_));
  OAI21_X1   g18143(.A1(new_n1239_), .A2(new_n15515_), .B(new_n18244_), .ZN(new_n18245_));
  AOI21_X1   g18144(.A1(new_n18245_), .A2(new_n68_), .B(new_n1239_), .ZN(new_n18246_));
  XOR2_X1    g18145(.A1(new_n15518_), .A2(new_n18246_), .Z(new_n18247_));
  INV_X1     g18146(.I(new_n18247_), .ZN(new_n18248_));
  NOR3_X1    g18147(.A1(new_n18243_), .A2(new_n18248_), .A3(new_n18183_), .ZN(new_n18249_));
  NOR2_X1    g18148(.A1(new_n18243_), .A2(new_n18183_), .ZN(new_n18250_));
  NOR2_X1    g18149(.A1(new_n18250_), .A2(new_n18247_), .ZN(new_n18251_));
  NOR2_X1    g18150(.A1(new_n18251_), .A2(new_n18249_), .ZN(new_n18252_));
  NOR2_X1    g18151(.A1(new_n18242_), .A2(new_n18252_), .ZN(new_n18253_));
  INV_X1     g18152(.I(new_n18242_), .ZN(new_n18254_));
  XOR2_X1    g18153(.A1(new_n18250_), .A2(new_n18248_), .Z(new_n18255_));
  NOR2_X1    g18154(.A1(new_n18254_), .A2(new_n18255_), .ZN(new_n18256_));
  NOR2_X1    g18155(.A1(new_n18256_), .A2(new_n18253_), .ZN(new_n18257_));
  NOR2_X1    g18156(.A1(new_n18192_), .A2(new_n18196_), .ZN(new_n18258_));
  NOR2_X1    g18157(.A1(new_n18258_), .A2(new_n18193_), .ZN(new_n18259_));
  NAND2_X1   g18158(.A1(new_n18257_), .A2(new_n18259_), .ZN(new_n18260_));
  INV_X1     g18159(.I(new_n18260_), .ZN(new_n18261_));
  NOR2_X1    g18160(.A1(new_n18257_), .A2(new_n18259_), .ZN(new_n18262_));
  NOR2_X1    g18161(.A1(new_n18261_), .A2(new_n18262_), .ZN(new_n18263_));
  XOR2_X1    g18162(.A1(new_n18199_), .A2(new_n18201_), .Z(new_n18264_));
  NOR2_X1    g18163(.A1(new_n18264_), .A2(new_n18263_), .ZN(new_n18265_));
  XOR2_X1    g18164(.A1(new_n18265_), .A2(new_n18202_), .Z(new_n18266_));
  XNOR2_X1   g18165(.A1(new_n18140_), .A2(new_n18266_), .ZN(new_n18267_));
  INV_X1     g18166(.I(new_n18267_), .ZN(new_n18268_));
  XOR2_X1    g18167(.A1(new_n18207_), .A2(new_n18268_), .Z(\result[26] ));
  NAND2_X1   g18168(.A1(new_n18263_), .A2(new_n18199_), .ZN(new_n18270_));
  OAI21_X1   g18169(.A1(new_n18263_), .A2(new_n18199_), .B(new_n18142_), .ZN(new_n18271_));
  NAND2_X1   g18170(.A1(new_n18271_), .A2(new_n18270_), .ZN(new_n18272_));
  OAI21_X1   g18171(.A1(new_n18209_), .A2(new_n18235_), .B(new_n18237_), .ZN(new_n18273_));
  INV_X1     g18172(.I(new_n18273_), .ZN(new_n18274_));
  INV_X1     g18173(.I(new_n18226_), .ZN(new_n18275_));
  AOI21_X1   g18174(.A1(new_n18275_), .A2(new_n18214_), .B(new_n18227_), .ZN(new_n18276_));
  NOR2_X1    g18175(.A1(new_n10577_), .A2(new_n88_), .ZN(new_n18277_));
  INV_X1     g18176(.I(new_n18277_), .ZN(new_n18278_));
  AOI22_X1   g18177(.A1(new_n10962_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n10949_), .ZN(new_n18279_));
  AOI21_X1   g18178(.A1(new_n18278_), .A2(new_n18279_), .B(new_n82_), .ZN(new_n18280_));
  NAND2_X1   g18179(.A1(new_n15071_), .A2(new_n18280_), .ZN(new_n18281_));
  INV_X1     g18180(.I(new_n18281_), .ZN(new_n18282_));
  XOR2_X1    g18181(.A1(new_n18276_), .A2(new_n18282_), .Z(new_n18283_));
  NOR2_X1    g18182(.A1(new_n18283_), .A2(new_n18215_), .ZN(new_n18284_));
  AND2_X2    g18183(.A1(new_n18276_), .A2(new_n18281_), .Z(new_n18285_));
  NOR2_X1    g18184(.A1(new_n18276_), .A2(new_n18281_), .ZN(new_n18286_));
  NOR2_X1    g18185(.A1(new_n18285_), .A2(new_n18286_), .ZN(new_n18287_));
  NOR2_X1    g18186(.A1(new_n18287_), .A2(new_n18214_), .ZN(new_n18288_));
  NOR2_X1    g18187(.A1(new_n18288_), .A2(new_n18284_), .ZN(new_n18289_));
  AOI22_X1   g18188(.A1(new_n14888_), .A2(new_n4767_), .B1(new_n4613_), .B2(new_n14603_), .ZN(new_n18290_));
  AOI21_X1   g18189(.A1(new_n117_), .A2(new_n15115_), .B(new_n18290_), .ZN(new_n18291_));
  OAI21_X1   g18190(.A1(new_n18291_), .A2(\a[26] ), .B(new_n117_), .ZN(new_n18292_));
  XNOR2_X1   g18191(.A1(new_n15125_), .A2(new_n18292_), .ZN(new_n18293_));
  AOI22_X1   g18192(.A1(new_n10971_), .A2(new_n4526_), .B1(new_n4570_), .B2(new_n10571_), .ZN(new_n18294_));
  AOI21_X1   g18193(.A1(new_n101_), .A2(new_n14274_), .B(new_n18294_), .ZN(new_n18295_));
  OAI21_X1   g18194(.A1(new_n18295_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n18296_));
  XOR2_X1    g18195(.A1(new_n14280_), .A2(new_n18296_), .Z(new_n18297_));
  INV_X1     g18196(.I(new_n18297_), .ZN(new_n18298_));
  XOR2_X1    g18197(.A1(new_n18293_), .A2(new_n18298_), .Z(new_n18299_));
  NOR2_X1    g18198(.A1(new_n18289_), .A2(new_n18299_), .ZN(new_n18300_));
  AND2_X2    g18199(.A1(new_n18293_), .A2(new_n18297_), .Z(new_n18301_));
  NOR2_X1    g18200(.A1(new_n18293_), .A2(new_n18297_), .ZN(new_n18302_));
  NOR2_X1    g18201(.A1(new_n18301_), .A2(new_n18302_), .ZN(new_n18303_));
  NOR3_X1    g18202(.A1(new_n18303_), .A2(new_n18284_), .A3(new_n18288_), .ZN(new_n18304_));
  NOR2_X1    g18203(.A1(new_n18300_), .A2(new_n18304_), .ZN(new_n18305_));
  INV_X1     g18204(.I(new_n18305_), .ZN(new_n18306_));
  NAND2_X1   g18205(.A1(new_n15515_), .A2(new_n4412_), .ZN(new_n18307_));
  NOR2_X1    g18206(.A1(new_n4410_), .A2(new_n247_), .ZN(new_n18308_));
  AOI21_X1   g18207(.A1(new_n15675_), .A2(new_n18308_), .B(\a[23] ), .ZN(new_n18309_));
  AOI21_X1   g18208(.A1(new_n18309_), .A2(new_n18307_), .B(new_n1239_), .ZN(new_n18310_));
  XNOR2_X1   g18209(.A1(new_n15678_), .A2(new_n18310_), .ZN(new_n18311_));
  INV_X1     g18210(.I(new_n18311_), .ZN(new_n18312_));
  NOR2_X1    g18211(.A1(new_n18306_), .A2(new_n18312_), .ZN(new_n18313_));
  NOR2_X1    g18212(.A1(new_n18305_), .A2(new_n18311_), .ZN(new_n18314_));
  NOR2_X1    g18213(.A1(new_n18313_), .A2(new_n18314_), .ZN(new_n18315_));
  NOR2_X1    g18214(.A1(new_n18315_), .A2(new_n18274_), .ZN(new_n18316_));
  XOR2_X1    g18215(.A1(new_n18305_), .A2(new_n18312_), .Z(new_n18317_));
  NOR2_X1    g18216(.A1(new_n18317_), .A2(new_n18273_), .ZN(new_n18318_));
  NOR2_X1    g18217(.A1(new_n18316_), .A2(new_n18318_), .ZN(new_n18319_));
  NOR2_X1    g18218(.A1(new_n18242_), .A2(new_n18249_), .ZN(new_n18320_));
  NOR2_X1    g18219(.A1(new_n18320_), .A2(new_n18251_), .ZN(new_n18321_));
  NOR2_X1    g18220(.A1(new_n18319_), .A2(new_n18321_), .ZN(new_n18322_));
  OAI21_X1   g18221(.A1(new_n18140_), .A2(new_n18272_), .B(new_n18322_), .ZN(new_n18323_));
  NOR3_X1    g18222(.A1(new_n18140_), .A2(new_n18272_), .A3(new_n18322_), .ZN(new_n18324_));
  INV_X1     g18223(.I(new_n18324_), .ZN(new_n18325_));
  AOI21_X1   g18224(.A1(new_n18325_), .A2(new_n18323_), .B(new_n18261_), .ZN(new_n18326_));
  INV_X1     g18225(.I(new_n18323_), .ZN(new_n18327_));
  NOR3_X1    g18226(.A1(new_n18327_), .A2(new_n18260_), .A3(new_n18324_), .ZN(new_n18328_));
  NOR2_X1    g18227(.A1(new_n18326_), .A2(new_n18328_), .ZN(new_n18329_));
  NAND4_X1   g18228(.A1(\result[24] ), .A2(new_n18203_), .A3(new_n18268_), .A4(new_n18329_), .ZN(new_n18330_));
  AOI21_X1   g18229(.A1(new_n17976_), .A2(new_n18043_), .B(new_n18131_), .ZN(new_n18331_));
  NOR3_X1    g18230(.A1(new_n18047_), .A2(new_n18132_), .A3(new_n18042_), .ZN(new_n18332_));
  OAI21_X1   g18231(.A1(new_n18332_), .A2(new_n18331_), .B(new_n18203_), .ZN(new_n18333_));
  OAI21_X1   g18232(.A1(new_n18327_), .A2(new_n18324_), .B(new_n18260_), .ZN(new_n18334_));
  NAND3_X1   g18233(.A1(new_n18325_), .A2(new_n18261_), .A3(new_n18323_), .ZN(new_n18335_));
  NAND2_X1   g18234(.A1(new_n18334_), .A2(new_n18335_), .ZN(new_n18336_));
  OAI21_X1   g18235(.A1(new_n18333_), .A2(new_n18267_), .B(new_n18336_), .ZN(new_n18337_));
  NAND2_X1   g18236(.A1(new_n18337_), .A2(new_n18330_), .ZN(\result[27] ));
  NOR2_X1    g18237(.A1(new_n18333_), .A2(new_n18267_), .ZN(new_n18339_));
  NOR2_X1    g18238(.A1(new_n18140_), .A2(new_n18272_), .ZN(new_n18340_));
  INV_X1     g18239(.I(new_n18319_), .ZN(new_n18341_));
  AOI21_X1   g18240(.A1(new_n18319_), .A2(new_n18260_), .B(new_n18321_), .ZN(new_n18342_));
  AOI22_X1   g18241(.A1(new_n18340_), .A2(new_n18342_), .B1(new_n18261_), .B2(new_n18341_), .ZN(new_n18343_));
  INV_X1     g18242(.I(new_n18314_), .ZN(new_n18344_));
  OAI21_X1   g18243(.A1(new_n18274_), .A2(new_n18313_), .B(new_n18344_), .ZN(new_n18345_));
  INV_X1     g18244(.I(new_n18301_), .ZN(new_n18346_));
  AOI21_X1   g18245(.A1(new_n18289_), .A2(new_n18346_), .B(new_n18302_), .ZN(new_n18347_));
  NOR2_X1    g18246(.A1(new_n15515_), .A2(new_n4413_), .ZN(new_n18348_));
  OAI22_X1   g18247(.A1(new_n18348_), .A2(\a[23] ), .B1(new_n4415_), .B2(new_n15515_), .ZN(new_n18349_));
  INV_X1     g18248(.I(new_n18349_), .ZN(new_n18350_));
  NAND2_X1   g18249(.A1(new_n10962_), .A2(new_n87_), .ZN(new_n18351_));
  AOI22_X1   g18250(.A1(new_n10958_), .A2(new_n4406_), .B1(new_n962_), .B2(new_n10571_), .ZN(new_n18352_));
  AOI21_X1   g18251(.A1(new_n18352_), .A2(new_n18351_), .B(new_n82_), .ZN(new_n18353_));
  AOI21_X1   g18252(.A1(new_n14077_), .A2(new_n18353_), .B(new_n18350_), .ZN(new_n18354_));
  NAND2_X1   g18253(.A1(new_n14077_), .A2(new_n18353_), .ZN(new_n18355_));
  NOR2_X1    g18254(.A1(new_n18355_), .A2(new_n18349_), .ZN(new_n18356_));
  NOR2_X1    g18255(.A1(new_n18356_), .A2(new_n18354_), .ZN(new_n18357_));
  NOR2_X1    g18256(.A1(new_n18357_), .A2(new_n18214_), .ZN(new_n18358_));
  XOR2_X1    g18257(.A1(new_n18355_), .A2(new_n18350_), .Z(new_n18359_));
  NOR2_X1    g18258(.A1(new_n18359_), .A2(new_n18215_), .ZN(new_n18360_));
  NOR2_X1    g18259(.A1(new_n18360_), .A2(new_n18358_), .ZN(new_n18361_));
  INV_X1     g18260(.I(new_n18285_), .ZN(new_n18362_));
  AOI21_X1   g18261(.A1(new_n18362_), .A2(new_n18214_), .B(new_n18286_), .ZN(new_n18363_));
  AOI22_X1   g18262(.A1(new_n10971_), .A2(new_n4570_), .B1(new_n4526_), .B2(new_n14274_), .ZN(new_n18364_));
  AOI21_X1   g18263(.A1(new_n101_), .A2(new_n14603_), .B(new_n18364_), .ZN(new_n18365_));
  OAI21_X1   g18264(.A1(new_n18365_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n18366_));
  XNOR2_X1   g18265(.A1(new_n14601_), .A2(new_n18366_), .ZN(new_n18367_));
  AND2_X2    g18266(.A1(new_n18363_), .A2(new_n18367_), .Z(new_n18368_));
  INV_X1     g18267(.I(new_n18368_), .ZN(new_n18369_));
  NOR2_X1    g18268(.A1(new_n18363_), .A2(new_n18367_), .ZN(new_n18370_));
  INV_X1     g18269(.I(new_n18370_), .ZN(new_n18371_));
  AOI21_X1   g18270(.A1(new_n18369_), .A2(new_n18371_), .B(new_n18361_), .ZN(new_n18372_));
  INV_X1     g18271(.I(new_n18361_), .ZN(new_n18373_));
  XNOR2_X1   g18272(.A1(new_n18363_), .A2(new_n18367_), .ZN(new_n18374_));
  NOR2_X1    g18273(.A1(new_n18374_), .A2(new_n18373_), .ZN(new_n18375_));
  OAI22_X1   g18274(.A1(new_n4612_), .A2(new_n14886_), .B1(new_n15114_), .B2(new_n4781_), .ZN(new_n18376_));
  OAI21_X1   g18275(.A1(new_n1128_), .A2(new_n15305_), .B(new_n18376_), .ZN(new_n18377_));
  AOI21_X1   g18276(.A1(new_n18377_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n18378_));
  XNOR2_X1   g18277(.A1(new_n15312_), .A2(new_n18378_), .ZN(new_n18379_));
  INV_X1     g18278(.I(new_n18379_), .ZN(new_n18380_));
  NOR3_X1    g18279(.A1(new_n18372_), .A2(new_n18375_), .A3(new_n18380_), .ZN(new_n18381_));
  NOR2_X1    g18280(.A1(new_n18372_), .A2(new_n18375_), .ZN(new_n18382_));
  NOR2_X1    g18281(.A1(new_n18382_), .A2(new_n18379_), .ZN(new_n18383_));
  NOR2_X1    g18282(.A1(new_n18383_), .A2(new_n18381_), .ZN(new_n18384_));
  NOR2_X1    g18283(.A1(new_n18384_), .A2(new_n18347_), .ZN(new_n18385_));
  INV_X1     g18284(.I(new_n18347_), .ZN(new_n18386_));
  XOR2_X1    g18285(.A1(new_n18382_), .A2(new_n18380_), .Z(new_n18387_));
  NOR2_X1    g18286(.A1(new_n18387_), .A2(new_n18386_), .ZN(new_n18388_));
  NOR2_X1    g18287(.A1(new_n18388_), .A2(new_n18385_), .ZN(new_n18389_));
  XOR2_X1    g18288(.A1(new_n18389_), .A2(new_n18345_), .Z(new_n18390_));
  NOR2_X1    g18289(.A1(new_n18343_), .A2(new_n18390_), .ZN(new_n18391_));
  XOR2_X1    g18290(.A1(new_n18336_), .A2(new_n18391_), .Z(new_n18392_));
  XOR2_X1    g18291(.A1(new_n18392_), .A2(new_n18339_), .Z(\result[28] ));
  INV_X1     g18292(.I(new_n18391_), .ZN(new_n18394_));
  AOI21_X1   g18293(.A1(new_n18337_), .A2(new_n18330_), .B(new_n18394_), .ZN(new_n18395_));
  OAI21_X1   g18294(.A1(new_n18388_), .A2(new_n18385_), .B(new_n18345_), .ZN(new_n18396_));
  NAND2_X1   g18295(.A1(new_n18369_), .A2(new_n18373_), .ZN(new_n18397_));
  NAND2_X1   g18296(.A1(new_n18397_), .A2(new_n18371_), .ZN(new_n18398_));
  INV_X1     g18297(.I(new_n18354_), .ZN(new_n18399_));
  AOI21_X1   g18298(.A1(new_n18399_), .A2(new_n18215_), .B(new_n18356_), .ZN(new_n18400_));
  NOR2_X1    g18299(.A1(new_n10564_), .A2(new_n511_), .ZN(new_n18401_));
  OAI21_X1   g18300(.A1(new_n10570_), .A2(new_n10961_), .B(new_n14580_), .ZN(new_n18402_));
  OAI21_X1   g18301(.A1(new_n18401_), .A2(new_n18402_), .B(new_n961_), .ZN(new_n18403_));
  NOR2_X1    g18302(.A1(new_n10976_), .A2(new_n18403_), .ZN(new_n18404_));
  INV_X1     g18303(.I(new_n18404_), .ZN(new_n18405_));
  OAI22_X1   g18304(.A1(new_n14886_), .A2(new_n79_), .B1(new_n4530_), .B2(new_n14598_), .ZN(new_n18406_));
  AOI21_X1   g18305(.A1(new_n18406_), .A2(new_n72_), .B(new_n79_), .ZN(new_n18407_));
  XOR2_X1    g18306(.A1(new_n14891_), .A2(new_n18407_), .Z(new_n18408_));
  XOR2_X1    g18307(.A1(new_n18408_), .A2(new_n18405_), .Z(new_n18409_));
  NOR2_X1    g18308(.A1(new_n18409_), .A2(new_n18400_), .ZN(new_n18410_));
  INV_X1     g18309(.I(new_n18400_), .ZN(new_n18411_));
  AND2_X2    g18310(.A1(new_n18408_), .A2(new_n18404_), .Z(new_n18412_));
  NOR2_X1    g18311(.A1(new_n18408_), .A2(new_n18404_), .ZN(new_n18413_));
  NOR2_X1    g18312(.A1(new_n18412_), .A2(new_n18413_), .ZN(new_n18414_));
  NOR2_X1    g18313(.A1(new_n18414_), .A2(new_n18411_), .ZN(new_n18415_));
  NOR2_X1    g18314(.A1(new_n18415_), .A2(new_n18410_), .ZN(new_n18416_));
  NOR2_X1    g18315(.A1(new_n15305_), .A2(new_n15114_), .ZN(new_n18417_));
  OAI22_X1   g18316(.A1(new_n18417_), .A2(new_n4782_), .B1(new_n1128_), .B2(new_n15515_), .ZN(new_n18418_));
  AOI21_X1   g18317(.A1(new_n18418_), .A2(new_n65_), .B(new_n1128_), .ZN(new_n18419_));
  XOR2_X1    g18318(.A1(new_n15518_), .A2(new_n18419_), .Z(new_n18420_));
  INV_X1     g18319(.I(new_n18420_), .ZN(new_n18421_));
  NOR2_X1    g18320(.A1(new_n18421_), .A2(new_n18416_), .ZN(new_n18422_));
  INV_X1     g18321(.I(new_n18422_), .ZN(new_n18423_));
  NAND2_X1   g18322(.A1(new_n18421_), .A2(new_n18416_), .ZN(new_n18424_));
  NAND2_X1   g18323(.A1(new_n18423_), .A2(new_n18424_), .ZN(new_n18425_));
  XOR2_X1    g18324(.A1(new_n18416_), .A2(new_n18420_), .Z(new_n18426_));
  NOR2_X1    g18325(.A1(new_n18398_), .A2(new_n18426_), .ZN(new_n18427_));
  AOI21_X1   g18326(.A1(new_n18398_), .A2(new_n18425_), .B(new_n18427_), .ZN(new_n18428_));
  NOR2_X1    g18327(.A1(new_n18381_), .A2(new_n18347_), .ZN(new_n18429_));
  NOR2_X1    g18328(.A1(new_n18429_), .A2(new_n18383_), .ZN(new_n18430_));
  NAND2_X1   g18329(.A1(new_n18430_), .A2(new_n18428_), .ZN(new_n18431_));
  INV_X1     g18330(.I(new_n18431_), .ZN(new_n18432_));
  NOR2_X1    g18331(.A1(new_n18430_), .A2(new_n18428_), .ZN(new_n18433_));
  NOR2_X1    g18332(.A1(new_n18432_), .A2(new_n18433_), .ZN(new_n18434_));
  NOR2_X1    g18333(.A1(new_n18390_), .A2(new_n18434_), .ZN(new_n18435_));
  XOR2_X1    g18334(.A1(new_n18435_), .A2(new_n18396_), .Z(new_n18436_));
  XNOR2_X1   g18335(.A1(new_n18343_), .A2(new_n18436_), .ZN(new_n18437_));
  INV_X1     g18336(.I(new_n18437_), .ZN(new_n18438_));
  XOR2_X1    g18337(.A1(new_n18395_), .A2(new_n18438_), .Z(\result[29] ));
  NAND2_X1   g18338(.A1(new_n18395_), .A2(new_n18438_), .ZN(new_n18440_));
  NAND2_X1   g18339(.A1(new_n18434_), .A2(new_n18389_), .ZN(new_n18441_));
  NOR2_X1    g18340(.A1(new_n18434_), .A2(new_n18389_), .ZN(new_n18442_));
  OAI21_X1   g18341(.A1(new_n18345_), .A2(new_n18442_), .B(new_n18441_), .ZN(new_n18443_));
  NOR2_X1    g18342(.A1(new_n18343_), .A2(new_n18443_), .ZN(new_n18444_));
  NOR2_X1    g18343(.A1(new_n18412_), .A2(new_n18400_), .ZN(new_n18445_));
  NOR2_X1    g18344(.A1(new_n18445_), .A2(new_n18413_), .ZN(new_n18446_));
  INV_X1     g18345(.I(new_n18446_), .ZN(new_n18447_));
  NAND2_X1   g18346(.A1(new_n10971_), .A2(new_n87_), .ZN(new_n18448_));
  AOI22_X1   g18347(.A1(new_n14274_), .A2(new_n962_), .B1(new_n4406_), .B2(new_n10571_), .ZN(new_n18449_));
  AOI21_X1   g18348(.A1(new_n18448_), .A2(new_n18449_), .B(new_n82_), .ZN(new_n18450_));
  NAND2_X1   g18349(.A1(new_n14280_), .A2(new_n18450_), .ZN(new_n18451_));
  XNOR2_X1   g18350(.A1(new_n18451_), .A2(new_n18404_), .ZN(new_n18452_));
  INV_X1     g18351(.I(new_n18452_), .ZN(new_n18453_));
  XOR2_X1    g18352(.A1(new_n18451_), .A2(new_n18404_), .Z(new_n18454_));
  NOR2_X1    g18353(.A1(new_n18447_), .A2(new_n18454_), .ZN(new_n18455_));
  AOI21_X1   g18354(.A1(new_n18447_), .A2(new_n18453_), .B(new_n18455_), .ZN(new_n18456_));
  INV_X1     g18355(.I(new_n18456_), .ZN(new_n18457_));
  NOR2_X1    g18356(.A1(new_n15511_), .A2(new_n4781_), .ZN(new_n18458_));
  INV_X1     g18357(.I(new_n18458_), .ZN(new_n18459_));
  NOR2_X1    g18358(.A1(new_n4613_), .A2(new_n117_), .ZN(new_n18460_));
  AOI21_X1   g18359(.A1(new_n15675_), .A2(new_n18460_), .B(\a[26] ), .ZN(new_n18461_));
  AOI21_X1   g18360(.A1(new_n18461_), .A2(new_n18459_), .B(new_n1128_), .ZN(new_n18462_));
  INV_X1     g18361(.I(new_n18462_), .ZN(new_n18463_));
  NOR2_X1    g18362(.A1(new_n15678_), .A2(new_n18463_), .ZN(new_n18464_));
  NAND2_X1   g18363(.A1(new_n15678_), .A2(new_n18463_), .ZN(new_n18465_));
  INV_X1     g18364(.I(new_n18465_), .ZN(new_n18466_));
  AOI22_X1   g18365(.A1(new_n14888_), .A2(new_n4526_), .B1(new_n4570_), .B2(new_n14603_), .ZN(new_n18467_));
  AOI21_X1   g18366(.A1(new_n101_), .A2(new_n15115_), .B(new_n18467_), .ZN(new_n18468_));
  OAI21_X1   g18367(.A1(new_n18468_), .A2(\a[29] ), .B(new_n101_), .ZN(new_n18469_));
  XNOR2_X1   g18368(.A1(new_n15125_), .A2(new_n18469_), .ZN(new_n18470_));
  INV_X1     g18369(.I(new_n18470_), .ZN(new_n18471_));
  NOR3_X1    g18370(.A1(new_n18471_), .A2(new_n18464_), .A3(new_n18466_), .ZN(new_n18472_));
  NOR2_X1    g18371(.A1(new_n18466_), .A2(new_n18464_), .ZN(new_n18473_));
  NOR2_X1    g18372(.A1(new_n18473_), .A2(new_n18470_), .ZN(new_n18474_));
  OAI21_X1   g18373(.A1(new_n18472_), .A2(new_n18474_), .B(new_n18457_), .ZN(new_n18475_));
  XNOR2_X1   g18374(.A1(new_n18473_), .A2(new_n18470_), .ZN(new_n18476_));
  OAI21_X1   g18375(.A1(new_n18457_), .A2(new_n18476_), .B(new_n18475_), .ZN(new_n18477_));
  INV_X1     g18376(.I(new_n18477_), .ZN(new_n18478_));
  NAND2_X1   g18377(.A1(new_n18398_), .A2(new_n18423_), .ZN(new_n18479_));
  NAND2_X1   g18378(.A1(new_n18479_), .A2(new_n18424_), .ZN(new_n18480_));
  INV_X1     g18379(.I(new_n18480_), .ZN(new_n18481_));
  NOR2_X1    g18380(.A1(new_n18481_), .A2(new_n18478_), .ZN(new_n18482_));
  INV_X1     g18381(.I(new_n18482_), .ZN(new_n18483_));
  NOR2_X1    g18382(.A1(new_n18444_), .A2(new_n18483_), .ZN(new_n18484_));
  INV_X1     g18383(.I(new_n18484_), .ZN(new_n18485_));
  NAND2_X1   g18384(.A1(new_n18444_), .A2(new_n18483_), .ZN(new_n18486_));
  AOI21_X1   g18385(.A1(new_n18485_), .A2(new_n18486_), .B(new_n18432_), .ZN(new_n18487_));
  NAND3_X1   g18386(.A1(new_n18485_), .A2(new_n18432_), .A3(new_n18486_), .ZN(new_n18488_));
  INV_X1     g18387(.I(new_n18488_), .ZN(new_n18489_));
  NOR2_X1    g18388(.A1(new_n18489_), .A2(new_n18487_), .ZN(new_n18490_));
  XOR2_X1    g18389(.A1(new_n18440_), .A2(new_n18490_), .Z(\result[30] ));
  NOR2_X1    g18390(.A1(new_n18431_), .A2(new_n18478_), .ZN(new_n18492_));
  NOR2_X1    g18391(.A1(new_n18432_), .A2(new_n18477_), .ZN(new_n18493_));
  NOR4_X1    g18392(.A1(new_n18343_), .A2(new_n18443_), .A3(new_n18481_), .A4(new_n18493_), .ZN(new_n18494_));
  NOR2_X1    g18393(.A1(new_n18494_), .A2(new_n18492_), .ZN(new_n18495_));
  NOR2_X1    g18394(.A1(new_n18451_), .A2(new_n18404_), .ZN(new_n18496_));
  NOR2_X1    g18395(.A1(new_n18452_), .A2(new_n72_), .ZN(new_n18497_));
  XNOR2_X1   g18396(.A1(new_n18497_), .A2(new_n18496_), .ZN(new_n18498_));
  NAND2_X1   g18397(.A1(new_n18498_), .A2(new_n18447_), .ZN(new_n18499_));
  OAI22_X1   g18398(.A1(new_n4529_), .A2(new_n14886_), .B1(new_n15114_), .B2(new_n4527_), .ZN(new_n18500_));
  OAI21_X1   g18399(.A1(new_n79_), .A2(new_n15305_), .B(new_n18500_), .ZN(new_n18501_));
  OR2_X2     g18400(.A1(new_n18498_), .A2(new_n18447_), .Z(new_n18502_));
  NAND3_X1   g18401(.A1(new_n18502_), .A2(new_n18499_), .A3(new_n18501_), .ZN(new_n18503_));
  NAND2_X1   g18402(.A1(new_n18503_), .A2(new_n101_), .ZN(new_n18504_));
  XNOR2_X1   g18403(.A1(new_n18504_), .A2(new_n15312_), .ZN(new_n18505_));
  XOR2_X1    g18404(.A1(new_n15511_), .A2(new_n10539_), .Z(new_n18506_));
  NOR2_X1    g18405(.A1(new_n18476_), .A2(new_n18506_), .ZN(new_n18507_));
  XNOR2_X1   g18406(.A1(new_n18507_), .A2(new_n18474_), .ZN(new_n18508_));
  XOR2_X1    g18407(.A1(new_n18508_), .A2(new_n18457_), .Z(new_n18509_));
  XOR2_X1    g18408(.A1(new_n18509_), .A2(new_n18404_), .Z(new_n18510_));
  INV_X1     g18409(.I(new_n18510_), .ZN(new_n18511_));
  XOR2_X1    g18410(.A1(new_n18509_), .A2(new_n18405_), .Z(new_n18512_));
  NOR2_X1    g18411(.A1(new_n18512_), .A2(new_n18505_), .ZN(new_n18513_));
  AOI21_X1   g18412(.A1(new_n18505_), .A2(new_n18511_), .B(new_n18513_), .ZN(new_n18514_));
  NOR2_X1    g18413(.A1(new_n18495_), .A2(new_n18514_), .ZN(new_n18515_));
  INV_X1     g18414(.I(new_n18515_), .ZN(new_n18516_));
  AOI21_X1   g18415(.A1(new_n18395_), .A2(new_n18438_), .B(new_n18516_), .ZN(new_n18517_));
  NOR3_X1    g18416(.A1(new_n18333_), .A2(new_n18267_), .A3(new_n18336_), .ZN(new_n18518_));
  AOI21_X1   g18417(.A1(new_n18207_), .A2(new_n18268_), .B(new_n18329_), .ZN(new_n18519_));
  OAI21_X1   g18418(.A1(new_n18518_), .A2(new_n18519_), .B(new_n18391_), .ZN(new_n18520_));
  NOR3_X1    g18419(.A1(new_n18520_), .A2(new_n18437_), .A3(new_n18515_), .ZN(new_n18521_));
  OAI21_X1   g18420(.A1(new_n18521_), .A2(new_n18517_), .B(new_n18490_), .ZN(new_n18522_));
  INV_X1     g18421(.I(new_n18487_), .ZN(new_n18523_));
  NAND2_X1   g18422(.A1(new_n18523_), .A2(new_n18488_), .ZN(new_n18524_));
  OAI21_X1   g18423(.A1(new_n18520_), .A2(new_n18437_), .B(new_n18515_), .ZN(new_n18525_));
  NAND4_X1   g18424(.A1(\result[27] ), .A2(new_n18391_), .A3(new_n18438_), .A4(new_n18516_), .ZN(new_n18526_));
  NAND3_X1   g18425(.A1(new_n18525_), .A2(new_n18526_), .A3(new_n18524_), .ZN(new_n18527_));
  NAND2_X1   g18426(.A1(new_n18522_), .A2(new_n18527_), .ZN(\result[31] ));
endmodule


