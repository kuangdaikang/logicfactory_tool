// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:35 2022

module ts10  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21,
    \v22.0 , \v22.1 , \v22.2 , \v22.3 , \v22.4 , \v22.5 , \v22.6 , \v22.7 ,
    \v22.8 , \v22.9 , \v22.10 , \v22.11 , \v22.12 , \v22.13 , \v22.14 ,
    \v22.15   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21;
  output \v22.0 , \v22.1 , \v22.2 , \v22.3 , \v22.4 , \v22.5 , \v22.6 ,
    \v22.7 , \v22.8 , \v22.9 , \v22.10 , \v22.11 , \v22.12 , \v22.13 ,
    \v22.14 , \v22.15 ;
  wire new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_, new_n45_,
    new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_,
    new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_,
    new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_,
    new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_,
    new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_,
    new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_,
    new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n113_, new_n114_, new_n115_,
    new_n116_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n129_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n244_, new_n245_, new_n246_, new_n247_;
  assign new_n39_ = ~v18 & v21;
  assign new_n40_ = v10 & new_n39_;
  assign new_n41_ = v18 & ~v21;
  assign new_n42_ = v9 & new_n41_;
  assign new_n43_ = ~new_n40_ & ~new_n42_;
  assign new_n44_ = ~v20 & ~new_n43_;
  assign new_n45_ = v17 & new_n44_;
  assign new_n46_ = v12 & new_n39_;
  assign new_n47_ = v11 & new_n41_;
  assign new_n48_ = ~new_n46_ & ~new_n47_;
  assign new_n49_ = v20 & ~new_n48_;
  assign new_n50_ = ~v17 & new_n49_;
  assign new_n51_ = ~new_n45_ & ~new_n50_;
  assign new_n52_ = ~v19 & ~new_n51_;
  assign new_n53_ = v16 & new_n52_;
  assign new_n54_ = v14 & new_n39_;
  assign new_n55_ = v13 & new_n41_;
  assign new_n56_ = ~new_n54_ & ~new_n55_;
  assign new_n57_ = ~v20 & ~new_n56_;
  assign new_n58_ = v17 & new_n57_;
  assign new_n59_ = v0 & new_n39_;
  assign new_n60_ = v15 & new_n41_;
  assign new_n61_ = ~new_n59_ & ~new_n60_;
  assign new_n62_ = v20 & ~new_n61_;
  assign new_n63_ = ~v17 & new_n62_;
  assign new_n64_ = ~new_n58_ & ~new_n63_;
  assign new_n65_ = v19 & ~new_n64_;
  assign new_n66_ = ~v16 & new_n65_;
  assign \v22.0  = new_n53_ | new_n66_;
  assign new_n68_ = v11 & new_n39_;
  assign new_n69_ = v10 & new_n41_;
  assign new_n70_ = ~new_n68_ & ~new_n69_;
  assign new_n71_ = ~v20 & ~new_n70_;
  assign new_n72_ = v17 & new_n71_;
  assign new_n73_ = v13 & new_n39_;
  assign new_n74_ = v12 & new_n41_;
  assign new_n75_ = ~new_n73_ & ~new_n74_;
  assign new_n76_ = v20 & ~new_n75_;
  assign new_n77_ = ~v17 & new_n76_;
  assign new_n78_ = ~new_n72_ & ~new_n77_;
  assign new_n79_ = ~v19 & ~new_n78_;
  assign new_n80_ = v16 & new_n79_;
  assign new_n81_ = v15 & new_n39_;
  assign new_n82_ = v14 & new_n41_;
  assign new_n83_ = ~new_n81_ & ~new_n82_;
  assign new_n84_ = ~v20 & ~new_n83_;
  assign new_n85_ = v17 & new_n84_;
  assign new_n86_ = v1 & new_n39_;
  assign new_n87_ = v0 & new_n41_;
  assign new_n88_ = ~new_n86_ & ~new_n87_;
  assign new_n89_ = v20 & ~new_n88_;
  assign new_n90_ = ~v17 & new_n89_;
  assign new_n91_ = ~new_n85_ & ~new_n90_;
  assign new_n92_ = v19 & ~new_n91_;
  assign new_n93_ = ~v16 & new_n92_;
  assign \v22.1  = new_n80_ | new_n93_;
  assign new_n95_ = ~v20 & ~new_n48_;
  assign new_n96_ = v17 & new_n95_;
  assign new_n97_ = v20 & ~new_n56_;
  assign new_n98_ = ~v17 & new_n97_;
  assign new_n99_ = ~new_n96_ & ~new_n98_;
  assign new_n100_ = ~v19 & ~new_n99_;
  assign new_n101_ = v16 & new_n100_;
  assign new_n102_ = ~v20 & ~new_n61_;
  assign new_n103_ = v17 & new_n102_;
  assign new_n104_ = v2 & new_n39_;
  assign new_n105_ = v1 & new_n41_;
  assign new_n106_ = ~new_n104_ & ~new_n105_;
  assign new_n107_ = v20 & ~new_n106_;
  assign new_n108_ = ~v17 & new_n107_;
  assign new_n109_ = ~new_n103_ & ~new_n108_;
  assign new_n110_ = v19 & ~new_n109_;
  assign new_n111_ = ~v16 & new_n110_;
  assign \v22.2  = new_n101_ | new_n111_;
  assign new_n113_ = ~v20 & ~new_n75_;
  assign new_n114_ = v17 & new_n113_;
  assign new_n115_ = v20 & ~new_n83_;
  assign new_n116_ = ~v17 & new_n115_;
  assign new_n117_ = ~new_n114_ & ~new_n116_;
  assign new_n118_ = ~v19 & ~new_n117_;
  assign new_n119_ = v16 & new_n118_;
  assign new_n120_ = ~v20 & ~new_n88_;
  assign new_n121_ = v17 & new_n120_;
  assign new_n122_ = v3 & new_n39_;
  assign new_n123_ = v2 & new_n41_;
  assign new_n124_ = ~new_n122_ & ~new_n123_;
  assign new_n125_ = v20 & ~new_n124_;
  assign new_n126_ = ~v17 & new_n125_;
  assign new_n127_ = ~new_n121_ & ~new_n126_;
  assign new_n128_ = v19 & ~new_n127_;
  assign new_n129_ = ~v16 & new_n128_;
  assign \v22.3  = new_n119_ | new_n129_;
  assign new_n131_ = ~v19 & ~new_n64_;
  assign new_n132_ = v16 & new_n131_;
  assign new_n133_ = ~v20 & ~new_n106_;
  assign new_n134_ = v17 & new_n133_;
  assign new_n135_ = v4 & new_n39_;
  assign new_n136_ = v3 & new_n41_;
  assign new_n137_ = ~new_n135_ & ~new_n136_;
  assign new_n138_ = v20 & ~new_n137_;
  assign new_n139_ = ~v17 & new_n138_;
  assign new_n140_ = ~new_n134_ & ~new_n139_;
  assign new_n141_ = v19 & ~new_n140_;
  assign new_n142_ = ~v16 & new_n141_;
  assign \v22.4  = new_n132_ | new_n142_;
  assign new_n144_ = ~v19 & ~new_n91_;
  assign new_n145_ = v16 & new_n144_;
  assign new_n146_ = ~v20 & ~new_n124_;
  assign new_n147_ = v17 & new_n146_;
  assign new_n148_ = v5 & new_n39_;
  assign new_n149_ = v4 & new_n41_;
  assign new_n150_ = ~new_n148_ & ~new_n149_;
  assign new_n151_ = v20 & ~new_n150_;
  assign new_n152_ = ~v17 & new_n151_;
  assign new_n153_ = ~new_n147_ & ~new_n152_;
  assign new_n154_ = v19 & ~new_n153_;
  assign new_n155_ = ~v16 & new_n154_;
  assign \v22.5  = new_n145_ | new_n155_;
  assign new_n157_ = ~v19 & ~new_n109_;
  assign new_n158_ = v16 & new_n157_;
  assign new_n159_ = ~v20 & ~new_n137_;
  assign new_n160_ = v17 & new_n159_;
  assign new_n161_ = v6 & new_n39_;
  assign new_n162_ = v5 & new_n41_;
  assign new_n163_ = ~new_n161_ & ~new_n162_;
  assign new_n164_ = v20 & ~new_n163_;
  assign new_n165_ = ~v17 & new_n164_;
  assign new_n166_ = ~new_n160_ & ~new_n165_;
  assign new_n167_ = v19 & ~new_n166_;
  assign new_n168_ = ~v16 & new_n167_;
  assign \v22.6  = new_n158_ | new_n168_;
  assign new_n170_ = ~v19 & ~new_n127_;
  assign new_n171_ = v16 & new_n170_;
  assign new_n172_ = ~v20 & ~new_n150_;
  assign new_n173_ = v17 & new_n172_;
  assign new_n174_ = v7 & new_n39_;
  assign new_n175_ = v6 & new_n41_;
  assign new_n176_ = ~new_n174_ & ~new_n175_;
  assign new_n177_ = v20 & ~new_n176_;
  assign new_n178_ = ~v17 & new_n177_;
  assign new_n179_ = ~new_n173_ & ~new_n178_;
  assign new_n180_ = v19 & ~new_n179_;
  assign new_n181_ = ~v16 & new_n180_;
  assign \v22.7  = new_n171_ | new_n181_;
  assign new_n183_ = ~v19 & ~new_n140_;
  assign new_n184_ = v16 & new_n183_;
  assign new_n185_ = ~v20 & ~new_n163_;
  assign new_n186_ = v17 & new_n185_;
  assign new_n187_ = v8 & new_n39_;
  assign new_n188_ = v7 & new_n41_;
  assign new_n189_ = ~new_n187_ & ~new_n188_;
  assign new_n190_ = v20 & ~new_n189_;
  assign new_n191_ = ~v17 & new_n190_;
  assign new_n192_ = ~new_n186_ & ~new_n191_;
  assign new_n193_ = v19 & ~new_n192_;
  assign new_n194_ = ~v16 & new_n193_;
  assign \v22.8  = new_n184_ | new_n194_;
  assign new_n196_ = ~v19 & ~new_n153_;
  assign new_n197_ = v16 & new_n196_;
  assign new_n198_ = ~v20 & ~new_n176_;
  assign new_n199_ = v17 & new_n198_;
  assign new_n200_ = v9 & new_n39_;
  assign new_n201_ = v8 & new_n41_;
  assign new_n202_ = ~new_n200_ & ~new_n201_;
  assign new_n203_ = v20 & ~new_n202_;
  assign new_n204_ = ~v17 & new_n203_;
  assign new_n205_ = ~new_n199_ & ~new_n204_;
  assign new_n206_ = v19 & ~new_n205_;
  assign new_n207_ = ~v16 & new_n206_;
  assign \v22.9  = new_n197_ | new_n207_;
  assign new_n209_ = ~v19 & ~new_n166_;
  assign new_n210_ = v16 & new_n209_;
  assign new_n211_ = ~v20 & ~new_n189_;
  assign new_n212_ = v17 & new_n211_;
  assign new_n213_ = v20 & ~new_n43_;
  assign new_n214_ = ~v17 & new_n213_;
  assign new_n215_ = ~new_n212_ & ~new_n214_;
  assign new_n216_ = v19 & ~new_n215_;
  assign new_n217_ = ~v16 & new_n216_;
  assign \v22.10  = new_n210_ | new_n217_;
  assign new_n219_ = ~v19 & ~new_n179_;
  assign new_n220_ = v16 & new_n219_;
  assign new_n221_ = ~v20 & ~new_n202_;
  assign new_n222_ = v17 & new_n221_;
  assign new_n223_ = v20 & ~new_n70_;
  assign new_n224_ = ~v17 & new_n223_;
  assign new_n225_ = ~new_n222_ & ~new_n224_;
  assign new_n226_ = v19 & ~new_n225_;
  assign new_n227_ = ~v16 & new_n226_;
  assign \v22.11  = new_n220_ | new_n227_;
  assign new_n229_ = ~v19 & ~new_n192_;
  assign new_n230_ = v16 & new_n229_;
  assign new_n231_ = v19 & ~new_n51_;
  assign new_n232_ = ~v16 & new_n231_;
  assign \v22.12  = new_n230_ | new_n232_;
  assign new_n234_ = ~v19 & ~new_n205_;
  assign new_n235_ = v16 & new_n234_;
  assign new_n236_ = v19 & ~new_n78_;
  assign new_n237_ = ~v16 & new_n236_;
  assign \v22.13  = new_n235_ | new_n237_;
  assign new_n239_ = ~v19 & ~new_n215_;
  assign new_n240_ = v16 & new_n239_;
  assign new_n241_ = v19 & ~new_n99_;
  assign new_n242_ = ~v16 & new_n241_;
  assign \v22.14  = new_n240_ | new_n242_;
  assign new_n244_ = ~v19 & ~new_n225_;
  assign new_n245_ = v16 & new_n244_;
  assign new_n246_ = v19 & ~new_n117_;
  assign new_n247_ = ~v16 & new_n246_;
  assign \v22.15  = new_n245_ | new_n247_;
endmodule


