// Benchmark "unreg" written by ABC on Fri Feb 25 15:12:35 2022

module unreg ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, s, t, u, v, w, x, y,
    z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0,
    l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, s, t, u, v,
    w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0;
  output l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1;
  wire new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n60_,
    new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n74_, new_n75_, new_n76_,
    new_n77_, new_n78_, new_n79_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n116_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_;
  assign new_n53_ = t & w;
  assign new_n54_ = ~d & ~t;
  assign new_n55_ = ~new_n53_ & ~new_n54_;
  assign new_n56_ = ~s & new_n55_;
  assign new_n57_ = ~u & ~v;
  assign new_n58_ = u & new_n56_;
  assign l0 = new_n57_ | new_n58_;
  assign new_n60_ = t & x;
  assign new_n61_ = ~c & ~t;
  assign new_n62_ = ~new_n60_ & ~new_n61_;
  assign new_n63_ = ~s & new_n62_;
  assign new_n64_ = ~u & ~w;
  assign new_n65_ = u & new_n63_;
  assign m0 = new_n64_ | new_n65_;
  assign new_n67_ = t & y;
  assign new_n68_ = ~b & ~t;
  assign new_n69_ = ~new_n67_ & ~new_n68_;
  assign new_n70_ = ~s & new_n69_;
  assign new_n71_ = ~u & ~x;
  assign new_n72_ = u & new_n70_;
  assign n0 = new_n71_ | new_n72_;
  assign new_n74_ = ~a & ~t;
  assign new_n75_ = ~q & t;
  assign new_n76_ = ~new_n74_ & ~new_n75_;
  assign new_n77_ = ~s & new_n76_;
  assign new_n78_ = ~u & ~y;
  assign new_n79_ = u & new_n77_;
  assign o0 = new_n78_ | new_n79_;
  assign new_n81_ = t & a0;
  assign new_n82_ = ~h & ~t;
  assign new_n83_ = ~new_n81_ & ~new_n82_;
  assign new_n84_ = ~s & new_n83_;
  assign new_n85_ = ~u & ~z;
  assign new_n86_ = u & new_n84_;
  assign p0 = new_n85_ | new_n86_;
  assign new_n88_ = t & b0;
  assign new_n89_ = ~g & ~t;
  assign new_n90_ = ~new_n88_ & ~new_n89_;
  assign new_n91_ = ~s & new_n90_;
  assign new_n92_ = ~u & ~a0;
  assign new_n93_ = u & new_n91_;
  assign q0 = new_n92_ | new_n93_;
  assign new_n95_ = t & c0;
  assign new_n96_ = ~f & ~t;
  assign new_n97_ = ~new_n95_ & ~new_n96_;
  assign new_n98_ = ~s & new_n97_;
  assign new_n99_ = ~u & ~b0;
  assign new_n100_ = u & new_n98_;
  assign r0 = new_n99_ | new_n100_;
  assign new_n102_ = t & v;
  assign new_n103_ = ~e & ~t;
  assign new_n104_ = ~new_n102_ & ~new_n103_;
  assign new_n105_ = ~s & new_n104_;
  assign new_n106_ = ~u & ~c0;
  assign new_n107_ = u & new_n105_;
  assign s0 = new_n106_ | new_n107_;
  assign new_n109_ = t & e0;
  assign new_n110_ = ~l & ~t;
  assign new_n111_ = ~new_n109_ & ~new_n110_;
  assign new_n112_ = ~s & new_n111_;
  assign new_n113_ = ~u & ~d0;
  assign new_n114_ = u & new_n112_;
  assign t0 = new_n113_ | new_n114_;
  assign new_n116_ = t & f0;
  assign new_n117_ = ~k & ~t;
  assign new_n118_ = ~new_n116_ & ~new_n117_;
  assign new_n119_ = ~s & new_n118_;
  assign new_n120_ = ~u & ~e0;
  assign new_n121_ = u & new_n119_;
  assign u0 = new_n120_ | new_n121_;
  assign new_n123_ = t & g0;
  assign new_n124_ = ~j & ~t;
  assign new_n125_ = ~new_n123_ & ~new_n124_;
  assign new_n126_ = ~s & new_n125_;
  assign new_n127_ = ~u & ~f0;
  assign new_n128_ = u & new_n126_;
  assign v0 = new_n127_ | new_n128_;
  assign new_n130_ = t & z;
  assign new_n131_ = ~i & ~t;
  assign new_n132_ = ~new_n130_ & ~new_n131_;
  assign new_n133_ = ~s & new_n132_;
  assign new_n134_ = ~u & ~g0;
  assign new_n135_ = u & new_n133_;
  assign w0 = new_n134_ | new_n135_;
  assign new_n137_ = t & i0;
  assign new_n138_ = ~p & ~t;
  assign new_n139_ = ~new_n137_ & ~new_n138_;
  assign new_n140_ = ~s & new_n139_;
  assign new_n141_ = ~u & ~h0;
  assign new_n142_ = u & new_n140_;
  assign x0 = new_n141_ | new_n142_;
  assign new_n144_ = t & j0;
  assign new_n145_ = ~o & ~t;
  assign new_n146_ = ~new_n144_ & ~new_n145_;
  assign new_n147_ = ~s & new_n146_;
  assign new_n148_ = ~u & ~i0;
  assign new_n149_ = u & new_n147_;
  assign y0 = new_n148_ | new_n149_;
  assign new_n151_ = t & k0;
  assign new_n152_ = ~n & ~t;
  assign new_n153_ = ~new_n151_ & ~new_n152_;
  assign new_n154_ = ~s & new_n153_;
  assign new_n155_ = ~u & ~j0;
  assign new_n156_ = u & new_n154_;
  assign z0 = new_n155_ | new_n156_;
  assign new_n158_ = t & d0;
  assign new_n159_ = ~m & ~t;
  assign new_n160_ = ~new_n158_ & ~new_n159_;
  assign new_n161_ = ~s & new_n160_;
  assign new_n162_ = ~u & ~k0;
  assign new_n163_ = u & new_n161_;
  assign a1 = new_n162_ | new_n163_;
endmodule


