// Benchmark "i2c" written by ABC on Mon Sep 11 23:31:09 2023

module i2c ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n473_, new_n474_, new_n475_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n485_, new_n486_, new_n487_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n510_,
    new_n511_, new_n512_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n521_, new_n522_, new_n523_, new_n525_,
    new_n526_, new_n527_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n553_, new_n554_, new_n555_, new_n557_, new_n558_, new_n559_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n890_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n957_, new_n958_, new_n959_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_, new_n971_,
    new_n972_, new_n973_, new_n975_, new_n976_, new_n977_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n984_, new_n985_, new_n987_,
    new_n988_, new_n990_, new_n991_, new_n993_, new_n994_, new_n996_,
    new_n997_, new_n998_, new_n1000_, new_n1001_, new_n1002_, new_n1004_,
    new_n1005_, new_n1006_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1015_, new_n1016_, new_n1018_, new_n1019_,
    new_n1021_, new_n1022_, new_n1024_, new_n1025_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1043_, new_n1044_, new_n1046_, new_n1047_, new_n1048_,
    new_n1050_, new_n1051_, new_n1053_, new_n1054_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1062_, new_n1063_, new_n1065_,
    new_n1066_, new_n1068_, new_n1069_, new_n1071_, new_n1072_, new_n1074_,
    new_n1075_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1090_, new_n1092_, new_n1094_, new_n1095_, new_n1097_, new_n1098_,
    new_n1100_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1156_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1184_, new_n1185_, new_n1187_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1195_,
    new_n1196_, new_n1198_, new_n1199_, new_n1201_, new_n1202_, new_n1204_,
    new_n1207_, new_n1208_, new_n1211_, new_n1217_, new_n1219_;
  NOR2_X1    g000(.A1(pi005), .A2(pi022), .ZN(new_n291_));
  NOR2_X1    g001(.A1(pi009), .A2(pi011), .ZN(new_n292_));
  NOR2_X1    g002(.A1(pi013), .A2(pi014), .ZN(new_n293_));
  INV_X1     g003(.I(pi008), .ZN(new_n294_));
  INV_X1     g004(.I(pi017), .ZN(new_n295_));
  INV_X1     g005(.I(pi021), .ZN(new_n296_));
  NAND3_X1   g006(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1     g007(.I(pi006), .ZN(new_n298_));
  INV_X1     g008(.I(pi007), .ZN(new_n299_));
  INV_X1     g009(.I(pi012), .ZN(new_n300_));
  NOR4_X1    g010(.A1(pi004), .A2(pi016), .A3(pi018), .A4(pi019), .ZN(new_n301_));
  NAND4_X1   g011(.A1(new_n301_), .A2(new_n298_), .A3(new_n299_), .A4(new_n300_), .ZN(new_n302_));
  NOR2_X1    g012(.A1(new_n302_), .A2(new_n297_), .ZN(new_n303_));
  NAND4_X1   g013(.A1(new_n303_), .A2(new_n291_), .A3(new_n292_), .A4(new_n293_), .ZN(new_n304_));
  AOI21_X1   g014(.A1(new_n304_), .A2(pi054), .B(pi000), .ZN(new_n305_));
  INV_X1     g015(.I(pi054), .ZN(new_n306_));
  NOR2_X1    g016(.A1(new_n292_), .A2(pi056), .ZN(new_n307_));
  NAND2_X1   g017(.A1(new_n307_), .A2(new_n291_), .ZN(new_n308_));
  NOR2_X1    g018(.A1(pi008), .A2(pi021), .ZN(new_n309_));
  NAND4_X1   g019(.A1(new_n293_), .A2(new_n309_), .A3(new_n299_), .A4(pi010), .ZN(new_n310_));
  INV_X1     g020(.I(pi010), .ZN(new_n311_));
  NAND3_X1   g021(.A1(new_n309_), .A2(new_n299_), .A3(pi013), .ZN(new_n312_));
  OR3_X2     g022(.A1(pi007), .A2(pi008), .A3(pi021), .Z(new_n313_));
  OAI21_X1   g023(.A1(pi008), .A2(pi021), .B(pi007), .ZN(new_n314_));
  AOI21_X1   g024(.A1(pi008), .A2(pi021), .B(pi013), .ZN(new_n315_));
  NAND3_X1   g025(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1   g026(.A1(new_n316_), .A2(new_n312_), .B(pi014), .ZN(new_n317_));
  INV_X1     g027(.I(pi014), .ZN(new_n318_));
  NOR3_X1    g028(.A1(new_n313_), .A2(pi013), .A3(new_n318_), .ZN(new_n319_));
  OAI21_X1   g029(.A1(new_n317_), .A2(new_n319_), .B(new_n311_), .ZN(new_n320_));
  NOR2_X1    g030(.A1(pi006), .A2(pi012), .ZN(new_n321_));
  NAND4_X1   g031(.A1(new_n301_), .A2(new_n295_), .A3(new_n291_), .A4(new_n321_), .ZN(new_n322_));
  AOI21_X1   g032(.A1(new_n320_), .A2(new_n310_), .B(new_n322_), .ZN(new_n323_));
  NOR2_X1    g033(.A1(new_n291_), .A2(pi056), .ZN(new_n324_));
  OAI21_X1   g034(.A1(new_n323_), .A2(new_n324_), .B(new_n292_), .ZN(new_n325_));
  AOI21_X1   g035(.A1(new_n325_), .A2(new_n308_), .B(new_n306_), .ZN(new_n326_));
  NOR2_X1    g036(.A1(pi003), .A2(pi129), .ZN(new_n327_));
  OAI21_X1   g037(.A1(new_n326_), .A2(new_n305_), .B(new_n327_), .ZN(po015));
  INV_X1     g038(.I(pi009), .ZN(new_n329_));
  INV_X1     g039(.I(new_n321_), .ZN(new_n330_));
  NOR2_X1    g040(.A1(new_n330_), .A2(pi005), .ZN(new_n331_));
  INV_X1     g041(.I(new_n331_), .ZN(new_n332_));
  NAND2_X1   g042(.A1(new_n330_), .A2(pi005), .ZN(new_n333_));
  NAND2_X1   g043(.A1(pi006), .A2(pi012), .ZN(new_n334_));
  NAND4_X1   g044(.A1(new_n332_), .A2(new_n299_), .A3(new_n333_), .A4(new_n334_), .ZN(new_n335_));
  NAND2_X1   g045(.A1(new_n331_), .A2(pi007), .ZN(new_n336_));
  AOI21_X1   g046(.A1(new_n335_), .A2(new_n336_), .B(pi013), .ZN(new_n337_));
  INV_X1     g047(.I(pi013), .ZN(new_n338_));
  NOR3_X1    g048(.A1(new_n332_), .A2(pi007), .A3(new_n338_), .ZN(new_n339_));
  OAI21_X1   g049(.A1(new_n337_), .A2(new_n339_), .B(new_n329_), .ZN(new_n340_));
  NOR2_X1    g050(.A1(pi007), .A2(pi013), .ZN(new_n341_));
  INV_X1     g051(.I(new_n341_), .ZN(new_n342_));
  NOR2_X1    g052(.A1(new_n332_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1   g053(.A1(new_n343_), .A2(pi009), .ZN(new_n344_));
  NOR2_X1    g054(.A1(pi010), .A2(pi022), .ZN(new_n345_));
  INV_X1     g055(.I(new_n345_), .ZN(new_n346_));
  NOR3_X1    g056(.A1(new_n346_), .A2(pi014), .A3(new_n306_), .ZN(new_n347_));
  INV_X1     g057(.I(pi011), .ZN(new_n348_));
  NAND2_X1   g058(.A1(new_n294_), .A2(new_n348_), .ZN(new_n349_));
  NOR3_X1    g059(.A1(new_n349_), .A2(pi017), .A3(pi021), .ZN(new_n350_));
  NAND3_X1   g060(.A1(new_n347_), .A2(new_n350_), .A3(new_n301_), .ZN(new_n351_));
  AOI21_X1   g061(.A1(new_n340_), .A2(new_n344_), .B(new_n351_), .ZN(new_n352_));
  NOR3_X1    g062(.A1(pi008), .A2(pi014), .A3(pi021), .ZN(new_n353_));
  NOR2_X1    g063(.A1(pi011), .A2(pi012), .ZN(new_n354_));
  INV_X1     g064(.I(new_n354_), .ZN(new_n355_));
  NOR2_X1    g065(.A1(new_n346_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1     g066(.I(pi005), .ZN(new_n357_));
  NAND2_X1   g067(.A1(new_n357_), .A2(new_n298_), .ZN(new_n358_));
  NOR2_X1    g068(.A1(new_n342_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1   g069(.A1(new_n356_), .A2(new_n359_), .A3(new_n301_), .A4(new_n353_), .ZN(new_n360_));
  NOR2_X1    g070(.A1(new_n306_), .A2(pi017), .ZN(new_n361_));
  AOI21_X1   g071(.A1(new_n360_), .A2(new_n361_), .B(pi001), .ZN(new_n362_));
  OAI21_X1   g072(.A1(new_n352_), .A2(new_n362_), .B(new_n327_), .ZN(po016));
  INV_X1     g073(.I(pi082), .ZN(new_n364_));
  INV_X1     g074(.I(pi002), .ZN(new_n365_));
  NOR2_X1    g075(.A1(pi043), .A2(pi047), .ZN(new_n366_));
  NOR2_X1    g076(.A1(pi045), .A2(pi048), .ZN(new_n367_));
  NAND3_X1   g077(.A1(new_n366_), .A2(new_n367_), .A3(new_n365_), .ZN(new_n368_));
  NOR2_X1    g078(.A1(pi041), .A2(pi046), .ZN(new_n369_));
  NOR2_X1    g079(.A1(pi038), .A2(pi050), .ZN(new_n370_));
  NAND2_X1   g080(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1    g081(.A1(pi042), .A2(pi044), .ZN(new_n372_));
  INV_X1     g082(.I(new_n372_), .ZN(new_n373_));
  NOR2_X1    g083(.A1(new_n373_), .A2(pi040), .ZN(new_n374_));
  INV_X1     g084(.I(new_n374_), .ZN(new_n375_));
  NOR2_X1    g085(.A1(pi024), .A2(pi049), .ZN(new_n376_));
  INV_X1     g086(.I(new_n376_), .ZN(new_n377_));
  NOR2_X1    g087(.A1(pi015), .A2(pi020), .ZN(new_n378_));
  INV_X1     g088(.I(new_n378_), .ZN(new_n379_));
  NOR2_X1    g089(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1     g090(.I(new_n380_), .ZN(new_n381_));
  NOR4_X1    g091(.A1(new_n381_), .A2(new_n375_), .A3(new_n368_), .A4(new_n371_), .ZN(new_n382_));
  NAND2_X1   g092(.A1(pi122), .A2(pi127), .ZN(new_n383_));
  INV_X1     g093(.I(new_n383_), .ZN(new_n384_));
  NOR2_X1    g094(.A1(new_n384_), .A2(pi065), .ZN(new_n385_));
  OAI21_X1   g095(.A1(new_n382_), .A2(new_n364_), .B(new_n385_), .ZN(new_n386_));
  NOR2_X1    g096(.A1(new_n383_), .A2(pi082), .ZN(new_n387_));
  NOR2_X1    g097(.A1(pi038), .A2(pi040), .ZN(new_n388_));
  NOR3_X1    g098(.A1(pi041), .A2(pi046), .A3(pi050), .ZN(new_n389_));
  NAND3_X1   g099(.A1(new_n389_), .A2(new_n372_), .A3(new_n388_), .ZN(new_n390_));
  NOR2_X1    g100(.A1(new_n390_), .A2(pi043), .ZN(new_n391_));
  INV_X1     g101(.I(new_n391_), .ZN(new_n392_));
  NOR2_X1    g102(.A1(new_n379_), .A2(pi049), .ZN(new_n393_));
  INV_X1     g103(.I(new_n393_), .ZN(new_n394_));
  NOR2_X1    g104(.A1(pi047), .A2(pi048), .ZN(new_n395_));
  INV_X1     g105(.I(new_n395_), .ZN(new_n396_));
  NOR2_X1    g106(.A1(pi024), .A2(pi045), .ZN(new_n397_));
  INV_X1     g107(.I(new_n397_), .ZN(new_n398_));
  NOR4_X1    g108(.A1(new_n392_), .A2(new_n394_), .A3(new_n396_), .A4(new_n398_), .ZN(new_n399_));
  NOR2_X1    g109(.A1(new_n399_), .A2(new_n364_), .ZN(new_n400_));
  OAI21_X1   g110(.A1(new_n400_), .A2(new_n387_), .B(pi002), .ZN(new_n401_));
  AOI21_X1   g111(.A1(new_n401_), .A2(new_n386_), .B(pi129), .ZN(po017));
  INV_X1     g112(.I(pi113), .ZN(new_n403_));
  INV_X1     g113(.I(pi123), .ZN(new_n404_));
  NAND3_X1   g114(.A1(new_n403_), .A2(new_n404_), .A3(pi000), .ZN(new_n405_));
  NOR3_X1    g115(.A1(new_n346_), .A2(pi009), .A3(pi014), .ZN(new_n406_));
  NAND2_X1   g116(.A1(new_n406_), .A2(new_n359_), .ZN(new_n407_));
  NOR2_X1    g117(.A1(pi008), .A2(pi017), .ZN(new_n408_));
  NAND4_X1   g118(.A1(new_n301_), .A2(new_n296_), .A3(new_n354_), .A4(new_n408_), .ZN(new_n409_));
  NOR2_X1    g119(.A1(pi061), .A2(pi118), .ZN(new_n410_));
  OAI21_X1   g120(.A1(new_n407_), .A2(new_n409_), .B(new_n410_), .ZN(new_n411_));
  AOI21_X1   g121(.A1(new_n411_), .A2(new_n405_), .B(pi129), .ZN(po018));
  INV_X1     g122(.I(new_n327_), .ZN(new_n413_));
  AND3_X2    g123(.A1(new_n350_), .A2(pi054), .A3(new_n301_), .Z(new_n414_));
  NOR4_X1    g124(.A1(new_n311_), .A2(pi009), .A3(pi014), .A4(pi022), .ZN(new_n415_));
  NAND3_X1   g125(.A1(new_n414_), .A2(new_n343_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1   g126(.A1(new_n306_), .A2(pi004), .ZN(new_n417_));
  AOI21_X1   g127(.A1(new_n416_), .A2(new_n417_), .B(new_n413_), .ZN(po019));
  INV_X1     g128(.I(pi059), .ZN(new_n419_));
  NAND2_X1   g129(.A1(new_n406_), .A2(new_n338_), .ZN(new_n420_));
  INV_X1     g130(.I(new_n420_), .ZN(new_n421_));
  AND3_X2    g131(.A1(new_n421_), .A2(new_n419_), .A3(new_n350_), .Z(new_n422_));
  INV_X1     g132(.I(pi016), .ZN(new_n423_));
  NAND2_X1   g133(.A1(new_n423_), .A2(pi054), .ZN(new_n424_));
  NAND2_X1   g134(.A1(new_n357_), .A2(new_n299_), .ZN(new_n425_));
  NOR3_X1    g135(.A1(new_n330_), .A2(new_n425_), .A3(new_n424_), .ZN(new_n426_));
  INV_X1     g136(.I(pi028), .ZN(new_n427_));
  INV_X1     g137(.I(pi018), .ZN(new_n428_));
  NOR2_X1    g138(.A1(pi004), .A2(pi019), .ZN(new_n429_));
  NAND2_X1   g139(.A1(new_n429_), .A2(new_n428_), .ZN(new_n430_));
  NOR4_X1    g140(.A1(new_n430_), .A2(pi025), .A3(new_n427_), .A4(pi029), .ZN(new_n431_));
  NAND3_X1   g141(.A1(new_n422_), .A2(new_n426_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1   g142(.A1(new_n306_), .A2(pi005), .ZN(new_n433_));
  AOI21_X1   g143(.A1(new_n432_), .A2(new_n433_), .B(new_n413_), .ZN(po020));
  INV_X1     g144(.I(pi025), .ZN(new_n435_));
  NOR4_X1    g145(.A1(new_n430_), .A2(new_n435_), .A3(pi028), .A4(pi029), .ZN(new_n436_));
  NAND3_X1   g146(.A1(new_n422_), .A2(new_n426_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1   g147(.A1(new_n306_), .A2(pi006), .ZN(new_n438_));
  AOI21_X1   g148(.A1(new_n437_), .A2(new_n438_), .B(new_n413_), .ZN(po021));
  NAND2_X1   g149(.A1(new_n295_), .A2(pi008), .ZN(new_n440_));
  NOR4_X1    g150(.A1(new_n425_), .A2(new_n440_), .A3(pi018), .A4(pi021), .ZN(new_n441_));
  INV_X1     g151(.I(new_n429_), .ZN(new_n442_));
  NOR2_X1    g152(.A1(new_n442_), .A2(new_n424_), .ZN(new_n443_));
  NOR2_X1    g153(.A1(new_n355_), .A2(pi006), .ZN(new_n444_));
  NAND4_X1   g154(.A1(new_n421_), .A2(new_n441_), .A3(new_n443_), .A4(new_n444_), .ZN(new_n445_));
  NAND2_X1   g155(.A1(new_n306_), .A2(pi007), .ZN(new_n446_));
  AOI21_X1   g156(.A1(new_n445_), .A2(new_n446_), .B(new_n413_), .ZN(po022));
  AND2_X2    g157(.A1(new_n406_), .A2(new_n343_), .Z(new_n448_));
  NAND2_X1   g158(.A1(new_n295_), .A2(new_n428_), .ZN(new_n449_));
  NOR3_X1    g159(.A1(new_n349_), .A2(new_n449_), .A3(new_n296_), .ZN(new_n450_));
  NAND3_X1   g160(.A1(new_n448_), .A2(new_n443_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1   g161(.A1(new_n306_), .A2(pi008), .ZN(new_n452_));
  AOI21_X1   g162(.A1(new_n451_), .A2(new_n452_), .B(new_n413_), .ZN(po023));
  NOR2_X1    g163(.A1(new_n330_), .A2(new_n425_), .ZN(new_n454_));
  INV_X1     g164(.I(new_n293_), .ZN(new_n455_));
  NOR4_X1    g165(.A1(new_n455_), .A2(new_n346_), .A3(pi009), .A4(new_n348_), .ZN(new_n456_));
  NAND3_X1   g166(.A1(new_n408_), .A2(new_n428_), .A3(new_n296_), .ZN(new_n457_));
  INV_X1     g167(.I(new_n457_), .ZN(new_n458_));
  NAND4_X1   g168(.A1(new_n456_), .A2(new_n454_), .A3(new_n458_), .A4(new_n443_), .ZN(new_n459_));
  NAND2_X1   g169(.A1(new_n306_), .A2(pi009), .ZN(new_n460_));
  AOI21_X1   g170(.A1(new_n459_), .A2(new_n460_), .B(new_n413_), .ZN(po024));
  NOR4_X1    g171(.A1(new_n457_), .A2(pi009), .A3(pi010), .A4(pi022), .ZN(new_n462_));
  NOR3_X1    g172(.A1(new_n355_), .A2(new_n425_), .A3(pi006), .ZN(new_n463_));
  NOR4_X1    g173(.A1(new_n442_), .A2(new_n424_), .A3(pi013), .A4(new_n318_), .ZN(new_n464_));
  NAND3_X1   g174(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1   g175(.A1(new_n306_), .A2(pi010), .ZN(new_n466_));
  AOI21_X1   g176(.A1(new_n465_), .A2(new_n466_), .B(new_n413_), .ZN(po025));
  NOR4_X1    g177(.A1(new_n442_), .A2(new_n424_), .A3(pi009), .A4(pi014), .ZN(new_n468_));
  AND3_X2    g178(.A1(new_n311_), .A2(new_n348_), .A3(pi022), .Z(new_n469_));
  NAND4_X1   g179(.A1(new_n343_), .A2(new_n458_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  NAND2_X1   g180(.A1(new_n306_), .A2(pi011), .ZN(new_n471_));
  AOI21_X1   g181(.A1(new_n470_), .A2(new_n471_), .B(new_n413_), .ZN(po026));
  NOR3_X1    g182(.A1(new_n297_), .A2(new_n355_), .A3(new_n428_), .ZN(new_n473_));
  NAND4_X1   g183(.A1(new_n473_), .A2(new_n406_), .A3(new_n359_), .A4(new_n443_), .ZN(new_n474_));
  NAND2_X1   g184(.A1(new_n306_), .A2(pi012), .ZN(new_n475_));
  AOI21_X1   g185(.A1(new_n474_), .A2(new_n475_), .B(new_n413_), .ZN(po027));
  INV_X1     g186(.I(new_n430_), .ZN(new_n477_));
  INV_X1     g187(.I(pi029), .ZN(new_n478_));
  NOR3_X1    g188(.A1(new_n478_), .A2(pi025), .A3(pi028), .ZN(new_n479_));
  AND3_X2    g189(.A1(new_n406_), .A2(new_n477_), .A3(new_n479_), .Z(new_n480_));
  NOR3_X1    g190(.A1(new_n332_), .A2(new_n342_), .A3(new_n424_), .ZN(new_n481_));
  NAND4_X1   g191(.A1(new_n480_), .A2(new_n481_), .A3(new_n419_), .A4(new_n350_), .ZN(new_n482_));
  NAND2_X1   g192(.A1(new_n306_), .A2(pi013), .ZN(new_n483_));
  AOI21_X1   g193(.A1(new_n482_), .A2(new_n483_), .B(new_n413_), .ZN(po028));
  NOR4_X1    g194(.A1(new_n442_), .A2(pi009), .A3(new_n338_), .A4(pi016), .ZN(new_n485_));
  NAND4_X1   g195(.A1(new_n485_), .A2(new_n463_), .A3(new_n347_), .A4(new_n458_), .ZN(new_n486_));
  NAND2_X1   g196(.A1(new_n306_), .A2(pi014), .ZN(new_n487_));
  AOI21_X1   g197(.A1(new_n486_), .A2(new_n487_), .B(new_n413_), .ZN(po029));
  INV_X1     g198(.I(pi015), .ZN(new_n489_));
  INV_X1     g199(.I(pi020), .ZN(new_n490_));
  NAND2_X1   g200(.A1(new_n365_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1   g201(.A1(new_n491_), .A2(new_n489_), .A3(new_n376_), .ZN(new_n492_));
  NOR4_X1    g202(.A1(new_n392_), .A2(pi045), .A3(new_n396_), .A4(new_n492_), .ZN(new_n493_));
  INV_X1     g203(.I(new_n366_), .ZN(new_n494_));
  NOR2_X1    g204(.A1(new_n494_), .A2(pi048), .ZN(new_n495_));
  INV_X1     g205(.I(new_n495_), .ZN(new_n496_));
  NOR4_X1    g206(.A1(new_n496_), .A2(pi045), .A3(new_n377_), .A4(new_n390_), .ZN(new_n497_));
  NOR2_X1    g207(.A1(new_n497_), .A2(new_n489_), .ZN(new_n498_));
  OAI21_X1   g208(.A1(new_n498_), .A2(new_n493_), .B(pi082), .ZN(new_n499_));
  INV_X1     g209(.I(new_n370_), .ZN(new_n500_));
  NOR2_X1    g210(.A1(new_n500_), .A2(pi046), .ZN(new_n501_));
  NAND2_X1   g211(.A1(new_n374_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1    g212(.A1(new_n377_), .A2(pi045), .ZN(new_n503_));
  NOR2_X1    g213(.A1(pi041), .A2(pi043), .ZN(new_n504_));
  NAND4_X1   g214(.A1(new_n503_), .A2(new_n489_), .A3(new_n395_), .A4(new_n504_), .ZN(new_n505_));
  OAI21_X1   g215(.A1(new_n505_), .A2(new_n502_), .B(pi082), .ZN(new_n506_));
  NOR2_X1    g216(.A1(new_n384_), .A2(pi070), .ZN(new_n507_));
  AOI22_X1   g217(.A1(new_n506_), .A2(new_n507_), .B1(pi015), .B2(new_n387_), .ZN(new_n508_));
  AOI21_X1   g218(.A1(new_n499_), .A2(new_n508_), .B(pi129), .ZN(po030));
  NOR4_X1    g219(.A1(new_n342_), .A2(pi005), .A3(new_n298_), .A4(pi012), .ZN(new_n510_));
  NAND3_X1   g220(.A1(new_n414_), .A2(new_n406_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1   g221(.A1(new_n306_), .A2(pi016), .ZN(new_n512_));
  AOI21_X1   g222(.A1(new_n511_), .A2(new_n512_), .B(new_n413_), .ZN(po031));
  NOR4_X1    g223(.A1(new_n430_), .A2(pi028), .A3(pi029), .A4(new_n419_), .ZN(new_n514_));
  INV_X1     g224(.I(new_n361_), .ZN(new_n515_));
  NAND4_X1   g225(.A1(new_n299_), .A2(new_n300_), .A3(new_n423_), .A4(new_n435_), .ZN(new_n516_));
  NOR4_X1    g226(.A1(new_n420_), .A2(new_n358_), .A3(new_n515_), .A4(new_n516_), .ZN(new_n517_));
  NAND4_X1   g227(.A1(new_n517_), .A2(new_n348_), .A3(new_n309_), .A4(new_n514_), .ZN(new_n518_));
  NAND2_X1   g228(.A1(new_n306_), .A2(pi017), .ZN(new_n519_));
  AOI21_X1   g229(.A1(new_n518_), .A2(new_n519_), .B(new_n413_), .ZN(po032));
  NOR2_X1    g230(.A1(new_n423_), .A2(new_n306_), .ZN(new_n521_));
  NAND4_X1   g231(.A1(new_n448_), .A2(new_n350_), .A3(new_n477_), .A4(new_n521_), .ZN(new_n522_));
  NAND2_X1   g232(.A1(new_n306_), .A2(pi018), .ZN(new_n523_));
  AOI21_X1   g233(.A1(new_n522_), .A2(new_n523_), .B(new_n413_), .ZN(po033));
  NOR4_X1    g234(.A1(new_n442_), .A2(new_n424_), .A3(new_n295_), .A4(pi018), .ZN(new_n525_));
  NAND4_X1   g235(.A1(new_n448_), .A2(new_n348_), .A3(new_n309_), .A4(new_n525_), .ZN(new_n526_));
  NAND2_X1   g236(.A1(new_n306_), .A2(pi019), .ZN(new_n527_));
  AOI21_X1   g237(.A1(new_n526_), .A2(new_n527_), .B(new_n413_), .ZN(po034));
  INV_X1     g238(.I(new_n367_), .ZN(new_n529_));
  NAND2_X1   g239(.A1(new_n366_), .A2(new_n369_), .ZN(new_n530_));
  NOR3_X1    g240(.A1(new_n530_), .A2(pi024), .A3(new_n529_), .ZN(new_n531_));
  INV_X1     g241(.I(pi050), .ZN(new_n532_));
  NAND2_X1   g242(.A1(new_n388_), .A2(new_n532_), .ZN(new_n533_));
  NOR4_X1    g243(.A1(new_n533_), .A2(new_n373_), .A3(pi015), .A4(pi049), .ZN(new_n534_));
  AOI21_X1   g244(.A1(new_n534_), .A2(new_n531_), .B(new_n490_), .ZN(new_n535_));
  INV_X1     g245(.I(pi044), .ZN(new_n536_));
  INV_X1     g246(.I(pi040), .ZN(new_n537_));
  INV_X1     g247(.I(pi042), .ZN(new_n538_));
  NAND2_X1   g248(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1    g249(.A1(new_n500_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1   g250(.A1(new_n531_), .A2(new_n536_), .A3(new_n393_), .A4(new_n540_), .ZN(new_n541_));
  NOR2_X1    g251(.A1(new_n541_), .A2(new_n365_), .ZN(new_n542_));
  OAI21_X1   g252(.A1(new_n542_), .A2(new_n535_), .B(pi082), .ZN(new_n543_));
  NAND2_X1   g253(.A1(new_n541_), .A2(pi082), .ZN(new_n544_));
  NOR2_X1    g254(.A1(new_n384_), .A2(pi071), .ZN(new_n545_));
  AOI22_X1   g255(.A1(new_n544_), .A2(new_n545_), .B1(pi020), .B2(new_n387_), .ZN(new_n546_));
  AOI21_X1   g256(.A1(new_n546_), .A2(new_n543_), .B(pi129), .ZN(po035));
  AND3_X2    g257(.A1(new_n296_), .A2(pi019), .A3(pi054), .Z(new_n548_));
  NOR4_X1    g258(.A1(new_n349_), .A2(new_n449_), .A3(pi004), .A4(pi016), .ZN(new_n549_));
  NAND3_X1   g259(.A1(new_n448_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1   g260(.A1(new_n306_), .A2(pi021), .ZN(new_n551_));
  AOI21_X1   g261(.A1(new_n550_), .A2(new_n551_), .B(new_n413_), .ZN(po036));
  NOR3_X1    g262(.A1(new_n455_), .A2(new_n357_), .A3(pi007), .ZN(new_n553_));
  NAND4_X1   g263(.A1(new_n462_), .A2(new_n443_), .A3(new_n444_), .A4(new_n553_), .ZN(new_n554_));
  NAND2_X1   g264(.A1(new_n306_), .A2(pi022), .ZN(new_n555_));
  AOI21_X1   g265(.A1(new_n554_), .A2(new_n555_), .B(new_n413_), .ZN(po037));
  INV_X1     g266(.I(pi023), .ZN(new_n557_));
  INV_X1     g267(.I(pi129), .ZN(new_n558_));
  NAND2_X1   g268(.A1(new_n558_), .A2(pi061), .ZN(new_n559_));
  AOI21_X1   g269(.A1(new_n557_), .A2(pi055), .B(new_n559_), .ZN(po038));
  INV_X1     g270(.I(new_n504_), .ZN(new_n561_));
  NOR2_X1    g271(.A1(new_n561_), .A2(pi047), .ZN(new_n562_));
  NAND2_X1   g272(.A1(new_n562_), .A2(new_n367_), .ZN(new_n563_));
  OAI21_X1   g273(.A1(new_n502_), .A2(new_n563_), .B(pi082), .ZN(new_n564_));
  INV_X1     g274(.I(pi049), .ZN(new_n565_));
  NAND4_X1   g275(.A1(new_n365_), .A2(new_n489_), .A3(new_n490_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1   g276(.A1(new_n566_), .A2(pi082), .ZN(new_n567_));
  NAND2_X1   g277(.A1(new_n567_), .A2(new_n384_), .ZN(new_n568_));
  AOI21_X1   g278(.A1(new_n564_), .A2(new_n568_), .B(pi024), .ZN(new_n569_));
  INV_X1     g279(.I(pi045), .ZN(new_n570_));
  NAND2_X1   g280(.A1(new_n365_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1     g281(.I(new_n571_), .ZN(new_n572_));
  NAND4_X1   g282(.A1(new_n391_), .A2(new_n393_), .A3(new_n395_), .A4(new_n572_), .ZN(new_n573_));
  NAND2_X1   g283(.A1(new_n383_), .A2(pi063), .ZN(new_n574_));
  AOI21_X1   g284(.A1(new_n573_), .A2(pi082), .B(new_n574_), .ZN(new_n575_));
  NOR3_X1    g285(.A1(pi041), .A2(pi043), .A3(pi046), .ZN(new_n576_));
  NAND3_X1   g286(.A1(new_n576_), .A2(new_n395_), .A3(new_n570_), .ZN(new_n577_));
  NAND2_X1   g287(.A1(pi024), .A2(pi082), .ZN(new_n578_));
  NOR4_X1    g288(.A1(new_n577_), .A2(new_n373_), .A3(new_n533_), .A4(new_n578_), .ZN(new_n579_));
  NOR4_X1    g289(.A1(new_n569_), .A2(pi129), .A3(new_n575_), .A4(new_n579_), .ZN(po039));
  INV_X1     g290(.I(pi026), .ZN(new_n581_));
  NOR2_X1    g291(.A1(new_n435_), .A2(pi116), .ZN(new_n582_));
  INV_X1     g292(.I(pi058), .ZN(new_n583_));
  NOR2_X1    g293(.A1(new_n583_), .A2(pi053), .ZN(new_n584_));
  NOR2_X1    g294(.A1(pi027), .A2(pi085), .ZN(new_n585_));
  NAND4_X1   g295(.A1(new_n582_), .A2(new_n584_), .A3(new_n581_), .A4(new_n585_), .ZN(new_n586_));
  INV_X1     g296(.I(new_n582_), .ZN(new_n587_));
  INV_X1     g297(.I(pi085), .ZN(new_n588_));
  NAND2_X1   g298(.A1(new_n588_), .A2(pi053), .ZN(new_n589_));
  NOR4_X1    g299(.A1(new_n587_), .A2(new_n589_), .A3(pi026), .A4(pi027), .ZN(new_n590_));
  INV_X1     g300(.I(pi027), .ZN(new_n591_));
  NOR3_X1    g301(.A1(pi039), .A2(pi051), .A3(pi052), .ZN(new_n592_));
  INV_X1     g302(.I(new_n592_), .ZN(new_n593_));
  INV_X1     g303(.I(pi116), .ZN(new_n594_));
  NOR2_X1    g304(.A1(new_n581_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1     g305(.I(pi110), .ZN(new_n596_));
  OR3_X2     g306(.A1(pi095), .A2(pi097), .A3(pi100), .Z(new_n597_));
  AOI21_X1   g307(.A1(new_n597_), .A2(new_n596_), .B(new_n435_), .ZN(new_n598_));
  OAI21_X1   g308(.A1(new_n598_), .A2(new_n595_), .B(new_n593_), .ZN(new_n599_));
  NAND2_X1   g309(.A1(new_n582_), .A2(pi026), .ZN(new_n600_));
  AOI21_X1   g310(.A1(new_n599_), .A2(new_n600_), .B(pi085), .ZN(new_n601_));
  NOR3_X1    g311(.A1(pi085), .A2(pi096), .A3(pi110), .ZN(new_n602_));
  NOR2_X1    g312(.A1(new_n588_), .A2(new_n594_), .ZN(new_n603_));
  OAI21_X1   g313(.A1(new_n603_), .A2(new_n602_), .B(pi100), .ZN(new_n604_));
  NAND2_X1   g314(.A1(new_n582_), .A2(pi085), .ZN(new_n605_));
  AOI21_X1   g315(.A1(new_n604_), .A2(new_n605_), .B(pi026), .ZN(new_n606_));
  OAI21_X1   g316(.A1(new_n601_), .A2(new_n606_), .B(new_n591_), .ZN(new_n607_));
  NOR3_X1    g317(.A1(pi039), .A2(pi051), .A3(pi052), .ZN(new_n608_));
  NAND2_X1   g318(.A1(new_n608_), .A2(pi116), .ZN(new_n609_));
  AOI21_X1   g319(.A1(new_n587_), .A2(new_n609_), .B(new_n591_), .ZN(new_n610_));
  AND2_X2    g320(.A1(new_n598_), .A2(new_n592_), .Z(new_n611_));
  NOR2_X1    g321(.A1(pi026), .A2(pi085), .ZN(new_n612_));
  OAI21_X1   g322(.A1(new_n611_), .A2(new_n610_), .B(new_n612_), .ZN(new_n613_));
  AOI21_X1   g323(.A1(new_n607_), .A2(new_n613_), .B(pi053), .ZN(new_n614_));
  OAI21_X1   g324(.A1(new_n614_), .A2(new_n590_), .B(new_n583_), .ZN(new_n615_));
  AOI21_X1   g325(.A1(new_n615_), .A2(new_n586_), .B(new_n413_), .ZN(po040));
  INV_X1     g326(.I(new_n603_), .ZN(new_n617_));
  NAND2_X1   g327(.A1(new_n594_), .A2(pi085), .ZN(new_n618_));
  NAND2_X1   g328(.A1(new_n618_), .A2(new_n596_), .ZN(new_n619_));
  INV_X1     g329(.I(pi096), .ZN(new_n620_));
  OAI21_X1   g330(.A1(new_n581_), .A2(new_n594_), .B(new_n620_), .ZN(new_n621_));
  OAI22_X1   g331(.A1(pi026), .A2(new_n617_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1   g332(.A1(new_n622_), .A2(pi100), .ZN(new_n623_));
  NAND3_X1   g333(.A1(new_n609_), .A2(pi026), .A3(new_n588_), .ZN(new_n624_));
  NOR3_X1    g334(.A1(pi027), .A2(pi053), .A3(pi058), .ZN(new_n625_));
  NAND2_X1   g335(.A1(new_n625_), .A2(new_n327_), .ZN(new_n626_));
  AOI21_X1   g336(.A1(new_n623_), .A2(new_n624_), .B(new_n626_), .ZN(po041));
  NAND3_X1   g337(.A1(new_n609_), .A2(pi027), .A3(new_n588_), .ZN(new_n628_));
  INV_X1     g338(.I(pi100), .ZN(new_n629_));
  INV_X1     g339(.I(pi095), .ZN(new_n630_));
  NOR2_X1    g340(.A1(new_n630_), .A2(pi096), .ZN(new_n631_));
  NAND2_X1   g341(.A1(pi027), .A2(pi116), .ZN(new_n632_));
  NAND2_X1   g342(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  OAI22_X1   g343(.A1(new_n619_), .A2(new_n633_), .B1(new_n617_), .B2(pi027), .ZN(new_n634_));
  NAND2_X1   g344(.A1(new_n634_), .A2(new_n629_), .ZN(new_n635_));
  NOR2_X1    g345(.A1(pi053), .A2(pi058), .ZN(new_n636_));
  NAND3_X1   g346(.A1(new_n327_), .A2(new_n636_), .A3(new_n581_), .ZN(new_n637_));
  AOI21_X1   g347(.A1(new_n635_), .A2(new_n628_), .B(new_n637_), .ZN(po042));
  NOR3_X1    g348(.A1(new_n427_), .A2(pi027), .A3(pi116), .ZN(new_n639_));
  NAND3_X1   g349(.A1(new_n639_), .A2(new_n584_), .A3(new_n612_), .ZN(new_n640_));
  INV_X1     g350(.I(new_n639_), .ZN(new_n641_));
  NOR3_X1    g351(.A1(new_n641_), .A2(pi026), .A3(new_n589_), .ZN(new_n642_));
  NAND2_X1   g352(.A1(new_n597_), .A2(new_n596_), .ZN(new_n643_));
  NOR2_X1    g353(.A1(new_n592_), .A2(pi026), .ZN(new_n644_));
  NOR4_X1    g354(.A1(pi027), .A2(pi039), .A3(pi051), .A4(pi052), .ZN(new_n645_));
  OAI21_X1   g355(.A1(new_n644_), .A2(new_n645_), .B(new_n643_), .ZN(new_n646_));
  NAND2_X1   g356(.A1(new_n581_), .A2(pi027), .ZN(new_n647_));
  NAND2_X1   g357(.A1(new_n591_), .A2(pi026), .ZN(new_n648_));
  NAND2_X1   g358(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1   g359(.A1(new_n649_), .A2(new_n594_), .ZN(new_n650_));
  AOI21_X1   g360(.A1(new_n646_), .A2(new_n650_), .B(new_n427_), .ZN(new_n651_));
  INV_X1     g361(.I(new_n644_), .ZN(new_n652_));
  NOR3_X1    g362(.A1(pi026), .A2(pi100), .A3(pi110), .ZN(new_n653_));
  AOI22_X1   g363(.A1(new_n595_), .A2(new_n608_), .B1(new_n631_), .B2(new_n653_), .ZN(new_n654_));
  OAI22_X1   g364(.A1(new_n654_), .A2(pi027), .B1(new_n652_), .B2(new_n632_), .ZN(new_n655_));
  OAI21_X1   g365(.A1(new_n651_), .A2(new_n655_), .B(new_n588_), .ZN(new_n656_));
  NOR2_X1    g366(.A1(new_n594_), .A2(pi100), .ZN(new_n657_));
  NOR2_X1    g367(.A1(new_n427_), .A2(pi116), .ZN(new_n658_));
  NOR3_X1    g368(.A1(new_n588_), .A2(pi026), .A3(pi027), .ZN(new_n659_));
  OAI21_X1   g369(.A1(new_n657_), .A2(new_n658_), .B(new_n659_), .ZN(new_n660_));
  AOI21_X1   g370(.A1(new_n656_), .A2(new_n660_), .B(pi053), .ZN(new_n661_));
  OAI21_X1   g371(.A1(new_n661_), .A2(new_n642_), .B(new_n583_), .ZN(new_n662_));
  AOI21_X1   g372(.A1(new_n662_), .A2(new_n640_), .B(new_n413_), .ZN(po043));
  NOR2_X1    g373(.A1(new_n478_), .A2(pi116), .ZN(new_n664_));
  AND3_X2    g374(.A1(new_n664_), .A2(pi085), .A3(new_n625_), .Z(new_n665_));
  NAND3_X1   g375(.A1(new_n664_), .A2(pi027), .A3(new_n636_), .ZN(new_n666_));
  NOR2_X1    g376(.A1(new_n478_), .A2(new_n596_), .ZN(new_n667_));
  OR2_X2     g377(.A1(pi095), .A2(pi100), .Z(new_n668_));
  NAND3_X1   g378(.A1(new_n620_), .A2(new_n596_), .A3(pi097), .ZN(new_n669_));
  INV_X1     g379(.I(pi097), .ZN(new_n670_));
  NAND2_X1   g380(.A1(new_n670_), .A2(pi029), .ZN(new_n671_));
  AOI21_X1   g381(.A1(new_n669_), .A2(new_n671_), .B(new_n668_), .ZN(new_n672_));
  OAI21_X1   g382(.A1(new_n672_), .A2(new_n667_), .B(new_n583_), .ZN(new_n673_));
  NOR2_X1    g383(.A1(new_n670_), .A2(new_n594_), .ZN(new_n674_));
  OAI21_X1   g384(.A1(new_n674_), .A2(new_n664_), .B(pi058), .ZN(new_n675_));
  AOI21_X1   g385(.A1(new_n673_), .A2(new_n675_), .B(pi053), .ZN(new_n676_));
  INV_X1     g386(.I(pi053), .ZN(new_n677_));
  NOR2_X1    g387(.A1(new_n677_), .A2(pi058), .ZN(new_n678_));
  INV_X1     g388(.I(new_n678_), .ZN(new_n679_));
  NOR3_X1    g389(.A1(new_n679_), .A2(new_n478_), .A3(pi116), .ZN(new_n680_));
  OAI21_X1   g390(.A1(new_n676_), .A2(new_n680_), .B(new_n591_), .ZN(new_n681_));
  AOI21_X1   g391(.A1(new_n681_), .A2(new_n666_), .B(pi085), .ZN(new_n682_));
  OAI21_X1   g392(.A1(new_n682_), .A2(new_n665_), .B(new_n581_), .ZN(new_n683_));
  NAND4_X1   g393(.A1(new_n664_), .A2(pi026), .A3(new_n585_), .A4(new_n636_), .ZN(new_n684_));
  AOI21_X1   g394(.A1(new_n683_), .A2(new_n684_), .B(new_n413_), .ZN(po044));
  INV_X1     g395(.I(pi106), .ZN(new_n686_));
  INV_X1     g396(.I(pi060), .ZN(new_n687_));
  INV_X1     g397(.I(pi109), .ZN(new_n688_));
  NOR2_X1    g398(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1     g399(.I(pi030), .ZN(new_n690_));
  NOR2_X1    g400(.A1(new_n690_), .A2(pi109), .ZN(new_n691_));
  OAI21_X1   g401(.A1(new_n689_), .A2(new_n691_), .B(new_n686_), .ZN(new_n692_));
  NAND2_X1   g402(.A1(pi088), .A2(pi106), .ZN(new_n693_));
  AOI21_X1   g403(.A1(new_n692_), .A2(new_n693_), .B(pi129), .ZN(po045));
  NOR2_X1    g404(.A1(new_n690_), .A2(new_n688_), .ZN(new_n695_));
  INV_X1     g405(.I(pi031), .ZN(new_n696_));
  NOR2_X1    g406(.A1(new_n696_), .A2(pi109), .ZN(new_n697_));
  OAI21_X1   g407(.A1(new_n695_), .A2(new_n697_), .B(new_n686_), .ZN(new_n698_));
  NAND2_X1   g408(.A1(pi089), .A2(pi106), .ZN(new_n699_));
  AOI21_X1   g409(.A1(new_n698_), .A2(new_n699_), .B(pi129), .ZN(po046));
  NOR2_X1    g410(.A1(new_n696_), .A2(new_n688_), .ZN(new_n701_));
  INV_X1     g411(.I(pi032), .ZN(new_n702_));
  NOR2_X1    g412(.A1(new_n702_), .A2(pi109), .ZN(new_n703_));
  OAI21_X1   g413(.A1(new_n701_), .A2(new_n703_), .B(new_n686_), .ZN(new_n704_));
  NAND2_X1   g414(.A1(pi099), .A2(pi106), .ZN(new_n705_));
  AOI21_X1   g415(.A1(new_n704_), .A2(new_n705_), .B(pi129), .ZN(po047));
  NOR2_X1    g416(.A1(new_n702_), .A2(new_n688_), .ZN(new_n707_));
  INV_X1     g417(.I(pi033), .ZN(new_n708_));
  NOR2_X1    g418(.A1(new_n708_), .A2(pi109), .ZN(new_n709_));
  OAI21_X1   g419(.A1(new_n707_), .A2(new_n709_), .B(new_n686_), .ZN(new_n710_));
  NAND2_X1   g420(.A1(pi090), .A2(pi106), .ZN(new_n711_));
  AOI21_X1   g421(.A1(new_n710_), .A2(new_n711_), .B(pi129), .ZN(po048));
  NOR2_X1    g422(.A1(new_n708_), .A2(new_n688_), .ZN(new_n713_));
  INV_X1     g423(.I(pi034), .ZN(new_n714_));
  NOR2_X1    g424(.A1(new_n714_), .A2(pi109), .ZN(new_n715_));
  OAI21_X1   g425(.A1(new_n713_), .A2(new_n715_), .B(new_n686_), .ZN(new_n716_));
  NAND2_X1   g426(.A1(pi091), .A2(pi106), .ZN(new_n717_));
  AOI21_X1   g427(.A1(new_n716_), .A2(new_n717_), .B(pi129), .ZN(po049));
  NOR2_X1    g428(.A1(new_n714_), .A2(new_n688_), .ZN(new_n719_));
  INV_X1     g429(.I(pi035), .ZN(new_n720_));
  NOR2_X1    g430(.A1(new_n720_), .A2(pi109), .ZN(new_n721_));
  OAI21_X1   g431(.A1(new_n719_), .A2(new_n721_), .B(new_n686_), .ZN(new_n722_));
  NAND2_X1   g432(.A1(pi092), .A2(pi106), .ZN(new_n723_));
  AOI21_X1   g433(.A1(new_n722_), .A2(new_n723_), .B(pi129), .ZN(po050));
  NOR2_X1    g434(.A1(new_n720_), .A2(new_n688_), .ZN(new_n725_));
  INV_X1     g435(.I(pi036), .ZN(new_n726_));
  NOR2_X1    g436(.A1(new_n726_), .A2(pi109), .ZN(new_n727_));
  OAI21_X1   g437(.A1(new_n725_), .A2(new_n727_), .B(new_n686_), .ZN(new_n728_));
  NAND2_X1   g438(.A1(pi098), .A2(pi106), .ZN(new_n729_));
  AOI21_X1   g439(.A1(new_n728_), .A2(new_n729_), .B(pi129), .ZN(po051));
  NOR2_X1    g440(.A1(new_n726_), .A2(new_n688_), .ZN(new_n731_));
  INV_X1     g441(.I(pi037), .ZN(new_n732_));
  NOR2_X1    g442(.A1(new_n732_), .A2(pi109), .ZN(new_n733_));
  OAI21_X1   g443(.A1(new_n731_), .A2(new_n733_), .B(new_n686_), .ZN(new_n734_));
  NAND2_X1   g444(.A1(pi093), .A2(pi106), .ZN(new_n735_));
  AOI21_X1   g445(.A1(new_n734_), .A2(new_n735_), .B(pi129), .ZN(po052));
  NAND2_X1   g446(.A1(new_n495_), .A2(new_n389_), .ZN(new_n737_));
  NAND2_X1   g447(.A1(new_n380_), .A2(new_n572_), .ZN(new_n738_));
  OAI21_X1   g448(.A1(new_n738_), .A2(new_n737_), .B(pi082), .ZN(new_n739_));
  AOI22_X1   g449(.A1(new_n739_), .A2(new_n384_), .B1(pi082), .B2(new_n375_), .ZN(new_n740_));
  NOR2_X1    g450(.A1(new_n740_), .A2(pi038), .ZN(new_n741_));
  INV_X1     g451(.I(pi074), .ZN(new_n742_));
  INV_X1     g452(.I(pi048), .ZN(new_n743_));
  NAND4_X1   g453(.A1(new_n393_), .A2(new_n365_), .A3(new_n743_), .A4(new_n397_), .ZN(new_n744_));
  NOR4_X1    g454(.A1(new_n744_), .A2(pi050), .A3(new_n375_), .A4(new_n530_), .ZN(new_n745_));
  NOR2_X1    g455(.A1(new_n745_), .A2(new_n364_), .ZN(new_n746_));
  NOR3_X1    g456(.A1(new_n746_), .A2(new_n742_), .A3(new_n384_), .ZN(new_n747_));
  INV_X1     g457(.I(new_n539_), .ZN(new_n748_));
  NOR2_X1    g458(.A1(new_n364_), .A2(pi044), .ZN(new_n749_));
  AND3_X2    g459(.A1(new_n748_), .A2(pi038), .A3(new_n749_), .Z(new_n750_));
  NOR4_X1    g460(.A1(new_n747_), .A2(new_n741_), .A3(pi129), .A4(new_n750_), .ZN(po053));
  NOR2_X1    g461(.A1(pi051), .A2(pi052), .ZN(new_n752_));
  NAND2_X1   g462(.A1(new_n752_), .A2(pi109), .ZN(new_n753_));
  NAND2_X1   g463(.A1(new_n753_), .A2(pi039), .ZN(new_n754_));
  NOR2_X1    g464(.A1(pi039), .A2(pi052), .ZN(new_n755_));
  NOR2_X1    g465(.A1(new_n688_), .A2(pi051), .ZN(new_n756_));
  AOI21_X1   g466(.A1(new_n756_), .A2(new_n755_), .B(pi106), .ZN(new_n757_));
  AOI21_X1   g467(.A1(new_n754_), .A2(new_n757_), .B(pi129), .ZN(po054));
  NOR3_X1    g468(.A1(new_n738_), .A2(new_n371_), .A3(new_n496_), .ZN(new_n759_));
  OAI21_X1   g469(.A1(new_n759_), .A2(new_n364_), .B(new_n384_), .ZN(new_n760_));
  NAND2_X1   g470(.A1(new_n373_), .A2(pi082), .ZN(new_n761_));
  AOI21_X1   g471(.A1(new_n760_), .A2(new_n761_), .B(pi040), .ZN(new_n762_));
  INV_X1     g472(.I(pi073), .ZN(new_n763_));
  NOR4_X1    g473(.A1(new_n744_), .A2(new_n500_), .A3(new_n373_), .A4(new_n530_), .ZN(new_n764_));
  NOR2_X1    g474(.A1(new_n764_), .A2(new_n364_), .ZN(new_n765_));
  NOR3_X1    g475(.A1(new_n765_), .A2(new_n763_), .A3(new_n384_), .ZN(new_n766_));
  NOR3_X1    g476(.A1(new_n373_), .A2(new_n537_), .A3(new_n364_), .ZN(new_n767_));
  NOR4_X1    g477(.A1(new_n766_), .A2(new_n762_), .A3(pi129), .A4(new_n767_), .ZN(po055));
  OAI21_X1   g478(.A1(new_n738_), .A2(new_n496_), .B(pi082), .ZN(new_n769_));
  AOI22_X1   g479(.A1(new_n769_), .A2(new_n384_), .B1(pi082), .B2(new_n502_), .ZN(new_n770_));
  NOR2_X1    g480(.A1(new_n770_), .A2(pi041), .ZN(new_n771_));
  INV_X1     g481(.I(new_n744_), .ZN(new_n772_));
  NAND2_X1   g482(.A1(new_n372_), .A2(new_n388_), .ZN(new_n773_));
  NOR4_X1    g483(.A1(new_n773_), .A2(pi046), .A3(new_n494_), .A4(pi050), .ZN(new_n774_));
  AOI21_X1   g484(.A1(new_n772_), .A2(new_n774_), .B(new_n364_), .ZN(new_n775_));
  NAND2_X1   g485(.A1(new_n383_), .A2(pi076), .ZN(new_n776_));
  NOR4_X1    g486(.A1(pi038), .A2(pi040), .A3(pi046), .A4(pi050), .ZN(new_n777_));
  AND3_X2    g487(.A1(new_n372_), .A2(pi041), .A3(pi082), .Z(new_n778_));
  AOI21_X1   g488(.A1(new_n778_), .A2(new_n777_), .B(pi129), .ZN(new_n779_));
  OAI21_X1   g489(.A1(new_n775_), .A2(new_n776_), .B(new_n779_), .ZN(new_n780_));
  NOR2_X1    g490(.A1(new_n771_), .A2(new_n780_), .ZN(po056));
  NAND2_X1   g491(.A1(new_n562_), .A2(new_n777_), .ZN(new_n782_));
  OAI21_X1   g492(.A1(new_n744_), .A2(new_n782_), .B(pi082), .ZN(new_n783_));
  AOI22_X1   g493(.A1(new_n783_), .A2(new_n384_), .B1(pi044), .B2(pi082), .ZN(new_n784_));
  NOR2_X1    g494(.A1(new_n784_), .A2(pi042), .ZN(new_n785_));
  INV_X1     g495(.I(pi072), .ZN(new_n786_));
  NOR2_X1    g496(.A1(new_n533_), .A2(pi044), .ZN(new_n787_));
  NOR2_X1    g497(.A1(new_n744_), .A2(new_n530_), .ZN(new_n788_));
  AOI21_X1   g498(.A1(new_n788_), .A2(new_n787_), .B(new_n364_), .ZN(new_n789_));
  NOR3_X1    g499(.A1(new_n789_), .A2(new_n786_), .A3(new_n384_), .ZN(new_n790_));
  INV_X1     g500(.I(new_n749_), .ZN(new_n791_));
  NOR2_X1    g501(.A1(new_n791_), .A2(new_n538_), .ZN(new_n792_));
  NOR4_X1    g502(.A1(new_n785_), .A2(new_n790_), .A3(pi129), .A4(new_n792_), .ZN(po057));
  OR3_X2     g503(.A1(new_n744_), .A2(pi047), .A3(new_n390_), .Z(new_n794_));
  NAND2_X1   g504(.A1(new_n383_), .A2(pi077), .ZN(new_n795_));
  AOI21_X1   g505(.A1(new_n794_), .A2(pi082), .B(new_n795_), .ZN(new_n796_));
  NAND2_X1   g506(.A1(new_n390_), .A2(pi082), .ZN(new_n797_));
  NOR3_X1    g507(.A1(new_n381_), .A2(new_n396_), .A3(new_n571_), .ZN(new_n798_));
  OAI21_X1   g508(.A1(new_n798_), .A2(new_n364_), .B(new_n384_), .ZN(new_n799_));
  AOI21_X1   g509(.A1(new_n799_), .A2(new_n797_), .B(pi043), .ZN(new_n800_));
  INV_X1     g510(.I(pi043), .ZN(new_n801_));
  NOR4_X1    g511(.A1(new_n791_), .A2(new_n371_), .A3(new_n801_), .A4(new_n539_), .ZN(new_n802_));
  NOR4_X1    g512(.A1(new_n800_), .A2(new_n796_), .A3(pi129), .A4(new_n802_), .ZN(po058));
  NAND3_X1   g513(.A1(new_n540_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n804_));
  OAI21_X1   g514(.A1(new_n744_), .A2(new_n804_), .B(pi082), .ZN(new_n805_));
  NAND2_X1   g515(.A1(new_n383_), .A2(pi067), .ZN(new_n806_));
  OAI21_X1   g516(.A1(pi044), .A2(new_n383_), .B(new_n806_), .ZN(new_n807_));
  OAI21_X1   g517(.A1(new_n536_), .A2(new_n364_), .B(new_n558_), .ZN(new_n808_));
  AOI21_X1   g518(.A1(new_n805_), .A2(new_n807_), .B(new_n808_), .ZN(po059));
  OAI21_X1   g519(.A1(new_n566_), .A2(pi024), .B(pi082), .ZN(new_n810_));
  NAND2_X1   g520(.A1(new_n810_), .A2(new_n384_), .ZN(new_n811_));
  NAND2_X1   g521(.A1(new_n374_), .A2(new_n370_), .ZN(new_n812_));
  NAND2_X1   g522(.A1(new_n576_), .A2(new_n395_), .ZN(new_n813_));
  OAI21_X1   g523(.A1(new_n812_), .A2(new_n813_), .B(pi082), .ZN(new_n814_));
  AOI21_X1   g524(.A1(new_n814_), .A2(new_n811_), .B(pi045), .ZN(new_n815_));
  NAND4_X1   g525(.A1(new_n391_), .A2(new_n365_), .A3(new_n380_), .A4(new_n395_), .ZN(new_n816_));
  NAND2_X1   g526(.A1(new_n383_), .A2(pi068), .ZN(new_n817_));
  AOI21_X1   g527(.A1(new_n816_), .A2(pi082), .B(new_n817_), .ZN(new_n818_));
  NOR2_X1    g528(.A1(new_n539_), .A2(pi038), .ZN(new_n819_));
  NAND3_X1   g529(.A1(new_n819_), .A2(pi045), .A3(new_n749_), .ZN(new_n820_));
  NOR2_X1    g530(.A1(new_n820_), .A2(new_n737_), .ZN(new_n821_));
  NOR4_X1    g531(.A1(new_n815_), .A2(new_n818_), .A3(pi129), .A4(new_n821_), .ZN(po060));
  NAND2_X1   g532(.A1(new_n812_), .A2(pi082), .ZN(new_n823_));
  NOR3_X1    g533(.A1(new_n744_), .A2(pi047), .A3(new_n561_), .ZN(new_n824_));
  OAI21_X1   g534(.A1(new_n824_), .A2(new_n364_), .B(new_n384_), .ZN(new_n825_));
  AOI21_X1   g535(.A1(new_n825_), .A2(new_n823_), .B(pi046), .ZN(new_n826_));
  NOR2_X1    g536(.A1(new_n773_), .A2(pi050), .ZN(new_n827_));
  AOI21_X1   g537(.A1(new_n824_), .A2(new_n827_), .B(new_n364_), .ZN(new_n828_));
  NAND2_X1   g538(.A1(new_n383_), .A2(pi075), .ZN(new_n829_));
  AND2_X2    g539(.A1(pi046), .A2(pi082), .Z(new_n830_));
  AOI21_X1   g540(.A1(new_n827_), .A2(new_n830_), .B(pi129), .ZN(new_n831_));
  OAI21_X1   g541(.A1(new_n828_), .A2(new_n829_), .B(new_n831_), .ZN(new_n832_));
  NOR2_X1    g542(.A1(new_n826_), .A2(new_n832_), .ZN(po061));
  INV_X1     g543(.I(pi064), .ZN(new_n834_));
  AOI21_X1   g544(.A1(new_n772_), .A2(new_n391_), .B(new_n364_), .ZN(new_n835_));
  NOR3_X1    g545(.A1(new_n835_), .A2(new_n834_), .A3(new_n384_), .ZN(new_n836_));
  NAND2_X1   g546(.A1(new_n392_), .A2(pi082), .ZN(new_n837_));
  OAI21_X1   g547(.A1(new_n772_), .A2(new_n364_), .B(new_n384_), .ZN(new_n838_));
  AOI21_X1   g548(.A1(new_n838_), .A2(new_n837_), .B(pi047), .ZN(new_n839_));
  NOR2_X1    g549(.A1(new_n791_), .A2(new_n539_), .ZN(new_n840_));
  NAND4_X1   g550(.A1(new_n840_), .A2(pi047), .A3(new_n501_), .A4(new_n504_), .ZN(new_n841_));
  NAND2_X1   g551(.A1(new_n841_), .A2(new_n558_), .ZN(new_n842_));
  NOR3_X1    g552(.A1(new_n836_), .A2(new_n839_), .A3(new_n842_), .ZN(po062));
  OAI21_X1   g553(.A1(new_n812_), .A2(new_n530_), .B(pi082), .ZN(new_n844_));
  NAND2_X1   g554(.A1(new_n738_), .A2(pi082), .ZN(new_n845_));
  NAND2_X1   g555(.A1(new_n845_), .A2(new_n384_), .ZN(new_n846_));
  AOI21_X1   g556(.A1(new_n846_), .A2(new_n844_), .B(pi048), .ZN(new_n847_));
  INV_X1     g557(.I(pi062), .ZN(new_n848_));
  NAND2_X1   g558(.A1(new_n393_), .A2(new_n397_), .ZN(new_n849_));
  NOR3_X1    g559(.A1(new_n849_), .A2(pi002), .A3(pi047), .ZN(new_n850_));
  AOI21_X1   g560(.A1(new_n850_), .A2(new_n391_), .B(new_n364_), .ZN(new_n851_));
  NOR3_X1    g561(.A1(new_n851_), .A2(new_n848_), .A3(new_n384_), .ZN(new_n852_));
  NAND2_X1   g562(.A1(new_n819_), .A2(new_n389_), .ZN(new_n853_));
  NOR4_X1    g563(.A1(new_n853_), .A2(new_n743_), .A3(new_n494_), .A4(new_n791_), .ZN(new_n854_));
  NOR4_X1    g564(.A1(new_n852_), .A2(pi129), .A3(new_n847_), .A4(new_n854_), .ZN(po063));
  NOR3_X1    g565(.A1(new_n577_), .A2(pi024), .A3(pi042), .ZN(new_n856_));
  AOI21_X1   g566(.A1(new_n856_), .A2(new_n787_), .B(new_n565_), .ZN(new_n857_));
  NAND2_X1   g567(.A1(new_n827_), .A2(new_n376_), .ZN(new_n858_));
  NOR2_X1    g568(.A1(new_n379_), .A2(pi002), .ZN(new_n859_));
  NOR4_X1    g569(.A1(new_n858_), .A2(new_n529_), .A3(new_n530_), .A4(new_n859_), .ZN(new_n860_));
  OAI21_X1   g570(.A1(new_n860_), .A2(new_n857_), .B(pi082), .ZN(new_n861_));
  OAI21_X1   g571(.A1(new_n858_), .A2(new_n577_), .B(pi082), .ZN(new_n862_));
  NOR2_X1    g572(.A1(new_n384_), .A2(pi069), .ZN(new_n863_));
  AOI22_X1   g573(.A1(new_n862_), .A2(new_n863_), .B1(pi049), .B2(new_n387_), .ZN(new_n864_));
  AOI21_X1   g574(.A1(new_n864_), .A2(new_n861_), .B(pi129), .ZN(po064));
  NAND3_X1   g575(.A1(new_n576_), .A2(new_n395_), .A3(new_n365_), .ZN(new_n866_));
  OAI21_X1   g576(.A1(new_n849_), .A2(new_n866_), .B(pi082), .ZN(new_n867_));
  AOI22_X1   g577(.A1(new_n867_), .A2(new_n384_), .B1(pi082), .B2(new_n773_), .ZN(new_n868_));
  NOR2_X1    g578(.A1(new_n868_), .A2(pi050), .ZN(new_n869_));
  INV_X1     g579(.I(pi066), .ZN(new_n870_));
  NOR2_X1    g580(.A1(new_n773_), .A2(new_n530_), .ZN(new_n871_));
  AOI21_X1   g581(.A1(new_n772_), .A2(new_n871_), .B(new_n364_), .ZN(new_n872_));
  NOR3_X1    g582(.A1(new_n872_), .A2(new_n870_), .A3(new_n384_), .ZN(new_n873_));
  NOR4_X1    g583(.A1(new_n791_), .A2(pi038), .A3(new_n532_), .A4(new_n539_), .ZN(new_n874_));
  NOR4_X1    g584(.A1(new_n869_), .A2(new_n873_), .A3(pi129), .A4(new_n874_), .ZN(po065));
  NAND2_X1   g585(.A1(new_n688_), .A2(pi051), .ZN(new_n876_));
  NOR2_X1    g586(.A1(new_n756_), .A2(pi106), .ZN(new_n877_));
  AOI21_X1   g587(.A1(new_n877_), .A2(new_n876_), .B(pi129), .ZN(po066));
  OAI21_X1   g588(.A1(new_n688_), .A2(pi051), .B(pi052), .ZN(new_n879_));
  AOI21_X1   g589(.A1(new_n752_), .A2(pi109), .B(pi106), .ZN(new_n880_));
  AOI21_X1   g590(.A1(new_n880_), .A2(new_n879_), .B(pi129), .ZN(po067));
  NAND3_X1   g591(.A1(new_n583_), .A2(new_n620_), .A3(new_n596_), .ZN(new_n882_));
  OAI22_X1   g592(.A1(new_n882_), .A2(new_n668_), .B1(new_n583_), .B2(new_n594_), .ZN(new_n883_));
  NAND3_X1   g593(.A1(new_n883_), .A2(new_n677_), .A3(pi097), .ZN(new_n884_));
  NAND2_X1   g594(.A1(new_n678_), .A2(new_n594_), .ZN(new_n885_));
  NAND3_X1   g595(.A1(new_n327_), .A2(new_n585_), .A3(new_n581_), .ZN(new_n886_));
  AOI21_X1   g596(.A1(new_n884_), .A2(new_n885_), .B(new_n886_), .ZN(po068));
  AOI21_X1   g597(.A1(new_n798_), .A2(new_n391_), .B(new_n364_), .ZN(new_n888_));
  OAI21_X1   g598(.A1(new_n888_), .A2(new_n384_), .B(new_n558_), .ZN(po069));
  INV_X1     g599(.I(pi114), .ZN(new_n890_));
  NAND2_X1   g600(.A1(new_n404_), .A2(new_n558_), .ZN(po129));
  NOR3_X1    g601(.A1(po129), .A2(new_n890_), .A3(pi122), .ZN(po070));
  NOR2_X1    g602(.A1(new_n732_), .A2(pi026), .ZN(new_n893_));
  NAND3_X1   g603(.A1(new_n893_), .A2(new_n588_), .A3(new_n636_), .ZN(new_n894_));
  INV_X1     g604(.I(pi094), .ZN(new_n895_));
  NAND2_X1   g605(.A1(new_n581_), .A2(pi058), .ZN(new_n896_));
  NAND2_X1   g606(.A1(new_n595_), .A2(new_n583_), .ZN(new_n897_));
  AOI21_X1   g607(.A1(new_n897_), .A2(new_n896_), .B(new_n895_), .ZN(new_n898_));
  NAND2_X1   g608(.A1(new_n594_), .A2(pi037), .ZN(new_n899_));
  AOI22_X1   g609(.A1(new_n896_), .A2(new_n899_), .B1(pi058), .B2(new_n594_), .ZN(new_n900_));
  OAI21_X1   g610(.A1(new_n898_), .A2(new_n900_), .B(new_n677_), .ZN(new_n901_));
  NAND2_X1   g611(.A1(new_n893_), .A2(new_n583_), .ZN(new_n902_));
  AOI21_X1   g612(.A1(new_n901_), .A2(new_n902_), .B(pi085), .ZN(new_n903_));
  INV_X1     g613(.I(new_n636_), .ZN(new_n904_));
  NOR3_X1    g614(.A1(new_n904_), .A2(pi026), .A3(new_n732_), .ZN(new_n905_));
  OAI21_X1   g615(.A1(new_n903_), .A2(new_n905_), .B(new_n591_), .ZN(new_n906_));
  AOI21_X1   g616(.A1(new_n906_), .A2(new_n894_), .B(new_n413_), .ZN(po071));
  NOR2_X1    g617(.A1(pi026), .A2(pi053), .ZN(new_n908_));
  NAND2_X1   g618(.A1(new_n908_), .A2(new_n588_), .ZN(new_n909_));
  INV_X1     g619(.I(new_n909_), .ZN(new_n910_));
  NAND3_X1   g620(.A1(new_n910_), .A2(pi057), .A3(new_n583_), .ZN(new_n911_));
  INV_X1     g621(.I(pi057), .ZN(new_n912_));
  AOI21_X1   g622(.A1(pi026), .A2(pi053), .B(pi085), .ZN(new_n913_));
  OAI21_X1   g623(.A1(new_n913_), .A2(new_n908_), .B(new_n583_), .ZN(new_n914_));
  NAND2_X1   g624(.A1(new_n910_), .A2(new_n594_), .ZN(new_n915_));
  AOI21_X1   g625(.A1(new_n915_), .A2(new_n914_), .B(new_n912_), .ZN(new_n916_));
  NOR4_X1    g626(.A1(new_n909_), .A2(new_n583_), .A3(new_n687_), .A4(new_n594_), .ZN(new_n917_));
  OAI21_X1   g627(.A1(new_n916_), .A2(new_n917_), .B(new_n591_), .ZN(new_n918_));
  AOI21_X1   g628(.A1(new_n918_), .A2(new_n911_), .B(new_n413_), .ZN(po072));
  NAND4_X1   g629(.A1(new_n581_), .A2(new_n591_), .A3(new_n594_), .A4(pi058), .ZN(new_n920_));
  NAND4_X1   g630(.A1(new_n649_), .A2(new_n583_), .A3(pi116), .A4(new_n608_), .ZN(new_n921_));
  NAND3_X1   g631(.A1(new_n327_), .A2(new_n677_), .A3(new_n588_), .ZN(new_n922_));
  AOI21_X1   g632(.A1(new_n921_), .A2(new_n920_), .B(new_n922_), .ZN(po073));
  NOR2_X1    g633(.A1(new_n419_), .A2(pi116), .ZN(new_n924_));
  NAND4_X1   g634(.A1(new_n924_), .A2(pi026), .A3(new_n585_), .A4(new_n636_), .ZN(new_n925_));
  INV_X1     g635(.I(new_n924_), .ZN(new_n926_));
  NOR4_X1    g636(.A1(new_n926_), .A2(new_n591_), .A3(pi085), .A4(new_n904_), .ZN(new_n927_));
  NOR3_X1    g637(.A1(new_n643_), .A2(new_n620_), .A3(new_n904_), .ZN(new_n928_));
  NAND2_X1   g638(.A1(new_n643_), .A2(new_n636_), .ZN(new_n929_));
  OAI21_X1   g639(.A1(new_n584_), .A2(new_n678_), .B(new_n594_), .ZN(new_n930_));
  AOI21_X1   g640(.A1(new_n929_), .A2(new_n930_), .B(new_n419_), .ZN(new_n931_));
  OAI21_X1   g641(.A1(new_n931_), .A2(new_n928_), .B(new_n588_), .ZN(new_n932_));
  NAND3_X1   g642(.A1(new_n924_), .A2(pi085), .A3(new_n636_), .ZN(new_n933_));
  AOI21_X1   g643(.A1(new_n932_), .A2(new_n933_), .B(pi027), .ZN(new_n934_));
  OAI21_X1   g644(.A1(new_n934_), .A2(new_n927_), .B(new_n581_), .ZN(new_n935_));
  AOI21_X1   g645(.A1(new_n935_), .A2(new_n925_), .B(new_n413_), .ZN(po074));
  NOR2_X1    g646(.A1(pi117), .A2(pi122), .ZN(new_n937_));
  MUX2_X1    g647(.I0(pi060), .I1(pi123), .S(new_n937_), .Z(po075));
  NOR4_X1    g648(.A1(new_n404_), .A2(pi114), .A3(pi122), .A4(pi129), .ZN(po076));
  NAND3_X1   g649(.A1(pi131), .A2(pi132), .A3(pi133), .ZN(new_n940_));
  NOR2_X1    g650(.A1(new_n940_), .A2(pi138), .ZN(new_n941_));
  INV_X1     g651(.I(new_n941_), .ZN(new_n942_));
  INV_X1     g652(.I(pi136), .ZN(new_n943_));
  NOR2_X1    g653(.A1(new_n943_), .A2(pi137), .ZN(new_n944_));
  INV_X1     g654(.I(new_n944_), .ZN(new_n945_));
  NOR3_X1    g655(.A1(new_n942_), .A2(pi140), .A3(new_n945_), .ZN(new_n946_));
  NOR3_X1    g656(.A1(new_n945_), .A2(pi138), .A3(new_n940_), .ZN(new_n947_));
  NOR2_X1    g657(.A1(new_n947_), .A2(new_n848_), .ZN(new_n948_));
  OAI21_X1   g658(.A1(new_n948_), .A2(new_n946_), .B(new_n558_), .ZN(po077));
  NOR3_X1    g659(.A1(new_n942_), .A2(pi142), .A3(new_n945_), .ZN(new_n950_));
  INV_X1     g660(.I(pi063), .ZN(new_n951_));
  NOR2_X1    g661(.A1(new_n947_), .A2(new_n951_), .ZN(new_n952_));
  OAI21_X1   g662(.A1(new_n952_), .A2(new_n950_), .B(new_n558_), .ZN(po078));
  NOR3_X1    g663(.A1(new_n942_), .A2(pi139), .A3(new_n945_), .ZN(new_n954_));
  NOR2_X1    g664(.A1(new_n947_), .A2(new_n834_), .ZN(new_n955_));
  OAI21_X1   g665(.A1(new_n955_), .A2(new_n954_), .B(new_n558_), .ZN(po079));
  NOR3_X1    g666(.A1(new_n942_), .A2(pi146), .A3(new_n945_), .ZN(new_n957_));
  INV_X1     g667(.I(pi065), .ZN(new_n958_));
  NOR2_X1    g668(.A1(new_n947_), .A2(new_n958_), .ZN(new_n959_));
  OAI21_X1   g669(.A1(new_n959_), .A2(new_n957_), .B(new_n558_), .ZN(po080));
  NOR2_X1    g670(.A1(pi136), .A2(pi137), .ZN(new_n961_));
  NAND2_X1   g671(.A1(new_n941_), .A2(new_n961_), .ZN(new_n962_));
  INV_X1     g672(.I(new_n962_), .ZN(new_n963_));
  NOR2_X1    g673(.A1(new_n963_), .A2(new_n870_), .ZN(new_n964_));
  NOR2_X1    g674(.A1(new_n962_), .A2(pi143), .ZN(new_n965_));
  OAI21_X1   g675(.A1(new_n964_), .A2(new_n965_), .B(new_n558_), .ZN(po081));
  INV_X1     g676(.I(pi067), .ZN(new_n967_));
  NOR2_X1    g677(.A1(new_n963_), .A2(new_n967_), .ZN(new_n968_));
  NOR2_X1    g678(.A1(new_n962_), .A2(pi139), .ZN(new_n969_));
  OAI21_X1   g679(.A1(new_n968_), .A2(new_n969_), .B(new_n558_), .ZN(po082));
  NOR3_X1    g680(.A1(new_n942_), .A2(pi141), .A3(new_n945_), .ZN(new_n971_));
  INV_X1     g681(.I(pi068), .ZN(new_n972_));
  NOR2_X1    g682(.A1(new_n947_), .A2(new_n972_), .ZN(new_n973_));
  OAI21_X1   g683(.A1(new_n973_), .A2(new_n971_), .B(new_n558_), .ZN(po083));
  NOR3_X1    g684(.A1(new_n942_), .A2(pi143), .A3(new_n945_), .ZN(new_n975_));
  INV_X1     g685(.I(pi069), .ZN(new_n976_));
  NOR2_X1    g686(.A1(new_n947_), .A2(new_n976_), .ZN(new_n977_));
  OAI21_X1   g687(.A1(new_n977_), .A2(new_n975_), .B(new_n558_), .ZN(po084));
  NOR3_X1    g688(.A1(new_n942_), .A2(pi144), .A3(new_n945_), .ZN(new_n979_));
  INV_X1     g689(.I(pi070), .ZN(new_n980_));
  NOR2_X1    g690(.A1(new_n947_), .A2(new_n980_), .ZN(new_n981_));
  OAI21_X1   g691(.A1(new_n981_), .A2(new_n979_), .B(new_n558_), .ZN(po085));
  NOR3_X1    g692(.A1(new_n942_), .A2(pi145), .A3(new_n945_), .ZN(new_n983_));
  INV_X1     g693(.I(pi071), .ZN(new_n984_));
  NOR2_X1    g694(.A1(new_n947_), .A2(new_n984_), .ZN(new_n985_));
  OAI21_X1   g695(.A1(new_n985_), .A2(new_n983_), .B(new_n558_), .ZN(po086));
  NOR2_X1    g696(.A1(new_n963_), .A2(new_n786_), .ZN(new_n987_));
  NOR2_X1    g697(.A1(new_n962_), .A2(pi140), .ZN(new_n988_));
  OAI21_X1   g698(.A1(new_n987_), .A2(new_n988_), .B(new_n558_), .ZN(po087));
  NOR2_X1    g699(.A1(new_n963_), .A2(new_n763_), .ZN(new_n990_));
  NOR2_X1    g700(.A1(new_n962_), .A2(pi141), .ZN(new_n991_));
  OAI21_X1   g701(.A1(new_n990_), .A2(new_n991_), .B(new_n558_), .ZN(po088));
  NOR2_X1    g702(.A1(new_n963_), .A2(new_n742_), .ZN(new_n993_));
  NOR2_X1    g703(.A1(new_n962_), .A2(pi142), .ZN(new_n994_));
  OAI21_X1   g704(.A1(new_n993_), .A2(new_n994_), .B(new_n558_), .ZN(po089));
  INV_X1     g705(.I(pi075), .ZN(new_n996_));
  NOR2_X1    g706(.A1(new_n963_), .A2(new_n996_), .ZN(new_n997_));
  NOR2_X1    g707(.A1(new_n962_), .A2(pi144), .ZN(new_n998_));
  OAI21_X1   g708(.A1(new_n997_), .A2(new_n998_), .B(new_n558_), .ZN(po090));
  INV_X1     g709(.I(pi076), .ZN(new_n1000_));
  NOR2_X1    g710(.A1(new_n963_), .A2(new_n1000_), .ZN(new_n1001_));
  NOR2_X1    g711(.A1(new_n962_), .A2(pi145), .ZN(new_n1002_));
  OAI21_X1   g712(.A1(new_n1001_), .A2(new_n1002_), .B(new_n558_), .ZN(po091));
  INV_X1     g713(.I(pi077), .ZN(new_n1004_));
  NOR2_X1    g714(.A1(new_n963_), .A2(new_n1004_), .ZN(new_n1005_));
  NOR2_X1    g715(.A1(new_n962_), .A2(pi146), .ZN(new_n1006_));
  OAI21_X1   g716(.A1(new_n1005_), .A2(new_n1006_), .B(new_n558_), .ZN(po092));
  INV_X1     g717(.I(pi137), .ZN(new_n1008_));
  NOR2_X1    g718(.A1(new_n1008_), .A2(pi136), .ZN(new_n1009_));
  NAND2_X1   g719(.A1(new_n941_), .A2(new_n1009_), .ZN(new_n1010_));
  NAND2_X1   g720(.A1(new_n1010_), .A2(pi078), .ZN(new_n1011_));
  INV_X1     g721(.I(new_n1010_), .ZN(new_n1012_));
  NAND2_X1   g722(.A1(new_n1012_), .A2(pi142), .ZN(new_n1013_));
  AOI21_X1   g723(.A1(new_n1013_), .A2(new_n1011_), .B(pi129), .ZN(po093));
  NAND2_X1   g724(.A1(new_n1010_), .A2(pi079), .ZN(new_n1015_));
  NAND2_X1   g725(.A1(new_n1012_), .A2(pi143), .ZN(new_n1016_));
  AOI21_X1   g726(.A1(new_n1016_), .A2(new_n1015_), .B(pi129), .ZN(po094));
  NAND2_X1   g727(.A1(new_n1010_), .A2(pi080), .ZN(new_n1018_));
  NAND2_X1   g728(.A1(new_n1012_), .A2(pi144), .ZN(new_n1019_));
  AOI21_X1   g729(.A1(new_n1019_), .A2(new_n1018_), .B(pi129), .ZN(po095));
  NAND2_X1   g730(.A1(new_n1010_), .A2(pi081), .ZN(new_n1021_));
  NAND2_X1   g731(.A1(new_n1012_), .A2(pi145), .ZN(new_n1022_));
  AOI21_X1   g732(.A1(new_n1022_), .A2(new_n1021_), .B(pi129), .ZN(po096));
  NAND2_X1   g733(.A1(new_n1010_), .A2(pi082), .ZN(new_n1024_));
  NAND2_X1   g734(.A1(new_n1012_), .A2(pi146), .ZN(new_n1025_));
  AOI21_X1   g735(.A1(new_n1025_), .A2(new_n1024_), .B(pi129), .ZN(po097));
  INV_X1     g736(.I(pi115), .ZN(new_n1027_));
  NAND2_X1   g737(.A1(new_n1027_), .A2(pi138), .ZN(new_n1028_));
  INV_X1     g738(.I(pi138), .ZN(new_n1029_));
  NAND2_X1   g739(.A1(new_n1029_), .A2(pi087), .ZN(new_n1030_));
  AOI21_X1   g740(.A1(new_n1028_), .A2(new_n1030_), .B(pi136), .ZN(new_n1031_));
  NAND2_X1   g741(.A1(new_n1029_), .A2(pi136), .ZN(new_n1032_));
  NOR2_X1    g742(.A1(new_n1032_), .A2(new_n696_), .ZN(new_n1033_));
  OAI21_X1   g743(.A1(new_n1031_), .A2(new_n1033_), .B(pi137), .ZN(new_n1034_));
  NAND2_X1   g744(.A1(pi089), .A2(pi138), .ZN(new_n1035_));
  NAND2_X1   g745(.A1(new_n848_), .A2(new_n1029_), .ZN(new_n1036_));
  AOI21_X1   g746(.A1(new_n1036_), .A2(new_n1035_), .B(new_n943_), .ZN(new_n1037_));
  NAND2_X1   g747(.A1(pi119), .A2(pi138), .ZN(new_n1038_));
  NAND2_X1   g748(.A1(new_n786_), .A2(new_n1029_), .ZN(new_n1039_));
  AOI21_X1   g749(.A1(new_n1039_), .A2(new_n1038_), .B(pi136), .ZN(new_n1040_));
  OAI21_X1   g750(.A1(new_n1037_), .A2(new_n1040_), .B(new_n1008_), .ZN(new_n1041_));
  NAND2_X1   g751(.A1(new_n1041_), .A2(new_n1034_), .ZN(po098));
  NAND2_X1   g752(.A1(new_n1010_), .A2(pi084), .ZN(new_n1043_));
  NAND2_X1   g753(.A1(new_n1012_), .A2(pi141), .ZN(new_n1044_));
  AOI21_X1   g754(.A1(new_n1044_), .A2(new_n1043_), .B(pi129), .ZN(po099));
  AND3_X2    g755(.A1(new_n597_), .A2(new_n588_), .A3(new_n596_), .Z(new_n1046_));
  NAND2_X1   g756(.A1(new_n1046_), .A2(pi096), .ZN(new_n1047_));
  NAND3_X1   g757(.A1(new_n625_), .A2(new_n327_), .A3(new_n581_), .ZN(new_n1048_));
  AOI21_X1   g758(.A1(new_n1047_), .A2(new_n618_), .B(new_n1048_), .ZN(po100));
  NAND2_X1   g759(.A1(new_n1010_), .A2(pi086), .ZN(new_n1050_));
  NAND2_X1   g760(.A1(new_n1012_), .A2(pi139), .ZN(new_n1051_));
  AOI21_X1   g761(.A1(new_n1051_), .A2(new_n1050_), .B(pi129), .ZN(po101));
  NAND2_X1   g762(.A1(new_n1010_), .A2(pi087), .ZN(new_n1053_));
  NAND2_X1   g763(.A1(new_n1012_), .A2(pi140), .ZN(new_n1054_));
  AOI21_X1   g764(.A1(new_n1054_), .A2(new_n1053_), .B(pi129), .ZN(po102));
  NOR2_X1    g765(.A1(new_n943_), .A2(new_n1008_), .ZN(new_n1056_));
  NAND2_X1   g766(.A1(new_n941_), .A2(new_n1056_), .ZN(new_n1057_));
  NAND2_X1   g767(.A1(new_n1057_), .A2(pi088), .ZN(new_n1058_));
  INV_X1     g768(.I(new_n1057_), .ZN(new_n1059_));
  NAND2_X1   g769(.A1(new_n1059_), .A2(pi139), .ZN(new_n1060_));
  AOI21_X1   g770(.A1(new_n1060_), .A2(new_n1058_), .B(pi129), .ZN(po103));
  NAND2_X1   g771(.A1(new_n1057_), .A2(pi089), .ZN(new_n1062_));
  NAND2_X1   g772(.A1(new_n1059_), .A2(pi140), .ZN(new_n1063_));
  AOI21_X1   g773(.A1(new_n1063_), .A2(new_n1062_), .B(pi129), .ZN(po104));
  NAND2_X1   g774(.A1(new_n1057_), .A2(pi090), .ZN(new_n1065_));
  NAND2_X1   g775(.A1(new_n1059_), .A2(pi142), .ZN(new_n1066_));
  AOI21_X1   g776(.A1(new_n1066_), .A2(new_n1065_), .B(pi129), .ZN(po105));
  NAND2_X1   g777(.A1(new_n1057_), .A2(pi091), .ZN(new_n1068_));
  NAND2_X1   g778(.A1(new_n1059_), .A2(pi143), .ZN(new_n1069_));
  AOI21_X1   g779(.A1(new_n1069_), .A2(new_n1068_), .B(pi129), .ZN(po106));
  NAND2_X1   g780(.A1(new_n1057_), .A2(pi092), .ZN(new_n1071_));
  NAND2_X1   g781(.A1(new_n1059_), .A2(pi144), .ZN(new_n1072_));
  AOI21_X1   g782(.A1(new_n1072_), .A2(new_n1071_), .B(pi129), .ZN(po107));
  NAND2_X1   g783(.A1(new_n1057_), .A2(pi093), .ZN(new_n1074_));
  NAND2_X1   g784(.A1(new_n1059_), .A2(pi146), .ZN(new_n1075_));
  AOI21_X1   g785(.A1(new_n1075_), .A2(new_n1074_), .B(pi129), .ZN(po108));
  INV_X1     g786(.I(new_n940_), .ZN(new_n1077_));
  NOR3_X1    g787(.A1(new_n364_), .A2(pi136), .A3(pi137), .ZN(new_n1078_));
  NAND3_X1   g788(.A1(new_n1077_), .A2(new_n1078_), .A3(pi138), .ZN(new_n1079_));
  NAND2_X1   g789(.A1(new_n1079_), .A2(pi094), .ZN(new_n1080_));
  INV_X1     g790(.I(new_n1079_), .ZN(new_n1081_));
  NAND2_X1   g791(.A1(new_n1081_), .A2(pi142), .ZN(new_n1082_));
  AOI21_X1   g792(.A1(new_n1082_), .A2(new_n1080_), .B(pi129), .ZN(po109));
  NOR4_X1    g793(.A1(new_n364_), .A2(new_n1029_), .A3(pi136), .A4(pi137), .ZN(new_n1084_));
  INV_X1     g794(.I(pi003), .ZN(new_n1085_));
  NAND3_X1   g795(.A1(new_n940_), .A2(new_n1085_), .A3(new_n596_), .ZN(new_n1086_));
  OAI21_X1   g796(.A1(new_n940_), .A2(new_n1084_), .B(new_n1086_), .ZN(new_n1087_));
  AOI22_X1   g797(.A1(new_n1081_), .A2(pi143), .B1(new_n1087_), .B2(pi095), .ZN(new_n1088_));
  NOR2_X1    g798(.A1(new_n1088_), .A2(pi129), .ZN(po110));
  AOI22_X1   g799(.A1(new_n1081_), .A2(pi146), .B1(new_n1087_), .B2(pi096), .ZN(new_n1090_));
  NOR2_X1    g800(.A1(new_n1090_), .A2(pi129), .ZN(po111));
  AOI22_X1   g801(.A1(new_n1081_), .A2(pi145), .B1(new_n1087_), .B2(pi097), .ZN(new_n1092_));
  NOR2_X1    g802(.A1(new_n1092_), .A2(pi129), .ZN(po112));
  NAND2_X1   g803(.A1(new_n1057_), .A2(pi098), .ZN(new_n1094_));
  NAND2_X1   g804(.A1(new_n1059_), .A2(pi145), .ZN(new_n1095_));
  AOI21_X1   g805(.A1(new_n1095_), .A2(new_n1094_), .B(pi129), .ZN(po113));
  NAND2_X1   g806(.A1(new_n1057_), .A2(pi099), .ZN(new_n1097_));
  NAND2_X1   g807(.A1(new_n1059_), .A2(pi141), .ZN(new_n1098_));
  AOI21_X1   g808(.A1(new_n1098_), .A2(new_n1097_), .B(pi129), .ZN(po114));
  AOI22_X1   g809(.A1(new_n1081_), .A2(pi144), .B1(new_n1087_), .B2(pi100), .ZN(new_n1100_));
  NOR2_X1    g810(.A1(new_n1100_), .A2(pi129), .ZN(po115));
  NAND2_X1   g811(.A1(pi096), .A2(pi138), .ZN(new_n1102_));
  NAND2_X1   g812(.A1(new_n1029_), .A2(pi082), .ZN(new_n1103_));
  AOI21_X1   g813(.A1(new_n1103_), .A2(new_n1102_), .B(pi136), .ZN(new_n1104_));
  NOR2_X1    g814(.A1(new_n1032_), .A2(new_n732_), .ZN(new_n1105_));
  OAI21_X1   g815(.A1(new_n1104_), .A2(new_n1105_), .B(pi137), .ZN(new_n1106_));
  NAND2_X1   g816(.A1(pi124), .A2(pi138), .ZN(new_n1107_));
  NAND2_X1   g817(.A1(new_n1004_), .A2(new_n1029_), .ZN(new_n1108_));
  AOI21_X1   g818(.A1(new_n1108_), .A2(new_n1107_), .B(pi136), .ZN(new_n1109_));
  NAND2_X1   g819(.A1(pi093), .A2(pi138), .ZN(new_n1110_));
  NAND2_X1   g820(.A1(new_n958_), .A2(new_n1029_), .ZN(new_n1111_));
  AOI21_X1   g821(.A1(new_n1111_), .A2(new_n1110_), .B(new_n943_), .ZN(new_n1112_));
  OAI21_X1   g822(.A1(new_n1109_), .A2(new_n1112_), .B(new_n1008_), .ZN(new_n1113_));
  NAND2_X1   g823(.A1(new_n1113_), .A2(new_n1106_), .ZN(po116));
  AOI22_X1   g824(.A1(pi091), .A2(new_n944_), .B1(new_n1009_), .B2(pi095), .ZN(new_n1115_));
  NAND2_X1   g825(.A1(pi034), .A2(pi136), .ZN(new_n1116_));
  NAND2_X1   g826(.A1(new_n943_), .A2(pi079), .ZN(new_n1117_));
  AOI21_X1   g827(.A1(new_n1117_), .A2(new_n1116_), .B(new_n1008_), .ZN(new_n1118_));
  NAND2_X1   g828(.A1(new_n870_), .A2(new_n943_), .ZN(new_n1119_));
  NAND2_X1   g829(.A1(new_n976_), .A2(pi136), .ZN(new_n1120_));
  AOI21_X1   g830(.A1(new_n1119_), .A2(new_n1120_), .B(pi137), .ZN(new_n1121_));
  OAI21_X1   g831(.A1(new_n1121_), .A2(new_n1118_), .B(new_n1029_), .ZN(new_n1122_));
  OAI21_X1   g832(.A1(new_n1029_), .A2(new_n1115_), .B(new_n1122_), .ZN(po117));
  AOI22_X1   g833(.A1(pi090), .A2(new_n944_), .B1(new_n1009_), .B2(pi094), .ZN(new_n1124_));
  NAND2_X1   g834(.A1(pi033), .A2(pi136), .ZN(new_n1125_));
  NAND2_X1   g835(.A1(new_n943_), .A2(pi078), .ZN(new_n1126_));
  AOI21_X1   g836(.A1(new_n1126_), .A2(new_n1125_), .B(new_n1008_), .ZN(new_n1127_));
  NAND2_X1   g837(.A1(new_n742_), .A2(new_n943_), .ZN(new_n1128_));
  NAND2_X1   g838(.A1(new_n951_), .A2(pi136), .ZN(new_n1129_));
  AOI21_X1   g839(.A1(new_n1128_), .A2(new_n1129_), .B(pi137), .ZN(new_n1130_));
  OAI21_X1   g840(.A1(new_n1130_), .A2(new_n1127_), .B(new_n1029_), .ZN(new_n1131_));
  OAI21_X1   g841(.A1(new_n1029_), .A2(new_n1124_), .B(new_n1131_), .ZN(po118));
  INV_X1     g842(.I(pi112), .ZN(new_n1133_));
  AOI22_X1   g843(.A1(pi099), .A2(new_n944_), .B1(new_n1009_), .B2(new_n1133_), .ZN(new_n1134_));
  NAND2_X1   g844(.A1(new_n763_), .A2(new_n943_), .ZN(new_n1135_));
  NAND2_X1   g845(.A1(new_n972_), .A2(pi136), .ZN(new_n1136_));
  AOI21_X1   g846(.A1(new_n1135_), .A2(new_n1136_), .B(pi137), .ZN(new_n1137_));
  NAND2_X1   g847(.A1(pi032), .A2(pi136), .ZN(new_n1138_));
  NAND2_X1   g848(.A1(new_n943_), .A2(pi084), .ZN(new_n1139_));
  AOI21_X1   g849(.A1(new_n1139_), .A2(new_n1138_), .B(new_n1008_), .ZN(new_n1140_));
  OAI21_X1   g850(.A1(new_n1137_), .A2(new_n1140_), .B(new_n1029_), .ZN(new_n1141_));
  OAI21_X1   g851(.A1(new_n1029_), .A2(new_n1134_), .B(new_n1141_), .ZN(po119));
  NAND2_X1   g852(.A1(pi100), .A2(pi138), .ZN(new_n1143_));
  NAND2_X1   g853(.A1(new_n1029_), .A2(pi080), .ZN(new_n1144_));
  AOI21_X1   g854(.A1(new_n1144_), .A2(new_n1143_), .B(pi136), .ZN(new_n1145_));
  NOR2_X1    g855(.A1(new_n1032_), .A2(new_n720_), .ZN(new_n1146_));
  OAI21_X1   g856(.A1(new_n1145_), .A2(new_n1146_), .B(pi137), .ZN(new_n1147_));
  NAND2_X1   g857(.A1(pi092), .A2(pi138), .ZN(new_n1148_));
  NAND2_X1   g858(.A1(new_n980_), .A2(new_n1029_), .ZN(new_n1149_));
  AOI21_X1   g859(.A1(new_n1149_), .A2(new_n1148_), .B(new_n943_), .ZN(new_n1150_));
  NAND2_X1   g860(.A1(pi125), .A2(pi138), .ZN(new_n1151_));
  NAND2_X1   g861(.A1(new_n996_), .A2(new_n1029_), .ZN(new_n1152_));
  AOI21_X1   g862(.A1(new_n1152_), .A2(new_n1151_), .B(pi136), .ZN(new_n1153_));
  OAI21_X1   g863(.A1(new_n1150_), .A2(new_n1153_), .B(new_n1008_), .ZN(new_n1154_));
  NAND2_X1   g864(.A1(new_n1154_), .A2(new_n1147_), .ZN(po120));
  NAND4_X1   g865(.A1(new_n1046_), .A2(new_n581_), .A3(new_n591_), .A4(new_n636_), .ZN(new_n1156_));
  AOI21_X1   g866(.A1(new_n1156_), .A2(new_n617_), .B(new_n413_), .ZN(po121));
  NAND2_X1   g867(.A1(pi097), .A2(pi138), .ZN(new_n1158_));
  NAND2_X1   g868(.A1(new_n1029_), .A2(pi081), .ZN(new_n1159_));
  AOI21_X1   g869(.A1(new_n1159_), .A2(new_n1158_), .B(pi136), .ZN(new_n1160_));
  NOR2_X1    g870(.A1(new_n1032_), .A2(new_n726_), .ZN(new_n1161_));
  OAI21_X1   g871(.A1(new_n1160_), .A2(new_n1161_), .B(pi137), .ZN(new_n1162_));
  NAND2_X1   g872(.A1(pi098), .A2(pi138), .ZN(new_n1163_));
  NAND2_X1   g873(.A1(new_n984_), .A2(new_n1029_), .ZN(new_n1164_));
  AOI21_X1   g874(.A1(new_n1164_), .A2(new_n1163_), .B(new_n943_), .ZN(new_n1165_));
  NAND2_X1   g875(.A1(new_n1000_), .A2(new_n1029_), .ZN(new_n1166_));
  NAND2_X1   g876(.A1(pi023), .A2(pi138), .ZN(new_n1167_));
  AOI21_X1   g877(.A1(new_n1166_), .A2(new_n1167_), .B(pi136), .ZN(new_n1168_));
  OAI21_X1   g878(.A1(new_n1165_), .A2(new_n1168_), .B(new_n1008_), .ZN(new_n1169_));
  NAND2_X1   g879(.A1(new_n1169_), .A2(new_n1162_), .ZN(po122));
  NAND2_X1   g880(.A1(pi111), .A2(pi138), .ZN(new_n1171_));
  NAND2_X1   g881(.A1(new_n1029_), .A2(pi086), .ZN(new_n1172_));
  AOI21_X1   g882(.A1(new_n1172_), .A2(new_n1171_), .B(pi136), .ZN(new_n1173_));
  NOR2_X1    g883(.A1(new_n1032_), .A2(new_n690_), .ZN(new_n1174_));
  OAI21_X1   g884(.A1(new_n1173_), .A2(new_n1174_), .B(pi137), .ZN(new_n1175_));
  NAND2_X1   g885(.A1(pi088), .A2(pi138), .ZN(new_n1176_));
  NAND2_X1   g886(.A1(new_n834_), .A2(new_n1029_), .ZN(new_n1177_));
  AOI21_X1   g887(.A1(new_n1177_), .A2(new_n1176_), .B(new_n943_), .ZN(new_n1178_));
  NAND2_X1   g888(.A1(pi120), .A2(pi138), .ZN(new_n1179_));
  NAND2_X1   g889(.A1(new_n967_), .A2(new_n1029_), .ZN(new_n1180_));
  AOI21_X1   g890(.A1(new_n1180_), .A2(new_n1179_), .B(pi136), .ZN(new_n1181_));
  OAI21_X1   g891(.A1(new_n1178_), .A2(new_n1181_), .B(new_n1008_), .ZN(new_n1182_));
  NAND2_X1   g892(.A1(new_n1182_), .A2(new_n1175_), .ZN(po123));
  NAND2_X1   g893(.A1(new_n327_), .A2(pi116), .ZN(new_n1184_));
  OR2_X2     g894(.A1(new_n647_), .A2(new_n608_), .Z(new_n1185_));
  AOI21_X1   g895(.A1(new_n1185_), .A2(new_n648_), .B(new_n1184_), .ZN(po124));
  NAND2_X1   g896(.A1(new_n584_), .A2(new_n670_), .ZN(new_n1187_));
  AOI21_X1   g897(.A1(new_n1187_), .A2(new_n679_), .B(new_n1184_), .ZN(po125));
  NAND2_X1   g898(.A1(new_n1077_), .A2(new_n558_), .ZN(new_n1189_));
  NOR3_X1    g899(.A1(new_n364_), .A2(new_n1029_), .A3(pi137), .ZN(new_n1190_));
  NAND3_X1   g900(.A1(new_n1190_), .A2(new_n943_), .A3(pi139), .ZN(new_n1191_));
  INV_X1     g901(.I(new_n1084_), .ZN(new_n1192_));
  NAND2_X1   g902(.A1(new_n1192_), .A2(pi111), .ZN(new_n1193_));
  AOI21_X1   g903(.A1(new_n1193_), .A2(new_n1191_), .B(new_n1189_), .ZN(po126));
  NAND3_X1   g904(.A1(new_n1190_), .A2(new_n943_), .A3(pi141), .ZN(new_n1195_));
  NAND2_X1   g905(.A1(new_n1192_), .A2(new_n1133_), .ZN(new_n1196_));
  AOI21_X1   g906(.A1(new_n1196_), .A2(new_n1195_), .B(new_n1189_), .ZN(po127));
  NAND2_X1   g907(.A1(new_n306_), .A2(new_n403_), .ZN(new_n1198_));
  OAI21_X1   g908(.A1(pi011), .A2(pi022), .B(pi054), .ZN(new_n1199_));
  AOI21_X1   g909(.A1(new_n1198_), .A2(new_n1199_), .B(new_n413_), .ZN(po128));
  NAND3_X1   g910(.A1(new_n1190_), .A2(new_n943_), .A3(pi140), .ZN(new_n1201_));
  NAND2_X1   g911(.A1(new_n1192_), .A2(new_n1027_), .ZN(new_n1202_));
  AOI21_X1   g912(.A1(new_n1202_), .A2(new_n1201_), .B(new_n1189_), .ZN(po130));
  NOR4_X1    g913(.A1(pi004), .A2(pi007), .A3(pi009), .A4(pi012), .ZN(new_n1204_));
  NOR3_X1    g914(.A1(new_n413_), .A2(new_n1204_), .A3(new_n306_), .ZN(po131));
  NAND2_X1   g915(.A1(new_n558_), .A2(pi122), .ZN(po132));
  NAND2_X1   g916(.A1(new_n306_), .A2(pi118), .ZN(new_n1207_));
  NAND3_X1   g917(.A1(new_n479_), .A2(pi054), .A3(new_n419_), .ZN(new_n1208_));
  AOI21_X1   g918(.A1(new_n1208_), .A2(new_n1207_), .B(pi129), .ZN(po133));
  AOI21_X1   g919(.A1(new_n630_), .A2(new_n629_), .B(pi129), .ZN(po134));
  NOR3_X1    g920(.A1(pi003), .A2(pi110), .A3(pi120), .ZN(new_n1211_));
  NOR3_X1    g921(.A1(new_n1211_), .A2(pi111), .A3(pi129), .ZN(po135));
  AND3_X2    g922(.A1(new_n558_), .A2(pi081), .A3(pi120), .Z(po136));
  OR2_X2     g923(.A1(pi129), .A2(pi134), .Z(po137));
  OR2_X2     g924(.A1(pi129), .A2(pi135), .Z(po138));
  NOR2_X1    g925(.A1(new_n912_), .A2(pi129), .ZN(po139));
  NAND2_X1   g926(.A1(new_n620_), .A2(pi125), .ZN(new_n1217_));
  AOI21_X1   g927(.A1(new_n1217_), .A2(new_n1085_), .B(pi129), .ZN(po140));
  INV_X1     g928(.I(pi126), .ZN(new_n1219_));
  AND3_X2    g929(.A1(new_n1219_), .A2(pi132), .A3(pi133), .Z(po141));
  assign     po012 = 1'b1;
  BUF_X16    g930(.I(pi108), .Z(po000));
  BUF_X16    g931(.I(pi083), .Z(po001));
  BUF_X16    g932(.I(pi104), .Z(po002));
  BUF_X16    g933(.I(pi103), .Z(po003));
  BUF_X16    g934(.I(pi102), .Z(po004));
  BUF_X16    g935(.I(pi105), .Z(po005));
  BUF_X16    g936(.I(pi107), .Z(po006));
  BUF_X16    g937(.I(pi101), .Z(po007));
  BUF_X16    g938(.I(pi126), .Z(po008));
  BUF_X16    g939(.I(pi121), .Z(po009));
  BUF_X16    g940(.I(pi001), .Z(po010));
  BUF_X16    g941(.I(pi000), .Z(po011));
  BUF_X16    g942(.I(pi130), .Z(po013));
  BUF_X16    g943(.I(pi128), .Z(po014));
endmodule


