module top(a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_, a_31_, a_32_, a_33_, a_34_, a_35_, a_36_, a_37_, a_38_, a_39_, a_40_, a_41_, a_42_, a_43_, a_44_, a_45_, a_46_, a_47_, a_48_, a_49_, a_50_, a_51_, a_52_, a_53_, a_54_, a_55_, a_56_, a_57_, a_58_, a_59_, a_60_, a_61_, a_62_, a_63_, a_64_, a_65_, a_66_, a_67_, a_68_, a_69_, a_70_, a_71_, a_72_, a_73_, a_74_, a_75_, a_76_, a_77_, a_78_, a_79_, a_80_, a_81_, a_82_, a_83_, a_84_, a_85_, a_86_, a_87_, a_88_, a_89_, a_90_, a_91_, a_92_, a_93_, a_94_, a_95_, a_96_, a_97_, a_98_, a_99_, a_100_, a_101_, a_102_, a_103_, a_104_, a_105_, a_106_, a_107_, a_108_, a_109_, a_110_, a_111_, a_112_, a_113_, a_114_, a_115_, a_116_, a_117_, a_118_, a_119_, a_120_, a_121_, a_122_, a_123_, a_124_, a_125_, a_126_, a_127_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_, b_30_, b_31_, b_32_, b_33_, b_34_, b_35_, b_36_, b_37_, b_38_, b_39_, b_40_, b_41_, b_42_, b_43_, b_44_, b_45_, b_46_, b_47_, b_48_, b_49_, b_50_, b_51_, b_52_, b_53_, b_54_, b_55_, b_56_, b_57_, b_58_, b_59_, b_60_, b_61_, b_62_, b_63_, b_64_, b_65_, b_66_, b_67_, b_68_, b_69_, b_70_, b_71_, b_72_, b_73_, b_74_, b_75_, b_76_, b_77_, b_78_, b_79_, b_80_, b_81_, b_82_, b_83_, b_84_, b_85_, b_86_, b_87_, b_88_, b_89_, b_90_, b_91_, b_92_, b_93_, b_94_, b_95_, b_96_, b_97_, b_98_, b_99_, b_100_, b_101_, b_102_, b_103_, b_104_, b_105_, b_106_, b_107_, b_108_, b_109_, b_110_, b_111_, b_112_, b_113_, b_114_, b_115_, b_116_, b_117_, b_118_, b_119_, b_120_, b_121_, b_122_, b_123_, b_124_, b_125_, b_126_, b_127_, f_0_, f_1_, f_2_, f_3_, f_4_, f_5_, f_6_, f_7_, f_8_, f_9_, f_10_, f_11_, f_12_, f_13_, f_14_, f_15_, f_16_, f_17_, f_18_, f_19_, f_20_, f_21_, f_22_, f_23_, f_24_, f_25_, f_26_, f_27_, f_28_, f_29_, f_30_, f_31_, f_32_, f_33_, f_34_, f_35_, f_36_, f_37_, f_38_, f_39_, f_40_, f_41_, f_42_, f_43_, f_44_, f_45_, f_46_, f_47_, f_48_, f_49_, f_50_, f_51_, f_52_, f_53_, f_54_, f_55_, f_56_, f_57_, f_58_, f_59_, f_60_, f_61_, f_62_, f_63_, f_64_, f_65_, f_66_, f_67_, f_68_, f_69_, f_70_, f_71_, f_72_, f_73_, f_74_, f_75_, f_76_, f_77_, f_78_, f_79_, f_80_, f_81_, f_82_, f_83_, f_84_, f_85_, f_86_, f_87_, f_88_, f_89_, f_90_, f_91_, f_92_, f_93_, f_94_, f_95_, f_96_, f_97_, f_98_, f_99_, f_100_, f_101_, f_102_, f_103_, f_104_, f_105_, f_106_, f_107_, f_108_, f_109_, f_110_, f_111_, f_112_, f_113_, f_114_, f_115_, f_116_, f_117_, f_118_, f_119_, f_120_, f_121_, f_122_, f_123_, f_124_, f_125_, f_126_, f_127_, cOut);
  wire n392;
  wire n391;
  wire n396;
  wire n400;
  wire n399;
  wire n404;
  wire n408;
  wire n407;
  wire n412;
  wire n416;
  wire n415;
  wire n420;
  wire n424;
  wire n423;
  wire n428;
  wire n432;
  wire n431;
  wire n436;
  wire n440;
  wire n439;
  wire n444;
  wire n448;
  wire n447;
  wire n452;
  wire n456;
  wire n455;
  wire n460;
  wire n464;
  wire n463;
  wire n468;
  wire n472;
  wire n471;
  wire n476;
  wire n480;
  wire n479;
  wire n484;
  wire n488;
  wire n487;
  wire n492;
  wire n496;
  wire n495;
  wire n500;
  wire n504;
  wire n503;
  wire n508;
  wire n512;
  wire n511;
  wire n516;
  wire n520;
  wire n519;
  wire n524;
  wire n528;
  wire n527;
  wire n532;
  wire n536;
  wire n535;
  wire n540;
  wire n544;
  wire n543;
  wire n548;
  wire n552;
  wire n551;
  wire n556;
  wire n560;
  wire n559;
  wire n564;
  wire n568;
  wire n567;
  wire n572;
  wire n576;
  wire n575;
  wire n580;
  wire n584;
  wire n583;
  wire n588;
  wire n592;
  wire n591;
  wire n596;
  wire n600;
  wire n599;
  wire n604;
  wire n608;
  wire n607;
  wire n612;
  wire n616;
  wire n615;
  wire n620;
  wire n624;
  wire n623;
  wire n628;
  wire n632;
  wire n631;
  wire n636;
  wire n640;
  wire n639;
  wire n644;
  wire n648;
  wire n647;
  wire n652;
  wire n656;
  wire n655;
  wire n660;
  wire n664;
  wire n663;
  wire n668;
  wire n672;
  wire n671;
  wire n676;
  wire n680;
  wire n679;
  wire n684;
  wire n688;
  wire n687;
  wire n692;
  wire n696;
  wire n695;
  wire n700;
  wire n704;
  wire n703;
  wire n708;
  wire n712;
  wire n711;
  wire n716;
  wire n720;
  wire n719;
  wire n724;
  wire n728;
  wire n727;
  wire n732;
  wire n736;
  wire n735;
  wire n740;
  wire n744;
  wire n743;
  wire n748;
  wire n752;
  wire n751;
  wire n756;
  wire n760;
  wire n759;
  wire n764;
  wire n768;
  wire n767;
  wire n772;
  wire n776;
  wire n775;
  wire n780;
  wire n784;
  wire n783;
  wire n788;
  wire n792;
  wire n791;
  wire n796;
  wire n800;
  wire n799;
  wire n804;
  wire n808;
  wire n807;
  wire n812;
  wire n816;
  wire n815;
  wire n820;
  wire n824;
  wire n823;
  wire n828;
  wire n832;
  wire n831;
  wire n836;
  wire n840;
  wire n839;
  wire n844;
  wire n848;
  wire n847;
  wire n852;
  wire n856;
  wire n855;
  wire n860;
  wire n864;
  wire n863;
  wire n868;
  wire n872;
  wire n871;
  wire n876;
  wire n880;
  wire n879;
  wire n884;
  wire n888;
  wire n887;
  wire n892;
  wire n896;
  wire n895;
  wire n900;
  wire n904;
  wire n903;
  wire n908;
  wire n912;
  wire n911;
  wire n916;
  wire n920;
  wire n919;
  wire n924;
  wire n928;
  wire n927;
  wire n932;
  wire n936;
  wire n935;
  wire n940;
  wire n944;
  wire n943;
  wire n948;
  wire n952;
  wire n951;
  wire n956;
  wire n960;
  wire n959;
  wire n964;
  wire n968;
  wire n967;
  wire n972;
  wire n976;
  wire n975;
  wire n980;
  wire n984;
  wire n983;
  wire n988;
  wire n992;
  wire n1000;
  wire n991;
  wire n996;
  wire n1004;
  wire n1008;
  wire n999;
  wire n1007;
  wire n1012;
  wire n1016;
  wire n1015;
  wire n1020;
  wire n1024;
  wire n1023;
  wire n1028;
  wire n1032;
  wire n1031;
  wire n1036;
  wire n1040;
  wire n1039;
  wire n1044;
  wire n1048;
  wire n1047;
  wire n1052;
  wire n1056;
  wire n1055;
  wire n1060;
  wire n1064;
  wire n1063;
  wire n1068;
  wire n1072;
  wire n1071;
  wire n1076;
  wire n1080;
  wire n1079;
  wire n1084;
  wire n1088;
  wire n1087;
  wire n1092;
  wire n1096;
  wire n1095;
  wire n1100;
  wire n1104;
  wire n1103;
  wire n1108;
  wire n1112;
  wire n1111;
  wire n1116;
  wire n1120;
  wire n1119;
  wire n1124;
  wire n1128;
  wire n1127;
  wire n1132;
  wire n1136;
  wire n1135;
  wire n1140;
  wire n1144;
  wire n1143;
  wire n1148;
  wire n1152;
  wire n1151;
  wire n1156;
  wire n1160;
  wire n1159;
  wire n1164;
  wire n1168;
  wire n1167;
  wire n1172;
  wire n1176;
  wire n1175;
  wire n1180;
  wire n1184;
  wire n1183;
  wire n1188;
  wire n1192;
  wire n1191;
  wire n1196;
  wire n1200;
  wire n1199;
  wire n1204;
  wire n1208;
  wire n1207;
  wire n1212;
  wire n1216;
  wire n1215;
  wire n1220;
  wire n1224;
  wire n1223;
  wire n1228;
  wire n1232;
  wire n1231;
  wire n1236;
  wire n1240;
  wire n1239;
  wire n1244;
  wire n1248;
  wire n1247;
  wire n1252;
  wire n1256;
  wire n1255;
  wire n1260;
  wire n1264;
  wire n1263;
  wire n1268;
  wire n1272;
  wire n1271;
  wire n1276;
  wire n1280;
  wire n1279;
  wire n1284;
  wire n1288;
  wire n1287;
  wire n1292;
  wire n1296;
  wire n1295;
  wire n1300;
  wire n1304;
  wire n1303;
  wire n1308;
  wire n1312;
  wire n1311;
  wire n1316;
  wire n1320;
  wire n1319;
  wire n1324;
  wire n1328;
  wire n1327;
  wire n1332;
  wire n1336;
  wire n1335;
  wire n1340;
  wire n1344;
  wire n1343;
  wire n1348;
  wire n1352;
  wire n1351;
  wire n1356;
  wire n1360;
  wire n1359;
  wire n1364;
  wire n1368;
  wire n1367;
  wire n1372;
  wire n1376;
  wire n1375;
  wire n1380;
  wire n1384;
  wire n1383;
  wire n1388;
  wire n1392;
  wire n1391;
  wire n1396;
  wire n1400;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n390;
  wire n1389;
  wire n1390;
  wire n1381;
  wire n1382;
  wire n1373;
  wire n1374;
  wire n1365;
  wire n1366;
  wire n1357;
  wire n1358;
  wire n1349;
  wire n1350;
  wire n1341;
  wire n1342;
  wire n1333;
  wire n1334;
  wire n1325;
  wire n1326;
  wire n1317;
  wire n1318;
  wire n1309;
  wire n1310;
  wire n1301;
  wire n1302;
  wire n1293;
  wire n1294;
  wire n1285;
  wire n1286;
  wire n1277;
  wire n1278;
  wire n1269;
  wire n1270;
  wire n1261;
  wire n1262;
  wire n1253;
  wire n1254;
  wire n1245;
  wire n1246;
  wire n1237;
  wire n1238;
  wire n1229;
  wire n1230;
  wire n1221;
  wire n1222;
  wire n1213;
  wire n1214;
  wire n1205;
  wire n1206;
  wire n1197;
  wire n1198;
  wire n1189;
  wire n1190;
  wire n1181;
  wire n1182;
  wire n1173;
  wire n1174;
  wire n1165;
  wire n1166;
  wire n1157;
  wire n1158;
  wire n1149;
  wire n1150;
  wire n1141;
  wire n1142;
  wire n1133;
  wire n1134;
  wire n1125;
  wire n1126;
  wire n1117;
  wire n1118;
  wire n1109;
  wire n1110;
  wire n1101;
  wire n1102;
  wire n1093;
  wire n1094;
  wire n1085;
  wire n1086;
  wire n1077;
  wire n1078;
  wire n1069;
  wire n1070;
  wire n1061;
  wire n1062;
  wire n1053;
  wire n1054;
  wire n1045;
  wire n1046;
  wire n1037;
  wire n1038;
  wire n1029;
  wire n1030;
  wire n1021;
  wire n1022;
  wire n1013;
  wire n1014;
  wire n1005;
  wire n1006;
  wire n997;
  wire n998;
  wire n989;
  wire n990;
  wire n981;
  wire n982;
  wire n973;
  wire n974;
  wire n965;
  wire n966;
  wire n957;
  wire n958;
  wire n949;
  wire n950;
  wire n941;
  wire n942;
  wire n933;
  wire n934;
  wire n925;
  wire n926;
  wire n917;
  wire n918;
  wire n909;
  wire n910;
  wire n901;
  wire n902;
  wire n893;
  wire n894;
  wire n885;
  wire n886;
  wire n877;
  wire n878;
  wire n869;
  wire n870;
  wire n861;
  wire n862;
  wire n853;
  wire n854;
  wire n845;
  wire n846;
  wire n837;
  wire n838;
  wire n829;
  wire n830;
  wire n821;
  wire n822;
  wire n813;
  wire n814;
  wire n805;
  wire n806;
  wire n797;
  wire n798;
  wire n789;
  wire n790;
  wire n781;
  wire n782;
  wire n773;
  wire n774;
  wire n765;
  wire n766;
  wire n757;
  wire n758;
  wire n749;
  wire n750;
  wire n741;
  wire n742;
  wire n733;
  wire n734;
  wire n725;
  wire n726;
  wire n717;
  wire n718;
  wire n709;
  wire n710;
  wire n701;
  wire n702;
  wire n693;
  wire n694;
  wire n685;
  wire n686;
  wire n677;
  wire n678;
  wire n669;
  wire n670;
  wire n661;
  wire n662;
  wire n653;
  wire n654;
  wire n645;
  wire n646;
  wire n637;
  wire n638;
  wire n629;
  wire n630;
  wire n621;
  wire n622;
  wire n613;
  wire n614;
  wire n605;
  wire n606;
  wire n597;
  wire n598;
  wire n589;
  wire n590;
  wire n581;
  wire n582;
  wire n573;
  wire n574;
  wire n565;
  wire n566;
  wire n557;
  wire n558;
  wire n549;
  wire n550;
  wire n541;
  wire n542;
  wire n533;
  wire n534;
  wire n525;
  wire n526;
  wire n517;
  wire n518;
  wire n509;
  wire n510;
  wire n501;
  wire n502;
  wire n493;
  wire n494;
  wire n485;
  wire n486;
  wire n477;
  wire n478;
  wire n469;
  wire n470;
  wire n461;
  wire n462;
  wire n453;
  wire n454;
  wire n445;
  wire n446;
  wire n437;
  wire n438;
  wire n429;
  wire n430;
  wire n421;
  wire n422;
  wire n413;
  wire n414;
  wire n405;
  wire n406;
  wire n397;
  wire n398;
  wire n389;
  input a_0_;
  input a_1_;
  input a_2_;
  input a_3_;
  input a_4_;
  input a_5_;
  input a_6_;
  input a_7_;
  input a_8_;
  input a_9_;
  input a_10_;
  input a_11_;
  input a_12_;
  input a_13_;
  input a_14_;
  input a_15_;
  input a_16_;
  input a_17_;
  input a_18_;
  input a_19_;
  input a_20_;
  input a_21_;
  input a_22_;
  input a_23_;
  input a_24_;
  input a_25_;
  input a_26_;
  input a_27_;
  input a_28_;
  input a_29_;
  input a_30_;
  input a_31_;
  input a_32_;
  input a_33_;
  input a_34_;
  input a_35_;
  input a_36_;
  input a_37_;
  input a_38_;
  input a_39_;
  input a_40_;
  input a_41_;
  input a_42_;
  input a_43_;
  input a_44_;
  input a_45_;
  input a_46_;
  input a_47_;
  input a_48_;
  input a_49_;
  input a_50_;
  input a_51_;
  input a_52_;
  input a_53_;
  input a_54_;
  input a_55_;
  input a_56_;
  input a_57_;
  input a_58_;
  input a_59_;
  input a_60_;
  input a_61_;
  input a_62_;
  input a_63_;
  input a_64_;
  input a_65_;
  input a_66_;
  input a_67_;
  input a_68_;
  input a_69_;
  input a_70_;
  input a_71_;
  input a_72_;
  input a_73_;
  input a_74_;
  input a_75_;
  input a_76_;
  input a_77_;
  input a_78_;
  input a_79_;
  input a_80_;
  input a_81_;
  input a_82_;
  input a_83_;
  input a_84_;
  input a_85_;
  input a_86_;
  input a_87_;
  input a_88_;
  input a_89_;
  input a_90_;
  input a_91_;
  input a_92_;
  input a_93_;
  input a_94_;
  input a_95_;
  input a_96_;
  input a_97_;
  input a_98_;
  input a_99_;
  input a_100_;
  input a_101_;
  input a_102_;
  input a_103_;
  input a_104_;
  input a_105_;
  input a_106_;
  input a_107_;
  input a_108_;
  input a_109_;
  input a_110_;
  input a_111_;
  input a_112_;
  input a_113_;
  input a_114_;
  input a_115_;
  input a_116_;
  input a_117_;
  input a_118_;
  input a_119_;
  input a_120_;
  input a_121_;
  input a_122_;
  input a_123_;
  input a_124_;
  input a_125_;
  input a_126_;
  input a_127_;
  input b_0_;
  input b_1_;
  input b_2_;
  input b_3_;
  input b_4_;
  input b_5_;
  input b_6_;
  input b_7_;
  input b_8_;
  input b_9_;
  input b_10_;
  input b_11_;
  input b_12_;
  input b_13_;
  input b_14_;
  input b_15_;
  input b_16_;
  input b_17_;
  input b_18_;
  input b_19_;
  input b_20_;
  input b_21_;
  input b_22_;
  input b_23_;
  input b_24_;
  input b_25_;
  input b_26_;
  input b_27_;
  input b_28_;
  input b_29_;
  input b_30_;
  input b_31_;
  input b_32_;
  input b_33_;
  input b_34_;
  input b_35_;
  input b_36_;
  input b_37_;
  input b_38_;
  input b_39_;
  input b_40_;
  input b_41_;
  input b_42_;
  input b_43_;
  input b_44_;
  input b_45_;
  input b_46_;
  input b_47_;
  input b_48_;
  input b_49_;
  input b_50_;
  input b_51_;
  input b_52_;
  input b_53_;
  input b_54_;
  input b_55_;
  input b_56_;
  input b_57_;
  input b_58_;
  input b_59_;
  input b_60_;
  input b_61_;
  input b_62_;
  input b_63_;
  input b_64_;
  input b_65_;
  input b_66_;
  input b_67_;
  input b_68_;
  input b_69_;
  input b_70_;
  input b_71_;
  input b_72_;
  input b_73_;
  input b_74_;
  input b_75_;
  input b_76_;
  input b_77_;
  input b_78_;
  input b_79_;
  input b_80_;
  input b_81_;
  input b_82_;
  input b_83_;
  input b_84_;
  input b_85_;
  input b_86_;
  input b_87_;
  input b_88_;
  input b_89_;
  input b_90_;
  input b_91_;
  input b_92_;
  input b_93_;
  input b_94_;
  input b_95_;
  input b_96_;
  input b_97_;
  input b_98_;
  input b_99_;
  input b_100_;
  input b_101_;
  input b_102_;
  input b_103_;
  input b_104_;
  input b_105_;
  input b_106_;
  input b_107_;
  input b_108_;
  input b_109_;
  input b_110_;
  input b_111_;
  input b_112_;
  input b_113_;
  input b_114_;
  input b_115_;
  input b_116_;
  input b_117_;
  input b_118_;
  input b_119_;
  input b_120_;
  input b_121_;
  input b_122_;
  input b_123_;
  input b_124_;
  input b_125_;
  input b_126_;
  input b_127_;
  output f_0_;
  output f_1_;
  output f_2_;
  output f_3_;
  output f_4_;
  output f_5_;
  output f_6_;
  output f_7_;
  output f_8_;
  output f_9_;
  output f_10_;
  output f_11_;
  output f_12_;
  output f_13_;
  output f_14_;
  output f_15_;
  output f_16_;
  output f_17_;
  output f_18_;
  output f_19_;
  output f_20_;
  output f_21_;
  output f_22_;
  output f_23_;
  output f_24_;
  output f_25_;
  output f_26_;
  output f_27_;
  output f_28_;
  output f_29_;
  output f_30_;
  output f_31_;
  output f_32_;
  output f_33_;
  output f_34_;
  output f_35_;
  output f_36_;
  output f_37_;
  output f_38_;
  output f_39_;
  output f_40_;
  output f_41_;
  output f_42_;
  output f_43_;
  output f_44_;
  output f_45_;
  output f_46_;
  output f_47_;
  output f_48_;
  output f_49_;
  output f_50_;
  output f_51_;
  output f_52_;
  output f_53_;
  output f_54_;
  output f_55_;
  output f_56_;
  output f_57_;
  output f_58_;
  output f_59_;
  output f_60_;
  output f_61_;
  output f_62_;
  output f_63_;
  output f_64_;
  output f_65_;
  output f_66_;
  output f_67_;
  output f_68_;
  output f_69_;
  output f_70_;
  output f_71_;
  output f_72_;
  output f_73_;
  output f_74_;
  output f_75_;
  output f_76_;
  output f_77_;
  output f_78_;
  output f_79_;
  output f_80_;
  output f_81_;
  output f_82_;
  output f_83_;
  output f_84_;
  output f_85_;
  output f_86_;
  output f_87_;
  output f_88_;
  output f_89_;
  output f_90_;
  output f_91_;
  output f_92_;
  output f_93_;
  output f_94_;
  output f_95_;
  output f_96_;
  output f_97_;
  output f_98_;
  output f_99_;
  output f_100_;
  output f_101_;
  output f_102_;
  output f_103_;
  output f_104_;
  output f_105_;
  output f_106_;
  output f_107_;
  output f_108_;
  output f_109_;
  output f_110_;
  output f_111_;
  output f_112_;
  output f_113_;
  output f_114_;
  output f_115_;
  output f_116_;
  output f_117_;
  output f_118_;
  output f_119_;
  output f_120_;
  output f_121_;
  output f_122_;
  output f_123_;
  output f_124_;
  output f_125_;
  output f_126_;
  output f_127_;
  output cOut;
  AND2_X2 n_n0 (
    .A1(a_0_),
    .A2(b_0_),
    .Z(f_0_)
  );
  OAI21_X1 n_n1 (
    .A1(a_0_),
    .A2(b_0_),
    .B(n392),
    .ZN(f_1_)
  );
  AOI21_X1 n_n2 (
    .A1(n391),
    .A2(n396),
    .B(n400),
    .ZN(f_2_)
  );
  AOI21_X1 n_n3 (
    .A1(n399),
    .A2(n404),
    .B(n408),
    .ZN(f_3_)
  );
  AOI21_X1 n_n4 (
    .A1(n407),
    .A2(n412),
    .B(n416),
    .ZN(f_4_)
  );
  AOI21_X1 n_n5 (
    .A1(n415),
    .A2(n420),
    .B(n424),
    .ZN(f_5_)
  );
  AOI21_X1 n_n6 (
    .A1(n423),
    .A2(n428),
    .B(n432),
    .ZN(f_6_)
  );
  AOI21_X1 n_n7 (
    .A1(n431),
    .A2(n436),
    .B(n440),
    .ZN(f_7_)
  );
  AOI21_X1 n_n8 (
    .A1(n439),
    .A2(n444),
    .B(n448),
    .ZN(f_8_)
  );
  AOI21_X1 n_n9 (
    .A1(n447),
    .A2(n452),
    .B(n456),
    .ZN(f_9_)
  );
  AOI21_X1 n_n10 (
    .A1(n455),
    .A2(n460),
    .B(n464),
    .ZN(f_10_)
  );
  AOI21_X1 n_n11 (
    .A1(n463),
    .A2(n468),
    .B(n472),
    .ZN(f_11_)
  );
  AOI21_X1 n_n12 (
    .A1(n471),
    .A2(n476),
    .B(n480),
    .ZN(f_12_)
  );
  AOI21_X1 n_n13 (
    .A1(n479),
    .A2(n484),
    .B(n488),
    .ZN(f_13_)
  );
  AOI21_X1 n_n14 (
    .A1(n487),
    .A2(n492),
    .B(n496),
    .ZN(f_14_)
  );
  AOI21_X1 n_n15 (
    .A1(n495),
    .A2(n500),
    .B(n504),
    .ZN(f_15_)
  );
  AOI21_X1 n_n16 (
    .A1(n503),
    .A2(n508),
    .B(n512),
    .ZN(f_16_)
  );
  AOI21_X1 n_n17 (
    .A1(n511),
    .A2(n516),
    .B(n520),
    .ZN(f_17_)
  );
  AOI21_X1 n_n18 (
    .A1(n519),
    .A2(n524),
    .B(n528),
    .ZN(f_18_)
  );
  AOI21_X1 n_n19 (
    .A1(n527),
    .A2(n532),
    .B(n536),
    .ZN(f_19_)
  );
  AOI21_X1 n_n20 (
    .A1(n535),
    .A2(n540),
    .B(n544),
    .ZN(f_20_)
  );
  AOI21_X1 n_n21 (
    .A1(n543),
    .A2(n548),
    .B(n552),
    .ZN(f_21_)
  );
  AOI21_X1 n_n22 (
    .A1(n551),
    .A2(n556),
    .B(n560),
    .ZN(f_22_)
  );
  AOI21_X1 n_n23 (
    .A1(n559),
    .A2(n564),
    .B(n568),
    .ZN(f_23_)
  );
  AOI21_X1 n_n24 (
    .A1(n567),
    .A2(n572),
    .B(n576),
    .ZN(f_24_)
  );
  AOI21_X1 n_n25 (
    .A1(n575),
    .A2(n580),
    .B(n584),
    .ZN(f_25_)
  );
  AOI21_X1 n_n26 (
    .A1(n583),
    .A2(n588),
    .B(n592),
    .ZN(f_26_)
  );
  AOI21_X1 n_n27 (
    .A1(n591),
    .A2(n596),
    .B(n600),
    .ZN(f_27_)
  );
  AOI21_X1 n_n28 (
    .A1(n599),
    .A2(n604),
    .B(n608),
    .ZN(f_28_)
  );
  AOI21_X1 n_n29 (
    .A1(n607),
    .A2(n612),
    .B(n616),
    .ZN(f_29_)
  );
  AOI21_X1 n_n30 (
    .A1(n615),
    .A2(n620),
    .B(n624),
    .ZN(f_30_)
  );
  AOI21_X1 n_n31 (
    .A1(n623),
    .A2(n628),
    .B(n632),
    .ZN(f_31_)
  );
  AOI21_X1 n_n32 (
    .A1(n631),
    .A2(n636),
    .B(n640),
    .ZN(f_32_)
  );
  AOI21_X1 n_n33 (
    .A1(n639),
    .A2(n644),
    .B(n648),
    .ZN(f_33_)
  );
  AOI21_X1 n_n34 (
    .A1(n647),
    .A2(n652),
    .B(n656),
    .ZN(f_34_)
  );
  AOI21_X1 n_n35 (
    .A1(n655),
    .A2(n660),
    .B(n664),
    .ZN(f_35_)
  );
  AOI21_X1 n_n36 (
    .A1(n663),
    .A2(n668),
    .B(n672),
    .ZN(f_36_)
  );
  AOI21_X1 n_n37 (
    .A1(n671),
    .A2(n676),
    .B(n680),
    .ZN(f_37_)
  );
  AOI21_X1 n_n38 (
    .A1(n679),
    .A2(n684),
    .B(n688),
    .ZN(f_38_)
  );
  AOI21_X1 n_n39 (
    .A1(n687),
    .A2(n692),
    .B(n696),
    .ZN(f_39_)
  );
  AOI21_X1 n_n40 (
    .A1(n695),
    .A2(n700),
    .B(n704),
    .ZN(f_40_)
  );
  AOI21_X1 n_n41 (
    .A1(n703),
    .A2(n708),
    .B(n712),
    .ZN(f_41_)
  );
  AOI21_X1 n_n42 (
    .A1(n711),
    .A2(n716),
    .B(n720),
    .ZN(f_42_)
  );
  AOI21_X1 n_n43 (
    .A1(n719),
    .A2(n724),
    .B(n728),
    .ZN(f_43_)
  );
  AOI21_X1 n_n44 (
    .A1(n727),
    .A2(n732),
    .B(n736),
    .ZN(f_44_)
  );
  AOI21_X1 n_n45 (
    .A1(n735),
    .A2(n740),
    .B(n744),
    .ZN(f_45_)
  );
  AOI21_X1 n_n46 (
    .A1(n743),
    .A2(n748),
    .B(n752),
    .ZN(f_46_)
  );
  AOI21_X1 n_n47 (
    .A1(n751),
    .A2(n756),
    .B(n760),
    .ZN(f_47_)
  );
  AOI21_X1 n_n48 (
    .A1(n759),
    .A2(n764),
    .B(n768),
    .ZN(f_48_)
  );
  AOI21_X1 n_n49 (
    .A1(n767),
    .A2(n772),
    .B(n776),
    .ZN(f_49_)
  );
  AOI21_X1 n_n50 (
    .A1(n775),
    .A2(n780),
    .B(n784),
    .ZN(f_50_)
  );
  AOI21_X1 n_n51 (
    .A1(n783),
    .A2(n788),
    .B(n792),
    .ZN(f_51_)
  );
  AOI21_X1 n_n52 (
    .A1(n791),
    .A2(n796),
    .B(n800),
    .ZN(f_52_)
  );
  AOI21_X1 n_n53 (
    .A1(n799),
    .A2(n804),
    .B(n808),
    .ZN(f_53_)
  );
  AOI21_X1 n_n54 (
    .A1(n807),
    .A2(n812),
    .B(n816),
    .ZN(f_54_)
  );
  AOI21_X1 n_n55 (
    .A1(n815),
    .A2(n820),
    .B(n824),
    .ZN(f_55_)
  );
  AOI21_X1 n_n56 (
    .A1(n823),
    .A2(n828),
    .B(n832),
    .ZN(f_56_)
  );
  AOI21_X1 n_n57 (
    .A1(n831),
    .A2(n836),
    .B(n840),
    .ZN(f_57_)
  );
  AOI21_X1 n_n58 (
    .A1(n839),
    .A2(n844),
    .B(n848),
    .ZN(f_58_)
  );
  AOI21_X1 n_n59 (
    .A1(n847),
    .A2(n852),
    .B(n856),
    .ZN(f_59_)
  );
  AOI21_X1 n_n60 (
    .A1(n855),
    .A2(n860),
    .B(n864),
    .ZN(f_60_)
  );
  AOI21_X1 n_n61 (
    .A1(n863),
    .A2(n868),
    .B(n872),
    .ZN(f_61_)
  );
  AOI21_X1 n_n62 (
    .A1(n871),
    .A2(n876),
    .B(n880),
    .ZN(f_62_)
  );
  AOI21_X1 n_n63 (
    .A1(n879),
    .A2(n884),
    .B(n888),
    .ZN(f_63_)
  );
  AOI21_X1 n_n64 (
    .A1(n887),
    .A2(n892),
    .B(n896),
    .ZN(f_64_)
  );
  AOI21_X1 n_n65 (
    .A1(n895),
    .A2(n900),
    .B(n904),
    .ZN(f_65_)
  );
  AOI21_X1 n_n66 (
    .A1(n903),
    .A2(n908),
    .B(n912),
    .ZN(f_66_)
  );
  AOI21_X1 n_n67 (
    .A1(n911),
    .A2(n916),
    .B(n920),
    .ZN(f_67_)
  );
  AOI21_X1 n_n68 (
    .A1(n919),
    .A2(n924),
    .B(n928),
    .ZN(f_68_)
  );
  AOI21_X1 n_n69 (
    .A1(n927),
    .A2(n932),
    .B(n936),
    .ZN(f_69_)
  );
  AOI21_X1 n_n70 (
    .A1(n935),
    .A2(n940),
    .B(n944),
    .ZN(f_70_)
  );
  AOI21_X1 n_n71 (
    .A1(n943),
    .A2(n948),
    .B(n952),
    .ZN(f_71_)
  );
  AOI21_X1 n_n72 (
    .A1(n951),
    .A2(n956),
    .B(n960),
    .ZN(f_72_)
  );
  AOI21_X1 n_n73 (
    .A1(n959),
    .A2(n964),
    .B(n968),
    .ZN(f_73_)
  );
  AOI21_X1 n_n74 (
    .A1(n967),
    .A2(n972),
    .B(n976),
    .ZN(f_74_)
  );
  AOI21_X1 n_n75 (
    .A1(n975),
    .A2(n980),
    .B(n984),
    .ZN(f_75_)
  );
  AOI21_X1 n_n76 (
    .A1(n983),
    .A2(n988),
    .B(n992),
    .ZN(f_76_)
  );
  OAI21_X1 n_n77 (
    .A1(n1000),
    .A2(n991),
    .B(n996),
    .ZN(f_77_)
  );
  OAI21_X1 n_n78 (
    .A1(n1004),
    .A2(n1008),
    .B(n999),
    .ZN(f_78_)
  );
  AOI21_X1 n_n79 (
    .A1(n1007),
    .A2(n1012),
    .B(n1016),
    .ZN(f_79_)
  );
  AOI21_X1 n_n80 (
    .A1(n1015),
    .A2(n1020),
    .B(n1024),
    .ZN(f_80_)
  );
  AOI21_X1 n_n81 (
    .A1(n1023),
    .A2(n1028),
    .B(n1032),
    .ZN(f_81_)
  );
  AOI21_X1 n_n82 (
    .A1(n1031),
    .A2(n1036),
    .B(n1040),
    .ZN(f_82_)
  );
  AOI21_X1 n_n83 (
    .A1(n1039),
    .A2(n1044),
    .B(n1048),
    .ZN(f_83_)
  );
  AOI21_X1 n_n84 (
    .A1(n1047),
    .A2(n1052),
    .B(n1056),
    .ZN(f_84_)
  );
  AOI21_X1 n_n85 (
    .A1(n1055),
    .A2(n1060),
    .B(n1064),
    .ZN(f_85_)
  );
  AOI21_X1 n_n86 (
    .A1(n1063),
    .A2(n1068),
    .B(n1072),
    .ZN(f_86_)
  );
  AOI21_X1 n_n87 (
    .A1(n1071),
    .A2(n1076),
    .B(n1080),
    .ZN(f_87_)
  );
  AOI21_X1 n_n88 (
    .A1(n1079),
    .A2(n1084),
    .B(n1088),
    .ZN(f_88_)
  );
  AOI21_X1 n_n89 (
    .A1(n1087),
    .A2(n1092),
    .B(n1096),
    .ZN(f_89_)
  );
  AOI21_X1 n_n90 (
    .A1(n1095),
    .A2(n1100),
    .B(n1104),
    .ZN(f_90_)
  );
  AOI21_X1 n_n91 (
    .A1(n1103),
    .A2(n1108),
    .B(n1112),
    .ZN(f_91_)
  );
  AOI21_X1 n_n92 (
    .A1(n1111),
    .A2(n1116),
    .B(n1120),
    .ZN(f_92_)
  );
  AOI21_X1 n_n93 (
    .A1(n1119),
    .A2(n1124),
    .B(n1128),
    .ZN(f_93_)
  );
  AOI21_X1 n_n94 (
    .A1(n1127),
    .A2(n1132),
    .B(n1136),
    .ZN(f_94_)
  );
  AOI21_X1 n_n95 (
    .A1(n1135),
    .A2(n1140),
    .B(n1144),
    .ZN(f_95_)
  );
  AOI21_X1 n_n96 (
    .A1(n1143),
    .A2(n1148),
    .B(n1152),
    .ZN(f_96_)
  );
  AOI21_X1 n_n97 (
    .A1(n1151),
    .A2(n1156),
    .B(n1160),
    .ZN(f_97_)
  );
  AOI21_X1 n_n98 (
    .A1(n1159),
    .A2(n1164),
    .B(n1168),
    .ZN(f_98_)
  );
  AOI21_X1 n_n99 (
    .A1(n1167),
    .A2(n1172),
    .B(n1176),
    .ZN(f_99_)
  );
  AOI21_X1 n_n100 (
    .A1(n1175),
    .A2(n1180),
    .B(n1184),
    .ZN(f_100_)
  );
  AOI21_X1 n_n101 (
    .A1(n1183),
    .A2(n1188),
    .B(n1192),
    .ZN(f_101_)
  );
  AOI21_X1 n_n102 (
    .A1(n1191),
    .A2(n1196),
    .B(n1200),
    .ZN(f_102_)
  );
  AOI21_X1 n_n103 (
    .A1(n1199),
    .A2(n1204),
    .B(n1208),
    .ZN(f_103_)
  );
  AOI21_X1 n_n104 (
    .A1(n1207),
    .A2(n1212),
    .B(n1216),
    .ZN(f_104_)
  );
  AOI21_X1 n_n105 (
    .A1(n1215),
    .A2(n1220),
    .B(n1224),
    .ZN(f_105_)
  );
  AOI21_X1 n_n106 (
    .A1(n1223),
    .A2(n1228),
    .B(n1232),
    .ZN(f_106_)
  );
  AOI21_X1 n_n107 (
    .A1(n1231),
    .A2(n1236),
    .B(n1240),
    .ZN(f_107_)
  );
  AOI21_X1 n_n108 (
    .A1(n1239),
    .A2(n1244),
    .B(n1248),
    .ZN(f_108_)
  );
  AOI21_X1 n_n109 (
    .A1(n1247),
    .A2(n1252),
    .B(n1256),
    .ZN(f_109_)
  );
  AOI21_X1 n_n110 (
    .A1(n1255),
    .A2(n1260),
    .B(n1264),
    .ZN(f_110_)
  );
  AOI21_X1 n_n111 (
    .A1(n1263),
    .A2(n1268),
    .B(n1272),
    .ZN(f_111_)
  );
  AOI21_X1 n_n112 (
    .A1(n1271),
    .A2(n1276),
    .B(n1280),
    .ZN(f_112_)
  );
  AOI21_X1 n_n113 (
    .A1(n1279),
    .A2(n1284),
    .B(n1288),
    .ZN(f_113_)
  );
  AOI21_X1 n_n114 (
    .A1(n1287),
    .A2(n1292),
    .B(n1296),
    .ZN(f_114_)
  );
  AOI21_X1 n_n115 (
    .A1(n1295),
    .A2(n1300),
    .B(n1304),
    .ZN(f_115_)
  );
  AOI21_X1 n_n116 (
    .A1(n1303),
    .A2(n1308),
    .B(n1312),
    .ZN(f_116_)
  );
  AOI21_X1 n_n117 (
    .A1(n1311),
    .A2(n1316),
    .B(n1320),
    .ZN(f_117_)
  );
  AOI21_X1 n_n118 (
    .A1(n1319),
    .A2(n1324),
    .B(n1328),
    .ZN(f_118_)
  );
  AOI21_X1 n_n119 (
    .A1(n1327),
    .A2(n1332),
    .B(n1336),
    .ZN(f_119_)
  );
  AOI21_X1 n_n120 (
    .A1(n1335),
    .A2(n1340),
    .B(n1344),
    .ZN(f_120_)
  );
  AOI21_X1 n_n121 (
    .A1(n1343),
    .A2(n1348),
    .B(n1352),
    .ZN(f_121_)
  );
  AOI21_X1 n_n122 (
    .A1(n1351),
    .A2(n1356),
    .B(n1360),
    .ZN(f_122_)
  );
  AOI21_X1 n_n123 (
    .A1(n1359),
    .A2(n1364),
    .B(n1368),
    .ZN(f_123_)
  );
  AOI21_X1 n_n124 (
    .A1(n1367),
    .A2(n1372),
    .B(n1376),
    .ZN(f_124_)
  );
  AOI21_X1 n_n125 (
    .A1(n1375),
    .A2(n1380),
    .B(n1384),
    .ZN(f_125_)
  );
  AOI21_X1 n_n126 (
    .A1(n1383),
    .A2(n1388),
    .B(n1392),
    .ZN(f_126_)
  );
  AOI21_X1 n_n127 (
    .A1(n1391),
    .A2(n1396),
    .B(n1400),
    .ZN(f_127_)
  );
  AOI21_X1 n_n128 (
    .A1(n1397),
    .A2(n1398),
    .B(n1399),
    .ZN(cOut)
  );
  XOR2_X1 n_n129 (
    .A1(a_1_),
    .A2(b_1_),
    .Z(n392)
  );
  AND2_X2 n_n130 (
    .A1(a_1_),
    .A2(b_1_),
    .Z(n391)
  );
  OAI21_X1 n_n131 (
    .A1(a_0_),
    .A2(b_0_),
    .B(n390),
    .ZN(n396)
  );
  XOR2_X1 n_n132 (
    .A1(a_2_),
    .A2(b_2_),
    .Z(n400)
  );
  AND2_X2 n_n133 (
    .A1(a_2_),
    .A2(b_2_),
    .Z(n399)
  );
  AOI22_X1 n_n134 (
    .A1(a_2_),
    .A2(b_2_),
    .B1(n391),
    .B2(n396),
    .ZN(n404)
  );
  XOR2_X1 n_n135 (
    .A1(a_3_),
    .A2(b_3_),
    .Z(n408)
  );
  AND2_X2 n_n136 (
    .A1(a_3_),
    .A2(b_3_),
    .Z(n407)
  );
  AOI22_X1 n_n137 (
    .A1(a_3_),
    .A2(b_3_),
    .B1(n399),
    .B2(n404),
    .ZN(n412)
  );
  XOR2_X1 n_n138 (
    .A1(a_4_),
    .A2(b_4_),
    .Z(n416)
  );
  AND2_X2 n_n139 (
    .A1(a_4_),
    .A2(b_4_),
    .Z(n415)
  );
  AOI22_X1 n_n140 (
    .A1(a_4_),
    .A2(b_4_),
    .B1(n407),
    .B2(n412),
    .ZN(n420)
  );
  XOR2_X1 n_n141 (
    .A1(a_5_),
    .A2(b_5_),
    .Z(n424)
  );
  AND2_X2 n_n142 (
    .A1(a_5_),
    .A2(b_5_),
    .Z(n423)
  );
  AOI22_X1 n_n143 (
    .A1(a_5_),
    .A2(b_5_),
    .B1(n415),
    .B2(n420),
    .ZN(n428)
  );
  XOR2_X1 n_n144 (
    .A1(a_6_),
    .A2(b_6_),
    .Z(n432)
  );
  AND2_X2 n_n145 (
    .A1(a_6_),
    .A2(b_6_),
    .Z(n431)
  );
  AOI22_X1 n_n146 (
    .A1(a_6_),
    .A2(b_6_),
    .B1(n423),
    .B2(n428),
    .ZN(n436)
  );
  XOR2_X1 n_n147 (
    .A1(a_7_),
    .A2(b_7_),
    .Z(n440)
  );
  AND2_X2 n_n148 (
    .A1(a_7_),
    .A2(b_7_),
    .Z(n439)
  );
  AOI22_X1 n_n149 (
    .A1(a_7_),
    .A2(b_7_),
    .B1(n431),
    .B2(n436),
    .ZN(n444)
  );
  XOR2_X1 n_n150 (
    .A1(a_8_),
    .A2(b_8_),
    .Z(n448)
  );
  AND2_X2 n_n151 (
    .A1(a_8_),
    .A2(b_8_),
    .Z(n447)
  );
  AOI22_X1 n_n152 (
    .A1(a_8_),
    .A2(b_8_),
    .B1(n439),
    .B2(n444),
    .ZN(n452)
  );
  XOR2_X1 n_n153 (
    .A1(a_9_),
    .A2(b_9_),
    .Z(n456)
  );
  AND2_X2 n_n154 (
    .A1(a_9_),
    .A2(b_9_),
    .Z(n455)
  );
  AOI22_X1 n_n155 (
    .A1(a_9_),
    .A2(b_9_),
    .B1(n447),
    .B2(n452),
    .ZN(n460)
  );
  XOR2_X1 n_n156 (
    .A1(a_10_),
    .A2(b_10_),
    .Z(n464)
  );
  AND2_X2 n_n157 (
    .A1(a_10_),
    .A2(b_10_),
    .Z(n463)
  );
  AOI22_X1 n_n158 (
    .A1(a_10_),
    .A2(b_10_),
    .B1(n455),
    .B2(n460),
    .ZN(n468)
  );
  XOR2_X1 n_n159 (
    .A1(a_11_),
    .A2(b_11_),
    .Z(n472)
  );
  AND2_X2 n_n160 (
    .A1(a_11_),
    .A2(b_11_),
    .Z(n471)
  );
  AOI22_X1 n_n161 (
    .A1(a_11_),
    .A2(b_11_),
    .B1(n463),
    .B2(n468),
    .ZN(n476)
  );
  XOR2_X1 n_n162 (
    .A1(a_12_),
    .A2(b_12_),
    .Z(n480)
  );
  AND2_X2 n_n163 (
    .A1(a_12_),
    .A2(b_12_),
    .Z(n479)
  );
  AOI22_X1 n_n164 (
    .A1(a_12_),
    .A2(b_12_),
    .B1(n471),
    .B2(n476),
    .ZN(n484)
  );
  XOR2_X1 n_n165 (
    .A1(a_13_),
    .A2(b_13_),
    .Z(n488)
  );
  AND2_X2 n_n166 (
    .A1(a_13_),
    .A2(b_13_),
    .Z(n487)
  );
  AOI22_X1 n_n167 (
    .A1(a_13_),
    .A2(b_13_),
    .B1(n479),
    .B2(n484),
    .ZN(n492)
  );
  XOR2_X1 n_n168 (
    .A1(a_14_),
    .A2(b_14_),
    .Z(n496)
  );
  AND2_X2 n_n169 (
    .A1(a_14_),
    .A2(b_14_),
    .Z(n495)
  );
  AOI22_X1 n_n170 (
    .A1(a_14_),
    .A2(b_14_),
    .B1(n487),
    .B2(n492),
    .ZN(n500)
  );
  XOR2_X1 n_n171 (
    .A1(a_15_),
    .A2(b_15_),
    .Z(n504)
  );
  AND2_X2 n_n172 (
    .A1(a_15_),
    .A2(b_15_),
    .Z(n503)
  );
  AOI22_X1 n_n173 (
    .A1(a_15_),
    .A2(b_15_),
    .B1(n495),
    .B2(n500),
    .ZN(n508)
  );
  XOR2_X1 n_n174 (
    .A1(a_16_),
    .A2(b_16_),
    .Z(n512)
  );
  AND2_X2 n_n175 (
    .A1(a_16_),
    .A2(b_16_),
    .Z(n511)
  );
  AOI22_X1 n_n176 (
    .A1(a_16_),
    .A2(b_16_),
    .B1(n503),
    .B2(n508),
    .ZN(n516)
  );
  XOR2_X1 n_n177 (
    .A1(a_17_),
    .A2(b_17_),
    .Z(n520)
  );
  AND2_X2 n_n178 (
    .A1(a_17_),
    .A2(b_17_),
    .Z(n519)
  );
  AOI22_X1 n_n179 (
    .A1(a_17_),
    .A2(b_17_),
    .B1(n511),
    .B2(n516),
    .ZN(n524)
  );
  XOR2_X1 n_n180 (
    .A1(a_18_),
    .A2(b_18_),
    .Z(n528)
  );
  AND2_X2 n_n181 (
    .A1(a_18_),
    .A2(b_18_),
    .Z(n527)
  );
  AOI22_X1 n_n182 (
    .A1(a_18_),
    .A2(b_18_),
    .B1(n519),
    .B2(n524),
    .ZN(n532)
  );
  XOR2_X1 n_n183 (
    .A1(a_19_),
    .A2(b_19_),
    .Z(n536)
  );
  AND2_X2 n_n184 (
    .A1(a_19_),
    .A2(b_19_),
    .Z(n535)
  );
  AOI22_X1 n_n185 (
    .A1(a_19_),
    .A2(b_19_),
    .B1(n527),
    .B2(n532),
    .ZN(n540)
  );
  XOR2_X1 n_n186 (
    .A1(a_20_),
    .A2(b_20_),
    .Z(n544)
  );
  AND2_X2 n_n187 (
    .A1(a_20_),
    .A2(b_20_),
    .Z(n543)
  );
  AOI22_X1 n_n188 (
    .A1(a_20_),
    .A2(b_20_),
    .B1(n535),
    .B2(n540),
    .ZN(n548)
  );
  XOR2_X1 n_n189 (
    .A1(a_21_),
    .A2(b_21_),
    .Z(n552)
  );
  AND2_X2 n_n190 (
    .A1(a_21_),
    .A2(b_21_),
    .Z(n551)
  );
  AOI22_X1 n_n191 (
    .A1(a_21_),
    .A2(b_21_),
    .B1(n543),
    .B2(n548),
    .ZN(n556)
  );
  XOR2_X1 n_n192 (
    .A1(a_22_),
    .A2(b_22_),
    .Z(n560)
  );
  AND2_X2 n_n193 (
    .A1(a_22_),
    .A2(b_22_),
    .Z(n559)
  );
  AOI22_X1 n_n194 (
    .A1(a_22_),
    .A2(b_22_),
    .B1(n551),
    .B2(n556),
    .ZN(n564)
  );
  XOR2_X1 n_n195 (
    .A1(a_23_),
    .A2(b_23_),
    .Z(n568)
  );
  AND2_X2 n_n196 (
    .A1(a_23_),
    .A2(b_23_),
    .Z(n567)
  );
  AOI22_X1 n_n197 (
    .A1(a_23_),
    .A2(b_23_),
    .B1(n559),
    .B2(n564),
    .ZN(n572)
  );
  XOR2_X1 n_n198 (
    .A1(a_24_),
    .A2(b_24_),
    .Z(n576)
  );
  AND2_X2 n_n199 (
    .A1(a_24_),
    .A2(b_24_),
    .Z(n575)
  );
  AOI22_X1 n_n200 (
    .A1(a_24_),
    .A2(b_24_),
    .B1(n567),
    .B2(n572),
    .ZN(n580)
  );
  XOR2_X1 n_n201 (
    .A1(a_25_),
    .A2(b_25_),
    .Z(n584)
  );
  AND2_X2 n_n202 (
    .A1(a_25_),
    .A2(b_25_),
    .Z(n583)
  );
  AOI22_X1 n_n203 (
    .A1(a_25_),
    .A2(b_25_),
    .B1(n575),
    .B2(n580),
    .ZN(n588)
  );
  XOR2_X1 n_n204 (
    .A1(a_26_),
    .A2(b_26_),
    .Z(n592)
  );
  AND2_X2 n_n205 (
    .A1(a_26_),
    .A2(b_26_),
    .Z(n591)
  );
  AOI22_X1 n_n206 (
    .A1(a_26_),
    .A2(b_26_),
    .B1(n583),
    .B2(n588),
    .ZN(n596)
  );
  XOR2_X1 n_n207 (
    .A1(a_27_),
    .A2(b_27_),
    .Z(n600)
  );
  AND2_X2 n_n208 (
    .A1(a_27_),
    .A2(b_27_),
    .Z(n599)
  );
  AOI22_X1 n_n209 (
    .A1(a_27_),
    .A2(b_27_),
    .B1(n591),
    .B2(n596),
    .ZN(n604)
  );
  XOR2_X1 n_n210 (
    .A1(a_28_),
    .A2(b_28_),
    .Z(n608)
  );
  AND2_X2 n_n211 (
    .A1(a_28_),
    .A2(b_28_),
    .Z(n607)
  );
  AOI22_X1 n_n212 (
    .A1(a_28_),
    .A2(b_28_),
    .B1(n599),
    .B2(n604),
    .ZN(n612)
  );
  XOR2_X1 n_n213 (
    .A1(a_29_),
    .A2(b_29_),
    .Z(n616)
  );
  AND2_X2 n_n214 (
    .A1(a_29_),
    .A2(b_29_),
    .Z(n615)
  );
  AOI22_X1 n_n215 (
    .A1(a_29_),
    .A2(b_29_),
    .B1(n607),
    .B2(n612),
    .ZN(n620)
  );
  XOR2_X1 n_n216 (
    .A1(a_30_),
    .A2(b_30_),
    .Z(n624)
  );
  AND2_X2 n_n217 (
    .A1(a_30_),
    .A2(b_30_),
    .Z(n623)
  );
  AOI22_X1 n_n218 (
    .A1(a_30_),
    .A2(b_30_),
    .B1(n615),
    .B2(n620),
    .ZN(n628)
  );
  XOR2_X1 n_n219 (
    .A1(a_31_),
    .A2(b_31_),
    .Z(n632)
  );
  AND2_X2 n_n220 (
    .A1(a_31_),
    .A2(b_31_),
    .Z(n631)
  );
  AOI22_X1 n_n221 (
    .A1(a_31_),
    .A2(b_31_),
    .B1(n623),
    .B2(n628),
    .ZN(n636)
  );
  XOR2_X1 n_n222 (
    .A1(a_32_),
    .A2(b_32_),
    .Z(n640)
  );
  AND2_X2 n_n223 (
    .A1(a_32_),
    .A2(b_32_),
    .Z(n639)
  );
  AOI22_X1 n_n224 (
    .A1(a_32_),
    .A2(b_32_),
    .B1(n631),
    .B2(n636),
    .ZN(n644)
  );
  XOR2_X1 n_n225 (
    .A1(a_33_),
    .A2(b_33_),
    .Z(n648)
  );
  AND2_X2 n_n226 (
    .A1(a_33_),
    .A2(b_33_),
    .Z(n647)
  );
  AOI22_X1 n_n227 (
    .A1(a_33_),
    .A2(b_33_),
    .B1(n639),
    .B2(n644),
    .ZN(n652)
  );
  XOR2_X1 n_n228 (
    .A1(a_34_),
    .A2(b_34_),
    .Z(n656)
  );
  AND2_X2 n_n229 (
    .A1(a_34_),
    .A2(b_34_),
    .Z(n655)
  );
  AOI22_X1 n_n230 (
    .A1(a_34_),
    .A2(b_34_),
    .B1(n647),
    .B2(n652),
    .ZN(n660)
  );
  XOR2_X1 n_n231 (
    .A1(a_35_),
    .A2(b_35_),
    .Z(n664)
  );
  AND2_X2 n_n232 (
    .A1(a_35_),
    .A2(b_35_),
    .Z(n663)
  );
  AOI22_X1 n_n233 (
    .A1(a_35_),
    .A2(b_35_),
    .B1(n655),
    .B2(n660),
    .ZN(n668)
  );
  XOR2_X1 n_n234 (
    .A1(a_36_),
    .A2(b_36_),
    .Z(n672)
  );
  AND2_X2 n_n235 (
    .A1(a_36_),
    .A2(b_36_),
    .Z(n671)
  );
  AOI22_X1 n_n236 (
    .A1(a_36_),
    .A2(b_36_),
    .B1(n663),
    .B2(n668),
    .ZN(n676)
  );
  XOR2_X1 n_n237 (
    .A1(a_37_),
    .A2(b_37_),
    .Z(n680)
  );
  AND2_X2 n_n238 (
    .A1(a_37_),
    .A2(b_37_),
    .Z(n679)
  );
  AOI22_X1 n_n239 (
    .A1(a_37_),
    .A2(b_37_),
    .B1(n671),
    .B2(n676),
    .ZN(n684)
  );
  XOR2_X1 n_n240 (
    .A1(a_38_),
    .A2(b_38_),
    .Z(n688)
  );
  AND2_X2 n_n241 (
    .A1(a_38_),
    .A2(b_38_),
    .Z(n687)
  );
  AOI22_X1 n_n242 (
    .A1(a_38_),
    .A2(b_38_),
    .B1(n679),
    .B2(n684),
    .ZN(n692)
  );
  XOR2_X1 n_n243 (
    .A1(a_39_),
    .A2(b_39_),
    .Z(n696)
  );
  AND2_X2 n_n244 (
    .A1(a_39_),
    .A2(b_39_),
    .Z(n695)
  );
  AOI22_X1 n_n245 (
    .A1(a_39_),
    .A2(b_39_),
    .B1(n687),
    .B2(n692),
    .ZN(n700)
  );
  XOR2_X1 n_n246 (
    .A1(a_40_),
    .A2(b_40_),
    .Z(n704)
  );
  AND2_X2 n_n247 (
    .A1(a_40_),
    .A2(b_40_),
    .Z(n703)
  );
  AOI22_X1 n_n248 (
    .A1(a_40_),
    .A2(b_40_),
    .B1(n695),
    .B2(n700),
    .ZN(n708)
  );
  XOR2_X1 n_n249 (
    .A1(a_41_),
    .A2(b_41_),
    .Z(n712)
  );
  AND2_X2 n_n250 (
    .A1(a_41_),
    .A2(b_41_),
    .Z(n711)
  );
  AOI22_X1 n_n251 (
    .A1(a_41_),
    .A2(b_41_),
    .B1(n703),
    .B2(n708),
    .ZN(n716)
  );
  XOR2_X1 n_n252 (
    .A1(a_42_),
    .A2(b_42_),
    .Z(n720)
  );
  AND2_X2 n_n253 (
    .A1(a_42_),
    .A2(b_42_),
    .Z(n719)
  );
  AOI22_X1 n_n254 (
    .A1(a_42_),
    .A2(b_42_),
    .B1(n711),
    .B2(n716),
    .ZN(n724)
  );
  XOR2_X1 n_n255 (
    .A1(a_43_),
    .A2(b_43_),
    .Z(n728)
  );
  AND2_X2 n_n256 (
    .A1(a_43_),
    .A2(b_43_),
    .Z(n727)
  );
  AOI22_X1 n_n257 (
    .A1(a_43_),
    .A2(b_43_),
    .B1(n719),
    .B2(n724),
    .ZN(n732)
  );
  XOR2_X1 n_n258 (
    .A1(a_44_),
    .A2(b_44_),
    .Z(n736)
  );
  AND2_X2 n_n259 (
    .A1(a_44_),
    .A2(b_44_),
    .Z(n735)
  );
  AOI22_X1 n_n260 (
    .A1(a_44_),
    .A2(b_44_),
    .B1(n727),
    .B2(n732),
    .ZN(n740)
  );
  XOR2_X1 n_n261 (
    .A1(a_45_),
    .A2(b_45_),
    .Z(n744)
  );
  AND2_X2 n_n262 (
    .A1(a_45_),
    .A2(b_45_),
    .Z(n743)
  );
  AOI22_X1 n_n263 (
    .A1(a_45_),
    .A2(b_45_),
    .B1(n735),
    .B2(n740),
    .ZN(n748)
  );
  XOR2_X1 n_n264 (
    .A1(a_46_),
    .A2(b_46_),
    .Z(n752)
  );
  AND2_X2 n_n265 (
    .A1(a_46_),
    .A2(b_46_),
    .Z(n751)
  );
  AOI22_X1 n_n266 (
    .A1(a_46_),
    .A2(b_46_),
    .B1(n743),
    .B2(n748),
    .ZN(n756)
  );
  XOR2_X1 n_n267 (
    .A1(a_47_),
    .A2(b_47_),
    .Z(n760)
  );
  AND2_X2 n_n268 (
    .A1(a_47_),
    .A2(b_47_),
    .Z(n759)
  );
  AOI22_X1 n_n269 (
    .A1(a_47_),
    .A2(b_47_),
    .B1(n751),
    .B2(n756),
    .ZN(n764)
  );
  XOR2_X1 n_n270 (
    .A1(a_48_),
    .A2(b_48_),
    .Z(n768)
  );
  AND2_X2 n_n271 (
    .A1(a_48_),
    .A2(b_48_),
    .Z(n767)
  );
  AOI22_X1 n_n272 (
    .A1(a_48_),
    .A2(b_48_),
    .B1(n759),
    .B2(n764),
    .ZN(n772)
  );
  XOR2_X1 n_n273 (
    .A1(a_49_),
    .A2(b_49_),
    .Z(n776)
  );
  AND2_X2 n_n274 (
    .A1(a_49_),
    .A2(b_49_),
    .Z(n775)
  );
  AOI22_X1 n_n275 (
    .A1(a_49_),
    .A2(b_49_),
    .B1(n767),
    .B2(n772),
    .ZN(n780)
  );
  XOR2_X1 n_n276 (
    .A1(a_50_),
    .A2(b_50_),
    .Z(n784)
  );
  AND2_X2 n_n277 (
    .A1(a_50_),
    .A2(b_50_),
    .Z(n783)
  );
  AOI22_X1 n_n278 (
    .A1(a_50_),
    .A2(b_50_),
    .B1(n775),
    .B2(n780),
    .ZN(n788)
  );
  XOR2_X1 n_n279 (
    .A1(a_51_),
    .A2(b_51_),
    .Z(n792)
  );
  AND2_X2 n_n280 (
    .A1(a_51_),
    .A2(b_51_),
    .Z(n791)
  );
  AOI22_X1 n_n281 (
    .A1(a_51_),
    .A2(b_51_),
    .B1(n783),
    .B2(n788),
    .ZN(n796)
  );
  XOR2_X1 n_n282 (
    .A1(a_52_),
    .A2(b_52_),
    .Z(n800)
  );
  AND2_X2 n_n283 (
    .A1(a_52_),
    .A2(b_52_),
    .Z(n799)
  );
  AOI22_X1 n_n284 (
    .A1(a_52_),
    .A2(b_52_),
    .B1(n791),
    .B2(n796),
    .ZN(n804)
  );
  XOR2_X1 n_n285 (
    .A1(a_53_),
    .A2(b_53_),
    .Z(n808)
  );
  AND2_X2 n_n286 (
    .A1(a_53_),
    .A2(b_53_),
    .Z(n807)
  );
  AOI22_X1 n_n287 (
    .A1(a_53_),
    .A2(b_53_),
    .B1(n799),
    .B2(n804),
    .ZN(n812)
  );
  XOR2_X1 n_n288 (
    .A1(a_54_),
    .A2(b_54_),
    .Z(n816)
  );
  AND2_X2 n_n289 (
    .A1(a_54_),
    .A2(b_54_),
    .Z(n815)
  );
  AOI22_X1 n_n290 (
    .A1(a_54_),
    .A2(b_54_),
    .B1(n807),
    .B2(n812),
    .ZN(n820)
  );
  XOR2_X1 n_n291 (
    .A1(a_55_),
    .A2(b_55_),
    .Z(n824)
  );
  AND2_X2 n_n292 (
    .A1(a_55_),
    .A2(b_55_),
    .Z(n823)
  );
  AOI22_X1 n_n293 (
    .A1(a_55_),
    .A2(b_55_),
    .B1(n815),
    .B2(n820),
    .ZN(n828)
  );
  XOR2_X1 n_n294 (
    .A1(a_56_),
    .A2(b_56_),
    .Z(n832)
  );
  AND2_X2 n_n295 (
    .A1(a_56_),
    .A2(b_56_),
    .Z(n831)
  );
  AOI22_X1 n_n296 (
    .A1(a_56_),
    .A2(b_56_),
    .B1(n823),
    .B2(n828),
    .ZN(n836)
  );
  XOR2_X1 n_n297 (
    .A1(a_57_),
    .A2(b_57_),
    .Z(n840)
  );
  AND2_X2 n_n298 (
    .A1(a_57_),
    .A2(b_57_),
    .Z(n839)
  );
  AOI22_X1 n_n299 (
    .A1(a_57_),
    .A2(b_57_),
    .B1(n831),
    .B2(n836),
    .ZN(n844)
  );
  XOR2_X1 n_n300 (
    .A1(a_58_),
    .A2(b_58_),
    .Z(n848)
  );
  AND2_X2 n_n301 (
    .A1(a_58_),
    .A2(b_58_),
    .Z(n847)
  );
  AOI22_X1 n_n302 (
    .A1(a_58_),
    .A2(b_58_),
    .B1(n839),
    .B2(n844),
    .ZN(n852)
  );
  XOR2_X1 n_n303 (
    .A1(a_59_),
    .A2(b_59_),
    .Z(n856)
  );
  AND2_X2 n_n304 (
    .A1(a_59_),
    .A2(b_59_),
    .Z(n855)
  );
  AOI22_X1 n_n305 (
    .A1(a_59_),
    .A2(b_59_),
    .B1(n847),
    .B2(n852),
    .ZN(n860)
  );
  XOR2_X1 n_n306 (
    .A1(a_60_),
    .A2(b_60_),
    .Z(n864)
  );
  AND2_X2 n_n307 (
    .A1(a_60_),
    .A2(b_60_),
    .Z(n863)
  );
  AOI22_X1 n_n308 (
    .A1(a_60_),
    .A2(b_60_),
    .B1(n855),
    .B2(n860),
    .ZN(n868)
  );
  XOR2_X1 n_n309 (
    .A1(a_61_),
    .A2(b_61_),
    .Z(n872)
  );
  AND2_X2 n_n310 (
    .A1(a_61_),
    .A2(b_61_),
    .Z(n871)
  );
  AOI22_X1 n_n311 (
    .A1(a_61_),
    .A2(b_61_),
    .B1(n863),
    .B2(n868),
    .ZN(n876)
  );
  XOR2_X1 n_n312 (
    .A1(a_62_),
    .A2(b_62_),
    .Z(n880)
  );
  AND2_X2 n_n313 (
    .A1(a_62_),
    .A2(b_62_),
    .Z(n879)
  );
  AOI22_X1 n_n314 (
    .A1(a_62_),
    .A2(b_62_),
    .B1(n871),
    .B2(n876),
    .ZN(n884)
  );
  XOR2_X1 n_n315 (
    .A1(a_63_),
    .A2(b_63_),
    .Z(n888)
  );
  AND2_X2 n_n316 (
    .A1(a_63_),
    .A2(b_63_),
    .Z(n887)
  );
  AOI22_X1 n_n317 (
    .A1(a_63_),
    .A2(b_63_),
    .B1(n879),
    .B2(n884),
    .ZN(n892)
  );
  XOR2_X1 n_n318 (
    .A1(a_64_),
    .A2(b_64_),
    .Z(n896)
  );
  AND2_X2 n_n319 (
    .A1(a_64_),
    .A2(b_64_),
    .Z(n895)
  );
  AOI22_X1 n_n320 (
    .A1(a_64_),
    .A2(b_64_),
    .B1(n887),
    .B2(n892),
    .ZN(n900)
  );
  XOR2_X1 n_n321 (
    .A1(a_65_),
    .A2(b_65_),
    .Z(n904)
  );
  AND2_X2 n_n322 (
    .A1(a_65_),
    .A2(b_65_),
    .Z(n903)
  );
  AOI22_X1 n_n323 (
    .A1(a_65_),
    .A2(b_65_),
    .B1(n895),
    .B2(n900),
    .ZN(n908)
  );
  XOR2_X1 n_n324 (
    .A1(a_66_),
    .A2(b_66_),
    .Z(n912)
  );
  AND2_X2 n_n325 (
    .A1(a_66_),
    .A2(b_66_),
    .Z(n911)
  );
  AOI22_X1 n_n326 (
    .A1(a_66_),
    .A2(b_66_),
    .B1(n903),
    .B2(n908),
    .ZN(n916)
  );
  XOR2_X1 n_n327 (
    .A1(a_67_),
    .A2(b_67_),
    .Z(n920)
  );
  AND2_X2 n_n328 (
    .A1(a_67_),
    .A2(b_67_),
    .Z(n919)
  );
  AOI22_X1 n_n329 (
    .A1(a_67_),
    .A2(b_67_),
    .B1(n911),
    .B2(n916),
    .ZN(n924)
  );
  XOR2_X1 n_n330 (
    .A1(a_68_),
    .A2(b_68_),
    .Z(n928)
  );
  AND2_X2 n_n331 (
    .A1(a_68_),
    .A2(b_68_),
    .Z(n927)
  );
  AOI22_X1 n_n332 (
    .A1(a_68_),
    .A2(b_68_),
    .B1(n919),
    .B2(n924),
    .ZN(n932)
  );
  XOR2_X1 n_n333 (
    .A1(a_69_),
    .A2(b_69_),
    .Z(n936)
  );
  AND2_X2 n_n334 (
    .A1(a_69_),
    .A2(b_69_),
    .Z(n935)
  );
  AOI22_X1 n_n335 (
    .A1(a_69_),
    .A2(b_69_),
    .B1(n927),
    .B2(n932),
    .ZN(n940)
  );
  XOR2_X1 n_n336 (
    .A1(a_70_),
    .A2(b_70_),
    .Z(n944)
  );
  AND2_X2 n_n337 (
    .A1(a_70_),
    .A2(b_70_),
    .Z(n943)
  );
  AOI22_X1 n_n338 (
    .A1(a_70_),
    .A2(b_70_),
    .B1(n935),
    .B2(n940),
    .ZN(n948)
  );
  XOR2_X1 n_n339 (
    .A1(a_71_),
    .A2(b_71_),
    .Z(n952)
  );
  AND2_X2 n_n340 (
    .A1(a_71_),
    .A2(b_71_),
    .Z(n951)
  );
  AOI22_X1 n_n341 (
    .A1(a_71_),
    .A2(b_71_),
    .B1(n943),
    .B2(n948),
    .ZN(n956)
  );
  XOR2_X1 n_n342 (
    .A1(a_72_),
    .A2(b_72_),
    .Z(n960)
  );
  AND2_X2 n_n343 (
    .A1(a_72_),
    .A2(b_72_),
    .Z(n959)
  );
  AOI22_X1 n_n344 (
    .A1(a_72_),
    .A2(b_72_),
    .B1(n951),
    .B2(n956),
    .ZN(n964)
  );
  XOR2_X1 n_n345 (
    .A1(a_73_),
    .A2(b_73_),
    .Z(n968)
  );
  AND2_X2 n_n346 (
    .A1(a_73_),
    .A2(b_73_),
    .Z(n967)
  );
  AOI22_X1 n_n347 (
    .A1(a_73_),
    .A2(b_73_),
    .B1(n959),
    .B2(n964),
    .ZN(n972)
  );
  XOR2_X1 n_n348 (
    .A1(a_74_),
    .A2(b_74_),
    .Z(n976)
  );
  AND2_X2 n_n349 (
    .A1(a_74_),
    .A2(b_74_),
    .Z(n975)
  );
  AOI22_X1 n_n350 (
    .A1(a_74_),
    .A2(b_74_),
    .B1(n967),
    .B2(n972),
    .ZN(n980)
  );
  XOR2_X1 n_n351 (
    .A1(a_75_),
    .A2(b_75_),
    .Z(n984)
  );
  AND2_X2 n_n352 (
    .A1(a_75_),
    .A2(b_75_),
    .Z(n983)
  );
  AOI22_X1 n_n353 (
    .A1(a_75_),
    .A2(b_75_),
    .B1(n975),
    .B2(n980),
    .ZN(n988)
  );
  XOR2_X1 n_n354 (
    .A1(a_76_),
    .A2(b_76_),
    .Z(n992)
  );
  XOR2_X1 n_n355 (
    .A1(a_77_),
    .A2(b_77_),
    .Z(n1000)
  );
  AND2_X2 n_n356 (
    .A1(a_76_),
    .A2(b_76_),
    .Z(n991)
  );
  AOI22_X1 n_n357 (
    .A1(a_76_),
    .A2(b_76_),
    .B1(n983),
    .B2(n988),
    .ZN(n996)
  );
  AOI22_X1 n_n358 (
    .A1(a_77_),
    .A2(b_77_),
    .B1(n991),
    .B2(n996),
    .ZN(n1004)
  );
  XOR2_X1 n_n359 (
    .A1(a_78_),
    .A2(b_78_),
    .Z(n1008)
  );
  AND2_X2 n_n360 (
    .A1(a_77_),
    .A2(b_77_),
    .Z(n999)
  );
  AND2_X2 n_n361 (
    .A1(a_78_),
    .A2(b_78_),
    .Z(n1007)
  );
  AOI22_X1 n_n362 (
    .A1(a_78_),
    .A2(b_78_),
    .B1(n1004),
    .B2(n999),
    .ZN(n1012)
  );
  XOR2_X1 n_n363 (
    .A1(a_79_),
    .A2(b_79_),
    .Z(n1016)
  );
  AND2_X2 n_n364 (
    .A1(a_79_),
    .A2(b_79_),
    .Z(n1015)
  );
  AOI22_X1 n_n365 (
    .A1(a_79_),
    .A2(b_79_),
    .B1(n1007),
    .B2(n1012),
    .ZN(n1020)
  );
  XOR2_X1 n_n366 (
    .A1(a_80_),
    .A2(b_80_),
    .Z(n1024)
  );
  AND2_X2 n_n367 (
    .A1(a_80_),
    .A2(b_80_),
    .Z(n1023)
  );
  AOI22_X1 n_n368 (
    .A1(a_80_),
    .A2(b_80_),
    .B1(n1015),
    .B2(n1020),
    .ZN(n1028)
  );
  XOR2_X1 n_n369 (
    .A1(a_81_),
    .A2(b_81_),
    .Z(n1032)
  );
  AND2_X2 n_n370 (
    .A1(a_81_),
    .A2(b_81_),
    .Z(n1031)
  );
  AOI22_X1 n_n371 (
    .A1(a_81_),
    .A2(b_81_),
    .B1(n1023),
    .B2(n1028),
    .ZN(n1036)
  );
  XOR2_X1 n_n372 (
    .A1(a_82_),
    .A2(b_82_),
    .Z(n1040)
  );
  AND2_X2 n_n373 (
    .A1(a_82_),
    .A2(b_82_),
    .Z(n1039)
  );
  AOI22_X1 n_n374 (
    .A1(a_82_),
    .A2(b_82_),
    .B1(n1031),
    .B2(n1036),
    .ZN(n1044)
  );
  XOR2_X1 n_n375 (
    .A1(a_83_),
    .A2(b_83_),
    .Z(n1048)
  );
  AND2_X2 n_n376 (
    .A1(a_83_),
    .A2(b_83_),
    .Z(n1047)
  );
  AOI22_X1 n_n377 (
    .A1(a_83_),
    .A2(b_83_),
    .B1(n1039),
    .B2(n1044),
    .ZN(n1052)
  );
  XOR2_X1 n_n378 (
    .A1(a_84_),
    .A2(b_84_),
    .Z(n1056)
  );
  AND2_X2 n_n379 (
    .A1(a_84_),
    .A2(b_84_),
    .Z(n1055)
  );
  AOI22_X1 n_n380 (
    .A1(a_84_),
    .A2(b_84_),
    .B1(n1047),
    .B2(n1052),
    .ZN(n1060)
  );
  XOR2_X1 n_n381 (
    .A1(a_85_),
    .A2(b_85_),
    .Z(n1064)
  );
  AND2_X2 n_n382 (
    .A1(a_85_),
    .A2(b_85_),
    .Z(n1063)
  );
  AOI22_X1 n_n383 (
    .A1(a_85_),
    .A2(b_85_),
    .B1(n1055),
    .B2(n1060),
    .ZN(n1068)
  );
  XOR2_X1 n_n384 (
    .A1(a_86_),
    .A2(b_86_),
    .Z(n1072)
  );
  AND2_X2 n_n385 (
    .A1(a_86_),
    .A2(b_86_),
    .Z(n1071)
  );
  AOI22_X1 n_n386 (
    .A1(a_86_),
    .A2(b_86_),
    .B1(n1063),
    .B2(n1068),
    .ZN(n1076)
  );
  XOR2_X1 n_n387 (
    .A1(a_87_),
    .A2(b_87_),
    .Z(n1080)
  );
  AND2_X2 n_n388 (
    .A1(a_87_),
    .A2(b_87_),
    .Z(n1079)
  );
  AOI22_X1 n_n389 (
    .A1(a_87_),
    .A2(b_87_),
    .B1(n1071),
    .B2(n1076),
    .ZN(n1084)
  );
  XOR2_X1 n_n390 (
    .A1(a_88_),
    .A2(b_88_),
    .Z(n1088)
  );
  AND2_X2 n_n391 (
    .A1(a_88_),
    .A2(b_88_),
    .Z(n1087)
  );
  AOI22_X1 n_n392 (
    .A1(a_88_),
    .A2(b_88_),
    .B1(n1079),
    .B2(n1084),
    .ZN(n1092)
  );
  XOR2_X1 n_n393 (
    .A1(a_89_),
    .A2(b_89_),
    .Z(n1096)
  );
  AND2_X2 n_n394 (
    .A1(a_89_),
    .A2(b_89_),
    .Z(n1095)
  );
  AOI22_X1 n_n395 (
    .A1(a_89_),
    .A2(b_89_),
    .B1(n1087),
    .B2(n1092),
    .ZN(n1100)
  );
  XOR2_X1 n_n396 (
    .A1(a_90_),
    .A2(b_90_),
    .Z(n1104)
  );
  AND2_X2 n_n397 (
    .A1(a_90_),
    .A2(b_90_),
    .Z(n1103)
  );
  AOI22_X1 n_n398 (
    .A1(a_90_),
    .A2(b_90_),
    .B1(n1095),
    .B2(n1100),
    .ZN(n1108)
  );
  XOR2_X1 n_n399 (
    .A1(a_91_),
    .A2(b_91_),
    .Z(n1112)
  );
  AND2_X2 n_n400 (
    .A1(a_91_),
    .A2(b_91_),
    .Z(n1111)
  );
  AOI22_X1 n_n401 (
    .A1(a_91_),
    .A2(b_91_),
    .B1(n1103),
    .B2(n1108),
    .ZN(n1116)
  );
  XOR2_X1 n_n402 (
    .A1(a_92_),
    .A2(b_92_),
    .Z(n1120)
  );
  AND2_X2 n_n403 (
    .A1(a_92_),
    .A2(b_92_),
    .Z(n1119)
  );
  AOI22_X1 n_n404 (
    .A1(a_92_),
    .A2(b_92_),
    .B1(n1111),
    .B2(n1116),
    .ZN(n1124)
  );
  XOR2_X1 n_n405 (
    .A1(a_93_),
    .A2(b_93_),
    .Z(n1128)
  );
  AND2_X2 n_n406 (
    .A1(a_93_),
    .A2(b_93_),
    .Z(n1127)
  );
  AOI22_X1 n_n407 (
    .A1(a_93_),
    .A2(b_93_),
    .B1(n1119),
    .B2(n1124),
    .ZN(n1132)
  );
  XOR2_X1 n_n408 (
    .A1(a_94_),
    .A2(b_94_),
    .Z(n1136)
  );
  AND2_X2 n_n409 (
    .A1(a_94_),
    .A2(b_94_),
    .Z(n1135)
  );
  AOI22_X1 n_n410 (
    .A1(a_94_),
    .A2(b_94_),
    .B1(n1127),
    .B2(n1132),
    .ZN(n1140)
  );
  XOR2_X1 n_n411 (
    .A1(a_95_),
    .A2(b_95_),
    .Z(n1144)
  );
  AND2_X2 n_n412 (
    .A1(a_95_),
    .A2(b_95_),
    .Z(n1143)
  );
  AOI22_X1 n_n413 (
    .A1(a_95_),
    .A2(b_95_),
    .B1(n1135),
    .B2(n1140),
    .ZN(n1148)
  );
  XOR2_X1 n_n414 (
    .A1(a_96_),
    .A2(b_96_),
    .Z(n1152)
  );
  AND2_X2 n_n415 (
    .A1(a_96_),
    .A2(b_96_),
    .Z(n1151)
  );
  AOI22_X1 n_n416 (
    .A1(a_96_),
    .A2(b_96_),
    .B1(n1143),
    .B2(n1148),
    .ZN(n1156)
  );
  XOR2_X1 n_n417 (
    .A1(a_97_),
    .A2(b_97_),
    .Z(n1160)
  );
  AND2_X2 n_n418 (
    .A1(a_97_),
    .A2(b_97_),
    .Z(n1159)
  );
  AOI22_X1 n_n419 (
    .A1(a_97_),
    .A2(b_97_),
    .B1(n1151),
    .B2(n1156),
    .ZN(n1164)
  );
  XOR2_X1 n_n420 (
    .A1(a_98_),
    .A2(b_98_),
    .Z(n1168)
  );
  AND2_X2 n_n421 (
    .A1(a_98_),
    .A2(b_98_),
    .Z(n1167)
  );
  AOI22_X1 n_n422 (
    .A1(a_98_),
    .A2(b_98_),
    .B1(n1159),
    .B2(n1164),
    .ZN(n1172)
  );
  XOR2_X1 n_n423 (
    .A1(a_99_),
    .A2(b_99_),
    .Z(n1176)
  );
  AND2_X2 n_n424 (
    .A1(a_99_),
    .A2(b_99_),
    .Z(n1175)
  );
  AOI22_X1 n_n425 (
    .A1(a_99_),
    .A2(b_99_),
    .B1(n1167),
    .B2(n1172),
    .ZN(n1180)
  );
  XOR2_X1 n_n426 (
    .A1(a_100_),
    .A2(b_100_),
    .Z(n1184)
  );
  AND2_X2 n_n427 (
    .A1(a_100_),
    .A2(b_100_),
    .Z(n1183)
  );
  AOI22_X1 n_n428 (
    .A1(a_100_),
    .A2(b_100_),
    .B1(n1175),
    .B2(n1180),
    .ZN(n1188)
  );
  XOR2_X1 n_n429 (
    .A1(a_101_),
    .A2(b_101_),
    .Z(n1192)
  );
  AND2_X2 n_n430 (
    .A1(a_101_),
    .A2(b_101_),
    .Z(n1191)
  );
  AOI22_X1 n_n431 (
    .A1(a_101_),
    .A2(b_101_),
    .B1(n1183),
    .B2(n1188),
    .ZN(n1196)
  );
  XOR2_X1 n_n432 (
    .A1(a_102_),
    .A2(b_102_),
    .Z(n1200)
  );
  AND2_X2 n_n433 (
    .A1(a_102_),
    .A2(b_102_),
    .Z(n1199)
  );
  AOI22_X1 n_n434 (
    .A1(a_102_),
    .A2(b_102_),
    .B1(n1191),
    .B2(n1196),
    .ZN(n1204)
  );
  XOR2_X1 n_n435 (
    .A1(a_103_),
    .A2(b_103_),
    .Z(n1208)
  );
  AND2_X2 n_n436 (
    .A1(a_103_),
    .A2(b_103_),
    .Z(n1207)
  );
  AOI22_X1 n_n437 (
    .A1(a_103_),
    .A2(b_103_),
    .B1(n1199),
    .B2(n1204),
    .ZN(n1212)
  );
  XOR2_X1 n_n438 (
    .A1(a_104_),
    .A2(b_104_),
    .Z(n1216)
  );
  AND2_X2 n_n439 (
    .A1(a_104_),
    .A2(b_104_),
    .Z(n1215)
  );
  AOI22_X1 n_n440 (
    .A1(a_104_),
    .A2(b_104_),
    .B1(n1207),
    .B2(n1212),
    .ZN(n1220)
  );
  XOR2_X1 n_n441 (
    .A1(a_105_),
    .A2(b_105_),
    .Z(n1224)
  );
  AND2_X2 n_n442 (
    .A1(a_105_),
    .A2(b_105_),
    .Z(n1223)
  );
  AOI22_X1 n_n443 (
    .A1(a_105_),
    .A2(b_105_),
    .B1(n1215),
    .B2(n1220),
    .ZN(n1228)
  );
  XOR2_X1 n_n444 (
    .A1(a_106_),
    .A2(b_106_),
    .Z(n1232)
  );
  AND2_X2 n_n445 (
    .A1(a_106_),
    .A2(b_106_),
    .Z(n1231)
  );
  AOI22_X1 n_n446 (
    .A1(a_106_),
    .A2(b_106_),
    .B1(n1223),
    .B2(n1228),
    .ZN(n1236)
  );
  XOR2_X1 n_n447 (
    .A1(a_107_),
    .A2(b_107_),
    .Z(n1240)
  );
  AND2_X2 n_n448 (
    .A1(a_107_),
    .A2(b_107_),
    .Z(n1239)
  );
  AOI22_X1 n_n449 (
    .A1(a_107_),
    .A2(b_107_),
    .B1(n1231),
    .B2(n1236),
    .ZN(n1244)
  );
  XOR2_X1 n_n450 (
    .A1(a_108_),
    .A2(b_108_),
    .Z(n1248)
  );
  AND2_X2 n_n451 (
    .A1(a_108_),
    .A2(b_108_),
    .Z(n1247)
  );
  AOI22_X1 n_n452 (
    .A1(a_108_),
    .A2(b_108_),
    .B1(n1239),
    .B2(n1244),
    .ZN(n1252)
  );
  XOR2_X1 n_n453 (
    .A1(a_109_),
    .A2(b_109_),
    .Z(n1256)
  );
  AND2_X2 n_n454 (
    .A1(a_109_),
    .A2(b_109_),
    .Z(n1255)
  );
  AOI22_X1 n_n455 (
    .A1(a_109_),
    .A2(b_109_),
    .B1(n1247),
    .B2(n1252),
    .ZN(n1260)
  );
  XOR2_X1 n_n456 (
    .A1(a_110_),
    .A2(b_110_),
    .Z(n1264)
  );
  AND2_X2 n_n457 (
    .A1(a_110_),
    .A2(b_110_),
    .Z(n1263)
  );
  AOI22_X1 n_n458 (
    .A1(a_110_),
    .A2(b_110_),
    .B1(n1255),
    .B2(n1260),
    .ZN(n1268)
  );
  XOR2_X1 n_n459 (
    .A1(a_111_),
    .A2(b_111_),
    .Z(n1272)
  );
  AND2_X2 n_n460 (
    .A1(a_111_),
    .A2(b_111_),
    .Z(n1271)
  );
  AOI22_X1 n_n461 (
    .A1(a_111_),
    .A2(b_111_),
    .B1(n1263),
    .B2(n1268),
    .ZN(n1276)
  );
  XOR2_X1 n_n462 (
    .A1(a_112_),
    .A2(b_112_),
    .Z(n1280)
  );
  AND2_X2 n_n463 (
    .A1(a_112_),
    .A2(b_112_),
    .Z(n1279)
  );
  AOI22_X1 n_n464 (
    .A1(a_112_),
    .A2(b_112_),
    .B1(n1271),
    .B2(n1276),
    .ZN(n1284)
  );
  XOR2_X1 n_n465 (
    .A1(a_113_),
    .A2(b_113_),
    .Z(n1288)
  );
  AND2_X2 n_n466 (
    .A1(a_113_),
    .A2(b_113_),
    .Z(n1287)
  );
  AOI22_X1 n_n467 (
    .A1(a_113_),
    .A2(b_113_),
    .B1(n1279),
    .B2(n1284),
    .ZN(n1292)
  );
  XOR2_X1 n_n468 (
    .A1(a_114_),
    .A2(b_114_),
    .Z(n1296)
  );
  AND2_X2 n_n469 (
    .A1(a_114_),
    .A2(b_114_),
    .Z(n1295)
  );
  AOI22_X1 n_n470 (
    .A1(a_114_),
    .A2(b_114_),
    .B1(n1287),
    .B2(n1292),
    .ZN(n1300)
  );
  XOR2_X1 n_n471 (
    .A1(a_115_),
    .A2(b_115_),
    .Z(n1304)
  );
  AND2_X2 n_n472 (
    .A1(a_115_),
    .A2(b_115_),
    .Z(n1303)
  );
  AOI22_X1 n_n473 (
    .A1(a_115_),
    .A2(b_115_),
    .B1(n1295),
    .B2(n1300),
    .ZN(n1308)
  );
  XOR2_X1 n_n474 (
    .A1(a_116_),
    .A2(b_116_),
    .Z(n1312)
  );
  AND2_X2 n_n475 (
    .A1(a_116_),
    .A2(b_116_),
    .Z(n1311)
  );
  AOI22_X1 n_n476 (
    .A1(a_116_),
    .A2(b_116_),
    .B1(n1303),
    .B2(n1308),
    .ZN(n1316)
  );
  XOR2_X1 n_n477 (
    .A1(a_117_),
    .A2(b_117_),
    .Z(n1320)
  );
  AND2_X2 n_n478 (
    .A1(a_117_),
    .A2(b_117_),
    .Z(n1319)
  );
  AOI22_X1 n_n479 (
    .A1(a_117_),
    .A2(b_117_),
    .B1(n1311),
    .B2(n1316),
    .ZN(n1324)
  );
  XOR2_X1 n_n480 (
    .A1(a_118_),
    .A2(b_118_),
    .Z(n1328)
  );
  AND2_X2 n_n481 (
    .A1(a_118_),
    .A2(b_118_),
    .Z(n1327)
  );
  AOI22_X1 n_n482 (
    .A1(a_118_),
    .A2(b_118_),
    .B1(n1319),
    .B2(n1324),
    .ZN(n1332)
  );
  XOR2_X1 n_n483 (
    .A1(a_119_),
    .A2(b_119_),
    .Z(n1336)
  );
  AND2_X2 n_n484 (
    .A1(a_119_),
    .A2(b_119_),
    .Z(n1335)
  );
  AOI22_X1 n_n485 (
    .A1(a_119_),
    .A2(b_119_),
    .B1(n1327),
    .B2(n1332),
    .ZN(n1340)
  );
  XOR2_X1 n_n486 (
    .A1(a_120_),
    .A2(b_120_),
    .Z(n1344)
  );
  AND2_X2 n_n487 (
    .A1(a_120_),
    .A2(b_120_),
    .Z(n1343)
  );
  AOI22_X1 n_n488 (
    .A1(a_120_),
    .A2(b_120_),
    .B1(n1335),
    .B2(n1340),
    .ZN(n1348)
  );
  XOR2_X1 n_n489 (
    .A1(a_121_),
    .A2(b_121_),
    .Z(n1352)
  );
  AND2_X2 n_n490 (
    .A1(a_121_),
    .A2(b_121_),
    .Z(n1351)
  );
  AOI22_X1 n_n491 (
    .A1(a_121_),
    .A2(b_121_),
    .B1(n1343),
    .B2(n1348),
    .ZN(n1356)
  );
  XOR2_X1 n_n492 (
    .A1(a_122_),
    .A2(b_122_),
    .Z(n1360)
  );
  AND2_X2 n_n493 (
    .A1(a_122_),
    .A2(b_122_),
    .Z(n1359)
  );
  AOI22_X1 n_n494 (
    .A1(a_122_),
    .A2(b_122_),
    .B1(n1351),
    .B2(n1356),
    .ZN(n1364)
  );
  XOR2_X1 n_n495 (
    .A1(a_123_),
    .A2(b_123_),
    .Z(n1368)
  );
  AND2_X2 n_n496 (
    .A1(a_123_),
    .A2(b_123_),
    .Z(n1367)
  );
  AOI22_X1 n_n497 (
    .A1(a_123_),
    .A2(b_123_),
    .B1(n1359),
    .B2(n1364),
    .ZN(n1372)
  );
  XOR2_X1 n_n498 (
    .A1(a_124_),
    .A2(b_124_),
    .Z(n1376)
  );
  AND2_X2 n_n499 (
    .A1(a_124_),
    .A2(b_124_),
    .Z(n1375)
  );
  AOI22_X1 n_n500 (
    .A1(a_124_),
    .A2(b_124_),
    .B1(n1367),
    .B2(n1372),
    .ZN(n1380)
  );
  XOR2_X1 n_n501 (
    .A1(a_125_),
    .A2(b_125_),
    .Z(n1384)
  );
  AND2_X2 n_n502 (
    .A1(a_125_),
    .A2(b_125_),
    .Z(n1383)
  );
  AOI22_X1 n_n503 (
    .A1(a_125_),
    .A2(b_125_),
    .B1(n1375),
    .B2(n1380),
    .ZN(n1388)
  );
  XOR2_X1 n_n504 (
    .A1(a_126_),
    .A2(b_126_),
    .Z(n1392)
  );
  AND2_X2 n_n505 (
    .A1(a_126_),
    .A2(b_126_),
    .Z(n1391)
  );
  AOI22_X1 n_n506 (
    .A1(a_126_),
    .A2(b_126_),
    .B1(n1383),
    .B2(n1388),
    .ZN(n1396)
  );
  XOR2_X1 n_n507 (
    .A1(a_127_),
    .A2(b_127_),
    .Z(n1400)
  );
  AOI21_X1 n_n508 (
    .A1(n1389),
    .A2(n1390),
    .B(n1391),
    .ZN(n1397)
  );
  AND2_X2 n_n509 (
    .A1(a_127_),
    .A2(b_127_),
    .Z(n1398)
  );
  AND2_X2 n_n510 (
    .A1(a_127_),
    .A2(b_127_),
    .Z(n1399)
  );
  AND2_X2 n_n511 (
    .A1(a_1_),
    .A2(b_1_),
    .Z(n390)
  );
  AOI21_X1 n_n512 (
    .A1(n1381),
    .A2(n1382),
    .B(n1383),
    .ZN(n1389)
  );
  AND2_X2 n_n513 (
    .A1(a_126_),
    .A2(b_126_),
    .Z(n1390)
  );
  AOI21_X1 n_n514 (
    .A1(n1373),
    .A2(n1374),
    .B(n1375),
    .ZN(n1381)
  );
  AND2_X2 n_n515 (
    .A1(a_125_),
    .A2(b_125_),
    .Z(n1382)
  );
  AOI21_X1 n_n516 (
    .A1(n1365),
    .A2(n1366),
    .B(n1367),
    .ZN(n1373)
  );
  AND2_X2 n_n517 (
    .A1(a_124_),
    .A2(b_124_),
    .Z(n1374)
  );
  AOI21_X1 n_n518 (
    .A1(n1357),
    .A2(n1358),
    .B(n1359),
    .ZN(n1365)
  );
  AND2_X2 n_n519 (
    .A1(a_123_),
    .A2(b_123_),
    .Z(n1366)
  );
  AOI21_X1 n_n520 (
    .A1(n1349),
    .A2(n1350),
    .B(n1351),
    .ZN(n1357)
  );
  AND2_X2 n_n521 (
    .A1(a_122_),
    .A2(b_122_),
    .Z(n1358)
  );
  AOI21_X1 n_n522 (
    .A1(n1341),
    .A2(n1342),
    .B(n1343),
    .ZN(n1349)
  );
  AND2_X2 n_n523 (
    .A1(a_121_),
    .A2(b_121_),
    .Z(n1350)
  );
  AOI21_X1 n_n524 (
    .A1(n1333),
    .A2(n1334),
    .B(n1335),
    .ZN(n1341)
  );
  AND2_X2 n_n525 (
    .A1(a_120_),
    .A2(b_120_),
    .Z(n1342)
  );
  AOI21_X1 n_n526 (
    .A1(n1325),
    .A2(n1326),
    .B(n1327),
    .ZN(n1333)
  );
  AND2_X2 n_n527 (
    .A1(a_119_),
    .A2(b_119_),
    .Z(n1334)
  );
  AOI21_X1 n_n528 (
    .A1(n1317),
    .A2(n1318),
    .B(n1319),
    .ZN(n1325)
  );
  AND2_X2 n_n529 (
    .A1(a_118_),
    .A2(b_118_),
    .Z(n1326)
  );
  AOI21_X1 n_n530 (
    .A1(n1309),
    .A2(n1310),
    .B(n1311),
    .ZN(n1317)
  );
  AND2_X2 n_n531 (
    .A1(a_117_),
    .A2(b_117_),
    .Z(n1318)
  );
  AOI21_X1 n_n532 (
    .A1(n1301),
    .A2(n1302),
    .B(n1303),
    .ZN(n1309)
  );
  AND2_X2 n_n533 (
    .A1(a_116_),
    .A2(b_116_),
    .Z(n1310)
  );
  AOI21_X1 n_n534 (
    .A1(n1293),
    .A2(n1294),
    .B(n1295),
    .ZN(n1301)
  );
  AND2_X2 n_n535 (
    .A1(a_115_),
    .A2(b_115_),
    .Z(n1302)
  );
  AOI21_X1 n_n536 (
    .A1(n1285),
    .A2(n1286),
    .B(n1287),
    .ZN(n1293)
  );
  AND2_X2 n_n537 (
    .A1(a_114_),
    .A2(b_114_),
    .Z(n1294)
  );
  AOI21_X1 n_n538 (
    .A1(n1277),
    .A2(n1278),
    .B(n1279),
    .ZN(n1285)
  );
  AND2_X2 n_n539 (
    .A1(a_113_),
    .A2(b_113_),
    .Z(n1286)
  );
  AOI21_X1 n_n540 (
    .A1(n1269),
    .A2(n1270),
    .B(n1271),
    .ZN(n1277)
  );
  AND2_X2 n_n541 (
    .A1(a_112_),
    .A2(b_112_),
    .Z(n1278)
  );
  AOI21_X1 n_n542 (
    .A1(n1261),
    .A2(n1262),
    .B(n1263),
    .ZN(n1269)
  );
  AND2_X2 n_n543 (
    .A1(a_111_),
    .A2(b_111_),
    .Z(n1270)
  );
  AOI21_X1 n_n544 (
    .A1(n1253),
    .A2(n1254),
    .B(n1255),
    .ZN(n1261)
  );
  AND2_X2 n_n545 (
    .A1(a_110_),
    .A2(b_110_),
    .Z(n1262)
  );
  AOI21_X1 n_n546 (
    .A1(n1245),
    .A2(n1246),
    .B(n1247),
    .ZN(n1253)
  );
  AND2_X2 n_n547 (
    .A1(a_109_),
    .A2(b_109_),
    .Z(n1254)
  );
  AOI21_X1 n_n548 (
    .A1(n1237),
    .A2(n1238),
    .B(n1239),
    .ZN(n1245)
  );
  AND2_X2 n_n549 (
    .A1(a_108_),
    .A2(b_108_),
    .Z(n1246)
  );
  AOI21_X1 n_n550 (
    .A1(n1229),
    .A2(n1230),
    .B(n1231),
    .ZN(n1237)
  );
  AND2_X2 n_n551 (
    .A1(a_107_),
    .A2(b_107_),
    .Z(n1238)
  );
  AOI21_X1 n_n552 (
    .A1(n1221),
    .A2(n1222),
    .B(n1223),
    .ZN(n1229)
  );
  AND2_X2 n_n553 (
    .A1(a_106_),
    .A2(b_106_),
    .Z(n1230)
  );
  AOI21_X1 n_n554 (
    .A1(n1213),
    .A2(n1214),
    .B(n1215),
    .ZN(n1221)
  );
  AND2_X2 n_n555 (
    .A1(a_105_),
    .A2(b_105_),
    .Z(n1222)
  );
  AOI21_X1 n_n556 (
    .A1(n1205),
    .A2(n1206),
    .B(n1207),
    .ZN(n1213)
  );
  AND2_X2 n_n557 (
    .A1(a_104_),
    .A2(b_104_),
    .Z(n1214)
  );
  AOI21_X1 n_n558 (
    .A1(n1197),
    .A2(n1198),
    .B(n1199),
    .ZN(n1205)
  );
  AND2_X2 n_n559 (
    .A1(a_103_),
    .A2(b_103_),
    .Z(n1206)
  );
  AOI21_X1 n_n560 (
    .A1(n1189),
    .A2(n1190),
    .B(n1191),
    .ZN(n1197)
  );
  AND2_X2 n_n561 (
    .A1(a_102_),
    .A2(b_102_),
    .Z(n1198)
  );
  AOI21_X1 n_n562 (
    .A1(n1181),
    .A2(n1182),
    .B(n1183),
    .ZN(n1189)
  );
  AND2_X2 n_n563 (
    .A1(a_101_),
    .A2(b_101_),
    .Z(n1190)
  );
  AOI21_X1 n_n564 (
    .A1(n1173),
    .A2(n1174),
    .B(n1175),
    .ZN(n1181)
  );
  AND2_X2 n_n565 (
    .A1(a_100_),
    .A2(b_100_),
    .Z(n1182)
  );
  AOI21_X1 n_n566 (
    .A1(n1165),
    .A2(n1166),
    .B(n1167),
    .ZN(n1173)
  );
  AND2_X2 n_n567 (
    .A1(a_99_),
    .A2(b_99_),
    .Z(n1174)
  );
  AOI21_X1 n_n568 (
    .A1(n1157),
    .A2(n1158),
    .B(n1159),
    .ZN(n1165)
  );
  AND2_X2 n_n569 (
    .A1(a_98_),
    .A2(b_98_),
    .Z(n1166)
  );
  AOI21_X1 n_n570 (
    .A1(n1149),
    .A2(n1150),
    .B(n1151),
    .ZN(n1157)
  );
  AND2_X2 n_n571 (
    .A1(a_97_),
    .A2(b_97_),
    .Z(n1158)
  );
  AOI21_X1 n_n572 (
    .A1(n1141),
    .A2(n1142),
    .B(n1143),
    .ZN(n1149)
  );
  AND2_X2 n_n573 (
    .A1(a_96_),
    .A2(b_96_),
    .Z(n1150)
  );
  AOI21_X1 n_n574 (
    .A1(n1133),
    .A2(n1134),
    .B(n1135),
    .ZN(n1141)
  );
  AND2_X2 n_n575 (
    .A1(a_95_),
    .A2(b_95_),
    .Z(n1142)
  );
  AOI21_X1 n_n576 (
    .A1(n1125),
    .A2(n1126),
    .B(n1127),
    .ZN(n1133)
  );
  AND2_X2 n_n577 (
    .A1(a_94_),
    .A2(b_94_),
    .Z(n1134)
  );
  AOI21_X1 n_n578 (
    .A1(n1117),
    .A2(n1118),
    .B(n1119),
    .ZN(n1125)
  );
  AND2_X2 n_n579 (
    .A1(a_93_),
    .A2(b_93_),
    .Z(n1126)
  );
  AOI21_X1 n_n580 (
    .A1(n1109),
    .A2(n1110),
    .B(n1111),
    .ZN(n1117)
  );
  AND2_X2 n_n581 (
    .A1(a_92_),
    .A2(b_92_),
    .Z(n1118)
  );
  AOI21_X1 n_n582 (
    .A1(n1101),
    .A2(n1102),
    .B(n1103),
    .ZN(n1109)
  );
  AND2_X2 n_n583 (
    .A1(a_91_),
    .A2(b_91_),
    .Z(n1110)
  );
  AOI21_X1 n_n584 (
    .A1(n1093),
    .A2(n1094),
    .B(n1095),
    .ZN(n1101)
  );
  AND2_X2 n_n585 (
    .A1(a_90_),
    .A2(b_90_),
    .Z(n1102)
  );
  AOI21_X1 n_n586 (
    .A1(n1085),
    .A2(n1086),
    .B(n1087),
    .ZN(n1093)
  );
  AND2_X2 n_n587 (
    .A1(a_89_),
    .A2(b_89_),
    .Z(n1094)
  );
  AOI21_X1 n_n588 (
    .A1(n1077),
    .A2(n1078),
    .B(n1079),
    .ZN(n1085)
  );
  AND2_X2 n_n589 (
    .A1(a_88_),
    .A2(b_88_),
    .Z(n1086)
  );
  AOI21_X1 n_n590 (
    .A1(n1069),
    .A2(n1070),
    .B(n1071),
    .ZN(n1077)
  );
  AND2_X2 n_n591 (
    .A1(a_87_),
    .A2(b_87_),
    .Z(n1078)
  );
  AOI21_X1 n_n592 (
    .A1(n1061),
    .A2(n1062),
    .B(n1063),
    .ZN(n1069)
  );
  AND2_X2 n_n593 (
    .A1(a_86_),
    .A2(b_86_),
    .Z(n1070)
  );
  AOI21_X1 n_n594 (
    .A1(n1053),
    .A2(n1054),
    .B(n1055),
    .ZN(n1061)
  );
  AND2_X2 n_n595 (
    .A1(a_85_),
    .A2(b_85_),
    .Z(n1062)
  );
  AOI21_X1 n_n596 (
    .A1(n1045),
    .A2(n1046),
    .B(n1047),
    .ZN(n1053)
  );
  AND2_X2 n_n597 (
    .A1(a_84_),
    .A2(b_84_),
    .Z(n1054)
  );
  AOI21_X1 n_n598 (
    .A1(n1037),
    .A2(n1038),
    .B(n1039),
    .ZN(n1045)
  );
  AND2_X2 n_n599 (
    .A1(a_83_),
    .A2(b_83_),
    .Z(n1046)
  );
  AOI21_X1 n_n600 (
    .A1(n1029),
    .A2(n1030),
    .B(n1031),
    .ZN(n1037)
  );
  AND2_X2 n_n601 (
    .A1(a_82_),
    .A2(b_82_),
    .Z(n1038)
  );
  AOI21_X1 n_n602 (
    .A1(n1021),
    .A2(n1022),
    .B(n1023),
    .ZN(n1029)
  );
  AND2_X2 n_n603 (
    .A1(a_81_),
    .A2(b_81_),
    .Z(n1030)
  );
  AOI21_X1 n_n604 (
    .A1(n1013),
    .A2(n1014),
    .B(n1015),
    .ZN(n1021)
  );
  AND2_X2 n_n605 (
    .A1(a_80_),
    .A2(b_80_),
    .Z(n1022)
  );
  AOI21_X1 n_n606 (
    .A1(n1005),
    .A2(n1006),
    .B(n1007),
    .ZN(n1013)
  );
  AND2_X2 n_n607 (
    .A1(a_79_),
    .A2(b_79_),
    .Z(n1014)
  );
  AOI21_X1 n_n608 (
    .A1(n997),
    .A2(n998),
    .B(n999),
    .ZN(n1005)
  );
  AND2_X2 n_n609 (
    .A1(a_78_),
    .A2(b_78_),
    .Z(n1006)
  );
  AOI21_X1 n_n610 (
    .A1(n989),
    .A2(n990),
    .B(n991),
    .ZN(n997)
  );
  AND2_X2 n_n611 (
    .A1(a_77_),
    .A2(b_77_),
    .Z(n998)
  );
  AOI21_X1 n_n612 (
    .A1(n981),
    .A2(n982),
    .B(n983),
    .ZN(n989)
  );
  AND2_X2 n_n613 (
    .A1(a_76_),
    .A2(b_76_),
    .Z(n990)
  );
  AOI21_X1 n_n614 (
    .A1(n973),
    .A2(n974),
    .B(n975),
    .ZN(n981)
  );
  AND2_X2 n_n615 (
    .A1(a_75_),
    .A2(b_75_),
    .Z(n982)
  );
  AOI21_X1 n_n616 (
    .A1(n965),
    .A2(n966),
    .B(n967),
    .ZN(n973)
  );
  AND2_X2 n_n617 (
    .A1(a_74_),
    .A2(b_74_),
    .Z(n974)
  );
  AOI21_X1 n_n618 (
    .A1(n957),
    .A2(n958),
    .B(n959),
    .ZN(n965)
  );
  AND2_X2 n_n619 (
    .A1(a_73_),
    .A2(b_73_),
    .Z(n966)
  );
  AOI21_X1 n_n620 (
    .A1(n949),
    .A2(n950),
    .B(n951),
    .ZN(n957)
  );
  AND2_X2 n_n621 (
    .A1(a_72_),
    .A2(b_72_),
    .Z(n958)
  );
  AOI21_X1 n_n622 (
    .A1(n941),
    .A2(n942),
    .B(n943),
    .ZN(n949)
  );
  AND2_X2 n_n623 (
    .A1(a_71_),
    .A2(b_71_),
    .Z(n950)
  );
  AOI21_X1 n_n624 (
    .A1(n933),
    .A2(n934),
    .B(n935),
    .ZN(n941)
  );
  AND2_X2 n_n625 (
    .A1(a_70_),
    .A2(b_70_),
    .Z(n942)
  );
  AOI21_X1 n_n626 (
    .A1(n925),
    .A2(n926),
    .B(n927),
    .ZN(n933)
  );
  AND2_X2 n_n627 (
    .A1(a_69_),
    .A2(b_69_),
    .Z(n934)
  );
  AOI21_X1 n_n628 (
    .A1(n917),
    .A2(n918),
    .B(n919),
    .ZN(n925)
  );
  AND2_X2 n_n629 (
    .A1(a_68_),
    .A2(b_68_),
    .Z(n926)
  );
  AOI21_X1 n_n630 (
    .A1(n909),
    .A2(n910),
    .B(n911),
    .ZN(n917)
  );
  AND2_X2 n_n631 (
    .A1(a_67_),
    .A2(b_67_),
    .Z(n918)
  );
  AOI21_X1 n_n632 (
    .A1(n901),
    .A2(n902),
    .B(n903),
    .ZN(n909)
  );
  AND2_X2 n_n633 (
    .A1(a_66_),
    .A2(b_66_),
    .Z(n910)
  );
  AOI21_X1 n_n634 (
    .A1(n893),
    .A2(n894),
    .B(n895),
    .ZN(n901)
  );
  AND2_X2 n_n635 (
    .A1(a_65_),
    .A2(b_65_),
    .Z(n902)
  );
  AOI21_X1 n_n636 (
    .A1(n885),
    .A2(n886),
    .B(n887),
    .ZN(n893)
  );
  AND2_X2 n_n637 (
    .A1(a_64_),
    .A2(b_64_),
    .Z(n894)
  );
  AOI21_X1 n_n638 (
    .A1(n877),
    .A2(n878),
    .B(n879),
    .ZN(n885)
  );
  AND2_X2 n_n639 (
    .A1(a_63_),
    .A2(b_63_),
    .Z(n886)
  );
  AOI21_X1 n_n640 (
    .A1(n869),
    .A2(n870),
    .B(n871),
    .ZN(n877)
  );
  AND2_X2 n_n641 (
    .A1(a_62_),
    .A2(b_62_),
    .Z(n878)
  );
  AOI21_X1 n_n642 (
    .A1(n861),
    .A2(n862),
    .B(n863),
    .ZN(n869)
  );
  AND2_X2 n_n643 (
    .A1(a_61_),
    .A2(b_61_),
    .Z(n870)
  );
  AOI21_X1 n_n644 (
    .A1(n853),
    .A2(n854),
    .B(n855),
    .ZN(n861)
  );
  AND2_X2 n_n645 (
    .A1(a_60_),
    .A2(b_60_),
    .Z(n862)
  );
  AOI21_X1 n_n646 (
    .A1(n845),
    .A2(n846),
    .B(n847),
    .ZN(n853)
  );
  AND2_X2 n_n647 (
    .A1(a_59_),
    .A2(b_59_),
    .Z(n854)
  );
  AOI21_X1 n_n648 (
    .A1(n837),
    .A2(n838),
    .B(n839),
    .ZN(n845)
  );
  AND2_X2 n_n649 (
    .A1(a_58_),
    .A2(b_58_),
    .Z(n846)
  );
  AOI21_X1 n_n650 (
    .A1(n829),
    .A2(n830),
    .B(n831),
    .ZN(n837)
  );
  AND2_X2 n_n651 (
    .A1(a_57_),
    .A2(b_57_),
    .Z(n838)
  );
  AOI21_X1 n_n652 (
    .A1(n821),
    .A2(n822),
    .B(n823),
    .ZN(n829)
  );
  AND2_X2 n_n653 (
    .A1(a_56_),
    .A2(b_56_),
    .Z(n830)
  );
  AOI21_X1 n_n654 (
    .A1(n813),
    .A2(n814),
    .B(n815),
    .ZN(n821)
  );
  AND2_X2 n_n655 (
    .A1(a_55_),
    .A2(b_55_),
    .Z(n822)
  );
  AOI21_X1 n_n656 (
    .A1(n805),
    .A2(n806),
    .B(n807),
    .ZN(n813)
  );
  AND2_X2 n_n657 (
    .A1(a_54_),
    .A2(b_54_),
    .Z(n814)
  );
  AOI21_X1 n_n658 (
    .A1(n797),
    .A2(n798),
    .B(n799),
    .ZN(n805)
  );
  AND2_X2 n_n659 (
    .A1(a_53_),
    .A2(b_53_),
    .Z(n806)
  );
  AOI21_X1 n_n660 (
    .A1(n789),
    .A2(n790),
    .B(n791),
    .ZN(n797)
  );
  AND2_X2 n_n661 (
    .A1(a_52_),
    .A2(b_52_),
    .Z(n798)
  );
  AOI21_X1 n_n662 (
    .A1(n781),
    .A2(n782),
    .B(n783),
    .ZN(n789)
  );
  AND2_X2 n_n663 (
    .A1(a_51_),
    .A2(b_51_),
    .Z(n790)
  );
  AOI21_X1 n_n664 (
    .A1(n773),
    .A2(n774),
    .B(n775),
    .ZN(n781)
  );
  AND2_X2 n_n665 (
    .A1(a_50_),
    .A2(b_50_),
    .Z(n782)
  );
  AOI21_X1 n_n666 (
    .A1(n765),
    .A2(n766),
    .B(n767),
    .ZN(n773)
  );
  AND2_X2 n_n667 (
    .A1(a_49_),
    .A2(b_49_),
    .Z(n774)
  );
  AOI21_X1 n_n668 (
    .A1(n757),
    .A2(n758),
    .B(n759),
    .ZN(n765)
  );
  AND2_X2 n_n669 (
    .A1(a_48_),
    .A2(b_48_),
    .Z(n766)
  );
  AOI21_X1 n_n670 (
    .A1(n749),
    .A2(n750),
    .B(n751),
    .ZN(n757)
  );
  AND2_X2 n_n671 (
    .A1(a_47_),
    .A2(b_47_),
    .Z(n758)
  );
  AOI21_X1 n_n672 (
    .A1(n741),
    .A2(n742),
    .B(n743),
    .ZN(n749)
  );
  AND2_X2 n_n673 (
    .A1(a_46_),
    .A2(b_46_),
    .Z(n750)
  );
  AOI21_X1 n_n674 (
    .A1(n733),
    .A2(n734),
    .B(n735),
    .ZN(n741)
  );
  AND2_X2 n_n675 (
    .A1(a_45_),
    .A2(b_45_),
    .Z(n742)
  );
  AOI21_X1 n_n676 (
    .A1(n725),
    .A2(n726),
    .B(n727),
    .ZN(n733)
  );
  AND2_X2 n_n677 (
    .A1(a_44_),
    .A2(b_44_),
    .Z(n734)
  );
  AOI21_X1 n_n678 (
    .A1(n717),
    .A2(n718),
    .B(n719),
    .ZN(n725)
  );
  AND2_X2 n_n679 (
    .A1(a_43_),
    .A2(b_43_),
    .Z(n726)
  );
  AOI21_X1 n_n680 (
    .A1(n709),
    .A2(n710),
    .B(n711),
    .ZN(n717)
  );
  AND2_X2 n_n681 (
    .A1(a_42_),
    .A2(b_42_),
    .Z(n718)
  );
  AOI21_X1 n_n682 (
    .A1(n701),
    .A2(n702),
    .B(n703),
    .ZN(n709)
  );
  AND2_X2 n_n683 (
    .A1(a_41_),
    .A2(b_41_),
    .Z(n710)
  );
  AOI21_X1 n_n684 (
    .A1(n693),
    .A2(n694),
    .B(n695),
    .ZN(n701)
  );
  AND2_X2 n_n685 (
    .A1(a_40_),
    .A2(b_40_),
    .Z(n702)
  );
  AOI21_X1 n_n686 (
    .A1(n685),
    .A2(n686),
    .B(n687),
    .ZN(n693)
  );
  AND2_X2 n_n687 (
    .A1(a_39_),
    .A2(b_39_),
    .Z(n694)
  );
  AOI21_X1 n_n688 (
    .A1(n677),
    .A2(n678),
    .B(n679),
    .ZN(n685)
  );
  AND2_X2 n_n689 (
    .A1(a_38_),
    .A2(b_38_),
    .Z(n686)
  );
  AOI21_X1 n_n690 (
    .A1(n669),
    .A2(n670),
    .B(n671),
    .ZN(n677)
  );
  AND2_X2 n_n691 (
    .A1(a_37_),
    .A2(b_37_),
    .Z(n678)
  );
  AOI21_X1 n_n692 (
    .A1(n661),
    .A2(n662),
    .B(n663),
    .ZN(n669)
  );
  AND2_X2 n_n693 (
    .A1(a_36_),
    .A2(b_36_),
    .Z(n670)
  );
  AOI21_X1 n_n694 (
    .A1(n653),
    .A2(n654),
    .B(n655),
    .ZN(n661)
  );
  AND2_X2 n_n695 (
    .A1(a_35_),
    .A2(b_35_),
    .Z(n662)
  );
  AOI21_X1 n_n696 (
    .A1(n645),
    .A2(n646),
    .B(n647),
    .ZN(n653)
  );
  AND2_X2 n_n697 (
    .A1(a_34_),
    .A2(b_34_),
    .Z(n654)
  );
  AOI21_X1 n_n698 (
    .A1(n637),
    .A2(n638),
    .B(n639),
    .ZN(n645)
  );
  AND2_X2 n_n699 (
    .A1(a_33_),
    .A2(b_33_),
    .Z(n646)
  );
  AOI21_X1 n_n700 (
    .A1(n629),
    .A2(n630),
    .B(n631),
    .ZN(n637)
  );
  AND2_X2 n_n701 (
    .A1(a_32_),
    .A2(b_32_),
    .Z(n638)
  );
  AOI21_X1 n_n702 (
    .A1(n621),
    .A2(n622),
    .B(n623),
    .ZN(n629)
  );
  AND2_X2 n_n703 (
    .A1(a_31_),
    .A2(b_31_),
    .Z(n630)
  );
  AOI21_X1 n_n704 (
    .A1(n613),
    .A2(n614),
    .B(n615),
    .ZN(n621)
  );
  AND2_X2 n_n705 (
    .A1(a_30_),
    .A2(b_30_),
    .Z(n622)
  );
  AOI21_X1 n_n706 (
    .A1(n605),
    .A2(n606),
    .B(n607),
    .ZN(n613)
  );
  AND2_X2 n_n707 (
    .A1(a_29_),
    .A2(b_29_),
    .Z(n614)
  );
  AOI21_X1 n_n708 (
    .A1(n597),
    .A2(n598),
    .B(n599),
    .ZN(n605)
  );
  AND2_X2 n_n709 (
    .A1(a_28_),
    .A2(b_28_),
    .Z(n606)
  );
  AOI21_X1 n_n710 (
    .A1(n589),
    .A2(n590),
    .B(n591),
    .ZN(n597)
  );
  AND2_X2 n_n711 (
    .A1(a_27_),
    .A2(b_27_),
    .Z(n598)
  );
  AOI21_X1 n_n712 (
    .A1(n581),
    .A2(n582),
    .B(n583),
    .ZN(n589)
  );
  AND2_X2 n_n713 (
    .A1(a_26_),
    .A2(b_26_),
    .Z(n590)
  );
  AOI21_X1 n_n714 (
    .A1(n573),
    .A2(n574),
    .B(n575),
    .ZN(n581)
  );
  AND2_X2 n_n715 (
    .A1(a_25_),
    .A2(b_25_),
    .Z(n582)
  );
  AOI21_X1 n_n716 (
    .A1(n565),
    .A2(n566),
    .B(n567),
    .ZN(n573)
  );
  AND2_X2 n_n717 (
    .A1(a_24_),
    .A2(b_24_),
    .Z(n574)
  );
  AOI21_X1 n_n718 (
    .A1(n557),
    .A2(n558),
    .B(n559),
    .ZN(n565)
  );
  AND2_X2 n_n719 (
    .A1(a_23_),
    .A2(b_23_),
    .Z(n566)
  );
  AOI21_X1 n_n720 (
    .A1(n549),
    .A2(n550),
    .B(n551),
    .ZN(n557)
  );
  AND2_X2 n_n721 (
    .A1(a_22_),
    .A2(b_22_),
    .Z(n558)
  );
  AOI21_X1 n_n722 (
    .A1(n541),
    .A2(n542),
    .B(n543),
    .ZN(n549)
  );
  AND2_X2 n_n723 (
    .A1(a_21_),
    .A2(b_21_),
    .Z(n550)
  );
  AOI21_X1 n_n724 (
    .A1(n533),
    .A2(n534),
    .B(n535),
    .ZN(n541)
  );
  AND2_X2 n_n725 (
    .A1(a_20_),
    .A2(b_20_),
    .Z(n542)
  );
  AOI21_X1 n_n726 (
    .A1(n525),
    .A2(n526),
    .B(n527),
    .ZN(n533)
  );
  AND2_X2 n_n727 (
    .A1(a_19_),
    .A2(b_19_),
    .Z(n534)
  );
  AOI21_X1 n_n728 (
    .A1(n517),
    .A2(n518),
    .B(n519),
    .ZN(n525)
  );
  AND2_X2 n_n729 (
    .A1(a_18_),
    .A2(b_18_),
    .Z(n526)
  );
  AOI21_X1 n_n730 (
    .A1(n509),
    .A2(n510),
    .B(n511),
    .ZN(n517)
  );
  AND2_X2 n_n731 (
    .A1(a_17_),
    .A2(b_17_),
    .Z(n518)
  );
  AOI21_X1 n_n732 (
    .A1(n501),
    .A2(n502),
    .B(n503),
    .ZN(n509)
  );
  AND2_X2 n_n733 (
    .A1(a_16_),
    .A2(b_16_),
    .Z(n510)
  );
  AOI21_X1 n_n734 (
    .A1(n493),
    .A2(n494),
    .B(n495),
    .ZN(n501)
  );
  AND2_X2 n_n735 (
    .A1(a_15_),
    .A2(b_15_),
    .Z(n502)
  );
  AOI21_X1 n_n736 (
    .A1(n485),
    .A2(n486),
    .B(n487),
    .ZN(n493)
  );
  AND2_X2 n_n737 (
    .A1(a_14_),
    .A2(b_14_),
    .Z(n494)
  );
  AOI21_X1 n_n738 (
    .A1(n477),
    .A2(n478),
    .B(n479),
    .ZN(n485)
  );
  AND2_X2 n_n739 (
    .A1(a_13_),
    .A2(b_13_),
    .Z(n486)
  );
  AOI21_X1 n_n740 (
    .A1(n469),
    .A2(n470),
    .B(n471),
    .ZN(n477)
  );
  AND2_X2 n_n741 (
    .A1(a_12_),
    .A2(b_12_),
    .Z(n478)
  );
  AOI21_X1 n_n742 (
    .A1(n461),
    .A2(n462),
    .B(n463),
    .ZN(n469)
  );
  AND2_X2 n_n743 (
    .A1(a_11_),
    .A2(b_11_),
    .Z(n470)
  );
  AOI21_X1 n_n744 (
    .A1(n453),
    .A2(n454),
    .B(n455),
    .ZN(n461)
  );
  AND2_X2 n_n745 (
    .A1(a_10_),
    .A2(b_10_),
    .Z(n462)
  );
  AOI21_X1 n_n746 (
    .A1(n445),
    .A2(n446),
    .B(n447),
    .ZN(n453)
  );
  AND2_X2 n_n747 (
    .A1(a_9_),
    .A2(b_9_),
    .Z(n454)
  );
  AOI21_X1 n_n748 (
    .A1(n437),
    .A2(n438),
    .B(n439),
    .ZN(n445)
  );
  AND2_X2 n_n749 (
    .A1(a_8_),
    .A2(b_8_),
    .Z(n446)
  );
  AOI21_X1 n_n750 (
    .A1(n429),
    .A2(n430),
    .B(n431),
    .ZN(n437)
  );
  AND2_X2 n_n751 (
    .A1(a_7_),
    .A2(b_7_),
    .Z(n438)
  );
  AOI21_X1 n_n752 (
    .A1(n421),
    .A2(n422),
    .B(n423),
    .ZN(n429)
  );
  AND2_X2 n_n753 (
    .A1(a_6_),
    .A2(b_6_),
    .Z(n430)
  );
  AOI21_X1 n_n754 (
    .A1(n413),
    .A2(n414),
    .B(n415),
    .ZN(n421)
  );
  AND2_X2 n_n755 (
    .A1(a_5_),
    .A2(b_5_),
    .Z(n422)
  );
  AOI21_X1 n_n756 (
    .A1(n405),
    .A2(n406),
    .B(n407),
    .ZN(n413)
  );
  AND2_X2 n_n757 (
    .A1(a_4_),
    .A2(b_4_),
    .Z(n414)
  );
  AOI21_X1 n_n758 (
    .A1(n397),
    .A2(n398),
    .B(n399),
    .ZN(n405)
  );
  AND2_X2 n_n759 (
    .A1(a_3_),
    .A2(b_3_),
    .Z(n406)
  );
  AOI21_X1 n_n760 (
    .A1(n389),
    .A2(n390),
    .B(n391),
    .ZN(n397)
  );
  AND2_X2 n_n761 (
    .A1(a_2_),
    .A2(b_2_),
    .Z(n398)
  );
  AND2_X2 n_n762 (
    .A1(a_0_),
    .A2(b_0_),
    .Z(n389)
  );
endmodule
