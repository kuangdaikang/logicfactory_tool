// Benchmark "dalu" written by ABC on Fri Feb 25 15:12:52 2022

module dalu ( 
    inA15, inA14, inA13, inA12, inA11, inA10, inA9, inA8, inA7, inA6, inA5,
    inA4, inA3, inA2, inA1, inA0, inB15, inB14, inB13, inB12, inB11, inB10,
    inB9, inB8, inB7, inB6, inB5, inB4, inB3, inB2, inB1, inB0, inC15,
    inC14, inC13, inC12, inC11, inC10, inC9, inC8, inC7, inC6, inC5, inC4,
    inC3, inC2, inC1, inC0, inD15, inD14, inD13, inD12, inD11, inD10, inD9,
    inD8, inD7, inD6, inD5, inD4, inD3, inD2, inD1, inD0, opsel3, opsel2,
    opsel1, opsel0, musel4, musel3, musel2, musel1, sh2, sh1, sh0,
    O15, O14, O13, O12, O11, O10, O9, O8, O7, O6, O5, O4, O3, O2, O1, O0  );
  input  inA15, inA14, inA13, inA12, inA11, inA10, inA9, inA8, inA7,
    inA6, inA5, inA4, inA3, inA2, inA1, inA0, inB15, inB14, inB13, inB12,
    inB11, inB10, inB9, inB8, inB7, inB6, inB5, inB4, inB3, inB2, inB1,
    inB0, inC15, inC14, inC13, inC12, inC11, inC10, inC9, inC8, inC7, inC6,
    inC5, inC4, inC3, inC2, inC1, inC0, inD15, inD14, inD13, inD12, inD11,
    inD10, inD9, inD8, inD7, inD6, inD5, inD4, inD3, inD2, inD1, inD0,
    opsel3, opsel2, opsel1, opsel0, musel4, musel3, musel2, musel1, sh2,
    sh1, sh0;
  output O15, O14, O13, O12, O11, O10, O9, O8, O7, O6, O5, O4, O3, O2, O1, O0;
  wire new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_;
  assign new_n92_ = ~opsel1 & ~opsel0;
  assign new_n93_ = inC14 & musel2;
  assign new_n94_ = ~musel2 & musel1;
  assign new_n95_ = inA14 & new_n94_;
  assign new_n96_ = ~musel1 & new_n93_;
  assign new_n97_ = ~new_n95_ & ~new_n96_;
  assign new_n98_ = ~musel3 & ~new_n97_;
  assign new_n99_ = musel4 & new_n98_;
  assign new_n100_ = inC15 & musel2;
  assign new_n101_ = inA15 & new_n94_;
  assign new_n102_ = ~musel1 & new_n100_;
  assign new_n103_ = ~new_n101_ & ~new_n102_;
  assign new_n104_ = ~musel3 & ~new_n103_;
  assign new_n105_ = musel4 & new_n104_;
  assign new_n106_ = ~new_n99_ & new_n105_;
  assign new_n107_ = new_n99_ & ~new_n105_;
  assign new_n108_ = ~new_n106_ & ~new_n107_;
  assign new_n109_ = inC13 & musel2;
  assign new_n110_ = inA13 & new_n94_;
  assign new_n111_ = ~musel1 & new_n109_;
  assign new_n112_ = ~new_n110_ & ~new_n111_;
  assign new_n113_ = ~musel3 & ~new_n112_;
  assign new_n114_ = musel4 & new_n113_;
  assign new_n115_ = new_n105_ & ~new_n114_;
  assign new_n116_ = ~new_n105_ & new_n114_;
  assign new_n117_ = ~new_n115_ & ~new_n116_;
  assign new_n118_ = inC12 & musel2;
  assign new_n119_ = inA12 & new_n94_;
  assign new_n120_ = ~musel1 & new_n118_;
  assign new_n121_ = ~new_n119_ & ~new_n120_;
  assign new_n122_ = ~musel3 & ~new_n121_;
  assign new_n123_ = musel4 & new_n122_;
  assign new_n124_ = new_n105_ & ~new_n123_;
  assign new_n125_ = ~new_n105_ & new_n123_;
  assign new_n126_ = ~new_n124_ & ~new_n125_;
  assign new_n127_ = inC7 & musel2;
  assign new_n128_ = inA7 & new_n94_;
  assign new_n129_ = ~musel1 & new_n127_;
  assign new_n130_ = ~new_n128_ & ~new_n129_;
  assign new_n131_ = ~musel3 & ~new_n130_;
  assign new_n132_ = musel4 & new_n131_;
  assign new_n133_ = new_n105_ & ~new_n132_;
  assign new_n134_ = ~new_n105_ & new_n132_;
  assign new_n135_ = ~new_n133_ & ~new_n134_;
  assign new_n136_ = inC6 & musel2;
  assign new_n137_ = inA6 & new_n94_;
  assign new_n138_ = ~musel1 & new_n136_;
  assign new_n139_ = ~new_n137_ & ~new_n138_;
  assign new_n140_ = ~musel3 & ~new_n139_;
  assign new_n141_ = musel4 & new_n140_;
  assign new_n142_ = new_n105_ & ~new_n141_;
  assign new_n143_ = ~new_n105_ & new_n141_;
  assign new_n144_ = ~new_n142_ & ~new_n143_;
  assign new_n145_ = inC5 & musel2;
  assign new_n146_ = inA5 & new_n94_;
  assign new_n147_ = ~musel1 & new_n145_;
  assign new_n148_ = ~new_n146_ & ~new_n147_;
  assign new_n149_ = ~musel3 & ~new_n148_;
  assign new_n150_ = musel4 & new_n149_;
  assign new_n151_ = new_n105_ & ~new_n150_;
  assign new_n152_ = ~new_n105_ & new_n150_;
  assign new_n153_ = ~new_n151_ & ~new_n152_;
  assign new_n154_ = inC4 & musel2;
  assign new_n155_ = inA4 & new_n94_;
  assign new_n156_ = ~musel1 & new_n154_;
  assign new_n157_ = ~new_n155_ & ~new_n156_;
  assign new_n158_ = ~musel3 & ~new_n157_;
  assign new_n159_ = musel4 & new_n158_;
  assign new_n160_ = new_n105_ & ~new_n159_;
  assign new_n161_ = ~new_n105_ & new_n159_;
  assign new_n162_ = ~new_n160_ & ~new_n161_;
  assign new_n163_ = ~new_n135_ & ~new_n144_;
  assign new_n164_ = ~new_n153_ & ~new_n162_;
  assign new_n165_ = new_n163_ & new_n164_;
  assign new_n166_ = inC11 & musel2;
  assign new_n167_ = inA11 & new_n94_;
  assign new_n168_ = ~musel1 & new_n166_;
  assign new_n169_ = ~new_n167_ & ~new_n168_;
  assign new_n170_ = ~musel3 & ~new_n169_;
  assign new_n171_ = musel4 & new_n170_;
  assign new_n172_ = new_n105_ & ~new_n171_;
  assign new_n173_ = ~new_n105_ & new_n171_;
  assign new_n174_ = ~new_n172_ & ~new_n173_;
  assign new_n175_ = inC10 & musel2;
  assign new_n176_ = inA10 & new_n94_;
  assign new_n177_ = ~musel1 & new_n175_;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign new_n179_ = ~musel3 & ~new_n178_;
  assign new_n180_ = musel4 & new_n179_;
  assign new_n181_ = new_n105_ & ~new_n180_;
  assign new_n182_ = ~new_n105_ & new_n180_;
  assign new_n183_ = ~new_n181_ & ~new_n182_;
  assign new_n184_ = inC9 & musel2;
  assign new_n185_ = inA9 & new_n94_;
  assign new_n186_ = ~musel1 & new_n184_;
  assign new_n187_ = ~new_n185_ & ~new_n186_;
  assign new_n188_ = ~musel3 & ~new_n187_;
  assign new_n189_ = musel4 & new_n188_;
  assign new_n190_ = new_n105_ & ~new_n189_;
  assign new_n191_ = ~new_n105_ & new_n189_;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign new_n193_ = inC8 & musel2;
  assign new_n194_ = inA8 & new_n94_;
  assign new_n195_ = ~musel1 & new_n193_;
  assign new_n196_ = ~new_n194_ & ~new_n195_;
  assign new_n197_ = ~musel3 & ~new_n196_;
  assign new_n198_ = musel4 & new_n197_;
  assign new_n199_ = new_n105_ & ~new_n198_;
  assign new_n200_ = ~new_n105_ & new_n198_;
  assign new_n201_ = ~new_n199_ & ~new_n200_;
  assign new_n202_ = ~new_n174_ & ~new_n183_;
  assign new_n203_ = ~new_n192_ & ~new_n201_;
  assign new_n204_ = new_n202_ & new_n203_;
  assign new_n205_ = inC3 & musel2;
  assign new_n206_ = inA3 & new_n94_;
  assign new_n207_ = ~musel1 & new_n205_;
  assign new_n208_ = ~new_n206_ & ~new_n207_;
  assign new_n209_ = ~musel3 & ~new_n208_;
  assign new_n210_ = musel4 & new_n209_;
  assign new_n211_ = new_n105_ & ~new_n210_;
  assign new_n212_ = ~new_n105_ & new_n210_;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = inC2 & musel2;
  assign new_n215_ = inA2 & new_n94_;
  assign new_n216_ = ~musel1 & new_n214_;
  assign new_n217_ = ~new_n215_ & ~new_n216_;
  assign new_n218_ = ~musel3 & ~new_n217_;
  assign new_n219_ = musel4 & new_n218_;
  assign new_n220_ = new_n105_ & ~new_n219_;
  assign new_n221_ = ~new_n105_ & new_n219_;
  assign new_n222_ = ~new_n220_ & ~new_n221_;
  assign new_n223_ = inC1 & musel2;
  assign new_n224_ = inA1 & new_n94_;
  assign new_n225_ = ~musel1 & new_n223_;
  assign new_n226_ = ~new_n224_ & ~new_n225_;
  assign new_n227_ = ~musel3 & ~new_n226_;
  assign new_n228_ = musel4 & new_n227_;
  assign new_n229_ = new_n105_ & ~new_n228_;
  assign new_n230_ = ~new_n105_ & new_n228_;
  assign new_n231_ = ~new_n229_ & ~new_n230_;
  assign new_n232_ = inC0 & musel2;
  assign new_n233_ = inA0 & new_n94_;
  assign new_n234_ = ~musel1 & new_n232_;
  assign new_n235_ = ~new_n233_ & ~new_n234_;
  assign new_n236_ = ~musel3 & ~new_n235_;
  assign new_n237_ = musel4 & new_n236_;
  assign new_n238_ = new_n105_ & ~new_n237_;
  assign new_n239_ = ~new_n105_ & new_n237_;
  assign new_n240_ = ~new_n238_ & ~new_n239_;
  assign new_n241_ = ~new_n213_ & ~new_n222_;
  assign new_n242_ = ~new_n231_ & ~new_n240_;
  assign new_n243_ = new_n241_ & new_n242_;
  assign new_n244_ = new_n165_ & new_n204_;
  assign new_n245_ = new_n105_ & new_n244_;
  assign new_n246_ = new_n243_ & new_n245_;
  assign new_n247_ = ~new_n108_ & ~new_n117_;
  assign new_n248_ = ~new_n126_ & new_n246_;
  assign new_n249_ = new_n247_ & new_n248_;
  assign new_n250_ = inD15 & musel2;
  assign new_n251_ = musel2 & ~musel1;
  assign new_n252_ = ~new_n94_ & ~new_n251_;
  assign new_n253_ = musel1 & new_n250_;
  assign new_n254_ = inB15 & ~new_n252_;
  assign new_n255_ = ~new_n253_ & ~new_n254_;
  assign new_n256_ = ~musel4 & musel3;
  assign new_n257_ = ~musel2 & ~musel1;
  assign new_n258_ = ~musel3 & new_n257_;
  assign new_n259_ = inD15 & musel4;
  assign new_n260_ = new_n258_ & new_n259_;
  assign new_n261_ = ~new_n255_ & new_n256_;
  assign new_n262_ = ~new_n260_ & ~new_n261_;
  assign new_n263_ = opsel2 & ~new_n262_;
  assign new_n264_ = ~opsel2 & new_n249_;
  assign new_n265_ = ~new_n263_ & ~new_n264_;
  assign new_n266_ = opsel2 & new_n92_;
  assign new_n267_ = new_n249_ & new_n266_;
  assign new_n268_ = ~new_n92_ & ~new_n265_;
  assign new_n269_ = ~new_n267_ & ~new_n268_;
  assign new_n270_ = inA15 & ~musel2;
  assign new_n271_ = ~new_n100_ & ~new_n270_;
  assign new_n272_ = ~musel3 & ~new_n271_;
  assign new_n273_ = musel1 & new_n272_;
  assign new_n274_ = musel3 & ~musel2;
  assign new_n275_ = inD15 & new_n274_;
  assign new_n276_ = ~musel3 & musel2;
  assign new_n277_ = inB15 & new_n276_;
  assign new_n278_ = ~new_n275_ & ~new_n277_;
  assign new_n279_ = ~musel1 & ~new_n278_;
  assign new_n280_ = ~new_n273_ & ~new_n279_;
  assign new_n281_ = ~musel4 & ~new_n280_;
  assign new_n282_ = inC15 & musel4;
  assign new_n283_ = ~musel3 & new_n282_;
  assign new_n284_ = ~musel2 & new_n283_;
  assign new_n285_ = ~musel1 & new_n284_;
  assign new_n286_ = musel1 & new_n100_;
  assign new_n287_ = inA15 & ~new_n252_;
  assign new_n288_ = ~new_n286_ & ~new_n287_;
  assign new_n289_ = ~musel4 & ~new_n288_;
  assign new_n290_ = musel3 & new_n289_;
  assign new_n291_ = ~new_n285_ & ~new_n290_;
  assign new_n292_ = ~opsel3 & ~opsel1;
  assign new_n293_ = ~opsel2 & opsel1;
  assign new_n294_ = ~new_n292_ & ~new_n293_;
  assign new_n295_ = opsel3 & opsel2;
  assign new_n296_ = ~opsel0 & new_n294_;
  assign new_n297_ = ~new_n295_ & new_n296_;
  assign new_n298_ = new_n291_ & new_n297_;
  assign new_n299_ = ~new_n291_ & ~new_n297_;
  assign new_n300_ = ~new_n298_ & ~new_n299_;
  assign new_n301_ = ~new_n281_ & ~new_n300_;
  assign new_n302_ = new_n281_ & new_n300_;
  assign new_n303_ = ~new_n301_ & ~new_n302_;
  assign new_n304_ = inC14 & musel4;
  assign new_n305_ = ~musel3 & new_n304_;
  assign new_n306_ = ~musel2 & new_n305_;
  assign new_n307_ = ~musel1 & new_n306_;
  assign new_n308_ = musel1 & new_n93_;
  assign new_n309_ = inA14 & ~new_n252_;
  assign new_n310_ = ~new_n308_ & ~new_n309_;
  assign new_n311_ = ~musel4 & ~new_n310_;
  assign new_n312_ = musel3 & new_n311_;
  assign new_n313_ = ~new_n307_ & ~new_n312_;
  assign new_n314_ = new_n297_ & new_n313_;
  assign new_n315_ = ~new_n297_ & ~new_n313_;
  assign new_n316_ = ~new_n314_ & ~new_n315_;
  assign new_n317_ = inA14 & ~musel2;
  assign new_n318_ = ~new_n93_ & ~new_n317_;
  assign new_n319_ = ~musel3 & ~new_n318_;
  assign new_n320_ = musel1 & new_n319_;
  assign new_n321_ = inD14 & new_n274_;
  assign new_n322_ = inB14 & new_n276_;
  assign new_n323_ = ~new_n321_ & ~new_n322_;
  assign new_n324_ = ~musel1 & ~new_n323_;
  assign new_n325_ = ~new_n320_ & ~new_n324_;
  assign new_n326_ = ~musel4 & ~new_n325_;
  assign new_n327_ = ~new_n316_ & new_n326_;
  assign new_n328_ = inC13 & musel4;
  assign new_n329_ = ~musel3 & new_n328_;
  assign new_n330_ = ~musel2 & new_n329_;
  assign new_n331_ = ~musel1 & new_n330_;
  assign new_n332_ = musel1 & new_n109_;
  assign new_n333_ = inA13 & ~new_n252_;
  assign new_n334_ = ~new_n332_ & ~new_n333_;
  assign new_n335_ = ~musel4 & ~new_n334_;
  assign new_n336_ = musel3 & new_n335_;
  assign new_n337_ = ~new_n331_ & ~new_n336_;
  assign new_n338_ = new_n297_ & new_n337_;
  assign new_n339_ = ~new_n297_ & ~new_n337_;
  assign new_n340_ = ~new_n338_ & ~new_n339_;
  assign new_n341_ = inA13 & ~musel2;
  assign new_n342_ = ~new_n109_ & ~new_n341_;
  assign new_n343_ = ~musel3 & ~new_n342_;
  assign new_n344_ = musel1 & new_n343_;
  assign new_n345_ = inD13 & new_n274_;
  assign new_n346_ = inB13 & new_n276_;
  assign new_n347_ = ~new_n345_ & ~new_n346_;
  assign new_n348_ = ~musel1 & ~new_n347_;
  assign new_n349_ = ~new_n344_ & ~new_n348_;
  assign new_n350_ = ~musel4 & ~new_n349_;
  assign new_n351_ = ~new_n340_ & new_n350_;
  assign new_n352_ = inC12 & musel4;
  assign new_n353_ = ~musel3 & new_n352_;
  assign new_n354_ = ~musel2 & new_n353_;
  assign new_n355_ = ~musel1 & new_n354_;
  assign new_n356_ = musel1 & new_n118_;
  assign new_n357_ = inA12 & ~new_n252_;
  assign new_n358_ = ~new_n356_ & ~new_n357_;
  assign new_n359_ = ~musel4 & ~new_n358_;
  assign new_n360_ = musel3 & new_n359_;
  assign new_n361_ = ~new_n355_ & ~new_n360_;
  assign new_n362_ = new_n297_ & new_n361_;
  assign new_n363_ = ~new_n297_ & ~new_n361_;
  assign new_n364_ = ~new_n362_ & ~new_n363_;
  assign new_n365_ = inA12 & ~musel2;
  assign new_n366_ = ~new_n118_ & ~new_n365_;
  assign new_n367_ = ~musel3 & ~new_n366_;
  assign new_n368_ = musel1 & new_n367_;
  assign new_n369_ = inD12 & new_n274_;
  assign new_n370_ = inB12 & new_n276_;
  assign new_n371_ = ~new_n369_ & ~new_n370_;
  assign new_n372_ = ~musel1 & ~new_n371_;
  assign new_n373_ = ~new_n368_ & ~new_n372_;
  assign new_n374_ = ~musel4 & ~new_n373_;
  assign new_n375_ = ~new_n364_ & new_n374_;
  assign new_n376_ = ~opsel2 & ~opsel1;
  assign new_n377_ = opsel3 & new_n376_;
  assign new_n378_ = ~opsel3 & opsel1;
  assign new_n379_ = opsel2 & new_n378_;
  assign new_n380_ = ~new_n377_ & ~new_n379_;
  assign new_n381_ = ~opsel0 & ~new_n380_;
  assign new_n382_ = inA3 & ~musel2;
  assign new_n383_ = ~new_n205_ & ~new_n382_;
  assign new_n384_ = ~musel3 & ~new_n383_;
  assign new_n385_ = musel1 & new_n384_;
  assign new_n386_ = inD3 & new_n274_;
  assign new_n387_ = inB3 & new_n276_;
  assign new_n388_ = ~new_n386_ & ~new_n387_;
  assign new_n389_ = ~musel1 & ~new_n388_;
  assign new_n390_ = ~new_n385_ & ~new_n389_;
  assign new_n391_ = ~musel4 & ~new_n390_;
  assign new_n392_ = inC3 & musel4;
  assign new_n393_ = ~musel3 & new_n392_;
  assign new_n394_ = ~musel2 & new_n393_;
  assign new_n395_ = ~musel1 & new_n394_;
  assign new_n396_ = musel1 & new_n205_;
  assign new_n397_ = inA3 & ~new_n252_;
  assign new_n398_ = ~new_n396_ & ~new_n397_;
  assign new_n399_ = ~musel4 & ~new_n398_;
  assign new_n400_ = musel3 & new_n399_;
  assign new_n401_ = ~new_n395_ & ~new_n400_;
  assign new_n402_ = new_n297_ & new_n401_;
  assign new_n403_ = ~new_n297_ & ~new_n401_;
  assign new_n404_ = ~new_n402_ & ~new_n403_;
  assign new_n405_ = inA2 & ~musel2;
  assign new_n406_ = ~new_n214_ & ~new_n405_;
  assign new_n407_ = ~musel3 & ~new_n406_;
  assign new_n408_ = musel1 & new_n407_;
  assign new_n409_ = inD2 & new_n274_;
  assign new_n410_ = inB2 & new_n276_;
  assign new_n411_ = ~new_n409_ & ~new_n410_;
  assign new_n412_ = ~musel1 & ~new_n411_;
  assign new_n413_ = ~new_n408_ & ~new_n412_;
  assign new_n414_ = ~musel4 & ~new_n413_;
  assign new_n415_ = inC2 & musel4;
  assign new_n416_ = ~musel3 & new_n415_;
  assign new_n417_ = ~musel2 & new_n416_;
  assign new_n418_ = ~musel1 & new_n417_;
  assign new_n419_ = musel1 & new_n214_;
  assign new_n420_ = inA2 & ~new_n252_;
  assign new_n421_ = ~new_n419_ & ~new_n420_;
  assign new_n422_ = ~musel4 & ~new_n421_;
  assign new_n423_ = musel3 & new_n422_;
  assign new_n424_ = ~new_n418_ & ~new_n423_;
  assign new_n425_ = new_n297_ & new_n424_;
  assign new_n426_ = ~new_n297_ & ~new_n424_;
  assign new_n427_ = ~new_n425_ & ~new_n426_;
  assign new_n428_ = ~new_n391_ & new_n404_;
  assign new_n429_ = ~new_n414_ & new_n427_;
  assign new_n430_ = ~new_n428_ & ~new_n429_;
  assign new_n431_ = inA1 & ~musel2;
  assign new_n432_ = ~new_n223_ & ~new_n431_;
  assign new_n433_ = ~musel3 & ~new_n432_;
  assign new_n434_ = musel1 & new_n433_;
  assign new_n435_ = inD1 & new_n274_;
  assign new_n436_ = inB1 & new_n276_;
  assign new_n437_ = ~new_n435_ & ~new_n436_;
  assign new_n438_ = ~musel1 & ~new_n437_;
  assign new_n439_ = ~new_n434_ & ~new_n438_;
  assign new_n440_ = ~musel4 & ~new_n439_;
  assign new_n441_ = inC1 & musel4;
  assign new_n442_ = ~musel3 & new_n441_;
  assign new_n443_ = ~musel2 & new_n442_;
  assign new_n444_ = ~musel1 & new_n443_;
  assign new_n445_ = musel1 & new_n223_;
  assign new_n446_ = inA1 & ~new_n252_;
  assign new_n447_ = ~new_n445_ & ~new_n446_;
  assign new_n448_ = ~musel4 & ~new_n447_;
  assign new_n449_ = musel3 & new_n448_;
  assign new_n450_ = ~new_n444_ & ~new_n449_;
  assign new_n451_ = new_n297_ & new_n450_;
  assign new_n452_ = ~new_n297_ & ~new_n450_;
  assign new_n453_ = ~new_n451_ & ~new_n452_;
  assign new_n454_ = inA0 & ~musel2;
  assign new_n455_ = ~new_n232_ & ~new_n454_;
  assign new_n456_ = ~musel3 & ~new_n455_;
  assign new_n457_ = musel1 & new_n456_;
  assign new_n458_ = inD0 & new_n274_;
  assign new_n459_ = inB0 & new_n276_;
  assign new_n460_ = ~new_n458_ & ~new_n459_;
  assign new_n461_ = ~musel1 & ~new_n460_;
  assign new_n462_ = ~new_n457_ & ~new_n461_;
  assign new_n463_ = ~musel4 & ~new_n462_;
  assign new_n464_ = inC0 & musel4;
  assign new_n465_ = ~musel3 & new_n464_;
  assign new_n466_ = ~musel2 & new_n465_;
  assign new_n467_ = ~musel1 & new_n466_;
  assign new_n468_ = musel1 & new_n232_;
  assign new_n469_ = inA0 & ~new_n252_;
  assign new_n470_ = ~new_n468_ & ~new_n469_;
  assign new_n471_ = ~musel4 & ~new_n470_;
  assign new_n472_ = musel3 & new_n471_;
  assign new_n473_ = ~new_n467_ & ~new_n472_;
  assign new_n474_ = new_n297_ & new_n473_;
  assign new_n475_ = ~new_n297_ & ~new_n473_;
  assign new_n476_ = ~new_n474_ & ~new_n475_;
  assign new_n477_ = ~new_n440_ & new_n453_;
  assign new_n478_ = ~new_n463_ & new_n476_;
  assign new_n479_ = ~new_n477_ & ~new_n478_;
  assign new_n480_ = new_n430_ & new_n479_;
  assign new_n481_ = new_n381_ & new_n480_;
  assign new_n482_ = new_n463_ & ~new_n476_;
  assign new_n483_ = new_n440_ & ~new_n453_;
  assign new_n484_ = ~new_n477_ & new_n482_;
  assign new_n485_ = ~new_n483_ & ~new_n484_;
  assign new_n486_ = ~new_n429_ & ~new_n485_;
  assign new_n487_ = new_n414_ & ~new_n427_;
  assign new_n488_ = ~new_n486_ & ~new_n487_;
  assign new_n489_ = ~new_n428_ & ~new_n488_;
  assign new_n490_ = new_n391_ & ~new_n404_;
  assign new_n491_ = ~new_n489_ & ~new_n490_;
  assign new_n492_ = ~new_n481_ & new_n491_;
  assign new_n493_ = inA7 & ~musel2;
  assign new_n494_ = ~new_n127_ & ~new_n493_;
  assign new_n495_ = ~musel3 & ~new_n494_;
  assign new_n496_ = musel1 & new_n495_;
  assign new_n497_ = inD7 & new_n274_;
  assign new_n498_ = inB7 & new_n276_;
  assign new_n499_ = ~new_n497_ & ~new_n498_;
  assign new_n500_ = ~musel1 & ~new_n499_;
  assign new_n501_ = ~new_n496_ & ~new_n500_;
  assign new_n502_ = ~musel4 & ~new_n501_;
  assign new_n503_ = inC7 & musel4;
  assign new_n504_ = ~musel3 & new_n503_;
  assign new_n505_ = ~musel2 & new_n504_;
  assign new_n506_ = ~musel1 & new_n505_;
  assign new_n507_ = musel1 & new_n127_;
  assign new_n508_ = inA7 & ~new_n252_;
  assign new_n509_ = ~new_n507_ & ~new_n508_;
  assign new_n510_ = ~musel4 & ~new_n509_;
  assign new_n511_ = musel3 & new_n510_;
  assign new_n512_ = ~new_n506_ & ~new_n511_;
  assign new_n513_ = new_n297_ & new_n512_;
  assign new_n514_ = ~new_n297_ & ~new_n512_;
  assign new_n515_ = ~new_n513_ & ~new_n514_;
  assign new_n516_ = inA6 & ~musel2;
  assign new_n517_ = ~new_n136_ & ~new_n516_;
  assign new_n518_ = ~musel3 & ~new_n517_;
  assign new_n519_ = musel1 & new_n518_;
  assign new_n520_ = inD6 & new_n274_;
  assign new_n521_ = inB6 & new_n276_;
  assign new_n522_ = ~new_n520_ & ~new_n521_;
  assign new_n523_ = ~musel1 & ~new_n522_;
  assign new_n524_ = ~new_n519_ & ~new_n523_;
  assign new_n525_ = ~musel4 & ~new_n524_;
  assign new_n526_ = inC6 & musel4;
  assign new_n527_ = ~musel3 & new_n526_;
  assign new_n528_ = ~musel2 & new_n527_;
  assign new_n529_ = ~musel1 & new_n528_;
  assign new_n530_ = musel1 & new_n136_;
  assign new_n531_ = inA6 & ~new_n252_;
  assign new_n532_ = ~new_n530_ & ~new_n531_;
  assign new_n533_ = ~musel4 & ~new_n532_;
  assign new_n534_ = musel3 & new_n533_;
  assign new_n535_ = ~new_n529_ & ~new_n534_;
  assign new_n536_ = new_n297_ & new_n535_;
  assign new_n537_ = ~new_n297_ & ~new_n535_;
  assign new_n538_ = ~new_n536_ & ~new_n537_;
  assign new_n539_ = ~new_n502_ & new_n515_;
  assign new_n540_ = ~new_n525_ & new_n538_;
  assign new_n541_ = ~new_n539_ & ~new_n540_;
  assign new_n542_ = inA5 & ~musel2;
  assign new_n543_ = ~new_n145_ & ~new_n542_;
  assign new_n544_ = ~musel3 & ~new_n543_;
  assign new_n545_ = musel1 & new_n544_;
  assign new_n546_ = inD5 & new_n274_;
  assign new_n547_ = inB5 & new_n276_;
  assign new_n548_ = ~new_n546_ & ~new_n547_;
  assign new_n549_ = ~musel1 & ~new_n548_;
  assign new_n550_ = ~new_n545_ & ~new_n549_;
  assign new_n551_ = ~musel4 & ~new_n550_;
  assign new_n552_ = inC5 & musel4;
  assign new_n553_ = ~musel3 & new_n552_;
  assign new_n554_ = ~musel2 & new_n553_;
  assign new_n555_ = ~musel1 & new_n554_;
  assign new_n556_ = musel1 & new_n145_;
  assign new_n557_ = inA5 & ~new_n252_;
  assign new_n558_ = ~new_n556_ & ~new_n557_;
  assign new_n559_ = ~musel4 & ~new_n558_;
  assign new_n560_ = musel3 & new_n559_;
  assign new_n561_ = ~new_n555_ & ~new_n560_;
  assign new_n562_ = new_n297_ & new_n561_;
  assign new_n563_ = ~new_n297_ & ~new_n561_;
  assign new_n564_ = ~new_n562_ & ~new_n563_;
  assign new_n565_ = inA4 & ~musel2;
  assign new_n566_ = ~new_n154_ & ~new_n565_;
  assign new_n567_ = ~musel3 & ~new_n566_;
  assign new_n568_ = musel1 & new_n567_;
  assign new_n569_ = inD4 & new_n274_;
  assign new_n570_ = inB4 & new_n276_;
  assign new_n571_ = ~new_n569_ & ~new_n570_;
  assign new_n572_ = ~musel1 & ~new_n571_;
  assign new_n573_ = ~new_n568_ & ~new_n572_;
  assign new_n574_ = ~musel4 & ~new_n573_;
  assign new_n575_ = inC4 & musel4;
  assign new_n576_ = ~musel3 & new_n575_;
  assign new_n577_ = ~musel2 & new_n576_;
  assign new_n578_ = ~musel1 & new_n577_;
  assign new_n579_ = musel1 & new_n154_;
  assign new_n580_ = inA4 & ~new_n252_;
  assign new_n581_ = ~new_n579_ & ~new_n580_;
  assign new_n582_ = ~musel4 & ~new_n581_;
  assign new_n583_ = musel3 & new_n582_;
  assign new_n584_ = ~new_n578_ & ~new_n583_;
  assign new_n585_ = new_n297_ & new_n584_;
  assign new_n586_ = ~new_n297_ & ~new_n584_;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = ~new_n551_ & new_n564_;
  assign new_n589_ = ~new_n574_ & new_n587_;
  assign new_n590_ = ~new_n588_ & ~new_n589_;
  assign new_n591_ = new_n541_ & new_n590_;
  assign new_n592_ = new_n574_ & ~new_n587_;
  assign new_n593_ = new_n551_ & ~new_n564_;
  assign new_n594_ = ~new_n588_ & new_n592_;
  assign new_n595_ = ~new_n593_ & ~new_n594_;
  assign new_n596_ = ~new_n540_ & ~new_n595_;
  assign new_n597_ = new_n525_ & ~new_n538_;
  assign new_n598_ = ~new_n596_ & ~new_n597_;
  assign new_n599_ = ~new_n539_ & ~new_n598_;
  assign new_n600_ = new_n502_ & ~new_n515_;
  assign new_n601_ = ~new_n599_ & ~new_n600_;
  assign new_n602_ = ~new_n492_ & new_n591_;
  assign new_n603_ = new_n601_ & ~new_n602_;
  assign new_n604_ = inA11 & ~musel2;
  assign new_n605_ = ~new_n166_ & ~new_n604_;
  assign new_n606_ = ~musel3 & ~new_n605_;
  assign new_n607_ = musel1 & new_n606_;
  assign new_n608_ = inD11 & new_n274_;
  assign new_n609_ = inB11 & new_n276_;
  assign new_n610_ = ~new_n608_ & ~new_n609_;
  assign new_n611_ = ~musel1 & ~new_n610_;
  assign new_n612_ = ~new_n607_ & ~new_n611_;
  assign new_n613_ = ~musel4 & ~new_n612_;
  assign new_n614_ = inC11 & musel4;
  assign new_n615_ = ~musel3 & new_n614_;
  assign new_n616_ = ~musel2 & new_n615_;
  assign new_n617_ = ~musel1 & new_n616_;
  assign new_n618_ = musel1 & new_n166_;
  assign new_n619_ = inA11 & ~new_n252_;
  assign new_n620_ = ~new_n618_ & ~new_n619_;
  assign new_n621_ = ~musel4 & ~new_n620_;
  assign new_n622_ = musel3 & new_n621_;
  assign new_n623_ = ~new_n617_ & ~new_n622_;
  assign new_n624_ = new_n297_ & new_n623_;
  assign new_n625_ = ~new_n297_ & ~new_n623_;
  assign new_n626_ = ~new_n624_ & ~new_n625_;
  assign new_n627_ = inA10 & ~musel2;
  assign new_n628_ = ~new_n175_ & ~new_n627_;
  assign new_n629_ = ~musel3 & ~new_n628_;
  assign new_n630_ = musel1 & new_n629_;
  assign new_n631_ = inD10 & new_n274_;
  assign new_n632_ = inB10 & new_n276_;
  assign new_n633_ = ~new_n631_ & ~new_n632_;
  assign new_n634_ = ~musel1 & ~new_n633_;
  assign new_n635_ = ~new_n630_ & ~new_n634_;
  assign new_n636_ = ~musel4 & ~new_n635_;
  assign new_n637_ = inC10 & musel4;
  assign new_n638_ = ~musel3 & new_n637_;
  assign new_n639_ = ~musel2 & new_n638_;
  assign new_n640_ = ~musel1 & new_n639_;
  assign new_n641_ = musel1 & new_n175_;
  assign new_n642_ = inA10 & ~new_n252_;
  assign new_n643_ = ~new_n641_ & ~new_n642_;
  assign new_n644_ = ~musel4 & ~new_n643_;
  assign new_n645_ = musel3 & new_n644_;
  assign new_n646_ = ~new_n640_ & ~new_n645_;
  assign new_n647_ = new_n297_ & new_n646_;
  assign new_n648_ = ~new_n297_ & ~new_n646_;
  assign new_n649_ = ~new_n647_ & ~new_n648_;
  assign new_n650_ = ~new_n613_ & new_n626_;
  assign new_n651_ = ~new_n636_ & new_n649_;
  assign new_n652_ = ~new_n650_ & ~new_n651_;
  assign new_n653_ = inA9 & ~musel2;
  assign new_n654_ = ~new_n184_ & ~new_n653_;
  assign new_n655_ = ~musel3 & ~new_n654_;
  assign new_n656_ = musel1 & new_n655_;
  assign new_n657_ = inD9 & new_n274_;
  assign new_n658_ = inB9 & new_n276_;
  assign new_n659_ = ~new_n657_ & ~new_n658_;
  assign new_n660_ = ~musel1 & ~new_n659_;
  assign new_n661_ = ~new_n656_ & ~new_n660_;
  assign new_n662_ = ~musel4 & ~new_n661_;
  assign new_n663_ = inC9 & musel4;
  assign new_n664_ = ~musel3 & new_n663_;
  assign new_n665_ = ~musel2 & new_n664_;
  assign new_n666_ = ~musel1 & new_n665_;
  assign new_n667_ = musel1 & new_n184_;
  assign new_n668_ = inA9 & ~new_n252_;
  assign new_n669_ = ~new_n667_ & ~new_n668_;
  assign new_n670_ = ~musel4 & ~new_n669_;
  assign new_n671_ = musel3 & new_n670_;
  assign new_n672_ = ~new_n666_ & ~new_n671_;
  assign new_n673_ = new_n297_ & new_n672_;
  assign new_n674_ = ~new_n297_ & ~new_n672_;
  assign new_n675_ = ~new_n673_ & ~new_n674_;
  assign new_n676_ = inA8 & ~musel2;
  assign new_n677_ = ~new_n193_ & ~new_n676_;
  assign new_n678_ = ~musel3 & ~new_n677_;
  assign new_n679_ = musel1 & new_n678_;
  assign new_n680_ = inD8 & new_n274_;
  assign new_n681_ = inB8 & new_n276_;
  assign new_n682_ = ~new_n680_ & ~new_n681_;
  assign new_n683_ = ~musel1 & ~new_n682_;
  assign new_n684_ = ~new_n679_ & ~new_n683_;
  assign new_n685_ = ~musel4 & ~new_n684_;
  assign new_n686_ = inC8 & musel4;
  assign new_n687_ = ~musel3 & new_n686_;
  assign new_n688_ = ~musel2 & new_n687_;
  assign new_n689_ = ~musel1 & new_n688_;
  assign new_n690_ = musel1 & new_n193_;
  assign new_n691_ = inA8 & ~new_n252_;
  assign new_n692_ = ~new_n690_ & ~new_n691_;
  assign new_n693_ = ~musel4 & ~new_n692_;
  assign new_n694_ = musel3 & new_n693_;
  assign new_n695_ = ~new_n689_ & ~new_n694_;
  assign new_n696_ = new_n297_ & new_n695_;
  assign new_n697_ = ~new_n297_ & ~new_n695_;
  assign new_n698_ = ~new_n696_ & ~new_n697_;
  assign new_n699_ = ~new_n662_ & new_n675_;
  assign new_n700_ = ~new_n685_ & new_n698_;
  assign new_n701_ = ~new_n699_ & ~new_n700_;
  assign new_n702_ = ~new_n603_ & new_n652_;
  assign new_n703_ = new_n701_ & new_n702_;
  assign new_n704_ = new_n685_ & ~new_n698_;
  assign new_n705_ = ~new_n699_ & new_n704_;
  assign new_n706_ = new_n662_ & ~new_n675_;
  assign new_n707_ = ~new_n705_ & ~new_n706_;
  assign new_n708_ = ~new_n651_ & ~new_n707_;
  assign new_n709_ = new_n636_ & ~new_n649_;
  assign new_n710_ = ~new_n708_ & ~new_n709_;
  assign new_n711_ = ~new_n650_ & ~new_n710_;
  assign new_n712_ = new_n613_ & ~new_n626_;
  assign new_n713_ = ~new_n711_ & ~new_n712_;
  assign new_n714_ = ~new_n703_ & new_n713_;
  assign new_n715_ = new_n364_ & ~new_n374_;
  assign new_n716_ = ~new_n375_ & new_n714_;
  assign new_n717_ = ~new_n715_ & ~new_n716_;
  assign new_n718_ = new_n340_ & ~new_n350_;
  assign new_n719_ = ~new_n351_ & ~new_n717_;
  assign new_n720_ = ~new_n718_ & ~new_n719_;
  assign new_n721_ = new_n316_ & ~new_n326_;
  assign new_n722_ = ~new_n327_ & ~new_n720_;
  assign new_n723_ = ~new_n721_ & ~new_n722_;
  assign new_n724_ = ~new_n714_ & ~new_n715_;
  assign new_n725_ = ~new_n375_ & ~new_n724_;
  assign new_n726_ = ~new_n718_ & ~new_n725_;
  assign new_n727_ = ~new_n351_ & ~new_n726_;
  assign new_n728_ = ~new_n721_ & ~new_n727_;
  assign new_n729_ = ~new_n327_ & ~new_n728_;
  assign new_n730_ = new_n303_ & ~new_n729_;
  assign new_n731_ = ~new_n303_ & ~new_n723_;
  assign new_n732_ = ~new_n730_ & ~new_n731_;
  assign new_n733_ = opsel1 & ~opsel0;
  assign new_n734_ = ~opsel1 & opsel0;
  assign new_n735_ = ~new_n733_ & ~new_n734_;
  assign new_n736_ = new_n92_ & ~new_n262_;
  assign new_n737_ = ~new_n732_ & ~new_n735_;
  assign new_n738_ = ~new_n736_ & ~new_n737_;
  assign new_n739_ = ~opsel2 & ~new_n738_;
  assign new_n740_ = opsel3 & new_n739_;
  assign new_n741_ = ~opsel3 & ~new_n269_;
  assign O15 = new_n740_ | new_n741_;
  assign new_n743_ = inD14 & musel2;
  assign new_n744_ = musel1 & new_n743_;
  assign new_n745_ = inB14 & ~new_n252_;
  assign new_n746_ = ~new_n744_ & ~new_n745_;
  assign new_n747_ = inD14 & musel4;
  assign new_n748_ = new_n258_ & new_n747_;
  assign new_n749_ = new_n256_ & ~new_n746_;
  assign new_n750_ = ~new_n748_ & ~new_n749_;
  assign new_n751_ = sh2 & ~sh0;
  assign new_n752_ = ~sh1 & sh0;
  assign new_n753_ = ~new_n751_ & ~new_n752_;
  assign new_n754_ = ~sh2 & sh1;
  assign new_n755_ = new_n753_ & ~new_n754_;
  assign new_n756_ = ~new_n262_ & ~new_n755_;
  assign new_n757_ = ~new_n750_ & new_n755_;
  assign new_n758_ = ~new_n756_ & ~new_n757_;
  assign new_n759_ = ~new_n117_ & new_n246_;
  assign new_n760_ = ~new_n126_ & new_n759_;
  assign new_n761_ = ~new_n108_ & ~new_n760_;
  assign new_n762_ = new_n108_ & new_n760_;
  assign new_n763_ = ~new_n761_ & ~new_n762_;
  assign new_n764_ = opsel2 & ~new_n758_;
  assign new_n765_ = ~opsel2 & ~new_n763_;
  assign new_n766_ = ~new_n764_ & ~new_n765_;
  assign new_n767_ = opsel2 & ~new_n763_;
  assign new_n768_ = new_n92_ & new_n767_;
  assign new_n769_ = ~new_n92_ & ~new_n766_;
  assign new_n770_ = ~new_n768_ & ~new_n769_;
  assign new_n771_ = new_n316_ & new_n326_;
  assign new_n772_ = ~new_n316_ & ~new_n326_;
  assign new_n773_ = ~new_n771_ & ~new_n772_;
  assign new_n774_ = ~new_n727_ & new_n773_;
  assign new_n775_ = ~new_n720_ & ~new_n773_;
  assign new_n776_ = ~new_n774_ & ~new_n775_;
  assign new_n777_ = new_n92_ & ~new_n758_;
  assign new_n778_ = ~new_n735_ & ~new_n776_;
  assign new_n779_ = ~new_n777_ & ~new_n778_;
  assign new_n780_ = ~opsel2 & ~new_n779_;
  assign new_n781_ = opsel3 & new_n780_;
  assign new_n782_ = ~opsel3 & ~new_n770_;
  assign O14 = new_n781_ | new_n782_;
  assign new_n784_ = sh2 & sh0;
  assign new_n785_ = inD13 & musel2;
  assign new_n786_ = musel1 & new_n785_;
  assign new_n787_ = inB13 & ~new_n252_;
  assign new_n788_ = ~new_n786_ & ~new_n787_;
  assign new_n789_ = inD13 & musel4;
  assign new_n790_ = new_n258_ & new_n789_;
  assign new_n791_ = new_n256_ & ~new_n788_;
  assign new_n792_ = ~new_n790_ & ~new_n791_;
  assign new_n793_ = sh1 & ~new_n792_;
  assign new_n794_ = sh1 & ~new_n784_;
  assign new_n795_ = sh2 & ~sh1;
  assign new_n796_ = ~new_n794_ & ~new_n795_;
  assign new_n797_ = ~sh0 & ~new_n792_;
  assign new_n798_ = sh0 & ~new_n750_;
  assign new_n799_ = ~new_n797_ & ~new_n798_;
  assign new_n800_ = ~sh2 & ~sh1;
  assign new_n801_ = ~new_n262_ & ~new_n796_;
  assign new_n802_ = ~new_n799_ & new_n800_;
  assign new_n803_ = ~new_n801_ & ~new_n802_;
  assign new_n804_ = new_n784_ & new_n793_;
  assign new_n805_ = new_n803_ & ~new_n804_;
  assign new_n806_ = ~new_n117_ & ~new_n248_;
  assign new_n807_ = new_n117_ & new_n248_;
  assign new_n808_ = ~new_n806_ & ~new_n807_;
  assign new_n809_ = opsel2 & ~new_n805_;
  assign new_n810_ = ~opsel2 & ~new_n808_;
  assign new_n811_ = ~new_n809_ & ~new_n810_;
  assign new_n812_ = opsel2 & ~new_n808_;
  assign new_n813_ = new_n92_ & new_n812_;
  assign new_n814_ = ~new_n92_ & ~new_n811_;
  assign new_n815_ = ~new_n813_ & ~new_n814_;
  assign new_n816_ = new_n340_ & new_n350_;
  assign new_n817_ = ~new_n340_ & ~new_n350_;
  assign new_n818_ = ~new_n816_ & ~new_n817_;
  assign new_n819_ = ~new_n725_ & new_n818_;
  assign new_n820_ = ~new_n717_ & ~new_n818_;
  assign new_n821_ = ~new_n819_ & ~new_n820_;
  assign new_n822_ = new_n92_ & ~new_n805_;
  assign new_n823_ = ~new_n735_ & ~new_n821_;
  assign new_n824_ = ~new_n822_ & ~new_n823_;
  assign new_n825_ = ~opsel2 & ~new_n824_;
  assign new_n826_ = opsel3 & new_n825_;
  assign new_n827_ = ~opsel3 & ~new_n815_;
  assign O13 = new_n826_ | new_n827_;
  assign new_n829_ = inD12 & musel2;
  assign new_n830_ = musel1 & new_n829_;
  assign new_n831_ = inB12 & ~new_n252_;
  assign new_n832_ = ~new_n830_ & ~new_n831_;
  assign new_n833_ = inD12 & musel4;
  assign new_n834_ = new_n258_ & new_n833_;
  assign new_n835_ = new_n256_ & ~new_n832_;
  assign new_n836_ = ~new_n834_ & ~new_n835_;
  assign new_n837_ = sh1 & sh0;
  assign new_n838_ = ~new_n836_ & new_n837_;
  assign new_n839_ = ~new_n262_ & ~new_n837_;
  assign new_n840_ = ~new_n838_ & ~new_n839_;
  assign new_n841_ = ~sh1 & ~new_n836_;
  assign new_n842_ = sh1 & ~new_n750_;
  assign new_n843_ = ~new_n841_ & ~new_n842_;
  assign new_n844_ = new_n752_ & ~new_n792_;
  assign new_n845_ = ~new_n262_ & new_n837_;
  assign new_n846_ = ~new_n844_ & ~new_n845_;
  assign new_n847_ = ~sh0 & ~new_n843_;
  assign new_n848_ = new_n846_ & ~new_n847_;
  assign new_n849_ = sh2 & ~new_n840_;
  assign new_n850_ = ~sh2 & ~new_n848_;
  assign new_n851_ = ~new_n849_ & ~new_n850_;
  assign new_n852_ = ~new_n364_ & ~new_n374_;
  assign new_n853_ = new_n364_ & new_n374_;
  assign new_n854_ = ~new_n852_ & ~new_n853_;
  assign new_n855_ = ~new_n714_ & new_n854_;
  assign new_n856_ = new_n714_ & ~new_n854_;
  assign new_n857_ = ~new_n855_ & ~new_n856_;
  assign new_n858_ = new_n92_ & ~new_n851_;
  assign new_n859_ = ~new_n735_ & ~new_n857_;
  assign new_n860_ = ~new_n858_ & ~new_n859_;
  assign new_n861_ = opsel3 & ~opsel2;
  assign new_n862_ = ~new_n126_ & ~new_n246_;
  assign new_n863_ = new_n126_ & new_n246_;
  assign new_n864_ = ~new_n862_ & ~new_n863_;
  assign new_n865_ = opsel2 & ~new_n851_;
  assign new_n866_ = ~opsel2 & ~new_n864_;
  assign new_n867_ = ~new_n865_ & ~new_n866_;
  assign new_n868_ = opsel2 & ~new_n864_;
  assign new_n869_ = new_n92_ & new_n868_;
  assign new_n870_ = ~new_n92_ & ~new_n867_;
  assign new_n871_ = ~new_n869_ & ~new_n870_;
  assign new_n872_ = ~new_n860_ & new_n861_;
  assign new_n873_ = ~opsel3 & ~new_n871_;
  assign O12 = new_n872_ | new_n873_;
  assign new_n875_ = inD11 & musel2;
  assign new_n876_ = musel1 & new_n875_;
  assign new_n877_ = inB11 & ~new_n252_;
  assign new_n878_ = ~new_n876_ & ~new_n877_;
  assign new_n879_ = inD11 & musel4;
  assign new_n880_ = new_n258_ & new_n879_;
  assign new_n881_ = new_n256_ & ~new_n878_;
  assign new_n882_ = ~new_n880_ & ~new_n881_;
  assign new_n883_ = ~sh2 & ~new_n750_;
  assign new_n884_ = sh2 & ~new_n882_;
  assign new_n885_ = ~new_n883_ & ~new_n884_;
  assign new_n886_ = sh2 & ~new_n262_;
  assign new_n887_ = ~sh1 & ~new_n882_;
  assign new_n888_ = ~new_n793_ & ~new_n887_;
  assign new_n889_ = new_n752_ & ~new_n836_;
  assign new_n890_ = ~sh0 & ~new_n888_;
  assign new_n891_ = ~new_n889_ & ~new_n890_;
  assign new_n892_ = ~new_n837_ & new_n886_;
  assign new_n893_ = ~sh2 & ~new_n891_;
  assign new_n894_ = ~new_n892_ & ~new_n893_;
  assign new_n895_ = new_n837_ & ~new_n885_;
  assign new_n896_ = new_n894_ & ~new_n895_;
  assign new_n897_ = new_n204_ & new_n243_;
  assign new_n898_ = new_n105_ & new_n897_;
  assign new_n899_ = ~new_n183_ & ~new_n192_;
  assign new_n900_ = ~new_n201_ & new_n898_;
  assign new_n901_ = new_n899_ & new_n900_;
  assign new_n902_ = ~new_n174_ & ~new_n901_;
  assign new_n903_ = new_n174_ & new_n901_;
  assign new_n904_ = ~new_n902_ & ~new_n903_;
  assign new_n905_ = opsel2 & ~new_n896_;
  assign new_n906_ = ~opsel2 & ~new_n904_;
  assign new_n907_ = ~new_n905_ & ~new_n906_;
  assign new_n908_ = opsel2 & ~new_n904_;
  assign new_n909_ = new_n92_ & new_n908_;
  assign new_n910_ = ~new_n92_ & ~new_n907_;
  assign new_n911_ = ~new_n909_ & ~new_n910_;
  assign new_n912_ = new_n613_ & new_n626_;
  assign new_n913_ = ~new_n613_ & ~new_n626_;
  assign new_n914_ = ~new_n912_ & ~new_n913_;
  assign new_n915_ = new_n603_ & ~new_n704_;
  assign new_n916_ = ~new_n700_ & ~new_n915_;
  assign new_n917_ = ~new_n706_ & ~new_n916_;
  assign new_n918_ = ~new_n699_ & ~new_n917_;
  assign new_n919_ = ~new_n709_ & ~new_n918_;
  assign new_n920_ = ~new_n651_ & ~new_n919_;
  assign new_n921_ = ~new_n603_ & ~new_n700_;
  assign new_n922_ = ~new_n704_ & ~new_n921_;
  assign new_n923_ = ~new_n699_ & ~new_n922_;
  assign new_n924_ = ~new_n706_ & ~new_n923_;
  assign new_n925_ = ~new_n651_ & ~new_n924_;
  assign new_n926_ = ~new_n709_ & ~new_n925_;
  assign new_n927_ = new_n914_ & ~new_n926_;
  assign new_n928_ = ~new_n914_ & ~new_n920_;
  assign new_n929_ = ~new_n927_ & ~new_n928_;
  assign new_n930_ = new_n92_ & ~new_n896_;
  assign new_n931_ = ~new_n735_ & ~new_n929_;
  assign new_n932_ = ~new_n930_ & ~new_n931_;
  assign new_n933_ = ~opsel2 & ~new_n932_;
  assign new_n934_ = opsel3 & new_n933_;
  assign new_n935_ = ~opsel3 & ~new_n911_;
  assign O11 = new_n934_ | new_n935_;
  assign new_n937_ = inD10 & musel2;
  assign new_n938_ = musel1 & new_n937_;
  assign new_n939_ = inB10 & ~new_n252_;
  assign new_n940_ = ~new_n938_ & ~new_n939_;
  assign new_n941_ = inD10 & musel4;
  assign new_n942_ = new_n258_ & new_n941_;
  assign new_n943_ = new_n256_ & ~new_n940_;
  assign new_n944_ = ~new_n942_ & ~new_n943_;
  assign new_n945_ = sh2 & ~new_n944_;
  assign new_n946_ = ~sh2 & ~new_n792_;
  assign new_n947_ = ~new_n945_ & ~new_n946_;
  assign new_n948_ = ~sh2 & ~new_n882_;
  assign new_n949_ = ~new_n886_ & ~new_n948_;
  assign new_n950_ = sh1 & ~new_n947_;
  assign new_n951_ = ~sh1 & ~new_n949_;
  assign new_n952_ = ~new_n950_ & ~new_n951_;
  assign new_n953_ = ~sh2 & ~new_n836_;
  assign new_n954_ = ~new_n886_ & ~new_n953_;
  assign new_n955_ = ~sh2 & ~new_n944_;
  assign new_n956_ = sh2 & ~new_n750_;
  assign new_n957_ = ~new_n955_ & ~new_n956_;
  assign new_n958_ = sh1 & ~new_n954_;
  assign new_n959_ = ~sh1 & ~new_n957_;
  assign new_n960_ = ~new_n958_ & ~new_n959_;
  assign new_n961_ = sh0 & ~new_n952_;
  assign new_n962_ = ~sh0 & ~new_n960_;
  assign new_n963_ = ~new_n961_ & ~new_n962_;
  assign new_n964_ = ~new_n192_ & new_n898_;
  assign new_n965_ = ~new_n201_ & new_n964_;
  assign new_n966_ = ~new_n183_ & ~new_n965_;
  assign new_n967_ = new_n183_ & new_n965_;
  assign new_n968_ = ~new_n966_ & ~new_n967_;
  assign new_n969_ = opsel2 & ~new_n963_;
  assign new_n970_ = ~opsel2 & ~new_n968_;
  assign new_n971_ = ~new_n969_ & ~new_n970_;
  assign new_n972_ = opsel2 & ~new_n968_;
  assign new_n973_ = new_n92_ & new_n972_;
  assign new_n974_ = ~new_n92_ & ~new_n971_;
  assign new_n975_ = ~new_n973_ & ~new_n974_;
  assign new_n976_ = new_n636_ & new_n649_;
  assign new_n977_ = ~new_n636_ & ~new_n649_;
  assign new_n978_ = ~new_n976_ & ~new_n977_;
  assign new_n979_ = ~new_n924_ & new_n978_;
  assign new_n980_ = ~new_n918_ & ~new_n978_;
  assign new_n981_ = ~new_n979_ & ~new_n980_;
  assign new_n982_ = new_n92_ & ~new_n963_;
  assign new_n983_ = ~new_n735_ & ~new_n981_;
  assign new_n984_ = ~new_n982_ & ~new_n983_;
  assign new_n985_ = ~opsel2 & ~new_n984_;
  assign new_n986_ = opsel3 & new_n985_;
  assign new_n987_ = ~opsel3 & ~new_n975_;
  assign O10 = new_n986_ | new_n987_;
  assign new_n989_ = inD9 & musel2;
  assign new_n990_ = musel1 & new_n989_;
  assign new_n991_ = inB9 & ~new_n252_;
  assign new_n992_ = ~new_n990_ & ~new_n991_;
  assign new_n993_ = inD9 & musel4;
  assign new_n994_ = new_n258_ & new_n993_;
  assign new_n995_ = new_n256_ & ~new_n992_;
  assign new_n996_ = ~new_n994_ & ~new_n995_;
  assign new_n997_ = sh2 & ~new_n996_;
  assign new_n998_ = ~new_n953_ & ~new_n997_;
  assign new_n999_ = sh1 & ~new_n998_;
  assign new_n1000_ = ~new_n959_ & ~new_n999_;
  assign new_n1001_ = ~sh2 & ~new_n996_;
  assign new_n1002_ = sh2 & ~new_n792_;
  assign new_n1003_ = ~new_n1001_ & ~new_n1002_;
  assign new_n1004_ = sh1 & ~new_n949_;
  assign new_n1005_ = ~sh1 & ~new_n1003_;
  assign new_n1006_ = ~new_n1004_ & ~new_n1005_;
  assign new_n1007_ = sh0 & ~new_n1000_;
  assign new_n1008_ = ~sh0 & ~new_n1006_;
  assign new_n1009_ = ~new_n1007_ & ~new_n1008_;
  assign new_n1010_ = ~new_n192_ & ~new_n900_;
  assign new_n1011_ = new_n192_ & new_n900_;
  assign new_n1012_ = ~new_n1010_ & ~new_n1011_;
  assign new_n1013_ = opsel2 & ~new_n1009_;
  assign new_n1014_ = ~opsel2 & ~new_n1012_;
  assign new_n1015_ = ~new_n1013_ & ~new_n1014_;
  assign new_n1016_ = opsel2 & ~new_n1012_;
  assign new_n1017_ = new_n92_ & new_n1016_;
  assign new_n1018_ = ~new_n92_ & ~new_n1015_;
  assign new_n1019_ = ~new_n1017_ & ~new_n1018_;
  assign new_n1020_ = new_n662_ & new_n675_;
  assign new_n1021_ = ~new_n662_ & ~new_n675_;
  assign new_n1022_ = ~new_n1020_ & ~new_n1021_;
  assign new_n1023_ = ~new_n922_ & new_n1022_;
  assign new_n1024_ = ~new_n916_ & ~new_n1022_;
  assign new_n1025_ = ~new_n1023_ & ~new_n1024_;
  assign new_n1026_ = new_n92_ & ~new_n1009_;
  assign new_n1027_ = ~new_n735_ & ~new_n1025_;
  assign new_n1028_ = ~new_n1026_ & ~new_n1027_;
  assign new_n1029_ = ~opsel2 & ~new_n1028_;
  assign new_n1030_ = opsel3 & new_n1029_;
  assign new_n1031_ = ~opsel3 & ~new_n1019_;
  assign O9 = new_n1030_ | new_n1031_;
  assign new_n1033_ = inD8 & musel2;
  assign new_n1034_ = musel1 & new_n1033_;
  assign new_n1035_ = inB8 & ~new_n252_;
  assign new_n1036_ = ~new_n1034_ & ~new_n1035_;
  assign new_n1037_ = inD8 & musel4;
  assign new_n1038_ = new_n258_ & new_n1037_;
  assign new_n1039_ = new_n256_ & ~new_n1036_;
  assign new_n1040_ = ~new_n1038_ & ~new_n1039_;
  assign new_n1041_ = sh2 & ~new_n1040_;
  assign new_n1042_ = ~new_n948_ & ~new_n1041_;
  assign new_n1043_ = sh1 & ~new_n1042_;
  assign new_n1044_ = ~new_n1005_ & ~new_n1043_;
  assign new_n1045_ = ~new_n886_ & ~new_n955_;
  assign new_n1046_ = ~sh2 & ~new_n1040_;
  assign new_n1047_ = sh2 & ~new_n836_;
  assign new_n1048_ = ~new_n1046_ & ~new_n1047_;
  assign new_n1049_ = sh1 & ~new_n1045_;
  assign new_n1050_ = ~sh1 & ~new_n1048_;
  assign new_n1051_ = ~new_n1049_ & ~new_n1050_;
  assign new_n1052_ = sh0 & ~new_n1044_;
  assign new_n1053_ = ~sh0 & ~new_n1051_;
  assign new_n1054_ = ~new_n1052_ & ~new_n1053_;
  assign new_n1055_ = new_n685_ & new_n698_;
  assign new_n1056_ = ~new_n685_ & ~new_n698_;
  assign new_n1057_ = ~new_n1055_ & ~new_n1056_;
  assign new_n1058_ = ~new_n603_ & new_n1057_;
  assign new_n1059_ = new_n603_ & ~new_n1057_;
  assign new_n1060_ = ~new_n1058_ & ~new_n1059_;
  assign new_n1061_ = new_n92_ & ~new_n1054_;
  assign new_n1062_ = ~new_n735_ & ~new_n1060_;
  assign new_n1063_ = ~new_n1061_ & ~new_n1062_;
  assign new_n1064_ = ~new_n201_ & ~new_n898_;
  assign new_n1065_ = new_n201_ & new_n898_;
  assign new_n1066_ = ~new_n1064_ & ~new_n1065_;
  assign new_n1067_ = opsel2 & ~new_n1054_;
  assign new_n1068_ = ~opsel2 & ~new_n1066_;
  assign new_n1069_ = ~new_n1067_ & ~new_n1068_;
  assign new_n1070_ = opsel2 & ~new_n1066_;
  assign new_n1071_ = new_n92_ & new_n1070_;
  assign new_n1072_ = ~new_n92_ & ~new_n1069_;
  assign new_n1073_ = ~new_n1071_ & ~new_n1072_;
  assign new_n1074_ = new_n861_ & ~new_n1063_;
  assign new_n1075_ = ~opsel3 & ~new_n1073_;
  assign O8 = new_n1074_ | new_n1075_;
  assign new_n1077_ = inD7 & musel2;
  assign new_n1078_ = musel1 & new_n1077_;
  assign new_n1079_ = inB7 & ~new_n252_;
  assign new_n1080_ = ~new_n1078_ & ~new_n1079_;
  assign new_n1081_ = inD7 & musel4;
  assign new_n1082_ = new_n258_ & new_n1081_;
  assign new_n1083_ = new_n256_ & ~new_n1080_;
  assign new_n1084_ = ~new_n1082_ & ~new_n1083_;
  assign new_n1085_ = sh2 & ~new_n1084_;
  assign new_n1086_ = ~new_n955_ & ~new_n1085_;
  assign new_n1087_ = sh1 & ~new_n1086_;
  assign new_n1088_ = ~new_n1050_ & ~new_n1087_;
  assign new_n1089_ = ~new_n886_ & ~new_n1001_;
  assign new_n1090_ = ~sh2 & ~new_n1084_;
  assign new_n1091_ = ~new_n884_ & ~new_n1090_;
  assign new_n1092_ = sh1 & ~new_n1089_;
  assign new_n1093_ = ~sh1 & ~new_n1091_;
  assign new_n1094_ = ~new_n1092_ & ~new_n1093_;
  assign new_n1095_ = sh0 & ~new_n1088_;
  assign new_n1096_ = ~sh0 & ~new_n1094_;
  assign new_n1097_ = ~new_n1095_ & ~new_n1096_;
  assign new_n1098_ = new_n105_ & new_n243_;
  assign new_n1099_ = ~new_n144_ & ~new_n153_;
  assign new_n1100_ = ~new_n162_ & new_n1098_;
  assign new_n1101_ = new_n1099_ & new_n1100_;
  assign new_n1102_ = ~new_n135_ & ~new_n1101_;
  assign new_n1103_ = new_n135_ & new_n1101_;
  assign new_n1104_ = ~new_n1102_ & ~new_n1103_;
  assign new_n1105_ = opsel2 & ~new_n1097_;
  assign new_n1106_ = ~opsel2 & ~new_n1104_;
  assign new_n1107_ = ~new_n1105_ & ~new_n1106_;
  assign new_n1108_ = opsel2 & ~new_n1104_;
  assign new_n1109_ = new_n92_ & new_n1108_;
  assign new_n1110_ = ~new_n92_ & ~new_n1107_;
  assign new_n1111_ = ~new_n1109_ & ~new_n1110_;
  assign new_n1112_ = new_n502_ & new_n515_;
  assign new_n1113_ = ~new_n502_ & ~new_n515_;
  assign new_n1114_ = ~new_n1112_ & ~new_n1113_;
  assign new_n1115_ = new_n492_ & ~new_n592_;
  assign new_n1116_ = ~new_n589_ & ~new_n1115_;
  assign new_n1117_ = ~new_n593_ & ~new_n1116_;
  assign new_n1118_ = ~new_n588_ & ~new_n1117_;
  assign new_n1119_ = ~new_n597_ & ~new_n1118_;
  assign new_n1120_ = ~new_n540_ & ~new_n1119_;
  assign new_n1121_ = ~new_n492_ & ~new_n589_;
  assign new_n1122_ = ~new_n592_ & ~new_n1121_;
  assign new_n1123_ = ~new_n588_ & ~new_n1122_;
  assign new_n1124_ = ~new_n593_ & ~new_n1123_;
  assign new_n1125_ = ~new_n540_ & ~new_n1124_;
  assign new_n1126_ = ~new_n597_ & ~new_n1125_;
  assign new_n1127_ = new_n1114_ & ~new_n1126_;
  assign new_n1128_ = ~new_n1114_ & ~new_n1120_;
  assign new_n1129_ = ~new_n1127_ & ~new_n1128_;
  assign new_n1130_ = new_n92_ & ~new_n1097_;
  assign new_n1131_ = ~new_n735_ & ~new_n1129_;
  assign new_n1132_ = ~new_n1130_ & ~new_n1131_;
  assign new_n1133_ = ~opsel2 & ~new_n1132_;
  assign new_n1134_ = opsel3 & new_n1133_;
  assign new_n1135_ = ~opsel3 & ~new_n1111_;
  assign O7 = new_n1134_ | new_n1135_;
  assign new_n1137_ = inD6 & musel2;
  assign new_n1138_ = musel1 & new_n1137_;
  assign new_n1139_ = inB6 & ~new_n252_;
  assign new_n1140_ = ~new_n1138_ & ~new_n1139_;
  assign new_n1141_ = inD6 & musel4;
  assign new_n1142_ = new_n258_ & new_n1141_;
  assign new_n1143_ = new_n256_ & ~new_n1140_;
  assign new_n1144_ = ~new_n1142_ & ~new_n1143_;
  assign new_n1145_ = sh2 & ~new_n1144_;
  assign new_n1146_ = ~new_n1001_ & ~new_n1145_;
  assign new_n1147_ = sh1 & ~new_n1146_;
  assign new_n1148_ = ~new_n1093_ & ~new_n1147_;
  assign new_n1149_ = ~new_n956_ & ~new_n1046_;
  assign new_n1150_ = ~sh2 & ~new_n1144_;
  assign new_n1151_ = ~new_n945_ & ~new_n1150_;
  assign new_n1152_ = sh1 & ~new_n1149_;
  assign new_n1153_ = ~sh1 & ~new_n1151_;
  assign new_n1154_ = ~new_n1152_ & ~new_n1153_;
  assign new_n1155_ = sh0 & ~new_n1148_;
  assign new_n1156_ = ~sh0 & ~new_n1154_;
  assign new_n1157_ = ~new_n1155_ & ~new_n1156_;
  assign new_n1158_ = ~new_n153_ & new_n1098_;
  assign new_n1159_ = ~new_n162_ & new_n1158_;
  assign new_n1160_ = ~new_n144_ & ~new_n1159_;
  assign new_n1161_ = new_n144_ & new_n1159_;
  assign new_n1162_ = ~new_n1160_ & ~new_n1161_;
  assign new_n1163_ = opsel2 & ~new_n1157_;
  assign new_n1164_ = ~opsel2 & ~new_n1162_;
  assign new_n1165_ = ~new_n1163_ & ~new_n1164_;
  assign new_n1166_ = opsel2 & ~new_n1162_;
  assign new_n1167_ = new_n92_ & new_n1166_;
  assign new_n1168_ = ~new_n92_ & ~new_n1165_;
  assign new_n1169_ = ~new_n1167_ & ~new_n1168_;
  assign new_n1170_ = new_n525_ & new_n538_;
  assign new_n1171_ = ~new_n525_ & ~new_n538_;
  assign new_n1172_ = ~new_n1170_ & ~new_n1171_;
  assign new_n1173_ = ~new_n1124_ & new_n1172_;
  assign new_n1174_ = ~new_n1118_ & ~new_n1172_;
  assign new_n1175_ = ~new_n1173_ & ~new_n1174_;
  assign new_n1176_ = new_n92_ & ~new_n1157_;
  assign new_n1177_ = ~new_n735_ & ~new_n1175_;
  assign new_n1178_ = ~new_n1176_ & ~new_n1177_;
  assign new_n1179_ = ~opsel2 & ~new_n1178_;
  assign new_n1180_ = opsel3 & new_n1179_;
  assign new_n1181_ = ~opsel3 & ~new_n1169_;
  assign O6 = new_n1180_ | new_n1181_;
  assign new_n1183_ = inD5 & musel2;
  assign new_n1184_ = musel1 & new_n1183_;
  assign new_n1185_ = inB5 & ~new_n252_;
  assign new_n1186_ = ~new_n1184_ & ~new_n1185_;
  assign new_n1187_ = inD5 & musel4;
  assign new_n1188_ = new_n258_ & new_n1187_;
  assign new_n1189_ = new_n256_ & ~new_n1186_;
  assign new_n1190_ = ~new_n1188_ & ~new_n1189_;
  assign new_n1191_ = sh2 & ~new_n1190_;
  assign new_n1192_ = ~new_n1046_ & ~new_n1191_;
  assign new_n1193_ = sh1 & ~new_n1192_;
  assign new_n1194_ = ~new_n1153_ & ~new_n1193_;
  assign new_n1195_ = ~new_n1002_ & ~new_n1090_;
  assign new_n1196_ = ~sh2 & ~new_n1190_;
  assign new_n1197_ = ~new_n997_ & ~new_n1196_;
  assign new_n1198_ = sh1 & ~new_n1195_;
  assign new_n1199_ = ~sh1 & ~new_n1197_;
  assign new_n1200_ = ~new_n1198_ & ~new_n1199_;
  assign new_n1201_ = sh0 & ~new_n1194_;
  assign new_n1202_ = ~sh0 & ~new_n1200_;
  assign new_n1203_ = ~new_n1201_ & ~new_n1202_;
  assign new_n1204_ = ~new_n153_ & ~new_n1100_;
  assign new_n1205_ = new_n153_ & new_n1100_;
  assign new_n1206_ = ~new_n1204_ & ~new_n1205_;
  assign new_n1207_ = opsel2 & ~new_n1203_;
  assign new_n1208_ = ~opsel2 & ~new_n1206_;
  assign new_n1209_ = ~new_n1207_ & ~new_n1208_;
  assign new_n1210_ = opsel2 & ~new_n1206_;
  assign new_n1211_ = new_n92_ & new_n1210_;
  assign new_n1212_ = ~new_n92_ & ~new_n1209_;
  assign new_n1213_ = ~new_n1211_ & ~new_n1212_;
  assign new_n1214_ = new_n551_ & new_n564_;
  assign new_n1215_ = ~new_n551_ & ~new_n564_;
  assign new_n1216_ = ~new_n1214_ & ~new_n1215_;
  assign new_n1217_ = ~new_n1122_ & new_n1216_;
  assign new_n1218_ = ~new_n1116_ & ~new_n1216_;
  assign new_n1219_ = ~new_n1217_ & ~new_n1218_;
  assign new_n1220_ = new_n92_ & ~new_n1203_;
  assign new_n1221_ = ~new_n735_ & ~new_n1219_;
  assign new_n1222_ = ~new_n1220_ & ~new_n1221_;
  assign new_n1223_ = ~opsel2 & ~new_n1222_;
  assign new_n1224_ = opsel3 & new_n1223_;
  assign new_n1225_ = ~opsel3 & ~new_n1213_;
  assign O5 = new_n1224_ | new_n1225_;
  assign new_n1227_ = inD4 & musel2;
  assign new_n1228_ = musel1 & new_n1227_;
  assign new_n1229_ = inB4 & ~new_n252_;
  assign new_n1230_ = ~new_n1228_ & ~new_n1229_;
  assign new_n1231_ = inD4 & musel4;
  assign new_n1232_ = new_n258_ & new_n1231_;
  assign new_n1233_ = new_n256_ & ~new_n1230_;
  assign new_n1234_ = ~new_n1232_ & ~new_n1233_;
  assign new_n1235_ = sh2 & ~new_n1234_;
  assign new_n1236_ = ~new_n1090_ & ~new_n1235_;
  assign new_n1237_ = sh1 & ~new_n1236_;
  assign new_n1238_ = ~new_n1199_ & ~new_n1237_;
  assign new_n1239_ = ~new_n1047_ & ~new_n1150_;
  assign new_n1240_ = ~sh2 & ~new_n1234_;
  assign new_n1241_ = ~new_n1041_ & ~new_n1240_;
  assign new_n1242_ = sh1 & ~new_n1239_;
  assign new_n1243_ = ~sh1 & ~new_n1241_;
  assign new_n1244_ = ~new_n1242_ & ~new_n1243_;
  assign new_n1245_ = sh0 & ~new_n1238_;
  assign new_n1246_ = ~sh0 & ~new_n1244_;
  assign new_n1247_ = ~new_n1245_ & ~new_n1246_;
  assign new_n1248_ = ~new_n574_ & ~new_n587_;
  assign new_n1249_ = new_n574_ & new_n587_;
  assign new_n1250_ = ~new_n1248_ & ~new_n1249_;
  assign new_n1251_ = ~new_n492_ & new_n1250_;
  assign new_n1252_ = new_n492_ & ~new_n1250_;
  assign new_n1253_ = ~new_n1251_ & ~new_n1252_;
  assign new_n1254_ = new_n92_ & ~new_n1247_;
  assign new_n1255_ = ~new_n735_ & ~new_n1253_;
  assign new_n1256_ = ~new_n1254_ & ~new_n1255_;
  assign new_n1257_ = ~new_n162_ & ~new_n1098_;
  assign new_n1258_ = new_n162_ & new_n1098_;
  assign new_n1259_ = ~new_n1257_ & ~new_n1258_;
  assign new_n1260_ = opsel2 & ~new_n1247_;
  assign new_n1261_ = ~opsel2 & ~new_n1259_;
  assign new_n1262_ = ~new_n1260_ & ~new_n1261_;
  assign new_n1263_ = opsel2 & ~new_n1259_;
  assign new_n1264_ = new_n92_ & new_n1263_;
  assign new_n1265_ = ~new_n92_ & ~new_n1262_;
  assign new_n1266_ = ~new_n1264_ & ~new_n1265_;
  assign new_n1267_ = new_n861_ & ~new_n1256_;
  assign new_n1268_ = ~opsel3 & ~new_n1266_;
  assign O4 = new_n1267_ | new_n1268_;
  assign new_n1270_ = inD3 & musel2;
  assign new_n1271_ = musel1 & new_n1270_;
  assign new_n1272_ = inB3 & ~new_n252_;
  assign new_n1273_ = ~new_n1271_ & ~new_n1272_;
  assign new_n1274_ = inD3 & musel4;
  assign new_n1275_ = new_n258_ & new_n1274_;
  assign new_n1276_ = new_n256_ & ~new_n1273_;
  assign new_n1277_ = ~new_n1275_ & ~new_n1276_;
  assign new_n1278_ = sh2 & ~new_n1277_;
  assign new_n1279_ = ~new_n1150_ & ~new_n1278_;
  assign new_n1280_ = sh1 & ~new_n1279_;
  assign new_n1281_ = ~new_n1243_ & ~new_n1280_;
  assign new_n1282_ = ~new_n884_ & ~new_n1196_;
  assign new_n1283_ = ~sh2 & ~new_n1277_;
  assign new_n1284_ = ~new_n1085_ & ~new_n1283_;
  assign new_n1285_ = sh1 & ~new_n1282_;
  assign new_n1286_ = ~sh1 & ~new_n1284_;
  assign new_n1287_ = ~new_n1285_ & ~new_n1286_;
  assign new_n1288_ = sh0 & ~new_n1281_;
  assign new_n1289_ = ~sh0 & ~new_n1287_;
  assign new_n1290_ = ~new_n1288_ & ~new_n1289_;
  assign new_n1291_ = ~new_n222_ & ~new_n231_;
  assign new_n1292_ = new_n105_ & ~new_n240_;
  assign new_n1293_ = new_n1291_ & new_n1292_;
  assign new_n1294_ = ~new_n213_ & ~new_n1293_;
  assign new_n1295_ = new_n213_ & new_n1293_;
  assign new_n1296_ = ~new_n1294_ & ~new_n1295_;
  assign new_n1297_ = opsel2 & ~new_n1290_;
  assign new_n1298_ = ~opsel2 & ~new_n1296_;
  assign new_n1299_ = ~new_n1297_ & ~new_n1298_;
  assign new_n1300_ = opsel2 & ~new_n1296_;
  assign new_n1301_ = new_n92_ & new_n1300_;
  assign new_n1302_ = ~new_n92_ & ~new_n1299_;
  assign new_n1303_ = ~new_n1301_ & ~new_n1302_;
  assign new_n1304_ = new_n391_ & new_n404_;
  assign new_n1305_ = ~new_n391_ & ~new_n404_;
  assign new_n1306_ = ~new_n1304_ & ~new_n1305_;
  assign new_n1307_ = ~new_n381_ & ~new_n482_;
  assign new_n1308_ = ~new_n478_ & ~new_n1307_;
  assign new_n1309_ = ~new_n483_ & ~new_n1308_;
  assign new_n1310_ = ~new_n477_ & ~new_n1309_;
  assign new_n1311_ = ~new_n487_ & ~new_n1310_;
  assign new_n1312_ = ~new_n429_ & ~new_n1311_;
  assign new_n1313_ = new_n381_ & ~new_n478_;
  assign new_n1314_ = ~new_n482_ & ~new_n1313_;
  assign new_n1315_ = ~new_n477_ & ~new_n1314_;
  assign new_n1316_ = ~new_n483_ & ~new_n1315_;
  assign new_n1317_ = ~new_n429_ & ~new_n1316_;
  assign new_n1318_ = ~new_n487_ & ~new_n1317_;
  assign new_n1319_ = new_n1306_ & ~new_n1318_;
  assign new_n1320_ = ~new_n1306_ & ~new_n1312_;
  assign new_n1321_ = ~new_n1319_ & ~new_n1320_;
  assign new_n1322_ = new_n92_ & ~new_n1290_;
  assign new_n1323_ = ~new_n735_ & ~new_n1321_;
  assign new_n1324_ = ~new_n1322_ & ~new_n1323_;
  assign new_n1325_ = ~opsel2 & ~new_n1324_;
  assign new_n1326_ = opsel3 & new_n1325_;
  assign new_n1327_ = ~opsel3 & ~new_n1303_;
  assign O3 = new_n1326_ | new_n1327_;
  assign new_n1329_ = inD2 & musel2;
  assign new_n1330_ = musel1 & new_n1329_;
  assign new_n1331_ = inB2 & ~new_n252_;
  assign new_n1332_ = ~new_n1330_ & ~new_n1331_;
  assign new_n1333_ = inD2 & musel4;
  assign new_n1334_ = new_n258_ & new_n1333_;
  assign new_n1335_ = new_n256_ & ~new_n1332_;
  assign new_n1336_ = ~new_n1334_ & ~new_n1335_;
  assign new_n1337_ = sh2 & ~new_n1336_;
  assign new_n1338_ = ~new_n1196_ & ~new_n1337_;
  assign new_n1339_ = sh1 & ~new_n1338_;
  assign new_n1340_ = ~new_n1286_ & ~new_n1339_;
  assign new_n1341_ = ~new_n945_ & ~new_n1240_;
  assign new_n1342_ = ~sh2 & ~new_n1336_;
  assign new_n1343_ = ~new_n1145_ & ~new_n1342_;
  assign new_n1344_ = sh1 & ~new_n1341_;
  assign new_n1345_ = ~sh1 & ~new_n1343_;
  assign new_n1346_ = ~new_n1344_ & ~new_n1345_;
  assign new_n1347_ = sh0 & ~new_n1340_;
  assign new_n1348_ = ~sh0 & ~new_n1346_;
  assign new_n1349_ = ~new_n1347_ & ~new_n1348_;
  assign new_n1350_ = new_n105_ & ~new_n231_;
  assign new_n1351_ = ~new_n240_ & new_n1350_;
  assign new_n1352_ = ~new_n222_ & ~new_n1351_;
  assign new_n1353_ = new_n222_ & new_n1351_;
  assign new_n1354_ = ~new_n1352_ & ~new_n1353_;
  assign new_n1355_ = opsel2 & ~new_n1349_;
  assign new_n1356_ = ~opsel2 & ~new_n1354_;
  assign new_n1357_ = ~new_n1355_ & ~new_n1356_;
  assign new_n1358_ = opsel2 & ~new_n1354_;
  assign new_n1359_ = new_n92_ & new_n1358_;
  assign new_n1360_ = ~new_n92_ & ~new_n1357_;
  assign new_n1361_ = ~new_n1359_ & ~new_n1360_;
  assign new_n1362_ = new_n414_ & new_n427_;
  assign new_n1363_ = ~new_n414_ & ~new_n427_;
  assign new_n1364_ = ~new_n1362_ & ~new_n1363_;
  assign new_n1365_ = ~new_n1316_ & new_n1364_;
  assign new_n1366_ = ~new_n1310_ & ~new_n1364_;
  assign new_n1367_ = ~new_n1365_ & ~new_n1366_;
  assign new_n1368_ = new_n92_ & ~new_n1349_;
  assign new_n1369_ = ~new_n735_ & ~new_n1367_;
  assign new_n1370_ = ~new_n1368_ & ~new_n1369_;
  assign new_n1371_ = ~opsel2 & ~new_n1370_;
  assign new_n1372_ = opsel3 & new_n1371_;
  assign new_n1373_ = ~opsel3 & ~new_n1361_;
  assign O2 = new_n1372_ | new_n1373_;
  assign new_n1375_ = inD1 & musel2;
  assign new_n1376_ = musel1 & new_n1375_;
  assign new_n1377_ = inB1 & ~new_n252_;
  assign new_n1378_ = ~new_n1376_ & ~new_n1377_;
  assign new_n1379_ = inD1 & musel4;
  assign new_n1380_ = new_n258_ & new_n1379_;
  assign new_n1381_ = new_n256_ & ~new_n1378_;
  assign new_n1382_ = ~new_n1380_ & ~new_n1381_;
  assign new_n1383_ = sh2 & ~new_n1382_;
  assign new_n1384_ = ~new_n1240_ & ~new_n1383_;
  assign new_n1385_ = sh1 & ~new_n1384_;
  assign new_n1386_ = ~new_n1345_ & ~new_n1385_;
  assign new_n1387_ = ~new_n997_ & ~new_n1283_;
  assign new_n1388_ = ~sh2 & ~new_n1382_;
  assign new_n1389_ = ~new_n1191_ & ~new_n1388_;
  assign new_n1390_ = sh1 & ~new_n1387_;
  assign new_n1391_ = ~sh1 & ~new_n1389_;
  assign new_n1392_ = ~new_n1390_ & ~new_n1391_;
  assign new_n1393_ = sh0 & ~new_n1386_;
  assign new_n1394_ = ~sh0 & ~new_n1392_;
  assign new_n1395_ = ~new_n1393_ & ~new_n1394_;
  assign new_n1396_ = ~new_n231_ & ~new_n1292_;
  assign new_n1397_ = new_n231_ & new_n1292_;
  assign new_n1398_ = ~new_n1396_ & ~new_n1397_;
  assign new_n1399_ = opsel2 & ~new_n1395_;
  assign new_n1400_ = ~opsel2 & ~new_n1398_;
  assign new_n1401_ = ~new_n1399_ & ~new_n1400_;
  assign new_n1402_ = opsel2 & ~new_n1398_;
  assign new_n1403_ = new_n92_ & new_n1402_;
  assign new_n1404_ = ~new_n92_ & ~new_n1401_;
  assign new_n1405_ = ~new_n1403_ & ~new_n1404_;
  assign new_n1406_ = new_n440_ & new_n453_;
  assign new_n1407_ = ~new_n440_ & ~new_n453_;
  assign new_n1408_ = ~new_n1406_ & ~new_n1407_;
  assign new_n1409_ = ~new_n1314_ & new_n1408_;
  assign new_n1410_ = ~new_n1308_ & ~new_n1408_;
  assign new_n1411_ = ~new_n1409_ & ~new_n1410_;
  assign new_n1412_ = new_n92_ & ~new_n1395_;
  assign new_n1413_ = ~new_n735_ & ~new_n1411_;
  assign new_n1414_ = ~new_n1412_ & ~new_n1413_;
  assign new_n1415_ = ~opsel2 & ~new_n1414_;
  assign new_n1416_ = opsel3 & new_n1415_;
  assign new_n1417_ = ~opsel3 & ~new_n1405_;
  assign O1 = new_n1416_ | new_n1417_;
  assign new_n1419_ = inD0 & musel2;
  assign new_n1420_ = musel1 & new_n1419_;
  assign new_n1421_ = inB0 & ~new_n252_;
  assign new_n1422_ = ~new_n1420_ & ~new_n1421_;
  assign new_n1423_ = inD0 & musel4;
  assign new_n1424_ = new_n258_ & new_n1423_;
  assign new_n1425_ = new_n256_ & ~new_n1422_;
  assign new_n1426_ = ~new_n1424_ & ~new_n1425_;
  assign new_n1427_ = sh2 & ~new_n1426_;
  assign new_n1428_ = ~new_n1283_ & ~new_n1427_;
  assign new_n1429_ = sh1 & ~new_n1428_;
  assign new_n1430_ = ~new_n1391_ & ~new_n1429_;
  assign new_n1431_ = ~new_n1041_ & ~new_n1342_;
  assign new_n1432_ = ~sh2 & ~new_n1426_;
  assign new_n1433_ = ~new_n1235_ & ~new_n1432_;
  assign new_n1434_ = sh1 & ~new_n1431_;
  assign new_n1435_ = ~sh1 & ~new_n1433_;
  assign new_n1436_ = ~new_n1434_ & ~new_n1435_;
  assign new_n1437_ = sh0 & ~new_n1430_;
  assign new_n1438_ = ~sh0 & ~new_n1436_;
  assign new_n1439_ = ~new_n1437_ & ~new_n1438_;
  assign new_n1440_ = ~new_n105_ & ~new_n240_;
  assign new_n1441_ = new_n105_ & new_n240_;
  assign new_n1442_ = ~new_n1440_ & ~new_n1441_;
  assign new_n1443_ = opsel2 & ~new_n1439_;
  assign new_n1444_ = ~opsel2 & ~new_n1442_;
  assign new_n1445_ = ~new_n1443_ & ~new_n1444_;
  assign new_n1446_ = opsel2 & ~new_n1442_;
  assign new_n1447_ = new_n92_ & new_n1446_;
  assign new_n1448_ = ~new_n92_ & ~new_n1445_;
  assign new_n1449_ = ~new_n1447_ & ~new_n1448_;
  assign new_n1450_ = ~new_n463_ & ~new_n476_;
  assign new_n1451_ = new_n463_ & new_n476_;
  assign new_n1452_ = ~new_n1450_ & ~new_n1451_;
  assign new_n1453_ = new_n381_ & new_n1452_;
  assign new_n1454_ = ~new_n381_ & ~new_n1452_;
  assign new_n1455_ = ~new_n1453_ & ~new_n1454_;
  assign new_n1456_ = new_n92_ & ~new_n1439_;
  assign new_n1457_ = ~new_n735_ & ~new_n1455_;
  assign new_n1458_ = ~new_n1456_ & ~new_n1457_;
  assign new_n1459_ = ~opsel2 & ~new_n1458_;
  assign new_n1460_ = opsel3 & new_n1459_;
  assign new_n1461_ = ~opsel3 & ~new_n1449_;
  assign O0 = new_n1460_ | new_n1461_;
endmodule


