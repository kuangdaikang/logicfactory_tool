// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:41 2022

module signet  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
    v30, v31, v32, v33, v34, v35, v36, v37, v38,
    \v39.0 , \v39.1 , \v39.2 , \v39.3 , \v39.4 , \v39.5 , \v39.6 , \v39.7   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28,
    v29, v30, v31, v32, v33, v34, v35, v36, v37, v38;
  output \v39.0 , \v39.1 , \v39.2 , \v39.3 , \v39.4 , \v39.5 , \v39.6 ,
    \v39.7 ;
  wire new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_,
    new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n335_,
    new_n336_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_;
  assign new_n48_ = v1 & v7;
  assign new_n49_ = ~v7 & v8;
  assign new_n50_ = ~new_n48_ & ~new_n49_;
  assign new_n51_ = v0 & ~new_n50_;
  assign new_n52_ = v1 & v9;
  assign new_n53_ = v8 & v11;
  assign new_n54_ = ~v22 & ~new_n53_;
  assign new_n55_ = ~new_n52_ & new_n54_;
  assign new_n56_ = ~new_n51_ & new_n55_;
  assign new_n57_ = ~v6 & ~new_n56_;
  assign new_n58_ = v10 & ~v14;
  assign new_n59_ = ~v17 & v18;
  assign new_n60_ = new_n58_ & new_n59_;
  assign new_n61_ = v15 & ~v24;
  assign new_n62_ = ~new_n60_ & ~new_n61_;
  assign new_n63_ = ~v1 & ~new_n62_;
  assign new_n64_ = v16 & v18;
  assign new_n65_ = ~v14 & new_n64_;
  assign new_n66_ = ~v27 & ~new_n65_;
  assign new_n67_ = ~new_n63_ & new_n66_;
  assign new_n68_ = ~new_n57_ & new_n67_;
  assign new_n69_ = ~v3 & ~new_n68_;
  assign new_n70_ = ~v2 & v3;
  assign new_n71_ = ~v1 & new_n70_;
  assign new_n72_ = v5 & v6;
  assign new_n73_ = v4 & new_n72_;
  assign new_n74_ = ~new_n71_ & ~new_n73_;
  assign new_n75_ = v0 & ~new_n74_;
  assign new_n76_ = ~v18 & ~v22;
  assign new_n77_ = v6 & ~v10;
  assign new_n78_ = ~new_n71_ & ~new_n77_;
  assign new_n79_ = ~new_n76_ & ~new_n78_;
  assign new_n80_ = v9 & v10;
  assign new_n81_ = ~v26 & ~new_n80_;
  assign new_n82_ = ~v8 & ~new_n81_;
  assign new_n83_ = v4 & v11;
  assign new_n84_ = v12 & v13;
  assign new_n85_ = new_n83_ & new_n84_;
  assign new_n86_ = ~new_n82_ & ~new_n85_;
  assign new_n87_ = ~v1 & ~new_n86_;
  assign new_n88_ = v4 & ~new_n84_;
  assign new_n89_ = ~v4 & ~v25;
  assign new_n90_ = ~new_n88_ & ~new_n89_;
  assign new_n91_ = v11 & ~new_n90_;
  assign new_n92_ = ~v15 & ~v26;
  assign new_n93_ = v10 & v12;
  assign new_n94_ = ~new_n92_ & ~new_n93_;
  assign new_n95_ = ~v17 & ~v20;
  assign new_n96_ = ~v21 & ~new_n95_;
  assign new_n97_ = v18 & ~new_n96_;
  assign new_n98_ = v9 & ~v10;
  assign new_n99_ = ~new_n97_ & ~new_n98_;
  assign new_n100_ = ~new_n94_ & new_n99_;
  assign new_n101_ = ~new_n91_ & new_n100_;
  assign new_n102_ = ~new_n87_ & new_n101_;
  assign new_n103_ = v6 & ~new_n102_;
  assign new_n104_ = v1 & ~v17;
  assign new_n105_ = ~v17 & ~new_n104_;
  assign new_n106_ = ~v16 & ~new_n105_;
  assign new_n107_ = ~v16 & ~new_n106_;
  assign new_n108_ = ~new_n92_ & ~new_n107_;
  assign new_n109_ = ~v16 & new_n59_;
  assign new_n110_ = ~v11 & ~new_n109_;
  assign new_n111_ = v1 & ~new_n110_;
  assign new_n112_ = ~v16 & v17;
  assign new_n113_ = ~v19 & ~new_n112_;
  assign new_n114_ = v18 & ~new_n113_;
  assign new_n115_ = ~v23 & v26;
  assign new_n116_ = v19 & new_n115_;
  assign new_n117_ = ~new_n114_ & ~new_n116_;
  assign new_n118_ = ~new_n111_ & new_n117_;
  assign new_n119_ = ~new_n108_ & new_n118_;
  assign new_n120_ = v24 & ~new_n119_;
  assign new_n121_ = ~v1 & ~v8;
  assign new_n122_ = ~v23 & ~new_n121_;
  assign new_n123_ = v11 & ~new_n122_;
  assign new_n124_ = v18 & v19;
  assign new_n125_ = ~new_n115_ & ~new_n124_;
  assign new_n126_ = ~v1 & ~new_n125_;
  assign new_n127_ = ~v17 & v20;
  assign new_n128_ = v1 & new_n127_;
  assign new_n129_ = ~v17 & ~new_n128_;
  assign new_n130_ = v18 & ~new_n129_;
  assign new_n131_ = ~new_n126_ & ~new_n130_;
  assign new_n132_ = ~new_n123_ & new_n131_;
  assign new_n133_ = v14 & ~new_n132_;
  assign new_n134_ = ~v14 & v22;
  assign new_n135_ = v23 & ~v24;
  assign new_n136_ = new_n134_ & new_n135_;
  assign new_n137_ = ~new_n133_ & ~new_n136_;
  assign new_n138_ = ~new_n120_ & new_n137_;
  assign new_n139_ = ~new_n103_ & new_n138_;
  assign new_n140_ = ~new_n79_ & new_n139_;
  assign new_n141_ = ~new_n75_ & new_n140_;
  assign \v39.0  = new_n69_ | ~new_n141_;
  assign new_n143_ = v2 & v3;
  assign new_n144_ = ~v1 & ~v3;
  assign new_n145_ = ~v6 & v7;
  assign new_n146_ = new_n144_ & new_n145_;
  assign new_n147_ = ~new_n143_ & ~new_n146_;
  assign new_n148_ = v0 & ~new_n147_;
  assign new_n149_ = v12 & v26;
  assign new_n150_ = ~v9 & ~new_n149_;
  assign new_n151_ = ~new_n121_ & ~new_n150_;
  assign new_n152_ = v12 & v15;
  assign new_n153_ = v1 & new_n152_;
  assign new_n154_ = v22 & v23;
  assign new_n155_ = ~new_n153_ & ~new_n154_;
  assign new_n156_ = ~new_n151_ & new_n155_;
  assign new_n157_ = v6 & ~new_n156_;
  assign new_n158_ = ~v3 & v18;
  assign new_n159_ = v24 & v26;
  assign new_n160_ = ~new_n158_ & ~new_n159_;
  assign new_n161_ = v17 & v33;
  assign new_n162_ = ~v20 & ~v34;
  assign new_n163_ = new_n104_ & new_n162_;
  assign new_n164_ = ~new_n161_ & ~new_n163_;
  assign new_n165_ = ~new_n160_ & ~new_n164_;
  assign new_n166_ = v1 & v33;
  assign new_n167_ = ~v16 & ~new_n166_;
  assign new_n168_ = v24 & ~new_n92_;
  assign new_n169_ = ~v14 & v18;
  assign new_n170_ = ~v3 & new_n169_;
  assign new_n171_ = ~new_n168_ & ~new_n170_;
  assign new_n172_ = ~new_n167_ & ~new_n171_;
  assign new_n173_ = ~v20 & ~v32;
  assign new_n174_ = new_n104_ & new_n173_;
  assign new_n175_ = ~new_n161_ & ~new_n174_;
  assign new_n176_ = v24 & ~new_n175_;
  assign new_n177_ = v15 & new_n176_;
  assign new_n178_ = v16 & v27;
  assign new_n179_ = ~v14 & new_n178_;
  assign new_n180_ = ~new_n177_ & ~new_n179_;
  assign new_n181_ = ~new_n172_ & new_n180_;
  assign new_n182_ = ~new_n165_ & new_n181_;
  assign new_n183_ = ~new_n157_ & new_n182_;
  assign new_n184_ = v10 & ~new_n183_;
  assign new_n185_ = v3 & v22;
  assign new_n186_ = v2 & new_n185_;
  assign new_n187_ = ~v1 & v15;
  assign new_n188_ = v23 & v24;
  assign new_n189_ = ~v17 & new_n188_;
  assign new_n190_ = new_n187_ & new_n189_;
  assign new_n191_ = ~new_n186_ & ~new_n190_;
  assign new_n192_ = v19 & ~new_n191_;
  assign new_n193_ = ~v15 & ~v18;
  assign new_n194_ = v2 & ~new_n193_;
  assign new_n195_ = v18 & ~v19;
  assign new_n196_ = ~v1 & new_n195_;
  assign new_n197_ = v15 & v31;
  assign new_n198_ = ~new_n196_ & ~new_n197_;
  assign new_n199_ = ~new_n194_ & new_n198_;
  assign new_n200_ = v3 & ~new_n199_;
  assign new_n201_ = v11 & v24;
  assign new_n202_ = ~v8 & new_n201_;
  assign new_n203_ = v9 & ~v28;
  assign new_n204_ = ~v3 & new_n203_;
  assign new_n205_ = ~new_n202_ & ~new_n204_;
  assign new_n206_ = ~v1 & ~new_n205_;
  assign new_n207_ = v1 & v4;
  assign new_n208_ = v6 & new_n84_;
  assign new_n209_ = new_n207_ & new_n208_;
  assign new_n210_ = ~v8 & v24;
  assign new_n211_ = v29 & ~v30;
  assign new_n212_ = new_n210_ & new_n211_;
  assign new_n213_ = ~new_n209_ & ~new_n212_;
  assign new_n214_ = v11 & ~new_n213_;
  assign new_n215_ = ~v22 & ~v27;
  assign new_n216_ = ~v8 & ~new_n215_;
  assign new_n217_ = v18 & v20;
  assign new_n218_ = ~new_n216_ & ~new_n217_;
  assign new_n219_ = ~v30 & ~new_n218_;
  assign new_n220_ = v20 & v33;
  assign new_n221_ = v18 & new_n220_;
  assign new_n222_ = ~v15 & ~new_n221_;
  assign new_n223_ = ~new_n219_ & new_n222_;
  assign new_n224_ = v1 & ~new_n223_;
  assign new_n225_ = v18 & ~v30;
  assign new_n226_ = v17 & new_n225_;
  assign new_n227_ = ~new_n224_ & ~new_n226_;
  assign new_n228_ = v14 & ~new_n227_;
  assign new_n229_ = ~v6 & new_n154_;
  assign new_n230_ = ~v8 & ~v16;
  assign new_n231_ = v24 & v27;
  assign new_n232_ = new_n230_ & new_n231_;
  assign new_n233_ = ~new_n229_ & ~new_n232_;
  assign new_n234_ = ~new_n228_ & new_n233_;
  assign new_n235_ = ~new_n214_ & new_n234_;
  assign new_n236_ = ~new_n206_ & new_n235_;
  assign new_n237_ = ~new_n200_ & new_n236_;
  assign new_n238_ = ~new_n192_ & new_n237_;
  assign new_n239_ = ~new_n184_ & new_n238_;
  assign \v39.1  = new_n148_ | ~new_n239_;
  assign new_n241_ = ~v20 & ~new_n92_;
  assign new_n242_ = v1 & new_n241_;
  assign new_n243_ = v15 & ~v23;
  assign new_n244_ = v23 & v26;
  assign new_n245_ = ~new_n243_ & ~new_n244_;
  assign new_n246_ = v19 & ~new_n245_;
  assign new_n247_ = ~v1 & new_n246_;
  assign new_n248_ = ~new_n242_ & ~new_n247_;
  assign new_n249_ = ~v17 & ~new_n248_;
  assign new_n250_ = ~v1 & ~v17;
  assign new_n251_ = ~v33 & ~new_n250_;
  assign new_n252_ = ~v16 & ~new_n251_;
  assign new_n253_ = ~new_n92_ & ~new_n252_;
  assign new_n254_ = v1 & v11;
  assign new_n255_ = ~new_n253_ & ~new_n254_;
  assign new_n256_ = ~new_n249_ & new_n255_;
  assign new_n257_ = v24 & ~new_n256_;
  assign new_n258_ = ~v9 & ~v26;
  assign new_n259_ = ~v8 & v10;
  assign new_n260_ = ~new_n258_ & ~new_n259_;
  assign new_n261_ = v15 & ~new_n93_;
  assign new_n262_ = ~v10 & ~new_n76_;
  assign new_n263_ = ~v26 & ~new_n83_;
  assign new_n264_ = ~v12 & ~new_n263_;
  assign new_n265_ = v0 & v5;
  assign new_n266_ = v11 & ~v13;
  assign new_n267_ = ~new_n265_ & ~new_n266_;
  assign new_n268_ = v4 & ~new_n267_;
  assign new_n269_ = v11 & ~v25;
  assign new_n270_ = ~v4 & new_n269_;
  assign new_n271_ = ~new_n268_ & ~new_n270_;
  assign new_n272_ = ~new_n264_ & new_n271_;
  assign new_n273_ = ~new_n262_ & new_n272_;
  assign new_n274_ = ~new_n261_ & new_n273_;
  assign new_n275_ = ~new_n260_ & new_n274_;
  assign new_n276_ = v6 & ~new_n275_;
  assign new_n277_ = ~v9 & ~new_n53_;
  assign new_n278_ = ~new_n51_ & new_n277_;
  assign new_n279_ = ~v6 & ~new_n278_;
  assign new_n280_ = v33 & ~new_n95_;
  assign new_n281_ = v1 & ~new_n280_;
  assign new_n282_ = ~v16 & ~new_n281_;
  assign new_n283_ = ~v14 & ~new_n282_;
  assign new_n284_ = v17 & ~v33;
  assign new_n285_ = ~new_n283_ & ~new_n284_;
  assign new_n286_ = v18 & ~new_n285_;
  assign new_n287_ = ~new_n279_ & ~new_n286_;
  assign new_n288_ = ~v3 & ~new_n287_;
  assign new_n289_ = v22 & ~v23;
  assign new_n290_ = ~v27 & ~new_n289_;
  assign new_n291_ = v14 & ~new_n121_;
  assign new_n292_ = v14 & ~new_n291_;
  assign new_n293_ = ~new_n290_ & ~new_n292_;
  assign new_n294_ = ~v1 & ~v23;
  assign new_n295_ = ~v11 & ~v26;
  assign new_n296_ = ~new_n294_ & ~new_n295_;
  assign new_n297_ = v20 & ~v33;
  assign new_n298_ = ~v20 & v34;
  assign new_n299_ = ~v17 & new_n298_;
  assign new_n300_ = ~new_n297_ & ~new_n299_;
  assign new_n301_ = v18 & ~new_n300_;
  assign new_n302_ = v1 & new_n301_;
  assign new_n303_ = ~new_n296_ & ~new_n302_;
  assign new_n304_ = v14 & ~new_n303_;
  assign new_n305_ = ~new_n293_ & ~new_n304_;
  assign new_n306_ = ~new_n288_ & new_n305_;
  assign new_n307_ = ~new_n276_ & new_n306_;
  assign \v39.2  = new_n257_ | ~new_n307_;
  assign new_n309_ = v10 & ~v16;
  assign new_n310_ = v6 & new_n309_;
  assign new_n311_ = ~v14 & ~new_n310_;
  assign new_n312_ = ~v17 & ~new_n311_;
  assign new_n313_ = v3 & v31;
  assign new_n314_ = ~v2 & new_n313_;
  assign new_n315_ = ~new_n312_ & ~new_n314_;
  assign new_n316_ = v18 & ~new_n315_;
  assign \v39.3  = v1 & new_n316_;
  assign new_n318_ = ~v16 & v24;
  assign new_n319_ = v10 & v35;
  assign new_n320_ = v6 & new_n319_;
  assign new_n321_ = ~new_n318_ & ~new_n320_;
  assign new_n322_ = v20 & ~new_n321_;
  assign new_n323_ = ~v17 & new_n322_;
  assign new_n324_ = v1 & new_n323_;
  assign new_n325_ = v6 & v10;
  assign new_n326_ = v17 & v35;
  assign new_n327_ = new_n325_ & new_n326_;
  assign new_n328_ = ~new_n324_ & ~new_n327_;
  assign new_n329_ = v18 & ~new_n328_;
  assign new_n330_ = v20 & new_n168_;
  assign new_n331_ = ~v17 & new_n330_;
  assign new_n332_ = ~v16 & new_n331_;
  assign new_n333_ = v1 & new_n332_;
  assign \v39.4  = new_n329_ | new_n333_;
  assign new_n335_ = v8 & ~v16;
  assign new_n336_ = v24 & new_n335_;
  assign \v39.5  = v27 & new_n336_;
  assign \v39.6  = v27 & new_n77_;
  assign new_n339_ = ~v6 & v18;
  assign new_n340_ = ~v3 & new_n339_;
  assign new_n341_ = ~new_n168_ & ~new_n340_;
  assign new_n342_ = v36 & ~new_n341_;
  assign new_n343_ = v37 & v38;
  assign \v39.7  = new_n342_ | new_n343_;
endmodule


