// Benchmark "testing" written by ABC on Fri Feb 25 15:12:36 2022

module g25 ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A142, A141, A140, A139, A138, A109, A108, A107, A106, A105, A76, A75,
    A74, A73, A72, A43, A42, A41, A40, A39, A6, A7, A8, A9, A10  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A142, A141, A140, A139, A138, A109, A108, A107, A106, A105, A76, A75,
    A74, A73, A72, A43, A42, A41, A40, A39, A6, A7, A8, A9, A10;
  wire new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_,
    new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_,
    new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n115_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n131_, new_n132_, new_n133_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n160_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n176_, new_n177_, new_n178_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n221_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n237_, new_n238_, new_n239_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n282_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n298_,
    new_n299_, new_n300_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n342_, new_n343_,
    new_n345_, new_n346_, new_n348_, new_n349_;
  assign new_n51_ = A169 & A170;
  assign new_n52_ = ~A169 & ~A170;
  assign new_n53_ = ~new_n51_ & ~new_n52_;
  assign new_n54_ = ~A166 & A167;
  assign new_n55_ = A166 & ~A167;
  assign new_n56_ = ~new_n54_ & ~new_n55_;
  assign new_n57_ = ~A169 & ~new_n56_;
  assign new_n58_ = A169 & new_n56_;
  assign new_n59_ = ~new_n57_ & ~new_n58_;
  assign new_n60_ = new_n53_ & ~new_n59_;
  assign new_n61_ = A168 & ~new_n60_;
  assign new_n62_ = ~A168 & new_n60_;
  assign new_n63_ = ~new_n61_ & ~new_n62_;
  assign new_n64_ = ~new_n56_ & ~new_n63_;
  assign new_n65_ = A200 & ~A199;
  assign new_n66_ = ~A200 & A199;
  assign new_n67_ = ~new_n65_ & ~new_n66_;
  assign new_n68_ = ~A202 & new_n67_;
  assign new_n69_ = ~A203 & ~A202;
  assign new_n70_ = ~new_n68_ & ~new_n69_;
  assign new_n71_ = A201 & new_n70_;
  assign new_n72_ = ~A201 & ~new_n70_;
  assign new_n73_ = ~new_n71_ & ~new_n72_;
  assign new_n74_ = ~new_n67_ & ~new_n73_;
  assign new_n75_ = ~new_n64_ & new_n74_;
  assign new_n76_ = new_n64_ & ~new_n74_;
  assign new_n77_ = ~new_n75_ & ~new_n76_;
  assign new_n78_ = A233 & ~A232;
  assign new_n79_ = ~A233 & A232;
  assign new_n80_ = ~new_n78_ & ~new_n79_;
  assign new_n81_ = ~A235 & new_n80_;
  assign new_n82_ = ~A236 & ~A235;
  assign new_n83_ = ~new_n81_ & ~new_n82_;
  assign new_n84_ = A234 & new_n83_;
  assign new_n85_ = ~A234 & ~new_n83_;
  assign new_n86_ = ~new_n84_ & ~new_n85_;
  assign new_n87_ = ~new_n80_ & ~new_n86_;
  assign new_n88_ = A266 & ~A265;
  assign new_n89_ = ~A266 & A265;
  assign new_n90_ = ~new_n88_ & ~new_n89_;
  assign new_n91_ = ~A268 & new_n90_;
  assign new_n92_ = ~A269 & ~A268;
  assign new_n93_ = ~new_n91_ & ~new_n92_;
  assign new_n94_ = A267 & new_n93_;
  assign new_n95_ = ~A267 & ~new_n93_;
  assign new_n96_ = ~new_n94_ & ~new_n95_;
  assign new_n97_ = ~new_n90_ & ~new_n96_;
  assign new_n98_ = new_n77_ & ~new_n97_;
  assign new_n99_ = A299 & ~A298;
  assign new_n100_ = ~A299 & A298;
  assign new_n101_ = ~new_n99_ & ~new_n100_;
  assign new_n102_ = ~A301 & new_n101_;
  assign new_n103_ = ~A302 & ~A301;
  assign new_n104_ = ~new_n102_ & ~new_n103_;
  assign new_n105_ = A300 & new_n104_;
  assign new_n106_ = ~A300 & ~new_n104_;
  assign new_n107_ = ~new_n105_ & ~new_n106_;
  assign new_n108_ = ~new_n101_ & ~new_n107_;
  assign new_n109_ = ~new_n97_ & ~new_n108_;
  assign new_n110_ = ~new_n98_ & ~new_n109_;
  assign new_n111_ = new_n87_ & new_n110_;
  assign new_n112_ = ~new_n87_ & ~new_n110_;
  assign new_n113_ = ~new_n111_ & ~new_n112_;
  assign A142 = ~new_n77_ & ~new_n113_;
  assign new_n115_ = ~new_n74_ & ~new_n111_;
  assign A141 = ~new_n77_ & ~new_n115_;
  assign new_n117_ = new_n74_ & new_n87_;
  assign new_n118_ = ~new_n77_ & ~new_n117_;
  assign new_n119_ = new_n77_ & ~new_n118_;
  assign new_n120_ = new_n77_ & new_n117_;
  assign new_n121_ = new_n119_ & ~new_n120_;
  assign new_n122_ = new_n87_ & ~new_n121_;
  assign A140 = new_n110_ | new_n122_;
  assign new_n124_ = new_n97_ & new_n108_;
  assign new_n125_ = ~new_n109_ & ~new_n124_;
  assign new_n126_ = ~new_n77_ & ~new_n97_;
  assign new_n127_ = new_n77_ & new_n97_;
  assign new_n128_ = ~new_n126_ & ~new_n127_;
  assign new_n129_ = new_n125_ & ~new_n128_;
  assign A139 = new_n122_ | new_n129_;
  assign new_n131_ = new_n87_ & ~new_n129_;
  assign new_n132_ = ~new_n87_ & new_n129_;
  assign new_n133_ = ~new_n131_ & ~new_n132_;
  assign A138 = ~new_n77_ & ~new_n133_;
  assign new_n135_ = A167 & A168;
  assign new_n136_ = ~new_n56_ & ~new_n135_;
  assign new_n137_ = new_n56_ & ~new_n136_;
  assign new_n138_ = new_n56_ & new_n135_;
  assign new_n139_ = new_n137_ & ~new_n138_;
  assign new_n140_ = A168 & ~new_n139_;
  assign new_n141_ = ~new_n60_ & ~new_n140_;
  assign new_n142_ = ~A200 & ~new_n71_;
  assign new_n143_ = ~new_n67_ & ~new_n142_;
  assign new_n144_ = new_n141_ & new_n143_;
  assign new_n145_ = ~new_n141_ & ~new_n143_;
  assign new_n146_ = ~new_n144_ & ~new_n145_;
  assign new_n147_ = ~A233 & ~new_n84_;
  assign new_n148_ = ~new_n80_ & ~new_n147_;
  assign new_n149_ = ~A266 & ~new_n94_;
  assign new_n150_ = ~new_n90_ & ~new_n149_;
  assign new_n151_ = new_n146_ & ~new_n150_;
  assign new_n152_ = ~A299 & ~new_n105_;
  assign new_n153_ = ~new_n101_ & ~new_n152_;
  assign new_n154_ = ~new_n150_ & ~new_n153_;
  assign new_n155_ = ~new_n151_ & ~new_n154_;
  assign new_n156_ = new_n148_ & new_n155_;
  assign new_n157_ = ~new_n148_ & ~new_n155_;
  assign new_n158_ = ~new_n156_ & ~new_n157_;
  assign A109 = ~new_n146_ & ~new_n158_;
  assign new_n160_ = ~new_n143_ & ~new_n156_;
  assign A108 = ~new_n146_ & ~new_n160_;
  assign new_n162_ = new_n143_ & new_n148_;
  assign new_n163_ = ~new_n146_ & ~new_n162_;
  assign new_n164_ = new_n146_ & ~new_n163_;
  assign new_n165_ = new_n146_ & new_n162_;
  assign new_n166_ = new_n164_ & ~new_n165_;
  assign new_n167_ = new_n148_ & ~new_n166_;
  assign A107 = new_n155_ | new_n167_;
  assign new_n169_ = new_n150_ & new_n153_;
  assign new_n170_ = ~new_n154_ & ~new_n169_;
  assign new_n171_ = ~new_n146_ & ~new_n150_;
  assign new_n172_ = new_n146_ & new_n150_;
  assign new_n173_ = ~new_n171_ & ~new_n172_;
  assign new_n174_ = new_n170_ & ~new_n173_;
  assign A106 = new_n167_ | new_n174_;
  assign new_n176_ = new_n148_ & ~new_n174_;
  assign new_n177_ = ~new_n148_ & new_n174_;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign A105 = ~new_n146_ & ~new_n178_;
  assign new_n180_ = ~A169 & new_n56_;
  assign new_n181_ = ~new_n52_ & ~new_n180_;
  assign new_n182_ = ~new_n140_ & ~new_n181_;
  assign new_n183_ = A201 & A200;
  assign new_n184_ = ~new_n67_ & ~new_n183_;
  assign new_n185_ = new_n67_ & ~new_n184_;
  assign new_n186_ = new_n67_ & new_n183_;
  assign new_n187_ = new_n185_ & ~new_n186_;
  assign new_n188_ = A201 & ~new_n187_;
  assign new_n189_ = ~new_n70_ & ~new_n188_;
  assign new_n190_ = new_n182_ & ~new_n189_;
  assign new_n191_ = ~new_n182_ & new_n189_;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign new_n193_ = A234 & A233;
  assign new_n194_ = ~new_n80_ & ~new_n193_;
  assign new_n195_ = new_n80_ & ~new_n194_;
  assign new_n196_ = new_n80_ & new_n193_;
  assign new_n197_ = new_n195_ & ~new_n196_;
  assign new_n198_ = A234 & ~new_n197_;
  assign new_n199_ = ~new_n83_ & ~new_n198_;
  assign new_n200_ = A267 & A266;
  assign new_n201_ = ~new_n90_ & ~new_n200_;
  assign new_n202_ = new_n90_ & ~new_n201_;
  assign new_n203_ = new_n90_ & new_n200_;
  assign new_n204_ = new_n202_ & ~new_n203_;
  assign new_n205_ = A267 & ~new_n204_;
  assign new_n206_ = ~new_n93_ & ~new_n205_;
  assign new_n207_ = new_n192_ & new_n206_;
  assign new_n208_ = A300 & A299;
  assign new_n209_ = ~new_n101_ & ~new_n208_;
  assign new_n210_ = new_n101_ & ~new_n209_;
  assign new_n211_ = new_n101_ & new_n208_;
  assign new_n212_ = new_n210_ & ~new_n211_;
  assign new_n213_ = A300 & ~new_n212_;
  assign new_n214_ = ~new_n104_ & ~new_n213_;
  assign new_n215_ = new_n206_ & new_n214_;
  assign new_n216_ = ~new_n207_ & ~new_n215_;
  assign new_n217_ = ~new_n199_ & new_n216_;
  assign new_n218_ = new_n199_ & ~new_n216_;
  assign new_n219_ = ~new_n217_ & ~new_n218_;
  assign A76 = ~new_n192_ & ~new_n219_;
  assign new_n221_ = new_n189_ & ~new_n217_;
  assign A75 = ~new_n192_ & ~new_n221_;
  assign new_n223_ = ~new_n189_ & ~new_n199_;
  assign new_n224_ = ~new_n192_ & ~new_n223_;
  assign new_n225_ = new_n192_ & ~new_n224_;
  assign new_n226_ = new_n192_ & new_n223_;
  assign new_n227_ = new_n225_ & ~new_n226_;
  assign new_n228_ = ~new_n199_ & ~new_n227_;
  assign A74 = new_n216_ | new_n228_;
  assign new_n230_ = ~new_n206_ & ~new_n214_;
  assign new_n231_ = ~new_n215_ & ~new_n230_;
  assign new_n232_ = ~new_n192_ & new_n206_;
  assign new_n233_ = new_n192_ & ~new_n206_;
  assign new_n234_ = ~new_n232_ & ~new_n233_;
  assign new_n235_ = new_n231_ & ~new_n234_;
  assign A73 = new_n228_ | new_n235_;
  assign new_n237_ = ~new_n199_ & ~new_n235_;
  assign new_n238_ = new_n199_ & new_n235_;
  assign new_n239_ = ~new_n237_ & ~new_n238_;
  assign A72 = ~new_n192_ & ~new_n239_;
  assign new_n241_ = A168 & new_n181_;
  assign new_n242_ = ~A167 & ~new_n241_;
  assign new_n243_ = ~new_n56_ & ~new_n242_;
  assign new_n244_ = A203 & A202;
  assign new_n245_ = ~new_n69_ & ~new_n244_;
  assign new_n246_ = ~A202 & ~new_n67_;
  assign new_n247_ = A202 & new_n67_;
  assign new_n248_ = ~new_n246_ & ~new_n247_;
  assign new_n249_ = new_n245_ & ~new_n248_;
  assign new_n250_ = ~new_n188_ & ~new_n249_;
  assign new_n251_ = ~new_n243_ & ~new_n250_;
  assign new_n252_ = new_n243_ & new_n250_;
  assign new_n253_ = ~new_n251_ & ~new_n252_;
  assign new_n254_ = A236 & A235;
  assign new_n255_ = ~new_n82_ & ~new_n254_;
  assign new_n256_ = ~A235 & ~new_n80_;
  assign new_n257_ = A235 & new_n80_;
  assign new_n258_ = ~new_n256_ & ~new_n257_;
  assign new_n259_ = new_n255_ & ~new_n258_;
  assign new_n260_ = ~new_n198_ & ~new_n259_;
  assign new_n261_ = A269 & A268;
  assign new_n262_ = ~new_n92_ & ~new_n261_;
  assign new_n263_ = ~A268 & ~new_n90_;
  assign new_n264_ = A268 & new_n90_;
  assign new_n265_ = ~new_n263_ & ~new_n264_;
  assign new_n266_ = new_n262_ & ~new_n265_;
  assign new_n267_ = ~new_n205_ & ~new_n266_;
  assign new_n268_ = new_n253_ & new_n267_;
  assign new_n269_ = A302 & A301;
  assign new_n270_ = ~new_n103_ & ~new_n269_;
  assign new_n271_ = ~A301 & ~new_n101_;
  assign new_n272_ = A301 & new_n101_;
  assign new_n273_ = ~new_n271_ & ~new_n272_;
  assign new_n274_ = new_n270_ & ~new_n273_;
  assign new_n275_ = ~new_n213_ & ~new_n274_;
  assign new_n276_ = new_n267_ & new_n275_;
  assign new_n277_ = ~new_n268_ & ~new_n276_;
  assign new_n278_ = ~new_n260_ & new_n277_;
  assign new_n279_ = new_n260_ & ~new_n277_;
  assign new_n280_ = ~new_n278_ & ~new_n279_;
  assign A43 = ~new_n253_ & ~new_n280_;
  assign new_n282_ = new_n250_ & ~new_n278_;
  assign A42 = ~new_n253_ & ~new_n282_;
  assign new_n284_ = ~new_n250_ & ~new_n260_;
  assign new_n285_ = ~new_n253_ & ~new_n284_;
  assign new_n286_ = new_n253_ & ~new_n285_;
  assign new_n287_ = new_n253_ & new_n284_;
  assign new_n288_ = new_n286_ & ~new_n287_;
  assign new_n289_ = ~new_n260_ & ~new_n288_;
  assign A41 = new_n277_ | new_n289_;
  assign new_n291_ = ~new_n267_ & ~new_n275_;
  assign new_n292_ = ~new_n276_ & ~new_n291_;
  assign new_n293_ = ~new_n253_ & new_n267_;
  assign new_n294_ = new_n253_ & ~new_n267_;
  assign new_n295_ = ~new_n293_ & ~new_n294_;
  assign new_n296_ = new_n292_ & ~new_n295_;
  assign A40 = new_n289_ | new_n296_;
  assign new_n298_ = ~new_n260_ & ~new_n296_;
  assign new_n299_ = new_n260_ & new_n296_;
  assign new_n300_ = ~new_n298_ & ~new_n299_;
  assign A39 = ~new_n253_ & ~new_n300_;
  assign new_n302_ = A201 & ~new_n249_;
  assign new_n303_ = ~A201 & new_n249_;
  assign new_n304_ = ~new_n302_ & ~new_n303_;
  assign new_n305_ = ~new_n67_ & ~new_n304_;
  assign new_n306_ = ~A168 & ~new_n181_;
  assign new_n307_ = ~new_n241_ & ~new_n306_;
  assign new_n308_ = ~new_n56_ & ~new_n307_;
  assign new_n309_ = new_n305_ & new_n308_;
  assign new_n310_ = ~new_n305_ & ~new_n308_;
  assign new_n311_ = ~new_n309_ & ~new_n310_;
  assign new_n312_ = A300 & ~new_n274_;
  assign new_n313_ = ~A300 & new_n274_;
  assign new_n314_ = ~new_n312_ & ~new_n313_;
  assign new_n315_ = ~new_n101_ & ~new_n314_;
  assign new_n316_ = A267 & ~new_n266_;
  assign new_n317_ = ~A267 & new_n266_;
  assign new_n318_ = ~new_n316_ & ~new_n317_;
  assign new_n319_ = ~new_n90_ & ~new_n318_;
  assign new_n320_ = ~new_n315_ & new_n319_;
  assign new_n321_ = new_n315_ & ~new_n319_;
  assign new_n322_ = ~new_n320_ & ~new_n321_;
  assign new_n323_ = ~new_n305_ & ~new_n322_;
  assign new_n324_ = new_n305_ & new_n322_;
  assign new_n325_ = ~new_n323_ & ~new_n324_;
  assign new_n326_ = new_n311_ & ~new_n325_;
  assign new_n327_ = A234 & ~new_n259_;
  assign new_n328_ = ~A234 & new_n259_;
  assign new_n329_ = ~new_n327_ & ~new_n328_;
  assign new_n330_ = ~new_n80_ & ~new_n329_;
  assign new_n331_ = ~new_n326_ & new_n330_;
  assign new_n332_ = new_n326_ & ~new_n330_;
  assign new_n333_ = ~new_n331_ & ~new_n332_;
  assign A6 = ~new_n322_ & ~new_n333_;
  assign new_n335_ = new_n319_ & new_n330_;
  assign new_n336_ = ~new_n322_ & ~new_n335_;
  assign new_n337_ = new_n322_ & ~new_n336_;
  assign new_n338_ = new_n322_ & new_n335_;
  assign new_n339_ = new_n337_ & ~new_n338_;
  assign new_n340_ = new_n330_ & ~new_n339_;
  assign A7 = new_n326_ | new_n340_;
  assign new_n342_ = ~new_n305_ & new_n322_;
  assign new_n343_ = ~new_n310_ & ~new_n342_;
  assign A8 = new_n340_ | new_n343_;
  assign new_n345_ = new_n330_ & new_n343_;
  assign new_n346_ = ~new_n319_ & ~new_n345_;
  assign A9 = ~new_n322_ & ~new_n346_;
  assign new_n348_ = ~new_n330_ & ~new_n343_;
  assign new_n349_ = ~new_n345_ & ~new_n348_;
  assign A10 = ~new_n322_ & ~new_n349_;
endmodule


