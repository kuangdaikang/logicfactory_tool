// Benchmark "arbiter" written by ABC on Thu Sep 14 22:38:55 2023

module arbiter ( 
    \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ,
    \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] , \grant[5] ,
    \grant[6] , \grant[7] , \grant[8] , \grant[9] , \grant[10] ,
    \grant[11] , \grant[12] , \grant[13] , \grant[14] , \grant[15] ,
    \grant[16] , \grant[17] , \grant[18] , \grant[19] , \grant[20] ,
    \grant[21] , \grant[22] , \grant[23] , \grant[24] , \grant[25] ,
    \grant[26] , \grant[27] , \grant[28] , \grant[29] , \grant[30] ,
    \grant[31] , \grant[32] , \grant[33] , \grant[34] , \grant[35] ,
    \grant[36] , \grant[37] , \grant[38] , \grant[39] , \grant[40] ,
    \grant[41] , \grant[42] , \grant[43] , \grant[44] , \grant[45] ,
    \grant[46] , \grant[47] , \grant[48] , \grant[49] , \grant[50] ,
    \grant[51] , \grant[52] , \grant[53] , \grant[54] , \grant[55] ,
    \grant[56] , \grant[57] , \grant[58] , \grant[59] , \grant[60] ,
    \grant[61] , \grant[62] , \grant[63] , \grant[64] , \grant[65] ,
    \grant[66] , \grant[67] , \grant[68] , \grant[69] , \grant[70] ,
    \grant[71] , \grant[72] , \grant[73] , \grant[74] , \grant[75] ,
    \grant[76] , \grant[77] , \grant[78] , \grant[79] , \grant[80] ,
    \grant[81] , \grant[82] , \grant[83] , \grant[84] , \grant[85] ,
    \grant[86] , \grant[87] , \grant[88] , \grant[89] , \grant[90] ,
    \grant[91] , \grant[92] , \grant[93] , \grant[94] , \grant[95] ,
    \grant[96] , \grant[97] , \grant[98] , \grant[99] , \grant[100] ,
    \grant[101] , \grant[102] , \grant[103] , \grant[104] , \grant[105] ,
    \grant[106] , \grant[107] , \grant[108] , \grant[109] , \grant[110] ,
    \grant[111] , \grant[112] , \grant[113] , \grant[114] , \grant[115] ,
    \grant[116] , \grant[117] , \grant[118] , \grant[119] , \grant[120] ,
    \grant[121] , \grant[122] , \grant[123] , \grant[124] , \grant[125] ,
    \grant[126] , \grant[127] , anyGrant  );
  input  \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ;
  output \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] ,
    \grant[5] , \grant[6] , \grant[7] , \grant[8] , \grant[9] ,
    \grant[10] , \grant[11] , \grant[12] , \grant[13] , \grant[14] ,
    \grant[15] , \grant[16] , \grant[17] , \grant[18] , \grant[19] ,
    \grant[20] , \grant[21] , \grant[22] , \grant[23] , \grant[24] ,
    \grant[25] , \grant[26] , \grant[27] , \grant[28] , \grant[29] ,
    \grant[30] , \grant[31] , \grant[32] , \grant[33] , \grant[34] ,
    \grant[35] , \grant[36] , \grant[37] , \grant[38] , \grant[39] ,
    \grant[40] , \grant[41] , \grant[42] , \grant[43] , \grant[44] ,
    \grant[45] , \grant[46] , \grant[47] , \grant[48] , \grant[49] ,
    \grant[50] , \grant[51] , \grant[52] , \grant[53] , \grant[54] ,
    \grant[55] , \grant[56] , \grant[57] , \grant[58] , \grant[59] ,
    \grant[60] , \grant[61] , \grant[62] , \grant[63] , \grant[64] ,
    \grant[65] , \grant[66] , \grant[67] , \grant[68] , \grant[69] ,
    \grant[70] , \grant[71] , \grant[72] , \grant[73] , \grant[74] ,
    \grant[75] , \grant[76] , \grant[77] , \grant[78] , \grant[79] ,
    \grant[80] , \grant[81] , \grant[82] , \grant[83] , \grant[84] ,
    \grant[85] , \grant[86] , \grant[87] , \grant[88] , \grant[89] ,
    \grant[90] , \grant[91] , \grant[92] , \grant[93] , \grant[94] ,
    \grant[95] , \grant[96] , \grant[97] , \grant[98] , \grant[99] ,
    \grant[100] , \grant[101] , \grant[102] , \grant[103] , \grant[104] ,
    \grant[105] , \grant[106] , \grant[107] , \grant[108] , \grant[109] ,
    \grant[110] , \grant[111] , \grant[112] , \grant[113] , \grant[114] ,
    \grant[115] , \grant[116] , \grant[117] , \grant[118] , \grant[119] ,
    \grant[120] , \grant[121] , \grant[122] , \grant[123] , \grant[124] ,
    \grant[125] , \grant[126] , \grant[127] , anyGrant;
  wire new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_,
    new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1739_, new_n1740_, new_n1741_,
    new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_,
    new_n1748_, new_n1749_, new_n1750_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1893_, new_n1894_,
    new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1949_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1960_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1968_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2020_, new_n2021_,
    new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_,
    new_n2028_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2058_, new_n2059_, new_n2060_, new_n2061_,
    new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2118_, new_n2119_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2186_, new_n2187_, new_n2188_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_,
    new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2234_, new_n2235_,
    new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_,
    new_n2242_, new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_,
    new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2294_, new_n2295_,
    new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_,
    new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_,
    new_n2309_, new_n2310_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2352_, new_n2353_, new_n2354_, new_n2355_,
    new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2408_, new_n2409_,
    new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_,
    new_n2416_, new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_,
    new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2448_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2466_, new_n2467_, new_n2468_, new_n2469_,
    new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2514_, new_n2515_, new_n2516_,
    new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_,
    new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_,
    new_n2530_, new_n2531_, new_n2532_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2562_, new_n2563_,
    new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2570_,
    new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_,
    new_n2577_, new_n2578_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2620_, new_n2621_, new_n2622_, new_n2623_,
    new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2630_,
    new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_,
    new_n2637_, new_n2638_, new_n2640_, new_n2641_, new_n2642_, new_n2643_,
    new_n2644_, new_n2645_, new_n2646_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2683_, new_n2684_,
    new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2735_, new_n2736_, new_n2737_, new_n2738_,
    new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2802_, new_n2803_, new_n2804_,
    new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_,
    new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_,
    new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_;
  INV_X1     g0000(.I(\req[0] ), .ZN(new_n386_));
  NOR2_X1    g0001(.A1(\priority[79] ), .A2(\priority[80] ), .ZN(new_n387_));
  NAND2_X1   g0002(.A1(\priority[78] ), .A2(\req[78] ), .ZN(new_n388_));
  NOR2_X1    g0003(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1    g0004(.A1(\req[80] ), .A2(\req[81] ), .ZN(new_n390_));
  NAND2_X1   g0005(.A1(\priority[80] ), .A2(\req[79] ), .ZN(new_n391_));
  NOR2_X1    g0006(.A1(\priority[82] ), .A2(\priority[83] ), .ZN(new_n392_));
  NAND2_X1   g0007(.A1(\priority[81] ), .A2(\req[81] ), .ZN(new_n393_));
  NOR4_X1    g0008(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .A4(new_n393_), .ZN(new_n394_));
  NOR2_X1    g0009(.A1(\req[83] ), .A2(\req[84] ), .ZN(new_n395_));
  NAND2_X1   g0010(.A1(\priority[83] ), .A2(\req[82] ), .ZN(new_n396_));
  NOR2_X1    g0011(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1    g0012(.A1(\priority[85] ), .A2(\priority[86] ), .ZN(new_n398_));
  NAND2_X1   g0013(.A1(\priority[84] ), .A2(\req[84] ), .ZN(new_n399_));
  NOR2_X1    g0014(.A1(\req[86] ), .A2(\req[87] ), .ZN(new_n400_));
  NAND2_X1   g0015(.A1(\priority[86] ), .A2(\req[85] ), .ZN(new_n401_));
  NOR4_X1    g0016(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  OAI22_X1   g0017(.A1(new_n389_), .A2(new_n394_), .B1(new_n402_), .B2(new_n397_), .ZN(new_n403_));
  NOR2_X1    g0018(.A1(\priority[88] ), .A2(\priority[89] ), .ZN(new_n404_));
  NAND2_X1   g0019(.A1(\priority[87] ), .A2(\req[87] ), .ZN(new_n405_));
  NOR2_X1    g0020(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1    g0021(.A1(\req[89] ), .A2(\req[90] ), .ZN(new_n407_));
  NAND2_X1   g0022(.A1(\priority[89] ), .A2(\req[88] ), .ZN(new_n408_));
  NOR2_X1    g0023(.A1(\priority[91] ), .A2(\priority[92] ), .ZN(new_n409_));
  NAND2_X1   g0024(.A1(\priority[90] ), .A2(\req[90] ), .ZN(new_n410_));
  NOR4_X1    g0025(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n411_));
  NOR2_X1    g0026(.A1(\req[92] ), .A2(\req[93] ), .ZN(new_n412_));
  NAND2_X1   g0027(.A1(\priority[92] ), .A2(\req[91] ), .ZN(new_n413_));
  NOR2_X1    g0028(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1    g0029(.A1(\priority[94] ), .A2(\priority[95] ), .ZN(new_n415_));
  NAND2_X1   g0030(.A1(\priority[93] ), .A2(\req[93] ), .ZN(new_n416_));
  NOR2_X1    g0031(.A1(\req[95] ), .A2(\req[96] ), .ZN(new_n417_));
  NAND2_X1   g0032(.A1(\priority[95] ), .A2(\req[94] ), .ZN(new_n418_));
  NOR4_X1    g0033(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n419_));
  OAI22_X1   g0034(.A1(new_n406_), .A2(new_n411_), .B1(new_n419_), .B2(new_n414_), .ZN(new_n420_));
  NOR2_X1    g0035(.A1(\priority[61] ), .A2(\priority[62] ), .ZN(new_n421_));
  NAND2_X1   g0036(.A1(\priority[60] ), .A2(\req[60] ), .ZN(new_n422_));
  NOR2_X1    g0037(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1    g0038(.A1(\req[62] ), .A2(\req[63] ), .ZN(new_n424_));
  NAND2_X1   g0039(.A1(\priority[62] ), .A2(\req[61] ), .ZN(new_n425_));
  NOR2_X1    g0040(.A1(\priority[64] ), .A2(\priority[65] ), .ZN(new_n426_));
  NAND2_X1   g0041(.A1(\priority[63] ), .A2(\req[63] ), .ZN(new_n427_));
  NOR4_X1    g0042(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .A4(new_n427_), .ZN(new_n428_));
  NOR2_X1    g0043(.A1(\req[65] ), .A2(\req[66] ), .ZN(new_n429_));
  NAND2_X1   g0044(.A1(\priority[65] ), .A2(\req[64] ), .ZN(new_n430_));
  NOR2_X1    g0045(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NOR2_X1    g0046(.A1(\priority[67] ), .A2(\priority[68] ), .ZN(new_n432_));
  NAND2_X1   g0047(.A1(\priority[66] ), .A2(\req[66] ), .ZN(new_n433_));
  NOR2_X1    g0048(.A1(\req[68] ), .A2(\req[69] ), .ZN(new_n434_));
  NAND2_X1   g0049(.A1(\priority[68] ), .A2(\req[67] ), .ZN(new_n435_));
  NOR4_X1    g0050(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .A4(new_n435_), .ZN(new_n436_));
  OAI22_X1   g0051(.A1(new_n423_), .A2(new_n428_), .B1(new_n436_), .B2(new_n431_), .ZN(new_n437_));
  NOR2_X1    g0052(.A1(\priority[70] ), .A2(\priority[71] ), .ZN(new_n438_));
  NAND2_X1   g0053(.A1(\priority[69] ), .A2(\req[69] ), .ZN(new_n439_));
  NOR2_X1    g0054(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1    g0055(.A1(\req[71] ), .A2(\req[72] ), .ZN(new_n441_));
  NAND2_X1   g0056(.A1(\priority[71] ), .A2(\req[70] ), .ZN(new_n442_));
  NOR2_X1    g0057(.A1(\priority[73] ), .A2(\priority[74] ), .ZN(new_n443_));
  NAND2_X1   g0058(.A1(\priority[72] ), .A2(\req[72] ), .ZN(new_n444_));
  NOR4_X1    g0059(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .A4(new_n444_), .ZN(new_n445_));
  NOR2_X1    g0060(.A1(\req[74] ), .A2(\req[75] ), .ZN(new_n446_));
  NAND2_X1   g0061(.A1(\priority[74] ), .A2(\req[73] ), .ZN(new_n447_));
  NOR2_X1    g0062(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1    g0063(.A1(\priority[76] ), .A2(\priority[77] ), .ZN(new_n449_));
  NAND2_X1   g0064(.A1(\priority[75] ), .A2(\req[75] ), .ZN(new_n450_));
  NOR2_X1    g0065(.A1(\req[77] ), .A2(\req[78] ), .ZN(new_n451_));
  NAND2_X1   g0066(.A1(\priority[77] ), .A2(\req[76] ), .ZN(new_n452_));
  NOR4_X1    g0067(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .A4(new_n452_), .ZN(new_n453_));
  OAI22_X1   g0068(.A1(new_n440_), .A2(new_n445_), .B1(new_n453_), .B2(new_n448_), .ZN(new_n454_));
  NOR4_X1    g0069(.A1(new_n403_), .A2(new_n420_), .A3(new_n437_), .A4(new_n454_), .ZN(new_n455_));
  NOR2_X1    g0070(.A1(\priority[124] ), .A2(\priority[125] ), .ZN(new_n456_));
  NAND2_X1   g0071(.A1(\priority[123] ), .A2(\req[123] ), .ZN(new_n457_));
  NOR2_X1    g0072(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1    g0073(.A1(\req[125] ), .A2(\req[126] ), .ZN(new_n459_));
  NAND2_X1   g0074(.A1(\priority[125] ), .A2(\req[124] ), .ZN(new_n460_));
  NOR2_X1    g0075(.A1(\priority[0] ), .A2(\priority[127] ), .ZN(new_n461_));
  NAND2_X1   g0076(.A1(\priority[126] ), .A2(\req[126] ), .ZN(new_n462_));
  NOR4_X1    g0077(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  NOR2_X1    g0078(.A1(new_n463_), .A2(new_n458_), .ZN(new_n464_));
  NOR2_X1    g0079(.A1(\priority[115] ), .A2(\priority[116] ), .ZN(new_n465_));
  NAND2_X1   g0080(.A1(\priority[114] ), .A2(\req[114] ), .ZN(new_n466_));
  NOR2_X1    g0081(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NOR2_X1    g0082(.A1(\req[116] ), .A2(\req[117] ), .ZN(new_n468_));
  NAND2_X1   g0083(.A1(\priority[116] ), .A2(\req[115] ), .ZN(new_n469_));
  NOR2_X1    g0084(.A1(\priority[118] ), .A2(\priority[119] ), .ZN(new_n470_));
  NAND2_X1   g0085(.A1(\priority[117] ), .A2(\req[117] ), .ZN(new_n471_));
  NOR4_X1    g0086(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .A4(new_n471_), .ZN(new_n472_));
  NOR2_X1    g0087(.A1(\req[119] ), .A2(\req[120] ), .ZN(new_n473_));
  NAND2_X1   g0088(.A1(\priority[119] ), .A2(\req[118] ), .ZN(new_n474_));
  NOR2_X1    g0089(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1    g0090(.A1(\priority[121] ), .A2(\priority[122] ), .ZN(new_n476_));
  NAND2_X1   g0091(.A1(\priority[120] ), .A2(\req[120] ), .ZN(new_n477_));
  NOR2_X1    g0092(.A1(\req[122] ), .A2(\req[123] ), .ZN(new_n478_));
  NAND2_X1   g0093(.A1(\priority[122] ), .A2(\req[121] ), .ZN(new_n479_));
  NOR4_X1    g0094(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .A4(new_n479_), .ZN(new_n480_));
  OAI22_X1   g0095(.A1(new_n467_), .A2(new_n472_), .B1(new_n480_), .B2(new_n475_), .ZN(new_n481_));
  NOR2_X1    g0096(.A1(\priority[97] ), .A2(\priority[98] ), .ZN(new_n482_));
  NAND2_X1   g0097(.A1(\priority[96] ), .A2(\req[96] ), .ZN(new_n483_));
  NOR2_X1    g0098(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NOR2_X1    g0099(.A1(\req[98] ), .A2(\req[99] ), .ZN(new_n485_));
  NAND2_X1   g0100(.A1(\priority[98] ), .A2(\req[97] ), .ZN(new_n486_));
  NOR2_X1    g0101(.A1(\priority[100] ), .A2(\priority[101] ), .ZN(new_n487_));
  NAND2_X1   g0102(.A1(\priority[99] ), .A2(\req[99] ), .ZN(new_n488_));
  NOR4_X1    g0103(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .A4(new_n488_), .ZN(new_n489_));
  NOR2_X1    g0104(.A1(\req[101] ), .A2(\req[102] ), .ZN(new_n490_));
  NAND2_X1   g0105(.A1(\priority[101] ), .A2(\req[100] ), .ZN(new_n491_));
  NOR2_X1    g0106(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1    g0107(.A1(\priority[103] ), .A2(\priority[104] ), .ZN(new_n493_));
  NAND2_X1   g0108(.A1(\priority[102] ), .A2(\req[102] ), .ZN(new_n494_));
  NOR2_X1    g0109(.A1(\req[104] ), .A2(\req[105] ), .ZN(new_n495_));
  NAND2_X1   g0110(.A1(\priority[104] ), .A2(\req[103] ), .ZN(new_n496_));
  NOR4_X1    g0111(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .A4(new_n496_), .ZN(new_n497_));
  OAI22_X1   g0112(.A1(new_n484_), .A2(new_n489_), .B1(new_n497_), .B2(new_n492_), .ZN(new_n498_));
  NOR2_X1    g0113(.A1(\priority[106] ), .A2(\priority[107] ), .ZN(new_n499_));
  NAND2_X1   g0114(.A1(\priority[105] ), .A2(\req[105] ), .ZN(new_n500_));
  NOR2_X1    g0115(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1    g0116(.A1(\req[107] ), .A2(\req[108] ), .ZN(new_n502_));
  NAND2_X1   g0117(.A1(\priority[107] ), .A2(\req[106] ), .ZN(new_n503_));
  NOR2_X1    g0118(.A1(\priority[109] ), .A2(\priority[110] ), .ZN(new_n504_));
  NAND2_X1   g0119(.A1(\priority[108] ), .A2(\req[108] ), .ZN(new_n505_));
  NOR4_X1    g0120(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  NOR2_X1    g0121(.A1(\req[110] ), .A2(\req[111] ), .ZN(new_n507_));
  NAND2_X1   g0122(.A1(\priority[110] ), .A2(\req[109] ), .ZN(new_n508_));
  NOR2_X1    g0123(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1    g0124(.A1(\priority[112] ), .A2(\priority[113] ), .ZN(new_n510_));
  NAND2_X1   g0125(.A1(\priority[111] ), .A2(\req[111] ), .ZN(new_n511_));
  NOR2_X1    g0126(.A1(\req[113] ), .A2(\req[114] ), .ZN(new_n512_));
  NAND2_X1   g0127(.A1(\priority[113] ), .A2(\req[112] ), .ZN(new_n513_));
  NOR4_X1    g0128(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n514_));
  OAI22_X1   g0129(.A1(new_n501_), .A2(new_n506_), .B1(new_n514_), .B2(new_n509_), .ZN(new_n515_));
  NOR4_X1    g0130(.A1(new_n481_), .A2(new_n498_), .A3(new_n515_), .A4(new_n464_), .ZN(new_n516_));
  NOR2_X1    g0131(.A1(\req[2] ), .A2(\req[3] ), .ZN(new_n517_));
  NOR2_X1    g0132(.A1(\priority[4] ), .A2(\priority[5] ), .ZN(new_n518_));
  NAND2_X1   g0133(.A1(\priority[3] ), .A2(\req[3] ), .ZN(new_n519_));
  NOR2_X1    g0134(.A1(\req[5] ), .A2(\req[6] ), .ZN(new_n520_));
  NAND2_X1   g0135(.A1(\priority[5] ), .A2(\req[4] ), .ZN(new_n521_));
  NOR4_X1    g0136(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .A4(new_n521_), .ZN(new_n522_));
  INV_X1     g0137(.I(\req[1] ), .ZN(new_n523_));
  AOI21_X1   g0138(.A1(new_n523_), .A2(\priority[1] ), .B(\priority[2] ), .ZN(new_n524_));
  OAI21_X1   g0139(.A1(new_n522_), .A2(new_n517_), .B(new_n524_), .ZN(new_n525_));
  NOR2_X1    g0140(.A1(\priority[7] ), .A2(\priority[8] ), .ZN(new_n526_));
  NAND2_X1   g0141(.A1(\priority[6] ), .A2(\req[6] ), .ZN(new_n527_));
  NOR2_X1    g0142(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1    g0143(.A1(\req[8] ), .A2(\req[9] ), .ZN(new_n529_));
  NAND2_X1   g0144(.A1(\priority[8] ), .A2(\req[7] ), .ZN(new_n530_));
  NOR2_X1    g0145(.A1(\priority[10] ), .A2(\priority[11] ), .ZN(new_n531_));
  NAND2_X1   g0146(.A1(\priority[9] ), .A2(\req[9] ), .ZN(new_n532_));
  NOR4_X1    g0147(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  NOR2_X1    g0148(.A1(\req[11] ), .A2(\req[12] ), .ZN(new_n534_));
  NAND2_X1   g0149(.A1(\priority[11] ), .A2(\req[10] ), .ZN(new_n535_));
  NOR2_X1    g0150(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1    g0151(.A1(\priority[13] ), .A2(\priority[14] ), .ZN(new_n537_));
  NAND2_X1   g0152(.A1(\priority[12] ), .A2(\req[12] ), .ZN(new_n538_));
  NOR2_X1    g0153(.A1(\req[14] ), .A2(\req[15] ), .ZN(new_n539_));
  NAND2_X1   g0154(.A1(\priority[14] ), .A2(\req[13] ), .ZN(new_n540_));
  NOR4_X1    g0155(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .A4(new_n540_), .ZN(new_n541_));
  OAI22_X1   g0156(.A1(new_n528_), .A2(new_n533_), .B1(new_n541_), .B2(new_n536_), .ZN(new_n542_));
  NOR2_X1    g0157(.A1(\priority[16] ), .A2(\priority[17] ), .ZN(new_n543_));
  NAND2_X1   g0158(.A1(\priority[15] ), .A2(\req[15] ), .ZN(new_n544_));
  NOR2_X1    g0159(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1    g0160(.A1(\req[17] ), .A2(\req[18] ), .ZN(new_n546_));
  NAND2_X1   g0161(.A1(\priority[17] ), .A2(\req[16] ), .ZN(new_n547_));
  NOR2_X1    g0162(.A1(\priority[19] ), .A2(\priority[20] ), .ZN(new_n548_));
  NAND2_X1   g0163(.A1(\priority[18] ), .A2(\req[18] ), .ZN(new_n549_));
  NOR4_X1    g0164(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .A4(new_n549_), .ZN(new_n550_));
  NOR2_X1    g0165(.A1(\req[20] ), .A2(\req[21] ), .ZN(new_n551_));
  NAND2_X1   g0166(.A1(\priority[20] ), .A2(\req[19] ), .ZN(new_n552_));
  NOR2_X1    g0167(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1    g0168(.A1(\priority[22] ), .A2(\priority[23] ), .ZN(new_n554_));
  NAND2_X1   g0169(.A1(\priority[21] ), .A2(\req[21] ), .ZN(new_n555_));
  NOR2_X1    g0170(.A1(\req[23] ), .A2(\req[24] ), .ZN(new_n556_));
  NAND2_X1   g0171(.A1(\priority[23] ), .A2(\req[22] ), .ZN(new_n557_));
  NOR4_X1    g0172(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .A4(new_n557_), .ZN(new_n558_));
  OAI22_X1   g0173(.A1(new_n545_), .A2(new_n550_), .B1(new_n558_), .B2(new_n553_), .ZN(new_n559_));
  NOR3_X1    g0174(.A1(new_n542_), .A2(new_n559_), .A3(new_n525_), .ZN(new_n560_));
  NOR2_X1    g0175(.A1(\priority[43] ), .A2(\priority[44] ), .ZN(new_n561_));
  NAND2_X1   g0176(.A1(\priority[42] ), .A2(\req[42] ), .ZN(new_n562_));
  NOR2_X1    g0177(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1    g0178(.A1(\req[44] ), .A2(\req[45] ), .ZN(new_n564_));
  NAND2_X1   g0179(.A1(\priority[44] ), .A2(\req[43] ), .ZN(new_n565_));
  NOR2_X1    g0180(.A1(\priority[46] ), .A2(\priority[47] ), .ZN(new_n566_));
  NAND2_X1   g0181(.A1(\priority[45] ), .A2(\req[45] ), .ZN(new_n567_));
  NOR4_X1    g0182(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n568_));
  NOR2_X1    g0183(.A1(\req[47] ), .A2(\req[48] ), .ZN(new_n569_));
  NAND2_X1   g0184(.A1(\priority[47] ), .A2(\req[46] ), .ZN(new_n570_));
  NOR2_X1    g0185(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1    g0186(.A1(\priority[49] ), .A2(\priority[50] ), .ZN(new_n572_));
  NAND2_X1   g0187(.A1(\priority[48] ), .A2(\req[48] ), .ZN(new_n573_));
  NOR2_X1    g0188(.A1(\req[50] ), .A2(\req[51] ), .ZN(new_n574_));
  NAND2_X1   g0189(.A1(\priority[50] ), .A2(\req[49] ), .ZN(new_n575_));
  NOR4_X1    g0190(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n576_));
  OAI22_X1   g0191(.A1(new_n563_), .A2(new_n568_), .B1(new_n576_), .B2(new_n571_), .ZN(new_n577_));
  NOR2_X1    g0192(.A1(\priority[52] ), .A2(\priority[53] ), .ZN(new_n578_));
  NAND2_X1   g0193(.A1(\priority[51] ), .A2(\req[51] ), .ZN(new_n579_));
  NOR2_X1    g0194(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1    g0195(.A1(\req[53] ), .A2(\req[54] ), .ZN(new_n581_));
  NAND2_X1   g0196(.A1(\priority[53] ), .A2(\req[52] ), .ZN(new_n582_));
  NOR2_X1    g0197(.A1(\priority[55] ), .A2(\priority[56] ), .ZN(new_n583_));
  NAND2_X1   g0198(.A1(\priority[54] ), .A2(\req[54] ), .ZN(new_n584_));
  NOR4_X1    g0199(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n585_));
  NOR2_X1    g0200(.A1(\req[56] ), .A2(\req[57] ), .ZN(new_n586_));
  NAND2_X1   g0201(.A1(\priority[56] ), .A2(\req[55] ), .ZN(new_n587_));
  NOR2_X1    g0202(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1    g0203(.A1(\priority[58] ), .A2(\priority[59] ), .ZN(new_n589_));
  NAND2_X1   g0204(.A1(\priority[57] ), .A2(\req[57] ), .ZN(new_n590_));
  NOR2_X1    g0205(.A1(\req[59] ), .A2(\req[60] ), .ZN(new_n591_));
  NAND2_X1   g0206(.A1(\priority[59] ), .A2(\req[58] ), .ZN(new_n592_));
  NOR4_X1    g0207(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .A4(new_n592_), .ZN(new_n593_));
  OAI22_X1   g0208(.A1(new_n580_), .A2(new_n585_), .B1(new_n593_), .B2(new_n588_), .ZN(new_n594_));
  NOR2_X1    g0209(.A1(\priority[25] ), .A2(\priority[26] ), .ZN(new_n595_));
  NAND2_X1   g0210(.A1(\priority[24] ), .A2(\req[24] ), .ZN(new_n596_));
  NOR2_X1    g0211(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1    g0212(.A1(\req[26] ), .A2(\req[27] ), .ZN(new_n598_));
  NAND2_X1   g0213(.A1(\priority[26] ), .A2(\req[25] ), .ZN(new_n599_));
  NOR2_X1    g0214(.A1(\priority[28] ), .A2(\priority[29] ), .ZN(new_n600_));
  NAND2_X1   g0215(.A1(\priority[27] ), .A2(\req[27] ), .ZN(new_n601_));
  NOR4_X1    g0216(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .A4(new_n601_), .ZN(new_n602_));
  NOR2_X1    g0217(.A1(\req[29] ), .A2(\req[30] ), .ZN(new_n603_));
  NAND2_X1   g0218(.A1(\priority[29] ), .A2(\req[28] ), .ZN(new_n604_));
  NOR2_X1    g0219(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1    g0220(.A1(\priority[31] ), .A2(\priority[32] ), .ZN(new_n606_));
  NAND2_X1   g0221(.A1(\priority[30] ), .A2(\req[30] ), .ZN(new_n607_));
  NOR2_X1    g0222(.A1(\req[32] ), .A2(\req[33] ), .ZN(new_n608_));
  NAND2_X1   g0223(.A1(\priority[32] ), .A2(\req[31] ), .ZN(new_n609_));
  NOR4_X1    g0224(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .A4(new_n609_), .ZN(new_n610_));
  OAI22_X1   g0225(.A1(new_n597_), .A2(new_n602_), .B1(new_n610_), .B2(new_n605_), .ZN(new_n611_));
  NOR2_X1    g0226(.A1(\priority[34] ), .A2(\priority[35] ), .ZN(new_n612_));
  NAND2_X1   g0227(.A1(\priority[33] ), .A2(\req[33] ), .ZN(new_n613_));
  NOR2_X1    g0228(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1    g0229(.A1(\req[35] ), .A2(\req[36] ), .ZN(new_n615_));
  NAND2_X1   g0230(.A1(\priority[35] ), .A2(\req[34] ), .ZN(new_n616_));
  NOR2_X1    g0231(.A1(\priority[37] ), .A2(\priority[38] ), .ZN(new_n617_));
  NAND2_X1   g0232(.A1(\priority[36] ), .A2(\req[36] ), .ZN(new_n618_));
  NOR4_X1    g0233(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .A4(new_n618_), .ZN(new_n619_));
  NOR2_X1    g0234(.A1(\req[38] ), .A2(\req[39] ), .ZN(new_n620_));
  NAND2_X1   g0235(.A1(\priority[38] ), .A2(\req[37] ), .ZN(new_n621_));
  NOR2_X1    g0236(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1    g0237(.A1(\priority[40] ), .A2(\priority[41] ), .ZN(new_n623_));
  NAND2_X1   g0238(.A1(\priority[39] ), .A2(\req[39] ), .ZN(new_n624_));
  NOR2_X1    g0239(.A1(\req[41] ), .A2(\req[42] ), .ZN(new_n625_));
  NAND2_X1   g0240(.A1(\priority[41] ), .A2(\req[40] ), .ZN(new_n626_));
  NOR4_X1    g0241(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .A4(new_n626_), .ZN(new_n627_));
  OAI22_X1   g0242(.A1(new_n614_), .A2(new_n619_), .B1(new_n627_), .B2(new_n622_), .ZN(new_n628_));
  NOR4_X1    g0243(.A1(new_n577_), .A2(new_n594_), .A3(new_n611_), .A4(new_n628_), .ZN(new_n629_));
  NAND4_X1   g0244(.A1(new_n455_), .A2(new_n629_), .A3(new_n516_), .A4(new_n560_), .ZN(new_n630_));
  NAND2_X1   g0245(.A1(\priority[0] ), .A2(\req[127] ), .ZN(new_n631_));
  AOI21_X1   g0246(.A1(new_n630_), .A2(new_n386_), .B(new_n631_), .ZN(\grant[0] ));
  NOR2_X1    g0247(.A1(\priority[80] ), .A2(\priority[81] ), .ZN(new_n633_));
  NAND2_X1   g0248(.A1(\priority[79] ), .A2(\req[79] ), .ZN(new_n634_));
  NOR2_X1    g0249(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1    g0250(.A1(\req[81] ), .A2(\req[82] ), .ZN(new_n636_));
  NAND2_X1   g0251(.A1(\priority[81] ), .A2(\req[80] ), .ZN(new_n637_));
  NOR2_X1    g0252(.A1(\priority[83] ), .A2(\priority[84] ), .ZN(new_n638_));
  NAND2_X1   g0253(.A1(\priority[82] ), .A2(\req[82] ), .ZN(new_n639_));
  NOR4_X1    g0254(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .A4(new_n639_), .ZN(new_n640_));
  NOR2_X1    g0255(.A1(\req[84] ), .A2(\req[85] ), .ZN(new_n641_));
  NAND2_X1   g0256(.A1(\priority[84] ), .A2(\req[83] ), .ZN(new_n642_));
  NOR2_X1    g0257(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1    g0258(.A1(\priority[86] ), .A2(\priority[87] ), .ZN(new_n644_));
  NAND2_X1   g0259(.A1(\priority[85] ), .A2(\req[85] ), .ZN(new_n645_));
  NOR2_X1    g0260(.A1(\req[87] ), .A2(\req[88] ), .ZN(new_n646_));
  NAND2_X1   g0261(.A1(\priority[87] ), .A2(\req[86] ), .ZN(new_n647_));
  NOR4_X1    g0262(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .A4(new_n647_), .ZN(new_n648_));
  OAI22_X1   g0263(.A1(new_n635_), .A2(new_n640_), .B1(new_n648_), .B2(new_n643_), .ZN(new_n649_));
  NOR2_X1    g0264(.A1(\priority[89] ), .A2(\priority[90] ), .ZN(new_n650_));
  NAND2_X1   g0265(.A1(\priority[88] ), .A2(\req[88] ), .ZN(new_n651_));
  NOR2_X1    g0266(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1    g0267(.A1(\req[90] ), .A2(\req[91] ), .ZN(new_n653_));
  NAND2_X1   g0268(.A1(\priority[90] ), .A2(\req[89] ), .ZN(new_n654_));
  NOR2_X1    g0269(.A1(\priority[92] ), .A2(\priority[93] ), .ZN(new_n655_));
  NAND2_X1   g0270(.A1(\priority[91] ), .A2(\req[91] ), .ZN(new_n656_));
  NOR4_X1    g0271(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .A4(new_n656_), .ZN(new_n657_));
  NOR2_X1    g0272(.A1(\req[93] ), .A2(\req[94] ), .ZN(new_n658_));
  NAND2_X1   g0273(.A1(\priority[93] ), .A2(\req[92] ), .ZN(new_n659_));
  NOR2_X1    g0274(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1    g0275(.A1(\priority[95] ), .A2(\priority[96] ), .ZN(new_n661_));
  NAND2_X1   g0276(.A1(\priority[94] ), .A2(\req[94] ), .ZN(new_n662_));
  NOR2_X1    g0277(.A1(\req[96] ), .A2(\req[97] ), .ZN(new_n663_));
  NAND2_X1   g0278(.A1(\priority[96] ), .A2(\req[95] ), .ZN(new_n664_));
  NOR4_X1    g0279(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .A4(new_n664_), .ZN(new_n665_));
  OAI22_X1   g0280(.A1(new_n652_), .A2(new_n657_), .B1(new_n665_), .B2(new_n660_), .ZN(new_n666_));
  NOR2_X1    g0281(.A1(\priority[62] ), .A2(\priority[63] ), .ZN(new_n667_));
  NAND2_X1   g0282(.A1(\priority[61] ), .A2(\req[61] ), .ZN(new_n668_));
  NOR2_X1    g0283(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1    g0284(.A1(\req[63] ), .A2(\req[64] ), .ZN(new_n670_));
  NAND2_X1   g0285(.A1(\priority[63] ), .A2(\req[62] ), .ZN(new_n671_));
  NOR2_X1    g0286(.A1(\priority[65] ), .A2(\priority[66] ), .ZN(new_n672_));
  NAND2_X1   g0287(.A1(\priority[64] ), .A2(\req[64] ), .ZN(new_n673_));
  NOR4_X1    g0288(.A1(new_n670_), .A2(new_n671_), .A3(new_n672_), .A4(new_n673_), .ZN(new_n674_));
  NOR2_X1    g0289(.A1(\req[66] ), .A2(\req[67] ), .ZN(new_n675_));
  NAND2_X1   g0290(.A1(\priority[66] ), .A2(\req[65] ), .ZN(new_n676_));
  NOR2_X1    g0291(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1    g0292(.A1(\priority[68] ), .A2(\priority[69] ), .ZN(new_n678_));
  NAND2_X1   g0293(.A1(\priority[67] ), .A2(\req[67] ), .ZN(new_n679_));
  NOR2_X1    g0294(.A1(\req[69] ), .A2(\req[70] ), .ZN(new_n680_));
  NAND2_X1   g0295(.A1(\priority[69] ), .A2(\req[68] ), .ZN(new_n681_));
  NOR4_X1    g0296(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .A4(new_n681_), .ZN(new_n682_));
  OAI22_X1   g0297(.A1(new_n669_), .A2(new_n674_), .B1(new_n682_), .B2(new_n677_), .ZN(new_n683_));
  NOR2_X1    g0298(.A1(\priority[71] ), .A2(\priority[72] ), .ZN(new_n684_));
  NAND2_X1   g0299(.A1(\priority[70] ), .A2(\req[70] ), .ZN(new_n685_));
  NOR2_X1    g0300(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NOR2_X1    g0301(.A1(\req[72] ), .A2(\req[73] ), .ZN(new_n687_));
  NAND2_X1   g0302(.A1(\priority[72] ), .A2(\req[71] ), .ZN(new_n688_));
  NOR2_X1    g0303(.A1(\priority[74] ), .A2(\priority[75] ), .ZN(new_n689_));
  NAND2_X1   g0304(.A1(\priority[73] ), .A2(\req[73] ), .ZN(new_n690_));
  NOR4_X1    g0305(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .A4(new_n690_), .ZN(new_n691_));
  NOR2_X1    g0306(.A1(\req[75] ), .A2(\req[76] ), .ZN(new_n692_));
  NAND2_X1   g0307(.A1(\priority[75] ), .A2(\req[74] ), .ZN(new_n693_));
  NOR2_X1    g0308(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1    g0309(.A1(\priority[77] ), .A2(\priority[78] ), .ZN(new_n695_));
  NAND2_X1   g0310(.A1(\priority[76] ), .A2(\req[76] ), .ZN(new_n696_));
  NOR2_X1    g0311(.A1(\req[78] ), .A2(\req[79] ), .ZN(new_n697_));
  NAND2_X1   g0312(.A1(\priority[78] ), .A2(\req[77] ), .ZN(new_n698_));
  NOR4_X1    g0313(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .A4(new_n698_), .ZN(new_n699_));
  OAI22_X1   g0314(.A1(new_n686_), .A2(new_n691_), .B1(new_n699_), .B2(new_n694_), .ZN(new_n700_));
  NOR4_X1    g0315(.A1(new_n649_), .A2(new_n666_), .A3(new_n683_), .A4(new_n700_), .ZN(new_n701_));
  NOR2_X1    g0316(.A1(\priority[125] ), .A2(\priority[126] ), .ZN(new_n702_));
  NAND2_X1   g0317(.A1(\priority[124] ), .A2(\req[124] ), .ZN(new_n703_));
  NOR2_X1    g0318(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NOR2_X1    g0319(.A1(\req[126] ), .A2(\req[127] ), .ZN(new_n705_));
  NAND2_X1   g0320(.A1(\priority[126] ), .A2(\req[125] ), .ZN(new_n706_));
  NOR2_X1    g0321(.A1(\priority[0] ), .A2(\priority[1] ), .ZN(new_n707_));
  NAND2_X1   g0322(.A1(\priority[127] ), .A2(\req[127] ), .ZN(new_n708_));
  NOR4_X1    g0323(.A1(new_n705_), .A2(new_n706_), .A3(new_n707_), .A4(new_n708_), .ZN(new_n709_));
  NOR2_X1    g0324(.A1(new_n709_), .A2(new_n704_), .ZN(new_n710_));
  NOR2_X1    g0325(.A1(\priority[116] ), .A2(\priority[117] ), .ZN(new_n711_));
  NAND2_X1   g0326(.A1(\priority[115] ), .A2(\req[115] ), .ZN(new_n712_));
  NOR2_X1    g0327(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NOR2_X1    g0328(.A1(\req[117] ), .A2(\req[118] ), .ZN(new_n714_));
  NAND2_X1   g0329(.A1(\priority[117] ), .A2(\req[116] ), .ZN(new_n715_));
  NOR2_X1    g0330(.A1(\priority[119] ), .A2(\priority[120] ), .ZN(new_n716_));
  NAND2_X1   g0331(.A1(\priority[118] ), .A2(\req[118] ), .ZN(new_n717_));
  NOR4_X1    g0332(.A1(new_n714_), .A2(new_n715_), .A3(new_n716_), .A4(new_n717_), .ZN(new_n718_));
  NOR2_X1    g0333(.A1(\req[120] ), .A2(\req[121] ), .ZN(new_n719_));
  NAND2_X1   g0334(.A1(\priority[120] ), .A2(\req[119] ), .ZN(new_n720_));
  NOR2_X1    g0335(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1    g0336(.A1(\priority[122] ), .A2(\priority[123] ), .ZN(new_n722_));
  NAND2_X1   g0337(.A1(\priority[121] ), .A2(\req[121] ), .ZN(new_n723_));
  NOR2_X1    g0338(.A1(\req[123] ), .A2(\req[124] ), .ZN(new_n724_));
  NAND2_X1   g0339(.A1(\priority[123] ), .A2(\req[122] ), .ZN(new_n725_));
  NOR4_X1    g0340(.A1(new_n722_), .A2(new_n723_), .A3(new_n724_), .A4(new_n725_), .ZN(new_n726_));
  OAI22_X1   g0341(.A1(new_n713_), .A2(new_n718_), .B1(new_n726_), .B2(new_n721_), .ZN(new_n727_));
  NOR2_X1    g0342(.A1(\priority[98] ), .A2(\priority[99] ), .ZN(new_n728_));
  NAND2_X1   g0343(.A1(\priority[97] ), .A2(\req[97] ), .ZN(new_n729_));
  NOR2_X1    g0344(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NOR2_X1    g0345(.A1(\req[99] ), .A2(\req[100] ), .ZN(new_n731_));
  NAND2_X1   g0346(.A1(\priority[99] ), .A2(\req[98] ), .ZN(new_n732_));
  NOR2_X1    g0347(.A1(\priority[101] ), .A2(\priority[102] ), .ZN(new_n733_));
  NAND2_X1   g0348(.A1(\priority[100] ), .A2(\req[100] ), .ZN(new_n734_));
  NOR4_X1    g0349(.A1(new_n731_), .A2(new_n732_), .A3(new_n733_), .A4(new_n734_), .ZN(new_n735_));
  NOR2_X1    g0350(.A1(\req[102] ), .A2(\req[103] ), .ZN(new_n736_));
  NAND2_X1   g0351(.A1(\priority[102] ), .A2(\req[101] ), .ZN(new_n737_));
  NOR2_X1    g0352(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NOR2_X1    g0353(.A1(\priority[104] ), .A2(\priority[105] ), .ZN(new_n739_));
  NAND2_X1   g0354(.A1(\priority[103] ), .A2(\req[103] ), .ZN(new_n740_));
  NOR2_X1    g0355(.A1(\req[105] ), .A2(\req[106] ), .ZN(new_n741_));
  NAND2_X1   g0356(.A1(\priority[105] ), .A2(\req[104] ), .ZN(new_n742_));
  NOR4_X1    g0357(.A1(new_n739_), .A2(new_n740_), .A3(new_n741_), .A4(new_n742_), .ZN(new_n743_));
  OAI22_X1   g0358(.A1(new_n730_), .A2(new_n735_), .B1(new_n743_), .B2(new_n738_), .ZN(new_n744_));
  NOR2_X1    g0359(.A1(\priority[107] ), .A2(\priority[108] ), .ZN(new_n745_));
  NAND2_X1   g0360(.A1(\priority[106] ), .A2(\req[106] ), .ZN(new_n746_));
  NOR2_X1    g0361(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1    g0362(.A1(\req[108] ), .A2(\req[109] ), .ZN(new_n748_));
  NAND2_X1   g0363(.A1(\priority[108] ), .A2(\req[107] ), .ZN(new_n749_));
  NOR2_X1    g0364(.A1(\priority[110] ), .A2(\priority[111] ), .ZN(new_n750_));
  NAND2_X1   g0365(.A1(\priority[109] ), .A2(\req[109] ), .ZN(new_n751_));
  NOR4_X1    g0366(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .A4(new_n751_), .ZN(new_n752_));
  NOR2_X1    g0367(.A1(\req[111] ), .A2(\req[112] ), .ZN(new_n753_));
  NAND2_X1   g0368(.A1(\priority[111] ), .A2(\req[110] ), .ZN(new_n754_));
  NOR2_X1    g0369(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NOR2_X1    g0370(.A1(\priority[113] ), .A2(\priority[114] ), .ZN(new_n756_));
  NAND2_X1   g0371(.A1(\priority[112] ), .A2(\req[112] ), .ZN(new_n757_));
  NOR2_X1    g0372(.A1(\req[114] ), .A2(\req[115] ), .ZN(new_n758_));
  NAND2_X1   g0373(.A1(\priority[114] ), .A2(\req[113] ), .ZN(new_n759_));
  NOR4_X1    g0374(.A1(new_n756_), .A2(new_n757_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n760_));
  OAI22_X1   g0375(.A1(new_n747_), .A2(new_n752_), .B1(new_n760_), .B2(new_n755_), .ZN(new_n761_));
  NOR4_X1    g0376(.A1(new_n727_), .A2(new_n744_), .A3(new_n761_), .A4(new_n710_), .ZN(new_n762_));
  NOR2_X1    g0377(.A1(\req[3] ), .A2(\req[4] ), .ZN(new_n763_));
  NOR2_X1    g0378(.A1(\priority[5] ), .A2(\priority[6] ), .ZN(new_n764_));
  NAND2_X1   g0379(.A1(\priority[4] ), .A2(\req[4] ), .ZN(new_n765_));
  NOR2_X1    g0380(.A1(\req[6] ), .A2(\req[7] ), .ZN(new_n766_));
  NAND2_X1   g0381(.A1(\priority[6] ), .A2(\req[5] ), .ZN(new_n767_));
  NOR4_X1    g0382(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .A4(new_n767_), .ZN(new_n768_));
  INV_X1     g0383(.I(\req[2] ), .ZN(new_n769_));
  AOI21_X1   g0384(.A1(new_n769_), .A2(\priority[2] ), .B(\priority[3] ), .ZN(new_n770_));
  OAI21_X1   g0385(.A1(new_n768_), .A2(new_n763_), .B(new_n770_), .ZN(new_n771_));
  NOR2_X1    g0386(.A1(\priority[8] ), .A2(\priority[9] ), .ZN(new_n772_));
  NAND2_X1   g0387(.A1(\priority[7] ), .A2(\req[7] ), .ZN(new_n773_));
  NOR2_X1    g0388(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NOR2_X1    g0389(.A1(\req[9] ), .A2(\req[10] ), .ZN(new_n775_));
  NAND2_X1   g0390(.A1(\priority[9] ), .A2(\req[8] ), .ZN(new_n776_));
  NOR2_X1    g0391(.A1(\priority[11] ), .A2(\priority[12] ), .ZN(new_n777_));
  NAND2_X1   g0392(.A1(\priority[10] ), .A2(\req[10] ), .ZN(new_n778_));
  NOR4_X1    g0393(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .A4(new_n778_), .ZN(new_n779_));
  NOR2_X1    g0394(.A1(\req[12] ), .A2(\req[13] ), .ZN(new_n780_));
  NAND2_X1   g0395(.A1(\priority[12] ), .A2(\req[11] ), .ZN(new_n781_));
  NOR2_X1    g0396(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NOR2_X1    g0397(.A1(\priority[14] ), .A2(\priority[15] ), .ZN(new_n783_));
  NAND2_X1   g0398(.A1(\priority[13] ), .A2(\req[13] ), .ZN(new_n784_));
  NOR2_X1    g0399(.A1(\req[15] ), .A2(\req[16] ), .ZN(new_n785_));
  NAND2_X1   g0400(.A1(\priority[15] ), .A2(\req[14] ), .ZN(new_n786_));
  NOR4_X1    g0401(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .A4(new_n786_), .ZN(new_n787_));
  OAI22_X1   g0402(.A1(new_n774_), .A2(new_n779_), .B1(new_n787_), .B2(new_n782_), .ZN(new_n788_));
  NOR2_X1    g0403(.A1(\priority[17] ), .A2(\priority[18] ), .ZN(new_n789_));
  NAND2_X1   g0404(.A1(\priority[16] ), .A2(\req[16] ), .ZN(new_n790_));
  NOR2_X1    g0405(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1    g0406(.A1(\req[18] ), .A2(\req[19] ), .ZN(new_n792_));
  NAND2_X1   g0407(.A1(\priority[18] ), .A2(\req[17] ), .ZN(new_n793_));
  NOR2_X1    g0408(.A1(\priority[20] ), .A2(\priority[21] ), .ZN(new_n794_));
  NAND2_X1   g0409(.A1(\priority[19] ), .A2(\req[19] ), .ZN(new_n795_));
  NOR4_X1    g0410(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .A4(new_n795_), .ZN(new_n796_));
  NOR2_X1    g0411(.A1(\req[21] ), .A2(\req[22] ), .ZN(new_n797_));
  NAND2_X1   g0412(.A1(\priority[21] ), .A2(\req[20] ), .ZN(new_n798_));
  NOR2_X1    g0413(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NOR2_X1    g0414(.A1(\priority[23] ), .A2(\priority[24] ), .ZN(new_n800_));
  NAND2_X1   g0415(.A1(\priority[22] ), .A2(\req[22] ), .ZN(new_n801_));
  NOR2_X1    g0416(.A1(\req[24] ), .A2(\req[25] ), .ZN(new_n802_));
  NAND2_X1   g0417(.A1(\priority[24] ), .A2(\req[23] ), .ZN(new_n803_));
  NOR4_X1    g0418(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .A4(new_n803_), .ZN(new_n804_));
  OAI22_X1   g0419(.A1(new_n791_), .A2(new_n796_), .B1(new_n804_), .B2(new_n799_), .ZN(new_n805_));
  NOR3_X1    g0420(.A1(new_n788_), .A2(new_n805_), .A3(new_n771_), .ZN(new_n806_));
  NOR2_X1    g0421(.A1(\priority[44] ), .A2(\priority[45] ), .ZN(new_n807_));
  NAND2_X1   g0422(.A1(\priority[43] ), .A2(\req[43] ), .ZN(new_n808_));
  NOR2_X1    g0423(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1    g0424(.A1(\req[45] ), .A2(\req[46] ), .ZN(new_n810_));
  NAND2_X1   g0425(.A1(\priority[45] ), .A2(\req[44] ), .ZN(new_n811_));
  NOR2_X1    g0426(.A1(\priority[47] ), .A2(\priority[48] ), .ZN(new_n812_));
  NAND2_X1   g0427(.A1(\priority[46] ), .A2(\req[46] ), .ZN(new_n813_));
  NOR4_X1    g0428(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .A4(new_n813_), .ZN(new_n814_));
  NOR2_X1    g0429(.A1(\req[48] ), .A2(\req[49] ), .ZN(new_n815_));
  NAND2_X1   g0430(.A1(\priority[48] ), .A2(\req[47] ), .ZN(new_n816_));
  NOR2_X1    g0431(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1    g0432(.A1(\priority[50] ), .A2(\priority[51] ), .ZN(new_n818_));
  NAND2_X1   g0433(.A1(\priority[49] ), .A2(\req[49] ), .ZN(new_n819_));
  NOR2_X1    g0434(.A1(\req[51] ), .A2(\req[52] ), .ZN(new_n820_));
  NAND2_X1   g0435(.A1(\priority[51] ), .A2(\req[50] ), .ZN(new_n821_));
  NOR4_X1    g0436(.A1(new_n818_), .A2(new_n819_), .A3(new_n820_), .A4(new_n821_), .ZN(new_n822_));
  OAI22_X1   g0437(.A1(new_n809_), .A2(new_n814_), .B1(new_n822_), .B2(new_n817_), .ZN(new_n823_));
  NOR2_X1    g0438(.A1(\priority[53] ), .A2(\priority[54] ), .ZN(new_n824_));
  NAND2_X1   g0439(.A1(\priority[52] ), .A2(\req[52] ), .ZN(new_n825_));
  NOR2_X1    g0440(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NOR2_X1    g0441(.A1(\req[54] ), .A2(\req[55] ), .ZN(new_n827_));
  NAND2_X1   g0442(.A1(\priority[54] ), .A2(\req[53] ), .ZN(new_n828_));
  NOR2_X1    g0443(.A1(\priority[56] ), .A2(\priority[57] ), .ZN(new_n829_));
  NAND2_X1   g0444(.A1(\priority[55] ), .A2(\req[55] ), .ZN(new_n830_));
  NOR4_X1    g0445(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .A4(new_n830_), .ZN(new_n831_));
  NOR2_X1    g0446(.A1(\req[57] ), .A2(\req[58] ), .ZN(new_n832_));
  NAND2_X1   g0447(.A1(\priority[57] ), .A2(\req[56] ), .ZN(new_n833_));
  NOR2_X1    g0448(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1    g0449(.A1(\priority[59] ), .A2(\priority[60] ), .ZN(new_n835_));
  NAND2_X1   g0450(.A1(\priority[58] ), .A2(\req[58] ), .ZN(new_n836_));
  NOR2_X1    g0451(.A1(\req[60] ), .A2(\req[61] ), .ZN(new_n837_));
  NAND2_X1   g0452(.A1(\priority[60] ), .A2(\req[59] ), .ZN(new_n838_));
  NOR4_X1    g0453(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .A4(new_n838_), .ZN(new_n839_));
  OAI22_X1   g0454(.A1(new_n826_), .A2(new_n831_), .B1(new_n839_), .B2(new_n834_), .ZN(new_n840_));
  NOR2_X1    g0455(.A1(\priority[26] ), .A2(\priority[27] ), .ZN(new_n841_));
  NAND2_X1   g0456(.A1(\priority[25] ), .A2(\req[25] ), .ZN(new_n842_));
  NOR2_X1    g0457(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1    g0458(.A1(\req[27] ), .A2(\req[28] ), .ZN(new_n844_));
  NAND2_X1   g0459(.A1(\priority[27] ), .A2(\req[26] ), .ZN(new_n845_));
  NOR2_X1    g0460(.A1(\priority[29] ), .A2(\priority[30] ), .ZN(new_n846_));
  NAND2_X1   g0461(.A1(\priority[28] ), .A2(\req[28] ), .ZN(new_n847_));
  NOR4_X1    g0462(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .A4(new_n847_), .ZN(new_n848_));
  NOR2_X1    g0463(.A1(\req[30] ), .A2(\req[31] ), .ZN(new_n849_));
  NAND2_X1   g0464(.A1(\priority[30] ), .A2(\req[29] ), .ZN(new_n850_));
  NOR2_X1    g0465(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1    g0466(.A1(\priority[32] ), .A2(\priority[33] ), .ZN(new_n852_));
  NAND2_X1   g0467(.A1(\priority[31] ), .A2(\req[31] ), .ZN(new_n853_));
  NOR2_X1    g0468(.A1(\req[33] ), .A2(\req[34] ), .ZN(new_n854_));
  NAND2_X1   g0469(.A1(\priority[33] ), .A2(\req[32] ), .ZN(new_n855_));
  NOR4_X1    g0470(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .A4(new_n855_), .ZN(new_n856_));
  OAI22_X1   g0471(.A1(new_n843_), .A2(new_n848_), .B1(new_n856_), .B2(new_n851_), .ZN(new_n857_));
  NOR2_X1    g0472(.A1(\priority[35] ), .A2(\priority[36] ), .ZN(new_n858_));
  NAND2_X1   g0473(.A1(\priority[34] ), .A2(\req[34] ), .ZN(new_n859_));
  NOR2_X1    g0474(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1    g0475(.A1(\req[36] ), .A2(\req[37] ), .ZN(new_n861_));
  NAND2_X1   g0476(.A1(\priority[36] ), .A2(\req[35] ), .ZN(new_n862_));
  NOR2_X1    g0477(.A1(\priority[38] ), .A2(\priority[39] ), .ZN(new_n863_));
  NAND2_X1   g0478(.A1(\priority[37] ), .A2(\req[37] ), .ZN(new_n864_));
  NOR4_X1    g0479(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .A4(new_n864_), .ZN(new_n865_));
  NOR2_X1    g0480(.A1(\req[39] ), .A2(\req[40] ), .ZN(new_n866_));
  NAND2_X1   g0481(.A1(\priority[39] ), .A2(\req[38] ), .ZN(new_n867_));
  NOR2_X1    g0482(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1    g0483(.A1(\priority[41] ), .A2(\priority[42] ), .ZN(new_n869_));
  NAND2_X1   g0484(.A1(\priority[40] ), .A2(\req[40] ), .ZN(new_n870_));
  NOR2_X1    g0485(.A1(\req[42] ), .A2(\req[43] ), .ZN(new_n871_));
  NAND2_X1   g0486(.A1(\priority[42] ), .A2(\req[41] ), .ZN(new_n872_));
  NOR4_X1    g0487(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .A4(new_n872_), .ZN(new_n873_));
  OAI22_X1   g0488(.A1(new_n860_), .A2(new_n865_), .B1(new_n873_), .B2(new_n868_), .ZN(new_n874_));
  NOR4_X1    g0489(.A1(new_n823_), .A2(new_n840_), .A3(new_n857_), .A4(new_n874_), .ZN(new_n875_));
  NAND4_X1   g0490(.A1(new_n701_), .A2(new_n875_), .A3(new_n762_), .A4(new_n806_), .ZN(new_n876_));
  NAND2_X1   g0491(.A1(\priority[1] ), .A2(\req[0] ), .ZN(new_n877_));
  AOI21_X1   g0492(.A1(new_n876_), .A2(new_n523_), .B(new_n877_), .ZN(\grant[1] ));
  NOR2_X1    g0493(.A1(\priority[81] ), .A2(\priority[82] ), .ZN(new_n879_));
  NAND2_X1   g0494(.A1(\priority[80] ), .A2(\req[80] ), .ZN(new_n880_));
  NOR2_X1    g0495(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NOR2_X1    g0496(.A1(\req[82] ), .A2(\req[83] ), .ZN(new_n882_));
  NAND2_X1   g0497(.A1(\priority[82] ), .A2(\req[81] ), .ZN(new_n883_));
  NOR2_X1    g0498(.A1(\priority[84] ), .A2(\priority[85] ), .ZN(new_n884_));
  NAND2_X1   g0499(.A1(\priority[83] ), .A2(\req[83] ), .ZN(new_n885_));
  NOR4_X1    g0500(.A1(new_n882_), .A2(new_n883_), .A3(new_n884_), .A4(new_n885_), .ZN(new_n886_));
  NOR2_X1    g0501(.A1(\req[85] ), .A2(\req[86] ), .ZN(new_n887_));
  NAND2_X1   g0502(.A1(\priority[85] ), .A2(\req[84] ), .ZN(new_n888_));
  NOR2_X1    g0503(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NOR2_X1    g0504(.A1(\priority[87] ), .A2(\priority[88] ), .ZN(new_n890_));
  NAND2_X1   g0505(.A1(\priority[86] ), .A2(\req[86] ), .ZN(new_n891_));
  NOR2_X1    g0506(.A1(\req[88] ), .A2(\req[89] ), .ZN(new_n892_));
  NAND2_X1   g0507(.A1(\priority[88] ), .A2(\req[87] ), .ZN(new_n893_));
  NOR4_X1    g0508(.A1(new_n890_), .A2(new_n891_), .A3(new_n892_), .A4(new_n893_), .ZN(new_n894_));
  OAI22_X1   g0509(.A1(new_n881_), .A2(new_n886_), .B1(new_n894_), .B2(new_n889_), .ZN(new_n895_));
  NOR2_X1    g0510(.A1(\priority[90] ), .A2(\priority[91] ), .ZN(new_n896_));
  NAND2_X1   g0511(.A1(\priority[89] ), .A2(\req[89] ), .ZN(new_n897_));
  NOR2_X1    g0512(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1    g0513(.A1(\req[91] ), .A2(\req[92] ), .ZN(new_n899_));
  NAND2_X1   g0514(.A1(\priority[91] ), .A2(\req[90] ), .ZN(new_n900_));
  NOR2_X1    g0515(.A1(\priority[93] ), .A2(\priority[94] ), .ZN(new_n901_));
  NAND2_X1   g0516(.A1(\priority[92] ), .A2(\req[92] ), .ZN(new_n902_));
  NOR4_X1    g0517(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .A4(new_n902_), .ZN(new_n903_));
  NOR2_X1    g0518(.A1(\req[94] ), .A2(\req[95] ), .ZN(new_n904_));
  NAND2_X1   g0519(.A1(\priority[94] ), .A2(\req[93] ), .ZN(new_n905_));
  NOR2_X1    g0520(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1    g0521(.A1(\priority[96] ), .A2(\priority[97] ), .ZN(new_n907_));
  NAND2_X1   g0522(.A1(\priority[95] ), .A2(\req[95] ), .ZN(new_n908_));
  NOR2_X1    g0523(.A1(\req[97] ), .A2(\req[98] ), .ZN(new_n909_));
  NAND2_X1   g0524(.A1(\priority[97] ), .A2(\req[96] ), .ZN(new_n910_));
  NOR4_X1    g0525(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .A4(new_n910_), .ZN(new_n911_));
  OAI22_X1   g0526(.A1(new_n898_), .A2(new_n903_), .B1(new_n911_), .B2(new_n906_), .ZN(new_n912_));
  NOR2_X1    g0527(.A1(\priority[63] ), .A2(\priority[64] ), .ZN(new_n913_));
  NAND2_X1   g0528(.A1(\priority[62] ), .A2(\req[62] ), .ZN(new_n914_));
  NOR2_X1    g0529(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1    g0530(.A1(\req[64] ), .A2(\req[65] ), .ZN(new_n916_));
  NAND2_X1   g0531(.A1(\priority[64] ), .A2(\req[63] ), .ZN(new_n917_));
  NOR2_X1    g0532(.A1(\priority[66] ), .A2(\priority[67] ), .ZN(new_n918_));
  NAND2_X1   g0533(.A1(\priority[65] ), .A2(\req[65] ), .ZN(new_n919_));
  NOR4_X1    g0534(.A1(new_n916_), .A2(new_n917_), .A3(new_n918_), .A4(new_n919_), .ZN(new_n920_));
  NOR2_X1    g0535(.A1(\req[67] ), .A2(\req[68] ), .ZN(new_n921_));
  NAND2_X1   g0536(.A1(\priority[67] ), .A2(\req[66] ), .ZN(new_n922_));
  NOR2_X1    g0537(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1    g0538(.A1(\priority[69] ), .A2(\priority[70] ), .ZN(new_n924_));
  NAND2_X1   g0539(.A1(\priority[68] ), .A2(\req[68] ), .ZN(new_n925_));
  NOR2_X1    g0540(.A1(\req[70] ), .A2(\req[71] ), .ZN(new_n926_));
  NAND2_X1   g0541(.A1(\priority[70] ), .A2(\req[69] ), .ZN(new_n927_));
  NOR4_X1    g0542(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .A4(new_n927_), .ZN(new_n928_));
  OAI22_X1   g0543(.A1(new_n915_), .A2(new_n920_), .B1(new_n928_), .B2(new_n923_), .ZN(new_n929_));
  NOR2_X1    g0544(.A1(\priority[72] ), .A2(\priority[73] ), .ZN(new_n930_));
  NAND2_X1   g0545(.A1(\priority[71] ), .A2(\req[71] ), .ZN(new_n931_));
  NOR2_X1    g0546(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1    g0547(.A1(\req[73] ), .A2(\req[74] ), .ZN(new_n933_));
  NAND2_X1   g0548(.A1(\priority[73] ), .A2(\req[72] ), .ZN(new_n934_));
  NOR2_X1    g0549(.A1(\priority[75] ), .A2(\priority[76] ), .ZN(new_n935_));
  NAND2_X1   g0550(.A1(\priority[74] ), .A2(\req[74] ), .ZN(new_n936_));
  NOR4_X1    g0551(.A1(new_n933_), .A2(new_n934_), .A3(new_n935_), .A4(new_n936_), .ZN(new_n937_));
  NOR2_X1    g0552(.A1(\req[76] ), .A2(\req[77] ), .ZN(new_n938_));
  NAND2_X1   g0553(.A1(\priority[76] ), .A2(\req[75] ), .ZN(new_n939_));
  NOR2_X1    g0554(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1    g0555(.A1(\priority[78] ), .A2(\priority[79] ), .ZN(new_n941_));
  NAND2_X1   g0556(.A1(\priority[77] ), .A2(\req[77] ), .ZN(new_n942_));
  NOR2_X1    g0557(.A1(\req[79] ), .A2(\req[80] ), .ZN(new_n943_));
  NAND2_X1   g0558(.A1(\priority[79] ), .A2(\req[78] ), .ZN(new_n944_));
  NOR4_X1    g0559(.A1(new_n941_), .A2(new_n942_), .A3(new_n943_), .A4(new_n944_), .ZN(new_n945_));
  OAI22_X1   g0560(.A1(new_n932_), .A2(new_n937_), .B1(new_n945_), .B2(new_n940_), .ZN(new_n946_));
  NOR4_X1    g0561(.A1(new_n895_), .A2(new_n912_), .A3(new_n929_), .A4(new_n946_), .ZN(new_n947_));
  NOR2_X1    g0562(.A1(\priority[126] ), .A2(\priority[127] ), .ZN(new_n948_));
  NAND2_X1   g0563(.A1(\priority[125] ), .A2(\req[125] ), .ZN(new_n949_));
  NOR2_X1    g0564(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  NOR2_X1    g0565(.A1(\req[0] ), .A2(\req[127] ), .ZN(new_n951_));
  NAND2_X1   g0566(.A1(\priority[127] ), .A2(\req[126] ), .ZN(new_n952_));
  NOR2_X1    g0567(.A1(\priority[1] ), .A2(\priority[2] ), .ZN(new_n953_));
  NAND2_X1   g0568(.A1(\priority[0] ), .A2(\req[0] ), .ZN(new_n954_));
  NOR4_X1    g0569(.A1(new_n951_), .A2(new_n952_), .A3(new_n953_), .A4(new_n954_), .ZN(new_n955_));
  NOR2_X1    g0570(.A1(new_n955_), .A2(new_n950_), .ZN(new_n956_));
  NOR2_X1    g0571(.A1(\priority[117] ), .A2(\priority[118] ), .ZN(new_n957_));
  NAND2_X1   g0572(.A1(\priority[116] ), .A2(\req[116] ), .ZN(new_n958_));
  NOR2_X1    g0573(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  NOR2_X1    g0574(.A1(\req[118] ), .A2(\req[119] ), .ZN(new_n960_));
  NAND2_X1   g0575(.A1(\priority[118] ), .A2(\req[117] ), .ZN(new_n961_));
  NOR2_X1    g0576(.A1(\priority[120] ), .A2(\priority[121] ), .ZN(new_n962_));
  NAND2_X1   g0577(.A1(\priority[119] ), .A2(\req[119] ), .ZN(new_n963_));
  NOR4_X1    g0578(.A1(new_n960_), .A2(new_n961_), .A3(new_n962_), .A4(new_n963_), .ZN(new_n964_));
  NOR2_X1    g0579(.A1(\req[121] ), .A2(\req[122] ), .ZN(new_n965_));
  NAND2_X1   g0580(.A1(\priority[121] ), .A2(\req[120] ), .ZN(new_n966_));
  NOR2_X1    g0581(.A1(new_n965_), .A2(new_n966_), .ZN(new_n967_));
  NOR2_X1    g0582(.A1(\priority[123] ), .A2(\priority[124] ), .ZN(new_n968_));
  NAND2_X1   g0583(.A1(\priority[122] ), .A2(\req[122] ), .ZN(new_n969_));
  NOR2_X1    g0584(.A1(\req[124] ), .A2(\req[125] ), .ZN(new_n970_));
  NAND2_X1   g0585(.A1(\priority[124] ), .A2(\req[123] ), .ZN(new_n971_));
  NOR4_X1    g0586(.A1(new_n968_), .A2(new_n969_), .A3(new_n970_), .A4(new_n971_), .ZN(new_n972_));
  OAI22_X1   g0587(.A1(new_n959_), .A2(new_n964_), .B1(new_n972_), .B2(new_n967_), .ZN(new_n973_));
  NOR2_X1    g0588(.A1(\priority[99] ), .A2(\priority[100] ), .ZN(new_n974_));
  NAND2_X1   g0589(.A1(\priority[98] ), .A2(\req[98] ), .ZN(new_n975_));
  NOR2_X1    g0590(.A1(new_n974_), .A2(new_n975_), .ZN(new_n976_));
  NOR2_X1    g0591(.A1(\req[100] ), .A2(\req[101] ), .ZN(new_n977_));
  NAND2_X1   g0592(.A1(\priority[100] ), .A2(\req[99] ), .ZN(new_n978_));
  NOR2_X1    g0593(.A1(\priority[102] ), .A2(\priority[103] ), .ZN(new_n979_));
  NAND2_X1   g0594(.A1(\priority[101] ), .A2(\req[101] ), .ZN(new_n980_));
  NOR4_X1    g0595(.A1(new_n977_), .A2(new_n978_), .A3(new_n979_), .A4(new_n980_), .ZN(new_n981_));
  NOR2_X1    g0596(.A1(\req[103] ), .A2(\req[104] ), .ZN(new_n982_));
  NAND2_X1   g0597(.A1(\priority[103] ), .A2(\req[102] ), .ZN(new_n983_));
  NOR2_X1    g0598(.A1(new_n982_), .A2(new_n983_), .ZN(new_n984_));
  NOR2_X1    g0599(.A1(\priority[105] ), .A2(\priority[106] ), .ZN(new_n985_));
  NAND2_X1   g0600(.A1(\priority[104] ), .A2(\req[104] ), .ZN(new_n986_));
  NOR2_X1    g0601(.A1(\req[106] ), .A2(\req[107] ), .ZN(new_n987_));
  NAND2_X1   g0602(.A1(\priority[106] ), .A2(\req[105] ), .ZN(new_n988_));
  NOR4_X1    g0603(.A1(new_n985_), .A2(new_n986_), .A3(new_n987_), .A4(new_n988_), .ZN(new_n989_));
  OAI22_X1   g0604(.A1(new_n976_), .A2(new_n981_), .B1(new_n989_), .B2(new_n984_), .ZN(new_n990_));
  NOR2_X1    g0605(.A1(\priority[108] ), .A2(\priority[109] ), .ZN(new_n991_));
  NAND2_X1   g0606(.A1(\priority[107] ), .A2(\req[107] ), .ZN(new_n992_));
  NOR2_X1    g0607(.A1(new_n991_), .A2(new_n992_), .ZN(new_n993_));
  NOR2_X1    g0608(.A1(\req[109] ), .A2(\req[110] ), .ZN(new_n994_));
  NAND2_X1   g0609(.A1(\priority[109] ), .A2(\req[108] ), .ZN(new_n995_));
  NOR2_X1    g0610(.A1(\priority[111] ), .A2(\priority[112] ), .ZN(new_n996_));
  NAND2_X1   g0611(.A1(\priority[110] ), .A2(\req[110] ), .ZN(new_n997_));
  NOR4_X1    g0612(.A1(new_n994_), .A2(new_n995_), .A3(new_n996_), .A4(new_n997_), .ZN(new_n998_));
  NOR2_X1    g0613(.A1(\req[112] ), .A2(\req[113] ), .ZN(new_n999_));
  NAND2_X1   g0614(.A1(\priority[112] ), .A2(\req[111] ), .ZN(new_n1000_));
  NOR2_X1    g0615(.A1(new_n999_), .A2(new_n1000_), .ZN(new_n1001_));
  NOR2_X1    g0616(.A1(\priority[114] ), .A2(\priority[115] ), .ZN(new_n1002_));
  NAND2_X1   g0617(.A1(\priority[113] ), .A2(\req[113] ), .ZN(new_n1003_));
  NOR2_X1    g0618(.A1(\req[115] ), .A2(\req[116] ), .ZN(new_n1004_));
  NAND2_X1   g0619(.A1(\priority[115] ), .A2(\req[114] ), .ZN(new_n1005_));
  NOR4_X1    g0620(.A1(new_n1002_), .A2(new_n1003_), .A3(new_n1004_), .A4(new_n1005_), .ZN(new_n1006_));
  OAI22_X1   g0621(.A1(new_n993_), .A2(new_n998_), .B1(new_n1006_), .B2(new_n1001_), .ZN(new_n1007_));
  NOR4_X1    g0622(.A1(new_n973_), .A2(new_n990_), .A3(new_n1007_), .A4(new_n956_), .ZN(new_n1008_));
  NOR2_X1    g0623(.A1(\req[4] ), .A2(\req[5] ), .ZN(new_n1009_));
  NOR2_X1    g0624(.A1(\priority[6] ), .A2(\priority[7] ), .ZN(new_n1010_));
  NAND2_X1   g0625(.A1(\priority[5] ), .A2(\req[5] ), .ZN(new_n1011_));
  NOR2_X1    g0626(.A1(\req[7] ), .A2(\req[8] ), .ZN(new_n1012_));
  NAND2_X1   g0627(.A1(\priority[7] ), .A2(\req[6] ), .ZN(new_n1013_));
  NOR4_X1    g0628(.A1(new_n1010_), .A2(new_n1011_), .A3(new_n1012_), .A4(new_n1013_), .ZN(new_n1014_));
  INV_X1     g0629(.I(\req[3] ), .ZN(new_n1015_));
  AOI21_X1   g0630(.A1(new_n1015_), .A2(\priority[3] ), .B(\priority[4] ), .ZN(new_n1016_));
  OAI21_X1   g0631(.A1(new_n1014_), .A2(new_n1009_), .B(new_n1016_), .ZN(new_n1017_));
  NOR2_X1    g0632(.A1(\priority[9] ), .A2(\priority[10] ), .ZN(new_n1018_));
  NAND2_X1   g0633(.A1(\priority[8] ), .A2(\req[8] ), .ZN(new_n1019_));
  NOR2_X1    g0634(.A1(new_n1018_), .A2(new_n1019_), .ZN(new_n1020_));
  NOR2_X1    g0635(.A1(\req[10] ), .A2(\req[11] ), .ZN(new_n1021_));
  NAND2_X1   g0636(.A1(\priority[10] ), .A2(\req[9] ), .ZN(new_n1022_));
  NOR2_X1    g0637(.A1(\priority[12] ), .A2(\priority[13] ), .ZN(new_n1023_));
  NAND2_X1   g0638(.A1(\priority[11] ), .A2(\req[11] ), .ZN(new_n1024_));
  NOR4_X1    g0639(.A1(new_n1021_), .A2(new_n1022_), .A3(new_n1023_), .A4(new_n1024_), .ZN(new_n1025_));
  NOR2_X1    g0640(.A1(\req[13] ), .A2(\req[14] ), .ZN(new_n1026_));
  NAND2_X1   g0641(.A1(\priority[13] ), .A2(\req[12] ), .ZN(new_n1027_));
  NOR2_X1    g0642(.A1(new_n1026_), .A2(new_n1027_), .ZN(new_n1028_));
  NOR2_X1    g0643(.A1(\priority[15] ), .A2(\priority[16] ), .ZN(new_n1029_));
  NAND2_X1   g0644(.A1(\priority[14] ), .A2(\req[14] ), .ZN(new_n1030_));
  NOR2_X1    g0645(.A1(\req[16] ), .A2(\req[17] ), .ZN(new_n1031_));
  NAND2_X1   g0646(.A1(\priority[16] ), .A2(\req[15] ), .ZN(new_n1032_));
  NOR4_X1    g0647(.A1(new_n1029_), .A2(new_n1030_), .A3(new_n1031_), .A4(new_n1032_), .ZN(new_n1033_));
  OAI22_X1   g0648(.A1(new_n1020_), .A2(new_n1025_), .B1(new_n1033_), .B2(new_n1028_), .ZN(new_n1034_));
  NOR2_X1    g0649(.A1(\priority[18] ), .A2(\priority[19] ), .ZN(new_n1035_));
  NAND2_X1   g0650(.A1(\priority[17] ), .A2(\req[17] ), .ZN(new_n1036_));
  NOR2_X1    g0651(.A1(new_n1035_), .A2(new_n1036_), .ZN(new_n1037_));
  NOR2_X1    g0652(.A1(\req[19] ), .A2(\req[20] ), .ZN(new_n1038_));
  NAND2_X1   g0653(.A1(\priority[19] ), .A2(\req[18] ), .ZN(new_n1039_));
  NOR2_X1    g0654(.A1(\priority[21] ), .A2(\priority[22] ), .ZN(new_n1040_));
  NAND2_X1   g0655(.A1(\priority[20] ), .A2(\req[20] ), .ZN(new_n1041_));
  NOR4_X1    g0656(.A1(new_n1038_), .A2(new_n1039_), .A3(new_n1040_), .A4(new_n1041_), .ZN(new_n1042_));
  NOR2_X1    g0657(.A1(\req[22] ), .A2(\req[23] ), .ZN(new_n1043_));
  NAND2_X1   g0658(.A1(\priority[22] ), .A2(\req[21] ), .ZN(new_n1044_));
  NOR2_X1    g0659(.A1(new_n1043_), .A2(new_n1044_), .ZN(new_n1045_));
  NOR2_X1    g0660(.A1(\priority[24] ), .A2(\priority[25] ), .ZN(new_n1046_));
  NAND2_X1   g0661(.A1(\priority[23] ), .A2(\req[23] ), .ZN(new_n1047_));
  NOR2_X1    g0662(.A1(\req[25] ), .A2(\req[26] ), .ZN(new_n1048_));
  NAND2_X1   g0663(.A1(\priority[25] ), .A2(\req[24] ), .ZN(new_n1049_));
  NOR4_X1    g0664(.A1(new_n1046_), .A2(new_n1047_), .A3(new_n1048_), .A4(new_n1049_), .ZN(new_n1050_));
  OAI22_X1   g0665(.A1(new_n1037_), .A2(new_n1042_), .B1(new_n1050_), .B2(new_n1045_), .ZN(new_n1051_));
  NOR3_X1    g0666(.A1(new_n1034_), .A2(new_n1051_), .A3(new_n1017_), .ZN(new_n1052_));
  NOR2_X1    g0667(.A1(\priority[45] ), .A2(\priority[46] ), .ZN(new_n1053_));
  NAND2_X1   g0668(.A1(\priority[44] ), .A2(\req[44] ), .ZN(new_n1054_));
  NOR2_X1    g0669(.A1(new_n1053_), .A2(new_n1054_), .ZN(new_n1055_));
  NOR2_X1    g0670(.A1(\req[46] ), .A2(\req[47] ), .ZN(new_n1056_));
  NAND2_X1   g0671(.A1(\priority[46] ), .A2(\req[45] ), .ZN(new_n1057_));
  NOR2_X1    g0672(.A1(\priority[48] ), .A2(\priority[49] ), .ZN(new_n1058_));
  NAND2_X1   g0673(.A1(\priority[47] ), .A2(\req[47] ), .ZN(new_n1059_));
  NOR4_X1    g0674(.A1(new_n1056_), .A2(new_n1057_), .A3(new_n1058_), .A4(new_n1059_), .ZN(new_n1060_));
  NOR2_X1    g0675(.A1(\req[49] ), .A2(\req[50] ), .ZN(new_n1061_));
  NAND2_X1   g0676(.A1(\priority[49] ), .A2(\req[48] ), .ZN(new_n1062_));
  NOR2_X1    g0677(.A1(new_n1061_), .A2(new_n1062_), .ZN(new_n1063_));
  NOR2_X1    g0678(.A1(\priority[51] ), .A2(\priority[52] ), .ZN(new_n1064_));
  NAND2_X1   g0679(.A1(\priority[50] ), .A2(\req[50] ), .ZN(new_n1065_));
  NOR2_X1    g0680(.A1(\req[52] ), .A2(\req[53] ), .ZN(new_n1066_));
  NAND2_X1   g0681(.A1(\priority[52] ), .A2(\req[51] ), .ZN(new_n1067_));
  NOR4_X1    g0682(.A1(new_n1064_), .A2(new_n1065_), .A3(new_n1066_), .A4(new_n1067_), .ZN(new_n1068_));
  OAI22_X1   g0683(.A1(new_n1055_), .A2(new_n1060_), .B1(new_n1068_), .B2(new_n1063_), .ZN(new_n1069_));
  NOR2_X1    g0684(.A1(\priority[54] ), .A2(\priority[55] ), .ZN(new_n1070_));
  NAND2_X1   g0685(.A1(\priority[53] ), .A2(\req[53] ), .ZN(new_n1071_));
  NOR2_X1    g0686(.A1(new_n1070_), .A2(new_n1071_), .ZN(new_n1072_));
  NOR2_X1    g0687(.A1(\req[55] ), .A2(\req[56] ), .ZN(new_n1073_));
  NAND2_X1   g0688(.A1(\priority[55] ), .A2(\req[54] ), .ZN(new_n1074_));
  NOR2_X1    g0689(.A1(\priority[57] ), .A2(\priority[58] ), .ZN(new_n1075_));
  NAND2_X1   g0690(.A1(\priority[56] ), .A2(\req[56] ), .ZN(new_n1076_));
  NOR4_X1    g0691(.A1(new_n1073_), .A2(new_n1074_), .A3(new_n1075_), .A4(new_n1076_), .ZN(new_n1077_));
  NOR2_X1    g0692(.A1(\req[58] ), .A2(\req[59] ), .ZN(new_n1078_));
  NAND2_X1   g0693(.A1(\priority[58] ), .A2(\req[57] ), .ZN(new_n1079_));
  NOR2_X1    g0694(.A1(new_n1078_), .A2(new_n1079_), .ZN(new_n1080_));
  NOR2_X1    g0695(.A1(\priority[60] ), .A2(\priority[61] ), .ZN(new_n1081_));
  NAND2_X1   g0696(.A1(\priority[59] ), .A2(\req[59] ), .ZN(new_n1082_));
  NOR2_X1    g0697(.A1(\req[61] ), .A2(\req[62] ), .ZN(new_n1083_));
  NAND2_X1   g0698(.A1(\priority[61] ), .A2(\req[60] ), .ZN(new_n1084_));
  NOR4_X1    g0699(.A1(new_n1081_), .A2(new_n1082_), .A3(new_n1083_), .A4(new_n1084_), .ZN(new_n1085_));
  OAI22_X1   g0700(.A1(new_n1072_), .A2(new_n1077_), .B1(new_n1085_), .B2(new_n1080_), .ZN(new_n1086_));
  NOR2_X1    g0701(.A1(\priority[27] ), .A2(\priority[28] ), .ZN(new_n1087_));
  NAND2_X1   g0702(.A1(\priority[26] ), .A2(\req[26] ), .ZN(new_n1088_));
  NOR2_X1    g0703(.A1(new_n1087_), .A2(new_n1088_), .ZN(new_n1089_));
  NOR2_X1    g0704(.A1(\req[28] ), .A2(\req[29] ), .ZN(new_n1090_));
  NAND2_X1   g0705(.A1(\priority[28] ), .A2(\req[27] ), .ZN(new_n1091_));
  NOR2_X1    g0706(.A1(\priority[30] ), .A2(\priority[31] ), .ZN(new_n1092_));
  NAND2_X1   g0707(.A1(\priority[29] ), .A2(\req[29] ), .ZN(new_n1093_));
  NOR4_X1    g0708(.A1(new_n1090_), .A2(new_n1091_), .A3(new_n1092_), .A4(new_n1093_), .ZN(new_n1094_));
  NOR2_X1    g0709(.A1(\req[31] ), .A2(\req[32] ), .ZN(new_n1095_));
  NAND2_X1   g0710(.A1(\priority[31] ), .A2(\req[30] ), .ZN(new_n1096_));
  NOR2_X1    g0711(.A1(new_n1095_), .A2(new_n1096_), .ZN(new_n1097_));
  NOR2_X1    g0712(.A1(\priority[33] ), .A2(\priority[34] ), .ZN(new_n1098_));
  NAND2_X1   g0713(.A1(\priority[32] ), .A2(\req[32] ), .ZN(new_n1099_));
  NOR2_X1    g0714(.A1(\req[34] ), .A2(\req[35] ), .ZN(new_n1100_));
  NAND2_X1   g0715(.A1(\priority[34] ), .A2(\req[33] ), .ZN(new_n1101_));
  NOR4_X1    g0716(.A1(new_n1098_), .A2(new_n1099_), .A3(new_n1100_), .A4(new_n1101_), .ZN(new_n1102_));
  OAI22_X1   g0717(.A1(new_n1089_), .A2(new_n1094_), .B1(new_n1102_), .B2(new_n1097_), .ZN(new_n1103_));
  NOR2_X1    g0718(.A1(\priority[36] ), .A2(\priority[37] ), .ZN(new_n1104_));
  NAND2_X1   g0719(.A1(\priority[35] ), .A2(\req[35] ), .ZN(new_n1105_));
  NOR2_X1    g0720(.A1(new_n1104_), .A2(new_n1105_), .ZN(new_n1106_));
  NOR2_X1    g0721(.A1(\req[37] ), .A2(\req[38] ), .ZN(new_n1107_));
  NAND2_X1   g0722(.A1(\priority[37] ), .A2(\req[36] ), .ZN(new_n1108_));
  NOR2_X1    g0723(.A1(\priority[39] ), .A2(\priority[40] ), .ZN(new_n1109_));
  NAND2_X1   g0724(.A1(\priority[38] ), .A2(\req[38] ), .ZN(new_n1110_));
  NOR4_X1    g0725(.A1(new_n1107_), .A2(new_n1108_), .A3(new_n1109_), .A4(new_n1110_), .ZN(new_n1111_));
  NOR2_X1    g0726(.A1(\req[40] ), .A2(\req[41] ), .ZN(new_n1112_));
  NAND2_X1   g0727(.A1(\priority[40] ), .A2(\req[39] ), .ZN(new_n1113_));
  NOR2_X1    g0728(.A1(new_n1112_), .A2(new_n1113_), .ZN(new_n1114_));
  NOR2_X1    g0729(.A1(\priority[42] ), .A2(\priority[43] ), .ZN(new_n1115_));
  NAND2_X1   g0730(.A1(\priority[41] ), .A2(\req[41] ), .ZN(new_n1116_));
  NOR2_X1    g0731(.A1(\req[43] ), .A2(\req[44] ), .ZN(new_n1117_));
  NAND2_X1   g0732(.A1(\priority[43] ), .A2(\req[42] ), .ZN(new_n1118_));
  NOR4_X1    g0733(.A1(new_n1115_), .A2(new_n1116_), .A3(new_n1117_), .A4(new_n1118_), .ZN(new_n1119_));
  OAI22_X1   g0734(.A1(new_n1106_), .A2(new_n1111_), .B1(new_n1119_), .B2(new_n1114_), .ZN(new_n1120_));
  NOR4_X1    g0735(.A1(new_n1069_), .A2(new_n1086_), .A3(new_n1103_), .A4(new_n1120_), .ZN(new_n1121_));
  NAND4_X1   g0736(.A1(new_n947_), .A2(new_n1121_), .A3(new_n1008_), .A4(new_n1052_), .ZN(new_n1122_));
  NAND2_X1   g0737(.A1(\priority[2] ), .A2(\req[1] ), .ZN(new_n1123_));
  AOI21_X1   g0738(.A1(new_n1122_), .A2(new_n769_), .B(new_n1123_), .ZN(\grant[2] ));
  NOR2_X1    g0739(.A1(new_n392_), .A2(new_n393_), .ZN(new_n1125_));
  NOR2_X1    g0740(.A1(new_n400_), .A2(new_n401_), .ZN(new_n1126_));
  NOR4_X1    g0741(.A1(new_n395_), .A2(new_n396_), .A3(new_n398_), .A4(new_n399_), .ZN(new_n1127_));
  NOR4_X1    g0742(.A1(new_n404_), .A2(new_n405_), .A3(new_n407_), .A4(new_n408_), .ZN(new_n1128_));
  OAI22_X1   g0743(.A1(new_n1125_), .A2(new_n1127_), .B1(new_n1128_), .B2(new_n1126_), .ZN(new_n1129_));
  NOR2_X1    g0744(.A1(new_n409_), .A2(new_n410_), .ZN(new_n1130_));
  NOR2_X1    g0745(.A1(new_n417_), .A2(new_n418_), .ZN(new_n1131_));
  NOR4_X1    g0746(.A1(new_n412_), .A2(new_n413_), .A3(new_n415_), .A4(new_n416_), .ZN(new_n1132_));
  NOR4_X1    g0747(.A1(new_n482_), .A2(new_n483_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n1133_));
  OAI22_X1   g0748(.A1(new_n1130_), .A2(new_n1132_), .B1(new_n1133_), .B2(new_n1131_), .ZN(new_n1134_));
  NOR2_X1    g0749(.A1(new_n426_), .A2(new_n427_), .ZN(new_n1135_));
  NOR2_X1    g0750(.A1(new_n434_), .A2(new_n435_), .ZN(new_n1136_));
  NOR4_X1    g0751(.A1(new_n429_), .A2(new_n430_), .A3(new_n432_), .A4(new_n433_), .ZN(new_n1137_));
  NOR4_X1    g0752(.A1(new_n438_), .A2(new_n439_), .A3(new_n441_), .A4(new_n442_), .ZN(new_n1138_));
  OAI22_X1   g0753(.A1(new_n1135_), .A2(new_n1137_), .B1(new_n1138_), .B2(new_n1136_), .ZN(new_n1139_));
  NOR2_X1    g0754(.A1(new_n443_), .A2(new_n444_), .ZN(new_n1140_));
  NOR2_X1    g0755(.A1(new_n451_), .A2(new_n452_), .ZN(new_n1141_));
  NOR4_X1    g0756(.A1(new_n446_), .A2(new_n447_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n1142_));
  NOR4_X1    g0757(.A1(new_n387_), .A2(new_n388_), .A3(new_n390_), .A4(new_n391_), .ZN(new_n1143_));
  OAI22_X1   g0758(.A1(new_n1140_), .A2(new_n1142_), .B1(new_n1143_), .B2(new_n1141_), .ZN(new_n1144_));
  NOR4_X1    g0759(.A1(new_n1129_), .A2(new_n1134_), .A3(new_n1139_), .A4(new_n1144_), .ZN(new_n1145_));
  NOR2_X1    g0760(.A1(new_n461_), .A2(new_n462_), .ZN(new_n1146_));
  NOR2_X1    g0761(.A1(\req[0] ), .A2(\req[1] ), .ZN(new_n1147_));
  NOR2_X1    g0762(.A1(\priority[2] ), .A2(\priority[3] ), .ZN(new_n1148_));
  NAND2_X1   g0763(.A1(\priority[1] ), .A2(\req[1] ), .ZN(new_n1149_));
  NOR4_X1    g0764(.A1(new_n631_), .A2(new_n1147_), .A3(new_n1148_), .A4(new_n1149_), .ZN(new_n1150_));
  NOR2_X1    g0765(.A1(new_n1150_), .A2(new_n1146_), .ZN(new_n1151_));
  NOR2_X1    g0766(.A1(new_n470_), .A2(new_n471_), .ZN(new_n1152_));
  NOR2_X1    g0767(.A1(new_n478_), .A2(new_n479_), .ZN(new_n1153_));
  NOR4_X1    g0768(.A1(new_n473_), .A2(new_n474_), .A3(new_n476_), .A4(new_n477_), .ZN(new_n1154_));
  NOR4_X1    g0769(.A1(new_n456_), .A2(new_n457_), .A3(new_n459_), .A4(new_n460_), .ZN(new_n1155_));
  OAI22_X1   g0770(.A1(new_n1152_), .A2(new_n1154_), .B1(new_n1155_), .B2(new_n1153_), .ZN(new_n1156_));
  NOR2_X1    g0771(.A1(new_n487_), .A2(new_n488_), .ZN(new_n1157_));
  NOR2_X1    g0772(.A1(new_n495_), .A2(new_n496_), .ZN(new_n1158_));
  NOR4_X1    g0773(.A1(new_n490_), .A2(new_n491_), .A3(new_n493_), .A4(new_n494_), .ZN(new_n1159_));
  NOR4_X1    g0774(.A1(new_n499_), .A2(new_n500_), .A3(new_n502_), .A4(new_n503_), .ZN(new_n1160_));
  OAI22_X1   g0775(.A1(new_n1157_), .A2(new_n1159_), .B1(new_n1160_), .B2(new_n1158_), .ZN(new_n1161_));
  NOR2_X1    g0776(.A1(new_n504_), .A2(new_n505_), .ZN(new_n1162_));
  NOR2_X1    g0777(.A1(new_n512_), .A2(new_n513_), .ZN(new_n1163_));
  NOR4_X1    g0778(.A1(new_n507_), .A2(new_n508_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n1164_));
  NOR4_X1    g0779(.A1(new_n465_), .A2(new_n466_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n1165_));
  OAI22_X1   g0780(.A1(new_n1162_), .A2(new_n1164_), .B1(new_n1165_), .B2(new_n1163_), .ZN(new_n1166_));
  NOR4_X1    g0781(.A1(new_n1156_), .A2(new_n1161_), .A3(new_n1166_), .A4(new_n1151_), .ZN(new_n1167_));
  NOR4_X1    g0782(.A1(new_n526_), .A2(new_n527_), .A3(new_n529_), .A4(new_n530_), .ZN(new_n1168_));
  INV_X1     g0783(.I(\req[4] ), .ZN(new_n1169_));
  AOI21_X1   g0784(.A1(new_n1169_), .A2(\priority[4] ), .B(\priority[5] ), .ZN(new_n1170_));
  OAI21_X1   g0785(.A1(new_n1168_), .A2(new_n520_), .B(new_n1170_), .ZN(new_n1171_));
  NOR2_X1    g0786(.A1(new_n531_), .A2(new_n532_), .ZN(new_n1172_));
  NOR2_X1    g0787(.A1(new_n539_), .A2(new_n540_), .ZN(new_n1173_));
  NOR4_X1    g0788(.A1(new_n534_), .A2(new_n535_), .A3(new_n537_), .A4(new_n538_), .ZN(new_n1174_));
  NOR4_X1    g0789(.A1(new_n543_), .A2(new_n544_), .A3(new_n546_), .A4(new_n547_), .ZN(new_n1175_));
  OAI22_X1   g0790(.A1(new_n1172_), .A2(new_n1174_), .B1(new_n1175_), .B2(new_n1173_), .ZN(new_n1176_));
  NOR2_X1    g0791(.A1(new_n548_), .A2(new_n549_), .ZN(new_n1177_));
  NOR2_X1    g0792(.A1(new_n556_), .A2(new_n557_), .ZN(new_n1178_));
  NOR4_X1    g0793(.A1(new_n551_), .A2(new_n552_), .A3(new_n554_), .A4(new_n555_), .ZN(new_n1179_));
  NOR4_X1    g0794(.A1(new_n595_), .A2(new_n596_), .A3(new_n598_), .A4(new_n599_), .ZN(new_n1180_));
  OAI22_X1   g0795(.A1(new_n1177_), .A2(new_n1179_), .B1(new_n1180_), .B2(new_n1178_), .ZN(new_n1181_));
  NOR3_X1    g0796(.A1(new_n1176_), .A2(new_n1181_), .A3(new_n1171_), .ZN(new_n1182_));
  NOR2_X1    g0797(.A1(new_n566_), .A2(new_n567_), .ZN(new_n1183_));
  NOR2_X1    g0798(.A1(new_n574_), .A2(new_n575_), .ZN(new_n1184_));
  NOR4_X1    g0799(.A1(new_n569_), .A2(new_n570_), .A3(new_n572_), .A4(new_n573_), .ZN(new_n1185_));
  NOR4_X1    g0800(.A1(new_n578_), .A2(new_n579_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n1186_));
  OAI22_X1   g0801(.A1(new_n1183_), .A2(new_n1185_), .B1(new_n1186_), .B2(new_n1184_), .ZN(new_n1187_));
  NOR2_X1    g0802(.A1(new_n583_), .A2(new_n584_), .ZN(new_n1188_));
  NOR2_X1    g0803(.A1(new_n591_), .A2(new_n592_), .ZN(new_n1189_));
  NOR4_X1    g0804(.A1(new_n586_), .A2(new_n587_), .A3(new_n589_), .A4(new_n590_), .ZN(new_n1190_));
  NOR4_X1    g0805(.A1(new_n421_), .A2(new_n422_), .A3(new_n424_), .A4(new_n425_), .ZN(new_n1191_));
  OAI22_X1   g0806(.A1(new_n1188_), .A2(new_n1190_), .B1(new_n1191_), .B2(new_n1189_), .ZN(new_n1192_));
  NOR2_X1    g0807(.A1(new_n600_), .A2(new_n601_), .ZN(new_n1193_));
  NOR2_X1    g0808(.A1(new_n608_), .A2(new_n609_), .ZN(new_n1194_));
  NOR4_X1    g0809(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .A4(new_n607_), .ZN(new_n1195_));
  NOR4_X1    g0810(.A1(new_n612_), .A2(new_n613_), .A3(new_n615_), .A4(new_n616_), .ZN(new_n1196_));
  OAI22_X1   g0811(.A1(new_n1193_), .A2(new_n1195_), .B1(new_n1196_), .B2(new_n1194_), .ZN(new_n1197_));
  NOR2_X1    g0812(.A1(new_n617_), .A2(new_n618_), .ZN(new_n1198_));
  NOR2_X1    g0813(.A1(new_n625_), .A2(new_n626_), .ZN(new_n1199_));
  NOR4_X1    g0814(.A1(new_n620_), .A2(new_n621_), .A3(new_n623_), .A4(new_n624_), .ZN(new_n1200_));
  NOR4_X1    g0815(.A1(new_n561_), .A2(new_n562_), .A3(new_n564_), .A4(new_n565_), .ZN(new_n1201_));
  OAI22_X1   g0816(.A1(new_n1198_), .A2(new_n1200_), .B1(new_n1201_), .B2(new_n1199_), .ZN(new_n1202_));
  NOR4_X1    g0817(.A1(new_n1187_), .A2(new_n1192_), .A3(new_n1197_), .A4(new_n1202_), .ZN(new_n1203_));
  NAND4_X1   g0818(.A1(new_n1145_), .A2(new_n1203_), .A3(new_n1167_), .A4(new_n1182_), .ZN(new_n1204_));
  NAND2_X1   g0819(.A1(\priority[3] ), .A2(\req[2] ), .ZN(new_n1205_));
  AOI21_X1   g0820(.A1(new_n1204_), .A2(new_n1015_), .B(new_n1205_), .ZN(\grant[3] ));
  NOR2_X1    g0821(.A1(new_n638_), .A2(new_n639_), .ZN(new_n1207_));
  NOR2_X1    g0822(.A1(new_n646_), .A2(new_n647_), .ZN(new_n1208_));
  NOR4_X1    g0823(.A1(new_n641_), .A2(new_n642_), .A3(new_n644_), .A4(new_n645_), .ZN(new_n1209_));
  NOR4_X1    g0824(.A1(new_n650_), .A2(new_n651_), .A3(new_n653_), .A4(new_n654_), .ZN(new_n1210_));
  OAI22_X1   g0825(.A1(new_n1207_), .A2(new_n1209_), .B1(new_n1210_), .B2(new_n1208_), .ZN(new_n1211_));
  NOR2_X1    g0826(.A1(new_n655_), .A2(new_n656_), .ZN(new_n1212_));
  NOR2_X1    g0827(.A1(new_n663_), .A2(new_n664_), .ZN(new_n1213_));
  NOR4_X1    g0828(.A1(new_n658_), .A2(new_n659_), .A3(new_n661_), .A4(new_n662_), .ZN(new_n1214_));
  NOR4_X1    g0829(.A1(new_n728_), .A2(new_n729_), .A3(new_n731_), .A4(new_n732_), .ZN(new_n1215_));
  OAI22_X1   g0830(.A1(new_n1212_), .A2(new_n1214_), .B1(new_n1215_), .B2(new_n1213_), .ZN(new_n1216_));
  NOR2_X1    g0831(.A1(new_n672_), .A2(new_n673_), .ZN(new_n1217_));
  NOR2_X1    g0832(.A1(new_n680_), .A2(new_n681_), .ZN(new_n1218_));
  NOR4_X1    g0833(.A1(new_n675_), .A2(new_n676_), .A3(new_n678_), .A4(new_n679_), .ZN(new_n1219_));
  NOR4_X1    g0834(.A1(new_n684_), .A2(new_n685_), .A3(new_n687_), .A4(new_n688_), .ZN(new_n1220_));
  OAI22_X1   g0835(.A1(new_n1217_), .A2(new_n1219_), .B1(new_n1220_), .B2(new_n1218_), .ZN(new_n1221_));
  NOR2_X1    g0836(.A1(new_n689_), .A2(new_n690_), .ZN(new_n1222_));
  NOR2_X1    g0837(.A1(new_n697_), .A2(new_n698_), .ZN(new_n1223_));
  NOR4_X1    g0838(.A1(new_n692_), .A2(new_n693_), .A3(new_n695_), .A4(new_n696_), .ZN(new_n1224_));
  NOR4_X1    g0839(.A1(new_n633_), .A2(new_n634_), .A3(new_n636_), .A4(new_n637_), .ZN(new_n1225_));
  OAI22_X1   g0840(.A1(new_n1222_), .A2(new_n1224_), .B1(new_n1225_), .B2(new_n1223_), .ZN(new_n1226_));
  NOR4_X1    g0841(.A1(new_n1211_), .A2(new_n1216_), .A3(new_n1221_), .A4(new_n1226_), .ZN(new_n1227_));
  NOR2_X1    g0842(.A1(new_n707_), .A2(new_n708_), .ZN(new_n1228_));
  NOR2_X1    g0843(.A1(\req[1] ), .A2(\req[2] ), .ZN(new_n1229_));
  NOR2_X1    g0844(.A1(\priority[3] ), .A2(\priority[4] ), .ZN(new_n1230_));
  NAND2_X1   g0845(.A1(\priority[2] ), .A2(\req[2] ), .ZN(new_n1231_));
  NOR4_X1    g0846(.A1(new_n877_), .A2(new_n1229_), .A3(new_n1230_), .A4(new_n1231_), .ZN(new_n1232_));
  NOR2_X1    g0847(.A1(new_n1232_), .A2(new_n1228_), .ZN(new_n1233_));
  NOR2_X1    g0848(.A1(new_n716_), .A2(new_n717_), .ZN(new_n1234_));
  NOR2_X1    g0849(.A1(new_n724_), .A2(new_n725_), .ZN(new_n1235_));
  NOR4_X1    g0850(.A1(new_n719_), .A2(new_n720_), .A3(new_n722_), .A4(new_n723_), .ZN(new_n1236_));
  NOR4_X1    g0851(.A1(new_n702_), .A2(new_n703_), .A3(new_n705_), .A4(new_n706_), .ZN(new_n1237_));
  OAI22_X1   g0852(.A1(new_n1234_), .A2(new_n1236_), .B1(new_n1237_), .B2(new_n1235_), .ZN(new_n1238_));
  NOR2_X1    g0853(.A1(new_n733_), .A2(new_n734_), .ZN(new_n1239_));
  NOR2_X1    g0854(.A1(new_n741_), .A2(new_n742_), .ZN(new_n1240_));
  NOR4_X1    g0855(.A1(new_n736_), .A2(new_n737_), .A3(new_n739_), .A4(new_n740_), .ZN(new_n1241_));
  NOR4_X1    g0856(.A1(new_n745_), .A2(new_n746_), .A3(new_n748_), .A4(new_n749_), .ZN(new_n1242_));
  OAI22_X1   g0857(.A1(new_n1239_), .A2(new_n1241_), .B1(new_n1242_), .B2(new_n1240_), .ZN(new_n1243_));
  NOR2_X1    g0858(.A1(new_n750_), .A2(new_n751_), .ZN(new_n1244_));
  NOR2_X1    g0859(.A1(new_n758_), .A2(new_n759_), .ZN(new_n1245_));
  NOR4_X1    g0860(.A1(new_n753_), .A2(new_n754_), .A3(new_n756_), .A4(new_n757_), .ZN(new_n1246_));
  NOR4_X1    g0861(.A1(new_n711_), .A2(new_n712_), .A3(new_n714_), .A4(new_n715_), .ZN(new_n1247_));
  OAI22_X1   g0862(.A1(new_n1244_), .A2(new_n1246_), .B1(new_n1247_), .B2(new_n1245_), .ZN(new_n1248_));
  NOR4_X1    g0863(.A1(new_n1238_), .A2(new_n1243_), .A3(new_n1248_), .A4(new_n1233_), .ZN(new_n1249_));
  NOR4_X1    g0864(.A1(new_n772_), .A2(new_n773_), .A3(new_n775_), .A4(new_n776_), .ZN(new_n1250_));
  INV_X1     g0865(.I(\req[5] ), .ZN(new_n1251_));
  AOI21_X1   g0866(.A1(new_n1251_), .A2(\priority[5] ), .B(\priority[6] ), .ZN(new_n1252_));
  OAI21_X1   g0867(.A1(new_n1250_), .A2(new_n766_), .B(new_n1252_), .ZN(new_n1253_));
  NOR2_X1    g0868(.A1(new_n777_), .A2(new_n778_), .ZN(new_n1254_));
  NOR2_X1    g0869(.A1(new_n785_), .A2(new_n786_), .ZN(new_n1255_));
  NOR4_X1    g0870(.A1(new_n780_), .A2(new_n781_), .A3(new_n783_), .A4(new_n784_), .ZN(new_n1256_));
  NOR4_X1    g0871(.A1(new_n789_), .A2(new_n790_), .A3(new_n792_), .A4(new_n793_), .ZN(new_n1257_));
  OAI22_X1   g0872(.A1(new_n1254_), .A2(new_n1256_), .B1(new_n1257_), .B2(new_n1255_), .ZN(new_n1258_));
  NOR2_X1    g0873(.A1(new_n794_), .A2(new_n795_), .ZN(new_n1259_));
  NOR2_X1    g0874(.A1(new_n802_), .A2(new_n803_), .ZN(new_n1260_));
  NOR4_X1    g0875(.A1(new_n797_), .A2(new_n798_), .A3(new_n800_), .A4(new_n801_), .ZN(new_n1261_));
  NOR4_X1    g0876(.A1(new_n841_), .A2(new_n842_), .A3(new_n844_), .A4(new_n845_), .ZN(new_n1262_));
  OAI22_X1   g0877(.A1(new_n1259_), .A2(new_n1261_), .B1(new_n1262_), .B2(new_n1260_), .ZN(new_n1263_));
  NOR3_X1    g0878(.A1(new_n1258_), .A2(new_n1263_), .A3(new_n1253_), .ZN(new_n1264_));
  NOR2_X1    g0879(.A1(new_n812_), .A2(new_n813_), .ZN(new_n1265_));
  NOR2_X1    g0880(.A1(new_n820_), .A2(new_n821_), .ZN(new_n1266_));
  NOR4_X1    g0881(.A1(new_n815_), .A2(new_n816_), .A3(new_n818_), .A4(new_n819_), .ZN(new_n1267_));
  NOR4_X1    g0882(.A1(new_n824_), .A2(new_n825_), .A3(new_n827_), .A4(new_n828_), .ZN(new_n1268_));
  OAI22_X1   g0883(.A1(new_n1265_), .A2(new_n1267_), .B1(new_n1268_), .B2(new_n1266_), .ZN(new_n1269_));
  NOR2_X1    g0884(.A1(new_n829_), .A2(new_n830_), .ZN(new_n1270_));
  NOR2_X1    g0885(.A1(new_n837_), .A2(new_n838_), .ZN(new_n1271_));
  NOR4_X1    g0886(.A1(new_n832_), .A2(new_n833_), .A3(new_n835_), .A4(new_n836_), .ZN(new_n1272_));
  NOR4_X1    g0887(.A1(new_n667_), .A2(new_n668_), .A3(new_n670_), .A4(new_n671_), .ZN(new_n1273_));
  OAI22_X1   g0888(.A1(new_n1270_), .A2(new_n1272_), .B1(new_n1273_), .B2(new_n1271_), .ZN(new_n1274_));
  NOR2_X1    g0889(.A1(new_n846_), .A2(new_n847_), .ZN(new_n1275_));
  NOR2_X1    g0890(.A1(new_n854_), .A2(new_n855_), .ZN(new_n1276_));
  NOR4_X1    g0891(.A1(new_n849_), .A2(new_n850_), .A3(new_n852_), .A4(new_n853_), .ZN(new_n1277_));
  NOR4_X1    g0892(.A1(new_n858_), .A2(new_n859_), .A3(new_n861_), .A4(new_n862_), .ZN(new_n1278_));
  OAI22_X1   g0893(.A1(new_n1275_), .A2(new_n1277_), .B1(new_n1278_), .B2(new_n1276_), .ZN(new_n1279_));
  NOR2_X1    g0894(.A1(new_n863_), .A2(new_n864_), .ZN(new_n1280_));
  NOR2_X1    g0895(.A1(new_n871_), .A2(new_n872_), .ZN(new_n1281_));
  NOR4_X1    g0896(.A1(new_n866_), .A2(new_n867_), .A3(new_n869_), .A4(new_n870_), .ZN(new_n1282_));
  NOR4_X1    g0897(.A1(new_n807_), .A2(new_n808_), .A3(new_n810_), .A4(new_n811_), .ZN(new_n1283_));
  OAI22_X1   g0898(.A1(new_n1280_), .A2(new_n1282_), .B1(new_n1283_), .B2(new_n1281_), .ZN(new_n1284_));
  NOR4_X1    g0899(.A1(new_n1269_), .A2(new_n1274_), .A3(new_n1279_), .A4(new_n1284_), .ZN(new_n1285_));
  NAND4_X1   g0900(.A1(new_n1227_), .A2(new_n1285_), .A3(new_n1249_), .A4(new_n1264_), .ZN(new_n1286_));
  NAND2_X1   g0901(.A1(\priority[4] ), .A2(\req[3] ), .ZN(new_n1287_));
  AOI21_X1   g0902(.A1(new_n1286_), .A2(new_n1169_), .B(new_n1287_), .ZN(\grant[4] ));
  NOR2_X1    g0903(.A1(new_n884_), .A2(new_n885_), .ZN(new_n1289_));
  NOR2_X1    g0904(.A1(new_n892_), .A2(new_n893_), .ZN(new_n1290_));
  NOR4_X1    g0905(.A1(new_n887_), .A2(new_n888_), .A3(new_n890_), .A4(new_n891_), .ZN(new_n1291_));
  NOR4_X1    g0906(.A1(new_n896_), .A2(new_n897_), .A3(new_n899_), .A4(new_n900_), .ZN(new_n1292_));
  OAI22_X1   g0907(.A1(new_n1289_), .A2(new_n1291_), .B1(new_n1292_), .B2(new_n1290_), .ZN(new_n1293_));
  NOR2_X1    g0908(.A1(new_n901_), .A2(new_n902_), .ZN(new_n1294_));
  NOR2_X1    g0909(.A1(new_n909_), .A2(new_n910_), .ZN(new_n1295_));
  NOR4_X1    g0910(.A1(new_n904_), .A2(new_n905_), .A3(new_n907_), .A4(new_n908_), .ZN(new_n1296_));
  NOR4_X1    g0911(.A1(new_n974_), .A2(new_n975_), .A3(new_n977_), .A4(new_n978_), .ZN(new_n1297_));
  OAI22_X1   g0912(.A1(new_n1294_), .A2(new_n1296_), .B1(new_n1297_), .B2(new_n1295_), .ZN(new_n1298_));
  NOR2_X1    g0913(.A1(new_n918_), .A2(new_n919_), .ZN(new_n1299_));
  NOR2_X1    g0914(.A1(new_n926_), .A2(new_n927_), .ZN(new_n1300_));
  NOR4_X1    g0915(.A1(new_n921_), .A2(new_n922_), .A3(new_n924_), .A4(new_n925_), .ZN(new_n1301_));
  NOR4_X1    g0916(.A1(new_n930_), .A2(new_n931_), .A3(new_n933_), .A4(new_n934_), .ZN(new_n1302_));
  OAI22_X1   g0917(.A1(new_n1299_), .A2(new_n1301_), .B1(new_n1302_), .B2(new_n1300_), .ZN(new_n1303_));
  NOR2_X1    g0918(.A1(new_n935_), .A2(new_n936_), .ZN(new_n1304_));
  NOR2_X1    g0919(.A1(new_n943_), .A2(new_n944_), .ZN(new_n1305_));
  NOR4_X1    g0920(.A1(new_n938_), .A2(new_n939_), .A3(new_n941_), .A4(new_n942_), .ZN(new_n1306_));
  NOR4_X1    g0921(.A1(new_n879_), .A2(new_n880_), .A3(new_n882_), .A4(new_n883_), .ZN(new_n1307_));
  OAI22_X1   g0922(.A1(new_n1304_), .A2(new_n1306_), .B1(new_n1307_), .B2(new_n1305_), .ZN(new_n1308_));
  NOR4_X1    g0923(.A1(new_n1293_), .A2(new_n1298_), .A3(new_n1303_), .A4(new_n1308_), .ZN(new_n1309_));
  NOR2_X1    g0924(.A1(new_n953_), .A2(new_n954_), .ZN(new_n1310_));
  NOR4_X1    g0925(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .A4(new_n1123_), .ZN(new_n1311_));
  NOR2_X1    g0926(.A1(new_n1311_), .A2(new_n1310_), .ZN(new_n1312_));
  NOR2_X1    g0927(.A1(new_n962_), .A2(new_n963_), .ZN(new_n1313_));
  NOR2_X1    g0928(.A1(new_n970_), .A2(new_n971_), .ZN(new_n1314_));
  NOR4_X1    g0929(.A1(new_n965_), .A2(new_n966_), .A3(new_n968_), .A4(new_n969_), .ZN(new_n1315_));
  NOR4_X1    g0930(.A1(new_n948_), .A2(new_n949_), .A3(new_n951_), .A4(new_n952_), .ZN(new_n1316_));
  OAI22_X1   g0931(.A1(new_n1313_), .A2(new_n1315_), .B1(new_n1316_), .B2(new_n1314_), .ZN(new_n1317_));
  NOR2_X1    g0932(.A1(new_n979_), .A2(new_n980_), .ZN(new_n1318_));
  NOR2_X1    g0933(.A1(new_n987_), .A2(new_n988_), .ZN(new_n1319_));
  NOR4_X1    g0934(.A1(new_n982_), .A2(new_n983_), .A3(new_n985_), .A4(new_n986_), .ZN(new_n1320_));
  NOR4_X1    g0935(.A1(new_n991_), .A2(new_n992_), .A3(new_n994_), .A4(new_n995_), .ZN(new_n1321_));
  OAI22_X1   g0936(.A1(new_n1318_), .A2(new_n1320_), .B1(new_n1321_), .B2(new_n1319_), .ZN(new_n1322_));
  NOR2_X1    g0937(.A1(new_n996_), .A2(new_n997_), .ZN(new_n1323_));
  NOR2_X1    g0938(.A1(new_n1004_), .A2(new_n1005_), .ZN(new_n1324_));
  NOR4_X1    g0939(.A1(new_n999_), .A2(new_n1000_), .A3(new_n1002_), .A4(new_n1003_), .ZN(new_n1325_));
  NOR4_X1    g0940(.A1(new_n957_), .A2(new_n958_), .A3(new_n960_), .A4(new_n961_), .ZN(new_n1326_));
  OAI22_X1   g0941(.A1(new_n1323_), .A2(new_n1325_), .B1(new_n1326_), .B2(new_n1324_), .ZN(new_n1327_));
  NOR4_X1    g0942(.A1(new_n1317_), .A2(new_n1322_), .A3(new_n1327_), .A4(new_n1312_), .ZN(new_n1328_));
  NOR4_X1    g0943(.A1(new_n1018_), .A2(new_n1019_), .A3(new_n1021_), .A4(new_n1022_), .ZN(new_n1329_));
  INV_X1     g0944(.I(\req[6] ), .ZN(new_n1330_));
  AOI21_X1   g0945(.A1(new_n1330_), .A2(\priority[6] ), .B(\priority[7] ), .ZN(new_n1331_));
  OAI21_X1   g0946(.A1(new_n1329_), .A2(new_n1012_), .B(new_n1331_), .ZN(new_n1332_));
  NOR2_X1    g0947(.A1(new_n1023_), .A2(new_n1024_), .ZN(new_n1333_));
  NOR2_X1    g0948(.A1(new_n1031_), .A2(new_n1032_), .ZN(new_n1334_));
  NOR4_X1    g0949(.A1(new_n1026_), .A2(new_n1027_), .A3(new_n1029_), .A4(new_n1030_), .ZN(new_n1335_));
  NOR4_X1    g0950(.A1(new_n1035_), .A2(new_n1036_), .A3(new_n1038_), .A4(new_n1039_), .ZN(new_n1336_));
  OAI22_X1   g0951(.A1(new_n1333_), .A2(new_n1335_), .B1(new_n1336_), .B2(new_n1334_), .ZN(new_n1337_));
  NOR2_X1    g0952(.A1(new_n1040_), .A2(new_n1041_), .ZN(new_n1338_));
  NOR2_X1    g0953(.A1(new_n1048_), .A2(new_n1049_), .ZN(new_n1339_));
  NOR4_X1    g0954(.A1(new_n1043_), .A2(new_n1044_), .A3(new_n1046_), .A4(new_n1047_), .ZN(new_n1340_));
  NOR4_X1    g0955(.A1(new_n1087_), .A2(new_n1088_), .A3(new_n1090_), .A4(new_n1091_), .ZN(new_n1341_));
  OAI22_X1   g0956(.A1(new_n1338_), .A2(new_n1340_), .B1(new_n1341_), .B2(new_n1339_), .ZN(new_n1342_));
  NOR3_X1    g0957(.A1(new_n1337_), .A2(new_n1342_), .A3(new_n1332_), .ZN(new_n1343_));
  NOR2_X1    g0958(.A1(new_n1058_), .A2(new_n1059_), .ZN(new_n1344_));
  NOR2_X1    g0959(.A1(new_n1066_), .A2(new_n1067_), .ZN(new_n1345_));
  NOR4_X1    g0960(.A1(new_n1061_), .A2(new_n1062_), .A3(new_n1064_), .A4(new_n1065_), .ZN(new_n1346_));
  NOR4_X1    g0961(.A1(new_n1070_), .A2(new_n1071_), .A3(new_n1073_), .A4(new_n1074_), .ZN(new_n1347_));
  OAI22_X1   g0962(.A1(new_n1344_), .A2(new_n1346_), .B1(new_n1347_), .B2(new_n1345_), .ZN(new_n1348_));
  NOR2_X1    g0963(.A1(new_n1075_), .A2(new_n1076_), .ZN(new_n1349_));
  NOR2_X1    g0964(.A1(new_n1083_), .A2(new_n1084_), .ZN(new_n1350_));
  NOR4_X1    g0965(.A1(new_n1078_), .A2(new_n1079_), .A3(new_n1081_), .A4(new_n1082_), .ZN(new_n1351_));
  NOR4_X1    g0966(.A1(new_n913_), .A2(new_n914_), .A3(new_n916_), .A4(new_n917_), .ZN(new_n1352_));
  OAI22_X1   g0967(.A1(new_n1349_), .A2(new_n1351_), .B1(new_n1352_), .B2(new_n1350_), .ZN(new_n1353_));
  NOR2_X1    g0968(.A1(new_n1092_), .A2(new_n1093_), .ZN(new_n1354_));
  NOR2_X1    g0969(.A1(new_n1100_), .A2(new_n1101_), .ZN(new_n1355_));
  NOR4_X1    g0970(.A1(new_n1095_), .A2(new_n1096_), .A3(new_n1098_), .A4(new_n1099_), .ZN(new_n1356_));
  NOR4_X1    g0971(.A1(new_n1104_), .A2(new_n1105_), .A3(new_n1107_), .A4(new_n1108_), .ZN(new_n1357_));
  OAI22_X1   g0972(.A1(new_n1354_), .A2(new_n1356_), .B1(new_n1357_), .B2(new_n1355_), .ZN(new_n1358_));
  NOR2_X1    g0973(.A1(new_n1109_), .A2(new_n1110_), .ZN(new_n1359_));
  NOR2_X1    g0974(.A1(new_n1117_), .A2(new_n1118_), .ZN(new_n1360_));
  NOR4_X1    g0975(.A1(new_n1112_), .A2(new_n1113_), .A3(new_n1115_), .A4(new_n1116_), .ZN(new_n1361_));
  NOR4_X1    g0976(.A1(new_n1053_), .A2(new_n1054_), .A3(new_n1056_), .A4(new_n1057_), .ZN(new_n1362_));
  OAI22_X1   g0977(.A1(new_n1359_), .A2(new_n1361_), .B1(new_n1362_), .B2(new_n1360_), .ZN(new_n1363_));
  NOR4_X1    g0978(.A1(new_n1348_), .A2(new_n1353_), .A3(new_n1358_), .A4(new_n1363_), .ZN(new_n1364_));
  NAND4_X1   g0979(.A1(new_n1309_), .A2(new_n1364_), .A3(new_n1328_), .A4(new_n1343_), .ZN(new_n1365_));
  AOI21_X1   g0980(.A1(new_n1365_), .A2(new_n1251_), .B(new_n521_), .ZN(\grant[5] ));
  NOR2_X1    g0981(.A1(new_n398_), .A2(new_n399_), .ZN(new_n1367_));
  NOR2_X1    g0982(.A1(new_n407_), .A2(new_n408_), .ZN(new_n1368_));
  NOR4_X1    g0983(.A1(new_n400_), .A2(new_n401_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n1369_));
  NOR4_X1    g0984(.A1(new_n409_), .A2(new_n410_), .A3(new_n412_), .A4(new_n413_), .ZN(new_n1370_));
  OAI22_X1   g0985(.A1(new_n1367_), .A2(new_n1369_), .B1(new_n1370_), .B2(new_n1368_), .ZN(new_n1371_));
  NOR2_X1    g0986(.A1(new_n415_), .A2(new_n416_), .ZN(new_n1372_));
  NOR2_X1    g0987(.A1(new_n485_), .A2(new_n486_), .ZN(new_n1373_));
  NOR4_X1    g0988(.A1(new_n417_), .A2(new_n418_), .A3(new_n482_), .A4(new_n483_), .ZN(new_n1374_));
  NOR4_X1    g0989(.A1(new_n487_), .A2(new_n488_), .A3(new_n490_), .A4(new_n491_), .ZN(new_n1375_));
  OAI22_X1   g0990(.A1(new_n1372_), .A2(new_n1374_), .B1(new_n1375_), .B2(new_n1373_), .ZN(new_n1376_));
  NOR2_X1    g0991(.A1(new_n432_), .A2(new_n433_), .ZN(new_n1377_));
  NOR2_X1    g0992(.A1(new_n441_), .A2(new_n442_), .ZN(new_n1378_));
  NOR4_X1    g0993(.A1(new_n434_), .A2(new_n435_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n1379_));
  NOR4_X1    g0994(.A1(new_n443_), .A2(new_n444_), .A3(new_n446_), .A4(new_n447_), .ZN(new_n1380_));
  OAI22_X1   g0995(.A1(new_n1377_), .A2(new_n1379_), .B1(new_n1380_), .B2(new_n1378_), .ZN(new_n1381_));
  NOR2_X1    g0996(.A1(new_n390_), .A2(new_n391_), .ZN(new_n1382_));
  NOR2_X1    g0997(.A1(new_n449_), .A2(new_n450_), .ZN(new_n1383_));
  NOR4_X1    g0998(.A1(new_n387_), .A2(new_n388_), .A3(new_n451_), .A4(new_n452_), .ZN(new_n1384_));
  NOR4_X1    g0999(.A1(new_n392_), .A2(new_n393_), .A3(new_n395_), .A4(new_n396_), .ZN(new_n1385_));
  OAI22_X1   g1000(.A1(new_n1382_), .A2(new_n1385_), .B1(new_n1384_), .B2(new_n1383_), .ZN(new_n1386_));
  NOR4_X1    g1001(.A1(new_n1371_), .A2(new_n1376_), .A3(new_n1381_), .A4(new_n1386_), .ZN(new_n1387_));
  NOR2_X1    g1002(.A1(new_n1148_), .A2(new_n1149_), .ZN(new_n1388_));
  NOR4_X1    g1003(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .A4(new_n1205_), .ZN(new_n1389_));
  NOR2_X1    g1004(.A1(new_n1389_), .A2(new_n1388_), .ZN(new_n1390_));
  NOR2_X1    g1005(.A1(new_n459_), .A2(new_n460_), .ZN(new_n1391_));
  NOR2_X1    g1006(.A1(new_n476_), .A2(new_n477_), .ZN(new_n1392_));
  NOR4_X1    g1007(.A1(new_n456_), .A2(new_n457_), .A3(new_n478_), .A4(new_n479_), .ZN(new_n1393_));
  NOR4_X1    g1008(.A1(new_n461_), .A2(new_n462_), .A3(new_n1147_), .A4(new_n631_), .ZN(new_n1394_));
  OAI22_X1   g1009(.A1(new_n1391_), .A2(new_n1394_), .B1(new_n1393_), .B2(new_n1392_), .ZN(new_n1395_));
  NOR2_X1    g1010(.A1(new_n493_), .A2(new_n494_), .ZN(new_n1396_));
  NOR2_X1    g1011(.A1(new_n502_), .A2(new_n503_), .ZN(new_n1397_));
  NOR4_X1    g1012(.A1(new_n495_), .A2(new_n496_), .A3(new_n499_), .A4(new_n500_), .ZN(new_n1398_));
  NOR4_X1    g1013(.A1(new_n504_), .A2(new_n505_), .A3(new_n507_), .A4(new_n508_), .ZN(new_n1399_));
  OAI22_X1   g1014(.A1(new_n1396_), .A2(new_n1398_), .B1(new_n1399_), .B2(new_n1397_), .ZN(new_n1400_));
  NOR2_X1    g1015(.A1(new_n468_), .A2(new_n469_), .ZN(new_n1401_));
  NOR2_X1    g1016(.A1(new_n510_), .A2(new_n511_), .ZN(new_n1402_));
  NOR4_X1    g1017(.A1(new_n465_), .A2(new_n466_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n1403_));
  NOR4_X1    g1018(.A1(new_n470_), .A2(new_n471_), .A3(new_n473_), .A4(new_n474_), .ZN(new_n1404_));
  OAI22_X1   g1019(.A1(new_n1401_), .A2(new_n1404_), .B1(new_n1403_), .B2(new_n1402_), .ZN(new_n1405_));
  NOR4_X1    g1020(.A1(new_n1395_), .A2(new_n1400_), .A3(new_n1405_), .A4(new_n1390_), .ZN(new_n1406_));
  NOR4_X1    g1021(.A1(new_n531_), .A2(new_n532_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n1407_));
  INV_X1     g1022(.I(\req[7] ), .ZN(new_n1408_));
  AOI21_X1   g1023(.A1(new_n1408_), .A2(\priority[7] ), .B(\priority[8] ), .ZN(new_n1409_));
  OAI21_X1   g1024(.A1(new_n1407_), .A2(new_n529_), .B(new_n1409_), .ZN(new_n1410_));
  NOR2_X1    g1025(.A1(new_n537_), .A2(new_n538_), .ZN(new_n1411_));
  NOR2_X1    g1026(.A1(new_n546_), .A2(new_n547_), .ZN(new_n1412_));
  NOR4_X1    g1027(.A1(new_n539_), .A2(new_n540_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n1413_));
  NOR4_X1    g1028(.A1(new_n548_), .A2(new_n549_), .A3(new_n551_), .A4(new_n552_), .ZN(new_n1414_));
  OAI22_X1   g1029(.A1(new_n1411_), .A2(new_n1413_), .B1(new_n1414_), .B2(new_n1412_), .ZN(new_n1415_));
  NOR2_X1    g1030(.A1(new_n554_), .A2(new_n555_), .ZN(new_n1416_));
  NOR2_X1    g1031(.A1(new_n598_), .A2(new_n599_), .ZN(new_n1417_));
  NOR4_X1    g1032(.A1(new_n556_), .A2(new_n557_), .A3(new_n595_), .A4(new_n596_), .ZN(new_n1418_));
  NOR4_X1    g1033(.A1(new_n600_), .A2(new_n601_), .A3(new_n603_), .A4(new_n604_), .ZN(new_n1419_));
  OAI22_X1   g1034(.A1(new_n1416_), .A2(new_n1418_), .B1(new_n1419_), .B2(new_n1417_), .ZN(new_n1420_));
  NOR3_X1    g1035(.A1(new_n1415_), .A2(new_n1420_), .A3(new_n1410_), .ZN(new_n1421_));
  NOR2_X1    g1036(.A1(new_n572_), .A2(new_n573_), .ZN(new_n1422_));
  NOR2_X1    g1037(.A1(new_n581_), .A2(new_n582_), .ZN(new_n1423_));
  NOR4_X1    g1038(.A1(new_n574_), .A2(new_n575_), .A3(new_n578_), .A4(new_n579_), .ZN(new_n1424_));
  NOR4_X1    g1039(.A1(new_n583_), .A2(new_n584_), .A3(new_n586_), .A4(new_n587_), .ZN(new_n1425_));
  OAI22_X1   g1040(.A1(new_n1422_), .A2(new_n1424_), .B1(new_n1425_), .B2(new_n1423_), .ZN(new_n1426_));
  NOR2_X1    g1041(.A1(new_n424_), .A2(new_n425_), .ZN(new_n1427_));
  NOR2_X1    g1042(.A1(new_n589_), .A2(new_n590_), .ZN(new_n1428_));
  NOR4_X1    g1043(.A1(new_n421_), .A2(new_n422_), .A3(new_n591_), .A4(new_n592_), .ZN(new_n1429_));
  NOR4_X1    g1044(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .A4(new_n430_), .ZN(new_n1430_));
  OAI22_X1   g1045(.A1(new_n1427_), .A2(new_n1430_), .B1(new_n1429_), .B2(new_n1428_), .ZN(new_n1431_));
  NOR2_X1    g1046(.A1(new_n606_), .A2(new_n607_), .ZN(new_n1432_));
  NOR2_X1    g1047(.A1(new_n615_), .A2(new_n616_), .ZN(new_n1433_));
  NOR4_X1    g1048(.A1(new_n608_), .A2(new_n609_), .A3(new_n612_), .A4(new_n613_), .ZN(new_n1434_));
  NOR4_X1    g1049(.A1(new_n617_), .A2(new_n618_), .A3(new_n620_), .A4(new_n621_), .ZN(new_n1435_));
  OAI22_X1   g1050(.A1(new_n1432_), .A2(new_n1434_), .B1(new_n1435_), .B2(new_n1433_), .ZN(new_n1436_));
  NOR2_X1    g1051(.A1(new_n564_), .A2(new_n565_), .ZN(new_n1437_));
  NOR2_X1    g1052(.A1(new_n623_), .A2(new_n624_), .ZN(new_n1438_));
  NOR4_X1    g1053(.A1(new_n561_), .A2(new_n562_), .A3(new_n625_), .A4(new_n626_), .ZN(new_n1439_));
  NOR4_X1    g1054(.A1(new_n566_), .A2(new_n567_), .A3(new_n569_), .A4(new_n570_), .ZN(new_n1440_));
  OAI22_X1   g1055(.A1(new_n1437_), .A2(new_n1440_), .B1(new_n1439_), .B2(new_n1438_), .ZN(new_n1441_));
  NOR4_X1    g1056(.A1(new_n1426_), .A2(new_n1431_), .A3(new_n1436_), .A4(new_n1441_), .ZN(new_n1442_));
  NAND4_X1   g1057(.A1(new_n1387_), .A2(new_n1442_), .A3(new_n1406_), .A4(new_n1421_), .ZN(new_n1443_));
  AOI21_X1   g1058(.A1(new_n1443_), .A2(new_n1330_), .B(new_n767_), .ZN(\grant[6] ));
  NOR2_X1    g1059(.A1(new_n644_), .A2(new_n645_), .ZN(new_n1445_));
  NOR2_X1    g1060(.A1(new_n653_), .A2(new_n654_), .ZN(new_n1446_));
  NOR4_X1    g1061(.A1(new_n646_), .A2(new_n647_), .A3(new_n650_), .A4(new_n651_), .ZN(new_n1447_));
  NOR4_X1    g1062(.A1(new_n655_), .A2(new_n656_), .A3(new_n658_), .A4(new_n659_), .ZN(new_n1448_));
  OAI22_X1   g1063(.A1(new_n1445_), .A2(new_n1447_), .B1(new_n1448_), .B2(new_n1446_), .ZN(new_n1449_));
  NOR2_X1    g1064(.A1(new_n661_), .A2(new_n662_), .ZN(new_n1450_));
  NOR2_X1    g1065(.A1(new_n731_), .A2(new_n732_), .ZN(new_n1451_));
  NOR4_X1    g1066(.A1(new_n663_), .A2(new_n664_), .A3(new_n728_), .A4(new_n729_), .ZN(new_n1452_));
  NOR4_X1    g1067(.A1(new_n733_), .A2(new_n734_), .A3(new_n736_), .A4(new_n737_), .ZN(new_n1453_));
  OAI22_X1   g1068(.A1(new_n1450_), .A2(new_n1452_), .B1(new_n1453_), .B2(new_n1451_), .ZN(new_n1454_));
  NOR2_X1    g1069(.A1(new_n678_), .A2(new_n679_), .ZN(new_n1455_));
  NOR2_X1    g1070(.A1(new_n687_), .A2(new_n688_), .ZN(new_n1456_));
  NOR4_X1    g1071(.A1(new_n680_), .A2(new_n681_), .A3(new_n684_), .A4(new_n685_), .ZN(new_n1457_));
  NOR4_X1    g1072(.A1(new_n689_), .A2(new_n690_), .A3(new_n692_), .A4(new_n693_), .ZN(new_n1458_));
  OAI22_X1   g1073(.A1(new_n1455_), .A2(new_n1457_), .B1(new_n1458_), .B2(new_n1456_), .ZN(new_n1459_));
  NOR2_X1    g1074(.A1(new_n636_), .A2(new_n637_), .ZN(new_n1460_));
  NOR2_X1    g1075(.A1(new_n695_), .A2(new_n696_), .ZN(new_n1461_));
  NOR4_X1    g1076(.A1(new_n633_), .A2(new_n634_), .A3(new_n697_), .A4(new_n698_), .ZN(new_n1462_));
  NOR4_X1    g1077(.A1(new_n638_), .A2(new_n639_), .A3(new_n641_), .A4(new_n642_), .ZN(new_n1463_));
  OAI22_X1   g1078(.A1(new_n1460_), .A2(new_n1463_), .B1(new_n1462_), .B2(new_n1461_), .ZN(new_n1464_));
  NOR4_X1    g1079(.A1(new_n1449_), .A2(new_n1454_), .A3(new_n1459_), .A4(new_n1464_), .ZN(new_n1465_));
  NOR2_X1    g1080(.A1(new_n1230_), .A2(new_n1231_), .ZN(new_n1466_));
  NOR4_X1    g1081(.A1(new_n1009_), .A2(new_n1010_), .A3(new_n1011_), .A4(new_n1287_), .ZN(new_n1467_));
  NOR2_X1    g1082(.A1(new_n1467_), .A2(new_n1466_), .ZN(new_n1468_));
  NOR2_X1    g1083(.A1(new_n705_), .A2(new_n706_), .ZN(new_n1469_));
  NOR2_X1    g1084(.A1(new_n722_), .A2(new_n723_), .ZN(new_n1470_));
  NOR4_X1    g1085(.A1(new_n702_), .A2(new_n703_), .A3(new_n724_), .A4(new_n725_), .ZN(new_n1471_));
  NOR4_X1    g1086(.A1(new_n707_), .A2(new_n708_), .A3(new_n1229_), .A4(new_n877_), .ZN(new_n1472_));
  OAI22_X1   g1087(.A1(new_n1469_), .A2(new_n1472_), .B1(new_n1471_), .B2(new_n1470_), .ZN(new_n1473_));
  NOR2_X1    g1088(.A1(new_n739_), .A2(new_n740_), .ZN(new_n1474_));
  NOR2_X1    g1089(.A1(new_n748_), .A2(new_n749_), .ZN(new_n1475_));
  NOR4_X1    g1090(.A1(new_n741_), .A2(new_n742_), .A3(new_n745_), .A4(new_n746_), .ZN(new_n1476_));
  NOR4_X1    g1091(.A1(new_n750_), .A2(new_n751_), .A3(new_n753_), .A4(new_n754_), .ZN(new_n1477_));
  OAI22_X1   g1092(.A1(new_n1474_), .A2(new_n1476_), .B1(new_n1477_), .B2(new_n1475_), .ZN(new_n1478_));
  NOR2_X1    g1093(.A1(new_n714_), .A2(new_n715_), .ZN(new_n1479_));
  NOR2_X1    g1094(.A1(new_n756_), .A2(new_n757_), .ZN(new_n1480_));
  NOR4_X1    g1095(.A1(new_n711_), .A2(new_n712_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n1481_));
  NOR4_X1    g1096(.A1(new_n716_), .A2(new_n717_), .A3(new_n719_), .A4(new_n720_), .ZN(new_n1482_));
  OAI22_X1   g1097(.A1(new_n1479_), .A2(new_n1482_), .B1(new_n1481_), .B2(new_n1480_), .ZN(new_n1483_));
  NOR4_X1    g1098(.A1(new_n1473_), .A2(new_n1478_), .A3(new_n1483_), .A4(new_n1468_), .ZN(new_n1484_));
  NOR4_X1    g1099(.A1(new_n777_), .A2(new_n778_), .A3(new_n780_), .A4(new_n781_), .ZN(new_n1485_));
  INV_X1     g1100(.I(\req[8] ), .ZN(new_n1486_));
  AOI21_X1   g1101(.A1(new_n1486_), .A2(\priority[8] ), .B(\priority[9] ), .ZN(new_n1487_));
  OAI21_X1   g1102(.A1(new_n1485_), .A2(new_n775_), .B(new_n1487_), .ZN(new_n1488_));
  NOR2_X1    g1103(.A1(new_n783_), .A2(new_n784_), .ZN(new_n1489_));
  NOR2_X1    g1104(.A1(new_n792_), .A2(new_n793_), .ZN(new_n1490_));
  NOR4_X1    g1105(.A1(new_n785_), .A2(new_n786_), .A3(new_n789_), .A4(new_n790_), .ZN(new_n1491_));
  NOR4_X1    g1106(.A1(new_n794_), .A2(new_n795_), .A3(new_n797_), .A4(new_n798_), .ZN(new_n1492_));
  OAI22_X1   g1107(.A1(new_n1489_), .A2(new_n1491_), .B1(new_n1492_), .B2(new_n1490_), .ZN(new_n1493_));
  NOR2_X1    g1108(.A1(new_n800_), .A2(new_n801_), .ZN(new_n1494_));
  NOR2_X1    g1109(.A1(new_n844_), .A2(new_n845_), .ZN(new_n1495_));
  NOR4_X1    g1110(.A1(new_n802_), .A2(new_n803_), .A3(new_n841_), .A4(new_n842_), .ZN(new_n1496_));
  NOR4_X1    g1111(.A1(new_n846_), .A2(new_n847_), .A3(new_n849_), .A4(new_n850_), .ZN(new_n1497_));
  OAI22_X1   g1112(.A1(new_n1494_), .A2(new_n1496_), .B1(new_n1497_), .B2(new_n1495_), .ZN(new_n1498_));
  NOR3_X1    g1113(.A1(new_n1493_), .A2(new_n1498_), .A3(new_n1488_), .ZN(new_n1499_));
  NOR2_X1    g1114(.A1(new_n818_), .A2(new_n819_), .ZN(new_n1500_));
  NOR2_X1    g1115(.A1(new_n827_), .A2(new_n828_), .ZN(new_n1501_));
  NOR4_X1    g1116(.A1(new_n820_), .A2(new_n821_), .A3(new_n824_), .A4(new_n825_), .ZN(new_n1502_));
  NOR4_X1    g1117(.A1(new_n829_), .A2(new_n830_), .A3(new_n832_), .A4(new_n833_), .ZN(new_n1503_));
  OAI22_X1   g1118(.A1(new_n1500_), .A2(new_n1502_), .B1(new_n1503_), .B2(new_n1501_), .ZN(new_n1504_));
  NOR2_X1    g1119(.A1(new_n670_), .A2(new_n671_), .ZN(new_n1505_));
  NOR2_X1    g1120(.A1(new_n835_), .A2(new_n836_), .ZN(new_n1506_));
  NOR4_X1    g1121(.A1(new_n667_), .A2(new_n668_), .A3(new_n837_), .A4(new_n838_), .ZN(new_n1507_));
  NOR4_X1    g1122(.A1(new_n672_), .A2(new_n673_), .A3(new_n675_), .A4(new_n676_), .ZN(new_n1508_));
  OAI22_X1   g1123(.A1(new_n1505_), .A2(new_n1508_), .B1(new_n1507_), .B2(new_n1506_), .ZN(new_n1509_));
  NOR2_X1    g1124(.A1(new_n852_), .A2(new_n853_), .ZN(new_n1510_));
  NOR2_X1    g1125(.A1(new_n861_), .A2(new_n862_), .ZN(new_n1511_));
  NOR4_X1    g1126(.A1(new_n854_), .A2(new_n855_), .A3(new_n858_), .A4(new_n859_), .ZN(new_n1512_));
  NOR4_X1    g1127(.A1(new_n863_), .A2(new_n864_), .A3(new_n866_), .A4(new_n867_), .ZN(new_n1513_));
  OAI22_X1   g1128(.A1(new_n1510_), .A2(new_n1512_), .B1(new_n1513_), .B2(new_n1511_), .ZN(new_n1514_));
  NOR2_X1    g1129(.A1(new_n810_), .A2(new_n811_), .ZN(new_n1515_));
  NOR2_X1    g1130(.A1(new_n869_), .A2(new_n870_), .ZN(new_n1516_));
  NOR4_X1    g1131(.A1(new_n807_), .A2(new_n808_), .A3(new_n871_), .A4(new_n872_), .ZN(new_n1517_));
  NOR4_X1    g1132(.A1(new_n812_), .A2(new_n813_), .A3(new_n815_), .A4(new_n816_), .ZN(new_n1518_));
  OAI22_X1   g1133(.A1(new_n1515_), .A2(new_n1518_), .B1(new_n1517_), .B2(new_n1516_), .ZN(new_n1519_));
  NOR4_X1    g1134(.A1(new_n1504_), .A2(new_n1509_), .A3(new_n1514_), .A4(new_n1519_), .ZN(new_n1520_));
  NAND4_X1   g1135(.A1(new_n1465_), .A2(new_n1520_), .A3(new_n1484_), .A4(new_n1499_), .ZN(new_n1521_));
  AOI21_X1   g1136(.A1(new_n1521_), .A2(new_n1408_), .B(new_n1013_), .ZN(\grant[7] ));
  NOR2_X1    g1137(.A1(new_n890_), .A2(new_n891_), .ZN(new_n1523_));
  NOR2_X1    g1138(.A1(new_n899_), .A2(new_n900_), .ZN(new_n1524_));
  NOR4_X1    g1139(.A1(new_n892_), .A2(new_n893_), .A3(new_n896_), .A4(new_n897_), .ZN(new_n1525_));
  NOR4_X1    g1140(.A1(new_n901_), .A2(new_n902_), .A3(new_n904_), .A4(new_n905_), .ZN(new_n1526_));
  OAI22_X1   g1141(.A1(new_n1523_), .A2(new_n1525_), .B1(new_n1526_), .B2(new_n1524_), .ZN(new_n1527_));
  NOR2_X1    g1142(.A1(new_n907_), .A2(new_n908_), .ZN(new_n1528_));
  NOR2_X1    g1143(.A1(new_n977_), .A2(new_n978_), .ZN(new_n1529_));
  NOR4_X1    g1144(.A1(new_n909_), .A2(new_n910_), .A3(new_n974_), .A4(new_n975_), .ZN(new_n1530_));
  NOR4_X1    g1145(.A1(new_n979_), .A2(new_n980_), .A3(new_n982_), .A4(new_n983_), .ZN(new_n1531_));
  OAI22_X1   g1146(.A1(new_n1528_), .A2(new_n1530_), .B1(new_n1531_), .B2(new_n1529_), .ZN(new_n1532_));
  NOR2_X1    g1147(.A1(new_n924_), .A2(new_n925_), .ZN(new_n1533_));
  NOR2_X1    g1148(.A1(new_n933_), .A2(new_n934_), .ZN(new_n1534_));
  NOR4_X1    g1149(.A1(new_n926_), .A2(new_n927_), .A3(new_n930_), .A4(new_n931_), .ZN(new_n1535_));
  NOR4_X1    g1150(.A1(new_n935_), .A2(new_n936_), .A3(new_n938_), .A4(new_n939_), .ZN(new_n1536_));
  OAI22_X1   g1151(.A1(new_n1533_), .A2(new_n1535_), .B1(new_n1536_), .B2(new_n1534_), .ZN(new_n1537_));
  NOR2_X1    g1152(.A1(new_n882_), .A2(new_n883_), .ZN(new_n1538_));
  NOR2_X1    g1153(.A1(new_n941_), .A2(new_n942_), .ZN(new_n1539_));
  NOR4_X1    g1154(.A1(new_n879_), .A2(new_n880_), .A3(new_n943_), .A4(new_n944_), .ZN(new_n1540_));
  NOR4_X1    g1155(.A1(new_n884_), .A2(new_n885_), .A3(new_n887_), .A4(new_n888_), .ZN(new_n1541_));
  OAI22_X1   g1156(.A1(new_n1538_), .A2(new_n1541_), .B1(new_n1540_), .B2(new_n1539_), .ZN(new_n1542_));
  NOR4_X1    g1157(.A1(new_n1527_), .A2(new_n1532_), .A3(new_n1537_), .A4(new_n1542_), .ZN(new_n1543_));
  NOR2_X1    g1158(.A1(new_n518_), .A2(new_n519_), .ZN(new_n1544_));
  NOR4_X1    g1159(.A1(new_n520_), .A2(new_n521_), .A3(new_n526_), .A4(new_n527_), .ZN(new_n1545_));
  NOR2_X1    g1160(.A1(new_n1545_), .A2(new_n1544_), .ZN(new_n1546_));
  NOR2_X1    g1161(.A1(new_n951_), .A2(new_n952_), .ZN(new_n1547_));
  NOR2_X1    g1162(.A1(new_n968_), .A2(new_n969_), .ZN(new_n1548_));
  NOR4_X1    g1163(.A1(new_n948_), .A2(new_n949_), .A3(new_n970_), .A4(new_n971_), .ZN(new_n1549_));
  NOR4_X1    g1164(.A1(new_n517_), .A2(new_n953_), .A3(new_n954_), .A4(new_n1123_), .ZN(new_n1550_));
  OAI22_X1   g1165(.A1(new_n1547_), .A2(new_n1550_), .B1(new_n1549_), .B2(new_n1548_), .ZN(new_n1551_));
  NOR2_X1    g1166(.A1(new_n985_), .A2(new_n986_), .ZN(new_n1552_));
  NOR2_X1    g1167(.A1(new_n994_), .A2(new_n995_), .ZN(new_n1553_));
  NOR4_X1    g1168(.A1(new_n987_), .A2(new_n988_), .A3(new_n991_), .A4(new_n992_), .ZN(new_n1554_));
  NOR4_X1    g1169(.A1(new_n996_), .A2(new_n997_), .A3(new_n999_), .A4(new_n1000_), .ZN(new_n1555_));
  OAI22_X1   g1170(.A1(new_n1552_), .A2(new_n1554_), .B1(new_n1555_), .B2(new_n1553_), .ZN(new_n1556_));
  NOR2_X1    g1171(.A1(new_n960_), .A2(new_n961_), .ZN(new_n1557_));
  NOR2_X1    g1172(.A1(new_n1002_), .A2(new_n1003_), .ZN(new_n1558_));
  NOR4_X1    g1173(.A1(new_n957_), .A2(new_n958_), .A3(new_n1004_), .A4(new_n1005_), .ZN(new_n1559_));
  NOR4_X1    g1174(.A1(new_n962_), .A2(new_n963_), .A3(new_n965_), .A4(new_n966_), .ZN(new_n1560_));
  OAI22_X1   g1175(.A1(new_n1557_), .A2(new_n1560_), .B1(new_n1559_), .B2(new_n1558_), .ZN(new_n1561_));
  NOR4_X1    g1176(.A1(new_n1551_), .A2(new_n1556_), .A3(new_n1561_), .A4(new_n1546_), .ZN(new_n1562_));
  NOR4_X1    g1177(.A1(new_n1023_), .A2(new_n1024_), .A3(new_n1026_), .A4(new_n1027_), .ZN(new_n1563_));
  INV_X1     g1178(.I(\req[9] ), .ZN(new_n1564_));
  AOI21_X1   g1179(.A1(new_n1564_), .A2(\priority[9] ), .B(\priority[10] ), .ZN(new_n1565_));
  OAI21_X1   g1180(.A1(new_n1563_), .A2(new_n1021_), .B(new_n1565_), .ZN(new_n1566_));
  NOR2_X1    g1181(.A1(new_n1029_), .A2(new_n1030_), .ZN(new_n1567_));
  NOR2_X1    g1182(.A1(new_n1038_), .A2(new_n1039_), .ZN(new_n1568_));
  NOR4_X1    g1183(.A1(new_n1031_), .A2(new_n1032_), .A3(new_n1035_), .A4(new_n1036_), .ZN(new_n1569_));
  NOR4_X1    g1184(.A1(new_n1040_), .A2(new_n1041_), .A3(new_n1043_), .A4(new_n1044_), .ZN(new_n1570_));
  OAI22_X1   g1185(.A1(new_n1567_), .A2(new_n1569_), .B1(new_n1570_), .B2(new_n1568_), .ZN(new_n1571_));
  NOR2_X1    g1186(.A1(new_n1046_), .A2(new_n1047_), .ZN(new_n1572_));
  NOR2_X1    g1187(.A1(new_n1090_), .A2(new_n1091_), .ZN(new_n1573_));
  NOR4_X1    g1188(.A1(new_n1048_), .A2(new_n1049_), .A3(new_n1087_), .A4(new_n1088_), .ZN(new_n1574_));
  NOR4_X1    g1189(.A1(new_n1092_), .A2(new_n1093_), .A3(new_n1095_), .A4(new_n1096_), .ZN(new_n1575_));
  OAI22_X1   g1190(.A1(new_n1572_), .A2(new_n1574_), .B1(new_n1575_), .B2(new_n1573_), .ZN(new_n1576_));
  NOR3_X1    g1191(.A1(new_n1571_), .A2(new_n1576_), .A3(new_n1566_), .ZN(new_n1577_));
  NOR2_X1    g1192(.A1(new_n1064_), .A2(new_n1065_), .ZN(new_n1578_));
  NOR2_X1    g1193(.A1(new_n1073_), .A2(new_n1074_), .ZN(new_n1579_));
  NOR4_X1    g1194(.A1(new_n1066_), .A2(new_n1067_), .A3(new_n1070_), .A4(new_n1071_), .ZN(new_n1580_));
  NOR4_X1    g1195(.A1(new_n1075_), .A2(new_n1076_), .A3(new_n1078_), .A4(new_n1079_), .ZN(new_n1581_));
  OAI22_X1   g1196(.A1(new_n1578_), .A2(new_n1580_), .B1(new_n1581_), .B2(new_n1579_), .ZN(new_n1582_));
  NOR2_X1    g1197(.A1(new_n916_), .A2(new_n917_), .ZN(new_n1583_));
  NOR2_X1    g1198(.A1(new_n1081_), .A2(new_n1082_), .ZN(new_n1584_));
  NOR4_X1    g1199(.A1(new_n913_), .A2(new_n914_), .A3(new_n1083_), .A4(new_n1084_), .ZN(new_n1585_));
  NOR4_X1    g1200(.A1(new_n918_), .A2(new_n919_), .A3(new_n921_), .A4(new_n922_), .ZN(new_n1586_));
  OAI22_X1   g1201(.A1(new_n1583_), .A2(new_n1586_), .B1(new_n1585_), .B2(new_n1584_), .ZN(new_n1587_));
  NOR2_X1    g1202(.A1(new_n1098_), .A2(new_n1099_), .ZN(new_n1588_));
  NOR2_X1    g1203(.A1(new_n1107_), .A2(new_n1108_), .ZN(new_n1589_));
  NOR4_X1    g1204(.A1(new_n1100_), .A2(new_n1101_), .A3(new_n1104_), .A4(new_n1105_), .ZN(new_n1590_));
  NOR4_X1    g1205(.A1(new_n1109_), .A2(new_n1110_), .A3(new_n1112_), .A4(new_n1113_), .ZN(new_n1591_));
  OAI22_X1   g1206(.A1(new_n1588_), .A2(new_n1590_), .B1(new_n1591_), .B2(new_n1589_), .ZN(new_n1592_));
  NOR2_X1    g1207(.A1(new_n1056_), .A2(new_n1057_), .ZN(new_n1593_));
  NOR2_X1    g1208(.A1(new_n1115_), .A2(new_n1116_), .ZN(new_n1594_));
  NOR4_X1    g1209(.A1(new_n1053_), .A2(new_n1054_), .A3(new_n1117_), .A4(new_n1118_), .ZN(new_n1595_));
  NOR4_X1    g1210(.A1(new_n1058_), .A2(new_n1059_), .A3(new_n1061_), .A4(new_n1062_), .ZN(new_n1596_));
  OAI22_X1   g1211(.A1(new_n1593_), .A2(new_n1596_), .B1(new_n1595_), .B2(new_n1594_), .ZN(new_n1597_));
  NOR4_X1    g1212(.A1(new_n1582_), .A2(new_n1587_), .A3(new_n1592_), .A4(new_n1597_), .ZN(new_n1598_));
  NAND4_X1   g1213(.A1(new_n1543_), .A2(new_n1598_), .A3(new_n1562_), .A4(new_n1577_), .ZN(new_n1599_));
  AOI21_X1   g1214(.A1(new_n1599_), .A2(new_n1486_), .B(new_n530_), .ZN(\grant[8] ));
  OAI22_X1   g1215(.A1(new_n414_), .A2(new_n419_), .B1(new_n489_), .B2(new_n484_), .ZN(new_n1601_));
  OAI22_X1   g1216(.A1(new_n492_), .A2(new_n497_), .B1(new_n506_), .B2(new_n501_), .ZN(new_n1602_));
  OAI22_X1   g1217(.A1(new_n389_), .A2(new_n394_), .B1(new_n453_), .B2(new_n448_), .ZN(new_n1603_));
  OAI22_X1   g1218(.A1(new_n397_), .A2(new_n402_), .B1(new_n411_), .B2(new_n406_), .ZN(new_n1604_));
  NOR4_X1    g1219(.A1(new_n1601_), .A2(new_n1602_), .A3(new_n1603_), .A4(new_n1604_), .ZN(new_n1605_));
  NOR2_X1    g1220(.A1(new_n764_), .A2(new_n765_), .ZN(new_n1606_));
  NOR4_X1    g1221(.A1(new_n766_), .A2(new_n767_), .A3(new_n772_), .A4(new_n773_), .ZN(new_n1607_));
  NOR2_X1    g1222(.A1(new_n1607_), .A2(new_n1606_), .ZN(new_n1608_));
  NOR2_X1    g1223(.A1(new_n1147_), .A2(new_n631_), .ZN(new_n1609_));
  NOR4_X1    g1224(.A1(new_n763_), .A2(new_n1148_), .A3(new_n1149_), .A4(new_n1205_), .ZN(new_n1610_));
  OAI22_X1   g1225(.A1(new_n534_), .A2(new_n541_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n1611_));
  OAI22_X1   g1226(.A1(new_n467_), .A2(new_n472_), .B1(new_n514_), .B2(new_n509_), .ZN(new_n1612_));
  OAI22_X1   g1227(.A1(new_n458_), .A2(new_n463_), .B1(new_n480_), .B2(new_n475_), .ZN(new_n1613_));
  NOR4_X1    g1228(.A1(new_n1611_), .A2(new_n1612_), .A3(new_n1613_), .A4(new_n1608_), .ZN(new_n1614_));
  INV_X1     g1229(.I(\req[10] ), .ZN(new_n1615_));
  AOI21_X1   g1230(.A1(new_n1615_), .A2(\priority[10] ), .B(\priority[11] ), .ZN(new_n1616_));
  OAI21_X1   g1231(.A1(new_n550_), .A2(new_n545_), .B(new_n1616_), .ZN(new_n1617_));
  OAI22_X1   g1232(.A1(new_n553_), .A2(new_n558_), .B1(new_n602_), .B2(new_n597_), .ZN(new_n1618_));
  OAI22_X1   g1233(.A1(new_n605_), .A2(new_n610_), .B1(new_n619_), .B2(new_n614_), .ZN(new_n1619_));
  NOR3_X1    g1234(.A1(new_n1618_), .A2(new_n1619_), .A3(new_n1617_), .ZN(new_n1620_));
  OAI22_X1   g1235(.A1(new_n423_), .A2(new_n428_), .B1(new_n593_), .B2(new_n588_), .ZN(new_n1621_));
  OAI22_X1   g1236(.A1(new_n431_), .A2(new_n436_), .B1(new_n445_), .B2(new_n440_), .ZN(new_n1622_));
  OAI22_X1   g1237(.A1(new_n563_), .A2(new_n568_), .B1(new_n627_), .B2(new_n622_), .ZN(new_n1623_));
  OAI22_X1   g1238(.A1(new_n571_), .A2(new_n576_), .B1(new_n585_), .B2(new_n580_), .ZN(new_n1624_));
  NOR4_X1    g1239(.A1(new_n1621_), .A2(new_n1622_), .A3(new_n1623_), .A4(new_n1624_), .ZN(new_n1625_));
  NAND4_X1   g1240(.A1(new_n1605_), .A2(new_n1625_), .A3(new_n1614_), .A4(new_n1620_), .ZN(new_n1626_));
  AOI21_X1   g1241(.A1(new_n1626_), .A2(new_n1564_), .B(new_n776_), .ZN(\grant[9] ));
  OAI22_X1   g1242(.A1(new_n660_), .A2(new_n665_), .B1(new_n735_), .B2(new_n730_), .ZN(new_n1628_));
  OAI22_X1   g1243(.A1(new_n738_), .A2(new_n743_), .B1(new_n752_), .B2(new_n747_), .ZN(new_n1629_));
  OAI22_X1   g1244(.A1(new_n635_), .A2(new_n640_), .B1(new_n699_), .B2(new_n694_), .ZN(new_n1630_));
  OAI22_X1   g1245(.A1(new_n643_), .A2(new_n648_), .B1(new_n657_), .B2(new_n652_), .ZN(new_n1631_));
  NOR4_X1    g1246(.A1(new_n1628_), .A2(new_n1629_), .A3(new_n1630_), .A4(new_n1631_), .ZN(new_n1632_));
  NOR2_X1    g1247(.A1(new_n1010_), .A2(new_n1011_), .ZN(new_n1633_));
  NOR4_X1    g1248(.A1(new_n1012_), .A2(new_n1013_), .A3(new_n1018_), .A4(new_n1019_), .ZN(new_n1634_));
  NOR2_X1    g1249(.A1(new_n1634_), .A2(new_n1633_), .ZN(new_n1635_));
  NOR2_X1    g1250(.A1(new_n1229_), .A2(new_n877_), .ZN(new_n1636_));
  NOR4_X1    g1251(.A1(new_n1009_), .A2(new_n1230_), .A3(new_n1231_), .A4(new_n1287_), .ZN(new_n1637_));
  OAI22_X1   g1252(.A1(new_n780_), .A2(new_n787_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n1638_));
  OAI22_X1   g1253(.A1(new_n713_), .A2(new_n718_), .B1(new_n760_), .B2(new_n755_), .ZN(new_n1639_));
  OAI22_X1   g1254(.A1(new_n704_), .A2(new_n709_), .B1(new_n726_), .B2(new_n721_), .ZN(new_n1640_));
  NOR4_X1    g1255(.A1(new_n1638_), .A2(new_n1639_), .A3(new_n1640_), .A4(new_n1635_), .ZN(new_n1641_));
  INV_X1     g1256(.I(\req[11] ), .ZN(new_n1642_));
  AOI21_X1   g1257(.A1(new_n1642_), .A2(\priority[11] ), .B(\priority[12] ), .ZN(new_n1643_));
  OAI21_X1   g1258(.A1(new_n796_), .A2(new_n791_), .B(new_n1643_), .ZN(new_n1644_));
  OAI22_X1   g1259(.A1(new_n799_), .A2(new_n804_), .B1(new_n848_), .B2(new_n843_), .ZN(new_n1645_));
  OAI22_X1   g1260(.A1(new_n851_), .A2(new_n856_), .B1(new_n865_), .B2(new_n860_), .ZN(new_n1646_));
  NOR3_X1    g1261(.A1(new_n1645_), .A2(new_n1646_), .A3(new_n1644_), .ZN(new_n1647_));
  OAI22_X1   g1262(.A1(new_n669_), .A2(new_n674_), .B1(new_n839_), .B2(new_n834_), .ZN(new_n1648_));
  OAI22_X1   g1263(.A1(new_n677_), .A2(new_n682_), .B1(new_n691_), .B2(new_n686_), .ZN(new_n1649_));
  OAI22_X1   g1264(.A1(new_n809_), .A2(new_n814_), .B1(new_n873_), .B2(new_n868_), .ZN(new_n1650_));
  OAI22_X1   g1265(.A1(new_n817_), .A2(new_n822_), .B1(new_n831_), .B2(new_n826_), .ZN(new_n1651_));
  NOR4_X1    g1266(.A1(new_n1648_), .A2(new_n1649_), .A3(new_n1650_), .A4(new_n1651_), .ZN(new_n1652_));
  NAND4_X1   g1267(.A1(new_n1632_), .A2(new_n1652_), .A3(new_n1641_), .A4(new_n1647_), .ZN(new_n1653_));
  AOI21_X1   g1268(.A1(new_n1653_), .A2(new_n1615_), .B(new_n1022_), .ZN(\grant[10] ));
  NOR4_X1    g1269(.A1(new_n895_), .A2(new_n912_), .A3(new_n946_), .A4(new_n990_), .ZN(new_n1655_));
  NOR2_X1    g1270(.A1(new_n517_), .A2(new_n1123_), .ZN(new_n1656_));
  NOR2_X1    g1271(.A1(new_n522_), .A2(new_n1656_), .ZN(new_n1657_));
  OAI22_X1   g1272(.A1(new_n950_), .A2(new_n955_), .B1(new_n1033_), .B2(new_n1026_), .ZN(new_n1658_));
  NOR4_X1    g1273(.A1(new_n973_), .A2(new_n1007_), .A3(new_n1658_), .A4(new_n1657_), .ZN(new_n1659_));
  INV_X1     g1274(.I(\req[12] ), .ZN(new_n1660_));
  AOI21_X1   g1275(.A1(new_n1660_), .A2(\priority[12] ), .B(\priority[13] ), .ZN(new_n1661_));
  OAI21_X1   g1276(.A1(new_n533_), .A2(new_n528_), .B(new_n1661_), .ZN(new_n1662_));
  NOR3_X1    g1277(.A1(new_n1051_), .A2(new_n1103_), .A3(new_n1662_), .ZN(new_n1663_));
  NOR4_X1    g1278(.A1(new_n929_), .A2(new_n1069_), .A3(new_n1086_), .A4(new_n1120_), .ZN(new_n1664_));
  NAND4_X1   g1279(.A1(new_n1655_), .A2(new_n1664_), .A3(new_n1659_), .A4(new_n1663_), .ZN(new_n1665_));
  AOI21_X1   g1280(.A1(new_n1665_), .A2(new_n1642_), .B(new_n535_), .ZN(\grant[11] ));
  NOR4_X1    g1281(.A1(new_n1129_), .A2(new_n1134_), .A3(new_n1144_), .A4(new_n1161_), .ZN(new_n1667_));
  NOR2_X1    g1282(.A1(new_n763_), .A2(new_n1205_), .ZN(new_n1668_));
  NOR2_X1    g1283(.A1(new_n768_), .A2(new_n1668_), .ZN(new_n1669_));
  OAI22_X1   g1284(.A1(new_n1146_), .A2(new_n1150_), .B1(new_n1175_), .B2(new_n539_), .ZN(new_n1670_));
  NOR4_X1    g1285(.A1(new_n1156_), .A2(new_n1166_), .A3(new_n1670_), .A4(new_n1669_), .ZN(new_n1671_));
  INV_X1     g1286(.I(\req[13] ), .ZN(new_n1672_));
  AOI21_X1   g1287(.A1(new_n1672_), .A2(\priority[13] ), .B(\priority[14] ), .ZN(new_n1673_));
  OAI21_X1   g1288(.A1(new_n779_), .A2(new_n774_), .B(new_n1673_), .ZN(new_n1674_));
  NOR3_X1    g1289(.A1(new_n1181_), .A2(new_n1197_), .A3(new_n1674_), .ZN(new_n1675_));
  NOR4_X1    g1290(.A1(new_n1139_), .A2(new_n1187_), .A3(new_n1192_), .A4(new_n1202_), .ZN(new_n1676_));
  NAND4_X1   g1291(.A1(new_n1667_), .A2(new_n1676_), .A3(new_n1671_), .A4(new_n1675_), .ZN(new_n1677_));
  AOI21_X1   g1292(.A1(new_n1677_), .A2(new_n1660_), .B(new_n781_), .ZN(\grant[12] ));
  NOR4_X1    g1293(.A1(new_n1211_), .A2(new_n1216_), .A3(new_n1226_), .A4(new_n1243_), .ZN(new_n1679_));
  NOR2_X1    g1294(.A1(new_n1009_), .A2(new_n1287_), .ZN(new_n1680_));
  NOR2_X1    g1295(.A1(new_n1014_), .A2(new_n1680_), .ZN(new_n1681_));
  OAI22_X1   g1296(.A1(new_n1228_), .A2(new_n1232_), .B1(new_n1257_), .B2(new_n785_), .ZN(new_n1682_));
  NOR4_X1    g1297(.A1(new_n1238_), .A2(new_n1248_), .A3(new_n1682_), .A4(new_n1681_), .ZN(new_n1683_));
  INV_X1     g1298(.I(\req[14] ), .ZN(new_n1684_));
  AOI21_X1   g1299(.A1(new_n1684_), .A2(\priority[14] ), .B(\priority[15] ), .ZN(new_n1685_));
  OAI21_X1   g1300(.A1(new_n1025_), .A2(new_n1020_), .B(new_n1685_), .ZN(new_n1686_));
  NOR3_X1    g1301(.A1(new_n1263_), .A2(new_n1279_), .A3(new_n1686_), .ZN(new_n1687_));
  NOR4_X1    g1302(.A1(new_n1221_), .A2(new_n1269_), .A3(new_n1274_), .A4(new_n1284_), .ZN(new_n1688_));
  NAND4_X1   g1303(.A1(new_n1679_), .A2(new_n1688_), .A3(new_n1683_), .A4(new_n1687_), .ZN(new_n1689_));
  AOI21_X1   g1304(.A1(new_n1689_), .A2(new_n1672_), .B(new_n1027_), .ZN(\grant[13] ));
  NOR4_X1    g1305(.A1(new_n1293_), .A2(new_n1298_), .A3(new_n1308_), .A4(new_n1322_), .ZN(new_n1691_));
  NOR2_X1    g1306(.A1(new_n520_), .A2(new_n521_), .ZN(new_n1692_));
  NOR2_X1    g1307(.A1(new_n1168_), .A2(new_n1692_), .ZN(new_n1693_));
  OAI22_X1   g1308(.A1(new_n1310_), .A2(new_n1311_), .B1(new_n1336_), .B2(new_n1031_), .ZN(new_n1694_));
  NOR4_X1    g1309(.A1(new_n1317_), .A2(new_n1327_), .A3(new_n1694_), .A4(new_n1693_), .ZN(new_n1695_));
  INV_X1     g1310(.I(\req[15] ), .ZN(new_n1696_));
  AOI21_X1   g1311(.A1(new_n1696_), .A2(\priority[15] ), .B(\priority[16] ), .ZN(new_n1697_));
  OAI21_X1   g1312(.A1(new_n1174_), .A2(new_n1172_), .B(new_n1697_), .ZN(new_n1698_));
  NOR3_X1    g1313(.A1(new_n1342_), .A2(new_n1358_), .A3(new_n1698_), .ZN(new_n1699_));
  NOR4_X1    g1314(.A1(new_n1303_), .A2(new_n1348_), .A3(new_n1353_), .A4(new_n1363_), .ZN(new_n1700_));
  NAND4_X1   g1315(.A1(new_n1691_), .A2(new_n1700_), .A3(new_n1695_), .A4(new_n1699_), .ZN(new_n1701_));
  AOI21_X1   g1316(.A1(new_n1701_), .A2(new_n1684_), .B(new_n540_), .ZN(\grant[14] ));
  NOR4_X1    g1317(.A1(new_n1371_), .A2(new_n1376_), .A3(new_n1386_), .A4(new_n1400_), .ZN(new_n1703_));
  NOR2_X1    g1318(.A1(new_n766_), .A2(new_n767_), .ZN(new_n1704_));
  NOR2_X1    g1319(.A1(new_n1250_), .A2(new_n1704_), .ZN(new_n1705_));
  OAI22_X1   g1320(.A1(new_n546_), .A2(new_n1414_), .B1(new_n1389_), .B2(new_n1388_), .ZN(new_n1706_));
  NOR4_X1    g1321(.A1(new_n1395_), .A2(new_n1405_), .A3(new_n1706_), .A4(new_n1705_), .ZN(new_n1707_));
  INV_X1     g1322(.I(\req[16] ), .ZN(new_n1708_));
  AOI21_X1   g1323(.A1(new_n1708_), .A2(\priority[16] ), .B(\priority[17] ), .ZN(new_n1709_));
  OAI21_X1   g1324(.A1(new_n1256_), .A2(new_n1254_), .B(new_n1709_), .ZN(new_n1710_));
  NOR3_X1    g1325(.A1(new_n1420_), .A2(new_n1436_), .A3(new_n1710_), .ZN(new_n1711_));
  NOR4_X1    g1326(.A1(new_n1381_), .A2(new_n1426_), .A3(new_n1431_), .A4(new_n1441_), .ZN(new_n1712_));
  NAND4_X1   g1327(.A1(new_n1703_), .A2(new_n1712_), .A3(new_n1707_), .A4(new_n1711_), .ZN(new_n1713_));
  AOI21_X1   g1328(.A1(new_n1713_), .A2(new_n1696_), .B(new_n786_), .ZN(\grant[15] ));
  NOR4_X1    g1329(.A1(new_n1449_), .A2(new_n1454_), .A3(new_n1464_), .A4(new_n1478_), .ZN(new_n1715_));
  NOR2_X1    g1330(.A1(new_n1012_), .A2(new_n1013_), .ZN(new_n1716_));
  NOR2_X1    g1331(.A1(new_n1329_), .A2(new_n1716_), .ZN(new_n1717_));
  OAI22_X1   g1332(.A1(new_n792_), .A2(new_n1492_), .B1(new_n1467_), .B2(new_n1466_), .ZN(new_n1718_));
  NOR4_X1    g1333(.A1(new_n1473_), .A2(new_n1483_), .A3(new_n1718_), .A4(new_n1717_), .ZN(new_n1719_));
  INV_X1     g1334(.I(\req[17] ), .ZN(new_n1720_));
  AOI21_X1   g1335(.A1(new_n1720_), .A2(\priority[17] ), .B(\priority[18] ), .ZN(new_n1721_));
  OAI21_X1   g1336(.A1(new_n1335_), .A2(new_n1333_), .B(new_n1721_), .ZN(new_n1722_));
  NOR3_X1    g1337(.A1(new_n1498_), .A2(new_n1514_), .A3(new_n1722_), .ZN(new_n1723_));
  NOR4_X1    g1338(.A1(new_n1459_), .A2(new_n1504_), .A3(new_n1509_), .A4(new_n1519_), .ZN(new_n1724_));
  NAND4_X1   g1339(.A1(new_n1715_), .A2(new_n1724_), .A3(new_n1719_), .A4(new_n1723_), .ZN(new_n1725_));
  AOI21_X1   g1340(.A1(new_n1725_), .A2(new_n1708_), .B(new_n1032_), .ZN(\grant[16] ));
  NOR4_X1    g1341(.A1(new_n1527_), .A2(new_n1532_), .A3(new_n1542_), .A4(new_n1556_), .ZN(new_n1727_));
  NOR2_X1    g1342(.A1(new_n529_), .A2(new_n530_), .ZN(new_n1728_));
  NOR2_X1    g1343(.A1(new_n1407_), .A2(new_n1728_), .ZN(new_n1729_));
  OAI22_X1   g1344(.A1(new_n1544_), .A2(new_n1545_), .B1(new_n1570_), .B2(new_n1038_), .ZN(new_n1730_));
  NOR4_X1    g1345(.A1(new_n1551_), .A2(new_n1561_), .A3(new_n1730_), .A4(new_n1729_), .ZN(new_n1731_));
  INV_X1     g1346(.I(\req[18] ), .ZN(new_n1732_));
  AOI21_X1   g1347(.A1(new_n1732_), .A2(\priority[18] ), .B(\priority[19] ), .ZN(new_n1733_));
  OAI21_X1   g1348(.A1(new_n1413_), .A2(new_n1411_), .B(new_n1733_), .ZN(new_n1734_));
  NOR3_X1    g1349(.A1(new_n1576_), .A2(new_n1592_), .A3(new_n1734_), .ZN(new_n1735_));
  NOR4_X1    g1350(.A1(new_n1537_), .A2(new_n1582_), .A3(new_n1587_), .A4(new_n1597_), .ZN(new_n1736_));
  NAND4_X1   g1351(.A1(new_n1727_), .A2(new_n1736_), .A3(new_n1731_), .A4(new_n1735_), .ZN(new_n1737_));
  AOI21_X1   g1352(.A1(new_n1737_), .A2(new_n1720_), .B(new_n547_), .ZN(\grant[17] ));
  NOR4_X1    g1353(.A1(new_n1601_), .A2(new_n1602_), .A3(new_n1604_), .A4(new_n1612_), .ZN(new_n1739_));
  NOR2_X1    g1354(.A1(new_n775_), .A2(new_n776_), .ZN(new_n1740_));
  NOR2_X1    g1355(.A1(new_n1485_), .A2(new_n1740_), .ZN(new_n1741_));
  OAI22_X1   g1356(.A1(new_n551_), .A2(new_n558_), .B1(new_n1607_), .B2(new_n1606_), .ZN(new_n1742_));
  OAI22_X1   g1357(.A1(new_n1489_), .A2(new_n1491_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n1743_));
  NOR4_X1    g1358(.A1(new_n1613_), .A2(new_n1742_), .A3(new_n1743_), .A4(new_n1741_), .ZN(new_n1744_));
  INV_X1     g1359(.I(\req[19] ), .ZN(new_n1745_));
  AOI21_X1   g1360(.A1(new_n1745_), .A2(\priority[19] ), .B(\priority[20] ), .ZN(new_n1746_));
  OAI21_X1   g1361(.A1(new_n602_), .A2(new_n597_), .B(new_n1746_), .ZN(new_n1747_));
  NOR3_X1    g1362(.A1(new_n1619_), .A2(new_n1623_), .A3(new_n1747_), .ZN(new_n1748_));
  NOR4_X1    g1363(.A1(new_n1603_), .A2(new_n1621_), .A3(new_n1622_), .A4(new_n1624_), .ZN(new_n1749_));
  NAND4_X1   g1364(.A1(new_n1739_), .A2(new_n1749_), .A3(new_n1744_), .A4(new_n1748_), .ZN(new_n1750_));
  AOI21_X1   g1365(.A1(new_n1750_), .A2(new_n1732_), .B(new_n793_), .ZN(\grant[18] ));
  NOR4_X1    g1366(.A1(new_n1628_), .A2(new_n1629_), .A3(new_n1631_), .A4(new_n1639_), .ZN(new_n1752_));
  NOR2_X1    g1367(.A1(new_n1021_), .A2(new_n1022_), .ZN(new_n1753_));
  NOR2_X1    g1368(.A1(new_n1563_), .A2(new_n1753_), .ZN(new_n1754_));
  OAI22_X1   g1369(.A1(new_n797_), .A2(new_n804_), .B1(new_n1634_), .B2(new_n1633_), .ZN(new_n1755_));
  OAI22_X1   g1370(.A1(new_n1567_), .A2(new_n1569_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n1756_));
  NOR4_X1    g1371(.A1(new_n1640_), .A2(new_n1755_), .A3(new_n1756_), .A4(new_n1754_), .ZN(new_n1757_));
  INV_X1     g1372(.I(\req[20] ), .ZN(new_n1758_));
  AOI21_X1   g1373(.A1(new_n1758_), .A2(\priority[20] ), .B(\priority[21] ), .ZN(new_n1759_));
  OAI21_X1   g1374(.A1(new_n848_), .A2(new_n843_), .B(new_n1759_), .ZN(new_n1760_));
  NOR3_X1    g1375(.A1(new_n1646_), .A2(new_n1650_), .A3(new_n1760_), .ZN(new_n1761_));
  NOR4_X1    g1376(.A1(new_n1630_), .A2(new_n1648_), .A3(new_n1649_), .A4(new_n1651_), .ZN(new_n1762_));
  NAND4_X1   g1377(.A1(new_n1752_), .A2(new_n1762_), .A3(new_n1757_), .A4(new_n1761_), .ZN(new_n1763_));
  AOI21_X1   g1378(.A1(new_n1763_), .A2(new_n1745_), .B(new_n1039_), .ZN(\grant[19] ));
  NOR2_X1    g1379(.A1(new_n1050_), .A2(new_n1043_), .ZN(new_n1765_));
  OAI22_X1   g1380(.A1(new_n522_), .A2(new_n1656_), .B1(new_n955_), .B2(new_n950_), .ZN(new_n1766_));
  NOR4_X1    g1381(.A1(new_n973_), .A2(new_n1007_), .A3(new_n1766_), .A4(new_n1765_), .ZN(new_n1767_));
  INV_X1     g1382(.I(\req[21] ), .ZN(new_n1768_));
  AOI21_X1   g1383(.A1(new_n1768_), .A2(\priority[21] ), .B(\priority[22] ), .ZN(new_n1769_));
  OAI21_X1   g1384(.A1(new_n533_), .A2(new_n528_), .B(new_n1769_), .ZN(new_n1770_));
  OAI22_X1   g1385(.A1(new_n536_), .A2(new_n541_), .B1(new_n550_), .B2(new_n545_), .ZN(new_n1771_));
  NOR3_X1    g1386(.A1(new_n1103_), .A2(new_n1771_), .A3(new_n1770_), .ZN(new_n1772_));
  NAND4_X1   g1387(.A1(new_n1655_), .A2(new_n1664_), .A3(new_n1767_), .A4(new_n1772_), .ZN(new_n1773_));
  AOI21_X1   g1388(.A1(new_n1773_), .A2(new_n1758_), .B(new_n552_), .ZN(\grant[20] ));
  NOR2_X1    g1389(.A1(new_n1180_), .A2(new_n556_), .ZN(new_n1775_));
  OAI22_X1   g1390(.A1(new_n1146_), .A2(new_n1150_), .B1(new_n768_), .B2(new_n1668_), .ZN(new_n1776_));
  NOR4_X1    g1391(.A1(new_n1156_), .A2(new_n1166_), .A3(new_n1776_), .A4(new_n1775_), .ZN(new_n1777_));
  INV_X1     g1392(.I(\req[22] ), .ZN(new_n1778_));
  AOI21_X1   g1393(.A1(new_n1778_), .A2(\priority[22] ), .B(\priority[23] ), .ZN(new_n1779_));
  OAI21_X1   g1394(.A1(new_n779_), .A2(new_n774_), .B(new_n1779_), .ZN(new_n1780_));
  OAI22_X1   g1395(.A1(new_n782_), .A2(new_n787_), .B1(new_n796_), .B2(new_n791_), .ZN(new_n1781_));
  NOR3_X1    g1396(.A1(new_n1197_), .A2(new_n1781_), .A3(new_n1780_), .ZN(new_n1782_));
  NAND4_X1   g1397(.A1(new_n1667_), .A2(new_n1676_), .A3(new_n1777_), .A4(new_n1782_), .ZN(new_n1783_));
  AOI21_X1   g1398(.A1(new_n1783_), .A2(new_n1768_), .B(new_n798_), .ZN(\grant[21] ));
  NOR2_X1    g1399(.A1(new_n1262_), .A2(new_n802_), .ZN(new_n1785_));
  OAI22_X1   g1400(.A1(new_n1228_), .A2(new_n1232_), .B1(new_n1014_), .B2(new_n1680_), .ZN(new_n1786_));
  NOR4_X1    g1401(.A1(new_n1238_), .A2(new_n1248_), .A3(new_n1786_), .A4(new_n1785_), .ZN(new_n1787_));
  INV_X1     g1402(.I(\req[23] ), .ZN(new_n1788_));
  AOI21_X1   g1403(.A1(new_n1788_), .A2(\priority[23] ), .B(\priority[24] ), .ZN(new_n1789_));
  OAI21_X1   g1404(.A1(new_n1025_), .A2(new_n1020_), .B(new_n1789_), .ZN(new_n1790_));
  OAI22_X1   g1405(.A1(new_n1028_), .A2(new_n1033_), .B1(new_n1042_), .B2(new_n1037_), .ZN(new_n1791_));
  NOR3_X1    g1406(.A1(new_n1279_), .A2(new_n1791_), .A3(new_n1790_), .ZN(new_n1792_));
  NAND4_X1   g1407(.A1(new_n1679_), .A2(new_n1688_), .A3(new_n1787_), .A4(new_n1792_), .ZN(new_n1793_));
  AOI21_X1   g1408(.A1(new_n1793_), .A2(new_n1778_), .B(new_n1044_), .ZN(\grant[22] ));
  NOR2_X1    g1409(.A1(new_n1341_), .A2(new_n1048_), .ZN(new_n1795_));
  OAI22_X1   g1410(.A1(new_n1692_), .A2(new_n1168_), .B1(new_n1311_), .B2(new_n1310_), .ZN(new_n1796_));
  NOR4_X1    g1411(.A1(new_n1317_), .A2(new_n1327_), .A3(new_n1796_), .A4(new_n1795_), .ZN(new_n1797_));
  INV_X1     g1412(.I(\req[24] ), .ZN(new_n1798_));
  AOI21_X1   g1413(.A1(new_n1798_), .A2(\priority[24] ), .B(\priority[25] ), .ZN(new_n1799_));
  OAI21_X1   g1414(.A1(new_n1174_), .A2(new_n1172_), .B(new_n1799_), .ZN(new_n1800_));
  OAI22_X1   g1415(.A1(new_n1173_), .A2(new_n1175_), .B1(new_n1179_), .B2(new_n1177_), .ZN(new_n1801_));
  NOR3_X1    g1416(.A1(new_n1358_), .A2(new_n1801_), .A3(new_n1800_), .ZN(new_n1802_));
  NAND4_X1   g1417(.A1(new_n1691_), .A2(new_n1700_), .A3(new_n1797_), .A4(new_n1802_), .ZN(new_n1803_));
  AOI21_X1   g1418(.A1(new_n1803_), .A2(new_n1788_), .B(new_n557_), .ZN(\grant[23] ));
  NOR2_X1    g1419(.A1(new_n1419_), .A2(new_n598_), .ZN(new_n1805_));
  OAI22_X1   g1420(.A1(new_n1704_), .A2(new_n1250_), .B1(new_n1389_), .B2(new_n1388_), .ZN(new_n1806_));
  NOR4_X1    g1421(.A1(new_n1395_), .A2(new_n1405_), .A3(new_n1806_), .A4(new_n1805_), .ZN(new_n1807_));
  INV_X1     g1422(.I(\req[25] ), .ZN(new_n1808_));
  AOI21_X1   g1423(.A1(new_n1808_), .A2(\priority[25] ), .B(\priority[26] ), .ZN(new_n1809_));
  OAI21_X1   g1424(.A1(new_n1256_), .A2(new_n1254_), .B(new_n1809_), .ZN(new_n1810_));
  OAI22_X1   g1425(.A1(new_n1255_), .A2(new_n1257_), .B1(new_n1261_), .B2(new_n1259_), .ZN(new_n1811_));
  NOR3_X1    g1426(.A1(new_n1436_), .A2(new_n1811_), .A3(new_n1810_), .ZN(new_n1812_));
  NAND4_X1   g1427(.A1(new_n1703_), .A2(new_n1712_), .A3(new_n1807_), .A4(new_n1812_), .ZN(new_n1813_));
  AOI21_X1   g1428(.A1(new_n1813_), .A2(new_n1798_), .B(new_n803_), .ZN(\grant[24] ));
  NOR2_X1    g1429(.A1(new_n1497_), .A2(new_n844_), .ZN(new_n1815_));
  OAI22_X1   g1430(.A1(new_n1716_), .A2(new_n1329_), .B1(new_n1467_), .B2(new_n1466_), .ZN(new_n1816_));
  NOR4_X1    g1431(.A1(new_n1473_), .A2(new_n1483_), .A3(new_n1816_), .A4(new_n1815_), .ZN(new_n1817_));
  INV_X1     g1432(.I(\req[26] ), .ZN(new_n1818_));
  AOI21_X1   g1433(.A1(new_n1818_), .A2(\priority[26] ), .B(\priority[27] ), .ZN(new_n1819_));
  OAI21_X1   g1434(.A1(new_n1335_), .A2(new_n1333_), .B(new_n1819_), .ZN(new_n1820_));
  OAI22_X1   g1435(.A1(new_n1334_), .A2(new_n1336_), .B1(new_n1340_), .B2(new_n1338_), .ZN(new_n1821_));
  NOR3_X1    g1436(.A1(new_n1514_), .A2(new_n1821_), .A3(new_n1820_), .ZN(new_n1822_));
  NAND4_X1   g1437(.A1(new_n1715_), .A2(new_n1724_), .A3(new_n1817_), .A4(new_n1822_), .ZN(new_n1823_));
  AOI21_X1   g1438(.A1(new_n1823_), .A2(new_n1808_), .B(new_n1049_), .ZN(\grant[25] ));
  NOR2_X1    g1439(.A1(new_n1575_), .A2(new_n1090_), .ZN(new_n1825_));
  OAI22_X1   g1440(.A1(new_n1544_), .A2(new_n1545_), .B1(new_n1407_), .B2(new_n1728_), .ZN(new_n1826_));
  NOR4_X1    g1441(.A1(new_n1551_), .A2(new_n1561_), .A3(new_n1826_), .A4(new_n1825_), .ZN(new_n1827_));
  INV_X1     g1442(.I(\req[27] ), .ZN(new_n1828_));
  AOI21_X1   g1443(.A1(new_n1828_), .A2(\priority[27] ), .B(\priority[28] ), .ZN(new_n1829_));
  OAI21_X1   g1444(.A1(new_n1413_), .A2(new_n1411_), .B(new_n1829_), .ZN(new_n1830_));
  OAI22_X1   g1445(.A1(new_n1412_), .A2(new_n1414_), .B1(new_n1418_), .B2(new_n1416_), .ZN(new_n1831_));
  NOR3_X1    g1446(.A1(new_n1592_), .A2(new_n1831_), .A3(new_n1830_), .ZN(new_n1832_));
  NAND4_X1   g1447(.A1(new_n1727_), .A2(new_n1736_), .A3(new_n1827_), .A4(new_n1832_), .ZN(new_n1833_));
  AOI21_X1   g1448(.A1(new_n1833_), .A2(new_n1818_), .B(new_n599_), .ZN(\grant[26] ));
  NOR4_X1    g1449(.A1(new_n1601_), .A2(new_n1602_), .A3(new_n1612_), .A4(new_n1613_), .ZN(new_n1835_));
  NOR2_X1    g1450(.A1(new_n610_), .A2(new_n603_), .ZN(new_n1836_));
  OAI22_X1   g1451(.A1(new_n1606_), .A2(new_n1607_), .B1(new_n1485_), .B2(new_n1740_), .ZN(new_n1837_));
  OAI22_X1   g1452(.A1(new_n1494_), .A2(new_n1496_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n1838_));
  NOR4_X1    g1453(.A1(new_n1493_), .A2(new_n1837_), .A3(new_n1838_), .A4(new_n1836_), .ZN(new_n1839_));
  INV_X1     g1454(.I(\req[28] ), .ZN(new_n1840_));
  AOI21_X1   g1455(.A1(new_n1840_), .A2(\priority[28] ), .B(\priority[29] ), .ZN(new_n1841_));
  OAI21_X1   g1456(.A1(new_n619_), .A2(new_n614_), .B(new_n1841_), .ZN(new_n1842_));
  NOR3_X1    g1457(.A1(new_n1623_), .A2(new_n1624_), .A3(new_n1842_), .ZN(new_n1843_));
  NOR4_X1    g1458(.A1(new_n1603_), .A2(new_n1604_), .A3(new_n1621_), .A4(new_n1622_), .ZN(new_n1844_));
  NAND4_X1   g1459(.A1(new_n1835_), .A2(new_n1844_), .A3(new_n1839_), .A4(new_n1843_), .ZN(new_n1845_));
  AOI21_X1   g1460(.A1(new_n1845_), .A2(new_n1828_), .B(new_n845_), .ZN(\grant[27] ));
  NOR4_X1    g1461(.A1(new_n1628_), .A2(new_n1629_), .A3(new_n1639_), .A4(new_n1640_), .ZN(new_n1847_));
  NOR2_X1    g1462(.A1(new_n856_), .A2(new_n849_), .ZN(new_n1848_));
  OAI22_X1   g1463(.A1(new_n1633_), .A2(new_n1634_), .B1(new_n1563_), .B2(new_n1753_), .ZN(new_n1849_));
  OAI22_X1   g1464(.A1(new_n1572_), .A2(new_n1574_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n1850_));
  NOR4_X1    g1465(.A1(new_n1571_), .A2(new_n1849_), .A3(new_n1850_), .A4(new_n1848_), .ZN(new_n1851_));
  INV_X1     g1466(.I(\req[29] ), .ZN(new_n1852_));
  AOI21_X1   g1467(.A1(new_n1852_), .A2(\priority[29] ), .B(\priority[30] ), .ZN(new_n1853_));
  OAI21_X1   g1468(.A1(new_n865_), .A2(new_n860_), .B(new_n1853_), .ZN(new_n1854_));
  NOR3_X1    g1469(.A1(new_n1650_), .A2(new_n1651_), .A3(new_n1854_), .ZN(new_n1855_));
  NOR4_X1    g1470(.A1(new_n1630_), .A2(new_n1631_), .A3(new_n1648_), .A4(new_n1649_), .ZN(new_n1856_));
  NAND4_X1   g1471(.A1(new_n1847_), .A2(new_n1856_), .A3(new_n1851_), .A4(new_n1855_), .ZN(new_n1857_));
  AOI21_X1   g1472(.A1(new_n1857_), .A2(new_n1840_), .B(new_n1091_), .ZN(\grant[28] ));
  NOR2_X1    g1473(.A1(new_n1102_), .A2(new_n1095_), .ZN(new_n1859_));
  NOR4_X1    g1474(.A1(new_n973_), .A2(new_n1007_), .A3(new_n1766_), .A4(new_n1859_), .ZN(new_n1860_));
  INV_X1     g1475(.I(\req[30] ), .ZN(new_n1861_));
  AOI21_X1   g1476(.A1(new_n1861_), .A2(\priority[30] ), .B(\priority[31] ), .ZN(new_n1862_));
  OAI21_X1   g1477(.A1(new_n533_), .A2(new_n528_), .B(new_n1862_), .ZN(new_n1863_));
  NOR3_X1    g1478(.A1(new_n1618_), .A2(new_n1771_), .A3(new_n1863_), .ZN(new_n1864_));
  NAND4_X1   g1479(.A1(new_n1655_), .A2(new_n1664_), .A3(new_n1860_), .A4(new_n1864_), .ZN(new_n1865_));
  AOI21_X1   g1480(.A1(new_n1865_), .A2(new_n1852_), .B(new_n604_), .ZN(\grant[29] ));
  NOR2_X1    g1481(.A1(new_n1196_), .A2(new_n608_), .ZN(new_n1867_));
  NOR4_X1    g1482(.A1(new_n1156_), .A2(new_n1166_), .A3(new_n1776_), .A4(new_n1867_), .ZN(new_n1868_));
  INV_X1     g1483(.I(\req[31] ), .ZN(new_n1869_));
  AOI21_X1   g1484(.A1(new_n1869_), .A2(\priority[31] ), .B(\priority[32] ), .ZN(new_n1870_));
  OAI21_X1   g1485(.A1(new_n779_), .A2(new_n774_), .B(new_n1870_), .ZN(new_n1871_));
  NOR3_X1    g1486(.A1(new_n1645_), .A2(new_n1781_), .A3(new_n1871_), .ZN(new_n1872_));
  NAND4_X1   g1487(.A1(new_n1667_), .A2(new_n1676_), .A3(new_n1868_), .A4(new_n1872_), .ZN(new_n1873_));
  AOI21_X1   g1488(.A1(new_n1873_), .A2(new_n1861_), .B(new_n850_), .ZN(\grant[30] ));
  NOR2_X1    g1489(.A1(new_n1278_), .A2(new_n854_), .ZN(new_n1875_));
  NOR4_X1    g1490(.A1(new_n1238_), .A2(new_n1248_), .A3(new_n1786_), .A4(new_n1875_), .ZN(new_n1876_));
  INV_X1     g1491(.I(\req[32] ), .ZN(new_n1877_));
  AOI21_X1   g1492(.A1(new_n1877_), .A2(\priority[32] ), .B(\priority[33] ), .ZN(new_n1878_));
  OAI21_X1   g1493(.A1(new_n1025_), .A2(new_n1020_), .B(new_n1878_), .ZN(new_n1879_));
  OAI22_X1   g1494(.A1(new_n1045_), .A2(new_n1050_), .B1(new_n1094_), .B2(new_n1089_), .ZN(new_n1880_));
  NOR3_X1    g1495(.A1(new_n1791_), .A2(new_n1880_), .A3(new_n1879_), .ZN(new_n1881_));
  NAND4_X1   g1496(.A1(new_n1679_), .A2(new_n1688_), .A3(new_n1876_), .A4(new_n1881_), .ZN(new_n1882_));
  AOI21_X1   g1497(.A1(new_n1882_), .A2(new_n1869_), .B(new_n1096_), .ZN(\grant[31] ));
  NOR2_X1    g1498(.A1(new_n1357_), .A2(new_n1100_), .ZN(new_n1884_));
  NOR4_X1    g1499(.A1(new_n1317_), .A2(new_n1327_), .A3(new_n1796_), .A4(new_n1884_), .ZN(new_n1885_));
  INV_X1     g1500(.I(\req[33] ), .ZN(new_n1886_));
  AOI21_X1   g1501(.A1(new_n1886_), .A2(\priority[33] ), .B(\priority[34] ), .ZN(new_n1887_));
  OAI21_X1   g1502(.A1(new_n1174_), .A2(new_n1172_), .B(new_n1887_), .ZN(new_n1888_));
  OAI22_X1   g1503(.A1(new_n1178_), .A2(new_n1180_), .B1(new_n1195_), .B2(new_n1193_), .ZN(new_n1889_));
  NOR3_X1    g1504(.A1(new_n1801_), .A2(new_n1889_), .A3(new_n1888_), .ZN(new_n1890_));
  NAND4_X1   g1505(.A1(new_n1691_), .A2(new_n1700_), .A3(new_n1885_), .A4(new_n1890_), .ZN(new_n1891_));
  AOI21_X1   g1506(.A1(new_n1891_), .A2(new_n1877_), .B(new_n609_), .ZN(\grant[32] ));
  NOR2_X1    g1507(.A1(new_n1435_), .A2(new_n615_), .ZN(new_n1893_));
  NOR4_X1    g1508(.A1(new_n1395_), .A2(new_n1405_), .A3(new_n1806_), .A4(new_n1893_), .ZN(new_n1894_));
  INV_X1     g1509(.I(\req[34] ), .ZN(new_n1895_));
  AOI21_X1   g1510(.A1(new_n1895_), .A2(\priority[34] ), .B(\priority[35] ), .ZN(new_n1896_));
  OAI21_X1   g1511(.A1(new_n1256_), .A2(new_n1254_), .B(new_n1896_), .ZN(new_n1897_));
  OAI22_X1   g1512(.A1(new_n1260_), .A2(new_n1262_), .B1(new_n1277_), .B2(new_n1275_), .ZN(new_n1898_));
  NOR3_X1    g1513(.A1(new_n1811_), .A2(new_n1898_), .A3(new_n1897_), .ZN(new_n1899_));
  NAND4_X1   g1514(.A1(new_n1703_), .A2(new_n1712_), .A3(new_n1894_), .A4(new_n1899_), .ZN(new_n1900_));
  AOI21_X1   g1515(.A1(new_n1900_), .A2(new_n1886_), .B(new_n855_), .ZN(\grant[33] ));
  NOR2_X1    g1516(.A1(new_n1513_), .A2(new_n861_), .ZN(new_n1902_));
  NOR4_X1    g1517(.A1(new_n1473_), .A2(new_n1483_), .A3(new_n1816_), .A4(new_n1902_), .ZN(new_n1903_));
  INV_X1     g1518(.I(\req[35] ), .ZN(new_n1904_));
  AOI21_X1   g1519(.A1(new_n1904_), .A2(\priority[35] ), .B(\priority[36] ), .ZN(new_n1905_));
  OAI21_X1   g1520(.A1(new_n1335_), .A2(new_n1333_), .B(new_n1905_), .ZN(new_n1906_));
  OAI22_X1   g1521(.A1(new_n1339_), .A2(new_n1341_), .B1(new_n1356_), .B2(new_n1354_), .ZN(new_n1907_));
  NOR3_X1    g1522(.A1(new_n1821_), .A2(new_n1907_), .A3(new_n1906_), .ZN(new_n1908_));
  NAND4_X1   g1523(.A1(new_n1715_), .A2(new_n1724_), .A3(new_n1903_), .A4(new_n1908_), .ZN(new_n1909_));
  AOI21_X1   g1524(.A1(new_n1909_), .A2(new_n1895_), .B(new_n1101_), .ZN(\grant[34] ));
  NOR2_X1    g1525(.A1(new_n1591_), .A2(new_n1107_), .ZN(new_n1911_));
  NOR4_X1    g1526(.A1(new_n1551_), .A2(new_n1561_), .A3(new_n1826_), .A4(new_n1911_), .ZN(new_n1912_));
  INV_X1     g1527(.I(\req[36] ), .ZN(new_n1913_));
  AOI21_X1   g1528(.A1(new_n1913_), .A2(\priority[36] ), .B(\priority[37] ), .ZN(new_n1914_));
  OAI21_X1   g1529(.A1(new_n1413_), .A2(new_n1411_), .B(new_n1914_), .ZN(new_n1915_));
  OAI22_X1   g1530(.A1(new_n1417_), .A2(new_n1419_), .B1(new_n1434_), .B2(new_n1432_), .ZN(new_n1916_));
  NOR3_X1    g1531(.A1(new_n1831_), .A2(new_n1916_), .A3(new_n1915_), .ZN(new_n1917_));
  NAND4_X1   g1532(.A1(new_n1727_), .A2(new_n1736_), .A3(new_n1912_), .A4(new_n1917_), .ZN(new_n1918_));
  AOI21_X1   g1533(.A1(new_n1918_), .A2(new_n1904_), .B(new_n616_), .ZN(\grant[35] ));
  NOR4_X1    g1534(.A1(new_n1493_), .A2(new_n1602_), .A3(new_n1612_), .A4(new_n1613_), .ZN(new_n1920_));
  NOR2_X1    g1535(.A1(new_n627_), .A2(new_n620_), .ZN(new_n1921_));
  OAI22_X1   g1536(.A1(new_n1510_), .A2(new_n1512_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n1922_));
  NOR4_X1    g1537(.A1(new_n1498_), .A2(new_n1837_), .A3(new_n1922_), .A4(new_n1921_), .ZN(new_n1923_));
  INV_X1     g1538(.I(\req[37] ), .ZN(new_n1924_));
  AOI21_X1   g1539(.A1(new_n1924_), .A2(\priority[37] ), .B(\priority[38] ), .ZN(new_n1925_));
  OAI21_X1   g1540(.A1(new_n568_), .A2(new_n563_), .B(new_n1925_), .ZN(new_n1926_));
  NOR3_X1    g1541(.A1(new_n1621_), .A2(new_n1624_), .A3(new_n1926_), .ZN(new_n1927_));
  NOR4_X1    g1542(.A1(new_n1601_), .A2(new_n1603_), .A3(new_n1604_), .A4(new_n1622_), .ZN(new_n1928_));
  NAND4_X1   g1543(.A1(new_n1920_), .A2(new_n1928_), .A3(new_n1923_), .A4(new_n1927_), .ZN(new_n1929_));
  AOI21_X1   g1544(.A1(new_n1929_), .A2(new_n1913_), .B(new_n862_), .ZN(\grant[36] ));
  NOR4_X1    g1545(.A1(new_n1571_), .A2(new_n1629_), .A3(new_n1639_), .A4(new_n1640_), .ZN(new_n1931_));
  NOR2_X1    g1546(.A1(new_n873_), .A2(new_n866_), .ZN(new_n1932_));
  OAI22_X1   g1547(.A1(new_n1588_), .A2(new_n1590_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n1933_));
  NOR4_X1    g1548(.A1(new_n1576_), .A2(new_n1849_), .A3(new_n1933_), .A4(new_n1932_), .ZN(new_n1934_));
  INV_X1     g1549(.I(\req[38] ), .ZN(new_n1935_));
  AOI21_X1   g1550(.A1(new_n1935_), .A2(\priority[38] ), .B(\priority[39] ), .ZN(new_n1936_));
  OAI21_X1   g1551(.A1(new_n814_), .A2(new_n809_), .B(new_n1936_), .ZN(new_n1937_));
  NOR3_X1    g1552(.A1(new_n1648_), .A2(new_n1651_), .A3(new_n1937_), .ZN(new_n1938_));
  NOR4_X1    g1553(.A1(new_n1628_), .A2(new_n1630_), .A3(new_n1631_), .A4(new_n1649_), .ZN(new_n1939_));
  NAND4_X1   g1554(.A1(new_n1931_), .A2(new_n1939_), .A3(new_n1934_), .A4(new_n1938_), .ZN(new_n1940_));
  AOI21_X1   g1555(.A1(new_n1940_), .A2(new_n1924_), .B(new_n1108_), .ZN(\grant[37] ));
  NOR2_X1    g1556(.A1(new_n1119_), .A2(new_n1112_), .ZN(new_n1942_));
  NOR4_X1    g1557(.A1(new_n973_), .A2(new_n1007_), .A3(new_n1766_), .A4(new_n1942_), .ZN(new_n1943_));
  INV_X1     g1558(.I(\req[39] ), .ZN(new_n1944_));
  AOI21_X1   g1559(.A1(new_n1944_), .A2(\priority[39] ), .B(\priority[40] ), .ZN(new_n1945_));
  OAI21_X1   g1560(.A1(new_n533_), .A2(new_n528_), .B(new_n1945_), .ZN(new_n1946_));
  NOR3_X1    g1561(.A1(new_n1618_), .A2(new_n1771_), .A3(new_n1946_), .ZN(new_n1947_));
  NOR4_X1    g1562(.A1(new_n929_), .A2(new_n1069_), .A3(new_n1086_), .A4(new_n1619_), .ZN(new_n1948_));
  NAND4_X1   g1563(.A1(new_n1655_), .A2(new_n1948_), .A3(new_n1943_), .A4(new_n1947_), .ZN(new_n1949_));
  AOI21_X1   g1564(.A1(new_n1949_), .A2(new_n1935_), .B(new_n621_), .ZN(\grant[38] ));
  NOR2_X1    g1565(.A1(new_n1201_), .A2(new_n625_), .ZN(new_n1951_));
  NOR4_X1    g1566(.A1(new_n1156_), .A2(new_n1166_), .A3(new_n1776_), .A4(new_n1951_), .ZN(new_n1952_));
  INV_X1     g1567(.I(\req[40] ), .ZN(new_n1953_));
  AOI21_X1   g1568(.A1(new_n1953_), .A2(\priority[40] ), .B(\priority[41] ), .ZN(new_n1954_));
  OAI21_X1   g1569(.A1(new_n779_), .A2(new_n774_), .B(new_n1954_), .ZN(new_n1955_));
  NOR3_X1    g1570(.A1(new_n1645_), .A2(new_n1781_), .A3(new_n1955_), .ZN(new_n1956_));
  NOR4_X1    g1571(.A1(new_n1139_), .A2(new_n1187_), .A3(new_n1192_), .A4(new_n1646_), .ZN(new_n1957_));
  NAND4_X1   g1572(.A1(new_n1667_), .A2(new_n1957_), .A3(new_n1952_), .A4(new_n1956_), .ZN(new_n1958_));
  AOI21_X1   g1573(.A1(new_n1958_), .A2(new_n1944_), .B(new_n867_), .ZN(\grant[39] ));
  NOR2_X1    g1574(.A1(new_n1283_), .A2(new_n871_), .ZN(new_n1960_));
  NOR4_X1    g1575(.A1(new_n1238_), .A2(new_n1248_), .A3(new_n1786_), .A4(new_n1960_), .ZN(new_n1961_));
  INV_X1     g1576(.I(\req[41] ), .ZN(new_n1962_));
  AOI21_X1   g1577(.A1(new_n1962_), .A2(\priority[41] ), .B(\priority[42] ), .ZN(new_n1963_));
  OAI21_X1   g1578(.A1(new_n1025_), .A2(new_n1020_), .B(new_n1963_), .ZN(new_n1964_));
  NOR3_X1    g1579(.A1(new_n1791_), .A2(new_n1880_), .A3(new_n1964_), .ZN(new_n1965_));
  OAI22_X1   g1580(.A1(new_n1097_), .A2(new_n1102_), .B1(new_n1111_), .B2(new_n1106_), .ZN(new_n1966_));
  NOR4_X1    g1581(.A1(new_n1221_), .A2(new_n1269_), .A3(new_n1274_), .A4(new_n1966_), .ZN(new_n1967_));
  NAND4_X1   g1582(.A1(new_n1679_), .A2(new_n1967_), .A3(new_n1961_), .A4(new_n1965_), .ZN(new_n1968_));
  AOI21_X1   g1583(.A1(new_n1968_), .A2(new_n1953_), .B(new_n1113_), .ZN(\grant[40] ));
  NOR2_X1    g1584(.A1(new_n1362_), .A2(new_n1117_), .ZN(new_n1970_));
  NOR4_X1    g1585(.A1(new_n1317_), .A2(new_n1327_), .A3(new_n1796_), .A4(new_n1970_), .ZN(new_n1971_));
  INV_X1     g1586(.I(\req[42] ), .ZN(new_n1972_));
  AOI21_X1   g1587(.A1(new_n1972_), .A2(\priority[42] ), .B(\priority[43] ), .ZN(new_n1973_));
  OAI21_X1   g1588(.A1(new_n1174_), .A2(new_n1172_), .B(new_n1973_), .ZN(new_n1974_));
  NOR3_X1    g1589(.A1(new_n1801_), .A2(new_n1889_), .A3(new_n1974_), .ZN(new_n1975_));
  OAI22_X1   g1590(.A1(new_n1194_), .A2(new_n1196_), .B1(new_n1200_), .B2(new_n1198_), .ZN(new_n1976_));
  NOR4_X1    g1591(.A1(new_n1303_), .A2(new_n1348_), .A3(new_n1353_), .A4(new_n1976_), .ZN(new_n1977_));
  NAND4_X1   g1592(.A1(new_n1691_), .A2(new_n1977_), .A3(new_n1971_), .A4(new_n1975_), .ZN(new_n1978_));
  AOI21_X1   g1593(.A1(new_n1978_), .A2(new_n1962_), .B(new_n626_), .ZN(\grant[41] ));
  NOR2_X1    g1594(.A1(new_n1440_), .A2(new_n564_), .ZN(new_n1980_));
  NOR4_X1    g1595(.A1(new_n1395_), .A2(new_n1405_), .A3(new_n1806_), .A4(new_n1980_), .ZN(new_n1981_));
  INV_X1     g1596(.I(\req[43] ), .ZN(new_n1982_));
  AOI21_X1   g1597(.A1(new_n1982_), .A2(\priority[43] ), .B(\priority[44] ), .ZN(new_n1983_));
  OAI21_X1   g1598(.A1(new_n1256_), .A2(new_n1254_), .B(new_n1983_), .ZN(new_n1984_));
  NOR3_X1    g1599(.A1(new_n1811_), .A2(new_n1898_), .A3(new_n1984_), .ZN(new_n1985_));
  OAI22_X1   g1600(.A1(new_n1276_), .A2(new_n1278_), .B1(new_n1282_), .B2(new_n1280_), .ZN(new_n1986_));
  NOR4_X1    g1601(.A1(new_n1381_), .A2(new_n1426_), .A3(new_n1431_), .A4(new_n1986_), .ZN(new_n1987_));
  NAND4_X1   g1602(.A1(new_n1703_), .A2(new_n1987_), .A3(new_n1981_), .A4(new_n1985_), .ZN(new_n1988_));
  AOI21_X1   g1603(.A1(new_n1988_), .A2(new_n1972_), .B(new_n872_), .ZN(\grant[42] ));
  NOR2_X1    g1604(.A1(new_n1518_), .A2(new_n810_), .ZN(new_n1990_));
  NOR4_X1    g1605(.A1(new_n1473_), .A2(new_n1483_), .A3(new_n1816_), .A4(new_n1990_), .ZN(new_n1991_));
  INV_X1     g1606(.I(\req[44] ), .ZN(new_n1992_));
  AOI21_X1   g1607(.A1(new_n1992_), .A2(\priority[44] ), .B(\priority[45] ), .ZN(new_n1993_));
  OAI21_X1   g1608(.A1(new_n1335_), .A2(new_n1333_), .B(new_n1993_), .ZN(new_n1994_));
  NOR3_X1    g1609(.A1(new_n1821_), .A2(new_n1907_), .A3(new_n1994_), .ZN(new_n1995_));
  OAI22_X1   g1610(.A1(new_n1355_), .A2(new_n1357_), .B1(new_n1361_), .B2(new_n1359_), .ZN(new_n1996_));
  NOR4_X1    g1611(.A1(new_n1459_), .A2(new_n1504_), .A3(new_n1509_), .A4(new_n1996_), .ZN(new_n1997_));
  NAND4_X1   g1612(.A1(new_n1715_), .A2(new_n1997_), .A3(new_n1991_), .A4(new_n1995_), .ZN(new_n1998_));
  AOI21_X1   g1613(.A1(new_n1998_), .A2(new_n1982_), .B(new_n1118_), .ZN(\grant[43] ));
  NOR2_X1    g1614(.A1(new_n1596_), .A2(new_n1056_), .ZN(new_n2000_));
  NOR4_X1    g1615(.A1(new_n1551_), .A2(new_n1561_), .A3(new_n1826_), .A4(new_n2000_), .ZN(new_n2001_));
  INV_X1     g1616(.I(\req[45] ), .ZN(new_n2002_));
  AOI21_X1   g1617(.A1(new_n2002_), .A2(\priority[45] ), .B(\priority[46] ), .ZN(new_n2003_));
  OAI21_X1   g1618(.A1(new_n1413_), .A2(new_n1411_), .B(new_n2003_), .ZN(new_n2004_));
  NOR3_X1    g1619(.A1(new_n1831_), .A2(new_n1916_), .A3(new_n2004_), .ZN(new_n2005_));
  OAI22_X1   g1620(.A1(new_n1433_), .A2(new_n1435_), .B1(new_n1439_), .B2(new_n1438_), .ZN(new_n2006_));
  NOR4_X1    g1621(.A1(new_n1537_), .A2(new_n1582_), .A3(new_n1587_), .A4(new_n2006_), .ZN(new_n2007_));
  NAND4_X1   g1622(.A1(new_n1727_), .A2(new_n2007_), .A3(new_n2001_), .A4(new_n2005_), .ZN(new_n2008_));
  AOI21_X1   g1623(.A1(new_n2008_), .A2(new_n1992_), .B(new_n565_), .ZN(\grant[44] ));
  NOR4_X1    g1624(.A1(new_n1493_), .A2(new_n1498_), .A3(new_n1612_), .A4(new_n1613_), .ZN(new_n2010_));
  NOR2_X1    g1625(.A1(new_n576_), .A2(new_n569_), .ZN(new_n2011_));
  OAI22_X1   g1626(.A1(new_n1516_), .A2(new_n1517_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n2012_));
  NOR4_X1    g1627(.A1(new_n1514_), .A2(new_n1837_), .A3(new_n2012_), .A4(new_n2011_), .ZN(new_n2013_));
  INV_X1     g1628(.I(\req[46] ), .ZN(new_n2014_));
  AOI21_X1   g1629(.A1(new_n2014_), .A2(\priority[46] ), .B(\priority[47] ), .ZN(new_n2015_));
  OAI21_X1   g1630(.A1(new_n585_), .A2(new_n580_), .B(new_n2015_), .ZN(new_n2016_));
  NOR3_X1    g1631(.A1(new_n1621_), .A2(new_n1622_), .A3(new_n2016_), .ZN(new_n2017_));
  NAND4_X1   g1632(.A1(new_n1605_), .A2(new_n2010_), .A3(new_n2013_), .A4(new_n2017_), .ZN(new_n2018_));
  AOI21_X1   g1633(.A1(new_n2018_), .A2(new_n2002_), .B(new_n811_), .ZN(\grant[45] ));
  NOR4_X1    g1634(.A1(new_n1571_), .A2(new_n1576_), .A3(new_n1639_), .A4(new_n1640_), .ZN(new_n2020_));
  NOR2_X1    g1635(.A1(new_n822_), .A2(new_n815_), .ZN(new_n2021_));
  OAI22_X1   g1636(.A1(new_n1594_), .A2(new_n1595_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n2022_));
  NOR4_X1    g1637(.A1(new_n1592_), .A2(new_n1849_), .A3(new_n2022_), .A4(new_n2021_), .ZN(new_n2023_));
  INV_X1     g1638(.I(\req[47] ), .ZN(new_n2024_));
  AOI21_X1   g1639(.A1(new_n2024_), .A2(\priority[47] ), .B(\priority[48] ), .ZN(new_n2025_));
  OAI21_X1   g1640(.A1(new_n831_), .A2(new_n826_), .B(new_n2025_), .ZN(new_n2026_));
  NOR3_X1    g1641(.A1(new_n1648_), .A2(new_n1649_), .A3(new_n2026_), .ZN(new_n2027_));
  NAND4_X1   g1642(.A1(new_n1632_), .A2(new_n2020_), .A3(new_n2023_), .A4(new_n2027_), .ZN(new_n2028_));
  AOI21_X1   g1643(.A1(new_n2028_), .A2(new_n2014_), .B(new_n1057_), .ZN(\grant[46] ));
  NOR2_X1    g1644(.A1(new_n1068_), .A2(new_n1061_), .ZN(new_n2030_));
  NOR4_X1    g1645(.A1(new_n973_), .A2(new_n1007_), .A3(new_n1766_), .A4(new_n2030_), .ZN(new_n2031_));
  INV_X1     g1646(.I(\req[48] ), .ZN(new_n2032_));
  AOI21_X1   g1647(.A1(new_n2032_), .A2(\priority[48] ), .B(\priority[49] ), .ZN(new_n2033_));
  OAI21_X1   g1648(.A1(new_n533_), .A2(new_n528_), .B(new_n2033_), .ZN(new_n2034_));
  NOR3_X1    g1649(.A1(new_n1618_), .A2(new_n1771_), .A3(new_n2034_), .ZN(new_n2035_));
  NOR4_X1    g1650(.A1(new_n929_), .A2(new_n1086_), .A3(new_n1619_), .A4(new_n1623_), .ZN(new_n2036_));
  NAND4_X1   g1651(.A1(new_n1655_), .A2(new_n2036_), .A3(new_n2031_), .A4(new_n2035_), .ZN(new_n2037_));
  AOI21_X1   g1652(.A1(new_n2037_), .A2(new_n2024_), .B(new_n570_), .ZN(\grant[47] ));
  NOR2_X1    g1653(.A1(new_n1186_), .A2(new_n574_), .ZN(new_n2039_));
  NOR4_X1    g1654(.A1(new_n1156_), .A2(new_n1166_), .A3(new_n1776_), .A4(new_n2039_), .ZN(new_n2040_));
  INV_X1     g1655(.I(\req[49] ), .ZN(new_n2041_));
  AOI21_X1   g1656(.A1(new_n2041_), .A2(\priority[49] ), .B(\priority[50] ), .ZN(new_n2042_));
  OAI21_X1   g1657(.A1(new_n779_), .A2(new_n774_), .B(new_n2042_), .ZN(new_n2043_));
  NOR3_X1    g1658(.A1(new_n1645_), .A2(new_n1781_), .A3(new_n2043_), .ZN(new_n2044_));
  NOR4_X1    g1659(.A1(new_n1139_), .A2(new_n1192_), .A3(new_n1646_), .A4(new_n1650_), .ZN(new_n2045_));
  NAND4_X1   g1660(.A1(new_n1667_), .A2(new_n2045_), .A3(new_n2040_), .A4(new_n2044_), .ZN(new_n2046_));
  AOI21_X1   g1661(.A1(new_n2046_), .A2(new_n2032_), .B(new_n816_), .ZN(\grant[48] ));
  NOR2_X1    g1662(.A1(new_n1268_), .A2(new_n820_), .ZN(new_n2048_));
  NOR4_X1    g1663(.A1(new_n1238_), .A2(new_n1248_), .A3(new_n1786_), .A4(new_n2048_), .ZN(new_n2049_));
  INV_X1     g1664(.I(\req[50] ), .ZN(new_n2050_));
  AOI21_X1   g1665(.A1(new_n2050_), .A2(\priority[50] ), .B(\priority[51] ), .ZN(new_n2051_));
  OAI21_X1   g1666(.A1(new_n1025_), .A2(new_n1020_), .B(new_n2051_), .ZN(new_n2052_));
  NOR3_X1    g1667(.A1(new_n1791_), .A2(new_n1880_), .A3(new_n2052_), .ZN(new_n2053_));
  OAI22_X1   g1668(.A1(new_n1055_), .A2(new_n1060_), .B1(new_n1119_), .B2(new_n1114_), .ZN(new_n2054_));
  NOR4_X1    g1669(.A1(new_n1221_), .A2(new_n1274_), .A3(new_n1966_), .A4(new_n2054_), .ZN(new_n2055_));
  NAND4_X1   g1670(.A1(new_n1679_), .A2(new_n2055_), .A3(new_n2049_), .A4(new_n2053_), .ZN(new_n2056_));
  AOI21_X1   g1671(.A1(new_n2056_), .A2(new_n2041_), .B(new_n1062_), .ZN(\grant[49] ));
  NOR2_X1    g1672(.A1(new_n1347_), .A2(new_n1066_), .ZN(new_n2058_));
  NOR4_X1    g1673(.A1(new_n1317_), .A2(new_n1327_), .A3(new_n1796_), .A4(new_n2058_), .ZN(new_n2059_));
  INV_X1     g1674(.I(\req[51] ), .ZN(new_n2060_));
  AOI21_X1   g1675(.A1(new_n2060_), .A2(\priority[51] ), .B(\priority[52] ), .ZN(new_n2061_));
  OAI21_X1   g1676(.A1(new_n1174_), .A2(new_n1172_), .B(new_n2061_), .ZN(new_n2062_));
  NOR3_X1    g1677(.A1(new_n1801_), .A2(new_n1889_), .A3(new_n2062_), .ZN(new_n2063_));
  OAI22_X1   g1678(.A1(new_n1183_), .A2(new_n1185_), .B1(new_n1201_), .B2(new_n1199_), .ZN(new_n2064_));
  NOR4_X1    g1679(.A1(new_n1303_), .A2(new_n1353_), .A3(new_n1976_), .A4(new_n2064_), .ZN(new_n2065_));
  NAND4_X1   g1680(.A1(new_n1691_), .A2(new_n2065_), .A3(new_n2059_), .A4(new_n2063_), .ZN(new_n2066_));
  AOI21_X1   g1681(.A1(new_n2066_), .A2(new_n2050_), .B(new_n575_), .ZN(\grant[50] ));
  NOR2_X1    g1682(.A1(new_n1425_), .A2(new_n581_), .ZN(new_n2068_));
  NOR4_X1    g1683(.A1(new_n1395_), .A2(new_n1405_), .A3(new_n1806_), .A4(new_n2068_), .ZN(new_n2069_));
  INV_X1     g1684(.I(\req[52] ), .ZN(new_n2070_));
  AOI21_X1   g1685(.A1(new_n2070_), .A2(\priority[52] ), .B(\priority[53] ), .ZN(new_n2071_));
  OAI21_X1   g1686(.A1(new_n1256_), .A2(new_n1254_), .B(new_n2071_), .ZN(new_n2072_));
  NOR3_X1    g1687(.A1(new_n1811_), .A2(new_n1898_), .A3(new_n2072_), .ZN(new_n2073_));
  OAI22_X1   g1688(.A1(new_n1265_), .A2(new_n1267_), .B1(new_n1283_), .B2(new_n1281_), .ZN(new_n2074_));
  NOR4_X1    g1689(.A1(new_n1381_), .A2(new_n1431_), .A3(new_n1986_), .A4(new_n2074_), .ZN(new_n2075_));
  NAND4_X1   g1690(.A1(new_n1703_), .A2(new_n2075_), .A3(new_n2069_), .A4(new_n2073_), .ZN(new_n2076_));
  AOI21_X1   g1691(.A1(new_n2076_), .A2(new_n2060_), .B(new_n821_), .ZN(\grant[51] ));
  NOR2_X1    g1692(.A1(new_n1503_), .A2(new_n827_), .ZN(new_n2078_));
  NOR4_X1    g1693(.A1(new_n1473_), .A2(new_n1483_), .A3(new_n1816_), .A4(new_n2078_), .ZN(new_n2079_));
  INV_X1     g1694(.I(\req[53] ), .ZN(new_n2080_));
  AOI21_X1   g1695(.A1(new_n2080_), .A2(\priority[53] ), .B(\priority[54] ), .ZN(new_n2081_));
  OAI21_X1   g1696(.A1(new_n1335_), .A2(new_n1333_), .B(new_n2081_), .ZN(new_n2082_));
  NOR3_X1    g1697(.A1(new_n1821_), .A2(new_n1907_), .A3(new_n2082_), .ZN(new_n2083_));
  OAI22_X1   g1698(.A1(new_n1344_), .A2(new_n1346_), .B1(new_n1362_), .B2(new_n1360_), .ZN(new_n2084_));
  NOR4_X1    g1699(.A1(new_n1459_), .A2(new_n1509_), .A3(new_n1996_), .A4(new_n2084_), .ZN(new_n2085_));
  NAND4_X1   g1700(.A1(new_n1715_), .A2(new_n2085_), .A3(new_n2079_), .A4(new_n2083_), .ZN(new_n2086_));
  AOI21_X1   g1701(.A1(new_n2086_), .A2(new_n2070_), .B(new_n1067_), .ZN(\grant[52] ));
  NOR2_X1    g1702(.A1(new_n1581_), .A2(new_n1073_), .ZN(new_n2088_));
  NOR4_X1    g1703(.A1(new_n1551_), .A2(new_n1561_), .A3(new_n1826_), .A4(new_n2088_), .ZN(new_n2089_));
  INV_X1     g1704(.I(\req[54] ), .ZN(new_n2090_));
  AOI21_X1   g1705(.A1(new_n2090_), .A2(\priority[54] ), .B(\priority[55] ), .ZN(new_n2091_));
  OAI21_X1   g1706(.A1(new_n1413_), .A2(new_n1411_), .B(new_n2091_), .ZN(new_n2092_));
  NOR3_X1    g1707(.A1(new_n1831_), .A2(new_n1916_), .A3(new_n2092_), .ZN(new_n2093_));
  OAI22_X1   g1708(.A1(new_n1437_), .A2(new_n1440_), .B1(new_n1424_), .B2(new_n1422_), .ZN(new_n2094_));
  NOR4_X1    g1709(.A1(new_n1537_), .A2(new_n1587_), .A3(new_n2006_), .A4(new_n2094_), .ZN(new_n2095_));
  NAND4_X1   g1710(.A1(new_n1727_), .A2(new_n2095_), .A3(new_n2089_), .A4(new_n2093_), .ZN(new_n2096_));
  AOI21_X1   g1711(.A1(new_n2096_), .A2(new_n2080_), .B(new_n582_), .ZN(\grant[53] ));
  NOR4_X1    g1712(.A1(new_n1493_), .A2(new_n1498_), .A3(new_n1514_), .A4(new_n1613_), .ZN(new_n2098_));
  NOR2_X1    g1713(.A1(new_n593_), .A2(new_n586_), .ZN(new_n2099_));
  OAI22_X1   g1714(.A1(new_n1500_), .A2(new_n1502_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n2100_));
  NOR4_X1    g1715(.A1(new_n1519_), .A2(new_n1837_), .A3(new_n2100_), .A4(new_n2099_), .ZN(new_n2101_));
  INV_X1     g1716(.I(\req[55] ), .ZN(new_n2102_));
  AOI21_X1   g1717(.A1(new_n2102_), .A2(\priority[55] ), .B(\priority[56] ), .ZN(new_n2103_));
  OAI21_X1   g1718(.A1(new_n428_), .A2(new_n423_), .B(new_n2103_), .ZN(new_n2104_));
  NOR3_X1    g1719(.A1(new_n1603_), .A2(new_n1622_), .A3(new_n2104_), .ZN(new_n2105_));
  NAND4_X1   g1720(.A1(new_n1739_), .A2(new_n2098_), .A3(new_n2101_), .A4(new_n2105_), .ZN(new_n2106_));
  AOI21_X1   g1721(.A1(new_n2106_), .A2(new_n2090_), .B(new_n828_), .ZN(\grant[54] ));
  NOR4_X1    g1722(.A1(new_n1571_), .A2(new_n1576_), .A3(new_n1592_), .A4(new_n1640_), .ZN(new_n2108_));
  NOR2_X1    g1723(.A1(new_n839_), .A2(new_n832_), .ZN(new_n2109_));
  OAI22_X1   g1724(.A1(new_n1578_), .A2(new_n1580_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n2110_));
  NOR4_X1    g1725(.A1(new_n1597_), .A2(new_n1849_), .A3(new_n2110_), .A4(new_n2109_), .ZN(new_n2111_));
  INV_X1     g1726(.I(\req[56] ), .ZN(new_n2112_));
  AOI21_X1   g1727(.A1(new_n2112_), .A2(\priority[56] ), .B(\priority[57] ), .ZN(new_n2113_));
  OAI21_X1   g1728(.A1(new_n674_), .A2(new_n669_), .B(new_n2113_), .ZN(new_n2114_));
  NOR3_X1    g1729(.A1(new_n1630_), .A2(new_n1649_), .A3(new_n2114_), .ZN(new_n2115_));
  NAND4_X1   g1730(.A1(new_n1752_), .A2(new_n2108_), .A3(new_n2111_), .A4(new_n2115_), .ZN(new_n2116_));
  AOI21_X1   g1731(.A1(new_n2116_), .A2(new_n2102_), .B(new_n1074_), .ZN(\grant[55] ));
  NOR2_X1    g1732(.A1(new_n1085_), .A2(new_n1078_), .ZN(new_n2118_));
  NOR4_X1    g1733(.A1(new_n973_), .A2(new_n1007_), .A3(new_n1766_), .A4(new_n2118_), .ZN(new_n2119_));
  INV_X1     g1734(.I(\req[57] ), .ZN(new_n2120_));
  AOI21_X1   g1735(.A1(new_n2120_), .A2(\priority[57] ), .B(\priority[58] ), .ZN(new_n2121_));
  OAI21_X1   g1736(.A1(new_n533_), .A2(new_n528_), .B(new_n2121_), .ZN(new_n2122_));
  NOR3_X1    g1737(.A1(new_n1618_), .A2(new_n1771_), .A3(new_n2122_), .ZN(new_n2123_));
  NOR4_X1    g1738(.A1(new_n929_), .A2(new_n1619_), .A3(new_n1623_), .A4(new_n1624_), .ZN(new_n2124_));
  NAND4_X1   g1739(.A1(new_n1655_), .A2(new_n2124_), .A3(new_n2119_), .A4(new_n2123_), .ZN(new_n2125_));
  AOI21_X1   g1740(.A1(new_n2125_), .A2(new_n2112_), .B(new_n587_), .ZN(\grant[56] ));
  NOR2_X1    g1741(.A1(new_n1191_), .A2(new_n591_), .ZN(new_n2127_));
  NOR4_X1    g1742(.A1(new_n1156_), .A2(new_n1166_), .A3(new_n1776_), .A4(new_n2127_), .ZN(new_n2128_));
  INV_X1     g1743(.I(\req[58] ), .ZN(new_n2129_));
  AOI21_X1   g1744(.A1(new_n2129_), .A2(\priority[58] ), .B(\priority[59] ), .ZN(new_n2130_));
  OAI21_X1   g1745(.A1(new_n779_), .A2(new_n774_), .B(new_n2130_), .ZN(new_n2131_));
  NOR3_X1    g1746(.A1(new_n1645_), .A2(new_n1781_), .A3(new_n2131_), .ZN(new_n2132_));
  NOR4_X1    g1747(.A1(new_n1139_), .A2(new_n1646_), .A3(new_n1650_), .A4(new_n1651_), .ZN(new_n2133_));
  NAND4_X1   g1748(.A1(new_n1667_), .A2(new_n2133_), .A3(new_n2128_), .A4(new_n2132_), .ZN(new_n2134_));
  AOI21_X1   g1749(.A1(new_n2134_), .A2(new_n2120_), .B(new_n833_), .ZN(\grant[57] ));
  NOR2_X1    g1750(.A1(new_n1273_), .A2(new_n837_), .ZN(new_n2136_));
  NOR4_X1    g1751(.A1(new_n1238_), .A2(new_n1248_), .A3(new_n1786_), .A4(new_n2136_), .ZN(new_n2137_));
  INV_X1     g1752(.I(\req[59] ), .ZN(new_n2138_));
  AOI21_X1   g1753(.A1(new_n2138_), .A2(\priority[59] ), .B(\priority[60] ), .ZN(new_n2139_));
  OAI21_X1   g1754(.A1(new_n1025_), .A2(new_n1020_), .B(new_n2139_), .ZN(new_n2140_));
  NOR3_X1    g1755(.A1(new_n1791_), .A2(new_n1880_), .A3(new_n2140_), .ZN(new_n2141_));
  OAI22_X1   g1756(.A1(new_n1063_), .A2(new_n1068_), .B1(new_n1077_), .B2(new_n1072_), .ZN(new_n2142_));
  NOR4_X1    g1757(.A1(new_n1221_), .A2(new_n1966_), .A3(new_n2054_), .A4(new_n2142_), .ZN(new_n2143_));
  NAND4_X1   g1758(.A1(new_n1679_), .A2(new_n2143_), .A3(new_n2137_), .A4(new_n2141_), .ZN(new_n2144_));
  AOI21_X1   g1759(.A1(new_n2144_), .A2(new_n2129_), .B(new_n1079_), .ZN(\grant[58] ));
  NOR2_X1    g1760(.A1(new_n1352_), .A2(new_n1083_), .ZN(new_n2146_));
  NOR4_X1    g1761(.A1(new_n1317_), .A2(new_n1327_), .A3(new_n1796_), .A4(new_n2146_), .ZN(new_n2147_));
  INV_X1     g1762(.I(\req[60] ), .ZN(new_n2148_));
  AOI21_X1   g1763(.A1(new_n2148_), .A2(\priority[60] ), .B(\priority[61] ), .ZN(new_n2149_));
  OAI21_X1   g1764(.A1(new_n1174_), .A2(new_n1172_), .B(new_n2149_), .ZN(new_n2150_));
  NOR3_X1    g1765(.A1(new_n1801_), .A2(new_n1889_), .A3(new_n2150_), .ZN(new_n2151_));
  OAI22_X1   g1766(.A1(new_n1184_), .A2(new_n1186_), .B1(new_n1190_), .B2(new_n1188_), .ZN(new_n2152_));
  NOR4_X1    g1767(.A1(new_n1303_), .A2(new_n1976_), .A3(new_n2064_), .A4(new_n2152_), .ZN(new_n2153_));
  NAND4_X1   g1768(.A1(new_n1691_), .A2(new_n2153_), .A3(new_n2147_), .A4(new_n2151_), .ZN(new_n2154_));
  AOI21_X1   g1769(.A1(new_n2154_), .A2(new_n2138_), .B(new_n592_), .ZN(\grant[59] ));
  NOR2_X1    g1770(.A1(new_n1430_), .A2(new_n424_), .ZN(new_n2156_));
  NOR4_X1    g1771(.A1(new_n1395_), .A2(new_n1405_), .A3(new_n1806_), .A4(new_n2156_), .ZN(new_n2157_));
  INV_X1     g1772(.I(\req[61] ), .ZN(new_n2158_));
  AOI21_X1   g1773(.A1(new_n2158_), .A2(\priority[61] ), .B(\priority[62] ), .ZN(new_n2159_));
  OAI21_X1   g1774(.A1(new_n1256_), .A2(new_n1254_), .B(new_n2159_), .ZN(new_n2160_));
  NOR3_X1    g1775(.A1(new_n1811_), .A2(new_n1898_), .A3(new_n2160_), .ZN(new_n2161_));
  OAI22_X1   g1776(.A1(new_n1266_), .A2(new_n1268_), .B1(new_n1272_), .B2(new_n1270_), .ZN(new_n2162_));
  NOR4_X1    g1777(.A1(new_n1381_), .A2(new_n1986_), .A3(new_n2074_), .A4(new_n2162_), .ZN(new_n2163_));
  NAND4_X1   g1778(.A1(new_n1703_), .A2(new_n2163_), .A3(new_n2157_), .A4(new_n2161_), .ZN(new_n2164_));
  AOI21_X1   g1779(.A1(new_n2164_), .A2(new_n2148_), .B(new_n838_), .ZN(\grant[60] ));
  NOR2_X1    g1780(.A1(new_n1508_), .A2(new_n670_), .ZN(new_n2166_));
  NOR4_X1    g1781(.A1(new_n1473_), .A2(new_n1483_), .A3(new_n1816_), .A4(new_n2166_), .ZN(new_n2167_));
  INV_X1     g1782(.I(\req[62] ), .ZN(new_n2168_));
  AOI21_X1   g1783(.A1(new_n2168_), .A2(\priority[62] ), .B(\priority[63] ), .ZN(new_n2169_));
  OAI21_X1   g1784(.A1(new_n1335_), .A2(new_n1333_), .B(new_n2169_), .ZN(new_n2170_));
  NOR3_X1    g1785(.A1(new_n1821_), .A2(new_n1907_), .A3(new_n2170_), .ZN(new_n2171_));
  OAI22_X1   g1786(.A1(new_n1345_), .A2(new_n1347_), .B1(new_n1351_), .B2(new_n1349_), .ZN(new_n2172_));
  NOR4_X1    g1787(.A1(new_n1459_), .A2(new_n1996_), .A3(new_n2084_), .A4(new_n2172_), .ZN(new_n2173_));
  NAND4_X1   g1788(.A1(new_n1715_), .A2(new_n2173_), .A3(new_n2167_), .A4(new_n2171_), .ZN(new_n2174_));
  AOI21_X1   g1789(.A1(new_n2174_), .A2(new_n2158_), .B(new_n1084_), .ZN(\grant[61] ));
  NOR2_X1    g1790(.A1(new_n1586_), .A2(new_n916_), .ZN(new_n2176_));
  NOR4_X1    g1791(.A1(new_n1551_), .A2(new_n1561_), .A3(new_n1826_), .A4(new_n2176_), .ZN(new_n2177_));
  INV_X1     g1792(.I(\req[63] ), .ZN(new_n2178_));
  AOI21_X1   g1793(.A1(new_n2178_), .A2(\priority[63] ), .B(\priority[64] ), .ZN(new_n2179_));
  OAI21_X1   g1794(.A1(new_n1413_), .A2(new_n1411_), .B(new_n2179_), .ZN(new_n2180_));
  NOR3_X1    g1795(.A1(new_n1831_), .A2(new_n1916_), .A3(new_n2180_), .ZN(new_n2181_));
  OAI22_X1   g1796(.A1(new_n1423_), .A2(new_n1425_), .B1(new_n1429_), .B2(new_n1428_), .ZN(new_n2182_));
  NOR4_X1    g1797(.A1(new_n1537_), .A2(new_n2006_), .A3(new_n2094_), .A4(new_n2182_), .ZN(new_n2183_));
  NAND4_X1   g1798(.A1(new_n1727_), .A2(new_n2183_), .A3(new_n2177_), .A4(new_n2181_), .ZN(new_n2184_));
  AOI21_X1   g1799(.A1(new_n2184_), .A2(new_n2168_), .B(new_n425_), .ZN(\grant[62] ));
  NOR4_X1    g1800(.A1(new_n1493_), .A2(new_n1498_), .A3(new_n1514_), .A4(new_n1519_), .ZN(new_n2186_));
  NOR2_X1    g1801(.A1(new_n436_), .A2(new_n429_), .ZN(new_n2187_));
  OAI22_X1   g1802(.A1(new_n1506_), .A2(new_n1507_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n2188_));
  NOR4_X1    g1803(.A1(new_n1504_), .A2(new_n1837_), .A3(new_n2188_), .A4(new_n2187_), .ZN(new_n2189_));
  INV_X1     g1804(.I(\req[64] ), .ZN(new_n2190_));
  AOI21_X1   g1805(.A1(new_n2190_), .A2(\priority[64] ), .B(\priority[65] ), .ZN(new_n2191_));
  OAI21_X1   g1806(.A1(new_n445_), .A2(new_n440_), .B(new_n2191_), .ZN(new_n2192_));
  NOR3_X1    g1807(.A1(new_n1603_), .A2(new_n1604_), .A3(new_n2192_), .ZN(new_n2193_));
  NAND4_X1   g1808(.A1(new_n1835_), .A2(new_n2186_), .A3(new_n2189_), .A4(new_n2193_), .ZN(new_n2194_));
  AOI21_X1   g1809(.A1(new_n2194_), .A2(new_n2178_), .B(new_n671_), .ZN(\grant[63] ));
  NOR4_X1    g1810(.A1(new_n1571_), .A2(new_n1576_), .A3(new_n1592_), .A4(new_n1597_), .ZN(new_n2196_));
  NOR2_X1    g1811(.A1(new_n682_), .A2(new_n675_), .ZN(new_n2197_));
  OAI22_X1   g1812(.A1(new_n1584_), .A2(new_n1585_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n2198_));
  NOR4_X1    g1813(.A1(new_n1582_), .A2(new_n1849_), .A3(new_n2198_), .A4(new_n2197_), .ZN(new_n2199_));
  INV_X1     g1814(.I(\req[65] ), .ZN(new_n2200_));
  AOI21_X1   g1815(.A1(new_n2200_), .A2(\priority[65] ), .B(\priority[66] ), .ZN(new_n2201_));
  OAI21_X1   g1816(.A1(new_n691_), .A2(new_n686_), .B(new_n2201_), .ZN(new_n2202_));
  NOR3_X1    g1817(.A1(new_n1630_), .A2(new_n1631_), .A3(new_n2202_), .ZN(new_n2203_));
  NAND4_X1   g1818(.A1(new_n1847_), .A2(new_n2196_), .A3(new_n2199_), .A4(new_n2203_), .ZN(new_n2204_));
  AOI21_X1   g1819(.A1(new_n2204_), .A2(new_n2190_), .B(new_n917_), .ZN(\grant[64] ));
  NOR2_X1    g1820(.A1(new_n928_), .A2(new_n921_), .ZN(new_n2206_));
  NOR4_X1    g1821(.A1(new_n973_), .A2(new_n1007_), .A3(new_n1766_), .A4(new_n2206_), .ZN(new_n2207_));
  INV_X1     g1822(.I(\req[66] ), .ZN(new_n2208_));
  AOI21_X1   g1823(.A1(new_n2208_), .A2(\priority[66] ), .B(\priority[67] ), .ZN(new_n2209_));
  OAI21_X1   g1824(.A1(new_n533_), .A2(new_n528_), .B(new_n2209_), .ZN(new_n2210_));
  NOR3_X1    g1825(.A1(new_n1618_), .A2(new_n1771_), .A3(new_n2210_), .ZN(new_n2211_));
  NOR4_X1    g1826(.A1(new_n1619_), .A2(new_n1621_), .A3(new_n1623_), .A4(new_n1624_), .ZN(new_n2212_));
  NAND4_X1   g1827(.A1(new_n1655_), .A2(new_n2212_), .A3(new_n2207_), .A4(new_n2211_), .ZN(new_n2213_));
  AOI21_X1   g1828(.A1(new_n2213_), .A2(new_n2200_), .B(new_n430_), .ZN(\grant[65] ));
  NOR2_X1    g1829(.A1(new_n1138_), .A2(new_n434_), .ZN(new_n2215_));
  NOR4_X1    g1830(.A1(new_n1156_), .A2(new_n1166_), .A3(new_n1776_), .A4(new_n2215_), .ZN(new_n2216_));
  INV_X1     g1831(.I(\req[67] ), .ZN(new_n2217_));
  AOI21_X1   g1832(.A1(new_n2217_), .A2(\priority[67] ), .B(\priority[68] ), .ZN(new_n2218_));
  OAI21_X1   g1833(.A1(new_n779_), .A2(new_n774_), .B(new_n2218_), .ZN(new_n2219_));
  NOR3_X1    g1834(.A1(new_n1645_), .A2(new_n1781_), .A3(new_n2219_), .ZN(new_n2220_));
  NOR4_X1    g1835(.A1(new_n1646_), .A2(new_n1648_), .A3(new_n1650_), .A4(new_n1651_), .ZN(new_n2221_));
  NAND4_X1   g1836(.A1(new_n1667_), .A2(new_n2221_), .A3(new_n2216_), .A4(new_n2220_), .ZN(new_n2222_));
  AOI21_X1   g1837(.A1(new_n2222_), .A2(new_n2208_), .B(new_n676_), .ZN(\grant[66] ));
  NOR2_X1    g1838(.A1(new_n1220_), .A2(new_n680_), .ZN(new_n2224_));
  NOR4_X1    g1839(.A1(new_n1238_), .A2(new_n1248_), .A3(new_n1786_), .A4(new_n2224_), .ZN(new_n2225_));
  INV_X1     g1840(.I(\req[68] ), .ZN(new_n2226_));
  AOI21_X1   g1841(.A1(new_n2226_), .A2(\priority[68] ), .B(\priority[69] ), .ZN(new_n2227_));
  OAI21_X1   g1842(.A1(new_n1025_), .A2(new_n1020_), .B(new_n2227_), .ZN(new_n2228_));
  NOR3_X1    g1843(.A1(new_n1791_), .A2(new_n1880_), .A3(new_n2228_), .ZN(new_n2229_));
  OAI22_X1   g1844(.A1(new_n915_), .A2(new_n920_), .B1(new_n1085_), .B2(new_n1080_), .ZN(new_n2230_));
  NOR4_X1    g1845(.A1(new_n1966_), .A2(new_n2054_), .A3(new_n2142_), .A4(new_n2230_), .ZN(new_n2231_));
  NAND4_X1   g1846(.A1(new_n1679_), .A2(new_n2231_), .A3(new_n2225_), .A4(new_n2229_), .ZN(new_n2232_));
  AOI21_X1   g1847(.A1(new_n2232_), .A2(new_n2217_), .B(new_n922_), .ZN(\grant[67] ));
  NOR2_X1    g1848(.A1(new_n1302_), .A2(new_n926_), .ZN(new_n2234_));
  NOR4_X1    g1849(.A1(new_n1317_), .A2(new_n1327_), .A3(new_n1796_), .A4(new_n2234_), .ZN(new_n2235_));
  INV_X1     g1850(.I(\req[69] ), .ZN(new_n2236_));
  AOI21_X1   g1851(.A1(new_n2236_), .A2(\priority[69] ), .B(\priority[70] ), .ZN(new_n2237_));
  OAI21_X1   g1852(.A1(new_n1174_), .A2(new_n1172_), .B(new_n2237_), .ZN(new_n2238_));
  NOR3_X1    g1853(.A1(new_n1801_), .A2(new_n1889_), .A3(new_n2238_), .ZN(new_n2239_));
  OAI22_X1   g1854(.A1(new_n1135_), .A2(new_n1137_), .B1(new_n1191_), .B2(new_n1189_), .ZN(new_n2240_));
  NOR4_X1    g1855(.A1(new_n1976_), .A2(new_n2064_), .A3(new_n2152_), .A4(new_n2240_), .ZN(new_n2241_));
  NAND4_X1   g1856(.A1(new_n1691_), .A2(new_n2241_), .A3(new_n2235_), .A4(new_n2239_), .ZN(new_n2242_));
  AOI21_X1   g1857(.A1(new_n2242_), .A2(new_n2226_), .B(new_n435_), .ZN(\grant[68] ));
  NOR2_X1    g1858(.A1(new_n1380_), .A2(new_n441_), .ZN(new_n2244_));
  NOR4_X1    g1859(.A1(new_n1395_), .A2(new_n1405_), .A3(new_n1806_), .A4(new_n2244_), .ZN(new_n2245_));
  INV_X1     g1860(.I(\req[70] ), .ZN(new_n2246_));
  AOI21_X1   g1861(.A1(new_n2246_), .A2(\priority[70] ), .B(\priority[71] ), .ZN(new_n2247_));
  OAI21_X1   g1862(.A1(new_n1256_), .A2(new_n1254_), .B(new_n2247_), .ZN(new_n2248_));
  NOR3_X1    g1863(.A1(new_n1811_), .A2(new_n1898_), .A3(new_n2248_), .ZN(new_n2249_));
  OAI22_X1   g1864(.A1(new_n1217_), .A2(new_n1219_), .B1(new_n1273_), .B2(new_n1271_), .ZN(new_n2250_));
  NOR4_X1    g1865(.A1(new_n1986_), .A2(new_n2074_), .A3(new_n2162_), .A4(new_n2250_), .ZN(new_n2251_));
  NAND4_X1   g1866(.A1(new_n1703_), .A2(new_n2251_), .A3(new_n2245_), .A4(new_n2249_), .ZN(new_n2252_));
  AOI21_X1   g1867(.A1(new_n2252_), .A2(new_n2236_), .B(new_n681_), .ZN(\grant[69] ));
  NOR2_X1    g1868(.A1(new_n1458_), .A2(new_n687_), .ZN(new_n2254_));
  NOR4_X1    g1869(.A1(new_n1473_), .A2(new_n1483_), .A3(new_n1816_), .A4(new_n2254_), .ZN(new_n2255_));
  INV_X1     g1870(.I(\req[71] ), .ZN(new_n2256_));
  AOI21_X1   g1871(.A1(new_n2256_), .A2(\priority[71] ), .B(\priority[72] ), .ZN(new_n2257_));
  OAI21_X1   g1872(.A1(new_n1335_), .A2(new_n1333_), .B(new_n2257_), .ZN(new_n2258_));
  NOR3_X1    g1873(.A1(new_n1821_), .A2(new_n1907_), .A3(new_n2258_), .ZN(new_n2259_));
  OAI22_X1   g1874(.A1(new_n1299_), .A2(new_n1301_), .B1(new_n1352_), .B2(new_n1350_), .ZN(new_n2260_));
  NOR4_X1    g1875(.A1(new_n1996_), .A2(new_n2084_), .A3(new_n2172_), .A4(new_n2260_), .ZN(new_n2261_));
  NAND4_X1   g1876(.A1(new_n1715_), .A2(new_n2261_), .A3(new_n2255_), .A4(new_n2259_), .ZN(new_n2262_));
  AOI21_X1   g1877(.A1(new_n2262_), .A2(new_n2246_), .B(new_n927_), .ZN(\grant[70] ));
  NOR2_X1    g1878(.A1(new_n1536_), .A2(new_n933_), .ZN(new_n2264_));
  NOR4_X1    g1879(.A1(new_n1551_), .A2(new_n1561_), .A3(new_n1826_), .A4(new_n2264_), .ZN(new_n2265_));
  INV_X1     g1880(.I(\req[72] ), .ZN(new_n2266_));
  AOI21_X1   g1881(.A1(new_n2266_), .A2(\priority[72] ), .B(\priority[73] ), .ZN(new_n2267_));
  OAI21_X1   g1882(.A1(new_n1413_), .A2(new_n1411_), .B(new_n2267_), .ZN(new_n2268_));
  NOR3_X1    g1883(.A1(new_n1831_), .A2(new_n1916_), .A3(new_n2268_), .ZN(new_n2269_));
  OAI22_X1   g1884(.A1(new_n1427_), .A2(new_n1430_), .B1(new_n1379_), .B2(new_n1377_), .ZN(new_n2270_));
  NOR4_X1    g1885(.A1(new_n2006_), .A2(new_n2094_), .A3(new_n2182_), .A4(new_n2270_), .ZN(new_n2271_));
  NAND4_X1   g1886(.A1(new_n1727_), .A2(new_n2271_), .A3(new_n2265_), .A4(new_n2269_), .ZN(new_n2272_));
  AOI21_X1   g1887(.A1(new_n2272_), .A2(new_n2256_), .B(new_n442_), .ZN(\grant[71] ));
  NOR4_X1    g1888(.A1(new_n1498_), .A2(new_n1504_), .A3(new_n1514_), .A4(new_n1519_), .ZN(new_n2274_));
  NOR2_X1    g1889(.A1(new_n453_), .A2(new_n446_), .ZN(new_n2275_));
  OAI22_X1   g1890(.A1(new_n1455_), .A2(new_n1457_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n2276_));
  NOR4_X1    g1891(.A1(new_n1509_), .A2(new_n1837_), .A3(new_n2276_), .A4(new_n2275_), .ZN(new_n2277_));
  INV_X1     g1892(.I(\req[73] ), .ZN(new_n2278_));
  AOI21_X1   g1893(.A1(new_n2278_), .A2(\priority[73] ), .B(\priority[74] ), .ZN(new_n2279_));
  OAI21_X1   g1894(.A1(new_n394_), .A2(new_n389_), .B(new_n2279_), .ZN(new_n2280_));
  NOR3_X1    g1895(.A1(new_n1601_), .A2(new_n1604_), .A3(new_n2280_), .ZN(new_n2281_));
  NAND4_X1   g1896(.A1(new_n1920_), .A2(new_n2274_), .A3(new_n2277_), .A4(new_n2281_), .ZN(new_n2282_));
  AOI21_X1   g1897(.A1(new_n2282_), .A2(new_n2266_), .B(new_n688_), .ZN(\grant[72] ));
  NOR4_X1    g1898(.A1(new_n1576_), .A2(new_n1582_), .A3(new_n1592_), .A4(new_n1597_), .ZN(new_n2284_));
  NOR2_X1    g1899(.A1(new_n699_), .A2(new_n692_), .ZN(new_n2285_));
  OAI22_X1   g1900(.A1(new_n1533_), .A2(new_n1535_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n2286_));
  NOR4_X1    g1901(.A1(new_n1587_), .A2(new_n1849_), .A3(new_n2286_), .A4(new_n2285_), .ZN(new_n2287_));
  INV_X1     g1902(.I(\req[74] ), .ZN(new_n2288_));
  AOI21_X1   g1903(.A1(new_n2288_), .A2(\priority[74] ), .B(\priority[75] ), .ZN(new_n2289_));
  OAI21_X1   g1904(.A1(new_n640_), .A2(new_n635_), .B(new_n2289_), .ZN(new_n2290_));
  NOR3_X1    g1905(.A1(new_n1628_), .A2(new_n1631_), .A3(new_n2290_), .ZN(new_n2291_));
  NAND4_X1   g1906(.A1(new_n1931_), .A2(new_n2284_), .A3(new_n2287_), .A4(new_n2291_), .ZN(new_n2292_));
  AOI21_X1   g1907(.A1(new_n2292_), .A2(new_n2278_), .B(new_n934_), .ZN(\grant[73] ));
  NOR4_X1    g1908(.A1(new_n895_), .A2(new_n912_), .A3(new_n990_), .A4(new_n1622_), .ZN(new_n2294_));
  NOR2_X1    g1909(.A1(new_n945_), .A2(new_n938_), .ZN(new_n2295_));
  NOR4_X1    g1910(.A1(new_n973_), .A2(new_n1007_), .A3(new_n1766_), .A4(new_n2295_), .ZN(new_n2296_));
  INV_X1     g1911(.I(\req[75] ), .ZN(new_n2297_));
  AOI21_X1   g1912(.A1(new_n2297_), .A2(\priority[75] ), .B(\priority[76] ), .ZN(new_n2298_));
  OAI21_X1   g1913(.A1(new_n533_), .A2(new_n528_), .B(new_n2298_), .ZN(new_n2299_));
  NOR3_X1    g1914(.A1(new_n1618_), .A2(new_n1771_), .A3(new_n2299_), .ZN(new_n2300_));
  NAND4_X1   g1915(.A1(new_n2212_), .A2(new_n2294_), .A3(new_n2296_), .A4(new_n2300_), .ZN(new_n2301_));
  AOI21_X1   g1916(.A1(new_n2301_), .A2(new_n2288_), .B(new_n447_), .ZN(\grant[74] ));
  NOR4_X1    g1917(.A1(new_n1129_), .A2(new_n1134_), .A3(new_n1161_), .A4(new_n1649_), .ZN(new_n2303_));
  NOR2_X1    g1918(.A1(new_n1143_), .A2(new_n451_), .ZN(new_n2304_));
  NOR4_X1    g1919(.A1(new_n1156_), .A2(new_n1166_), .A3(new_n1776_), .A4(new_n2304_), .ZN(new_n2305_));
  INV_X1     g1920(.I(\req[76] ), .ZN(new_n2306_));
  AOI21_X1   g1921(.A1(new_n2306_), .A2(\priority[76] ), .B(\priority[77] ), .ZN(new_n2307_));
  OAI21_X1   g1922(.A1(new_n779_), .A2(new_n774_), .B(new_n2307_), .ZN(new_n2308_));
  NOR3_X1    g1923(.A1(new_n1645_), .A2(new_n1781_), .A3(new_n2308_), .ZN(new_n2309_));
  NAND4_X1   g1924(.A1(new_n2221_), .A2(new_n2303_), .A3(new_n2305_), .A4(new_n2309_), .ZN(new_n2310_));
  AOI21_X1   g1925(.A1(new_n2310_), .A2(new_n2297_), .B(new_n693_), .ZN(\grant[75] ));
  OAI22_X1   g1926(.A1(new_n923_), .A2(new_n928_), .B1(new_n937_), .B2(new_n932_), .ZN(new_n2312_));
  NOR4_X1    g1927(.A1(new_n1211_), .A2(new_n1216_), .A3(new_n1243_), .A4(new_n2312_), .ZN(new_n2313_));
  NOR2_X1    g1928(.A1(new_n1225_), .A2(new_n697_), .ZN(new_n2314_));
  NOR4_X1    g1929(.A1(new_n1238_), .A2(new_n1248_), .A3(new_n1786_), .A4(new_n2314_), .ZN(new_n2315_));
  INV_X1     g1930(.I(\req[77] ), .ZN(new_n2316_));
  AOI21_X1   g1931(.A1(new_n2316_), .A2(\priority[77] ), .B(\priority[78] ), .ZN(new_n2317_));
  OAI21_X1   g1932(.A1(new_n1025_), .A2(new_n1020_), .B(new_n2317_), .ZN(new_n2318_));
  NOR3_X1    g1933(.A1(new_n1791_), .A2(new_n1880_), .A3(new_n2318_), .ZN(new_n2319_));
  NAND4_X1   g1934(.A1(new_n2231_), .A2(new_n2313_), .A3(new_n2315_), .A4(new_n2319_), .ZN(new_n2320_));
  AOI21_X1   g1935(.A1(new_n2320_), .A2(new_n2306_), .B(new_n939_), .ZN(\grant[76] ));
  OAI22_X1   g1936(.A1(new_n1136_), .A2(new_n1138_), .B1(new_n1142_), .B2(new_n1140_), .ZN(new_n2322_));
  NOR4_X1    g1937(.A1(new_n1293_), .A2(new_n1298_), .A3(new_n1322_), .A4(new_n2322_), .ZN(new_n2323_));
  NOR2_X1    g1938(.A1(new_n1307_), .A2(new_n943_), .ZN(new_n2324_));
  NOR4_X1    g1939(.A1(new_n1317_), .A2(new_n1327_), .A3(new_n1796_), .A4(new_n2324_), .ZN(new_n2325_));
  INV_X1     g1940(.I(\req[78] ), .ZN(new_n2326_));
  AOI21_X1   g1941(.A1(new_n2326_), .A2(\priority[78] ), .B(\priority[79] ), .ZN(new_n2327_));
  OAI21_X1   g1942(.A1(new_n1174_), .A2(new_n1172_), .B(new_n2327_), .ZN(new_n2328_));
  NOR3_X1    g1943(.A1(new_n1801_), .A2(new_n1889_), .A3(new_n2328_), .ZN(new_n2329_));
  NAND4_X1   g1944(.A1(new_n2241_), .A2(new_n2323_), .A3(new_n2325_), .A4(new_n2329_), .ZN(new_n2330_));
  AOI21_X1   g1945(.A1(new_n2330_), .A2(new_n2316_), .B(new_n452_), .ZN(\grant[77] ));
  OAI22_X1   g1946(.A1(new_n1218_), .A2(new_n1220_), .B1(new_n1224_), .B2(new_n1222_), .ZN(new_n2332_));
  NOR4_X1    g1947(.A1(new_n1371_), .A2(new_n1376_), .A3(new_n1400_), .A4(new_n2332_), .ZN(new_n2333_));
  NOR2_X1    g1948(.A1(new_n1385_), .A2(new_n390_), .ZN(new_n2334_));
  NOR4_X1    g1949(.A1(new_n1395_), .A2(new_n1405_), .A3(new_n1806_), .A4(new_n2334_), .ZN(new_n2335_));
  INV_X1     g1950(.I(\req[79] ), .ZN(new_n2336_));
  AOI21_X1   g1951(.A1(new_n2336_), .A2(\priority[79] ), .B(\priority[80] ), .ZN(new_n2337_));
  OAI21_X1   g1952(.A1(new_n1256_), .A2(new_n1254_), .B(new_n2337_), .ZN(new_n2338_));
  NOR3_X1    g1953(.A1(new_n1811_), .A2(new_n1898_), .A3(new_n2338_), .ZN(new_n2339_));
  NAND4_X1   g1954(.A1(new_n2251_), .A2(new_n2333_), .A3(new_n2335_), .A4(new_n2339_), .ZN(new_n2340_));
  AOI21_X1   g1955(.A1(new_n2340_), .A2(new_n2326_), .B(new_n698_), .ZN(\grant[78] ));
  OAI22_X1   g1956(.A1(new_n1300_), .A2(new_n1302_), .B1(new_n1306_), .B2(new_n1304_), .ZN(new_n2342_));
  NOR4_X1    g1957(.A1(new_n1449_), .A2(new_n1454_), .A3(new_n1478_), .A4(new_n2342_), .ZN(new_n2343_));
  NOR2_X1    g1958(.A1(new_n1463_), .A2(new_n636_), .ZN(new_n2344_));
  NOR4_X1    g1959(.A1(new_n1473_), .A2(new_n1483_), .A3(new_n1816_), .A4(new_n2344_), .ZN(new_n2345_));
  INV_X1     g1960(.I(\req[80] ), .ZN(new_n2346_));
  AOI21_X1   g1961(.A1(new_n2346_), .A2(\priority[80] ), .B(\priority[81] ), .ZN(new_n2347_));
  OAI21_X1   g1962(.A1(new_n1335_), .A2(new_n1333_), .B(new_n2347_), .ZN(new_n2348_));
  NOR3_X1    g1963(.A1(new_n1821_), .A2(new_n1907_), .A3(new_n2348_), .ZN(new_n2349_));
  NAND4_X1   g1964(.A1(new_n2261_), .A2(new_n2343_), .A3(new_n2345_), .A4(new_n2349_), .ZN(new_n2350_));
  AOI21_X1   g1965(.A1(new_n2350_), .A2(new_n2336_), .B(new_n944_), .ZN(\grant[79] ));
  OAI22_X1   g1966(.A1(new_n1378_), .A2(new_n1380_), .B1(new_n1384_), .B2(new_n1383_), .ZN(new_n2352_));
  NOR4_X1    g1967(.A1(new_n1527_), .A2(new_n1532_), .A3(new_n1556_), .A4(new_n2352_), .ZN(new_n2353_));
  NOR2_X1    g1968(.A1(new_n1541_), .A2(new_n882_), .ZN(new_n2354_));
  NOR4_X1    g1969(.A1(new_n1551_), .A2(new_n1561_), .A3(new_n1826_), .A4(new_n2354_), .ZN(new_n2355_));
  INV_X1     g1970(.I(\req[81] ), .ZN(new_n2356_));
  AOI21_X1   g1971(.A1(new_n2356_), .A2(\priority[81] ), .B(\priority[82] ), .ZN(new_n2357_));
  OAI21_X1   g1972(.A1(new_n1413_), .A2(new_n1411_), .B(new_n2357_), .ZN(new_n2358_));
  NOR3_X1    g1973(.A1(new_n1831_), .A2(new_n1916_), .A3(new_n2358_), .ZN(new_n2359_));
  NAND4_X1   g1974(.A1(new_n2271_), .A2(new_n2353_), .A3(new_n2355_), .A4(new_n2359_), .ZN(new_n2360_));
  AOI21_X1   g1975(.A1(new_n2360_), .A2(new_n2346_), .B(new_n391_), .ZN(\grant[80] ));
  NOR2_X1    g1976(.A1(new_n402_), .A2(new_n395_), .ZN(new_n2362_));
  OAI22_X1   g1977(.A1(new_n1461_), .A2(new_n1462_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n2363_));
  NOR4_X1    g1978(.A1(new_n1459_), .A2(new_n1837_), .A3(new_n2363_), .A4(new_n2362_), .ZN(new_n2364_));
  INV_X1     g1979(.I(\req[82] ), .ZN(new_n2365_));
  AOI21_X1   g1980(.A1(new_n2365_), .A2(\priority[82] ), .B(\priority[83] ), .ZN(new_n2366_));
  OAI21_X1   g1981(.A1(new_n411_), .A2(new_n406_), .B(new_n2366_), .ZN(new_n2367_));
  NOR3_X1    g1982(.A1(new_n1601_), .A2(new_n1602_), .A3(new_n2367_), .ZN(new_n2368_));
  NAND4_X1   g1983(.A1(new_n1520_), .A2(new_n2010_), .A3(new_n2364_), .A4(new_n2368_), .ZN(new_n2369_));
  AOI21_X1   g1984(.A1(new_n2369_), .A2(new_n2356_), .B(new_n637_), .ZN(\grant[81] ));
  NOR2_X1    g1985(.A1(new_n648_), .A2(new_n641_), .ZN(new_n2371_));
  OAI22_X1   g1986(.A1(new_n1539_), .A2(new_n1540_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n2372_));
  NOR4_X1    g1987(.A1(new_n1537_), .A2(new_n1849_), .A3(new_n2372_), .A4(new_n2371_), .ZN(new_n2373_));
  INV_X1     g1988(.I(\req[83] ), .ZN(new_n2374_));
  AOI21_X1   g1989(.A1(new_n2374_), .A2(\priority[83] ), .B(\priority[84] ), .ZN(new_n2375_));
  OAI21_X1   g1990(.A1(new_n657_), .A2(new_n652_), .B(new_n2375_), .ZN(new_n2376_));
  NOR3_X1    g1991(.A1(new_n1628_), .A2(new_n1629_), .A3(new_n2376_), .ZN(new_n2377_));
  NAND4_X1   g1992(.A1(new_n1598_), .A2(new_n2020_), .A3(new_n2373_), .A4(new_n2377_), .ZN(new_n2378_));
  AOI21_X1   g1993(.A1(new_n2378_), .A2(new_n2365_), .B(new_n883_), .ZN(\grant[82] ));
  NOR4_X1    g1994(.A1(new_n912_), .A2(new_n990_), .A3(new_n1603_), .A4(new_n1622_), .ZN(new_n2380_));
  NOR2_X1    g1995(.A1(new_n894_), .A2(new_n887_), .ZN(new_n2381_));
  NOR4_X1    g1996(.A1(new_n973_), .A2(new_n1007_), .A3(new_n1766_), .A4(new_n2381_), .ZN(new_n2382_));
  INV_X1     g1997(.I(\req[84] ), .ZN(new_n2383_));
  AOI21_X1   g1998(.A1(new_n2383_), .A2(\priority[84] ), .B(\priority[85] ), .ZN(new_n2384_));
  OAI21_X1   g1999(.A1(new_n533_), .A2(new_n528_), .B(new_n2384_), .ZN(new_n2385_));
  NOR3_X1    g2000(.A1(new_n1618_), .A2(new_n1771_), .A3(new_n2385_), .ZN(new_n2386_));
  NAND4_X1   g2001(.A1(new_n2212_), .A2(new_n2380_), .A3(new_n2382_), .A4(new_n2386_), .ZN(new_n2387_));
  AOI21_X1   g2002(.A1(new_n2387_), .A2(new_n2374_), .B(new_n396_), .ZN(\grant[83] ));
  NOR4_X1    g2003(.A1(new_n1134_), .A2(new_n1161_), .A3(new_n1630_), .A4(new_n1649_), .ZN(new_n2389_));
  NOR2_X1    g2004(.A1(new_n1128_), .A2(new_n400_), .ZN(new_n2390_));
  NOR4_X1    g2005(.A1(new_n1156_), .A2(new_n1166_), .A3(new_n1776_), .A4(new_n2390_), .ZN(new_n2391_));
  INV_X1     g2006(.I(\req[85] ), .ZN(new_n2392_));
  AOI21_X1   g2007(.A1(new_n2392_), .A2(\priority[85] ), .B(\priority[86] ), .ZN(new_n2393_));
  OAI21_X1   g2008(.A1(new_n779_), .A2(new_n774_), .B(new_n2393_), .ZN(new_n2394_));
  NOR3_X1    g2009(.A1(new_n1645_), .A2(new_n1781_), .A3(new_n2394_), .ZN(new_n2395_));
  NAND4_X1   g2010(.A1(new_n2221_), .A2(new_n2389_), .A3(new_n2391_), .A4(new_n2395_), .ZN(new_n2396_));
  AOI21_X1   g2011(.A1(new_n2396_), .A2(new_n2383_), .B(new_n642_), .ZN(\grant[84] ));
  OAI22_X1   g2012(.A1(new_n881_), .A2(new_n886_), .B1(new_n945_), .B2(new_n940_), .ZN(new_n2398_));
  NOR4_X1    g2013(.A1(new_n1216_), .A2(new_n1243_), .A3(new_n2312_), .A4(new_n2398_), .ZN(new_n2399_));
  NOR2_X1    g2014(.A1(new_n1210_), .A2(new_n646_), .ZN(new_n2400_));
  NOR4_X1    g2015(.A1(new_n1238_), .A2(new_n1248_), .A3(new_n1786_), .A4(new_n2400_), .ZN(new_n2401_));
  INV_X1     g2016(.I(\req[86] ), .ZN(new_n2402_));
  AOI21_X1   g2017(.A1(new_n2402_), .A2(\priority[86] ), .B(\priority[87] ), .ZN(new_n2403_));
  OAI21_X1   g2018(.A1(new_n1025_), .A2(new_n1020_), .B(new_n2403_), .ZN(new_n2404_));
  NOR3_X1    g2019(.A1(new_n1791_), .A2(new_n1880_), .A3(new_n2404_), .ZN(new_n2405_));
  NAND4_X1   g2020(.A1(new_n2231_), .A2(new_n2399_), .A3(new_n2401_), .A4(new_n2405_), .ZN(new_n2406_));
  AOI21_X1   g2021(.A1(new_n2406_), .A2(new_n2392_), .B(new_n888_), .ZN(\grant[85] ));
  OAI22_X1   g2022(.A1(new_n1125_), .A2(new_n1127_), .B1(new_n1143_), .B2(new_n1141_), .ZN(new_n2408_));
  NOR4_X1    g2023(.A1(new_n1298_), .A2(new_n1322_), .A3(new_n2322_), .A4(new_n2408_), .ZN(new_n2409_));
  NOR2_X1    g2024(.A1(new_n1292_), .A2(new_n892_), .ZN(new_n2410_));
  NOR4_X1    g2025(.A1(new_n1317_), .A2(new_n1327_), .A3(new_n1796_), .A4(new_n2410_), .ZN(new_n2411_));
  INV_X1     g2026(.I(\req[87] ), .ZN(new_n2412_));
  AOI21_X1   g2027(.A1(new_n2412_), .A2(\priority[87] ), .B(\priority[88] ), .ZN(new_n2413_));
  OAI21_X1   g2028(.A1(new_n1174_), .A2(new_n1172_), .B(new_n2413_), .ZN(new_n2414_));
  NOR3_X1    g2029(.A1(new_n1801_), .A2(new_n1889_), .A3(new_n2414_), .ZN(new_n2415_));
  NAND4_X1   g2030(.A1(new_n2241_), .A2(new_n2409_), .A3(new_n2411_), .A4(new_n2415_), .ZN(new_n2416_));
  AOI21_X1   g2031(.A1(new_n2416_), .A2(new_n2402_), .B(new_n401_), .ZN(\grant[86] ));
  OAI22_X1   g2032(.A1(new_n1207_), .A2(new_n1209_), .B1(new_n1225_), .B2(new_n1223_), .ZN(new_n2418_));
  NOR4_X1    g2033(.A1(new_n1376_), .A2(new_n1400_), .A3(new_n2332_), .A4(new_n2418_), .ZN(new_n2419_));
  NOR2_X1    g2034(.A1(new_n1370_), .A2(new_n407_), .ZN(new_n2420_));
  NOR4_X1    g2035(.A1(new_n1395_), .A2(new_n1405_), .A3(new_n1806_), .A4(new_n2420_), .ZN(new_n2421_));
  INV_X1     g2036(.I(\req[88] ), .ZN(new_n2422_));
  AOI21_X1   g2037(.A1(new_n2422_), .A2(\priority[88] ), .B(\priority[89] ), .ZN(new_n2423_));
  OAI21_X1   g2038(.A1(new_n1256_), .A2(new_n1254_), .B(new_n2423_), .ZN(new_n2424_));
  NOR3_X1    g2039(.A1(new_n1811_), .A2(new_n1898_), .A3(new_n2424_), .ZN(new_n2425_));
  NAND4_X1   g2040(.A1(new_n2251_), .A2(new_n2419_), .A3(new_n2421_), .A4(new_n2425_), .ZN(new_n2426_));
  AOI21_X1   g2041(.A1(new_n2426_), .A2(new_n2412_), .B(new_n647_), .ZN(\grant[87] ));
  OAI22_X1   g2042(.A1(new_n1289_), .A2(new_n1291_), .B1(new_n1307_), .B2(new_n1305_), .ZN(new_n2428_));
  NOR4_X1    g2043(.A1(new_n1454_), .A2(new_n1478_), .A3(new_n2342_), .A4(new_n2428_), .ZN(new_n2429_));
  NOR2_X1    g2044(.A1(new_n1448_), .A2(new_n653_), .ZN(new_n2430_));
  NOR4_X1    g2045(.A1(new_n1473_), .A2(new_n1483_), .A3(new_n1816_), .A4(new_n2430_), .ZN(new_n2431_));
  INV_X1     g2046(.I(\req[89] ), .ZN(new_n2432_));
  AOI21_X1   g2047(.A1(new_n2432_), .A2(\priority[89] ), .B(\priority[90] ), .ZN(new_n2433_));
  OAI21_X1   g2048(.A1(new_n1335_), .A2(new_n1333_), .B(new_n2433_), .ZN(new_n2434_));
  NOR3_X1    g2049(.A1(new_n1821_), .A2(new_n1907_), .A3(new_n2434_), .ZN(new_n2435_));
  NAND4_X1   g2050(.A1(new_n2261_), .A2(new_n2429_), .A3(new_n2431_), .A4(new_n2435_), .ZN(new_n2436_));
  AOI21_X1   g2051(.A1(new_n2436_), .A2(new_n2422_), .B(new_n893_), .ZN(\grant[88] ));
  OAI22_X1   g2052(.A1(new_n1382_), .A2(new_n1385_), .B1(new_n1369_), .B2(new_n1367_), .ZN(new_n2438_));
  NOR4_X1    g2053(.A1(new_n1532_), .A2(new_n1556_), .A3(new_n2352_), .A4(new_n2438_), .ZN(new_n2439_));
  NOR2_X1    g2054(.A1(new_n1526_), .A2(new_n899_), .ZN(new_n2440_));
  NOR4_X1    g2055(.A1(new_n1551_), .A2(new_n1561_), .A3(new_n1826_), .A4(new_n2440_), .ZN(new_n2441_));
  INV_X1     g2056(.I(\req[90] ), .ZN(new_n2442_));
  AOI21_X1   g2057(.A1(new_n2442_), .A2(\priority[90] ), .B(\priority[91] ), .ZN(new_n2443_));
  OAI21_X1   g2058(.A1(new_n1413_), .A2(new_n1411_), .B(new_n2443_), .ZN(new_n2444_));
  NOR3_X1    g2059(.A1(new_n1831_), .A2(new_n1916_), .A3(new_n2444_), .ZN(new_n2445_));
  NAND4_X1   g2060(.A1(new_n2271_), .A2(new_n2439_), .A3(new_n2441_), .A4(new_n2445_), .ZN(new_n2446_));
  AOI21_X1   g2061(.A1(new_n2446_), .A2(new_n2432_), .B(new_n408_), .ZN(\grant[89] ));
  NOR2_X1    g2062(.A1(new_n419_), .A2(new_n412_), .ZN(new_n2448_));
  OAI22_X1   g2063(.A1(new_n1445_), .A2(new_n1447_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n2449_));
  NOR4_X1    g2064(.A1(new_n1464_), .A2(new_n1837_), .A3(new_n2449_), .A4(new_n2448_), .ZN(new_n2450_));
  INV_X1     g2065(.I(\req[91] ), .ZN(new_n2451_));
  AOI21_X1   g2066(.A1(new_n2451_), .A2(\priority[91] ), .B(\priority[92] ), .ZN(new_n2452_));
  OAI21_X1   g2067(.A1(new_n489_), .A2(new_n484_), .B(new_n2452_), .ZN(new_n2453_));
  NOR3_X1    g2068(.A1(new_n1602_), .A2(new_n1612_), .A3(new_n2453_), .ZN(new_n2454_));
  NAND4_X1   g2069(.A1(new_n1724_), .A2(new_n2098_), .A3(new_n2450_), .A4(new_n2454_), .ZN(new_n2455_));
  AOI21_X1   g2070(.A1(new_n2455_), .A2(new_n2442_), .B(new_n654_), .ZN(\grant[90] ));
  NOR2_X1    g2071(.A1(new_n665_), .A2(new_n658_), .ZN(new_n2457_));
  OAI22_X1   g2072(.A1(new_n1523_), .A2(new_n1525_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n2458_));
  NOR4_X1    g2073(.A1(new_n1542_), .A2(new_n1849_), .A3(new_n2458_), .A4(new_n2457_), .ZN(new_n2459_));
  INV_X1     g2074(.I(\req[92] ), .ZN(new_n2460_));
  AOI21_X1   g2075(.A1(new_n2460_), .A2(\priority[92] ), .B(\priority[93] ), .ZN(new_n2461_));
  OAI21_X1   g2076(.A1(new_n735_), .A2(new_n730_), .B(new_n2461_), .ZN(new_n2462_));
  NOR3_X1    g2077(.A1(new_n1629_), .A2(new_n1639_), .A3(new_n2462_), .ZN(new_n2463_));
  NAND4_X1   g2078(.A1(new_n1736_), .A2(new_n2108_), .A3(new_n2459_), .A4(new_n2463_), .ZN(new_n2464_));
  AOI21_X1   g2079(.A1(new_n2464_), .A2(new_n2451_), .B(new_n900_), .ZN(\grant[91] ));
  NOR4_X1    g2080(.A1(new_n990_), .A2(new_n1603_), .A3(new_n1604_), .A4(new_n1622_), .ZN(new_n2466_));
  NOR2_X1    g2081(.A1(new_n911_), .A2(new_n904_), .ZN(new_n2467_));
  NOR4_X1    g2082(.A1(new_n973_), .A2(new_n1007_), .A3(new_n1766_), .A4(new_n2467_), .ZN(new_n2468_));
  INV_X1     g2083(.I(\req[93] ), .ZN(new_n2469_));
  AOI21_X1   g2084(.A1(new_n2469_), .A2(\priority[93] ), .B(\priority[94] ), .ZN(new_n2470_));
  OAI21_X1   g2085(.A1(new_n533_), .A2(new_n528_), .B(new_n2470_), .ZN(new_n2471_));
  NOR3_X1    g2086(.A1(new_n1618_), .A2(new_n1771_), .A3(new_n2471_), .ZN(new_n2472_));
  NAND4_X1   g2087(.A1(new_n2212_), .A2(new_n2466_), .A3(new_n2468_), .A4(new_n2472_), .ZN(new_n2473_));
  AOI21_X1   g2088(.A1(new_n2473_), .A2(new_n2460_), .B(new_n413_), .ZN(\grant[92] ));
  NOR4_X1    g2089(.A1(new_n1161_), .A2(new_n1630_), .A3(new_n1631_), .A4(new_n1649_), .ZN(new_n2475_));
  NOR2_X1    g2090(.A1(new_n1133_), .A2(new_n417_), .ZN(new_n2476_));
  NOR4_X1    g2091(.A1(new_n1156_), .A2(new_n1166_), .A3(new_n1776_), .A4(new_n2476_), .ZN(new_n2477_));
  INV_X1     g2092(.I(\req[94] ), .ZN(new_n2478_));
  AOI21_X1   g2093(.A1(new_n2478_), .A2(\priority[94] ), .B(\priority[95] ), .ZN(new_n2479_));
  OAI21_X1   g2094(.A1(new_n779_), .A2(new_n774_), .B(new_n2479_), .ZN(new_n2480_));
  NOR3_X1    g2095(.A1(new_n1645_), .A2(new_n1781_), .A3(new_n2480_), .ZN(new_n2481_));
  NAND4_X1   g2096(.A1(new_n2221_), .A2(new_n2475_), .A3(new_n2477_), .A4(new_n2481_), .ZN(new_n2482_));
  AOI21_X1   g2097(.A1(new_n2482_), .A2(new_n2469_), .B(new_n659_), .ZN(\grant[93] ));
  OAI22_X1   g2098(.A1(new_n889_), .A2(new_n894_), .B1(new_n903_), .B2(new_n898_), .ZN(new_n2484_));
  NOR4_X1    g2099(.A1(new_n1243_), .A2(new_n2312_), .A3(new_n2398_), .A4(new_n2484_), .ZN(new_n2485_));
  NOR2_X1    g2100(.A1(new_n1215_), .A2(new_n663_), .ZN(new_n2486_));
  NOR4_X1    g2101(.A1(new_n1238_), .A2(new_n1248_), .A3(new_n1786_), .A4(new_n2486_), .ZN(new_n2487_));
  INV_X1     g2102(.I(\req[95] ), .ZN(new_n2488_));
  AOI21_X1   g2103(.A1(new_n2488_), .A2(\priority[95] ), .B(\priority[96] ), .ZN(new_n2489_));
  OAI21_X1   g2104(.A1(new_n1025_), .A2(new_n1020_), .B(new_n2489_), .ZN(new_n2490_));
  NOR3_X1    g2105(.A1(new_n1791_), .A2(new_n1880_), .A3(new_n2490_), .ZN(new_n2491_));
  NAND4_X1   g2106(.A1(new_n2231_), .A2(new_n2485_), .A3(new_n2487_), .A4(new_n2491_), .ZN(new_n2492_));
  AOI21_X1   g2107(.A1(new_n2492_), .A2(new_n2478_), .B(new_n905_), .ZN(\grant[94] ));
  OAI22_X1   g2108(.A1(new_n1126_), .A2(new_n1128_), .B1(new_n1132_), .B2(new_n1130_), .ZN(new_n2494_));
  NOR4_X1    g2109(.A1(new_n1322_), .A2(new_n2322_), .A3(new_n2408_), .A4(new_n2494_), .ZN(new_n2495_));
  NOR2_X1    g2110(.A1(new_n1297_), .A2(new_n909_), .ZN(new_n2496_));
  NOR4_X1    g2111(.A1(new_n1317_), .A2(new_n1327_), .A3(new_n1796_), .A4(new_n2496_), .ZN(new_n2497_));
  INV_X1     g2112(.I(\req[96] ), .ZN(new_n2498_));
  AOI21_X1   g2113(.A1(new_n2498_), .A2(\priority[96] ), .B(\priority[97] ), .ZN(new_n2499_));
  OAI21_X1   g2114(.A1(new_n1174_), .A2(new_n1172_), .B(new_n2499_), .ZN(new_n2500_));
  NOR3_X1    g2115(.A1(new_n1801_), .A2(new_n1889_), .A3(new_n2500_), .ZN(new_n2501_));
  NAND4_X1   g2116(.A1(new_n2241_), .A2(new_n2495_), .A3(new_n2497_), .A4(new_n2501_), .ZN(new_n2502_));
  AOI21_X1   g2117(.A1(new_n2502_), .A2(new_n2488_), .B(new_n418_), .ZN(\grant[95] ));
  OAI22_X1   g2118(.A1(new_n1208_), .A2(new_n1210_), .B1(new_n1214_), .B2(new_n1212_), .ZN(new_n2504_));
  NOR4_X1    g2119(.A1(new_n1400_), .A2(new_n2332_), .A3(new_n2418_), .A4(new_n2504_), .ZN(new_n2505_));
  NOR2_X1    g2120(.A1(new_n1375_), .A2(new_n485_), .ZN(new_n2506_));
  NOR4_X1    g2121(.A1(new_n1395_), .A2(new_n1405_), .A3(new_n1806_), .A4(new_n2506_), .ZN(new_n2507_));
  INV_X1     g2122(.I(\req[97] ), .ZN(new_n2508_));
  AOI21_X1   g2123(.A1(new_n2508_), .A2(\priority[97] ), .B(\priority[98] ), .ZN(new_n2509_));
  OAI21_X1   g2124(.A1(new_n1256_), .A2(new_n1254_), .B(new_n2509_), .ZN(new_n2510_));
  NOR3_X1    g2125(.A1(new_n1811_), .A2(new_n1898_), .A3(new_n2510_), .ZN(new_n2511_));
  NAND4_X1   g2126(.A1(new_n2251_), .A2(new_n2505_), .A3(new_n2507_), .A4(new_n2511_), .ZN(new_n2512_));
  AOI21_X1   g2127(.A1(new_n2512_), .A2(new_n2498_), .B(new_n664_), .ZN(\grant[96] ));
  OAI22_X1   g2128(.A1(new_n1290_), .A2(new_n1292_), .B1(new_n1296_), .B2(new_n1294_), .ZN(new_n2514_));
  NOR4_X1    g2129(.A1(new_n1478_), .A2(new_n2342_), .A3(new_n2428_), .A4(new_n2514_), .ZN(new_n2515_));
  NOR2_X1    g2130(.A1(new_n1453_), .A2(new_n731_), .ZN(new_n2516_));
  NOR4_X1    g2131(.A1(new_n1473_), .A2(new_n1483_), .A3(new_n1816_), .A4(new_n2516_), .ZN(new_n2517_));
  INV_X1     g2132(.I(\req[98] ), .ZN(new_n2518_));
  AOI21_X1   g2133(.A1(new_n2518_), .A2(\priority[98] ), .B(\priority[99] ), .ZN(new_n2519_));
  OAI21_X1   g2134(.A1(new_n1335_), .A2(new_n1333_), .B(new_n2519_), .ZN(new_n2520_));
  NOR3_X1    g2135(.A1(new_n1821_), .A2(new_n1907_), .A3(new_n2520_), .ZN(new_n2521_));
  NAND4_X1   g2136(.A1(new_n2261_), .A2(new_n2515_), .A3(new_n2517_), .A4(new_n2521_), .ZN(new_n2522_));
  AOI21_X1   g2137(.A1(new_n2522_), .A2(new_n2508_), .B(new_n910_), .ZN(\grant[97] ));
  OAI22_X1   g2138(.A1(new_n1368_), .A2(new_n1370_), .B1(new_n1374_), .B2(new_n1372_), .ZN(new_n2524_));
  NOR4_X1    g2139(.A1(new_n1556_), .A2(new_n2352_), .A3(new_n2438_), .A4(new_n2524_), .ZN(new_n2525_));
  NOR2_X1    g2140(.A1(new_n1531_), .A2(new_n977_), .ZN(new_n2526_));
  NOR4_X1    g2141(.A1(new_n1551_), .A2(new_n1561_), .A3(new_n1826_), .A4(new_n2526_), .ZN(new_n2527_));
  INV_X1     g2142(.I(\req[99] ), .ZN(new_n2528_));
  AOI21_X1   g2143(.A1(new_n2528_), .A2(\priority[99] ), .B(\priority[100] ), .ZN(new_n2529_));
  OAI21_X1   g2144(.A1(new_n1413_), .A2(new_n1411_), .B(new_n2529_), .ZN(new_n2530_));
  NOR3_X1    g2145(.A1(new_n1831_), .A2(new_n1916_), .A3(new_n2530_), .ZN(new_n2531_));
  NAND4_X1   g2146(.A1(new_n2271_), .A2(new_n2525_), .A3(new_n2527_), .A4(new_n2531_), .ZN(new_n2532_));
  AOI21_X1   g2147(.A1(new_n2532_), .A2(new_n2518_), .B(new_n486_), .ZN(\grant[98] ));
  NOR4_X1    g2148(.A1(new_n1459_), .A2(new_n1464_), .A3(new_n1504_), .A4(new_n1509_), .ZN(new_n2534_));
  NOR2_X1    g2149(.A1(new_n497_), .A2(new_n490_), .ZN(new_n2535_));
  OAI22_X1   g2150(.A1(new_n1450_), .A2(new_n1452_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n2536_));
  NOR4_X1    g2151(.A1(new_n1449_), .A2(new_n1837_), .A3(new_n2536_), .A4(new_n2535_), .ZN(new_n2537_));
  INV_X1     g2152(.I(\req[100] ), .ZN(new_n2538_));
  AOI21_X1   g2153(.A1(new_n2538_), .A2(\priority[100] ), .B(\priority[101] ), .ZN(new_n2539_));
  OAI21_X1   g2154(.A1(new_n506_), .A2(new_n501_), .B(new_n2539_), .ZN(new_n2540_));
  NOR3_X1    g2155(.A1(new_n1612_), .A2(new_n1613_), .A3(new_n2540_), .ZN(new_n2541_));
  NAND4_X1   g2156(.A1(new_n2186_), .A2(new_n2534_), .A3(new_n2537_), .A4(new_n2541_), .ZN(new_n2542_));
  AOI21_X1   g2157(.A1(new_n2542_), .A2(new_n2528_), .B(new_n732_), .ZN(\grant[99] ));
  NOR4_X1    g2158(.A1(new_n1537_), .A2(new_n1542_), .A3(new_n1582_), .A4(new_n1587_), .ZN(new_n2544_));
  NOR2_X1    g2159(.A1(new_n743_), .A2(new_n736_), .ZN(new_n2545_));
  OAI22_X1   g2160(.A1(new_n1528_), .A2(new_n1530_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n2546_));
  NOR4_X1    g2161(.A1(new_n1527_), .A2(new_n1849_), .A3(new_n2546_), .A4(new_n2545_), .ZN(new_n2547_));
  INV_X1     g2162(.I(\req[101] ), .ZN(new_n2548_));
  AOI21_X1   g2163(.A1(new_n2548_), .A2(\priority[101] ), .B(\priority[102] ), .ZN(new_n2549_));
  OAI21_X1   g2164(.A1(new_n752_), .A2(new_n747_), .B(new_n2549_), .ZN(new_n2550_));
  NOR3_X1    g2165(.A1(new_n1639_), .A2(new_n1640_), .A3(new_n2550_), .ZN(new_n2551_));
  NAND4_X1   g2166(.A1(new_n2196_), .A2(new_n2544_), .A3(new_n2547_), .A4(new_n2551_), .ZN(new_n2552_));
  AOI21_X1   g2167(.A1(new_n2552_), .A2(new_n2538_), .B(new_n978_), .ZN(\grant[100] ));
  NOR2_X1    g2168(.A1(new_n989_), .A2(new_n982_), .ZN(new_n2554_));
  NOR4_X1    g2169(.A1(new_n973_), .A2(new_n1007_), .A3(new_n1766_), .A4(new_n2554_), .ZN(new_n2555_));
  INV_X1     g2170(.I(\req[102] ), .ZN(new_n2556_));
  AOI21_X1   g2171(.A1(new_n2556_), .A2(\priority[102] ), .B(\priority[103] ), .ZN(new_n2557_));
  OAI21_X1   g2172(.A1(new_n533_), .A2(new_n528_), .B(new_n2557_), .ZN(new_n2558_));
  NOR3_X1    g2173(.A1(new_n1618_), .A2(new_n1771_), .A3(new_n2558_), .ZN(new_n2559_));
  NAND4_X1   g2174(.A1(new_n1928_), .A2(new_n2212_), .A3(new_n2555_), .A4(new_n2559_), .ZN(new_n2560_));
  AOI21_X1   g2175(.A1(new_n2560_), .A2(new_n2548_), .B(new_n491_), .ZN(\grant[101] ));
  NOR2_X1    g2176(.A1(new_n1160_), .A2(new_n495_), .ZN(new_n2562_));
  NOR4_X1    g2177(.A1(new_n1156_), .A2(new_n1166_), .A3(new_n1776_), .A4(new_n2562_), .ZN(new_n2563_));
  INV_X1     g2178(.I(\req[103] ), .ZN(new_n2564_));
  AOI21_X1   g2179(.A1(new_n2564_), .A2(\priority[103] ), .B(\priority[104] ), .ZN(new_n2565_));
  OAI21_X1   g2180(.A1(new_n779_), .A2(new_n774_), .B(new_n2565_), .ZN(new_n2566_));
  NOR3_X1    g2181(.A1(new_n1645_), .A2(new_n1781_), .A3(new_n2566_), .ZN(new_n2567_));
  NAND4_X1   g2182(.A1(new_n1939_), .A2(new_n2221_), .A3(new_n2563_), .A4(new_n2567_), .ZN(new_n2568_));
  AOI21_X1   g2183(.A1(new_n2568_), .A2(new_n2556_), .B(new_n737_), .ZN(\grant[102] ));
  OAI22_X1   g2184(.A1(new_n906_), .A2(new_n911_), .B1(new_n981_), .B2(new_n976_), .ZN(new_n2570_));
  NOR4_X1    g2185(.A1(new_n2312_), .A2(new_n2398_), .A3(new_n2484_), .A4(new_n2570_), .ZN(new_n2571_));
  NOR2_X1    g2186(.A1(new_n1242_), .A2(new_n741_), .ZN(new_n2572_));
  NOR4_X1    g2187(.A1(new_n1238_), .A2(new_n1248_), .A3(new_n1786_), .A4(new_n2572_), .ZN(new_n2573_));
  INV_X1     g2188(.I(\req[104] ), .ZN(new_n2574_));
  AOI21_X1   g2189(.A1(new_n2574_), .A2(\priority[104] ), .B(\priority[105] ), .ZN(new_n2575_));
  OAI21_X1   g2190(.A1(new_n1025_), .A2(new_n1020_), .B(new_n2575_), .ZN(new_n2576_));
  NOR3_X1    g2191(.A1(new_n1791_), .A2(new_n1880_), .A3(new_n2576_), .ZN(new_n2577_));
  NAND4_X1   g2192(.A1(new_n2231_), .A2(new_n2571_), .A3(new_n2573_), .A4(new_n2577_), .ZN(new_n2578_));
  AOI21_X1   g2193(.A1(new_n2578_), .A2(new_n2564_), .B(new_n983_), .ZN(\grant[103] ));
  OAI22_X1   g2194(.A1(new_n1131_), .A2(new_n1133_), .B1(new_n1159_), .B2(new_n1157_), .ZN(new_n2580_));
  NOR4_X1    g2195(.A1(new_n2322_), .A2(new_n2408_), .A3(new_n2494_), .A4(new_n2580_), .ZN(new_n2581_));
  NOR2_X1    g2196(.A1(new_n1321_), .A2(new_n987_), .ZN(new_n2582_));
  NOR4_X1    g2197(.A1(new_n1317_), .A2(new_n1327_), .A3(new_n1796_), .A4(new_n2582_), .ZN(new_n2583_));
  INV_X1     g2198(.I(\req[105] ), .ZN(new_n2584_));
  AOI21_X1   g2199(.A1(new_n2584_), .A2(\priority[105] ), .B(\priority[106] ), .ZN(new_n2585_));
  OAI21_X1   g2200(.A1(new_n1174_), .A2(new_n1172_), .B(new_n2585_), .ZN(new_n2586_));
  NOR3_X1    g2201(.A1(new_n1801_), .A2(new_n1889_), .A3(new_n2586_), .ZN(new_n2587_));
  NAND4_X1   g2202(.A1(new_n2241_), .A2(new_n2581_), .A3(new_n2583_), .A4(new_n2587_), .ZN(new_n2588_));
  AOI21_X1   g2203(.A1(new_n2588_), .A2(new_n2574_), .B(new_n496_), .ZN(\grant[104] ));
  OAI22_X1   g2204(.A1(new_n1213_), .A2(new_n1215_), .B1(new_n1241_), .B2(new_n1239_), .ZN(new_n2590_));
  NOR4_X1    g2205(.A1(new_n2332_), .A2(new_n2418_), .A3(new_n2504_), .A4(new_n2590_), .ZN(new_n2591_));
  NOR2_X1    g2206(.A1(new_n1399_), .A2(new_n502_), .ZN(new_n2592_));
  NOR4_X1    g2207(.A1(new_n1395_), .A2(new_n1405_), .A3(new_n1806_), .A4(new_n2592_), .ZN(new_n2593_));
  INV_X1     g2208(.I(\req[106] ), .ZN(new_n2594_));
  AOI21_X1   g2209(.A1(new_n2594_), .A2(\priority[106] ), .B(\priority[107] ), .ZN(new_n2595_));
  OAI21_X1   g2210(.A1(new_n1256_), .A2(new_n1254_), .B(new_n2595_), .ZN(new_n2596_));
  NOR3_X1    g2211(.A1(new_n1811_), .A2(new_n1898_), .A3(new_n2596_), .ZN(new_n2597_));
  NAND4_X1   g2212(.A1(new_n2251_), .A2(new_n2591_), .A3(new_n2593_), .A4(new_n2597_), .ZN(new_n2598_));
  AOI21_X1   g2213(.A1(new_n2598_), .A2(new_n2584_), .B(new_n742_), .ZN(\grant[105] ));
  OAI22_X1   g2214(.A1(new_n1295_), .A2(new_n1297_), .B1(new_n1320_), .B2(new_n1318_), .ZN(new_n2600_));
  NOR4_X1    g2215(.A1(new_n2342_), .A2(new_n2428_), .A3(new_n2514_), .A4(new_n2600_), .ZN(new_n2601_));
  NOR2_X1    g2216(.A1(new_n1477_), .A2(new_n748_), .ZN(new_n2602_));
  NOR4_X1    g2217(.A1(new_n1473_), .A2(new_n1483_), .A3(new_n1816_), .A4(new_n2602_), .ZN(new_n2603_));
  INV_X1     g2218(.I(\req[107] ), .ZN(new_n2604_));
  AOI21_X1   g2219(.A1(new_n2604_), .A2(\priority[107] ), .B(\priority[108] ), .ZN(new_n2605_));
  OAI21_X1   g2220(.A1(new_n1335_), .A2(new_n1333_), .B(new_n2605_), .ZN(new_n2606_));
  NOR3_X1    g2221(.A1(new_n1821_), .A2(new_n1907_), .A3(new_n2606_), .ZN(new_n2607_));
  NAND4_X1   g2222(.A1(new_n2261_), .A2(new_n2601_), .A3(new_n2603_), .A4(new_n2607_), .ZN(new_n2608_));
  AOI21_X1   g2223(.A1(new_n2608_), .A2(new_n2594_), .B(new_n988_), .ZN(\grant[106] ));
  OAI22_X1   g2224(.A1(new_n1373_), .A2(new_n1375_), .B1(new_n1398_), .B2(new_n1396_), .ZN(new_n2610_));
  NOR4_X1    g2225(.A1(new_n2352_), .A2(new_n2438_), .A3(new_n2524_), .A4(new_n2610_), .ZN(new_n2611_));
  NOR2_X1    g2226(.A1(new_n1555_), .A2(new_n994_), .ZN(new_n2612_));
  NOR4_X1    g2227(.A1(new_n1551_), .A2(new_n1561_), .A3(new_n1826_), .A4(new_n2612_), .ZN(new_n2613_));
  INV_X1     g2228(.I(\req[108] ), .ZN(new_n2614_));
  AOI21_X1   g2229(.A1(new_n2614_), .A2(\priority[108] ), .B(\priority[109] ), .ZN(new_n2615_));
  OAI21_X1   g2230(.A1(new_n1413_), .A2(new_n1411_), .B(new_n2615_), .ZN(new_n2616_));
  NOR3_X1    g2231(.A1(new_n1831_), .A2(new_n1916_), .A3(new_n2616_), .ZN(new_n2617_));
  NAND4_X1   g2232(.A1(new_n2271_), .A2(new_n2611_), .A3(new_n2613_), .A4(new_n2617_), .ZN(new_n2618_));
  AOI21_X1   g2233(.A1(new_n2618_), .A2(new_n2604_), .B(new_n503_), .ZN(\grant[107] ));
  NOR4_X1    g2234(.A1(new_n1449_), .A2(new_n1459_), .A3(new_n1464_), .A4(new_n1509_), .ZN(new_n2620_));
  NOR2_X1    g2235(.A1(new_n514_), .A2(new_n507_), .ZN(new_n2621_));
  OAI22_X1   g2236(.A1(new_n1474_), .A2(new_n1476_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n2622_));
  NOR4_X1    g2237(.A1(new_n1454_), .A2(new_n1837_), .A3(new_n2622_), .A4(new_n2621_), .ZN(new_n2623_));
  INV_X1     g2238(.I(\req[109] ), .ZN(new_n2624_));
  AOI21_X1   g2239(.A1(new_n2624_), .A2(\priority[109] ), .B(\priority[110] ), .ZN(new_n2625_));
  OAI21_X1   g2240(.A1(new_n472_), .A2(new_n467_), .B(new_n2625_), .ZN(new_n2626_));
  NOR3_X1    g2241(.A1(new_n1493_), .A2(new_n1613_), .A3(new_n2626_), .ZN(new_n2627_));
  NAND4_X1   g2242(.A1(new_n2274_), .A2(new_n2620_), .A3(new_n2623_), .A4(new_n2627_), .ZN(new_n2628_));
  AOI21_X1   g2243(.A1(new_n2628_), .A2(new_n2614_), .B(new_n749_), .ZN(\grant[108] ));
  NOR4_X1    g2244(.A1(new_n1527_), .A2(new_n1537_), .A3(new_n1542_), .A4(new_n1587_), .ZN(new_n2630_));
  NOR2_X1    g2245(.A1(new_n760_), .A2(new_n753_), .ZN(new_n2631_));
  OAI22_X1   g2246(.A1(new_n1552_), .A2(new_n1554_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n2632_));
  NOR4_X1    g2247(.A1(new_n1532_), .A2(new_n1849_), .A3(new_n2632_), .A4(new_n2631_), .ZN(new_n2633_));
  INV_X1     g2248(.I(\req[110] ), .ZN(new_n2634_));
  AOI21_X1   g2249(.A1(new_n2634_), .A2(\priority[110] ), .B(\priority[111] ), .ZN(new_n2635_));
  OAI21_X1   g2250(.A1(new_n718_), .A2(new_n713_), .B(new_n2635_), .ZN(new_n2636_));
  NOR3_X1    g2251(.A1(new_n1571_), .A2(new_n1640_), .A3(new_n2636_), .ZN(new_n2637_));
  NAND4_X1   g2252(.A1(new_n2284_), .A2(new_n2630_), .A3(new_n2633_), .A4(new_n2637_), .ZN(new_n2638_));
  AOI21_X1   g2253(.A1(new_n2638_), .A2(new_n2624_), .B(new_n995_), .ZN(\grant[109] ));
  NOR2_X1    g2254(.A1(new_n1006_), .A2(new_n999_), .ZN(new_n2640_));
  NOR4_X1    g2255(.A1(new_n973_), .A2(new_n1602_), .A3(new_n1766_), .A4(new_n2640_), .ZN(new_n2641_));
  INV_X1     g2256(.I(\req[111] ), .ZN(new_n2642_));
  AOI21_X1   g2257(.A1(new_n2642_), .A2(\priority[111] ), .B(\priority[112] ), .ZN(new_n2643_));
  OAI21_X1   g2258(.A1(new_n533_), .A2(new_n528_), .B(new_n2643_), .ZN(new_n2644_));
  NOR3_X1    g2259(.A1(new_n1618_), .A2(new_n1771_), .A3(new_n2644_), .ZN(new_n2645_));
  NAND4_X1   g2260(.A1(new_n1928_), .A2(new_n2212_), .A3(new_n2641_), .A4(new_n2645_), .ZN(new_n2646_));
  AOI21_X1   g2261(.A1(new_n2646_), .A2(new_n2634_), .B(new_n508_), .ZN(\grant[110] ));
  NOR2_X1    g2262(.A1(new_n1165_), .A2(new_n512_), .ZN(new_n2648_));
  NOR4_X1    g2263(.A1(new_n1156_), .A2(new_n1629_), .A3(new_n1776_), .A4(new_n2648_), .ZN(new_n2649_));
  INV_X1     g2264(.I(\req[112] ), .ZN(new_n2650_));
  AOI21_X1   g2265(.A1(new_n2650_), .A2(\priority[112] ), .B(\priority[113] ), .ZN(new_n2651_));
  OAI21_X1   g2266(.A1(new_n779_), .A2(new_n774_), .B(new_n2651_), .ZN(new_n2652_));
  NOR3_X1    g2267(.A1(new_n1645_), .A2(new_n1781_), .A3(new_n2652_), .ZN(new_n2653_));
  NAND4_X1   g2268(.A1(new_n1939_), .A2(new_n2221_), .A3(new_n2649_), .A4(new_n2653_), .ZN(new_n2654_));
  AOI21_X1   g2269(.A1(new_n2654_), .A2(new_n2642_), .B(new_n754_), .ZN(\grant[111] ));
  NOR2_X1    g2270(.A1(new_n1247_), .A2(new_n758_), .ZN(new_n2656_));
  OAI22_X1   g2271(.A1(new_n984_), .A2(new_n989_), .B1(new_n998_), .B2(new_n993_), .ZN(new_n2657_));
  NOR4_X1    g2272(.A1(new_n1238_), .A2(new_n1786_), .A3(new_n2657_), .A4(new_n2656_), .ZN(new_n2658_));
  INV_X1     g2273(.I(\req[113] ), .ZN(new_n2659_));
  AOI21_X1   g2274(.A1(new_n2659_), .A2(\priority[113] ), .B(\priority[114] ), .ZN(new_n2660_));
  OAI21_X1   g2275(.A1(new_n1025_), .A2(new_n1020_), .B(new_n2660_), .ZN(new_n2661_));
  NOR3_X1    g2276(.A1(new_n1791_), .A2(new_n1880_), .A3(new_n2661_), .ZN(new_n2662_));
  NAND4_X1   g2277(.A1(new_n2231_), .A2(new_n2571_), .A3(new_n2658_), .A4(new_n2662_), .ZN(new_n2663_));
  AOI21_X1   g2278(.A1(new_n2663_), .A2(new_n2650_), .B(new_n1000_), .ZN(\grant[112] ));
  NOR2_X1    g2279(.A1(new_n1326_), .A2(new_n1004_), .ZN(new_n2665_));
  OAI22_X1   g2280(.A1(new_n1158_), .A2(new_n1160_), .B1(new_n1164_), .B2(new_n1162_), .ZN(new_n2666_));
  NOR4_X1    g2281(.A1(new_n1317_), .A2(new_n1796_), .A3(new_n2666_), .A4(new_n2665_), .ZN(new_n2667_));
  INV_X1     g2282(.I(\req[114] ), .ZN(new_n2668_));
  AOI21_X1   g2283(.A1(new_n2668_), .A2(\priority[114] ), .B(\priority[115] ), .ZN(new_n2669_));
  OAI21_X1   g2284(.A1(new_n1174_), .A2(new_n1172_), .B(new_n2669_), .ZN(new_n2670_));
  NOR3_X1    g2285(.A1(new_n1801_), .A2(new_n1889_), .A3(new_n2670_), .ZN(new_n2671_));
  NAND4_X1   g2286(.A1(new_n2241_), .A2(new_n2581_), .A3(new_n2667_), .A4(new_n2671_), .ZN(new_n2672_));
  AOI21_X1   g2287(.A1(new_n2672_), .A2(new_n2659_), .B(new_n513_), .ZN(\grant[113] ));
  NOR2_X1    g2288(.A1(new_n1404_), .A2(new_n468_), .ZN(new_n2674_));
  OAI22_X1   g2289(.A1(new_n1240_), .A2(new_n1242_), .B1(new_n1246_), .B2(new_n1244_), .ZN(new_n2675_));
  NOR4_X1    g2290(.A1(new_n1395_), .A2(new_n1806_), .A3(new_n2675_), .A4(new_n2674_), .ZN(new_n2676_));
  INV_X1     g2291(.I(\req[115] ), .ZN(new_n2677_));
  AOI21_X1   g2292(.A1(new_n2677_), .A2(\priority[115] ), .B(\priority[116] ), .ZN(new_n2678_));
  OAI21_X1   g2293(.A1(new_n1256_), .A2(new_n1254_), .B(new_n2678_), .ZN(new_n2679_));
  NOR3_X1    g2294(.A1(new_n1811_), .A2(new_n1898_), .A3(new_n2679_), .ZN(new_n2680_));
  NAND4_X1   g2295(.A1(new_n2251_), .A2(new_n2591_), .A3(new_n2676_), .A4(new_n2680_), .ZN(new_n2681_));
  AOI21_X1   g2296(.A1(new_n2681_), .A2(new_n2668_), .B(new_n759_), .ZN(\grant[114] ));
  NOR2_X1    g2297(.A1(new_n1482_), .A2(new_n714_), .ZN(new_n2683_));
  OAI22_X1   g2298(.A1(new_n1319_), .A2(new_n1321_), .B1(new_n1325_), .B2(new_n1323_), .ZN(new_n2684_));
  NOR4_X1    g2299(.A1(new_n1473_), .A2(new_n1816_), .A3(new_n2684_), .A4(new_n2683_), .ZN(new_n2685_));
  INV_X1     g2300(.I(\req[116] ), .ZN(new_n2686_));
  AOI21_X1   g2301(.A1(new_n2686_), .A2(\priority[116] ), .B(\priority[117] ), .ZN(new_n2687_));
  OAI21_X1   g2302(.A1(new_n1335_), .A2(new_n1333_), .B(new_n2687_), .ZN(new_n2688_));
  NOR3_X1    g2303(.A1(new_n1821_), .A2(new_n1907_), .A3(new_n2688_), .ZN(new_n2689_));
  NAND4_X1   g2304(.A1(new_n2261_), .A2(new_n2601_), .A3(new_n2685_), .A4(new_n2689_), .ZN(new_n2690_));
  AOI21_X1   g2305(.A1(new_n2690_), .A2(new_n2677_), .B(new_n1005_), .ZN(\grant[115] ));
  NOR2_X1    g2306(.A1(new_n1560_), .A2(new_n960_), .ZN(new_n2692_));
  OAI22_X1   g2307(.A1(new_n1397_), .A2(new_n1399_), .B1(new_n1403_), .B2(new_n1402_), .ZN(new_n2693_));
  NOR4_X1    g2308(.A1(new_n1551_), .A2(new_n1826_), .A3(new_n2693_), .A4(new_n2692_), .ZN(new_n2694_));
  INV_X1     g2309(.I(\req[117] ), .ZN(new_n2695_));
  AOI21_X1   g2310(.A1(new_n2695_), .A2(\priority[117] ), .B(\priority[118] ), .ZN(new_n2696_));
  OAI21_X1   g2311(.A1(new_n1413_), .A2(new_n1411_), .B(new_n2696_), .ZN(new_n2697_));
  NOR3_X1    g2312(.A1(new_n1831_), .A2(new_n1916_), .A3(new_n2697_), .ZN(new_n2698_));
  NAND4_X1   g2313(.A1(new_n2271_), .A2(new_n2611_), .A3(new_n2694_), .A4(new_n2698_), .ZN(new_n2699_));
  AOI21_X1   g2314(.A1(new_n2699_), .A2(new_n2686_), .B(new_n469_), .ZN(\grant[116] ));
  NOR2_X1    g2315(.A1(new_n480_), .A2(new_n473_), .ZN(new_n2701_));
  OAI22_X1   g2316(.A1(new_n1480_), .A2(new_n1481_), .B1(new_n1610_), .B2(new_n1609_), .ZN(new_n2702_));
  NOR4_X1    g2317(.A1(new_n1478_), .A2(new_n1837_), .A3(new_n2702_), .A4(new_n2701_), .ZN(new_n2703_));
  INV_X1     g2318(.I(\req[118] ), .ZN(new_n2704_));
  AOI21_X1   g2319(.A1(new_n2704_), .A2(\priority[118] ), .B(\priority[119] ), .ZN(new_n2705_));
  OAI21_X1   g2320(.A1(new_n463_), .A2(new_n458_), .B(new_n2705_), .ZN(new_n2706_));
  NOR3_X1    g2321(.A1(new_n1493_), .A2(new_n1498_), .A3(new_n2706_), .ZN(new_n2707_));
  NAND4_X1   g2322(.A1(new_n1465_), .A2(new_n1520_), .A3(new_n2703_), .A4(new_n2707_), .ZN(new_n2708_));
  AOI21_X1   g2323(.A1(new_n2708_), .A2(new_n2695_), .B(new_n715_), .ZN(\grant[117] ));
  NOR2_X1    g2324(.A1(new_n726_), .A2(new_n719_), .ZN(new_n2710_));
  OAI22_X1   g2325(.A1(new_n1558_), .A2(new_n1559_), .B1(new_n1637_), .B2(new_n1636_), .ZN(new_n2711_));
  NOR4_X1    g2326(.A1(new_n1556_), .A2(new_n1849_), .A3(new_n2711_), .A4(new_n2710_), .ZN(new_n2712_));
  INV_X1     g2327(.I(\req[119] ), .ZN(new_n2713_));
  AOI21_X1   g2328(.A1(new_n2713_), .A2(\priority[119] ), .B(\priority[120] ), .ZN(new_n2714_));
  OAI21_X1   g2329(.A1(new_n709_), .A2(new_n704_), .B(new_n2714_), .ZN(new_n2715_));
  NOR3_X1    g2330(.A1(new_n1571_), .A2(new_n1576_), .A3(new_n2715_), .ZN(new_n2716_));
  NAND4_X1   g2331(.A1(new_n1543_), .A2(new_n1598_), .A3(new_n2712_), .A4(new_n2716_), .ZN(new_n2717_));
  AOI21_X1   g2332(.A1(new_n2717_), .A2(new_n2704_), .B(new_n961_), .ZN(\grant[118] ));
  NOR2_X1    g2333(.A1(new_n972_), .A2(new_n965_), .ZN(new_n2719_));
  NOR4_X1    g2334(.A1(new_n1602_), .A2(new_n1612_), .A3(new_n1766_), .A4(new_n2719_), .ZN(new_n2720_));
  INV_X1     g2335(.I(\req[120] ), .ZN(new_n2721_));
  AOI21_X1   g2336(.A1(new_n2721_), .A2(\priority[120] ), .B(\priority[121] ), .ZN(new_n2722_));
  OAI21_X1   g2337(.A1(new_n533_), .A2(new_n528_), .B(new_n2722_), .ZN(new_n2723_));
  NOR3_X1    g2338(.A1(new_n1618_), .A2(new_n1771_), .A3(new_n2723_), .ZN(new_n2724_));
  NAND4_X1   g2339(.A1(new_n1928_), .A2(new_n2212_), .A3(new_n2720_), .A4(new_n2724_), .ZN(new_n2725_));
  AOI21_X1   g2340(.A1(new_n2725_), .A2(new_n2713_), .B(new_n474_), .ZN(\grant[119] ));
  NOR2_X1    g2341(.A1(new_n1155_), .A2(new_n478_), .ZN(new_n2727_));
  NOR4_X1    g2342(.A1(new_n1629_), .A2(new_n1639_), .A3(new_n1776_), .A4(new_n2727_), .ZN(new_n2728_));
  INV_X1     g2343(.I(\req[121] ), .ZN(new_n2729_));
  AOI21_X1   g2344(.A1(new_n2729_), .A2(\priority[121] ), .B(\priority[122] ), .ZN(new_n2730_));
  OAI21_X1   g2345(.A1(new_n779_), .A2(new_n774_), .B(new_n2730_), .ZN(new_n2731_));
  NOR3_X1    g2346(.A1(new_n1645_), .A2(new_n1781_), .A3(new_n2731_), .ZN(new_n2732_));
  NAND4_X1   g2347(.A1(new_n1939_), .A2(new_n2221_), .A3(new_n2728_), .A4(new_n2732_), .ZN(new_n2733_));
  AOI21_X1   g2348(.A1(new_n2733_), .A2(new_n2721_), .B(new_n720_), .ZN(\grant[120] ));
  NOR2_X1    g2349(.A1(new_n1237_), .A2(new_n724_), .ZN(new_n2735_));
  OAI22_X1   g2350(.A1(new_n959_), .A2(new_n964_), .B1(new_n1006_), .B2(new_n1001_), .ZN(new_n2736_));
  NOR4_X1    g2351(.A1(new_n1786_), .A2(new_n2657_), .A3(new_n2736_), .A4(new_n2735_), .ZN(new_n2737_));
  INV_X1     g2352(.I(\req[122] ), .ZN(new_n2738_));
  AOI21_X1   g2353(.A1(new_n2738_), .A2(\priority[122] ), .B(\priority[123] ), .ZN(new_n2739_));
  OAI21_X1   g2354(.A1(new_n1025_), .A2(new_n1020_), .B(new_n2739_), .ZN(new_n2740_));
  NOR3_X1    g2355(.A1(new_n1791_), .A2(new_n1880_), .A3(new_n2740_), .ZN(new_n2741_));
  NAND4_X1   g2356(.A1(new_n2231_), .A2(new_n2571_), .A3(new_n2737_), .A4(new_n2741_), .ZN(new_n2742_));
  AOI21_X1   g2357(.A1(new_n2742_), .A2(new_n2729_), .B(new_n966_), .ZN(\grant[121] ));
  NOR2_X1    g2358(.A1(new_n1316_), .A2(new_n970_), .ZN(new_n2744_));
  OAI22_X1   g2359(.A1(new_n1152_), .A2(new_n1154_), .B1(new_n1165_), .B2(new_n1163_), .ZN(new_n2745_));
  NOR4_X1    g2360(.A1(new_n1796_), .A2(new_n2666_), .A3(new_n2745_), .A4(new_n2744_), .ZN(new_n2746_));
  INV_X1     g2361(.I(\req[123] ), .ZN(new_n2747_));
  AOI21_X1   g2362(.A1(new_n2747_), .A2(\priority[123] ), .B(\priority[124] ), .ZN(new_n2748_));
  OAI21_X1   g2363(.A1(new_n1174_), .A2(new_n1172_), .B(new_n2748_), .ZN(new_n2749_));
  NOR3_X1    g2364(.A1(new_n1801_), .A2(new_n1889_), .A3(new_n2749_), .ZN(new_n2750_));
  NAND4_X1   g2365(.A1(new_n2241_), .A2(new_n2581_), .A3(new_n2746_), .A4(new_n2750_), .ZN(new_n2751_));
  AOI21_X1   g2366(.A1(new_n2751_), .A2(new_n2738_), .B(new_n479_), .ZN(\grant[122] ));
  NOR2_X1    g2367(.A1(new_n1394_), .A2(new_n459_), .ZN(new_n2753_));
  OAI22_X1   g2368(.A1(new_n1234_), .A2(new_n1236_), .B1(new_n1247_), .B2(new_n1245_), .ZN(new_n2754_));
  NOR4_X1    g2369(.A1(new_n1806_), .A2(new_n2675_), .A3(new_n2754_), .A4(new_n2753_), .ZN(new_n2755_));
  INV_X1     g2370(.I(\req[124] ), .ZN(new_n2756_));
  AOI21_X1   g2371(.A1(new_n2756_), .A2(\priority[124] ), .B(\priority[125] ), .ZN(new_n2757_));
  OAI21_X1   g2372(.A1(new_n1256_), .A2(new_n1254_), .B(new_n2757_), .ZN(new_n2758_));
  NOR3_X1    g2373(.A1(new_n1811_), .A2(new_n1898_), .A3(new_n2758_), .ZN(new_n2759_));
  NAND4_X1   g2374(.A1(new_n2251_), .A2(new_n2591_), .A3(new_n2755_), .A4(new_n2759_), .ZN(new_n2760_));
  AOI21_X1   g2375(.A1(new_n2760_), .A2(new_n2747_), .B(new_n725_), .ZN(\grant[123] ));
  NOR2_X1    g2376(.A1(new_n1472_), .A2(new_n705_), .ZN(new_n2762_));
  OAI22_X1   g2377(.A1(new_n1313_), .A2(new_n1315_), .B1(new_n1326_), .B2(new_n1324_), .ZN(new_n2763_));
  NOR4_X1    g2378(.A1(new_n1816_), .A2(new_n2684_), .A3(new_n2763_), .A4(new_n2762_), .ZN(new_n2764_));
  INV_X1     g2379(.I(\req[125] ), .ZN(new_n2765_));
  AOI21_X1   g2380(.A1(new_n2765_), .A2(\priority[125] ), .B(\priority[126] ), .ZN(new_n2766_));
  OAI21_X1   g2381(.A1(new_n1335_), .A2(new_n1333_), .B(new_n2766_), .ZN(new_n2767_));
  NOR3_X1    g2382(.A1(new_n1821_), .A2(new_n1907_), .A3(new_n2767_), .ZN(new_n2768_));
  NAND4_X1   g2383(.A1(new_n2261_), .A2(new_n2601_), .A3(new_n2764_), .A4(new_n2768_), .ZN(new_n2769_));
  AOI21_X1   g2384(.A1(new_n2769_), .A2(new_n2756_), .B(new_n971_), .ZN(\grant[124] ));
  NOR2_X1    g2385(.A1(new_n1550_), .A2(new_n951_), .ZN(new_n2771_));
  OAI22_X1   g2386(.A1(new_n1401_), .A2(new_n1404_), .B1(new_n1393_), .B2(new_n1392_), .ZN(new_n2772_));
  NOR4_X1    g2387(.A1(new_n1826_), .A2(new_n2693_), .A3(new_n2772_), .A4(new_n2771_), .ZN(new_n2773_));
  INV_X1     g2388(.I(\req[126] ), .ZN(new_n2774_));
  AOI21_X1   g2389(.A1(new_n2774_), .A2(\priority[126] ), .B(\priority[127] ), .ZN(new_n2775_));
  OAI21_X1   g2390(.A1(new_n1413_), .A2(new_n1411_), .B(new_n2775_), .ZN(new_n2776_));
  NOR3_X1    g2391(.A1(new_n1831_), .A2(new_n1916_), .A3(new_n2776_), .ZN(new_n2777_));
  NAND4_X1   g2392(.A1(new_n2271_), .A2(new_n2611_), .A3(new_n2773_), .A4(new_n2777_), .ZN(new_n2778_));
  AOI21_X1   g2393(.A1(new_n2778_), .A2(new_n2765_), .B(new_n460_), .ZN(\grant[125] ));
  OAI22_X1   g2394(.A1(new_n1446_), .A2(new_n1448_), .B1(new_n1452_), .B2(new_n1450_), .ZN(new_n2780_));
  OAI22_X1   g2395(.A1(new_n1451_), .A2(new_n1453_), .B1(new_n1476_), .B2(new_n1474_), .ZN(new_n2781_));
  OAI22_X1   g2396(.A1(new_n1456_), .A2(new_n1458_), .B1(new_n1462_), .B2(new_n1461_), .ZN(new_n2782_));
  OAI22_X1   g2397(.A1(new_n1460_), .A2(new_n1463_), .B1(new_n1447_), .B2(new_n1445_), .ZN(new_n2783_));
  NOR4_X1    g2398(.A1(new_n2780_), .A2(new_n2781_), .A3(new_n2782_), .A4(new_n2783_), .ZN(new_n2784_));
  NOR2_X1    g2399(.A1(new_n1610_), .A2(new_n1147_), .ZN(new_n2785_));
  OAI22_X1   g2400(.A1(new_n1475_), .A2(new_n1477_), .B1(new_n1481_), .B2(new_n1480_), .ZN(new_n2786_));
  OAI22_X1   g2401(.A1(new_n1479_), .A2(new_n1482_), .B1(new_n1471_), .B2(new_n1470_), .ZN(new_n2787_));
  NOR4_X1    g2402(.A1(new_n1837_), .A2(new_n2786_), .A3(new_n2787_), .A4(new_n2785_), .ZN(new_n2788_));
  INV_X1     g2403(.I(\req[127] ), .ZN(new_n2789_));
  AOI21_X1   g2404(.A1(new_n2789_), .A2(\priority[127] ), .B(\priority[0] ), .ZN(new_n2790_));
  OAI21_X1   g2405(.A1(new_n1491_), .A2(new_n1489_), .B(new_n2790_), .ZN(new_n2791_));
  OAI22_X1   g2406(.A1(new_n1490_), .A2(new_n1492_), .B1(new_n1496_), .B2(new_n1494_), .ZN(new_n2792_));
  OAI22_X1   g2407(.A1(new_n1495_), .A2(new_n1497_), .B1(new_n1512_), .B2(new_n1510_), .ZN(new_n2793_));
  NOR3_X1    g2408(.A1(new_n2792_), .A2(new_n2793_), .A3(new_n2791_), .ZN(new_n2794_));
  OAI22_X1   g2409(.A1(new_n1501_), .A2(new_n1503_), .B1(new_n1507_), .B2(new_n1506_), .ZN(new_n2795_));
  OAI22_X1   g2410(.A1(new_n1505_), .A2(new_n1508_), .B1(new_n1457_), .B2(new_n1455_), .ZN(new_n2796_));
  OAI22_X1   g2411(.A1(new_n1511_), .A2(new_n1513_), .B1(new_n1517_), .B2(new_n1516_), .ZN(new_n2797_));
  OAI22_X1   g2412(.A1(new_n1515_), .A2(new_n1518_), .B1(new_n1502_), .B2(new_n1500_), .ZN(new_n2798_));
  NOR4_X1    g2413(.A1(new_n2795_), .A2(new_n2796_), .A3(new_n2797_), .A4(new_n2798_), .ZN(new_n2799_));
  NAND4_X1   g2414(.A1(new_n2784_), .A2(new_n2799_), .A3(new_n2788_), .A4(new_n2794_), .ZN(new_n2800_));
  AOI21_X1   g2415(.A1(new_n2800_), .A2(new_n2774_), .B(new_n706_), .ZN(\grant[126] ));
  OAI22_X1   g2416(.A1(new_n1524_), .A2(new_n1526_), .B1(new_n1530_), .B2(new_n1528_), .ZN(new_n2802_));
  OAI22_X1   g2417(.A1(new_n1529_), .A2(new_n1531_), .B1(new_n1554_), .B2(new_n1552_), .ZN(new_n2803_));
  OAI22_X1   g2418(.A1(new_n1534_), .A2(new_n1536_), .B1(new_n1540_), .B2(new_n1539_), .ZN(new_n2804_));
  OAI22_X1   g2419(.A1(new_n1538_), .A2(new_n1541_), .B1(new_n1525_), .B2(new_n1523_), .ZN(new_n2805_));
  NOR4_X1    g2420(.A1(new_n2802_), .A2(new_n2803_), .A3(new_n2804_), .A4(new_n2805_), .ZN(new_n2806_));
  NOR2_X1    g2421(.A1(new_n1637_), .A2(new_n1229_), .ZN(new_n2807_));
  OAI22_X1   g2422(.A1(new_n1553_), .A2(new_n1555_), .B1(new_n1559_), .B2(new_n1558_), .ZN(new_n2808_));
  OAI22_X1   g2423(.A1(new_n1557_), .A2(new_n1560_), .B1(new_n1549_), .B2(new_n1548_), .ZN(new_n2809_));
  NOR4_X1    g2424(.A1(new_n1849_), .A2(new_n2808_), .A3(new_n2809_), .A4(new_n2807_), .ZN(new_n2810_));
  AOI21_X1   g2425(.A1(new_n386_), .A2(\priority[0] ), .B(\priority[1] ), .ZN(new_n2811_));
  OAI21_X1   g2426(.A1(new_n1569_), .A2(new_n1567_), .B(new_n2811_), .ZN(new_n2812_));
  OAI22_X1   g2427(.A1(new_n1568_), .A2(new_n1570_), .B1(new_n1574_), .B2(new_n1572_), .ZN(new_n2813_));
  OAI22_X1   g2428(.A1(new_n1573_), .A2(new_n1575_), .B1(new_n1590_), .B2(new_n1588_), .ZN(new_n2814_));
  NOR3_X1    g2429(.A1(new_n2813_), .A2(new_n2814_), .A3(new_n2812_), .ZN(new_n2815_));
  OAI22_X1   g2430(.A1(new_n1579_), .A2(new_n1581_), .B1(new_n1585_), .B2(new_n1584_), .ZN(new_n2816_));
  OAI22_X1   g2431(.A1(new_n1583_), .A2(new_n1586_), .B1(new_n1535_), .B2(new_n1533_), .ZN(new_n2817_));
  OAI22_X1   g2432(.A1(new_n1589_), .A2(new_n1591_), .B1(new_n1595_), .B2(new_n1594_), .ZN(new_n2818_));
  OAI22_X1   g2433(.A1(new_n1593_), .A2(new_n1596_), .B1(new_n1580_), .B2(new_n1578_), .ZN(new_n2819_));
  NOR4_X1    g2434(.A1(new_n2816_), .A2(new_n2817_), .A3(new_n2818_), .A4(new_n2819_), .ZN(new_n2820_));
  NAND4_X1   g2435(.A1(new_n2806_), .A2(new_n2820_), .A3(new_n2810_), .A4(new_n2815_), .ZN(new_n2821_));
  AOI21_X1   g2436(.A1(new_n2821_), .A2(new_n2789_), .B(new_n952_), .ZN(\grant[127] ));
  NAND4_X1   g2437(.A1(new_n478_), .A2(new_n766_), .A3(new_n780_), .A4(new_n792_), .ZN(new_n2823_));
  NAND4_X1   g2438(.A1(new_n468_), .A2(new_n485_), .A3(new_n495_), .A4(new_n507_), .ZN(new_n2824_));
  NAND4_X1   g2439(.A1(new_n675_), .A2(new_n815_), .A3(new_n827_), .A4(new_n837_), .ZN(new_n2825_));
  NAND4_X1   g2440(.A1(new_n802_), .A2(new_n849_), .A3(new_n861_), .A4(new_n871_), .ZN(new_n2826_));
  NOR4_X1    g2441(.A1(new_n2823_), .A2(new_n2824_), .A3(new_n2825_), .A4(new_n2826_), .ZN(new_n2827_));
  NAND4_X1   g2442(.A1(new_n564_), .A2(new_n598_), .A3(new_n608_), .A4(new_n620_), .ZN(new_n2828_));
  NAND4_X1   g2443(.A1(new_n517_), .A2(new_n529_), .A3(new_n539_), .A4(new_n551_), .ZN(new_n2829_));
  NAND4_X1   g2444(.A1(new_n390_), .A2(new_n400_), .A3(new_n412_), .A4(new_n446_), .ZN(new_n2830_));
  NAND4_X1   g2445(.A1(new_n424_), .A2(new_n434_), .A3(new_n574_), .A4(new_n586_), .ZN(new_n2831_));
  NOR4_X1    g2446(.A1(new_n2828_), .A2(new_n2829_), .A3(new_n2830_), .A4(new_n2831_), .ZN(new_n2832_));
  NAND4_X1   g2447(.A1(new_n882_), .A2(new_n916_), .A3(new_n926_), .A4(new_n938_), .ZN(new_n2833_));
  NAND4_X1   g2448(.A1(new_n1056_), .A2(new_n1066_), .A3(new_n1078_), .A4(new_n1112_), .ZN(new_n2834_));
  NAND4_X1   g2449(.A1(new_n960_), .A2(new_n970_), .A3(new_n999_), .A4(new_n1147_), .ZN(new_n2835_));
  NAND4_X1   g2450(.A1(new_n892_), .A2(new_n904_), .A3(new_n977_), .A4(new_n987_), .ZN(new_n2836_));
  NOR4_X1    g2451(.A1(new_n2833_), .A2(new_n2834_), .A3(new_n2835_), .A4(new_n2836_), .ZN(new_n2837_));
  NAND4_X1   g2452(.A1(new_n663_), .A2(new_n736_), .A3(new_n748_), .A4(new_n758_), .ZN(new_n2838_));
  NAND4_X1   g2453(.A1(new_n641_), .A2(new_n653_), .A3(new_n687_), .A4(new_n697_), .ZN(new_n2839_));
  NAND4_X1   g2454(.A1(new_n1031_), .A2(new_n1043_), .A3(new_n1090_), .A4(new_n1100_), .ZN(new_n2840_));
  NAND4_X1   g2455(.A1(new_n705_), .A2(new_n719_), .A3(new_n1009_), .A4(new_n1021_), .ZN(new_n2841_));
  NOR4_X1    g2456(.A1(new_n2838_), .A2(new_n2839_), .A3(new_n2840_), .A4(new_n2841_), .ZN(new_n2842_));
  AND4_X2    g2457(.A1(new_n2827_), .A2(new_n2832_), .A3(new_n2837_), .A4(new_n2842_), .Z(anyGrant));
endmodule


