// Benchmark "sin" written by ABC on Thu Sep 14 20:28:55 2023

module sin ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ;
  output \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24] ;
  wire new_n50_, new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_,
    new_n57_, new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_,
    new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_,
    new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_,
    new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_,
    new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_,
    new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_,
    new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_,
    new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_,
    new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_,
    new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_,
    new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_,
    new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_,
    new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_,
    new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_,
    new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_,
    new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_,
    new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_,
    new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_,
    new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_,
    new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_,
    new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_,
    new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_,
    new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_,
    new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_,
    new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_,
    new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_,
    new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_,
    new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_,
    new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_,
    new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_,
    new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_,
    new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_,
    new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_,
    new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_,
    new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_,
    new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_,
    new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_,
    new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_,
    new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_,
    new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_,
    new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_,
    new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_,
    new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_,
    new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_,
    new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_,
    new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_,
    new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_,
    new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_,
    new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_,
    new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_,
    new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_,
    new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_,
    new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_,
    new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_,
    new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_,
    new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_,
    new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_,
    new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_,
    new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_,
    new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_,
    new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_,
    new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_,
    new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_,
    new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_,
    new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_,
    new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_,
    new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_,
    new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_,
    new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_,
    new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_,
    new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_,
    new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4445_, new_n4446_, new_n4447_, new_n4448_,
    new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_,
    new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_,
    new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_,
    new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_,
    new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_,
    new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_,
    new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_,
    new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_,
    new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_,
    new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_,
    new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_,
    new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_,
    new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_,
    new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4575_,
    new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_,
    new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_,
    new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_,
    new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_,
    new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4648_,
    new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_,
    new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_,
    new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_,
    new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_,
    new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_,
    new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_,
    new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_,
    new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_,
    new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_,
    new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_,
    new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_,
    new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_,
    new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_,
    new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_,
    new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4848_,
    new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_,
    new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_,
    new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_,
    new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_,
    new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_,
    new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4885_,
    new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_,
    new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_,
    new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_,
    new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_,
    new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_,
    new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_,
    new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_,
    new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_,
    new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_,
    new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_,
    new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_,
    new_n5018_, new_n5019_, new_n5021_, new_n5022_, new_n5023_, new_n5024_,
    new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_,
    new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_,
    new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_,
    new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_,
    new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_,
    new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_,
    new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_,
    new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_,
    new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_,
    new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_,
    new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_,
    new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_,
    new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_,
    new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_,
    new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_,
    new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_,
    new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_,
    new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_,
    new_n5133_, new_n5134_, new_n5135_, new_n5137_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_,
    new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5152_,
    new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_,
    new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_,
    new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_,
    new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_,
    new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_,
    new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_,
    new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_,
    new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_,
    new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_,
    new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_,
    new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_,
    new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_,
    new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_,
    new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_,
    new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_,
    new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_,
    new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_,
    new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_,
    new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_,
    new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_,
    new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_,
    new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_,
    new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_,
    new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_,
    new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_,
    new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_,
    new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_,
    new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_,
    new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_,
    new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_,
    new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_,
    new_n5424_, new_n5425_, new_n5426_, new_n5428_, new_n5429_, new_n5430_,
    new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_,
    new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_,
    new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_,
    new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_,
    new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_,
    new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_,
    new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_,
    new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_,
    new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_,
    new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_,
    new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_,
    new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_,
    new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_,
    new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_,
    new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_,
    new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_,
    new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_,
    new_n5533_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_,
    new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_,
    new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_,
    new_n5624_, new_n5625_, new_n5627_, new_n5628_, new_n5629_, new_n5630_,
    new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_,
    new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_,
    new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_,
    new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_,
    new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_,
    new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_,
    new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_,
    new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_,
    new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_,
    new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_,
    new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_,
    new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_,
    new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_,
    new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_,
    new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_,
    new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_, new_n5726_,
    new_n5727_, new_n5728_, new_n5729_, new_n5731_, new_n5732_, new_n5733_,
    new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_,
    new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_,
    new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_,
    new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_,
    new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_,
    new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_, new_n5769_,
    new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_,
    new_n5776_, new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_,
    new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_,
    new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_,
    new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_,
    new_n5800_, new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_,
    new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_,
    new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_,
    new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_,
    new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_,
    new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_,
    new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_,
    new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_,
    new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_,
    new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_,
    new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_,
    new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_,
    new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_,
    new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_,
    new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5940_,
    new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_,
    new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_,
    new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_,
    new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_,
    new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_,
    new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_,
    new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_,
    new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_,
    new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_,
    new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_,
    new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_,
    new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_,
    new_n6013_, new_n6014_, new_n6016_, new_n6017_, new_n6018_, new_n6019_,
    new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_,
    new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_,
    new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_,
    new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_,
    new_n6044_, new_n6045_, new_n6046_, new_n6048_, new_n6049_, new_n6050_,
    new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_,
    new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_,
    new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_,
    new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_,
    new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_,
    new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_,
    new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_,
    new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6099_,
    new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_,
    new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_,
    new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_,
    new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_,
    new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_,
    new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_,
    new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_,
    new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_,
    new_n6161_, new_n6162_, new_n6164_, new_n6165_, new_n6166_, new_n6167_,
    new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_,
    new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6180_,
    new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_,
    new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_,
    new_n6193_, new_n6194_, new_n6195_, new_n6200_, new_n6201_, new_n6202_,
    new_n6203_, new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_,
    new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_,
    new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6221_, new_n6222_,
    new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_,
    new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_,
    new_n6235_, new_n6236_, new_n6238_, new_n6239_, new_n6240_, new_n6241_,
    new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_,
    new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_;
  AND4_X2    g0000(.A1(\a[0] ), .A2(\a[1] ), .A3(\a[2] ), .A4(\a[3] ), .Z(new_n50_));
  AND3_X2    g0001(.A1(\a[4] ), .A2(\a[5] ), .A3(\a[6] ), .Z(new_n51_));
  NAND2_X1   g0002(.A1(new_n50_), .A2(new_n51_), .ZN(new_n52_));
  NAND3_X1   g0003(.A1(\a[7] ), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n53_));
  NAND3_X1   g0004(.A1(\a[10] ), .A2(\a[11] ), .A3(\a[12] ), .ZN(new_n54_));
  NOR2_X1    g0005(.A1(\a[13] ), .A2(\a[14] ), .ZN(new_n55_));
  INV_X1     g0006(.I(new_n55_), .ZN(new_n56_));
  NOR4_X1    g0007(.A1(new_n52_), .A2(new_n53_), .A3(new_n54_), .A4(new_n56_), .ZN(new_n57_));
  NAND4_X1   g0008(.A1(\a[0] ), .A2(\a[1] ), .A3(\a[2] ), .A4(\a[3] ), .ZN(new_n58_));
  NAND3_X1   g0009(.A1(\a[4] ), .A2(\a[5] ), .A3(\a[6] ), .ZN(new_n59_));
  NOR4_X1    g0010(.A1(new_n58_), .A2(new_n59_), .A3(new_n53_), .A4(new_n54_), .ZN(new_n60_));
  AOI21_X1   g0011(.A1(new_n60_), .A2(new_n55_), .B(\a[22] ), .ZN(new_n61_));
  INV_X1     g0012(.I(\a[22] ), .ZN(new_n62_));
  NAND2_X1   g0013(.A1(new_n62_), .A2(\a[15] ), .ZN(new_n63_));
  OAI22_X1   g0014(.A1(new_n57_), .A2(new_n63_), .B1(new_n61_), .B2(\a[15] ), .ZN(new_n64_));
  INV_X1     g0015(.I(\a[15] ), .ZN(new_n65_));
  INV_X1     g0016(.I(\a[16] ), .ZN(new_n66_));
  INV_X1     g0017(.I(\a[17] ), .ZN(new_n67_));
  NOR3_X1    g0018(.A1(new_n65_), .A2(new_n66_), .A3(new_n67_), .ZN(new_n68_));
  NOR2_X1    g0019(.A1(\a[18] ), .A2(\a[19] ), .ZN(new_n69_));
  NAND4_X1   g0020(.A1(new_n60_), .A2(new_n55_), .A3(new_n68_), .A4(new_n69_), .ZN(new_n70_));
  AOI21_X1   g0021(.A1(new_n70_), .A2(new_n62_), .B(\a[20] ), .ZN(new_n71_));
  AND3_X2    g0022(.A1(\a[7] ), .A2(\a[8] ), .A3(\a[9] ), .Z(new_n72_));
  NAND3_X1   g0023(.A1(new_n50_), .A2(new_n51_), .A3(new_n72_), .ZN(new_n73_));
  INV_X1     g0024(.I(new_n68_), .ZN(new_n74_));
  NOR4_X1    g0025(.A1(new_n73_), .A2(new_n54_), .A3(new_n56_), .A4(new_n74_), .ZN(new_n75_));
  NAND2_X1   g0026(.A1(new_n62_), .A2(\a[20] ), .ZN(new_n76_));
  AOI21_X1   g0027(.A1(new_n75_), .A2(new_n69_), .B(new_n76_), .ZN(new_n77_));
  OAI21_X1   g0028(.A1(new_n71_), .A2(new_n77_), .B(new_n64_), .ZN(new_n78_));
  INV_X1     g0029(.I(\a[21] ), .ZN(new_n79_));
  INV_X1     g0030(.I(\a[18] ), .ZN(new_n80_));
  INV_X1     g0031(.I(\a[19] ), .ZN(new_n81_));
  INV_X1     g0032(.I(\a[20] ), .ZN(new_n82_));
  NOR3_X1    g0033(.A1(new_n80_), .A2(new_n81_), .A3(new_n82_), .ZN(new_n83_));
  NAND4_X1   g0034(.A1(new_n60_), .A2(new_n55_), .A3(new_n68_), .A4(new_n83_), .ZN(new_n84_));
  NOR3_X1    g0035(.A1(new_n58_), .A2(new_n59_), .A3(new_n53_), .ZN(new_n85_));
  INV_X1     g0036(.I(new_n54_), .ZN(new_n86_));
  NAND4_X1   g0037(.A1(new_n85_), .A2(new_n86_), .A3(new_n55_), .A4(new_n68_), .ZN(new_n87_));
  INV_X1     g0038(.I(new_n83_), .ZN(new_n88_));
  OAI21_X1   g0039(.A1(new_n87_), .A2(new_n88_), .B(new_n62_), .ZN(new_n89_));
  NOR2_X1    g0040(.A1(new_n79_), .A2(\a[22] ), .ZN(new_n90_));
  AOI22_X1   g0041(.A1(new_n89_), .A2(new_n79_), .B1(new_n84_), .B2(new_n90_), .ZN(new_n91_));
  NAND2_X1   g0042(.A1(\a[0] ), .A2(\a[1] ), .ZN(new_n92_));
  NAND2_X1   g0043(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n93_));
  NOR3_X1    g0044(.A1(new_n59_), .A2(new_n92_), .A3(new_n93_), .ZN(new_n94_));
  NAND4_X1   g0045(.A1(new_n94_), .A2(new_n72_), .A3(new_n86_), .A4(new_n55_), .ZN(new_n95_));
  NOR2_X1    g0046(.A1(new_n81_), .A2(new_n62_), .ZN(new_n96_));
  OAI21_X1   g0047(.A1(new_n95_), .A2(new_n74_), .B(new_n96_), .ZN(new_n97_));
  INV_X1     g0048(.I(new_n96_), .ZN(new_n98_));
  NAND4_X1   g0049(.A1(new_n60_), .A2(new_n55_), .A3(new_n68_), .A4(new_n98_), .ZN(new_n99_));
  XNOR2_X1   g0050(.A1(\a[18] ), .A2(\a[22] ), .ZN(new_n100_));
  INV_X1     g0051(.I(new_n100_), .ZN(new_n101_));
  NAND3_X1   g0052(.A1(new_n97_), .A2(new_n99_), .A3(new_n101_), .ZN(new_n102_));
  NOR2_X1    g0053(.A1(new_n66_), .A2(new_n62_), .ZN(new_n103_));
  INV_X1     g0054(.I(new_n103_), .ZN(new_n104_));
  NAND4_X1   g0055(.A1(new_n60_), .A2(new_n65_), .A3(new_n55_), .A4(new_n104_), .ZN(new_n105_));
  OAI21_X1   g0056(.A1(new_n95_), .A2(\a[15] ), .B(new_n103_), .ZN(new_n106_));
  XNOR2_X1   g0057(.A1(\a[16] ), .A2(\a[17] ), .ZN(new_n107_));
  INV_X1     g0058(.I(new_n107_), .ZN(new_n108_));
  NAND3_X1   g0059(.A1(new_n106_), .A2(new_n105_), .A3(new_n108_), .ZN(new_n109_));
  NOR4_X1    g0060(.A1(new_n78_), .A2(new_n91_), .A3(new_n102_), .A4(new_n109_), .ZN(new_n110_));
  NAND2_X1   g0061(.A1(\a[21] ), .A2(\a[22] ), .ZN(new_n111_));
  INV_X1     g0062(.I(new_n111_), .ZN(new_n112_));
  NOR2_X1    g0063(.A1(new_n70_), .A2(new_n112_), .ZN(new_n113_));
  AOI21_X1   g0064(.A1(new_n75_), .A2(new_n69_), .B(new_n111_), .ZN(new_n114_));
  INV_X1     g0065(.I(new_n76_), .ZN(new_n115_));
  NOR2_X1    g0066(.A1(new_n62_), .A2(\a[20] ), .ZN(new_n116_));
  NOR2_X1    g0067(.A1(new_n115_), .A2(new_n116_), .ZN(new_n117_));
  NOR3_X1    g0068(.A1(new_n114_), .A2(new_n113_), .A3(new_n117_), .ZN(new_n118_));
  NAND2_X1   g0069(.A1(new_n95_), .A2(new_n62_), .ZN(new_n119_));
  AOI21_X1   g0070(.A1(new_n60_), .A2(new_n55_), .B(new_n63_), .ZN(new_n120_));
  AOI21_X1   g0071(.A1(new_n119_), .A2(new_n65_), .B(new_n120_), .ZN(new_n121_));
  NOR2_X1    g0072(.A1(new_n67_), .A2(new_n62_), .ZN(new_n122_));
  INV_X1     g0073(.I(new_n122_), .ZN(new_n123_));
  AOI21_X1   g0074(.A1(new_n57_), .A2(new_n65_), .B(new_n123_), .ZN(new_n124_));
  NAND4_X1   g0075(.A1(new_n60_), .A2(new_n65_), .A3(new_n55_), .A4(new_n123_), .ZN(new_n125_));
  INV_X1     g0076(.I(new_n125_), .ZN(new_n126_));
  XNOR2_X1   g0077(.A1(\a[16] ), .A2(\a[22] ), .ZN(new_n127_));
  NOR3_X1    g0078(.A1(new_n124_), .A2(new_n126_), .A3(new_n127_), .ZN(new_n128_));
  OAI21_X1   g0079(.A1(new_n95_), .A2(new_n74_), .B(\a[18] ), .ZN(new_n129_));
  NAND4_X1   g0080(.A1(new_n60_), .A2(new_n80_), .A3(new_n55_), .A4(new_n68_), .ZN(new_n130_));
  AOI22_X1   g0081(.A1(new_n97_), .A2(new_n99_), .B1(new_n129_), .B2(new_n130_), .ZN(new_n131_));
  NAND4_X1   g0082(.A1(new_n118_), .A2(new_n128_), .A3(new_n131_), .A4(new_n121_), .ZN(new_n132_));
  NAND4_X1   g0083(.A1(new_n85_), .A2(new_n65_), .A3(new_n86_), .A4(new_n55_), .ZN(new_n133_));
  NAND2_X1   g0084(.A1(new_n133_), .A2(new_n122_), .ZN(new_n134_));
  OAI21_X1   g0085(.A1(new_n95_), .A2(\a[15] ), .B(\a[16] ), .ZN(new_n135_));
  NAND4_X1   g0086(.A1(new_n60_), .A2(new_n65_), .A3(new_n66_), .A4(new_n55_), .ZN(new_n136_));
  AOI22_X1   g0087(.A1(new_n134_), .A2(new_n125_), .B1(new_n135_), .B2(new_n136_), .ZN(new_n137_));
  AOI21_X1   g0088(.A1(new_n70_), .A2(new_n112_), .B(new_n117_), .ZN(new_n138_));
  INV_X1     g0089(.I(new_n138_), .ZN(new_n139_));
  NOR3_X1    g0090(.A1(new_n139_), .A2(new_n113_), .A3(new_n64_), .ZN(new_n140_));
  NAND3_X1   g0091(.A1(new_n140_), .A2(new_n131_), .A3(new_n137_), .ZN(new_n141_));
  INV_X1     g0092(.I(new_n69_), .ZN(new_n142_));
  NOR3_X1    g0093(.A1(new_n95_), .A2(new_n74_), .A3(new_n142_), .ZN(new_n143_));
  OAI21_X1   g0094(.A1(new_n143_), .A2(\a[22] ), .B(new_n82_), .ZN(new_n144_));
  NAND2_X1   g0095(.A1(new_n70_), .A2(new_n115_), .ZN(new_n145_));
  AOI21_X1   g0096(.A1(new_n144_), .A2(new_n145_), .B(new_n121_), .ZN(new_n146_));
  AOI21_X1   g0097(.A1(new_n75_), .A2(new_n83_), .B(\a[22] ), .ZN(new_n147_));
  NAND2_X1   g0098(.A1(new_n84_), .A2(new_n90_), .ZN(new_n148_));
  OAI21_X1   g0099(.A1(new_n147_), .A2(\a[21] ), .B(new_n148_), .ZN(new_n149_));
  NOR2_X1    g0100(.A1(new_n102_), .A2(new_n109_), .ZN(new_n150_));
  NAND3_X1   g0101(.A1(new_n146_), .A2(new_n150_), .A3(new_n149_), .ZN(new_n151_));
  NAND3_X1   g0102(.A1(new_n141_), .A2(new_n151_), .A3(new_n132_), .ZN(new_n152_));
  NAND2_X1   g0103(.A1(new_n134_), .A2(new_n125_), .ZN(new_n153_));
  NAND2_X1   g0104(.A1(new_n135_), .A2(new_n136_), .ZN(new_n154_));
  NAND2_X1   g0105(.A1(new_n153_), .A2(new_n154_), .ZN(new_n155_));
  NOR4_X1    g0106(.A1(new_n78_), .A2(new_n155_), .A3(new_n91_), .A4(new_n102_), .ZN(new_n156_));
  NOR2_X1    g0107(.A1(new_n75_), .A2(new_n98_), .ZN(new_n157_));
  INV_X1     g0108(.I(new_n99_), .ZN(new_n158_));
  NOR3_X1    g0109(.A1(new_n157_), .A2(new_n158_), .A3(new_n100_), .ZN(new_n159_));
  NAND4_X1   g0110(.A1(new_n146_), .A2(new_n137_), .A3(new_n149_), .A4(new_n159_), .ZN(new_n160_));
  INV_X1     g0111(.I(new_n127_), .ZN(new_n161_));
  NAND3_X1   g0112(.A1(new_n134_), .A2(new_n125_), .A3(new_n161_), .ZN(new_n162_));
  NAND2_X1   g0113(.A1(new_n97_), .A2(new_n99_), .ZN(new_n163_));
  INV_X1     g0114(.I(new_n163_), .ZN(new_n164_));
  XOR2_X1    g0115(.A1(new_n87_), .A2(\a[18] ), .Z(new_n165_));
  NOR3_X1    g0116(.A1(new_n164_), .A2(new_n165_), .A3(new_n162_), .ZN(new_n166_));
  NOR3_X1    g0117(.A1(new_n139_), .A2(new_n113_), .A3(new_n121_), .ZN(new_n167_));
  NAND2_X1   g0118(.A1(new_n166_), .A2(new_n167_), .ZN(new_n168_));
  NAND2_X1   g0119(.A1(new_n128_), .A2(new_n131_), .ZN(new_n169_));
  NAND2_X1   g0120(.A1(new_n129_), .A2(new_n130_), .ZN(new_n170_));
  NAND4_X1   g0121(.A1(new_n153_), .A2(new_n163_), .A3(new_n170_), .A4(new_n154_), .ZN(new_n171_));
  NAND3_X1   g0122(.A1(new_n75_), .A2(new_n69_), .A3(new_n111_), .ZN(new_n172_));
  NAND3_X1   g0123(.A1(new_n64_), .A2(new_n172_), .A3(new_n138_), .ZN(new_n173_));
  NOR3_X1    g0124(.A1(new_n169_), .A2(new_n171_), .A3(new_n173_), .ZN(new_n174_));
  NAND3_X1   g0125(.A1(new_n174_), .A2(new_n168_), .A3(new_n160_), .ZN(new_n175_));
  NOR4_X1    g0126(.A1(new_n175_), .A2(new_n110_), .A3(new_n152_), .A4(new_n156_), .ZN(new_n176_));
  NOR2_X1    g0127(.A1(new_n124_), .A2(new_n126_), .ZN(new_n177_));
  XOR2_X1    g0128(.A1(new_n133_), .A2(\a[16] ), .Z(new_n178_));
  NOR2_X1    g0129(.A1(new_n80_), .A2(new_n62_), .ZN(new_n179_));
  INV_X1     g0130(.I(new_n179_), .ZN(new_n180_));
  NAND4_X1   g0131(.A1(new_n60_), .A2(new_n55_), .A3(new_n68_), .A4(new_n180_), .ZN(new_n181_));
  NAND2_X1   g0132(.A1(new_n87_), .A2(new_n179_), .ZN(new_n182_));
  XNOR2_X1   g0133(.A1(\a[18] ), .A2(\a[19] ), .ZN(new_n183_));
  INV_X1     g0134(.I(new_n183_), .ZN(new_n184_));
  NAND3_X1   g0135(.A1(new_n182_), .A2(new_n181_), .A3(new_n184_), .ZN(new_n185_));
  NOR3_X1    g0136(.A1(new_n177_), .A2(new_n178_), .A3(new_n185_), .ZN(new_n186_));
  NAND2_X1   g0137(.A1(new_n186_), .A2(new_n167_), .ZN(new_n187_));
  NOR2_X1    g0138(.A1(new_n77_), .A2(new_n71_), .ZN(new_n188_));
  NOR2_X1    g0139(.A1(new_n188_), .A2(new_n91_), .ZN(new_n189_));
  NOR3_X1    g0140(.A1(new_n164_), .A2(new_n165_), .A3(new_n109_), .ZN(new_n190_));
  NAND3_X1   g0141(.A1(new_n190_), .A2(new_n189_), .A3(new_n64_), .ZN(new_n191_));
  NOR2_X1    g0142(.A1(new_n191_), .A2(new_n187_), .ZN(new_n192_));
  NAND2_X1   g0143(.A1(new_n172_), .A2(new_n138_), .ZN(new_n193_));
  AOI21_X1   g0144(.A1(new_n87_), .A2(new_n179_), .B(new_n183_), .ZN(new_n194_));
  NAND4_X1   g0145(.A1(new_n153_), .A2(new_n154_), .A3(new_n181_), .A4(new_n194_), .ZN(new_n195_));
  NOR3_X1    g0146(.A1(new_n195_), .A2(new_n193_), .A3(new_n64_), .ZN(new_n196_));
  NOR3_X1    g0147(.A1(new_n173_), .A2(new_n162_), .A3(new_n185_), .ZN(new_n197_));
  NAND3_X1   g0148(.A1(new_n192_), .A2(new_n196_), .A3(new_n197_), .ZN(new_n198_));
  NAND3_X1   g0149(.A1(new_n121_), .A2(new_n172_), .A3(new_n138_), .ZN(new_n199_));
  NOR2_X1    g0150(.A1(new_n195_), .A2(new_n199_), .ZN(new_n200_));
  NAND4_X1   g0151(.A1(new_n146_), .A2(new_n131_), .A3(new_n149_), .A4(new_n137_), .ZN(new_n201_));
  NOR2_X1    g0152(.A1(new_n162_), .A2(new_n185_), .ZN(new_n202_));
  NAND2_X1   g0153(.A1(new_n140_), .A2(new_n202_), .ZN(new_n203_));
  NAND3_X1   g0154(.A1(new_n201_), .A2(new_n203_), .A3(new_n200_), .ZN(new_n204_));
  NOR4_X1    g0155(.A1(new_n171_), .A2(new_n121_), .A3(new_n188_), .A4(new_n91_), .ZN(new_n205_));
  NOR3_X1    g0156(.A1(new_n188_), .A2(new_n91_), .A3(new_n121_), .ZN(new_n206_));
  NAND2_X1   g0157(.A1(new_n206_), .A2(new_n190_), .ZN(new_n207_));
  NOR4_X1    g0158(.A1(new_n198_), .A2(new_n204_), .A3(new_n205_), .A4(new_n207_), .ZN(new_n208_));
  NAND2_X1   g0159(.A1(new_n140_), .A2(new_n150_), .ZN(new_n209_));
  AOI21_X1   g0160(.A1(new_n133_), .A2(new_n103_), .B(new_n107_), .ZN(new_n210_));
  NAND4_X1   g0161(.A1(new_n163_), .A2(new_n170_), .A3(new_n105_), .A4(new_n210_), .ZN(new_n211_));
  NOR2_X1    g0162(.A1(new_n211_), .A2(new_n199_), .ZN(new_n212_));
  INV_X1     g0163(.I(new_n212_), .ZN(new_n213_));
  NAND2_X1   g0164(.A1(new_n167_), .A2(new_n150_), .ZN(new_n214_));
  NOR2_X1    g0165(.A1(new_n162_), .A2(new_n102_), .ZN(new_n215_));
  AOI21_X1   g0166(.A1(new_n144_), .A2(new_n145_), .B(new_n64_), .ZN(new_n216_));
  NAND3_X1   g0167(.A1(new_n216_), .A2(new_n215_), .A3(new_n91_), .ZN(new_n217_));
  INV_X1     g0168(.I(new_n217_), .ZN(new_n218_));
  NOR3_X1    g0169(.A1(new_n155_), .A2(new_n173_), .A3(new_n102_), .ZN(new_n219_));
  NOR2_X1    g0170(.A1(new_n211_), .A2(new_n173_), .ZN(new_n220_));
  NAND4_X1   g0171(.A1(new_n118_), .A2(new_n131_), .A3(new_n137_), .A4(new_n64_), .ZN(new_n221_));
  NAND4_X1   g0172(.A1(new_n118_), .A2(new_n131_), .A3(new_n137_), .A4(new_n121_), .ZN(new_n222_));
  NOR2_X1    g0173(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND4_X1   g0174(.A1(new_n223_), .A2(new_n218_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n224_));
  NOR4_X1    g0175(.A1(new_n224_), .A2(new_n209_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n225_));
  NAND3_X1   g0176(.A1(new_n208_), .A2(new_n176_), .A3(new_n225_), .ZN(new_n226_));
  NAND3_X1   g0177(.A1(new_n166_), .A2(new_n91_), .A3(new_n216_), .ZN(new_n227_));
  NOR2_X1    g0178(.A1(new_n171_), .A2(new_n173_), .ZN(new_n228_));
  NAND2_X1   g0179(.A1(new_n163_), .A2(new_n170_), .ZN(new_n229_));
  NOR4_X1    g0180(.A1(new_n78_), .A2(new_n162_), .A3(new_n229_), .A4(new_n91_), .ZN(new_n230_));
  NOR2_X1    g0181(.A1(new_n230_), .A2(new_n228_), .ZN(new_n231_));
  NOR4_X1    g0182(.A1(new_n78_), .A2(new_n162_), .A3(new_n91_), .A4(new_n185_), .ZN(new_n232_));
  NOR3_X1    g0183(.A1(new_n195_), .A2(new_n78_), .A3(new_n91_), .ZN(new_n233_));
  NOR2_X1    g0184(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1   g0185(.A1(new_n234_), .A2(new_n231_), .A3(new_n227_), .ZN(new_n235_));
  AOI21_X1   g0186(.A1(new_n75_), .A2(new_n69_), .B(\a[22] ), .ZN(new_n236_));
  OAI21_X1   g0187(.A1(new_n236_), .A2(\a[20] ), .B(new_n145_), .ZN(new_n237_));
  NOR3_X1    g0188(.A1(new_n229_), .A2(new_n155_), .A3(new_n91_), .ZN(new_n238_));
  NAND4_X1   g0189(.A1(new_n210_), .A2(new_n194_), .A3(new_n105_), .A4(new_n181_), .ZN(new_n239_));
  NOR2_X1    g0190(.A1(new_n173_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1     g0191(.I(new_n240_), .ZN(new_n241_));
  NAND4_X1   g0192(.A1(new_n241_), .A2(new_n238_), .A3(new_n222_), .A4(new_n237_), .ZN(new_n242_));
  NAND3_X1   g0193(.A1(new_n146_), .A2(new_n202_), .A3(new_n149_), .ZN(new_n243_));
  NOR2_X1    g0194(.A1(new_n185_), .A2(new_n109_), .ZN(new_n244_));
  NAND2_X1   g0195(.A1(new_n140_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1   g0196(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1   g0197(.A1(new_n195_), .A2(new_n211_), .B(new_n173_), .ZN(new_n247_));
  NOR4_X1    g0198(.A1(new_n235_), .A2(new_n242_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n248_));
  INV_X1     g0199(.I(new_n215_), .ZN(new_n249_));
  NAND4_X1   g0200(.A1(new_n118_), .A2(new_n159_), .A3(new_n137_), .A4(new_n121_), .ZN(new_n250_));
  NAND4_X1   g0201(.A1(new_n118_), .A2(new_n159_), .A3(new_n137_), .A4(new_n64_), .ZN(new_n251_));
  NOR2_X1    g0202(.A1(new_n156_), .A2(new_n251_), .ZN(new_n252_));
  NAND4_X1   g0203(.A1(new_n146_), .A2(new_n137_), .A3(new_n91_), .A4(new_n159_), .ZN(new_n253_));
  INV_X1     g0204(.I(new_n253_), .ZN(new_n254_));
  NOR3_X1    g0205(.A1(new_n162_), .A2(new_n102_), .A3(new_n121_), .ZN(new_n255_));
  NAND2_X1   g0206(.A1(new_n189_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1   g0207(.A1(new_n166_), .A2(new_n140_), .ZN(new_n257_));
  NOR2_X1    g0208(.A1(new_n257_), .A2(new_n256_), .ZN(new_n258_));
  NAND4_X1   g0209(.A1(new_n258_), .A2(new_n252_), .A3(new_n250_), .A4(new_n254_), .ZN(new_n259_));
  NAND2_X1   g0210(.A1(new_n159_), .A2(new_n137_), .ZN(new_n260_));
  AOI21_X1   g0211(.A1(new_n260_), .A2(new_n211_), .B(new_n199_), .ZN(new_n261_));
  AND4_X2    g0212(.A1(new_n153_), .A2(new_n163_), .A3(new_n170_), .A4(new_n154_), .Z(new_n262_));
  NOR2_X1    g0213(.A1(new_n262_), .A2(new_n118_), .ZN(new_n263_));
  NOR4_X1    g0214(.A1(new_n259_), .A2(new_n249_), .A3(new_n261_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1   g0215(.A1(new_n264_), .A2(new_n248_), .ZN(new_n265_));
  NOR2_X1    g0216(.A1(new_n226_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1     g0217(.I(\a[7] ), .ZN(new_n267_));
  NOR2_X1    g0218(.A1(\a[8] ), .A2(\a[22] ), .ZN(new_n268_));
  AOI21_X1   g0219(.A1(new_n52_), .A2(new_n268_), .B(new_n267_), .ZN(new_n269_));
  XOR2_X1    g0220(.A1(new_n269_), .A2(\a[9] ), .Z(new_n270_));
  INV_X1     g0221(.I(new_n270_), .ZN(new_n271_));
  NOR2_X1    g0222(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  NOR4_X1    g0223(.A1(new_n193_), .A2(new_n64_), .A3(new_n162_), .A4(new_n102_), .ZN(new_n273_));
  AOI21_X1   g0224(.A1(new_n84_), .A2(new_n62_), .B(\a[21] ), .ZN(new_n274_));
  INV_X1     g0225(.I(new_n148_), .ZN(new_n275_));
  OAI22_X1   g0226(.A1(new_n275_), .A2(new_n274_), .B1(new_n77_), .B2(new_n71_), .ZN(new_n276_));
  NOR3_X1    g0227(.A1(new_n171_), .A2(new_n276_), .A3(new_n121_), .ZN(new_n277_));
  INV_X1     g0228(.I(new_n181_), .ZN(new_n278_));
  NOR2_X1    g0229(.A1(new_n75_), .A2(new_n180_), .ZN(new_n279_));
  NOR3_X1    g0230(.A1(new_n279_), .A2(new_n278_), .A3(new_n183_), .ZN(new_n280_));
  NAND4_X1   g0231(.A1(new_n146_), .A2(new_n137_), .A3(new_n149_), .A4(new_n280_), .ZN(new_n281_));
  NAND3_X1   g0232(.A1(new_n146_), .A2(new_n244_), .A3(new_n149_), .ZN(new_n282_));
  AOI21_X1   g0233(.A1(new_n171_), .A2(new_n195_), .B(new_n199_), .ZN(new_n283_));
  NOR4_X1    g0234(.A1(new_n257_), .A2(new_n283_), .A3(new_n281_), .A4(new_n282_), .ZN(new_n284_));
  NAND3_X1   g0235(.A1(new_n216_), .A2(new_n202_), .A3(new_n149_), .ZN(new_n285_));
  NAND2_X1   g0236(.A1(\a[20] ), .A2(\a[22] ), .ZN(new_n286_));
  NAND3_X1   g0237(.A1(new_n75_), .A2(new_n69_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1     g0238(.I(new_n286_), .ZN(new_n288_));
  XNOR2_X1   g0239(.A1(\a[20] ), .A2(\a[21] ), .ZN(new_n289_));
  AOI21_X1   g0240(.A1(new_n70_), .A2(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND3_X1   g0241(.A1(new_n64_), .A2(new_n287_), .A3(new_n290_), .ZN(new_n291_));
  NOR2_X1    g0242(.A1(new_n171_), .A2(new_n291_), .ZN(new_n292_));
  NOR3_X1    g0243(.A1(new_n156_), .A2(new_n292_), .A3(new_n285_), .ZN(new_n293_));
  NAND2_X1   g0244(.A1(new_n284_), .A2(new_n293_), .ZN(new_n294_));
  NOR2_X1    g0245(.A1(new_n70_), .A2(new_n288_), .ZN(new_n295_));
  INV_X1     g0246(.I(new_n289_), .ZN(new_n296_));
  OAI21_X1   g0247(.A1(new_n143_), .A2(new_n286_), .B(new_n296_), .ZN(new_n297_));
  NOR3_X1    g0248(.A1(new_n297_), .A2(new_n121_), .A3(new_n295_), .ZN(new_n298_));
  NAND2_X1   g0249(.A1(new_n202_), .A2(new_n298_), .ZN(new_n299_));
  NOR4_X1    g0250(.A1(new_n168_), .A2(new_n187_), .A3(new_n221_), .A4(new_n299_), .ZN(new_n300_));
  NAND3_X1   g0251(.A1(new_n216_), .A2(new_n244_), .A3(new_n91_), .ZN(new_n301_));
  NOR3_X1    g0252(.A1(new_n261_), .A2(new_n251_), .A3(new_n301_), .ZN(new_n302_));
  NAND3_X1   g0253(.A1(new_n121_), .A2(new_n287_), .A3(new_n290_), .ZN(new_n303_));
  NOR3_X1    g0254(.A1(new_n303_), .A2(new_n162_), .A3(new_n185_), .ZN(new_n304_));
  NOR2_X1    g0255(.A1(new_n292_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1   g0256(.A1(new_n237_), .A2(new_n149_), .A3(new_n64_), .ZN(new_n306_));
  NOR2_X1    g0257(.A1(new_n306_), .A2(new_n239_), .ZN(new_n307_));
  NAND4_X1   g0258(.A1(new_n300_), .A2(new_n302_), .A3(new_n305_), .A4(new_n307_), .ZN(new_n308_));
  NOR4_X1    g0259(.A1(new_n308_), .A2(new_n273_), .A3(new_n294_), .A4(new_n277_), .ZN(new_n309_));
  NOR2_X1    g0260(.A1(new_n260_), .A2(new_n303_), .ZN(new_n310_));
  NAND3_X1   g0261(.A1(new_n216_), .A2(new_n244_), .A3(new_n149_), .ZN(new_n311_));
  NAND2_X1   g0262(.A1(new_n201_), .A2(new_n311_), .ZN(new_n312_));
  NOR3_X1    g0263(.A1(new_n276_), .A2(new_n211_), .A3(new_n121_), .ZN(new_n313_));
  NAND2_X1   g0264(.A1(new_n298_), .A2(new_n244_), .ZN(new_n314_));
  NOR3_X1    g0265(.A1(new_n177_), .A2(new_n178_), .A3(new_n102_), .ZN(new_n315_));
  NOR3_X1    g0266(.A1(new_n297_), .A2(new_n64_), .A3(new_n295_), .ZN(new_n316_));
  NAND2_X1   g0267(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1    g0268(.A1(new_n317_), .A2(new_n314_), .ZN(new_n318_));
  NOR3_X1    g0269(.A1(new_n211_), .A2(new_n78_), .A3(new_n91_), .ZN(new_n319_));
  NOR2_X1    g0270(.A1(new_n230_), .A2(new_n319_), .ZN(new_n320_));
  NAND4_X1   g0271(.A1(new_n320_), .A2(new_n318_), .A3(new_n205_), .A4(new_n313_), .ZN(new_n321_));
  NAND2_X1   g0272(.A1(new_n287_), .A2(new_n290_), .ZN(new_n322_));
  NOR3_X1    g0273(.A1(new_n171_), .A2(new_n64_), .A3(new_n322_), .ZN(new_n323_));
  NOR4_X1    g0274(.A1(new_n321_), .A2(new_n310_), .A3(new_n312_), .A4(new_n323_), .ZN(new_n324_));
  NOR4_X1    g0275(.A1(new_n193_), .A2(new_n64_), .A3(new_n102_), .A4(new_n109_), .ZN(new_n325_));
  NOR3_X1    g0276(.A1(new_n155_), .A2(new_n291_), .A3(new_n102_), .ZN(new_n326_));
  NOR3_X1    g0277(.A1(new_n156_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1     g0278(.I(new_n327_), .ZN(new_n328_));
  NOR4_X1    g0279(.A1(new_n322_), .A2(new_n64_), .A3(new_n162_), .A4(new_n102_), .ZN(new_n329_));
  NOR3_X1    g0280(.A1(new_n219_), .A2(new_n212_), .A3(new_n329_), .ZN(new_n330_));
  NOR2_X1    g0281(.A1(new_n171_), .A2(new_n199_), .ZN(new_n331_));
  NOR3_X1    g0282(.A1(new_n171_), .A2(new_n78_), .A3(new_n149_), .ZN(new_n332_));
  NOR3_X1    g0283(.A1(new_n332_), .A2(new_n331_), .A3(new_n228_), .ZN(new_n333_));
  NAND2_X1   g0284(.A1(new_n333_), .A2(new_n330_), .ZN(new_n334_));
  INV_X1     g0285(.I(new_n105_), .ZN(new_n335_));
  AOI21_X1   g0286(.A1(new_n57_), .A2(new_n65_), .B(new_n104_), .ZN(new_n336_));
  NOR3_X1    g0287(.A1(new_n336_), .A2(new_n335_), .A3(new_n107_), .ZN(new_n337_));
  NAND3_X1   g0288(.A1(new_n316_), .A2(new_n131_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1   g0289(.A1(new_n298_), .A2(new_n215_), .ZN(new_n339_));
  NOR3_X1    g0290(.A1(new_n188_), .A2(new_n91_), .A3(new_n64_), .ZN(new_n340_));
  NAND2_X1   g0291(.A1(new_n340_), .A2(new_n190_), .ZN(new_n341_));
  NOR4_X1    g0292(.A1(new_n341_), .A2(new_n160_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n342_));
  INV_X1     g0293(.I(new_n342_), .ZN(new_n343_));
  NOR2_X1    g0294(.A1(new_n160_), .A2(new_n151_), .ZN(new_n344_));
  NAND3_X1   g0295(.A1(new_n298_), .A2(new_n128_), .A3(new_n131_), .ZN(new_n345_));
  NOR2_X1    g0296(.A1(new_n345_), .A2(new_n132_), .ZN(new_n346_));
  NOR3_X1    g0297(.A1(new_n260_), .A2(new_n121_), .A3(new_n276_), .ZN(new_n347_));
  NAND4_X1   g0298(.A1(new_n344_), .A2(new_n346_), .A3(new_n332_), .A4(new_n347_), .ZN(new_n348_));
  NOR4_X1    g0299(.A1(new_n343_), .A2(new_n334_), .A3(new_n348_), .A4(new_n328_), .ZN(new_n349_));
  NAND4_X1   g0300(.A1(new_n216_), .A2(new_n128_), .A3(new_n149_), .A4(new_n131_), .ZN(new_n350_));
  AOI21_X1   g0301(.A1(new_n75_), .A2(new_n69_), .B(new_n286_), .ZN(new_n351_));
  NOR3_X1    g0302(.A1(new_n351_), .A2(new_n295_), .A3(new_n289_), .ZN(new_n352_));
  NAND3_X1   g0303(.A1(new_n150_), .A2(new_n352_), .A3(new_n64_), .ZN(new_n353_));
  NOR4_X1    g0304(.A1(new_n253_), .A2(new_n350_), .A3(new_n151_), .A4(new_n353_), .ZN(new_n354_));
  INV_X1     g0305(.I(new_n354_), .ZN(new_n355_));
  NOR3_X1    g0306(.A1(new_n276_), .A2(new_n211_), .A3(new_n121_), .ZN(new_n356_));
  NOR2_X1    g0307(.A1(new_n110_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1     g0308(.I(new_n357_), .ZN(new_n358_));
  NOR3_X1    g0309(.A1(new_n195_), .A2(new_n64_), .A3(new_n322_), .ZN(new_n359_));
  NOR4_X1    g0310(.A1(new_n193_), .A2(new_n121_), .A3(new_n162_), .A4(new_n102_), .ZN(new_n360_));
  NOR2_X1    g0311(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1   g0312(.A1(new_n361_), .A2(new_n201_), .A3(new_n214_), .ZN(new_n362_));
  NOR3_X1    g0313(.A1(new_n229_), .A2(new_n155_), .A3(new_n303_), .ZN(new_n363_));
  NOR2_X1    g0314(.A1(new_n260_), .A2(new_n199_), .ZN(new_n364_));
  NOR2_X1    g0315(.A1(new_n364_), .A2(new_n313_), .ZN(new_n365_));
  NAND4_X1   g0316(.A1(new_n146_), .A2(new_n128_), .A3(new_n149_), .A4(new_n131_), .ZN(new_n366_));
  NAND3_X1   g0317(.A1(new_n298_), .A2(new_n131_), .A3(new_n137_), .ZN(new_n367_));
  NOR2_X1    g0318(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1   g0319(.A1(new_n365_), .A2(new_n368_), .A3(new_n363_), .A4(new_n319_), .ZN(new_n369_));
  NOR4_X1    g0320(.A1(new_n369_), .A2(new_n355_), .A3(new_n358_), .A4(new_n362_), .ZN(new_n370_));
  NAND4_X1   g0321(.A1(new_n309_), .A2(new_n324_), .A3(new_n349_), .A4(new_n370_), .ZN(new_n371_));
  NAND4_X1   g0322(.A1(new_n262_), .A2(new_n64_), .A3(new_n237_), .A4(new_n149_), .ZN(new_n372_));
  NAND2_X1   g0323(.A1(new_n156_), .A2(new_n228_), .ZN(new_n373_));
  NOR4_X1    g0324(.A1(new_n229_), .A2(new_n193_), .A3(new_n64_), .A4(new_n162_), .ZN(new_n374_));
  NOR2_X1    g0325(.A1(new_n195_), .A2(new_n291_), .ZN(new_n375_));
  NOR4_X1    g0326(.A1(new_n322_), .A2(new_n121_), .A3(new_n102_), .A4(new_n109_), .ZN(new_n376_));
  NAND4_X1   g0327(.A1(new_n374_), .A2(new_n220_), .A3(new_n375_), .A4(new_n376_), .ZN(new_n377_));
  NAND2_X1   g0328(.A1(new_n262_), .A2(new_n340_), .ZN(new_n378_));
  NOR4_X1    g0329(.A1(new_n377_), .A2(new_n373_), .A3(new_n372_), .A4(new_n378_), .ZN(new_n379_));
  NOR2_X1    g0330(.A1(new_n306_), .A2(new_n169_), .ZN(new_n380_));
  NAND3_X1   g0331(.A1(new_n216_), .A2(new_n215_), .A3(new_n149_), .ZN(new_n381_));
  NAND2_X1   g0332(.A1(new_n232_), .A2(new_n203_), .ZN(new_n382_));
  NOR3_X1    g0333(.A1(new_n229_), .A2(new_n291_), .A3(new_n162_), .ZN(new_n383_));
  NOR2_X1    g0334(.A1(new_n169_), .A2(new_n303_), .ZN(new_n384_));
  NAND2_X1   g0335(.A1(new_n384_), .A2(new_n383_), .ZN(new_n385_));
  NOR4_X1    g0336(.A1(new_n385_), .A2(new_n382_), .A3(new_n380_), .A4(new_n381_), .ZN(new_n386_));
  NOR4_X1    g0337(.A1(new_n160_), .A2(new_n187_), .A3(new_n253_), .A4(new_n350_), .ZN(new_n387_));
  NOR4_X1    g0338(.A1(new_n78_), .A2(new_n229_), .A3(new_n155_), .A4(new_n91_), .ZN(new_n388_));
  NOR3_X1    g0339(.A1(new_n211_), .A2(new_n78_), .A3(new_n149_), .ZN(new_n389_));
  NAND2_X1   g0340(.A1(new_n186_), .A2(new_n140_), .ZN(new_n390_));
  NAND2_X1   g0341(.A1(new_n186_), .A2(new_n316_), .ZN(new_n391_));
  NAND3_X1   g0342(.A1(new_n390_), .A2(new_n391_), .A3(new_n222_), .ZN(new_n392_));
  NOR4_X1    g0343(.A1(new_n392_), .A2(new_n110_), .A3(new_n388_), .A4(new_n389_), .ZN(new_n393_));
  NAND4_X1   g0344(.A1(new_n393_), .A2(new_n379_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n394_));
  NAND3_X1   g0345(.A1(new_n215_), .A2(new_n352_), .A3(new_n121_), .ZN(new_n395_));
  NAND2_X1   g0346(.A1(new_n151_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1   g0347(.A1(new_n205_), .A2(new_n313_), .ZN(new_n397_));
  NAND4_X1   g0348(.A1(new_n352_), .A2(new_n131_), .A3(new_n137_), .A4(new_n121_), .ZN(new_n398_));
  NAND4_X1   g0349(.A1(new_n216_), .A2(new_n137_), .A3(new_n149_), .A4(new_n280_), .ZN(new_n399_));
  NAND2_X1   g0350(.A1(new_n399_), .A2(new_n398_), .ZN(new_n400_));
  NOR2_X1    g0351(.A1(new_n169_), .A2(new_n173_), .ZN(new_n401_));
  NAND3_X1   g0352(.A1(new_n401_), .A2(new_n232_), .A3(new_n326_), .ZN(new_n402_));
  NOR4_X1    g0353(.A1(new_n402_), .A2(new_n397_), .A3(new_n396_), .A4(new_n400_), .ZN(new_n403_));
  NAND4_X1   g0354(.A1(new_n146_), .A2(new_n131_), .A3(new_n137_), .A4(new_n91_), .ZN(new_n404_));
  NAND3_X1   g0355(.A1(new_n281_), .A2(new_n399_), .A3(new_n311_), .ZN(new_n405_));
  NAND2_X1   g0356(.A1(new_n167_), .A2(new_n202_), .ZN(new_n406_));
  NOR2_X1    g0357(.A1(new_n291_), .A2(new_n239_), .ZN(new_n407_));
  NAND3_X1   g0358(.A1(new_n406_), .A2(new_n222_), .A3(new_n407_), .ZN(new_n408_));
  NOR4_X1    g0359(.A1(new_n260_), .A2(new_n78_), .A3(new_n91_), .A4(new_n195_), .ZN(new_n409_));
  INV_X1     g0360(.I(new_n409_), .ZN(new_n410_));
  NOR4_X1    g0361(.A1(new_n405_), .A2(new_n410_), .A3(new_n408_), .A4(new_n404_), .ZN(new_n411_));
  OAI21_X1   g0362(.A1(new_n71_), .A2(new_n77_), .B(new_n121_), .ZN(new_n412_));
  NOR4_X1    g0363(.A1(new_n412_), .A2(new_n229_), .A3(new_n149_), .A4(new_n162_), .ZN(new_n413_));
  NAND4_X1   g0364(.A1(new_n313_), .A2(new_n413_), .A3(new_n319_), .A4(new_n292_), .ZN(new_n414_));
  NAND3_X1   g0365(.A1(new_n323_), .A2(new_n310_), .A3(new_n304_), .ZN(new_n415_));
  NAND4_X1   g0366(.A1(new_n118_), .A2(new_n337_), .A3(new_n131_), .A4(new_n64_), .ZN(new_n416_));
  NAND2_X1   g0367(.A1(new_n206_), .A2(new_n315_), .ZN(new_n417_));
  NAND3_X1   g0368(.A1(new_n417_), .A2(new_n388_), .A3(new_n416_), .ZN(new_n418_));
  NOR3_X1    g0369(.A1(new_n414_), .A2(new_n418_), .A3(new_n415_), .ZN(new_n419_));
  NOR2_X1    g0370(.A1(new_n211_), .A2(new_n291_), .ZN(new_n420_));
  NOR3_X1    g0371(.A1(new_n211_), .A2(new_n64_), .A3(new_n322_), .ZN(new_n421_));
  NAND3_X1   g0372(.A1(new_n421_), .A2(new_n375_), .A3(new_n420_), .ZN(new_n422_));
  NAND3_X1   g0373(.A1(new_n277_), .A2(new_n160_), .A3(new_n221_), .ZN(new_n423_));
  NAND4_X1   g0374(.A1(new_n216_), .A2(new_n137_), .A3(new_n91_), .A4(new_n280_), .ZN(new_n424_));
  NAND3_X1   g0375(.A1(new_n424_), .A2(new_n301_), .A3(new_n398_), .ZN(new_n425_));
  NOR3_X1    g0376(.A1(new_n423_), .A2(new_n425_), .A3(new_n422_), .ZN(new_n426_));
  NAND4_X1   g0377(.A1(new_n419_), .A2(new_n403_), .A3(new_n411_), .A4(new_n426_), .ZN(new_n427_));
  NOR2_X1    g0378(.A1(new_n427_), .A2(new_n394_), .ZN(new_n428_));
  XOR2_X1    g0379(.A1(new_n371_), .A2(new_n428_), .Z(new_n429_));
  INV_X1     g0380(.I(\a[13] ), .ZN(new_n430_));
  INV_X1     g0381(.I(\a[14] ), .ZN(new_n431_));
  AOI21_X1   g0382(.A1(new_n431_), .A2(new_n62_), .B(new_n430_), .ZN(new_n432_));
  INV_X1     g0383(.I(new_n432_), .ZN(new_n433_));
  NOR2_X1    g0384(.A1(new_n60_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1     g0385(.I(new_n60_), .ZN(new_n435_));
  NOR2_X1    g0386(.A1(new_n435_), .A2(new_n432_), .ZN(new_n436_));
  NOR2_X1    g0387(.A1(new_n436_), .A2(new_n434_), .ZN(new_n437_));
  INV_X1     g0388(.I(new_n437_), .ZN(new_n438_));
  NOR2_X1    g0389(.A1(new_n211_), .A2(new_n303_), .ZN(new_n439_));
  NOR2_X1    g0390(.A1(new_n209_), .A2(new_n398_), .ZN(new_n440_));
  NAND2_X1   g0391(.A1(new_n440_), .A2(new_n439_), .ZN(new_n441_));
  NAND2_X1   g0392(.A1(new_n206_), .A2(new_n166_), .ZN(new_n442_));
  NAND2_X1   g0393(.A1(new_n281_), .A2(new_n251_), .ZN(new_n443_));
  NAND2_X1   g0394(.A1(new_n364_), .A2(new_n230_), .ZN(new_n444_));
  NOR4_X1    g0395(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .A4(new_n444_), .ZN(new_n445_));
  NAND2_X1   g0396(.A1(new_n366_), .A2(new_n151_), .ZN(new_n446_));
  NOR2_X1    g0397(.A1(new_n169_), .A2(new_n199_), .ZN(new_n447_));
  NAND3_X1   g0398(.A1(new_n447_), .A2(new_n331_), .A3(new_n273_), .ZN(new_n448_));
  NAND2_X1   g0399(.A1(new_n262_), .A2(new_n206_), .ZN(new_n449_));
  NAND2_X1   g0400(.A1(new_n233_), .A2(new_n219_), .ZN(new_n450_));
  NOR4_X1    g0401(.A1(new_n448_), .A2(new_n446_), .A3(new_n450_), .A4(new_n449_), .ZN(new_n451_));
  NAND2_X1   g0402(.A1(new_n206_), .A2(new_n186_), .ZN(new_n452_));
  NAND2_X1   g0403(.A1(new_n452_), .A2(new_n201_), .ZN(new_n453_));
  NOR2_X1    g0404(.A1(new_n199_), .A2(new_n239_), .ZN(new_n454_));
  NAND3_X1   g0405(.A1(new_n454_), .A2(new_n189_), .A3(new_n255_), .ZN(new_n455_));
  NAND4_X1   g0406(.A1(new_n352_), .A2(new_n128_), .A3(new_n131_), .A4(new_n121_), .ZN(new_n456_));
  NAND3_X1   g0407(.A1(new_n350_), .A2(new_n381_), .A3(new_n456_), .ZN(new_n457_));
  NOR4_X1    g0408(.A1(new_n453_), .A2(new_n457_), .A3(new_n241_), .A4(new_n455_), .ZN(new_n458_));
  NAND3_X1   g0409(.A1(new_n445_), .A2(new_n451_), .A3(new_n458_), .ZN(new_n459_));
  NAND3_X1   g0410(.A1(new_n262_), .A2(new_n166_), .A3(new_n167_), .ZN(new_n460_));
  NAND2_X1   g0411(.A1(new_n285_), .A2(new_n250_), .ZN(new_n461_));
  NOR4_X1    g0412(.A1(new_n461_), .A2(new_n460_), .A3(new_n407_), .A4(new_n310_), .ZN(new_n462_));
  NOR3_X1    g0413(.A1(new_n199_), .A2(new_n162_), .A3(new_n185_), .ZN(new_n463_));
  NOR4_X1    g0414(.A1(new_n160_), .A2(new_n197_), .A3(new_n212_), .A4(new_n463_), .ZN(new_n464_));
  NAND3_X1   g0415(.A1(new_n298_), .A2(new_n137_), .A3(new_n159_), .ZN(new_n465_));
  NAND2_X1   g0416(.A1(new_n214_), .A2(new_n465_), .ZN(new_n466_));
  NOR3_X1    g0417(.A1(new_n466_), .A2(new_n247_), .A3(new_n399_), .ZN(new_n467_));
  NOR4_X1    g0418(.A1(new_n229_), .A2(new_n155_), .A3(new_n193_), .A4(new_n64_), .ZN(new_n468_));
  NOR2_X1    g0419(.A1(new_n468_), .A2(new_n375_), .ZN(new_n469_));
  NAND4_X1   g0420(.A1(new_n462_), .A2(new_n467_), .A3(new_n464_), .A4(new_n469_), .ZN(new_n470_));
  NAND4_X1   g0421(.A1(new_n361_), .A2(new_n388_), .A3(new_n292_), .A4(new_n420_), .ZN(new_n471_));
  INV_X1     g0422(.I(new_n471_), .ZN(new_n472_));
  NAND2_X1   g0423(.A1(new_n316_), .A2(new_n150_), .ZN(new_n473_));
  NOR4_X1    g0424(.A1(new_n160_), .A2(new_n366_), .A3(new_n282_), .A4(new_n473_), .ZN(new_n474_));
  NOR3_X1    g0425(.A1(new_n291_), .A2(new_n162_), .A3(new_n102_), .ZN(new_n475_));
  NOR3_X1    g0426(.A1(new_n292_), .A2(new_n363_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1   g0427(.A1(new_n149_), .A2(new_n159_), .A3(new_n137_), .ZN(new_n477_));
  NAND3_X1   g0428(.A1(new_n149_), .A2(new_n128_), .A3(new_n131_), .ZN(new_n478_));
  AOI21_X1   g0429(.A1(new_n477_), .A2(new_n478_), .B(new_n78_), .ZN(new_n479_));
  NOR2_X1    g0430(.A1(new_n479_), .A2(new_n243_), .ZN(new_n480_));
  NAND4_X1   g0431(.A1(new_n472_), .A2(new_n474_), .A3(new_n476_), .A4(new_n480_), .ZN(new_n481_));
  NAND3_X1   g0432(.A1(new_n449_), .A2(new_n201_), .A3(new_n253_), .ZN(new_n482_));
  NAND2_X1   g0433(.A1(new_n301_), .A2(new_n367_), .ZN(new_n483_));
  NOR2_X1    g0434(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND4_X1   g0435(.A1(new_n118_), .A2(new_n280_), .A3(new_n137_), .A4(new_n121_), .ZN(new_n485_));
  NAND3_X1   g0436(.A1(new_n227_), .A2(new_n485_), .A3(new_n424_), .ZN(new_n486_));
  NOR4_X1    g0437(.A1(new_n486_), .A2(new_n227_), .A3(new_n373_), .A4(new_n395_), .ZN(new_n487_));
  NAND2_X1   g0438(.A1(new_n487_), .A2(new_n484_), .ZN(new_n488_));
  NOR4_X1    g0439(.A1(new_n459_), .A2(new_n481_), .A3(new_n470_), .A4(new_n488_), .ZN(new_n489_));
  OR2_X2     g0440(.A1(new_n429_), .A2(new_n489_), .Z(new_n490_));
  NAND2_X1   g0441(.A1(new_n490_), .A2(new_n438_), .ZN(new_n491_));
  OR2_X2     g0442(.A1(new_n490_), .A2(new_n438_), .Z(new_n492_));
  XNOR2_X1   g0443(.A1(new_n489_), .A2(new_n371_), .ZN(new_n493_));
  NAND4_X1   g0444(.A1(new_n492_), .A2(new_n429_), .A3(new_n491_), .A4(new_n493_), .ZN(new_n494_));
  XNOR2_X1   g0445(.A1(new_n494_), .A2(new_n272_), .ZN(new_n495_));
  INV_X1     g0446(.I(new_n495_), .ZN(new_n496_));
  NOR3_X1    g0447(.A1(new_n227_), .A2(new_n388_), .A3(new_n326_), .ZN(new_n497_));
  NOR2_X1    g0448(.A1(new_n205_), .A2(new_n404_), .ZN(new_n498_));
  NOR2_X1    g0449(.A1(new_n388_), .A2(new_n319_), .ZN(new_n499_));
  NOR2_X1    g0450(.A1(new_n233_), .A2(new_n475_), .ZN(new_n500_));
  NAND4_X1   g0451(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .A4(new_n500_), .ZN(new_n501_));
  NOR3_X1    g0452(.A1(new_n322_), .A2(new_n102_), .A3(new_n109_), .ZN(new_n502_));
  OAI21_X1   g0453(.A1(new_n502_), .A2(new_n315_), .B(new_n64_), .ZN(new_n503_));
  NOR3_X1    g0454(.A1(new_n385_), .A2(new_n317_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1     g0455(.I(new_n389_), .ZN(new_n505_));
  NOR2_X1    g0456(.A1(new_n326_), .A2(new_n329_), .ZN(new_n506_));
  NAND4_X1   g0457(.A1(new_n505_), .A2(new_n506_), .A3(new_n366_), .A4(new_n398_), .ZN(new_n507_));
  INV_X1     g0458(.I(new_n507_), .ZN(new_n508_));
  NAND2_X1   g0459(.A1(new_n508_), .A2(new_n504_), .ZN(new_n509_));
  NOR3_X1    g0460(.A1(new_n412_), .A2(new_n149_), .A3(new_n239_), .ZN(new_n510_));
  NOR3_X1    g0461(.A1(new_n195_), .A2(new_n412_), .A3(new_n149_), .ZN(new_n511_));
  NOR2_X1    g0462(.A1(new_n511_), .A2(new_n510_), .ZN(new_n512_));
  NAND2_X1   g0463(.A1(new_n280_), .A2(new_n128_), .ZN(new_n513_));
  NOR2_X1    g0464(.A1(new_n513_), .A2(new_n291_), .ZN(new_n514_));
  NOR2_X1    g0465(.A1(new_n303_), .A2(new_n239_), .ZN(new_n515_));
  NAND3_X1   g0466(.A1(new_n514_), .A2(new_n375_), .A3(new_n515_), .ZN(new_n516_));
  NOR2_X1    g0467(.A1(new_n195_), .A2(new_n303_), .ZN(new_n517_));
  NAND3_X1   g0468(.A1(new_n363_), .A2(new_n338_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1   g0469(.A1(new_n202_), .A2(new_n316_), .ZN(new_n519_));
  NAND3_X1   g0470(.A1(new_n367_), .A2(new_n519_), .A3(new_n420_), .ZN(new_n520_));
  NOR3_X1    g0471(.A1(new_n516_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n521_));
  NOR3_X1    g0472(.A1(new_n78_), .A2(new_n91_), .A3(new_n239_), .ZN(new_n522_));
  NOR2_X1    g0473(.A1(new_n233_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1   g0474(.A1(new_n521_), .A2(new_n512_), .A3(new_n523_), .ZN(new_n524_));
  NOR3_X1    g0475(.A1(new_n509_), .A2(new_n524_), .A3(new_n501_), .ZN(new_n525_));
  NOR2_X1    g0476(.A1(new_n359_), .A2(new_n420_), .ZN(new_n526_));
  NAND4_X1   g0477(.A1(new_n526_), .A2(new_n292_), .A3(new_n383_), .A4(new_n421_), .ZN(new_n527_));
  NAND3_X1   g0478(.A1(new_n128_), .A2(new_n131_), .A3(new_n121_), .ZN(new_n528_));
  NOR4_X1    g0479(.A1(new_n528_), .A2(new_n121_), .A3(new_n195_), .A4(new_n322_), .ZN(new_n529_));
  NAND2_X1   g0480(.A1(new_n529_), .A2(new_n323_), .ZN(new_n530_));
  NOR2_X1    g0481(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1   g0482(.A1(new_n531_), .A2(new_n314_), .ZN(new_n532_));
  INV_X1     g0483(.I(new_n532_), .ZN(new_n533_));
  NAND2_X1   g0484(.A1(new_n525_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1    g0485(.A1(new_n156_), .A2(new_n292_), .ZN(new_n535_));
  NAND3_X1   g0486(.A1(new_n535_), .A2(new_n523_), .A3(new_n347_), .ZN(new_n536_));
  NAND4_X1   g0487(.A1(new_n216_), .A2(new_n137_), .A3(new_n149_), .A4(new_n159_), .ZN(new_n537_));
  NAND2_X1   g0488(.A1(new_n537_), .A2(new_n151_), .ZN(new_n538_));
  NOR3_X1    g0489(.A1(new_n249_), .A2(new_n91_), .A3(new_n412_), .ZN(new_n539_));
  NOR2_X1    g0490(.A1(new_n256_), .A2(new_n151_), .ZN(new_n540_));
  NAND2_X1   g0491(.A1(new_n540_), .A2(new_n539_), .ZN(new_n541_));
  NOR4_X1    g0492(.A1(new_n536_), .A2(new_n541_), .A3(new_n425_), .A4(new_n538_), .ZN(new_n542_));
  NAND2_X1   g0493(.A1(new_n388_), .A2(new_n230_), .ZN(new_n543_));
  NOR3_X1    g0494(.A1(new_n543_), .A2(new_n160_), .A3(new_n442_), .ZN(new_n544_));
  NAND2_X1   g0495(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NOR3_X1    g0496(.A1(new_n211_), .A2(new_n412_), .A3(new_n91_), .ZN(new_n546_));
  NAND2_X1   g0497(.A1(new_n216_), .A2(new_n149_), .ZN(new_n547_));
  NOR2_X1    g0498(.A1(new_n547_), .A2(new_n171_), .ZN(new_n548_));
  NAND4_X1   g0499(.A1(new_n548_), .A2(new_n205_), .A3(new_n313_), .A4(new_n546_), .ZN(new_n549_));
  NOR4_X1    g0500(.A1(new_n545_), .A2(new_n501_), .A3(new_n509_), .A4(new_n549_), .ZN(new_n550_));
  NOR2_X1    g0501(.A1(new_n534_), .A2(new_n550_), .ZN(new_n551_));
  NOR4_X1    g0502(.A1(new_n532_), .A2(new_n509_), .A3(new_n524_), .A4(new_n501_), .ZN(new_n552_));
  NOR3_X1    g0503(.A1(new_n511_), .A2(new_n510_), .A3(new_n363_), .ZN(new_n553_));
  NOR3_X1    g0504(.A1(new_n417_), .A2(new_n156_), .A3(new_n292_), .ZN(new_n554_));
  NOR4_X1    g0505(.A1(new_n538_), .A2(new_n151_), .A3(new_n256_), .A4(new_n381_), .ZN(new_n555_));
  NAND4_X1   g0506(.A1(new_n555_), .A2(new_n553_), .A3(new_n523_), .A4(new_n554_), .ZN(new_n556_));
  NOR4_X1    g0507(.A1(new_n556_), .A2(new_n160_), .A3(new_n442_), .A4(new_n543_), .ZN(new_n557_));
  NOR3_X1    g0508(.A1(new_n509_), .A2(new_n501_), .A3(new_n549_), .ZN(new_n558_));
  NAND2_X1   g0509(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1    g0510(.A1(new_n559_), .A2(new_n552_), .ZN(new_n560_));
  OAI21_X1   g0511(.A1(new_n560_), .A2(new_n551_), .B(new_n266_), .ZN(new_n561_));
  INV_X1     g0512(.I(new_n561_), .ZN(new_n562_));
  NOR2_X1    g0513(.A1(new_n559_), .A2(new_n534_), .ZN(new_n563_));
  NOR2_X1    g0514(.A1(new_n550_), .A2(new_n552_), .ZN(new_n564_));
  NOR3_X1    g0515(.A1(new_n563_), .A2(new_n564_), .A3(new_n266_), .ZN(new_n565_));
  INV_X1     g0516(.I(new_n266_), .ZN(new_n566_));
  AOI21_X1   g0517(.A1(new_n566_), .A2(new_n564_), .B(new_n563_), .ZN(new_n567_));
  NAND2_X1   g0518(.A1(new_n567_), .A2(new_n270_), .ZN(new_n568_));
  NAND2_X1   g0519(.A1(new_n550_), .A2(new_n552_), .ZN(new_n569_));
  NOR2_X1    g0520(.A1(new_n569_), .A2(new_n566_), .ZN(new_n570_));
  NOR2_X1    g0521(.A1(new_n570_), .A2(new_n564_), .ZN(new_n571_));
  INV_X1     g0522(.I(new_n571_), .ZN(new_n572_));
  OAI21_X1   g0523(.A1(new_n572_), .A2(new_n270_), .B(new_n568_), .ZN(new_n573_));
  AOI21_X1   g0524(.A1(new_n73_), .A2(new_n62_), .B(\a[10] ), .ZN(new_n574_));
  AND3_X2    g0525(.A1(new_n73_), .A2(\a[10] ), .A3(new_n62_), .Z(new_n575_));
  NOR2_X1    g0526(.A1(new_n575_), .A2(new_n574_), .ZN(new_n576_));
  INV_X1     g0527(.I(new_n576_), .ZN(new_n577_));
  NAND3_X1   g0528(.A1(new_n573_), .A2(new_n565_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1   g0529(.A1(new_n559_), .A2(new_n534_), .ZN(new_n579_));
  NAND3_X1   g0530(.A1(new_n579_), .A2(new_n569_), .A3(new_n566_), .ZN(new_n580_));
  NAND3_X1   g0531(.A1(new_n573_), .A2(new_n580_), .A3(new_n576_), .ZN(new_n581_));
  NAND2_X1   g0532(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1   g0533(.A1(new_n582_), .A2(new_n562_), .ZN(new_n583_));
  INV_X1     g0534(.I(new_n459_), .ZN(new_n584_));
  NAND3_X1   g0535(.A1(new_n480_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n585_));
  NOR4_X1    g0536(.A1(new_n488_), .A2(new_n470_), .A3(new_n471_), .A4(new_n585_), .ZN(new_n586_));
  NAND2_X1   g0537(.A1(new_n586_), .A2(new_n584_), .ZN(new_n587_));
  NOR2_X1    g0538(.A1(new_n160_), .A2(new_n221_), .ZN(new_n588_));
  NAND3_X1   g0539(.A1(new_n298_), .A2(new_n137_), .A3(new_n280_), .ZN(new_n589_));
  NOR4_X1    g0540(.A1(new_n132_), .A2(new_n589_), .A3(new_n353_), .A4(new_n416_), .ZN(new_n590_));
  NAND4_X1   g0541(.A1(new_n590_), .A2(new_n205_), .A3(new_n588_), .A4(new_n548_), .ZN(new_n591_));
  NOR2_X1    g0542(.A1(new_n243_), .A2(new_n463_), .ZN(new_n592_));
  NAND2_X1   g0543(.A1(new_n166_), .A2(new_n316_), .ZN(new_n593_));
  NOR2_X1    g0544(.A1(new_n593_), .A2(new_n345_), .ZN(new_n594_));
  NAND4_X1   g0545(.A1(new_n594_), .A2(new_n592_), .A3(new_n442_), .A4(new_n539_), .ZN(new_n595_));
  NOR3_X1    g0546(.A1(new_n110_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n596_));
  NOR2_X1    g0547(.A1(new_n468_), .A2(new_n200_), .ZN(new_n597_));
  NAND4_X1   g0548(.A1(new_n387_), .A2(new_n596_), .A3(new_n391_), .A4(new_n597_), .ZN(new_n598_));
  NOR3_X1    g0549(.A1(new_n598_), .A2(new_n591_), .A3(new_n595_), .ZN(new_n599_));
  NOR2_X1    g0550(.A1(new_n110_), .A2(new_n329_), .ZN(new_n600_));
  NAND3_X1   g0551(.A1(new_n600_), .A2(new_n205_), .A3(new_n313_), .ZN(new_n601_));
  NOR3_X1    g0552(.A1(new_n195_), .A2(new_n412_), .A3(new_n91_), .ZN(new_n602_));
  NOR2_X1    g0553(.A1(new_n602_), .A2(new_n363_), .ZN(new_n603_));
  NAND4_X1   g0554(.A1(new_n603_), .A2(new_n401_), .A3(new_n232_), .A4(new_n326_), .ZN(new_n604_));
  NOR2_X1    g0555(.A1(new_n468_), .A2(new_n197_), .ZN(new_n605_));
  NAND4_X1   g0556(.A1(new_n605_), .A2(new_n407_), .A3(new_n332_), .A4(new_n409_), .ZN(new_n606_));
  NOR4_X1    g0557(.A1(new_n604_), .A2(new_n606_), .A3(new_n601_), .A4(new_n405_), .ZN(new_n607_));
  NAND4_X1   g0558(.A1(new_n352_), .A2(new_n337_), .A3(new_n131_), .A4(new_n64_), .ZN(new_n608_));
  NAND4_X1   g0559(.A1(new_n352_), .A2(new_n337_), .A3(new_n131_), .A4(new_n121_), .ZN(new_n609_));
  NOR3_X1    g0560(.A1(new_n589_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NOR2_X1    g0561(.A1(new_n156_), .A2(new_n228_), .ZN(new_n611_));
  NAND4_X1   g0562(.A1(new_n553_), .A2(new_n611_), .A3(new_n610_), .A4(new_n277_), .ZN(new_n612_));
  NOR4_X1    g0563(.A1(new_n612_), .A2(new_n414_), .A3(new_n415_), .A4(new_n418_), .ZN(new_n613_));
  NAND3_X1   g0564(.A1(new_n599_), .A2(new_n613_), .A3(new_n607_), .ZN(new_n614_));
  NAND2_X1   g0565(.A1(new_n371_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1     g0566(.I(new_n615_), .ZN(new_n616_));
  OAI21_X1   g0567(.A1(new_n262_), .A2(new_n186_), .B(new_n140_), .ZN(new_n617_));
  NAND4_X1   g0568(.A1(new_n617_), .A2(new_n233_), .A3(new_n447_), .A4(new_n522_), .ZN(new_n618_));
  NOR4_X1    g0569(.A1(new_n412_), .A2(new_n162_), .A3(new_n91_), .A4(new_n185_), .ZN(new_n619_));
  NAND3_X1   g0570(.A1(new_n619_), .A2(new_n160_), .A3(new_n367_), .ZN(new_n620_));
  NOR2_X1    g0571(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1   g0572(.A1(new_n190_), .A2(new_n315_), .B(new_n140_), .ZN(new_n622_));
  NAND2_X1   g0573(.A1(new_n622_), .A2(new_n219_), .ZN(new_n623_));
  NAND2_X1   g0574(.A1(new_n519_), .A2(new_n367_), .ZN(new_n624_));
  NAND2_X1   g0575(.A1(new_n206_), .A2(new_n244_), .ZN(new_n625_));
  NOR4_X1    g0576(.A1(new_n623_), .A2(new_n301_), .A3(new_n624_), .A4(new_n625_), .ZN(new_n626_));
  NOR2_X1    g0577(.A1(new_n277_), .A2(new_n273_), .ZN(new_n627_));
  NAND4_X1   g0578(.A1(new_n621_), .A2(new_n626_), .A3(new_n300_), .A4(new_n627_), .ZN(new_n628_));
  INV_X1     g0579(.I(new_n324_), .ZN(new_n629_));
  NOR2_X1    g0580(.A1(new_n331_), .A2(new_n228_), .ZN(new_n630_));
  AND3_X2    g0581(.A1(new_n630_), .A2(new_n330_), .A3(new_n404_), .Z(new_n631_));
  INV_X1     g0582(.I(new_n348_), .ZN(new_n632_));
  NAND4_X1   g0583(.A1(new_n632_), .A2(new_n631_), .A3(new_n327_), .A4(new_n342_), .ZN(new_n633_));
  NOR2_X1    g0584(.A1(new_n362_), .A2(new_n358_), .ZN(new_n634_));
  NAND3_X1   g0585(.A1(new_n190_), .A2(new_n146_), .A3(new_n149_), .ZN(new_n635_));
  NAND2_X1   g0586(.A1(new_n207_), .A2(new_n250_), .ZN(new_n636_));
  NAND2_X1   g0587(.A1(new_n230_), .A2(new_n292_), .ZN(new_n637_));
  NOR4_X1    g0588(.A1(new_n636_), .A2(new_n637_), .A3(new_n398_), .A4(new_n635_), .ZN(new_n638_));
  NAND3_X1   g0589(.A1(new_n634_), .A2(new_n354_), .A3(new_n638_), .ZN(new_n639_));
  NOR4_X1    g0590(.A1(new_n629_), .A2(new_n628_), .A3(new_n633_), .A4(new_n639_), .ZN(new_n640_));
  NAND2_X1   g0591(.A1(new_n640_), .A2(new_n428_), .ZN(new_n641_));
  INV_X1     g0592(.I(new_n641_), .ZN(new_n642_));
  AOI21_X1   g0593(.A1(new_n435_), .A2(new_n62_), .B(\a[13] ), .ZN(new_n643_));
  NOR3_X1    g0594(.A1(new_n60_), .A2(new_n430_), .A3(\a[22] ), .ZN(new_n644_));
  NOR2_X1    g0595(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR4_X1    g0596(.A1(new_n642_), .A2(new_n438_), .A3(new_n587_), .A4(new_n616_), .ZN(new_n646_));
  INV_X1     g0597(.I(new_n646_), .ZN(new_n647_));
  NAND2_X1   g0598(.A1(new_n583_), .A2(new_n647_), .ZN(new_n648_));
  NOR3_X1    g0599(.A1(new_n276_), .A2(new_n195_), .A3(new_n121_), .ZN(new_n649_));
  NOR2_X1    g0600(.A1(new_n589_), .A2(new_n398_), .ZN(new_n650_));
  NAND4_X1   g0601(.A1(new_n650_), .A2(new_n196_), .A3(new_n212_), .A4(new_n649_), .ZN(new_n651_));
  NOR2_X1    g0602(.A1(new_n347_), .A2(new_n602_), .ZN(new_n652_));
  INV_X1     g0603(.I(new_n652_), .ZN(new_n653_));
  OAI21_X1   g0604(.A1(new_n190_), .A2(new_n186_), .B(new_n167_), .ZN(new_n654_));
  NAND2_X1   g0605(.A1(new_n654_), .A2(new_n363_), .ZN(new_n655_));
  NOR3_X1    g0606(.A1(new_n651_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  NOR4_X1    g0607(.A1(new_n452_), .A2(new_n201_), .A3(new_n424_), .A4(new_n311_), .ZN(new_n657_));
  NAND3_X1   g0608(.A1(new_n221_), .A2(new_n367_), .A3(new_n416_), .ZN(new_n658_));
  NAND4_X1   g0609(.A1(new_n468_), .A2(new_n439_), .A3(new_n463_), .A4(new_n240_), .ZN(new_n659_));
  NAND2_X1   g0610(.A1(new_n366_), .A2(new_n537_), .ZN(new_n660_));
  NOR3_X1    g0611(.A1(new_n659_), .A2(new_n660_), .A3(new_n658_), .ZN(new_n661_));
  NAND3_X1   g0612(.A1(new_n656_), .A2(new_n657_), .A3(new_n661_), .ZN(new_n662_));
  NOR2_X1    g0613(.A1(new_n662_), .A2(new_n628_), .ZN(new_n663_));
  NOR4_X1    g0614(.A1(new_n399_), .A2(new_n381_), .A3(new_n214_), .A4(new_n245_), .ZN(new_n664_));
  NOR2_X1    g0615(.A1(new_n218_), .A2(new_n389_), .ZN(new_n665_));
  NAND3_X1   g0616(.A1(new_n665_), .A2(new_n664_), .A3(new_n333_), .ZN(new_n666_));
  NOR3_X1    g0617(.A1(new_n666_), .A2(new_n374_), .A3(new_n319_), .ZN(new_n667_));
  NAND2_X1   g0618(.A1(new_n255_), .A2(new_n118_), .ZN(new_n668_));
  NOR4_X1    g0619(.A1(new_n391_), .A2(new_n209_), .A3(new_n668_), .A4(new_n608_), .ZN(new_n669_));
  INV_X1     g0620(.I(new_n255_), .ZN(new_n670_));
  NOR2_X1    g0621(.A1(new_n670_), .A2(new_n276_), .ZN(new_n671_));
  NOR2_X1    g0622(.A1(new_n671_), .A2(new_n228_), .ZN(new_n672_));
  NOR2_X1    g0623(.A1(new_n201_), .A2(new_n250_), .ZN(new_n673_));
  NAND3_X1   g0624(.A1(new_n669_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1     g0625(.I(new_n515_), .ZN(new_n675_));
  NAND3_X1   g0626(.A1(new_n675_), .A2(new_n256_), .A3(new_n243_), .ZN(new_n676_));
  NAND3_X1   g0627(.A1(new_n227_), .A2(new_n251_), .A3(new_n281_), .ZN(new_n677_));
  AOI21_X1   g0628(.A1(new_n151_), .A2(new_n222_), .B(new_n406_), .ZN(new_n678_));
  NOR2_X1    g0629(.A1(new_n205_), .A2(new_n110_), .ZN(new_n679_));
  NAND2_X1   g0630(.A1(new_n679_), .A2(new_n678_), .ZN(new_n680_));
  NOR4_X1    g0631(.A1(new_n674_), .A2(new_n676_), .A3(new_n680_), .A4(new_n677_), .ZN(new_n681_));
  NAND2_X1   g0632(.A1(new_n681_), .A2(new_n667_), .ZN(new_n682_));
  INV_X1     g0633(.I(new_n682_), .ZN(new_n683_));
  NAND2_X1   g0634(.A1(new_n683_), .A2(new_n663_), .ZN(new_n684_));
  NAND2_X1   g0635(.A1(new_n684_), .A2(new_n587_), .ZN(new_n685_));
  NAND4_X1   g0636(.A1(new_n309_), .A2(new_n656_), .A3(new_n657_), .A4(new_n661_), .ZN(new_n686_));
  NOR2_X1    g0637(.A1(new_n686_), .A2(new_n682_), .ZN(new_n687_));
  NAND2_X1   g0638(.A1(new_n687_), .A2(new_n489_), .ZN(new_n688_));
  NAND2_X1   g0639(.A1(new_n685_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1    g0640(.A1(new_n687_), .A2(new_n489_), .ZN(new_n690_));
  NOR2_X1    g0641(.A1(new_n690_), .A2(new_n550_), .ZN(new_n691_));
  NOR2_X1    g0642(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1   g0643(.A1(new_n685_), .A2(new_n688_), .A3(new_n559_), .ZN(new_n693_));
  NOR3_X1    g0644(.A1(new_n587_), .A2(new_n686_), .A3(new_n682_), .ZN(new_n694_));
  NOR2_X1    g0645(.A1(new_n690_), .A2(new_n694_), .ZN(new_n695_));
  NOR2_X1    g0646(.A1(new_n695_), .A2(new_n691_), .ZN(new_n696_));
  INV_X1     g0647(.I(new_n696_), .ZN(new_n697_));
  INV_X1     g0648(.I(\a[11] ), .ZN(new_n698_));
  NOR2_X1    g0649(.A1(new_n73_), .A2(\a[10] ), .ZN(new_n699_));
  OAI21_X1   g0650(.A1(new_n699_), .A2(\a[22] ), .B(new_n698_), .ZN(new_n700_));
  OR3_X2     g0651(.A1(new_n699_), .A2(new_n698_), .A3(\a[22] ), .Z(new_n701_));
  NAND2_X1   g0652(.A1(new_n701_), .A2(new_n700_), .ZN(new_n702_));
  OAI21_X1   g0653(.A1(new_n685_), .A2(new_n550_), .B(new_n688_), .ZN(new_n703_));
  NOR2_X1    g0654(.A1(new_n703_), .A2(new_n702_), .ZN(new_n704_));
  AOI21_X1   g0655(.A1(new_n697_), .A2(new_n702_), .B(new_n704_), .ZN(new_n705_));
  NOR2_X1    g0656(.A1(\a[12] ), .A2(\a[22] ), .ZN(new_n706_));
  NOR2_X1    g0657(.A1(new_n706_), .A2(new_n698_), .ZN(new_n707_));
  XNOR2_X1   g0658(.A1(new_n699_), .A2(new_n707_), .ZN(new_n708_));
  NOR3_X1    g0659(.A1(new_n705_), .A2(new_n693_), .A3(new_n708_), .ZN(new_n709_));
  NOR3_X1    g0660(.A1(new_n690_), .A2(new_n694_), .A3(new_n550_), .ZN(new_n710_));
  INV_X1     g0661(.I(new_n708_), .ZN(new_n711_));
  NOR3_X1    g0662(.A1(new_n705_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  OAI21_X1   g0663(.A1(new_n712_), .A2(new_n709_), .B(new_n692_), .ZN(new_n713_));
  INV_X1     g0664(.I(new_n713_), .ZN(new_n714_));
  NOR2_X1    g0665(.A1(new_n583_), .A2(new_n647_), .ZN(new_n715_));
  OAI21_X1   g0666(.A1(new_n714_), .A2(new_n715_), .B(new_n648_), .ZN(new_n716_));
  INV_X1     g0667(.I(new_n716_), .ZN(new_n717_));
  NAND2_X1   g0668(.A1(new_n567_), .A2(new_n576_), .ZN(new_n718_));
  OAI21_X1   g0669(.A1(new_n572_), .A2(new_n576_), .B(new_n718_), .ZN(new_n719_));
  NAND3_X1   g0670(.A1(new_n719_), .A2(new_n565_), .A3(new_n702_), .ZN(new_n720_));
  INV_X1     g0671(.I(new_n702_), .ZN(new_n721_));
  NAND3_X1   g0672(.A1(new_n719_), .A2(new_n580_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1   g0673(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1   g0674(.A1(new_n723_), .A2(new_n562_), .ZN(new_n724_));
  NOR3_X1    g0675(.A1(new_n339_), .A2(new_n306_), .A3(new_n211_), .ZN(new_n725_));
  NAND3_X1   g0676(.A1(new_n237_), .A2(new_n64_), .A3(new_n91_), .ZN(new_n726_));
  NOR3_X1    g0677(.A1(new_n547_), .A2(new_n726_), .A3(new_n171_), .ZN(new_n727_));
  NAND3_X1   g0678(.A1(new_n280_), .A2(new_n137_), .A3(new_n121_), .ZN(new_n728_));
  NOR4_X1    g0679(.A1(new_n728_), .A2(new_n193_), .A3(new_n171_), .A4(new_n121_), .ZN(new_n729_));
  NAND4_X1   g0680(.A1(new_n725_), .A2(new_n727_), .A3(new_n729_), .A4(new_n546_), .ZN(new_n730_));
  NOR4_X1    g0681(.A1(new_n217_), .A2(new_n260_), .A3(new_n211_), .A4(new_n726_), .ZN(new_n731_));
  NOR2_X1    g0682(.A1(new_n151_), .A2(new_n222_), .ZN(new_n732_));
  NAND3_X1   g0683(.A1(new_n215_), .A2(new_n118_), .A3(new_n121_), .ZN(new_n733_));
  NOR2_X1    g0684(.A1(new_n118_), .A2(new_n64_), .ZN(new_n734_));
  NAND4_X1   g0685(.A1(new_n337_), .A2(new_n280_), .A3(new_n131_), .A4(new_n137_), .ZN(new_n735_));
  NOR3_X1    g0686(.A1(new_n733_), .A2(new_n735_), .A3(new_n734_), .ZN(new_n736_));
  NOR3_X1    g0687(.A1(new_n209_), .A2(new_n353_), .A3(new_n398_), .ZN(new_n737_));
  NAND4_X1   g0688(.A1(new_n731_), .A2(new_n737_), .A3(new_n736_), .A4(new_n732_), .ZN(new_n738_));
  NOR3_X1    g0689(.A1(new_n668_), .A2(new_n473_), .A3(new_n251_), .ZN(new_n739_));
  NOR3_X1    g0690(.A1(new_n243_), .A2(new_n221_), .A3(new_n250_), .ZN(new_n740_));
  NAND3_X1   g0691(.A1(new_n740_), .A2(new_n739_), .A3(new_n277_), .ZN(new_n741_));
  NOR3_X1    g0692(.A1(new_n738_), .A2(new_n741_), .A3(new_n730_), .ZN(new_n742_));
  NOR2_X1    g0693(.A1(new_n383_), .A2(new_n517_), .ZN(new_n743_));
  NAND4_X1   g0694(.A1(new_n743_), .A2(new_n230_), .A3(new_n380_), .A4(new_n511_), .ZN(new_n744_));
  NAND3_X1   g0695(.A1(new_n337_), .A2(new_n131_), .A3(new_n64_), .ZN(new_n745_));
  NOR3_X1    g0696(.A1(new_n670_), .A2(new_n276_), .A3(new_n745_), .ZN(new_n746_));
  NAND3_X1   g0697(.A1(new_n746_), .A2(new_n654_), .A3(new_n420_), .ZN(new_n747_));
  NOR4_X1    g0698(.A1(new_n744_), .A2(new_n618_), .A3(new_n747_), .A4(new_n620_), .ZN(new_n748_));
  NAND2_X1   g0699(.A1(new_n372_), .A2(new_n160_), .ZN(new_n749_));
  NOR4_X1    g0700(.A1(new_n513_), .A2(new_n171_), .A3(new_n78_), .A4(new_n91_), .ZN(new_n750_));
  NAND2_X1   g0701(.A1(new_n159_), .A2(new_n337_), .ZN(new_n751_));
  NOR4_X1    g0702(.A1(new_n751_), .A2(new_n169_), .A3(new_n173_), .A4(new_n291_), .ZN(new_n752_));
  NAND4_X1   g0703(.A1(new_n750_), .A2(new_n752_), .A3(new_n201_), .A4(new_n381_), .ZN(new_n753_));
  NAND3_X1   g0704(.A1(new_n227_), .A2(new_n593_), .A3(new_n338_), .ZN(new_n754_));
  NOR4_X1    g0705(.A1(new_n260_), .A2(new_n199_), .A3(new_n78_), .A4(new_n91_), .ZN(new_n755_));
  NAND4_X1   g0706(.A1(new_n529_), .A2(new_n755_), .A3(new_n514_), .A4(new_n332_), .ZN(new_n756_));
  NOR4_X1    g0707(.A1(new_n753_), .A2(new_n756_), .A3(new_n749_), .A4(new_n754_), .ZN(new_n757_));
  NAND3_X1   g0708(.A1(new_n742_), .A2(new_n748_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1     g0709(.I(new_n455_), .ZN(new_n759_));
  NOR3_X1    g0710(.A1(new_n233_), .A2(new_n468_), .A3(new_n219_), .ZN(new_n760_));
  NOR4_X1    g0711(.A1(new_n243_), .A2(new_n367_), .A3(new_n345_), .A4(new_n395_), .ZN(new_n761_));
  NAND3_X1   g0712(.A1(new_n761_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n762_));
  NAND4_X1   g0713(.A1(new_n352_), .A2(new_n280_), .A3(new_n137_), .A4(new_n64_), .ZN(new_n763_));
  NAND3_X1   g0714(.A1(new_n195_), .A2(new_n121_), .A3(new_n352_), .ZN(new_n764_));
  AOI21_X1   g0715(.A1(new_n764_), .A2(new_n763_), .B(new_n260_), .ZN(new_n765_));
  NOR3_X1    g0716(.A1(new_n519_), .A2(new_n668_), .A3(new_n609_), .ZN(new_n766_));
  NOR2_X1    g0717(.A1(new_n168_), .A2(new_n160_), .ZN(new_n767_));
  NAND4_X1   g0718(.A1(new_n767_), .A2(new_n766_), .A3(new_n765_), .A4(new_n619_), .ZN(new_n768_));
  NOR3_X1    g0719(.A1(new_n156_), .A2(new_n230_), .A3(new_n416_), .ZN(new_n769_));
  NOR3_X1    g0720(.A1(new_n214_), .A2(new_n465_), .A3(new_n353_), .ZN(new_n770_));
  NOR3_X1    g0721(.A1(new_n201_), .A2(new_n366_), .A3(new_n243_), .ZN(new_n771_));
  NAND4_X1   g0722(.A1(new_n771_), .A2(new_n769_), .A3(new_n770_), .A4(new_n727_), .ZN(new_n772_));
  NOR3_X1    g0723(.A1(new_n772_), .A2(new_n762_), .A3(new_n768_), .ZN(new_n773_));
  NAND4_X1   g0724(.A1(new_n548_), .A2(new_n332_), .A3(new_n313_), .A4(new_n475_), .ZN(new_n774_));
  NOR3_X1    g0725(.A1(new_n209_), .A2(new_n608_), .A3(new_n407_), .ZN(new_n775_));
  NOR3_X1    g0726(.A1(new_n91_), .A2(new_n162_), .A3(new_n185_), .ZN(new_n776_));
  AOI22_X1   g0727(.A1(new_n167_), .A2(new_n190_), .B1(new_n776_), .B2(new_n146_), .ZN(new_n777_));
  NOR2_X1    g0728(.A1(new_n356_), .A2(new_n374_), .ZN(new_n778_));
  NAND3_X1   g0729(.A1(new_n778_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n779_));
  NAND3_X1   g0730(.A1(new_n149_), .A2(new_n131_), .A3(new_n137_), .ZN(new_n780_));
  NOR4_X1    g0731(.A1(new_n780_), .A2(new_n513_), .A3(new_n199_), .A4(new_n78_), .ZN(new_n781_));
  NOR3_X1    g0732(.A1(new_n171_), .A2(new_n199_), .A3(new_n291_), .ZN(new_n782_));
  NOR4_X1    g0733(.A1(new_n670_), .A2(new_n478_), .A3(new_n78_), .A4(new_n276_), .ZN(new_n783_));
  NAND4_X1   g0734(.A1(new_n783_), .A2(new_n781_), .A3(new_n205_), .A4(new_n782_), .ZN(new_n784_));
  NOR4_X1    g0735(.A1(new_n784_), .A2(new_n779_), .A3(new_n457_), .A4(new_n774_), .ZN(new_n785_));
  OAI21_X1   g0736(.A1(new_n262_), .A2(new_n190_), .B(new_n206_), .ZN(new_n786_));
  NAND3_X1   g0737(.A1(new_n786_), .A2(new_n388_), .A3(new_n218_), .ZN(new_n787_));
  NOR3_X1    g0738(.A1(new_n156_), .A2(new_n273_), .A3(new_n383_), .ZN(new_n788_));
  NOR3_X1    g0739(.A1(new_n277_), .A2(new_n364_), .A3(new_n200_), .ZN(new_n789_));
  NAND2_X1   g0740(.A1(new_n789_), .A2(new_n788_), .ZN(new_n790_));
  NOR3_X1    g0741(.A1(new_n260_), .A2(new_n91_), .A3(new_n412_), .ZN(new_n791_));
  NOR2_X1    g0742(.A1(new_n201_), .A2(new_n222_), .ZN(new_n792_));
  NAND4_X1   g0743(.A1(new_n792_), .A2(new_n319_), .A3(new_n409_), .A4(new_n791_), .ZN(new_n793_));
  NOR3_X1    g0744(.A1(new_n413_), .A2(new_n511_), .A3(new_n196_), .ZN(new_n794_));
  NOR3_X1    g0745(.A1(new_n306_), .A2(new_n171_), .A3(new_n211_), .ZN(new_n795_));
  NAND3_X1   g0746(.A1(new_n794_), .A2(new_n526_), .A3(new_n795_), .ZN(new_n796_));
  NOR4_X1    g0747(.A1(new_n796_), .A2(new_n790_), .A3(new_n793_), .A4(new_n787_), .ZN(new_n797_));
  NAND3_X1   g0748(.A1(new_n773_), .A2(new_n797_), .A3(new_n785_), .ZN(new_n798_));
  NAND2_X1   g0749(.A1(new_n798_), .A2(new_n758_), .ZN(new_n799_));
  NAND2_X1   g0750(.A1(new_n799_), .A2(new_n614_), .ZN(new_n800_));
  NOR2_X1    g0751(.A1(new_n268_), .A2(new_n267_), .ZN(new_n801_));
  XNOR2_X1   g0752(.A1(new_n94_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1     g0753(.I(new_n802_), .ZN(new_n803_));
  NOR2_X1    g0754(.A1(new_n266_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1    g0755(.A1(new_n94_), .A2(\a[22] ), .ZN(new_n805_));
  INV_X1     g0756(.I(new_n805_), .ZN(new_n806_));
  NOR2_X1    g0757(.A1(new_n267_), .A2(\a[22] ), .ZN(new_n807_));
  AOI22_X1   g0758(.A1(new_n806_), .A2(new_n267_), .B1(new_n52_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1     g0759(.I(new_n808_), .ZN(new_n809_));
  AOI21_X1   g0760(.A1(new_n266_), .A2(new_n803_), .B(new_n809_), .ZN(new_n810_));
  NOR3_X1    g0761(.A1(new_n810_), .A2(new_n800_), .A3(new_n804_), .ZN(new_n811_));
  NAND2_X1   g0762(.A1(new_n724_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1    g0763(.A1(new_n724_), .A2(new_n811_), .ZN(new_n813_));
  INV_X1     g0764(.I(new_n813_), .ZN(new_n814_));
  AOI21_X1   g0765(.A1(new_n812_), .A2(new_n814_), .B(new_n717_), .ZN(new_n815_));
  XNOR2_X1   g0766(.A1(new_n724_), .A2(new_n811_), .ZN(new_n816_));
  NOR2_X1    g0767(.A1(new_n816_), .A2(new_n716_), .ZN(new_n817_));
  NOR2_X1    g0768(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  NOR2_X1    g0769(.A1(new_n266_), .A2(new_n809_), .ZN(new_n819_));
  NOR3_X1    g0770(.A1(new_n169_), .A2(new_n91_), .A3(new_n412_), .ZN(new_n820_));
  NOR2_X1    g0771(.A1(new_n528_), .A2(new_n322_), .ZN(new_n821_));
  NOR3_X1    g0772(.A1(new_n539_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND4_X1   g0773(.A1(new_n822_), .A2(new_n775_), .A3(new_n777_), .A4(new_n778_), .ZN(new_n823_));
  NAND4_X1   g0774(.A1(new_n140_), .A2(new_n298_), .A3(new_n131_), .A4(new_n137_), .ZN(new_n824_));
  NOR3_X1    g0775(.A1(new_n824_), .A2(new_n201_), .A3(new_n203_), .ZN(new_n825_));
  NAND4_X1   g0776(.A1(new_n237_), .A2(new_n149_), .A3(new_n131_), .A4(new_n137_), .ZN(new_n826_));
  NOR4_X1    g0777(.A1(new_n256_), .A2(new_n366_), .A3(new_n121_), .A4(new_n826_), .ZN(new_n827_));
  NAND4_X1   g0778(.A1(new_n827_), .A2(new_n825_), .A3(new_n725_), .A4(new_n727_), .ZN(new_n828_));
  NOR4_X1    g0779(.A1(new_n277_), .A2(new_n201_), .A3(new_n313_), .A4(new_n217_), .ZN(new_n829_));
  NAND3_X1   g0780(.A1(new_n829_), .A2(new_n789_), .A3(new_n788_), .ZN(new_n830_));
  NOR3_X1    g0781(.A1(new_n635_), .A2(new_n201_), .A3(new_n222_), .ZN(new_n831_));
  NOR3_X1    g0782(.A1(new_n160_), .A2(new_n281_), .A3(new_n537_), .ZN(new_n832_));
  OAI22_X1   g0783(.A1(new_n728_), .A2(new_n322_), .B1(new_n211_), .B2(new_n291_), .ZN(new_n833_));
  NAND3_X1   g0784(.A1(new_n262_), .A2(new_n206_), .A3(new_n190_), .ZN(new_n834_));
  NOR2_X1    g0785(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1   g0786(.A1(new_n835_), .A2(new_n831_), .A3(new_n832_), .A4(new_n794_), .ZN(new_n836_));
  NOR4_X1    g0787(.A1(new_n836_), .A2(new_n823_), .A3(new_n828_), .A4(new_n830_), .ZN(new_n837_));
  NAND3_X1   g0788(.A1(new_n758_), .A2(new_n773_), .A3(new_n837_), .ZN(new_n838_));
  NAND3_X1   g0789(.A1(new_n475_), .A2(new_n206_), .A3(new_n190_), .ZN(new_n839_));
  NAND4_X1   g0790(.A1(new_n262_), .A2(new_n340_), .A3(new_n146_), .A4(new_n91_), .ZN(new_n840_));
  NAND2_X1   g0791(.A1(new_n228_), .A2(new_n196_), .ZN(new_n841_));
  NOR4_X1    g0792(.A1(new_n841_), .A2(new_n840_), .A3(new_n839_), .A4(new_n341_), .ZN(new_n842_));
  NAND2_X1   g0793(.A1(new_n193_), .A2(new_n121_), .ZN(new_n843_));
  NAND4_X1   g0794(.A1(new_n273_), .A2(new_n190_), .A3(new_n186_), .A4(new_n843_), .ZN(new_n844_));
  NAND3_X1   g0795(.A1(new_n363_), .A2(new_n325_), .A3(new_n376_), .ZN(new_n845_));
  NOR4_X1    g0796(.A1(new_n845_), .A2(new_n844_), .A3(new_n151_), .A4(new_n222_), .ZN(new_n846_));
  NOR4_X1    g0797(.A1(new_n322_), .A2(new_n64_), .A3(new_n102_), .A4(new_n109_), .ZN(new_n847_));
  NAND3_X1   g0798(.A1(new_n219_), .A2(new_n360_), .A3(new_n847_), .ZN(new_n848_));
  NAND4_X1   g0799(.A1(new_n315_), .A2(new_n776_), .A3(new_n140_), .A4(new_n146_), .ZN(new_n849_));
  NOR4_X1    g0800(.A1(new_n848_), .A2(new_n221_), .A3(new_n849_), .A4(new_n449_), .ZN(new_n850_));
  NAND4_X1   g0801(.A1(new_n842_), .A2(new_n846_), .A3(new_n850_), .A4(new_n731_), .ZN(new_n851_));
  OAI22_X1   g0802(.A1(new_n169_), .A2(new_n291_), .B1(new_n195_), .B2(new_n303_), .ZN(new_n852_));
  NOR4_X1    g0803(.A1(new_n852_), .A2(new_n442_), .A3(new_n366_), .A4(new_n424_), .ZN(new_n853_));
  NOR4_X1    g0804(.A1(new_n191_), .A2(new_n247_), .A3(new_n256_), .A4(new_n608_), .ZN(new_n854_));
  NAND4_X1   g0805(.A1(new_n853_), .A2(new_n854_), .A3(new_n284_), .A4(new_n293_), .ZN(new_n855_));
  NOR2_X1    g0806(.A1(new_n205_), .A2(new_n156_), .ZN(new_n856_));
  NAND2_X1   g0807(.A1(new_n201_), .A2(new_n381_), .ZN(new_n857_));
  NAND3_X1   g0808(.A1(new_n238_), .A2(new_n146_), .A3(new_n776_), .ZN(new_n858_));
  NOR3_X1    g0809(.A1(new_n173_), .A2(new_n102_), .A3(new_n109_), .ZN(new_n859_));
  NAND2_X1   g0810(.A1(new_n383_), .A2(new_n859_), .ZN(new_n860_));
  NOR3_X1    g0811(.A1(new_n857_), .A2(new_n858_), .A3(new_n860_), .ZN(new_n861_));
  NOR3_X1    g0812(.A1(new_n384_), .A2(new_n413_), .A3(new_n439_), .ZN(new_n862_));
  NAND4_X1   g0813(.A1(new_n375_), .A2(new_n121_), .A3(new_n166_), .A4(new_n352_), .ZN(new_n863_));
  NAND4_X1   g0814(.A1(new_n315_), .A2(new_n140_), .A3(new_n146_), .A4(new_n149_), .ZN(new_n864_));
  NOR4_X1    g0815(.A1(new_n863_), .A2(new_n299_), .A3(new_n864_), .A4(new_n404_), .ZN(new_n865_));
  NAND4_X1   g0816(.A1(new_n865_), .A2(new_n861_), .A3(new_n856_), .A4(new_n862_), .ZN(new_n866_));
  NOR3_X1    g0817(.A1(new_n851_), .A2(new_n866_), .A3(new_n855_), .ZN(new_n867_));
  NAND2_X1   g0818(.A1(new_n798_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1   g0819(.A1(new_n868_), .A2(new_n838_), .B(new_n428_), .ZN(new_n869_));
  XOR2_X1    g0820(.A1(new_n428_), .A2(new_n867_), .Z(new_n870_));
  NAND3_X1   g0821(.A1(new_n870_), .A2(new_n838_), .A3(new_n868_), .ZN(new_n871_));
  AOI21_X1   g0822(.A1(new_n437_), .A2(new_n869_), .B(new_n871_), .ZN(new_n872_));
  OAI21_X1   g0823(.A1(new_n437_), .A2(new_n869_), .B(new_n872_), .ZN(new_n873_));
  AND2_X2    g0824(.A1(new_n873_), .A2(new_n819_), .Z(new_n874_));
  INV_X1     g0825(.I(new_n645_), .ZN(new_n875_));
  NOR4_X1    g0826(.A1(new_n642_), .A2(new_n587_), .A3(new_n616_), .A4(new_n875_), .ZN(new_n876_));
  NOR2_X1    g0827(.A1(new_n873_), .A2(new_n819_), .ZN(new_n877_));
  NOR2_X1    g0828(.A1(new_n877_), .A2(new_n876_), .ZN(new_n878_));
  NOR2_X1    g0829(.A1(new_n878_), .A2(new_n874_), .ZN(new_n879_));
  XOR2_X1    g0830(.A1(new_n800_), .A2(new_n802_), .Z(new_n880_));
  NAND2_X1   g0831(.A1(new_n880_), .A2(new_n809_), .ZN(new_n881_));
  XOR2_X1    g0832(.A1(new_n881_), .A2(new_n266_), .Z(new_n882_));
  NOR2_X1    g0833(.A1(new_n879_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1     g0834(.I(new_n883_), .ZN(new_n884_));
  NAND2_X1   g0835(.A1(new_n567_), .A2(new_n802_), .ZN(new_n885_));
  OAI21_X1   g0836(.A1(new_n572_), .A2(new_n802_), .B(new_n885_), .ZN(new_n886_));
  NAND3_X1   g0837(.A1(new_n886_), .A2(new_n271_), .A3(new_n565_), .ZN(new_n887_));
  NAND3_X1   g0838(.A1(new_n886_), .A2(new_n270_), .A3(new_n580_), .ZN(new_n888_));
  NAND2_X1   g0839(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1   g0840(.A1(new_n889_), .A2(new_n562_), .ZN(new_n890_));
  NOR3_X1    g0841(.A1(new_n211_), .A2(new_n193_), .A3(new_n64_), .ZN(new_n891_));
  INV_X1     g0842(.I(new_n891_), .ZN(new_n892_));
  NOR4_X1    g0843(.A1(new_n892_), .A2(new_n243_), .A3(new_n635_), .A4(new_n281_), .ZN(new_n893_));
  NAND2_X1   g0844(.A1(new_n228_), .A2(new_n468_), .ZN(new_n894_));
  NOR4_X1    g0845(.A1(new_n894_), .A2(new_n479_), .A3(new_n191_), .A4(new_n256_), .ZN(new_n895_));
  NAND2_X1   g0846(.A1(new_n424_), .A2(new_n301_), .ZN(new_n896_));
  NAND2_X1   g0847(.A1(new_n413_), .A2(new_n206_), .ZN(new_n897_));
  AOI21_X1   g0848(.A1(new_n388_), .A2(new_n262_), .B(new_n340_), .ZN(new_n898_));
  NOR4_X1    g0849(.A1(new_n446_), .A2(new_n898_), .A3(new_n897_), .A4(new_n896_), .ZN(new_n899_));
  NAND4_X1   g0850(.A1(new_n206_), .A2(new_n340_), .A3(new_n190_), .A4(new_n202_), .ZN(new_n900_));
  NOR4_X1    g0851(.A1(new_n900_), .A2(new_n156_), .A3(new_n205_), .A4(new_n399_), .ZN(new_n901_));
  NAND4_X1   g0852(.A1(new_n899_), .A2(new_n895_), .A3(new_n893_), .A4(new_n901_), .ZN(new_n902_));
  NOR2_X1    g0853(.A1(new_n313_), .A2(new_n602_), .ZN(new_n903_));
  NAND4_X1   g0854(.A1(new_n388_), .A2(new_n319_), .A3(new_n196_), .A4(new_n273_), .ZN(new_n904_));
  NOR3_X1    g0855(.A1(new_n904_), .A2(new_n636_), .A3(new_n903_), .ZN(new_n905_));
  OAI21_X1   g0856(.A1(new_n110_), .A2(new_n468_), .B(new_n197_), .ZN(new_n906_));
  NAND3_X1   g0857(.A1(new_n449_), .A2(new_n390_), .A3(new_n250_), .ZN(new_n907_));
  NAND3_X1   g0858(.A1(new_n228_), .A2(new_n383_), .A3(new_n439_), .ZN(new_n908_));
  NOR3_X1    g0859(.A1(new_n907_), .A2(new_n906_), .A3(new_n908_), .ZN(new_n909_));
  OAI21_X1   g0860(.A1(new_n169_), .A2(new_n322_), .B(new_n171_), .ZN(new_n910_));
  NAND4_X1   g0861(.A1(new_n910_), .A2(new_n205_), .A3(new_n156_), .A4(new_n359_), .ZN(new_n911_));
  INV_X1     g0862(.I(new_n911_), .ZN(new_n912_));
  NAND2_X1   g0863(.A1(new_n219_), .A2(new_n360_), .ZN(new_n913_));
  NOR4_X1    g0864(.A1(new_n246_), .A2(new_n372_), .A3(new_n913_), .A4(new_n625_), .ZN(new_n914_));
  NAND4_X1   g0865(.A1(new_n909_), .A2(new_n905_), .A3(new_n912_), .A4(new_n914_), .ZN(new_n915_));
  NAND3_X1   g0866(.A1(new_n244_), .A2(new_n352_), .A3(new_n121_), .ZN(new_n918_));
  NOR2_X1    g0867(.A1(new_n227_), .A2(new_n918_), .ZN(new_n919_));
  NOR4_X1    g0868(.A1(new_n624_), .A2(new_n396_), .A3(new_n247_), .A4(new_n503_), .ZN(new_n920_));
  NOR2_X1    g0869(.A1(new_n195_), .A2(new_n173_), .ZN(new_n921_));
  NAND3_X1   g0870(.A1(new_n326_), .A2(new_n921_), .A3(new_n240_), .ZN(new_n922_));
  NOR4_X1    g0871(.A1(new_n922_), .A2(new_n132_), .A3(new_n168_), .A4(new_n608_), .ZN(new_n923_));
  NAND3_X1   g0872(.A1(new_n920_), .A2(new_n923_), .A3(new_n919_), .ZN(new_n924_));
  NOR3_X1    g0873(.A1(new_n915_), .A2(new_n902_), .A3(new_n924_), .ZN(new_n925_));
  NAND2_X1   g0874(.A1(new_n925_), .A2(new_n798_), .ZN(new_n926_));
  NOR2_X1    g0875(.A1(new_n566_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1   g0876(.A1(new_n890_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1   g0877(.A1(new_n685_), .A2(new_n559_), .ZN(new_n929_));
  NAND2_X1   g0878(.A1(new_n929_), .A2(new_n695_), .ZN(new_n930_));
  OR2_X2     g0879(.A1(new_n703_), .A2(new_n577_), .Z(new_n931_));
  OAI21_X1   g0880(.A1(new_n576_), .A2(new_n696_), .B(new_n931_), .ZN(new_n932_));
  NAND3_X1   g0881(.A1(new_n932_), .A2(new_n710_), .A3(new_n702_), .ZN(new_n933_));
  NAND3_X1   g0882(.A1(new_n932_), .A2(new_n693_), .A3(new_n721_), .ZN(new_n934_));
  AOI21_X1   g0883(.A1(new_n933_), .A2(new_n934_), .B(new_n930_), .ZN(new_n935_));
  INV_X1     g0884(.I(new_n935_), .ZN(new_n936_));
  INV_X1     g0885(.I(new_n927_), .ZN(new_n937_));
  NAND3_X1   g0886(.A1(new_n889_), .A2(new_n562_), .A3(new_n937_), .ZN(new_n938_));
  NAND2_X1   g0887(.A1(new_n936_), .A2(new_n938_), .ZN(new_n939_));
  AND2_X2    g0888(.A1(new_n939_), .A2(new_n928_), .Z(new_n940_));
  INV_X1     g0889(.I(new_n940_), .ZN(new_n941_));
  NAND2_X1   g0890(.A1(new_n879_), .A2(new_n882_), .ZN(new_n942_));
  NAND2_X1   g0891(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1   g0892(.A1(new_n943_), .A2(new_n884_), .ZN(new_n944_));
  NOR4_X1    g0893(.A1(new_n690_), .A2(new_n559_), .A3(new_n694_), .A4(new_n875_), .ZN(new_n945_));
  INV_X1     g0894(.I(new_n945_), .ZN(new_n946_));
  NOR2_X1    g0895(.A1(new_n944_), .A2(new_n946_), .ZN(new_n947_));
  NAND2_X1   g0896(.A1(new_n944_), .A2(new_n946_), .ZN(new_n948_));
  INV_X1     g0897(.I(new_n948_), .ZN(new_n949_));
  OAI21_X1   g0898(.A1(new_n949_), .A2(new_n947_), .B(new_n818_), .ZN(new_n950_));
  INV_X1     g0899(.I(new_n818_), .ZN(new_n951_));
  INV_X1     g0900(.I(new_n947_), .ZN(new_n952_));
  NAND3_X1   g0901(.A1(new_n952_), .A2(new_n951_), .A3(new_n948_), .ZN(new_n953_));
  AOI21_X1   g0902(.A1(new_n950_), .A2(new_n953_), .B(new_n496_), .ZN(new_n954_));
  AOI21_X1   g0903(.A1(new_n952_), .A2(new_n948_), .B(new_n951_), .ZN(new_n955_));
  NOR3_X1    g0904(.A1(new_n949_), .A2(new_n818_), .A3(new_n947_), .ZN(new_n956_));
  NOR3_X1    g0905(.A1(new_n955_), .A2(new_n956_), .A3(new_n495_), .ZN(new_n957_));
  AOI21_X1   g0906(.A1(new_n884_), .A2(new_n942_), .B(new_n940_), .ZN(new_n958_));
  XNOR2_X1   g0907(.A1(new_n879_), .A2(new_n882_), .ZN(new_n959_));
  NOR2_X1    g0908(.A1(new_n941_), .A2(new_n959_), .ZN(new_n960_));
  NOR2_X1    g0909(.A1(new_n960_), .A2(new_n958_), .ZN(new_n961_));
  XOR2_X1    g0910(.A1(new_n583_), .A2(new_n647_), .Z(new_n962_));
  NAND2_X1   g0911(.A1(new_n962_), .A2(new_n714_), .ZN(new_n963_));
  INV_X1     g0912(.I(new_n648_), .ZN(new_n964_));
  OAI21_X1   g0913(.A1(new_n964_), .A2(new_n715_), .B(new_n713_), .ZN(new_n965_));
  NAND2_X1   g0914(.A1(new_n963_), .A2(new_n965_), .ZN(new_n966_));
  INV_X1     g0915(.I(new_n966_), .ZN(new_n967_));
  NOR2_X1    g0916(.A1(new_n961_), .A2(new_n967_), .ZN(new_n968_));
  NAND2_X1   g0917(.A1(new_n928_), .A2(new_n938_), .ZN(new_n969_));
  NAND2_X1   g0918(.A1(new_n969_), .A2(new_n935_), .ZN(new_n970_));
  XOR2_X1    g0919(.A1(new_n890_), .A2(new_n927_), .Z(new_n971_));
  NAND2_X1   g0920(.A1(new_n971_), .A2(new_n936_), .ZN(new_n972_));
  NAND2_X1   g0921(.A1(new_n972_), .A2(new_n970_), .ZN(new_n973_));
  OAI21_X1   g0922(.A1(new_n874_), .A2(new_n877_), .B(new_n876_), .ZN(new_n974_));
  XNOR2_X1   g0923(.A1(new_n873_), .A2(new_n819_), .ZN(new_n975_));
  OAI21_X1   g0924(.A1(new_n876_), .A2(new_n975_), .B(new_n974_), .ZN(new_n976_));
  NOR2_X1    g0925(.A1(new_n973_), .A2(new_n976_), .ZN(new_n977_));
  NAND2_X1   g0926(.A1(new_n567_), .A2(new_n808_), .ZN(new_n978_));
  OAI21_X1   g0927(.A1(new_n572_), .A2(new_n808_), .B(new_n978_), .ZN(new_n979_));
  NAND3_X1   g0928(.A1(new_n979_), .A2(new_n565_), .A3(new_n803_), .ZN(new_n980_));
  NAND3_X1   g0929(.A1(new_n979_), .A2(new_n580_), .A3(new_n802_), .ZN(new_n981_));
  NAND2_X1   g0930(.A1(new_n980_), .A2(new_n981_), .ZN(new_n982_));
  NAND2_X1   g0931(.A1(new_n982_), .A2(new_n562_), .ZN(new_n983_));
  NAND3_X1   g0932(.A1(new_n281_), .A2(new_n251_), .A3(new_n222_), .ZN(new_n984_));
  NAND4_X1   g0933(.A1(new_n232_), .A2(new_n292_), .A3(new_n383_), .A4(new_n329_), .ZN(new_n985_));
  NOR3_X1    g0934(.A1(new_n985_), .A2(new_n984_), .A3(new_n455_), .ZN(new_n986_));
  NAND3_X1   g0935(.A1(new_n421_), .A2(new_n360_), .A3(new_n304_), .ZN(new_n987_));
  NOR4_X1    g0936(.A1(new_n987_), .A2(new_n160_), .A3(new_n168_), .A4(new_n285_), .ZN(new_n988_));
  NAND3_X1   g0937(.A1(new_n160_), .A2(new_n366_), .A3(new_n220_), .ZN(new_n989_));
  NAND3_X1   g0938(.A1(new_n326_), .A2(new_n859_), .A3(new_n376_), .ZN(new_n990_));
  NOR3_X1    g0939(.A1(new_n229_), .A2(new_n162_), .A3(new_n91_), .ZN(new_n991_));
  NAND4_X1   g0940(.A1(new_n238_), .A2(new_n991_), .A3(new_n146_), .A4(new_n776_), .ZN(new_n992_));
  NOR4_X1    g0941(.A1(new_n989_), .A2(new_n840_), .A3(new_n992_), .A4(new_n990_), .ZN(new_n993_));
  NAND4_X1   g0942(.A1(new_n993_), .A2(new_n986_), .A3(new_n988_), .A4(new_n765_), .ZN(new_n994_));
  NOR2_X1    g0943(.A1(new_n840_), .A2(new_n839_), .ZN(new_n995_));
  NAND4_X1   g0944(.A1(new_n325_), .A2(new_n190_), .A3(new_n239_), .A4(new_n298_), .ZN(new_n996_));
  NAND2_X1   g0945(.A1(new_n243_), .A2(new_n416_), .ZN(new_n997_));
  OAI21_X1   g0946(.A1(new_n276_), .A2(new_n745_), .B(new_n132_), .ZN(new_n998_));
  NOR4_X1    g0947(.A1(new_n457_), .A2(new_n998_), .A3(new_n997_), .A4(new_n996_), .ZN(new_n999_));
  NAND2_X1   g0948(.A1(new_n388_), .A2(new_n463_), .ZN(new_n1000_));
  NAND4_X1   g0949(.A1(new_n991_), .A2(new_n146_), .A3(new_n189_), .A4(new_n255_), .ZN(new_n1001_));
  NOR4_X1    g0950(.A1(new_n1000_), .A2(new_n1001_), .A3(new_n372_), .A4(new_n824_), .ZN(new_n1002_));
  NAND3_X1   g0951(.A1(new_n999_), .A2(new_n1002_), .A3(new_n995_), .ZN(new_n1003_));
  NAND3_X1   g0952(.A1(new_n160_), .A2(new_n345_), .A3(new_n733_), .ZN(new_n1004_));
  NOR2_X1    g0953(.A1(new_n907_), .A2(new_n1004_), .ZN(new_n1005_));
  NOR3_X1    g0954(.A1(new_n229_), .A2(new_n91_), .A3(new_n109_), .ZN(new_n1006_));
  NAND4_X1   g0955(.A1(new_n468_), .A2(new_n238_), .A3(new_n1006_), .A4(new_n146_), .ZN(new_n1007_));
  NAND2_X1   g0956(.A1(new_n409_), .A2(new_n791_), .ZN(new_n1008_));
  NOR2_X1    g0957(.A1(new_n1008_), .A2(new_n1007_), .ZN(new_n1009_));
  NAND3_X1   g0958(.A1(new_n237_), .A2(new_n121_), .A3(new_n91_), .ZN(new_n1010_));
  OAI22_X1   g0959(.A1(new_n1010_), .A2(new_n169_), .B1(new_n728_), .B2(new_n193_), .ZN(new_n1011_));
  NOR4_X1    g0960(.A1(new_n1011_), .A2(new_n833_), .A3(new_n834_), .A4(new_n511_), .ZN(new_n1012_));
  NAND4_X1   g0961(.A1(new_n1005_), .A2(new_n1009_), .A3(new_n1012_), .A4(new_n829_), .ZN(new_n1013_));
  NOR3_X1    g0962(.A1(new_n994_), .A2(new_n1013_), .A3(new_n1003_), .ZN(new_n1014_));
  NAND2_X1   g0963(.A1(new_n1014_), .A2(new_n867_), .ZN(new_n1015_));
  OAI21_X1   g0964(.A1(new_n428_), .A2(new_n799_), .B(new_n1015_), .ZN(new_n1016_));
  OAI21_X1   g0965(.A1(new_n614_), .A2(new_n1015_), .B(new_n799_), .ZN(new_n1017_));
  INV_X1     g0966(.I(new_n1017_), .ZN(new_n1018_));
  AOI21_X1   g0967(.A1(new_n868_), .A2(new_n838_), .B(new_n614_), .ZN(new_n1019_));
  NOR2_X1    g0968(.A1(new_n1019_), .A2(new_n437_), .ZN(new_n1020_));
  NOR2_X1    g0969(.A1(new_n869_), .A2(new_n438_), .ZN(new_n1021_));
  OAI21_X1   g0970(.A1(new_n1020_), .A2(new_n1021_), .B(new_n1018_), .ZN(new_n1022_));
  OAI21_X1   g0971(.A1(new_n1020_), .A2(new_n1021_), .B(new_n875_), .ZN(new_n1023_));
  XOR2_X1    g0972(.A1(new_n1022_), .A2(new_n1023_), .Z(new_n1024_));
  NAND2_X1   g0973(.A1(new_n1024_), .A2(new_n1016_), .ZN(new_n1025_));
  NAND2_X1   g0974(.A1(new_n983_), .A2(new_n1025_), .ZN(new_n1026_));
  INV_X1     g0975(.I(new_n1026_), .ZN(new_n1027_));
  NOR2_X1    g0976(.A1(new_n703_), .A2(new_n271_), .ZN(new_n1028_));
  AOI21_X1   g0977(.A1(new_n271_), .A2(new_n697_), .B(new_n1028_), .ZN(new_n1029_));
  NOR3_X1    g0978(.A1(new_n1029_), .A2(new_n576_), .A3(new_n693_), .ZN(new_n1030_));
  NOR3_X1    g0979(.A1(new_n1029_), .A2(new_n577_), .A3(new_n710_), .ZN(new_n1031_));
  OAI21_X1   g0980(.A1(new_n1030_), .A2(new_n1031_), .B(new_n692_), .ZN(new_n1032_));
  AOI21_X1   g0981(.A1(new_n980_), .A2(new_n981_), .B(new_n561_), .ZN(new_n1033_));
  INV_X1     g0982(.I(new_n1025_), .ZN(new_n1034_));
  NAND2_X1   g0983(.A1(new_n1034_), .A2(new_n1033_), .ZN(new_n1035_));
  AOI21_X1   g0984(.A1(new_n1032_), .A2(new_n1035_), .B(new_n1027_), .ZN(new_n1036_));
  INV_X1     g0985(.I(new_n1036_), .ZN(new_n1037_));
  NAND2_X1   g0986(.A1(new_n973_), .A2(new_n976_), .ZN(new_n1038_));
  AOI21_X1   g0987(.A1(new_n1037_), .A2(new_n1038_), .B(new_n977_), .ZN(new_n1039_));
  INV_X1     g0988(.I(new_n1039_), .ZN(new_n1040_));
  NAND2_X1   g0989(.A1(new_n961_), .A2(new_n967_), .ZN(new_n1041_));
  AOI21_X1   g0990(.A1(new_n1040_), .A2(new_n1041_), .B(new_n968_), .ZN(new_n1042_));
  INV_X1     g0991(.I(new_n1042_), .ZN(new_n1043_));
  NOR3_X1    g0992(.A1(new_n954_), .A2(new_n957_), .A3(new_n1043_), .ZN(new_n1044_));
  NOR2_X1    g0993(.A1(new_n58_), .A2(\a[4] ), .ZN(new_n1045_));
  NOR2_X1    g0994(.A1(new_n1045_), .A2(\a[22] ), .ZN(new_n1046_));
  NOR2_X1    g0995(.A1(new_n1046_), .A2(\a[5] ), .ZN(new_n1047_));
  NAND2_X1   g0996(.A1(new_n62_), .A2(\a[5] ), .ZN(new_n1048_));
  NOR2_X1    g0997(.A1(new_n1045_), .A2(new_n1048_), .ZN(new_n1049_));
  NOR2_X1    g0998(.A1(new_n1047_), .A2(new_n1049_), .ZN(new_n1050_));
  INV_X1     g0999(.I(new_n1050_), .ZN(new_n1051_));
  NOR2_X1    g1000(.A1(new_n565_), .A2(new_n1051_), .ZN(new_n1052_));
  XOR2_X1    g1001(.A1(new_n550_), .A2(new_n552_), .Z(new_n1053_));
  AOI21_X1   g1002(.A1(new_n1053_), .A2(new_n266_), .B(new_n1050_), .ZN(new_n1054_));
  NOR2_X1    g1003(.A1(new_n1054_), .A2(new_n1052_), .ZN(new_n1055_));
  OAI21_X1   g1004(.A1(new_n579_), .A2(new_n266_), .B(new_n569_), .ZN(new_n1056_));
  INV_X1     g1005(.I(\a[4] ), .ZN(new_n1057_));
  NAND2_X1   g1006(.A1(new_n58_), .A2(new_n62_), .ZN(new_n1058_));
  NOR2_X1    g1007(.A1(new_n1057_), .A2(\a[22] ), .ZN(new_n1059_));
  AOI22_X1   g1008(.A1(new_n1058_), .A2(new_n1057_), .B1(new_n58_), .B2(new_n1059_), .ZN(new_n1060_));
  INV_X1     g1009(.I(new_n1060_), .ZN(new_n1061_));
  NOR2_X1    g1010(.A1(new_n1056_), .A2(new_n1061_), .ZN(new_n1062_));
  NOR3_X1    g1011(.A1(new_n570_), .A2(new_n564_), .A3(new_n1060_), .ZN(new_n1063_));
  NOR2_X1    g1012(.A1(new_n1062_), .A2(new_n1063_), .ZN(new_n1064_));
  NAND4_X1   g1013(.A1(new_n262_), .A2(new_n167_), .A3(new_n189_), .A4(new_n255_), .ZN(new_n1065_));
  NOR3_X1    g1014(.A1(new_n91_), .A2(new_n102_), .A3(new_n109_), .ZN(new_n1066_));
  NAND3_X1   g1015(.A1(new_n456_), .A2(new_n146_), .A3(new_n1066_), .ZN(new_n1067_));
  NOR4_X1    g1016(.A1(new_n1067_), .A2(new_n1065_), .A3(new_n468_), .A4(new_n261_), .ZN(new_n1068_));
  NAND4_X1   g1017(.A1(new_n166_), .A2(new_n315_), .A3(new_n146_), .A4(new_n149_), .ZN(new_n1069_));
  NOR2_X1    g1018(.A1(new_n239_), .A2(new_n91_), .ZN(new_n1070_));
  NAND4_X1   g1019(.A1(new_n1070_), .A2(new_n146_), .A3(new_n150_), .A4(new_n316_), .ZN(new_n1071_));
  NOR4_X1    g1020(.A1(new_n1069_), .A2(new_n1071_), .A3(new_n205_), .A4(new_n110_), .ZN(new_n1072_));
  NAND2_X1   g1021(.A1(new_n345_), .A2(new_n485_), .ZN(new_n1073_));
  NOR4_X1    g1022(.A1(new_n1073_), .A2(new_n156_), .A3(new_n205_), .A4(new_n332_), .ZN(new_n1074_));
  NAND3_X1   g1023(.A1(new_n1068_), .A2(new_n1074_), .A3(new_n1072_), .ZN(new_n1075_));
  NOR3_X1    g1024(.A1(new_n110_), .A2(new_n331_), .A3(new_n374_), .ZN(new_n1076_));
  NOR3_X1    g1025(.A1(new_n460_), .A2(new_n156_), .A3(new_n401_), .ZN(new_n1077_));
  NOR3_X1    g1026(.A1(new_n313_), .A2(new_n649_), .A3(new_n311_), .ZN(new_n1078_));
  NAND3_X1   g1027(.A1(new_n315_), .A2(new_n167_), .A3(new_n244_), .ZN(new_n1079_));
  NAND4_X1   g1028(.A1(new_n186_), .A2(new_n121_), .A3(new_n239_), .A4(new_n352_), .ZN(new_n1080_));
  NOR4_X1    g1029(.A1(new_n1080_), .A2(new_n1079_), .A3(new_n347_), .A4(new_n602_), .ZN(new_n1081_));
  NAND4_X1   g1030(.A1(new_n1081_), .A2(new_n1077_), .A3(new_n1076_), .A4(new_n1078_), .ZN(new_n1082_));
  NOR4_X1    g1031(.A1(new_n388_), .A2(new_n367_), .A3(new_n420_), .A4(new_n398_), .ZN(new_n1083_));
  NAND3_X1   g1032(.A1(new_n340_), .A2(new_n315_), .A3(new_n202_), .ZN(new_n1084_));
  NOR3_X1    g1033(.A1(new_n1084_), .A2(new_n449_), .A3(new_n413_), .ZN(new_n1085_));
  NOR4_X1    g1034(.A1(new_n201_), .A2(new_n366_), .A3(new_n339_), .A4(new_n395_), .ZN(new_n1086_));
  NAND3_X1   g1035(.A1(new_n149_), .A2(new_n337_), .A3(new_n131_), .ZN(new_n1087_));
  AOI21_X1   g1036(.A1(new_n478_), .A2(new_n1087_), .B(new_n78_), .ZN(new_n1088_));
  NAND3_X1   g1037(.A1(new_n454_), .A2(new_n776_), .A3(new_n146_), .ZN(new_n1089_));
  NOR4_X1    g1038(.A1(new_n1088_), .A2(new_n449_), .A3(new_n1089_), .A4(new_n207_), .ZN(new_n1090_));
  NAND4_X1   g1039(.A1(new_n1090_), .A2(new_n1083_), .A3(new_n1085_), .A4(new_n1086_), .ZN(new_n1091_));
  NOR3_X1    g1040(.A1(new_n1091_), .A2(new_n1075_), .A3(new_n1082_), .ZN(new_n1092_));
  NAND3_X1   g1041(.A1(new_n1092_), .A2(new_n437_), .A3(new_n875_), .ZN(new_n1093_));
  NOR2_X1    g1042(.A1(new_n256_), .A2(new_n221_), .ZN(new_n1094_));
  NOR2_X1    g1043(.A1(new_n821_), .A2(new_n151_), .ZN(new_n1095_));
  NAND4_X1   g1044(.A1(new_n1095_), .A2(new_n1094_), .A3(new_n222_), .A4(new_n622_), .ZN(new_n1096_));
  NAND2_X1   g1045(.A1(new_n474_), .A2(new_n679_), .ZN(new_n1097_));
  NOR2_X1    g1046(.A1(new_n196_), .A2(new_n383_), .ZN(new_n1098_));
  NAND4_X1   g1047(.A1(new_n1098_), .A2(new_n372_), .A3(new_n160_), .A4(new_n404_), .ZN(new_n1099_));
  NOR3_X1    g1048(.A1(new_n1096_), .A2(new_n1097_), .A3(new_n1099_), .ZN(new_n1100_));
  NOR3_X1    g1049(.A1(new_n412_), .A2(new_n91_), .A3(new_n239_), .ZN(new_n1101_));
  NAND3_X1   g1050(.A1(new_n207_), .A2(new_n452_), .A3(new_n1101_), .ZN(new_n1102_));
  NOR3_X1    g1051(.A1(new_n260_), .A2(new_n173_), .A3(new_n239_), .ZN(new_n1103_));
  NOR3_X1    g1052(.A1(new_n515_), .A2(new_n728_), .A3(new_n322_), .ZN(new_n1104_));
  NAND4_X1   g1053(.A1(new_n1104_), .A2(new_n417_), .A3(new_n1103_), .A4(new_n399_), .ZN(new_n1105_));
  NOR4_X1    g1054(.A1(new_n1105_), .A2(new_n152_), .A3(new_n1102_), .A4(new_n175_), .ZN(new_n1106_));
  NOR3_X1    g1055(.A1(new_n413_), .A2(new_n171_), .A3(new_n306_), .ZN(new_n1107_));
  NOR2_X1    g1056(.A1(new_n537_), .A2(new_n285_), .ZN(new_n1108_));
  NAND3_X1   g1057(.A1(new_n1083_), .A2(new_n1107_), .A3(new_n1108_), .ZN(new_n1109_));
  NOR4_X1    g1058(.A1(new_n243_), .A2(new_n245_), .A3(new_n306_), .A4(new_n211_), .ZN(new_n1110_));
  NOR4_X1    g1059(.A1(new_n230_), .A2(new_n319_), .A3(new_n171_), .A4(new_n306_), .ZN(new_n1111_));
  NAND3_X1   g1060(.A1(new_n1086_), .A2(new_n1111_), .A3(new_n1110_), .ZN(new_n1112_));
  NOR2_X1    g1061(.A1(new_n1112_), .A2(new_n1109_), .ZN(new_n1113_));
  NAND3_X1   g1062(.A1(new_n1100_), .A2(new_n1113_), .A3(new_n1106_), .ZN(new_n1114_));
  OAI21_X1   g1063(.A1(new_n1114_), .A2(new_n645_), .B(new_n438_), .ZN(new_n1115_));
  AOI21_X1   g1064(.A1(new_n1115_), .A2(new_n1093_), .B(new_n645_), .ZN(new_n1116_));
  INV_X1     g1065(.I(new_n1116_), .ZN(new_n1117_));
  INV_X1     g1066(.I(\a[1] ), .ZN(new_n1118_));
  NOR2_X1    g1067(.A1(\a[0] ), .A2(\a[2] ), .ZN(new_n1119_));
  AOI21_X1   g1068(.A1(new_n1119_), .A2(new_n62_), .B(new_n1118_), .ZN(new_n1120_));
  XOR2_X1    g1069(.A1(new_n1120_), .A2(\a[3] ), .Z(new_n1121_));
  INV_X1     g1070(.I(new_n1121_), .ZN(new_n1122_));
  AOI21_X1   g1071(.A1(new_n266_), .A2(new_n1122_), .B(new_n552_), .ZN(new_n1123_));
  NOR2_X1    g1072(.A1(new_n266_), .A2(new_n1122_), .ZN(new_n1124_));
  NOR3_X1    g1073(.A1(new_n1123_), .A2(new_n1124_), .A3(new_n559_), .ZN(new_n1125_));
  INV_X1     g1074(.I(new_n1125_), .ZN(new_n1126_));
  NOR2_X1    g1075(.A1(new_n1126_), .A2(new_n1117_), .ZN(new_n1127_));
  INV_X1     g1076(.I(new_n1127_), .ZN(new_n1128_));
  NOR3_X1    g1077(.A1(new_n1128_), .A2(new_n1055_), .A3(new_n1064_), .ZN(new_n1129_));
  INV_X1     g1078(.I(new_n1129_), .ZN(new_n1130_));
  NOR2_X1    g1079(.A1(new_n687_), .A2(new_n559_), .ZN(new_n1131_));
  NOR3_X1    g1080(.A1(new_n550_), .A2(new_n686_), .A3(new_n682_), .ZN(new_n1132_));
  NOR2_X1    g1081(.A1(new_n1131_), .A2(new_n1132_), .ZN(new_n1133_));
  AOI21_X1   g1082(.A1(new_n683_), .A2(new_n663_), .B(new_n1050_), .ZN(new_n1134_));
  NOR3_X1    g1083(.A1(new_n686_), .A2(new_n682_), .A3(new_n1051_), .ZN(new_n1135_));
  NOR2_X1    g1084(.A1(new_n364_), .A2(new_n619_), .ZN(new_n1136_));
  NOR2_X1    g1085(.A1(new_n310_), .A2(new_n407_), .ZN(new_n1137_));
  NAND3_X1   g1086(.A1(new_n1136_), .A2(new_n1137_), .A3(new_n174_), .ZN(new_n1138_));
  INV_X1     g1087(.I(new_n464_), .ZN(new_n1139_));
  NAND4_X1   g1088(.A1(new_n654_), .A2(new_n214_), .A3(new_n602_), .A4(new_n465_), .ZN(new_n1140_));
  INV_X1     g1089(.I(new_n469_), .ZN(new_n1141_));
  NOR4_X1    g1090(.A1(new_n1138_), .A2(new_n1139_), .A3(new_n1140_), .A4(new_n1141_), .ZN(new_n1142_));
  NOR2_X1    g1091(.A1(new_n585_), .A2(new_n471_), .ZN(new_n1143_));
  NAND4_X1   g1092(.A1(new_n1143_), .A2(new_n1142_), .A3(new_n484_), .A4(new_n487_), .ZN(new_n1144_));
  NOR3_X1    g1093(.A1(new_n1144_), .A2(new_n459_), .A3(new_n1051_), .ZN(new_n1145_));
  NOR2_X1    g1094(.A1(new_n489_), .A2(new_n1050_), .ZN(new_n1146_));
  NOR4_X1    g1095(.A1(new_n1134_), .A2(new_n1135_), .A3(new_n1146_), .A4(new_n1145_), .ZN(new_n1147_));
  OAI21_X1   g1096(.A1(\a[6] ), .A2(\a[22] ), .B(\a[5] ), .ZN(new_n1148_));
  XOR2_X1    g1097(.A1(new_n1045_), .A2(new_n1148_), .Z(new_n1149_));
  NOR4_X1    g1098(.A1(new_n693_), .A2(new_n1133_), .A3(new_n1147_), .A4(new_n1149_), .ZN(new_n1150_));
  INV_X1     g1099(.I(new_n1149_), .ZN(new_n1151_));
  NOR4_X1    g1100(.A1(new_n710_), .A2(new_n1133_), .A3(new_n1147_), .A4(new_n1151_), .ZN(new_n1152_));
  OAI21_X1   g1101(.A1(new_n1150_), .A2(new_n1152_), .B(new_n692_), .ZN(new_n1153_));
  MUX2_X1    g1102(.I0(new_n869_), .I1(new_n1019_), .S(new_n577_), .Z(new_n1154_));
  NOR3_X1    g1103(.A1(new_n1154_), .A2(new_n270_), .A3(new_n1018_), .ZN(new_n1155_));
  NOR3_X1    g1104(.A1(new_n1154_), .A2(new_n271_), .A3(new_n1017_), .ZN(new_n1156_));
  OAI21_X1   g1105(.A1(new_n1155_), .A2(new_n1156_), .B(new_n1016_), .ZN(new_n1157_));
  OAI21_X1   g1106(.A1(new_n1054_), .A2(new_n1052_), .B(new_n1116_), .ZN(new_n1158_));
  NAND2_X1   g1107(.A1(new_n567_), .A2(new_n1060_), .ZN(new_n1159_));
  NAND2_X1   g1108(.A1(new_n563_), .A2(new_n266_), .ZN(new_n1160_));
  NAND3_X1   g1109(.A1(new_n1160_), .A2(new_n579_), .A3(new_n1061_), .ZN(new_n1161_));
  AOI21_X1   g1110(.A1(new_n1159_), .A2(new_n1161_), .B(new_n1126_), .ZN(new_n1162_));
  NAND2_X1   g1111(.A1(new_n1158_), .A2(new_n1162_), .ZN(new_n1163_));
  NAND2_X1   g1112(.A1(new_n580_), .A2(new_n1050_), .ZN(new_n1164_));
  NAND2_X1   g1113(.A1(new_n561_), .A2(new_n1051_), .ZN(new_n1165_));
  AOI21_X1   g1114(.A1(new_n1165_), .A2(new_n1164_), .B(new_n1117_), .ZN(new_n1166_));
  OAI21_X1   g1115(.A1(new_n1062_), .A2(new_n1063_), .B(new_n1125_), .ZN(new_n1167_));
  NAND2_X1   g1116(.A1(new_n1166_), .A2(new_n1167_), .ZN(new_n1168_));
  AND2_X2    g1117(.A1(new_n1163_), .A2(new_n1168_), .Z(new_n1169_));
  OAI21_X1   g1118(.A1(new_n1169_), .A2(new_n1157_), .B(new_n1153_), .ZN(new_n1170_));
  NOR4_X1    g1119(.A1(new_n642_), .A2(new_n587_), .A3(new_n616_), .A4(new_n803_), .ZN(new_n1171_));
  INV_X1     g1120(.I(new_n1171_), .ZN(new_n1172_));
  AOI21_X1   g1121(.A1(new_n1169_), .A2(new_n1157_), .B(new_n1172_), .ZN(new_n1173_));
  AND2_X2    g1122(.A1(new_n1173_), .A2(new_n1170_), .Z(new_n1174_));
  NOR4_X1    g1123(.A1(new_n690_), .A2(new_n559_), .A3(new_n694_), .A4(new_n803_), .ZN(new_n1175_));
  INV_X1     g1124(.I(new_n1175_), .ZN(new_n1176_));
  NAND2_X1   g1125(.A1(new_n641_), .A2(new_n615_), .ZN(new_n1177_));
  NAND2_X1   g1126(.A1(new_n615_), .A2(new_n587_), .ZN(new_n1178_));
  INV_X1     g1127(.I(new_n1178_), .ZN(new_n1179_));
  NOR2_X1    g1128(.A1(new_n1179_), .A2(new_n1177_), .ZN(new_n1180_));
  NOR3_X1    g1129(.A1(new_n642_), .A2(new_n489_), .A3(new_n616_), .ZN(new_n1181_));
  INV_X1     g1130(.I(new_n1181_), .ZN(new_n1182_));
  AOI21_X1   g1131(.A1(new_n616_), .A2(new_n587_), .B(new_n642_), .ZN(new_n1183_));
  OAI21_X1   g1132(.A1(new_n641_), .A2(new_n587_), .B(new_n615_), .ZN(new_n1184_));
  NOR2_X1    g1133(.A1(new_n1184_), .A2(new_n270_), .ZN(new_n1185_));
  AOI21_X1   g1134(.A1(new_n270_), .A2(new_n1183_), .B(new_n1185_), .ZN(new_n1186_));
  NOR3_X1    g1135(.A1(new_n1186_), .A2(new_n576_), .A3(new_n1182_), .ZN(new_n1187_));
  NOR3_X1    g1136(.A1(new_n1186_), .A2(new_n577_), .A3(new_n1181_), .ZN(new_n1188_));
  OAI21_X1   g1137(.A1(new_n1187_), .A2(new_n1188_), .B(new_n1180_), .ZN(new_n1189_));
  NOR2_X1    g1138(.A1(new_n784_), .A2(new_n774_), .ZN(new_n1190_));
  INV_X1     g1139(.I(new_n830_), .ZN(new_n1191_));
  NAND2_X1   g1140(.A1(new_n526_), .A2(new_n795_), .ZN(new_n1192_));
  NOR4_X1    g1141(.A1(new_n1192_), .A2(new_n486_), .A3(new_n1008_), .A4(new_n1007_), .ZN(new_n1193_));
  NAND4_X1   g1142(.A1(new_n1191_), .A2(new_n1193_), .A3(new_n1190_), .A4(new_n999_), .ZN(new_n1194_));
  NOR3_X1    g1143(.A1(new_n867_), .A2(new_n1194_), .A3(new_n994_), .ZN(new_n1195_));
  NOR2_X1    g1144(.A1(new_n1014_), .A2(new_n758_), .ZN(new_n1196_));
  OAI21_X1   g1145(.A1(new_n1196_), .A2(new_n1195_), .B(new_n614_), .ZN(new_n1197_));
  NOR2_X1    g1146(.A1(new_n1019_), .A2(new_n708_), .ZN(new_n1198_));
  AOI21_X1   g1147(.A1(new_n708_), .A2(new_n1197_), .B(new_n1198_), .ZN(new_n1199_));
  NOR3_X1    g1148(.A1(new_n1199_), .A2(new_n721_), .A3(new_n1018_), .ZN(new_n1200_));
  NOR3_X1    g1149(.A1(new_n1199_), .A2(new_n702_), .A3(new_n1017_), .ZN(new_n1201_));
  OAI21_X1   g1150(.A1(new_n1200_), .A2(new_n1201_), .B(new_n1016_), .ZN(new_n1202_));
  INV_X1     g1151(.I(new_n1202_), .ZN(new_n1203_));
  NAND2_X1   g1152(.A1(new_n1189_), .A2(new_n1203_), .ZN(new_n1204_));
  INV_X1     g1153(.I(new_n1189_), .ZN(new_n1205_));
  NAND2_X1   g1154(.A1(new_n1205_), .A2(new_n1202_), .ZN(new_n1206_));
  AOI21_X1   g1155(.A1(new_n1206_), .A2(new_n1204_), .B(new_n1176_), .ZN(new_n1207_));
  NOR2_X1    g1156(.A1(new_n1189_), .A2(new_n1202_), .ZN(new_n1208_));
  INV_X1     g1157(.I(new_n1208_), .ZN(new_n1209_));
  NAND2_X1   g1158(.A1(new_n1189_), .A2(new_n1202_), .ZN(new_n1210_));
  AOI21_X1   g1159(.A1(new_n1209_), .A2(new_n1210_), .B(new_n1175_), .ZN(new_n1211_));
  NOR2_X1    g1160(.A1(new_n1211_), .A2(new_n1207_), .ZN(new_n1212_));
  XOR2_X1    g1161(.A1(new_n266_), .A2(new_n1060_), .Z(new_n1213_));
  NOR3_X1    g1162(.A1(new_n1212_), .A2(new_n1174_), .A3(new_n1213_), .ZN(new_n1214_));
  INV_X1     g1163(.I(new_n1174_), .ZN(new_n1215_));
  OR2_X2     g1164(.A1(new_n1211_), .A2(new_n1207_), .Z(new_n1216_));
  INV_X1     g1165(.I(new_n1213_), .ZN(new_n1217_));
  AOI21_X1   g1166(.A1(new_n1216_), .A2(new_n1217_), .B(new_n1215_), .ZN(new_n1218_));
  OAI21_X1   g1167(.A1(new_n1218_), .A2(new_n1214_), .B(new_n1130_), .ZN(new_n1219_));
  NAND3_X1   g1168(.A1(new_n1216_), .A2(new_n1215_), .A3(new_n1217_), .ZN(new_n1220_));
  OAI21_X1   g1169(.A1(new_n1212_), .A2(new_n1213_), .B(new_n1174_), .ZN(new_n1221_));
  NAND3_X1   g1170(.A1(new_n1220_), .A2(new_n1129_), .A3(new_n1221_), .ZN(new_n1222_));
  NOR2_X1    g1171(.A1(new_n925_), .A2(new_n1014_), .ZN(new_n1223_));
  NOR2_X1    g1172(.A1(new_n281_), .A2(new_n243_), .ZN(new_n1224_));
  NAND3_X1   g1173(.A1(new_n1224_), .A2(new_n319_), .A3(new_n891_), .ZN(new_n1225_));
  NOR2_X1    g1174(.A1(new_n156_), .A2(new_n230_), .ZN(new_n1226_));
  NAND3_X1   g1175(.A1(new_n1226_), .A2(new_n223_), .A3(new_n746_), .ZN(new_n1227_));
  OAI21_X1   g1176(.A1(new_n991_), .A2(new_n1066_), .B(new_n146_), .ZN(new_n1228_));
  NOR3_X1    g1177(.A1(new_n306_), .A2(new_n1010_), .A3(new_n169_), .ZN(new_n1229_));
  OAI21_X1   g1178(.A1(new_n201_), .A2(new_n171_), .B(new_n547_), .ZN(new_n1230_));
  NAND4_X1   g1179(.A1(new_n1230_), .A2(new_n512_), .A3(new_n1228_), .A4(new_n1229_), .ZN(new_n1231_));
  NOR3_X1    g1180(.A1(new_n207_), .A2(new_n285_), .A3(new_n399_), .ZN(new_n1232_));
  NAND2_X1   g1181(.A1(new_n1232_), .A2(new_n856_), .ZN(new_n1233_));
  NOR4_X1    g1182(.A1(new_n1231_), .A2(new_n1233_), .A3(new_n1227_), .A4(new_n1225_), .ZN(new_n1234_));
  NAND2_X1   g1183(.A1(new_n207_), .A2(new_n399_), .ZN(new_n1235_));
  NOR4_X1    g1184(.A1(new_n635_), .A2(new_n485_), .A3(new_n201_), .A4(new_n733_), .ZN(new_n1236_));
  NAND3_X1   g1185(.A1(new_n1236_), .A2(new_n365_), .A3(new_n1235_), .ZN(new_n1237_));
  NOR2_X1    g1186(.A1(new_n338_), .A2(new_n221_), .ZN(new_n1238_));
  NAND4_X1   g1187(.A1(new_n789_), .A2(new_n678_), .A3(new_n383_), .A4(new_n1238_), .ZN(new_n1239_));
  NOR2_X1    g1188(.A1(new_n232_), .A2(new_n454_), .ZN(new_n1240_));
  NOR2_X1    g1189(.A1(new_n668_), .A2(new_n251_), .ZN(new_n1241_));
  NAND4_X1   g1190(.A1(new_n1240_), .A2(new_n1241_), .A3(new_n205_), .A4(new_n307_), .ZN(new_n1242_));
  NOR4_X1    g1191(.A1(new_n1237_), .A2(new_n1239_), .A3(new_n911_), .A4(new_n1242_), .ZN(new_n1243_));
  INV_X1     g1192(.I(new_n919_), .ZN(new_n1244_));
  NAND2_X1   g1193(.A1(new_n150_), .A2(new_n352_), .ZN(new_n1245_));
  AOI21_X1   g1194(.A1(new_n1245_), .A2(new_n260_), .B(new_n121_), .ZN(new_n1246_));
  NAND4_X1   g1195(.A1(new_n600_), .A2(new_n305_), .A3(new_n1246_), .A4(new_n654_), .ZN(new_n1247_));
  NOR2_X1    g1196(.A1(new_n168_), .A2(new_n132_), .ZN(new_n1248_));
  NAND2_X1   g1197(.A1(new_n1248_), .A2(new_n420_), .ZN(new_n1249_));
  NOR4_X1    g1198(.A1(new_n1247_), .A2(new_n1244_), .A3(new_n1249_), .A4(new_n922_), .ZN(new_n1250_));
  NAND3_X1   g1199(.A1(new_n1243_), .A2(new_n1234_), .A3(new_n1250_), .ZN(new_n1251_));
  NOR2_X1    g1200(.A1(new_n1251_), .A2(new_n1014_), .ZN(new_n1252_));
  NAND2_X1   g1201(.A1(new_n925_), .A2(new_n1014_), .ZN(new_n1253_));
  NAND2_X1   g1202(.A1(new_n1253_), .A2(new_n875_), .ZN(new_n1254_));
  OAI21_X1   g1203(.A1(new_n875_), .A2(new_n1252_), .B(new_n1254_), .ZN(new_n1255_));
  NAND3_X1   g1204(.A1(new_n1255_), .A2(new_n711_), .A3(new_n1223_), .ZN(new_n1256_));
  INV_X1     g1205(.I(new_n1223_), .ZN(new_n1257_));
  NAND3_X1   g1206(.A1(new_n1255_), .A2(new_n708_), .A3(new_n1257_), .ZN(new_n1258_));
  AOI21_X1   g1207(.A1(new_n1256_), .A2(new_n1258_), .B(new_n925_), .ZN(new_n1259_));
  NOR2_X1    g1208(.A1(new_n1114_), .A2(new_n438_), .ZN(new_n1260_));
  INV_X1     g1209(.I(new_n1260_), .ZN(new_n1261_));
  NAND3_X1   g1210(.A1(new_n1259_), .A2(new_n566_), .A3(new_n1261_), .ZN(new_n1262_));
  AOI21_X1   g1211(.A1(new_n1259_), .A2(new_n1261_), .B(new_n566_), .ZN(new_n1263_));
  INV_X1     g1212(.I(new_n1263_), .ZN(new_n1264_));
  AOI21_X1   g1213(.A1(new_n1264_), .A2(new_n1262_), .B(new_n1122_), .ZN(new_n1265_));
  INV_X1     g1214(.I(new_n1262_), .ZN(new_n1266_));
  NOR3_X1    g1215(.A1(new_n1266_), .A2(new_n1121_), .A3(new_n1263_), .ZN(new_n1267_));
  NOR2_X1    g1216(.A1(new_n1265_), .A2(new_n1267_), .ZN(new_n1268_));
  NOR4_X1    g1217(.A1(new_n642_), .A2(new_n271_), .A3(new_n587_), .A4(new_n616_), .ZN(new_n1269_));
  NOR4_X1    g1218(.A1(new_n687_), .A2(new_n559_), .A3(new_n587_), .A4(new_n809_), .ZN(new_n1270_));
  INV_X1     g1219(.I(new_n1270_), .ZN(new_n1271_));
  MUX2_X1    g1220(.I0(new_n869_), .I1(new_n1019_), .S(new_n702_), .Z(new_n1272_));
  NOR3_X1    g1221(.A1(new_n1272_), .A2(new_n576_), .A3(new_n1018_), .ZN(new_n1273_));
  NOR3_X1    g1222(.A1(new_n1272_), .A2(new_n577_), .A3(new_n1017_), .ZN(new_n1274_));
  OAI21_X1   g1223(.A1(new_n1273_), .A2(new_n1274_), .B(new_n1016_), .ZN(new_n1275_));
  XOR2_X1    g1224(.A1(new_n1275_), .A2(new_n1271_), .Z(new_n1276_));
  NAND2_X1   g1225(.A1(new_n1276_), .A2(new_n1269_), .ZN(new_n1277_));
  INV_X1     g1226(.I(new_n1269_), .ZN(new_n1278_));
  NOR2_X1    g1227(.A1(new_n1275_), .A2(new_n1271_), .ZN(new_n1279_));
  NAND2_X1   g1228(.A1(new_n1275_), .A2(new_n1271_), .ZN(new_n1280_));
  INV_X1     g1229(.I(new_n1280_), .ZN(new_n1281_));
  OAI21_X1   g1230(.A1(new_n1281_), .A2(new_n1279_), .B(new_n1278_), .ZN(new_n1282_));
  NAND2_X1   g1231(.A1(new_n1277_), .A2(new_n1282_), .ZN(new_n1283_));
  NAND2_X1   g1232(.A1(new_n1283_), .A2(new_n1268_), .ZN(new_n1284_));
  XOR2_X1    g1233(.A1(new_n1125_), .A2(new_n1117_), .Z(new_n1285_));
  NAND2_X1   g1234(.A1(new_n1253_), .A2(new_n711_), .ZN(new_n1286_));
  OAI21_X1   g1235(.A1(new_n711_), .A2(new_n1252_), .B(new_n1286_), .ZN(new_n1287_));
  NAND3_X1   g1236(.A1(new_n1287_), .A2(new_n702_), .A3(new_n1223_), .ZN(new_n1288_));
  NAND3_X1   g1237(.A1(new_n1287_), .A2(new_n721_), .A3(new_n1257_), .ZN(new_n1289_));
  NAND2_X1   g1238(.A1(new_n1288_), .A2(new_n1289_), .ZN(new_n1290_));
  NAND2_X1   g1239(.A1(new_n1290_), .A2(new_n1251_), .ZN(new_n1291_));
  NAND2_X1   g1240(.A1(new_n1291_), .A2(new_n1285_), .ZN(new_n1292_));
  INV_X1     g1241(.I(new_n1292_), .ZN(new_n1293_));
  NAND2_X1   g1242(.A1(new_n567_), .A2(new_n1121_), .ZN(new_n1294_));
  OAI21_X1   g1243(.A1(new_n572_), .A2(new_n1121_), .B(new_n1294_), .ZN(new_n1295_));
  NAND3_X1   g1244(.A1(new_n1295_), .A2(new_n565_), .A3(new_n1061_), .ZN(new_n1296_));
  NAND3_X1   g1245(.A1(new_n1295_), .A2(new_n580_), .A3(new_n1060_), .ZN(new_n1297_));
  AOI21_X1   g1246(.A1(new_n1296_), .A2(new_n1297_), .B(new_n561_), .ZN(new_n1298_));
  INV_X1     g1247(.I(new_n1298_), .ZN(new_n1299_));
  NOR2_X1    g1248(.A1(new_n1291_), .A2(new_n1285_), .ZN(new_n1300_));
  INV_X1     g1249(.I(new_n1300_), .ZN(new_n1301_));
  AOI21_X1   g1250(.A1(new_n1299_), .A2(new_n1301_), .B(new_n1293_), .ZN(new_n1302_));
  INV_X1     g1251(.I(new_n1302_), .ZN(new_n1303_));
  OAI21_X1   g1252(.A1(new_n1266_), .A2(new_n1263_), .B(new_n1121_), .ZN(new_n1304_));
  NAND3_X1   g1253(.A1(new_n1264_), .A2(new_n1122_), .A3(new_n1262_), .ZN(new_n1305_));
  NAND2_X1   g1254(.A1(new_n1305_), .A2(new_n1304_), .ZN(new_n1306_));
  NAND3_X1   g1255(.A1(new_n1306_), .A2(new_n1277_), .A3(new_n1282_), .ZN(new_n1307_));
  NAND2_X1   g1256(.A1(new_n1307_), .A2(new_n1303_), .ZN(new_n1308_));
  NAND2_X1   g1257(.A1(new_n1308_), .A2(new_n1284_), .ZN(new_n1309_));
  OAI21_X1   g1258(.A1(new_n1269_), .A2(new_n1279_), .B(new_n1280_), .ZN(new_n1310_));
  INV_X1     g1259(.I(new_n1310_), .ZN(new_n1311_));
  NAND2_X1   g1260(.A1(new_n567_), .A2(new_n1050_), .ZN(new_n1312_));
  OAI21_X1   g1261(.A1(new_n572_), .A2(new_n1050_), .B(new_n1312_), .ZN(new_n1313_));
  NAND3_X1   g1262(.A1(new_n1313_), .A2(new_n565_), .A3(new_n1151_), .ZN(new_n1314_));
  NAND3_X1   g1263(.A1(new_n1313_), .A2(new_n580_), .A3(new_n1149_), .ZN(new_n1315_));
  AOI21_X1   g1264(.A1(new_n1314_), .A2(new_n1315_), .B(new_n561_), .ZN(new_n1316_));
  NAND2_X1   g1265(.A1(new_n1259_), .A2(new_n266_), .ZN(new_n1317_));
  NOR2_X1    g1266(.A1(new_n1260_), .A2(new_n1121_), .ZN(new_n1318_));
  OAI21_X1   g1267(.A1(new_n1259_), .A2(new_n266_), .B(new_n1318_), .ZN(new_n1319_));
  NAND2_X1   g1268(.A1(new_n1319_), .A2(new_n1317_), .ZN(new_n1320_));
  NAND2_X1   g1269(.A1(new_n1316_), .A2(new_n1320_), .ZN(new_n1321_));
  INV_X1     g1270(.I(new_n1316_), .ZN(new_n1322_));
  INV_X1     g1271(.I(new_n1320_), .ZN(new_n1323_));
  NAND2_X1   g1272(.A1(new_n1322_), .A2(new_n1323_), .ZN(new_n1324_));
  AOI21_X1   g1273(.A1(new_n1324_), .A2(new_n1321_), .B(new_n1311_), .ZN(new_n1325_));
  NAND2_X1   g1274(.A1(new_n1322_), .A2(new_n1320_), .ZN(new_n1326_));
  NAND2_X1   g1275(.A1(new_n1323_), .A2(new_n1316_), .ZN(new_n1327_));
  AOI21_X1   g1276(.A1(new_n1326_), .A2(new_n1327_), .B(new_n1310_), .ZN(new_n1328_));
  NOR2_X1    g1277(.A1(new_n1325_), .A2(new_n1328_), .ZN(new_n1329_));
  NOR2_X1    g1278(.A1(new_n1309_), .A2(new_n1329_), .ZN(new_n1330_));
  INV_X1     g1279(.I(new_n1330_), .ZN(new_n1331_));
  NAND2_X1   g1280(.A1(new_n1309_), .A2(new_n1329_), .ZN(new_n1332_));
  AOI22_X1   g1281(.A1(new_n1332_), .A2(new_n1331_), .B1(new_n1219_), .B2(new_n1222_), .ZN(new_n1333_));
  NAND2_X1   g1282(.A1(new_n1219_), .A2(new_n1222_), .ZN(new_n1334_));
  XNOR2_X1   g1283(.A1(new_n1309_), .A2(new_n1329_), .ZN(new_n1335_));
  NOR2_X1    g1284(.A1(new_n1334_), .A2(new_n1335_), .ZN(new_n1336_));
  NOR2_X1    g1285(.A1(new_n1336_), .A2(new_n1333_), .ZN(new_n1337_));
  INV_X1     g1286(.I(new_n1337_), .ZN(new_n1338_));
  INV_X1     g1287(.I(new_n1016_), .ZN(new_n1339_));
  OAI21_X1   g1288(.A1(new_n1196_), .A2(new_n1195_), .B(new_n428_), .ZN(new_n1340_));
  MUX2_X1    g1289(.I0(new_n1340_), .I1(new_n1197_), .S(new_n808_), .Z(new_n1341_));
  NAND3_X1   g1290(.A1(new_n1341_), .A2(new_n1017_), .A3(new_n1151_), .ZN(new_n1342_));
  NAND3_X1   g1291(.A1(new_n1341_), .A2(new_n1018_), .A3(new_n1149_), .ZN(new_n1343_));
  AOI21_X1   g1292(.A1(new_n1342_), .A2(new_n1343_), .B(new_n1339_), .ZN(new_n1344_));
  NOR2_X1    g1293(.A1(new_n1251_), .A2(new_n798_), .ZN(new_n1345_));
  MUX2_X1    g1294(.I0(new_n1252_), .I1(new_n1345_), .S(new_n271_), .Z(new_n1346_));
  NOR3_X1    g1295(.A1(new_n1346_), .A2(new_n802_), .A3(new_n1257_), .ZN(new_n1347_));
  NOR3_X1    g1296(.A1(new_n1346_), .A2(new_n803_), .A3(new_n1223_), .ZN(new_n1348_));
  OAI21_X1   g1297(.A1(new_n1347_), .A2(new_n1348_), .B(new_n1251_), .ZN(new_n1349_));
  NAND2_X1   g1298(.A1(new_n1092_), .A2(new_n577_), .ZN(new_n1350_));
  XOR2_X1    g1299(.A1(new_n1350_), .A2(new_n702_), .Z(new_n1351_));
  NOR2_X1    g1300(.A1(new_n1351_), .A2(new_n576_), .ZN(new_n1352_));
  INV_X1     g1301(.I(new_n1352_), .ZN(new_n1353_));
  NOR2_X1    g1302(.A1(new_n1349_), .A2(new_n1353_), .ZN(new_n1354_));
  NAND2_X1   g1303(.A1(new_n1253_), .A2(new_n271_), .ZN(new_n1355_));
  NAND2_X1   g1304(.A1(new_n926_), .A2(new_n270_), .ZN(new_n1356_));
  NAND2_X1   g1305(.A1(new_n1356_), .A2(new_n1355_), .ZN(new_n1357_));
  NAND3_X1   g1306(.A1(new_n1357_), .A2(new_n803_), .A3(new_n1223_), .ZN(new_n1358_));
  NAND3_X1   g1307(.A1(new_n1357_), .A2(new_n802_), .A3(new_n1257_), .ZN(new_n1359_));
  NAND2_X1   g1308(.A1(new_n1358_), .A2(new_n1359_), .ZN(new_n1360_));
  AOI21_X1   g1309(.A1(new_n1360_), .A2(new_n1251_), .B(new_n1352_), .ZN(new_n1361_));
  OAI21_X1   g1310(.A1(new_n1354_), .A2(new_n1361_), .B(new_n1344_), .ZN(new_n1362_));
  AOI21_X1   g1311(.A1(new_n1360_), .A2(new_n1251_), .B(new_n1353_), .ZN(new_n1363_));
  NOR2_X1    g1312(.A1(new_n1349_), .A2(new_n1352_), .ZN(new_n1364_));
  NOR2_X1    g1313(.A1(new_n1363_), .A2(new_n1364_), .ZN(new_n1365_));
  OAI21_X1   g1314(.A1(new_n1344_), .A2(new_n1365_), .B(new_n1362_), .ZN(new_n1366_));
  MUX2_X1    g1315(.I0(new_n1340_), .I1(new_n1197_), .S(new_n1149_), .Z(new_n1367_));
  NAND3_X1   g1316(.A1(new_n1367_), .A2(new_n1017_), .A3(new_n1051_), .ZN(new_n1368_));
  NAND3_X1   g1317(.A1(new_n1367_), .A2(new_n1018_), .A3(new_n1050_), .ZN(new_n1369_));
  AOI21_X1   g1318(.A1(new_n1368_), .A2(new_n1369_), .B(new_n1339_), .ZN(new_n1370_));
  NAND2_X1   g1319(.A1(new_n1253_), .A2(new_n803_), .ZN(new_n1371_));
  OAI21_X1   g1320(.A1(new_n803_), .A2(new_n1252_), .B(new_n1371_), .ZN(new_n1372_));
  NAND3_X1   g1321(.A1(new_n1372_), .A2(new_n809_), .A3(new_n1223_), .ZN(new_n1373_));
  NAND3_X1   g1322(.A1(new_n1372_), .A2(new_n808_), .A3(new_n1257_), .ZN(new_n1374_));
  AOI21_X1   g1323(.A1(new_n1373_), .A2(new_n1374_), .B(new_n925_), .ZN(new_n1375_));
  NOR2_X1    g1324(.A1(new_n1370_), .A2(new_n1375_), .ZN(new_n1376_));
  NOR4_X1    g1325(.A1(new_n587_), .A2(new_n640_), .A3(new_n614_), .A4(new_n1061_), .ZN(new_n1377_));
  INV_X1     g1326(.I(new_n1377_), .ZN(new_n1378_));
  NAND2_X1   g1327(.A1(new_n1370_), .A2(new_n1375_), .ZN(new_n1379_));
  AOI21_X1   g1328(.A1(new_n1378_), .A2(new_n1379_), .B(new_n1376_), .ZN(new_n1380_));
  NOR2_X1    g1329(.A1(new_n1366_), .A2(new_n1380_), .ZN(new_n1381_));
  NAND4_X1   g1330(.A1(new_n641_), .A2(new_n615_), .A3(new_n489_), .A4(new_n1050_), .ZN(new_n1382_));
  NOR3_X1    g1331(.A1(new_n1114_), .A2(new_n270_), .A3(new_n577_), .ZN(new_n1383_));
  AOI21_X1   g1332(.A1(new_n1092_), .A2(new_n271_), .B(new_n576_), .ZN(new_n1384_));
  OAI21_X1   g1333(.A1(new_n1383_), .A2(new_n1384_), .B(new_n271_), .ZN(new_n1385_));
  INV_X1     g1334(.I(new_n1385_), .ZN(new_n1386_));
  NAND2_X1   g1335(.A1(new_n371_), .A2(new_n1121_), .ZN(new_n1387_));
  NOR4_X1    g1336(.A1(new_n489_), .A2(new_n371_), .A3(new_n428_), .A4(new_n1121_), .ZN(new_n1388_));
  AOI21_X1   g1337(.A1(new_n586_), .A2(new_n584_), .B(new_n1121_), .ZN(new_n1389_));
  AOI21_X1   g1338(.A1(new_n1389_), .A2(new_n640_), .B(new_n614_), .ZN(new_n1390_));
  OAI21_X1   g1339(.A1(new_n1390_), .A2(new_n1388_), .B(new_n1387_), .ZN(new_n1391_));
  NOR2_X1    g1340(.A1(new_n1391_), .A2(new_n1178_), .ZN(new_n1392_));
  NAND2_X1   g1341(.A1(new_n1392_), .A2(new_n1386_), .ZN(new_n1393_));
  NOR3_X1    g1342(.A1(new_n1393_), .A2(new_n689_), .A3(new_n1382_), .ZN(new_n1394_));
  INV_X1     g1343(.I(new_n1394_), .ZN(new_n1395_));
  OAI21_X1   g1344(.A1(new_n1393_), .A2(new_n1382_), .B(new_n689_), .ZN(new_n1396_));
  AOI21_X1   g1345(.A1(new_n1395_), .A2(new_n1396_), .B(new_n1122_), .ZN(new_n1397_));
  INV_X1     g1346(.I(new_n1396_), .ZN(new_n1398_));
  NOR3_X1    g1347(.A1(new_n1398_), .A2(new_n1121_), .A3(new_n1394_), .ZN(new_n1399_));
  NOR2_X1    g1348(.A1(new_n1397_), .A2(new_n1399_), .ZN(new_n1400_));
  NAND2_X1   g1349(.A1(new_n1366_), .A2(new_n1380_), .ZN(new_n1401_));
  AOI21_X1   g1350(.A1(new_n1400_), .A2(new_n1401_), .B(new_n1381_), .ZN(new_n1402_));
  INV_X1     g1351(.I(new_n1402_), .ZN(new_n1403_));
  MUX2_X1    g1352(.I0(new_n1019_), .I1(new_n869_), .S(new_n1050_), .Z(new_n1404_));
  NOR3_X1    g1353(.A1(new_n1404_), .A2(new_n1018_), .A3(new_n1060_), .ZN(new_n1405_));
  NOR3_X1    g1354(.A1(new_n1404_), .A2(new_n1017_), .A3(new_n1061_), .ZN(new_n1406_));
  OAI21_X1   g1355(.A1(new_n1405_), .A2(new_n1406_), .B(new_n1016_), .ZN(new_n1407_));
  OAI21_X1   g1356(.A1(new_n1251_), .A2(new_n1014_), .B(new_n808_), .ZN(new_n1408_));
  OAI21_X1   g1357(.A1(new_n808_), .A2(new_n1345_), .B(new_n1408_), .ZN(new_n1409_));
  NAND3_X1   g1358(.A1(new_n1409_), .A2(new_n1151_), .A3(new_n1223_), .ZN(new_n1410_));
  NAND3_X1   g1359(.A1(new_n1409_), .A2(new_n1149_), .A3(new_n1257_), .ZN(new_n1411_));
  NAND2_X1   g1360(.A1(new_n1410_), .A2(new_n1411_), .ZN(new_n1412_));
  NAND2_X1   g1361(.A1(new_n1092_), .A2(new_n803_), .ZN(new_n1413_));
  XOR2_X1    g1362(.A1(new_n1413_), .A2(new_n270_), .Z(new_n1414_));
  NAND2_X1   g1363(.A1(new_n1414_), .A2(new_n803_), .ZN(new_n1415_));
  INV_X1     g1364(.I(new_n1415_), .ZN(new_n1416_));
  NAND3_X1   g1365(.A1(new_n1412_), .A2(new_n1416_), .A3(new_n1251_), .ZN(new_n1417_));
  AOI21_X1   g1366(.A1(new_n925_), .A2(new_n1014_), .B(new_n808_), .ZN(new_n1418_));
  AOI21_X1   g1367(.A1(new_n808_), .A2(new_n926_), .B(new_n1418_), .ZN(new_n1419_));
  NOR3_X1    g1368(.A1(new_n1419_), .A2(new_n1149_), .A3(new_n1257_), .ZN(new_n1420_));
  NOR3_X1    g1369(.A1(new_n1419_), .A2(new_n1151_), .A3(new_n1223_), .ZN(new_n1421_));
  OAI21_X1   g1370(.A1(new_n1420_), .A2(new_n1421_), .B(new_n1251_), .ZN(new_n1422_));
  NAND2_X1   g1371(.A1(new_n1422_), .A2(new_n1415_), .ZN(new_n1423_));
  AOI21_X1   g1372(.A1(new_n1417_), .A2(new_n1423_), .B(new_n1407_), .ZN(new_n1424_));
  MUX2_X1    g1373(.I0(new_n1197_), .I1(new_n1340_), .S(new_n1051_), .Z(new_n1425_));
  NAND3_X1   g1374(.A1(new_n1425_), .A2(new_n1017_), .A3(new_n1061_), .ZN(new_n1426_));
  NAND3_X1   g1375(.A1(new_n1425_), .A2(new_n1018_), .A3(new_n1060_), .ZN(new_n1427_));
  NAND2_X1   g1376(.A1(new_n1426_), .A2(new_n1427_), .ZN(new_n1428_));
  NAND2_X1   g1377(.A1(new_n1422_), .A2(new_n1416_), .ZN(new_n1429_));
  NAND3_X1   g1378(.A1(new_n1412_), .A2(new_n1251_), .A3(new_n1415_), .ZN(new_n1430_));
  AOI22_X1   g1379(.A1(new_n1428_), .A2(new_n1016_), .B1(new_n1429_), .B2(new_n1430_), .ZN(new_n1431_));
  NOR2_X1    g1380(.A1(new_n1424_), .A2(new_n1431_), .ZN(new_n1432_));
  NOR2_X1    g1381(.A1(new_n175_), .A2(new_n152_), .ZN(new_n1433_));
  NOR2_X1    g1382(.A1(new_n1105_), .A2(new_n1102_), .ZN(new_n1434_));
  NAND4_X1   g1383(.A1(new_n201_), .A2(new_n292_), .A3(new_n363_), .A4(new_n608_), .ZN(new_n1435_));
  NOR4_X1    g1384(.A1(new_n1435_), .A2(new_n413_), .A3(new_n449_), .A4(new_n1084_), .ZN(new_n1436_));
  NAND4_X1   g1385(.A1(new_n388_), .A2(new_n230_), .A3(new_n475_), .A4(new_n329_), .ZN(new_n1437_));
  NAND3_X1   g1386(.A1(new_n232_), .A2(new_n313_), .A3(new_n454_), .ZN(new_n1438_));
  NOR4_X1    g1387(.A1(new_n1437_), .A2(new_n1438_), .A3(new_n449_), .A4(new_n1088_), .ZN(new_n1439_));
  NAND4_X1   g1388(.A1(new_n1434_), .A2(new_n1439_), .A3(new_n1436_), .A4(new_n1433_), .ZN(new_n1440_));
  NOR4_X1    g1389(.A1(new_n1440_), .A2(new_n803_), .A3(new_n808_), .A4(new_n1075_), .ZN(new_n1441_));
  AOI21_X1   g1390(.A1(new_n1092_), .A2(new_n809_), .B(new_n802_), .ZN(new_n1442_));
  OAI21_X1   g1391(.A1(new_n1442_), .A2(new_n1441_), .B(new_n809_), .ZN(new_n1443_));
  AOI21_X1   g1392(.A1(new_n428_), .A2(new_n1122_), .B(new_n1014_), .ZN(new_n1444_));
  OAI21_X1   g1393(.A1(new_n428_), .A2(new_n1122_), .B(new_n867_), .ZN(new_n1445_));
  NOR2_X1    g1394(.A1(new_n1444_), .A2(new_n1445_), .ZN(new_n1446_));
  NOR2_X1    g1395(.A1(new_n1391_), .A2(new_n1179_), .ZN(new_n1447_));
  NAND3_X1   g1396(.A1(new_n1389_), .A2(new_n640_), .A3(new_n614_), .ZN(new_n1448_));
  OAI21_X1   g1397(.A1(new_n1144_), .A2(new_n459_), .B(new_n1122_), .ZN(new_n1449_));
  OAI21_X1   g1398(.A1(new_n1449_), .A2(new_n371_), .B(new_n428_), .ZN(new_n1450_));
  NAND2_X1   g1399(.A1(new_n1450_), .A2(new_n1448_), .ZN(new_n1451_));
  AOI21_X1   g1400(.A1(new_n1451_), .A2(new_n1387_), .B(new_n1178_), .ZN(new_n1452_));
  NOR2_X1    g1401(.A1(new_n1452_), .A2(new_n1447_), .ZN(new_n1453_));
  NOR4_X1    g1402(.A1(new_n428_), .A2(new_n1014_), .A3(new_n758_), .A4(new_n1061_), .ZN(new_n1454_));
  NOR2_X1    g1403(.A1(new_n1446_), .A2(new_n1443_), .ZN(new_n1455_));
  NAND3_X1   g1404(.A1(new_n1092_), .A2(new_n802_), .A3(new_n809_), .ZN(new_n1456_));
  NAND4_X1   g1405(.A1(new_n1100_), .A2(new_n1113_), .A3(new_n809_), .A4(new_n1106_), .ZN(new_n1457_));
  NAND2_X1   g1406(.A1(new_n1457_), .A2(new_n803_), .ZN(new_n1458_));
  AOI21_X1   g1407(.A1(new_n1458_), .A2(new_n1456_), .B(new_n808_), .ZN(new_n1459_));
  NOR3_X1    g1408(.A1(new_n1459_), .A2(new_n1444_), .A3(new_n1445_), .ZN(new_n1460_));
  NOR3_X1    g1409(.A1(new_n1455_), .A2(new_n1460_), .A3(new_n1454_), .ZN(new_n1461_));
  NOR3_X1    g1410(.A1(new_n925_), .A2(new_n1014_), .A3(new_n1050_), .ZN(new_n1462_));
  AOI21_X1   g1411(.A1(new_n925_), .A2(new_n1014_), .B(new_n1149_), .ZN(new_n1463_));
  AOI21_X1   g1412(.A1(new_n925_), .A2(new_n798_), .B(new_n1151_), .ZN(new_n1464_));
  NOR2_X1    g1413(.A1(new_n1464_), .A2(new_n1463_), .ZN(new_n1465_));
  NOR3_X1    g1414(.A1(new_n1465_), .A2(new_n1051_), .A3(new_n1223_), .ZN(new_n1466_));
  OAI21_X1   g1415(.A1(new_n1466_), .A2(new_n1462_), .B(new_n1251_), .ZN(new_n1467_));
  OAI21_X1   g1416(.A1(new_n1455_), .A2(new_n1460_), .B(new_n1454_), .ZN(new_n1468_));
  AOI21_X1   g1417(.A1(new_n1467_), .A2(new_n1468_), .B(new_n1461_), .ZN(new_n1469_));
  NOR3_X1    g1418(.A1(new_n1469_), .A2(new_n1453_), .A3(new_n1446_), .ZN(new_n1470_));
  NAND4_X1   g1419(.A1(new_n599_), .A2(new_n613_), .A3(new_n607_), .A4(new_n1122_), .ZN(new_n1471_));
  NAND2_X1   g1420(.A1(new_n1471_), .A2(new_n798_), .ZN(new_n1472_));
  AOI21_X1   g1421(.A1(new_n614_), .A2(new_n1121_), .B(new_n758_), .ZN(new_n1473_));
  NAND2_X1   g1422(.A1(new_n1473_), .A2(new_n1472_), .ZN(new_n1474_));
  NAND3_X1   g1423(.A1(new_n1451_), .A2(new_n1178_), .A3(new_n1387_), .ZN(new_n1475_));
  NAND2_X1   g1424(.A1(new_n1391_), .A2(new_n1179_), .ZN(new_n1476_));
  NAND2_X1   g1425(.A1(new_n1475_), .A2(new_n1476_), .ZN(new_n1477_));
  INV_X1     g1426(.I(new_n1454_), .ZN(new_n1478_));
  NAND2_X1   g1427(.A1(new_n1474_), .A2(new_n1459_), .ZN(new_n1479_));
  NAND3_X1   g1428(.A1(new_n1443_), .A2(new_n1472_), .A3(new_n1473_), .ZN(new_n1480_));
  NAND3_X1   g1429(.A1(new_n1479_), .A2(new_n1480_), .A3(new_n1478_), .ZN(new_n1481_));
  INV_X1     g1430(.I(new_n1462_), .ZN(new_n1482_));
  OAI21_X1   g1431(.A1(new_n1251_), .A2(new_n798_), .B(new_n1151_), .ZN(new_n1483_));
  OAI21_X1   g1432(.A1(new_n1251_), .A2(new_n1014_), .B(new_n1149_), .ZN(new_n1484_));
  NAND2_X1   g1433(.A1(new_n1483_), .A2(new_n1484_), .ZN(new_n1485_));
  NAND3_X1   g1434(.A1(new_n1485_), .A2(new_n1050_), .A3(new_n1257_), .ZN(new_n1486_));
  AOI21_X1   g1435(.A1(new_n1486_), .A2(new_n1482_), .B(new_n925_), .ZN(new_n1487_));
  AOI21_X1   g1436(.A1(new_n1479_), .A2(new_n1480_), .B(new_n1478_), .ZN(new_n1488_));
  OAI21_X1   g1437(.A1(new_n1487_), .A2(new_n1488_), .B(new_n1481_), .ZN(new_n1489_));
  AOI21_X1   g1438(.A1(new_n1489_), .A2(new_n1477_), .B(new_n1474_), .ZN(new_n1490_));
  OAI21_X1   g1439(.A1(new_n1470_), .A2(new_n1490_), .B(new_n1443_), .ZN(new_n1491_));
  NAND3_X1   g1440(.A1(new_n1489_), .A2(new_n1474_), .A3(new_n1477_), .ZN(new_n1492_));
  OAI21_X1   g1441(.A1(new_n1469_), .A2(new_n1453_), .B(new_n1446_), .ZN(new_n1493_));
  NAND3_X1   g1442(.A1(new_n1493_), .A2(new_n1492_), .A3(new_n1459_), .ZN(new_n1494_));
  NAND2_X1   g1443(.A1(new_n1491_), .A2(new_n1494_), .ZN(new_n1495_));
  NAND2_X1   g1444(.A1(new_n1495_), .A2(new_n1432_), .ZN(new_n1496_));
  AOI21_X1   g1445(.A1(new_n1479_), .A2(new_n1480_), .B(new_n1454_), .ZN(new_n1497_));
  INV_X1     g1446(.I(new_n1497_), .ZN(new_n1498_));
  NAND3_X1   g1447(.A1(new_n1479_), .A2(new_n1480_), .A3(new_n1454_), .ZN(new_n1499_));
  AOI21_X1   g1448(.A1(new_n1498_), .A2(new_n1499_), .B(new_n1467_), .ZN(new_n1500_));
  AOI21_X1   g1449(.A1(new_n1481_), .A2(new_n1468_), .B(new_n1487_), .ZN(new_n1501_));
  OAI21_X1   g1450(.A1(new_n925_), .A2(new_n1061_), .B(new_n1014_), .ZN(new_n1502_));
  NOR4_X1    g1451(.A1(new_n1502_), .A2(new_n1014_), .A3(new_n1251_), .A4(new_n1051_), .ZN(new_n1503_));
  NAND3_X1   g1452(.A1(new_n1092_), .A2(new_n808_), .A3(new_n1151_), .ZN(new_n1504_));
  OAI21_X1   g1453(.A1(new_n1114_), .A2(new_n1149_), .B(new_n809_), .ZN(new_n1505_));
  AOI21_X1   g1454(.A1(new_n1505_), .A2(new_n1504_), .B(new_n1149_), .ZN(new_n1506_));
  NOR2_X1    g1455(.A1(new_n1503_), .A2(new_n1506_), .ZN(new_n1507_));
  NAND3_X1   g1456(.A1(new_n925_), .A2(new_n798_), .A3(new_n1122_), .ZN(new_n1508_));
  NOR4_X1    g1457(.A1(new_n1440_), .A2(new_n1050_), .A3(new_n1075_), .A4(new_n1151_), .ZN(new_n1509_));
  AOI21_X1   g1458(.A1(new_n1092_), .A2(new_n1051_), .B(new_n1149_), .ZN(new_n1510_));
  OAI21_X1   g1459(.A1(new_n1510_), .A2(new_n1509_), .B(new_n1051_), .ZN(new_n1511_));
  NOR2_X1    g1460(.A1(new_n1511_), .A2(new_n1508_), .ZN(new_n1512_));
  INV_X1     g1461(.I(new_n1512_), .ZN(new_n1513_));
  NAND2_X1   g1462(.A1(new_n1503_), .A2(new_n1506_), .ZN(new_n1514_));
  AOI21_X1   g1463(.A1(new_n1513_), .A2(new_n1514_), .B(new_n1507_), .ZN(new_n1515_));
  INV_X1     g1464(.I(new_n1515_), .ZN(new_n1516_));
  OAI21_X1   g1465(.A1(new_n1500_), .A2(new_n1501_), .B(new_n1516_), .ZN(new_n1517_));
  NOR4_X1    g1466(.A1(new_n1114_), .A2(new_n1051_), .A3(new_n1060_), .A4(new_n1121_), .ZN(new_n1518_));
  INV_X1     g1467(.I(new_n1518_), .ZN(new_n1519_));
  NAND3_X1   g1468(.A1(new_n1092_), .A2(new_n1050_), .A3(new_n1061_), .ZN(new_n1520_));
  NAND4_X1   g1469(.A1(new_n1100_), .A2(new_n1113_), .A3(new_n1061_), .A4(new_n1106_), .ZN(new_n1521_));
  NAND2_X1   g1470(.A1(new_n1521_), .A2(new_n1051_), .ZN(new_n1522_));
  NAND2_X1   g1471(.A1(new_n1522_), .A2(new_n1520_), .ZN(new_n1523_));
  NOR2_X1    g1472(.A1(new_n1521_), .A2(new_n1121_), .ZN(new_n1524_));
  AOI21_X1   g1473(.A1(new_n1523_), .A2(new_n1061_), .B(new_n1524_), .ZN(new_n1525_));
  NOR3_X1    g1474(.A1(new_n1251_), .A2(new_n798_), .A3(new_n1121_), .ZN(new_n1526_));
  NOR3_X1    g1475(.A1(new_n1251_), .A2(new_n1014_), .A3(new_n1122_), .ZN(new_n1527_));
  NOR2_X1    g1476(.A1(new_n1526_), .A2(new_n1527_), .ZN(new_n1528_));
  OAI21_X1   g1477(.A1(new_n1525_), .A2(new_n1528_), .B(new_n1519_), .ZN(new_n1529_));
  OAI21_X1   g1478(.A1(new_n925_), .A2(new_n1122_), .B(new_n1014_), .ZN(new_n1530_));
  NOR4_X1    g1479(.A1(new_n1530_), .A2(new_n1014_), .A3(new_n1251_), .A4(new_n1061_), .ZN(new_n1531_));
  NAND2_X1   g1480(.A1(new_n1529_), .A2(new_n1531_), .ZN(new_n1532_));
  NAND3_X1   g1481(.A1(new_n1092_), .A2(new_n1051_), .A3(new_n1149_), .ZN(new_n1533_));
  NAND4_X1   g1482(.A1(new_n1100_), .A2(new_n1113_), .A3(new_n1051_), .A4(new_n1106_), .ZN(new_n1534_));
  NAND2_X1   g1483(.A1(new_n1534_), .A2(new_n1151_), .ZN(new_n1535_));
  NAND2_X1   g1484(.A1(new_n1535_), .A2(new_n1533_), .ZN(new_n1536_));
  NAND3_X1   g1485(.A1(new_n1536_), .A2(new_n1051_), .A3(new_n1508_), .ZN(new_n1537_));
  NOR3_X1    g1486(.A1(new_n1251_), .A2(new_n1014_), .A3(new_n1121_), .ZN(new_n1538_));
  NAND2_X1   g1487(.A1(new_n1511_), .A2(new_n1538_), .ZN(new_n1539_));
  NAND2_X1   g1488(.A1(new_n1537_), .A2(new_n1539_), .ZN(new_n1540_));
  OAI21_X1   g1489(.A1(new_n1529_), .A2(new_n1531_), .B(new_n1540_), .ZN(new_n1541_));
  NAND3_X1   g1490(.A1(new_n799_), .A2(new_n1015_), .A3(new_n1121_), .ZN(new_n1542_));
  AOI21_X1   g1491(.A1(new_n1541_), .A2(new_n1532_), .B(new_n1542_), .ZN(new_n1543_));
  NAND3_X1   g1492(.A1(new_n1541_), .A2(new_n1532_), .A3(new_n1542_), .ZN(new_n1544_));
  AOI21_X1   g1493(.A1(new_n1251_), .A2(new_n1060_), .B(new_n798_), .ZN(new_n1545_));
  NAND4_X1   g1494(.A1(new_n1545_), .A2(new_n798_), .A3(new_n925_), .A4(new_n1050_), .ZN(new_n1546_));
  INV_X1     g1495(.I(new_n1506_), .ZN(new_n1547_));
  NOR2_X1    g1496(.A1(new_n1547_), .A2(new_n1546_), .ZN(new_n1548_));
  OAI21_X1   g1497(.A1(new_n1548_), .A2(new_n1507_), .B(new_n1513_), .ZN(new_n1549_));
  NAND2_X1   g1498(.A1(new_n1547_), .A2(new_n1546_), .ZN(new_n1550_));
  NAND3_X1   g1499(.A1(new_n1550_), .A2(new_n1514_), .A3(new_n1512_), .ZN(new_n1551_));
  NAND2_X1   g1500(.A1(new_n1549_), .A2(new_n1551_), .ZN(new_n1552_));
  AOI21_X1   g1501(.A1(new_n1544_), .A2(new_n1552_), .B(new_n1543_), .ZN(new_n1553_));
  NOR3_X1    g1502(.A1(new_n1500_), .A2(new_n1501_), .A3(new_n1516_), .ZN(new_n1554_));
  OAI21_X1   g1503(.A1(new_n1553_), .A2(new_n1554_), .B(new_n1517_), .ZN(new_n1555_));
  OAI21_X1   g1504(.A1(new_n1495_), .A2(new_n1432_), .B(new_n1555_), .ZN(new_n1556_));
  NOR2_X1    g1505(.A1(new_n1469_), .A2(new_n1453_), .ZN(new_n1557_));
  NAND2_X1   g1506(.A1(new_n1446_), .A2(new_n1459_), .ZN(new_n1558_));
  AOI21_X1   g1507(.A1(new_n1469_), .A2(new_n1453_), .B(new_n1558_), .ZN(new_n1559_));
  NOR2_X1    g1508(.A1(new_n1559_), .A2(new_n1557_), .ZN(new_n1560_));
  AOI21_X1   g1509(.A1(new_n1556_), .A2(new_n1496_), .B(new_n1560_), .ZN(new_n1561_));
  NAND3_X1   g1510(.A1(new_n1556_), .A2(new_n1496_), .A3(new_n1560_), .ZN(new_n1562_));
  NOR2_X1    g1511(.A1(new_n1252_), .A2(new_n803_), .ZN(new_n1563_));
  AOI21_X1   g1512(.A1(new_n803_), .A2(new_n1253_), .B(new_n1563_), .ZN(new_n1564_));
  NOR3_X1    g1513(.A1(new_n1564_), .A2(new_n808_), .A3(new_n1257_), .ZN(new_n1565_));
  NOR3_X1    g1514(.A1(new_n1564_), .A2(new_n809_), .A3(new_n1223_), .ZN(new_n1566_));
  OAI21_X1   g1515(.A1(new_n1565_), .A2(new_n1566_), .B(new_n1251_), .ZN(new_n1567_));
  NOR2_X1    g1516(.A1(new_n1370_), .A2(new_n1567_), .ZN(new_n1568_));
  MUX2_X1    g1517(.I0(new_n1019_), .I1(new_n869_), .S(new_n1149_), .Z(new_n1569_));
  NOR3_X1    g1518(.A1(new_n1569_), .A2(new_n1018_), .A3(new_n1050_), .ZN(new_n1570_));
  NOR3_X1    g1519(.A1(new_n1569_), .A2(new_n1017_), .A3(new_n1051_), .ZN(new_n1571_));
  OAI21_X1   g1520(.A1(new_n1570_), .A2(new_n1571_), .B(new_n1016_), .ZN(new_n1572_));
  NOR2_X1    g1521(.A1(new_n1572_), .A2(new_n1375_), .ZN(new_n1573_));
  OAI21_X1   g1522(.A1(new_n1568_), .A2(new_n1573_), .B(new_n1377_), .ZN(new_n1574_));
  NOR2_X1    g1523(.A1(new_n1572_), .A2(new_n1567_), .ZN(new_n1575_));
  OAI21_X1   g1524(.A1(new_n1376_), .A2(new_n1575_), .B(new_n1378_), .ZN(new_n1576_));
  NAND2_X1   g1525(.A1(new_n1407_), .A2(new_n1417_), .ZN(new_n1577_));
  NAND2_X1   g1526(.A1(new_n1179_), .A2(new_n1385_), .ZN(new_n1578_));
  OAI22_X1   g1527(.A1(new_n1392_), .A2(new_n1385_), .B1(new_n1391_), .B2(new_n1578_), .ZN(new_n1579_));
  INV_X1     g1528(.I(new_n1579_), .ZN(new_n1580_));
  NAND3_X1   g1529(.A1(new_n1577_), .A2(new_n1423_), .A3(new_n1580_), .ZN(new_n1581_));
  AOI21_X1   g1530(.A1(new_n1426_), .A2(new_n1427_), .B(new_n1339_), .ZN(new_n1582_));
  NOR2_X1    g1531(.A1(new_n1422_), .A2(new_n1415_), .ZN(new_n1583_));
  OAI21_X1   g1532(.A1(new_n1582_), .A2(new_n1583_), .B(new_n1423_), .ZN(new_n1584_));
  NAND2_X1   g1533(.A1(new_n1584_), .A2(new_n1579_), .ZN(new_n1585_));
  NAND2_X1   g1534(.A1(new_n1585_), .A2(new_n1581_), .ZN(new_n1586_));
  NAND3_X1   g1535(.A1(new_n1586_), .A2(new_n1574_), .A3(new_n1576_), .ZN(new_n1587_));
  NAND2_X1   g1536(.A1(new_n1574_), .A2(new_n1576_), .ZN(new_n1588_));
  NOR2_X1    g1537(.A1(new_n1584_), .A2(new_n1579_), .ZN(new_n1589_));
  AOI21_X1   g1538(.A1(new_n1577_), .A2(new_n1423_), .B(new_n1580_), .ZN(new_n1590_));
  NOR2_X1    g1539(.A1(new_n1589_), .A2(new_n1590_), .ZN(new_n1591_));
  NAND2_X1   g1540(.A1(new_n1588_), .A2(new_n1591_), .ZN(new_n1592_));
  NAND2_X1   g1541(.A1(new_n1592_), .A2(new_n1587_), .ZN(new_n1593_));
  AOI21_X1   g1542(.A1(new_n1593_), .A2(new_n1562_), .B(new_n1561_), .ZN(new_n1594_));
  INV_X1     g1543(.I(new_n1584_), .ZN(new_n1595_));
  NOR2_X1    g1544(.A1(new_n1595_), .A2(new_n1579_), .ZN(new_n1596_));
  NAND2_X1   g1545(.A1(new_n1595_), .A2(new_n1579_), .ZN(new_n1597_));
  AOI21_X1   g1546(.A1(new_n1588_), .A2(new_n1597_), .B(new_n1596_), .ZN(new_n1598_));
  NOR2_X1    g1547(.A1(new_n1594_), .A2(new_n1598_), .ZN(new_n1599_));
  INV_X1     g1548(.I(new_n1344_), .ZN(new_n1600_));
  OAI21_X1   g1549(.A1(new_n1363_), .A2(new_n1364_), .B(new_n1600_), .ZN(new_n1601_));
  NAND2_X1   g1550(.A1(new_n1572_), .A2(new_n1567_), .ZN(new_n1602_));
  OAI21_X1   g1551(.A1(new_n1377_), .A2(new_n1575_), .B(new_n1602_), .ZN(new_n1603_));
  NAND3_X1   g1552(.A1(new_n1603_), .A2(new_n1601_), .A3(new_n1362_), .ZN(new_n1604_));
  OR2_X2     g1553(.A1(new_n1397_), .A2(new_n1399_), .Z(new_n1605_));
  AOI21_X1   g1554(.A1(new_n1401_), .A2(new_n1604_), .B(new_n1605_), .ZN(new_n1606_));
  AOI21_X1   g1555(.A1(new_n1362_), .A2(new_n1601_), .B(new_n1603_), .ZN(new_n1607_));
  NOR3_X1    g1556(.A1(new_n1381_), .A2(new_n1607_), .A3(new_n1400_), .ZN(new_n1608_));
  NOR2_X1    g1557(.A1(new_n1606_), .A2(new_n1608_), .ZN(new_n1609_));
  AOI21_X1   g1558(.A1(new_n1594_), .A2(new_n1598_), .B(new_n1609_), .ZN(new_n1610_));
  OAI21_X1   g1559(.A1(new_n1610_), .A2(new_n1599_), .B(new_n1403_), .ZN(new_n1611_));
  NOR3_X1    g1560(.A1(new_n1610_), .A2(new_n1599_), .A3(new_n1403_), .ZN(new_n1612_));
  NOR2_X1    g1561(.A1(new_n695_), .A2(new_n1382_), .ZN(new_n1613_));
  NAND2_X1   g1562(.A1(new_n695_), .A2(new_n1382_), .ZN(new_n1614_));
  NOR2_X1    g1563(.A1(new_n1393_), .A2(new_n1121_), .ZN(new_n1615_));
  AOI21_X1   g1564(.A1(new_n1615_), .A2(new_n1614_), .B(new_n1613_), .ZN(new_n1616_));
  NOR2_X1    g1565(.A1(new_n1184_), .A2(new_n1050_), .ZN(new_n1617_));
  AOI21_X1   g1566(.A1(new_n1183_), .A2(new_n1050_), .B(new_n1617_), .ZN(new_n1618_));
  NOR3_X1    g1567(.A1(new_n1618_), .A2(new_n1182_), .A3(new_n1149_), .ZN(new_n1619_));
  NOR3_X1    g1568(.A1(new_n1618_), .A2(new_n1181_), .A3(new_n1151_), .ZN(new_n1620_));
  OAI21_X1   g1569(.A1(new_n1619_), .A2(new_n1620_), .B(new_n1180_), .ZN(new_n1621_));
  INV_X1     g1570(.I(new_n1621_), .ZN(new_n1622_));
  NOR2_X1    g1571(.A1(new_n1019_), .A2(new_n802_), .ZN(new_n1623_));
  AOI21_X1   g1572(.A1(new_n802_), .A2(new_n1197_), .B(new_n1623_), .ZN(new_n1624_));
  NOR3_X1    g1573(.A1(new_n1624_), .A2(new_n808_), .A3(new_n1018_), .ZN(new_n1625_));
  NOR3_X1    g1574(.A1(new_n1624_), .A2(new_n809_), .A3(new_n1017_), .ZN(new_n1626_));
  OAI21_X1   g1575(.A1(new_n1625_), .A2(new_n1626_), .B(new_n1016_), .ZN(new_n1627_));
  NAND2_X1   g1576(.A1(new_n1253_), .A2(new_n577_), .ZN(new_n1628_));
  OAI21_X1   g1577(.A1(new_n577_), .A2(new_n1252_), .B(new_n1628_), .ZN(new_n1629_));
  NAND3_X1   g1578(.A1(new_n1629_), .A2(new_n271_), .A3(new_n1223_), .ZN(new_n1630_));
  NAND3_X1   g1579(.A1(new_n1629_), .A2(new_n270_), .A3(new_n1257_), .ZN(new_n1631_));
  AOI21_X1   g1580(.A1(new_n1630_), .A2(new_n1631_), .B(new_n925_), .ZN(new_n1632_));
  INV_X1     g1581(.I(new_n1632_), .ZN(new_n1633_));
  NOR2_X1    g1582(.A1(new_n1627_), .A2(new_n1633_), .ZN(new_n1634_));
  NAND2_X1   g1583(.A1(new_n1627_), .A2(new_n1633_), .ZN(new_n1635_));
  INV_X1     g1584(.I(new_n1635_), .ZN(new_n1636_));
  OAI21_X1   g1585(.A1(new_n1636_), .A2(new_n1634_), .B(new_n1622_), .ZN(new_n1637_));
  NAND2_X1   g1586(.A1(new_n1627_), .A2(new_n1632_), .ZN(new_n1638_));
  INV_X1     g1587(.I(new_n1638_), .ZN(new_n1639_));
  NOR2_X1    g1588(.A1(new_n1627_), .A2(new_n1632_), .ZN(new_n1640_));
  OAI21_X1   g1589(.A1(new_n1639_), .A2(new_n1640_), .B(new_n1621_), .ZN(new_n1641_));
  NAND3_X1   g1590(.A1(new_n1637_), .A2(new_n1641_), .A3(new_n1616_), .ZN(new_n1642_));
  INV_X1     g1591(.I(new_n1616_), .ZN(new_n1643_));
  NAND2_X1   g1592(.A1(new_n1637_), .A2(new_n1641_), .ZN(new_n1644_));
  NAND2_X1   g1593(.A1(new_n1644_), .A2(new_n1643_), .ZN(new_n1645_));
  NAND2_X1   g1594(.A1(new_n1645_), .A2(new_n1642_), .ZN(new_n1646_));
  NOR4_X1    g1595(.A1(new_n690_), .A2(new_n559_), .A3(new_n694_), .A4(new_n1061_), .ZN(new_n1647_));
  INV_X1     g1596(.I(new_n1647_), .ZN(new_n1648_));
  INV_X1     g1597(.I(new_n1361_), .ZN(new_n1649_));
  OR2_X2     g1598(.A1(new_n1344_), .A2(new_n1354_), .Z(new_n1650_));
  OAI21_X1   g1599(.A1(new_n559_), .A2(new_n1121_), .B(new_n587_), .ZN(new_n1651_));
  NAND2_X1   g1600(.A1(new_n559_), .A2(new_n1121_), .ZN(new_n1652_));
  NAND3_X1   g1601(.A1(new_n1651_), .A2(new_n687_), .A3(new_n1652_), .ZN(new_n1653_));
  NAND2_X1   g1602(.A1(new_n1092_), .A2(new_n702_), .ZN(new_n1654_));
  XOR2_X1    g1603(.A1(new_n1654_), .A2(new_n708_), .Z(new_n1655_));
  NAND2_X1   g1604(.A1(new_n1655_), .A2(new_n702_), .ZN(new_n1656_));
  XNOR2_X1   g1605(.A1(new_n1656_), .A2(new_n1653_), .ZN(new_n1657_));
  INV_X1     g1606(.I(new_n1657_), .ZN(new_n1658_));
  NAND3_X1   g1607(.A1(new_n1650_), .A2(new_n1649_), .A3(new_n1658_), .ZN(new_n1659_));
  AOI21_X1   g1608(.A1(new_n1650_), .A2(new_n1649_), .B(new_n1658_), .ZN(new_n1660_));
  INV_X1     g1609(.I(new_n1660_), .ZN(new_n1661_));
  AOI21_X1   g1610(.A1(new_n1661_), .A2(new_n1659_), .B(new_n1648_), .ZN(new_n1662_));
  NAND2_X1   g1611(.A1(new_n1650_), .A2(new_n1649_), .ZN(new_n1663_));
  XOR2_X1    g1612(.A1(new_n1663_), .A2(new_n1657_), .Z(new_n1664_));
  AOI21_X1   g1613(.A1(new_n1664_), .A2(new_n1648_), .B(new_n1662_), .ZN(new_n1665_));
  XOR2_X1    g1614(.A1(new_n1665_), .A2(new_n1646_), .Z(new_n1666_));
  OAI21_X1   g1615(.A1(new_n1612_), .A2(new_n1666_), .B(new_n1611_), .ZN(new_n1667_));
  NOR2_X1    g1616(.A1(new_n1644_), .A2(new_n1616_), .ZN(new_n1668_));
  NAND2_X1   g1617(.A1(new_n1644_), .A2(new_n1616_), .ZN(new_n1669_));
  AOI21_X1   g1618(.A1(new_n1665_), .A2(new_n1669_), .B(new_n1668_), .ZN(new_n1670_));
  INV_X1     g1619(.I(new_n1670_), .ZN(new_n1671_));
  NAND2_X1   g1620(.A1(new_n1667_), .A2(new_n1671_), .ZN(new_n1672_));
  NAND2_X1   g1621(.A1(new_n1659_), .A2(new_n1648_), .ZN(new_n1673_));
  NAND2_X1   g1622(.A1(new_n1673_), .A2(new_n1661_), .ZN(new_n1674_));
  NOR4_X1    g1623(.A1(new_n687_), .A2(new_n559_), .A3(new_n587_), .A4(new_n1051_), .ZN(new_n1675_));
  NAND2_X1   g1624(.A1(new_n1253_), .A2(new_n702_), .ZN(new_n1676_));
  OAI21_X1   g1625(.A1(new_n702_), .A2(new_n1252_), .B(new_n1676_), .ZN(new_n1677_));
  NAND3_X1   g1626(.A1(new_n1677_), .A2(new_n577_), .A3(new_n1223_), .ZN(new_n1678_));
  NAND3_X1   g1627(.A1(new_n1677_), .A2(new_n576_), .A3(new_n1257_), .ZN(new_n1679_));
  AOI21_X1   g1628(.A1(new_n1678_), .A2(new_n1679_), .B(new_n925_), .ZN(new_n1680_));
  NAND2_X1   g1629(.A1(new_n1092_), .A2(new_n711_), .ZN(new_n1681_));
  XOR2_X1    g1630(.A1(new_n1681_), .A2(new_n875_), .Z(new_n1682_));
  NOR2_X1    g1631(.A1(new_n1682_), .A2(new_n708_), .ZN(new_n1683_));
  XOR2_X1    g1632(.A1(new_n1680_), .A2(new_n1683_), .Z(new_n1684_));
  NAND2_X1   g1633(.A1(new_n1684_), .A2(new_n1675_), .ZN(new_n1685_));
  INV_X1     g1634(.I(new_n1675_), .ZN(new_n1686_));
  NAND2_X1   g1635(.A1(new_n1680_), .A2(new_n1683_), .ZN(new_n1687_));
  NOR2_X1    g1636(.A1(new_n1680_), .A2(new_n1683_), .ZN(new_n1688_));
  INV_X1     g1637(.I(new_n1688_), .ZN(new_n1689_));
  NAND2_X1   g1638(.A1(new_n1689_), .A2(new_n1687_), .ZN(new_n1690_));
  NAND2_X1   g1639(.A1(new_n1690_), .A2(new_n1686_), .ZN(new_n1691_));
  NAND2_X1   g1640(.A1(new_n1691_), .A2(new_n1685_), .ZN(new_n1692_));
  XOR2_X1    g1641(.A1(new_n1674_), .A2(new_n1692_), .Z(new_n1693_));
  INV_X1     g1642(.I(new_n1634_), .ZN(new_n1694_));
  AOI21_X1   g1643(.A1(new_n1621_), .A2(new_n1694_), .B(new_n1636_), .ZN(new_n1695_));
  NOR4_X1    g1644(.A1(new_n642_), .A2(new_n587_), .A3(new_n616_), .A4(new_n809_), .ZN(new_n1696_));
  INV_X1     g1645(.I(new_n1696_), .ZN(new_n1697_));
  NOR2_X1    g1646(.A1(new_n1656_), .A2(new_n1653_), .ZN(new_n1698_));
  NAND2_X1   g1647(.A1(new_n1340_), .A2(new_n271_), .ZN(new_n1699_));
  NAND2_X1   g1648(.A1(new_n1197_), .A2(new_n270_), .ZN(new_n1700_));
  NAND2_X1   g1649(.A1(new_n1699_), .A2(new_n1700_), .ZN(new_n1701_));
  NAND3_X1   g1650(.A1(new_n1701_), .A2(new_n803_), .A3(new_n1017_), .ZN(new_n1702_));
  NAND3_X1   g1651(.A1(new_n1701_), .A2(new_n802_), .A3(new_n1018_), .ZN(new_n1703_));
  NAND2_X1   g1652(.A1(new_n1702_), .A2(new_n1703_), .ZN(new_n1704_));
  NAND3_X1   g1653(.A1(new_n1704_), .A2(new_n1016_), .A3(new_n1698_), .ZN(new_n1705_));
  INV_X1     g1654(.I(new_n1698_), .ZN(new_n1706_));
  MUX2_X1    g1655(.I0(new_n869_), .I1(new_n1019_), .S(new_n271_), .Z(new_n1707_));
  NOR3_X1    g1656(.A1(new_n1707_), .A2(new_n802_), .A3(new_n1018_), .ZN(new_n1708_));
  NOR3_X1    g1657(.A1(new_n1707_), .A2(new_n803_), .A3(new_n1017_), .ZN(new_n1709_));
  OAI21_X1   g1658(.A1(new_n1708_), .A2(new_n1709_), .B(new_n1016_), .ZN(new_n1710_));
  NAND2_X1   g1659(.A1(new_n1710_), .A2(new_n1706_), .ZN(new_n1711_));
  AOI21_X1   g1660(.A1(new_n1705_), .A2(new_n1711_), .B(new_n1697_), .ZN(new_n1712_));
  NAND3_X1   g1661(.A1(new_n1704_), .A2(new_n1706_), .A3(new_n1016_), .ZN(new_n1713_));
  NAND2_X1   g1662(.A1(new_n1710_), .A2(new_n1698_), .ZN(new_n1714_));
  AOI21_X1   g1663(.A1(new_n1713_), .A2(new_n1714_), .B(new_n1696_), .ZN(new_n1715_));
  NOR2_X1    g1664(.A1(new_n559_), .A2(new_n1122_), .ZN(new_n1716_));
  NOR2_X1    g1665(.A1(new_n550_), .A2(new_n1121_), .ZN(new_n1717_));
  OAI21_X1   g1666(.A1(new_n1716_), .A2(new_n1717_), .B(new_n266_), .ZN(new_n1718_));
  INV_X1     g1667(.I(new_n1718_), .ZN(new_n1719_));
  OAI21_X1   g1668(.A1(new_n1712_), .A2(new_n1715_), .B(new_n1719_), .ZN(new_n1720_));
  NOR2_X1    g1669(.A1(new_n1710_), .A2(new_n1706_), .ZN(new_n1721_));
  AOI21_X1   g1670(.A1(new_n1704_), .A2(new_n1016_), .B(new_n1698_), .ZN(new_n1722_));
  OAI21_X1   g1671(.A1(new_n1722_), .A2(new_n1721_), .B(new_n1696_), .ZN(new_n1723_));
  NOR2_X1    g1672(.A1(new_n1710_), .A2(new_n1698_), .ZN(new_n1724_));
  AOI21_X1   g1673(.A1(new_n1704_), .A2(new_n1016_), .B(new_n1706_), .ZN(new_n1725_));
  OAI21_X1   g1674(.A1(new_n1725_), .A2(new_n1724_), .B(new_n1697_), .ZN(new_n1726_));
  NAND3_X1   g1675(.A1(new_n1723_), .A2(new_n1726_), .A3(new_n1718_), .ZN(new_n1727_));
  AOI21_X1   g1676(.A1(new_n1720_), .A2(new_n1727_), .B(new_n1695_), .ZN(new_n1728_));
  OAI21_X1   g1677(.A1(new_n1622_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n1729_));
  NAND3_X1   g1678(.A1(new_n1723_), .A2(new_n1726_), .A3(new_n1719_), .ZN(new_n1730_));
  OAI21_X1   g1679(.A1(new_n1712_), .A2(new_n1715_), .B(new_n1718_), .ZN(new_n1731_));
  AOI21_X1   g1680(.A1(new_n1731_), .A2(new_n1730_), .B(new_n1729_), .ZN(new_n1732_));
  NOR2_X1    g1681(.A1(new_n1728_), .A2(new_n1732_), .ZN(new_n1733_));
  XOR2_X1    g1682(.A1(new_n1693_), .A2(new_n1733_), .Z(new_n1734_));
  OAI21_X1   g1683(.A1(new_n1667_), .A2(new_n1671_), .B(new_n1734_), .ZN(new_n1735_));
  NAND2_X1   g1684(.A1(new_n1735_), .A2(new_n1672_), .ZN(new_n1736_));
  NOR3_X1    g1685(.A1(new_n1712_), .A2(new_n1715_), .A3(new_n1719_), .ZN(new_n1737_));
  AOI21_X1   g1686(.A1(new_n1729_), .A2(new_n1720_), .B(new_n1737_), .ZN(new_n1738_));
  AOI21_X1   g1687(.A1(new_n1697_), .A2(new_n1705_), .B(new_n1722_), .ZN(new_n1739_));
  INV_X1     g1688(.I(new_n1739_), .ZN(new_n1740_));
  AOI21_X1   g1689(.A1(new_n1680_), .A2(new_n1683_), .B(new_n1675_), .ZN(new_n1741_));
  NOR2_X1    g1690(.A1(new_n1741_), .A2(new_n1688_), .ZN(new_n1742_));
  NAND2_X1   g1691(.A1(new_n684_), .A2(new_n550_), .ZN(new_n1743_));
  NAND2_X1   g1692(.A1(new_n687_), .A2(new_n559_), .ZN(new_n1744_));
  NAND2_X1   g1693(.A1(new_n1743_), .A2(new_n1744_), .ZN(new_n1745_));
  OAI21_X1   g1694(.A1(new_n686_), .A2(new_n682_), .B(new_n1051_), .ZN(new_n1746_));
  NAND3_X1   g1695(.A1(new_n683_), .A2(new_n663_), .A3(new_n1050_), .ZN(new_n1747_));
  NAND2_X1   g1696(.A1(new_n489_), .A2(new_n1050_), .ZN(new_n1748_));
  NAND2_X1   g1697(.A1(new_n587_), .A2(new_n1051_), .ZN(new_n1749_));
  NAND4_X1   g1698(.A1(new_n1749_), .A2(new_n1747_), .A3(new_n1746_), .A4(new_n1748_), .ZN(new_n1750_));
  NAND4_X1   g1699(.A1(new_n710_), .A2(new_n1745_), .A3(new_n1750_), .A4(new_n1151_), .ZN(new_n1751_));
  NAND4_X1   g1700(.A1(new_n693_), .A2(new_n1745_), .A3(new_n1750_), .A4(new_n1149_), .ZN(new_n1752_));
  AOI21_X1   g1701(.A1(new_n1752_), .A2(new_n1751_), .B(new_n930_), .ZN(new_n1753_));
  NOR2_X1    g1702(.A1(new_n1157_), .A2(new_n1753_), .ZN(new_n1754_));
  MUX2_X1    g1703(.I0(new_n1197_), .I1(new_n1340_), .S(new_n577_), .Z(new_n1755_));
  NAND3_X1   g1704(.A1(new_n1755_), .A2(new_n271_), .A3(new_n1017_), .ZN(new_n1756_));
  NAND3_X1   g1705(.A1(new_n1755_), .A2(new_n270_), .A3(new_n1018_), .ZN(new_n1757_));
  AOI21_X1   g1706(.A1(new_n1756_), .A2(new_n1757_), .B(new_n1339_), .ZN(new_n1758_));
  NOR2_X1    g1707(.A1(new_n1758_), .A2(new_n1153_), .ZN(new_n1759_));
  OAI21_X1   g1708(.A1(new_n1759_), .A2(new_n1754_), .B(new_n1171_), .ZN(new_n1760_));
  NOR2_X1    g1709(.A1(new_n1157_), .A2(new_n1153_), .ZN(new_n1761_));
  NOR2_X1    g1710(.A1(new_n1758_), .A2(new_n1753_), .ZN(new_n1762_));
  OAI21_X1   g1711(.A1(new_n1762_), .A2(new_n1761_), .B(new_n1172_), .ZN(new_n1763_));
  AOI21_X1   g1712(.A1(new_n1760_), .A2(new_n1763_), .B(new_n1742_), .ZN(new_n1764_));
  INV_X1     g1713(.I(new_n1742_), .ZN(new_n1765_));
  NAND2_X1   g1714(.A1(new_n1758_), .A2(new_n1153_), .ZN(new_n1766_));
  NAND2_X1   g1715(.A1(new_n1157_), .A2(new_n1753_), .ZN(new_n1767_));
  AOI21_X1   g1716(.A1(new_n1766_), .A2(new_n1767_), .B(new_n1172_), .ZN(new_n1768_));
  NAND2_X1   g1717(.A1(new_n1758_), .A2(new_n1753_), .ZN(new_n1769_));
  NAND2_X1   g1718(.A1(new_n1157_), .A2(new_n1153_), .ZN(new_n1770_));
  AOI21_X1   g1719(.A1(new_n1769_), .A2(new_n1770_), .B(new_n1171_), .ZN(new_n1771_));
  NOR3_X1    g1720(.A1(new_n1765_), .A2(new_n1768_), .A3(new_n1771_), .ZN(new_n1772_));
  OAI21_X1   g1721(.A1(new_n1772_), .A2(new_n1764_), .B(new_n1740_), .ZN(new_n1773_));
  AOI21_X1   g1722(.A1(new_n1760_), .A2(new_n1763_), .B(new_n1765_), .ZN(new_n1774_));
  NOR3_X1    g1723(.A1(new_n1768_), .A2(new_n1771_), .A3(new_n1742_), .ZN(new_n1775_));
  OAI21_X1   g1724(.A1(new_n1774_), .A2(new_n1775_), .B(new_n1739_), .ZN(new_n1776_));
  XOR2_X1    g1725(.A1(new_n1291_), .A2(new_n1285_), .Z(new_n1777_));
  NAND2_X1   g1726(.A1(new_n1777_), .A2(new_n1298_), .ZN(new_n1778_));
  AOI21_X1   g1727(.A1(new_n1301_), .A2(new_n1292_), .B(new_n1298_), .ZN(new_n1779_));
  INV_X1     g1728(.I(new_n1779_), .ZN(new_n1780_));
  NAND2_X1   g1729(.A1(new_n1780_), .A2(new_n1778_), .ZN(new_n1781_));
  NAND3_X1   g1730(.A1(new_n1773_), .A2(new_n1776_), .A3(new_n1781_), .ZN(new_n1782_));
  OAI21_X1   g1731(.A1(new_n1768_), .A2(new_n1771_), .B(new_n1765_), .ZN(new_n1783_));
  NAND3_X1   g1732(.A1(new_n1760_), .A2(new_n1763_), .A3(new_n1742_), .ZN(new_n1784_));
  AOI21_X1   g1733(.A1(new_n1783_), .A2(new_n1784_), .B(new_n1739_), .ZN(new_n1785_));
  OAI21_X1   g1734(.A1(new_n1768_), .A2(new_n1771_), .B(new_n1742_), .ZN(new_n1786_));
  NAND3_X1   g1735(.A1(new_n1765_), .A2(new_n1760_), .A3(new_n1763_), .ZN(new_n1787_));
  AOI21_X1   g1736(.A1(new_n1787_), .A2(new_n1786_), .B(new_n1740_), .ZN(new_n1788_));
  AOI21_X1   g1737(.A1(new_n1777_), .A2(new_n1298_), .B(new_n1779_), .ZN(new_n1789_));
  OAI21_X1   g1738(.A1(new_n1788_), .A2(new_n1785_), .B(new_n1789_), .ZN(new_n1790_));
  AOI21_X1   g1739(.A1(new_n1790_), .A2(new_n1782_), .B(new_n1738_), .ZN(new_n1791_));
  INV_X1     g1740(.I(new_n1738_), .ZN(new_n1792_));
  OAI21_X1   g1741(.A1(new_n1788_), .A2(new_n1785_), .B(new_n1781_), .ZN(new_n1793_));
  NAND3_X1   g1742(.A1(new_n1773_), .A2(new_n1776_), .A3(new_n1789_), .ZN(new_n1794_));
  AOI21_X1   g1743(.A1(new_n1793_), .A2(new_n1794_), .B(new_n1792_), .ZN(new_n1795_));
  NOR2_X1    g1744(.A1(new_n1791_), .A2(new_n1795_), .ZN(new_n1796_));
  AOI21_X1   g1745(.A1(new_n1773_), .A2(new_n1776_), .B(new_n1789_), .ZN(new_n1797_));
  AOI21_X1   g1746(.A1(new_n1792_), .A2(new_n1794_), .B(new_n1797_), .ZN(new_n1798_));
  AOI21_X1   g1747(.A1(new_n1284_), .A2(new_n1307_), .B(new_n1302_), .ZN(new_n1799_));
  XOR2_X1    g1748(.A1(new_n1275_), .A2(new_n1270_), .Z(new_n1800_));
  NOR2_X1    g1749(.A1(new_n1800_), .A2(new_n1278_), .ZN(new_n1801_));
  INV_X1     g1750(.I(new_n1282_), .ZN(new_n1802_));
  OAI21_X1   g1751(.A1(new_n1801_), .A2(new_n1802_), .B(new_n1306_), .ZN(new_n1803_));
  NAND3_X1   g1752(.A1(new_n1268_), .A2(new_n1277_), .A3(new_n1282_), .ZN(new_n1804_));
  AOI21_X1   g1753(.A1(new_n1803_), .A2(new_n1804_), .B(new_n1303_), .ZN(new_n1805_));
  NOR2_X1    g1754(.A1(new_n1799_), .A2(new_n1805_), .ZN(new_n1806_));
  NOR2_X1    g1755(.A1(new_n1774_), .A2(new_n1775_), .ZN(new_n1807_));
  NAND2_X1   g1756(.A1(new_n1163_), .A2(new_n1168_), .ZN(new_n1808_));
  NAND2_X1   g1757(.A1(new_n1766_), .A2(new_n1767_), .ZN(new_n1809_));
  NAND3_X1   g1758(.A1(new_n1809_), .A2(new_n1808_), .A3(new_n1769_), .ZN(new_n1810_));
  NOR2_X1    g1759(.A1(new_n1157_), .A2(new_n1153_), .ZN(new_n1811_));
  INV_X1     g1760(.I(new_n1811_), .ZN(new_n1812_));
  AOI21_X1   g1761(.A1(new_n1810_), .A2(new_n1812_), .B(new_n1171_), .ZN(new_n1813_));
  NOR2_X1    g1762(.A1(new_n1759_), .A2(new_n1754_), .ZN(new_n1814_));
  NOR3_X1    g1763(.A1(new_n1814_), .A2(new_n1169_), .A3(new_n1761_), .ZN(new_n1815_));
  NOR3_X1    g1764(.A1(new_n1815_), .A2(new_n1172_), .A3(new_n1811_), .ZN(new_n1816_));
  NOR2_X1    g1765(.A1(new_n1816_), .A2(new_n1813_), .ZN(new_n1817_));
  NOR3_X1    g1766(.A1(new_n1817_), .A2(new_n1764_), .A3(new_n1807_), .ZN(new_n1818_));
  AOI21_X1   g1767(.A1(new_n1760_), .A2(new_n1763_), .B(new_n1742_), .ZN(new_n1819_));
  OAI21_X1   g1768(.A1(new_n1818_), .A2(new_n1819_), .B(new_n1739_), .ZN(new_n1820_));
  NAND2_X1   g1769(.A1(new_n1787_), .A2(new_n1786_), .ZN(new_n1821_));
  OAI21_X1   g1770(.A1(new_n1815_), .A2(new_n1811_), .B(new_n1172_), .ZN(new_n1822_));
  NAND3_X1   g1771(.A1(new_n1810_), .A2(new_n1171_), .A3(new_n1812_), .ZN(new_n1823_));
  NAND2_X1   g1772(.A1(new_n1822_), .A2(new_n1823_), .ZN(new_n1824_));
  NAND3_X1   g1773(.A1(new_n1824_), .A2(new_n1783_), .A3(new_n1821_), .ZN(new_n1825_));
  INV_X1     g1774(.I(new_n1819_), .ZN(new_n1826_));
  NAND3_X1   g1775(.A1(new_n1825_), .A2(new_n1826_), .A3(new_n1740_), .ZN(new_n1827_));
  NAND3_X1   g1776(.A1(new_n1820_), .A2(new_n1827_), .A3(new_n1806_), .ZN(new_n1828_));
  AOI21_X1   g1777(.A1(new_n1277_), .A2(new_n1282_), .B(new_n1306_), .ZN(new_n1829_));
  INV_X1     g1778(.I(new_n1307_), .ZN(new_n1830_));
  OAI21_X1   g1779(.A1(new_n1830_), .A2(new_n1829_), .B(new_n1303_), .ZN(new_n1831_));
  AOI21_X1   g1780(.A1(new_n1277_), .A2(new_n1282_), .B(new_n1268_), .ZN(new_n1832_));
  NOR3_X1    g1781(.A1(new_n1802_), .A2(new_n1306_), .A3(new_n1801_), .ZN(new_n1833_));
  OAI21_X1   g1782(.A1(new_n1832_), .A2(new_n1833_), .B(new_n1302_), .ZN(new_n1834_));
  NAND2_X1   g1783(.A1(new_n1831_), .A2(new_n1834_), .ZN(new_n1835_));
  AOI21_X1   g1784(.A1(new_n1825_), .A2(new_n1826_), .B(new_n1740_), .ZN(new_n1836_));
  NOR3_X1    g1785(.A1(new_n1818_), .A2(new_n1739_), .A3(new_n1819_), .ZN(new_n1837_));
  OAI21_X1   g1786(.A1(new_n1837_), .A2(new_n1836_), .B(new_n1835_), .ZN(new_n1838_));
  NAND3_X1   g1787(.A1(new_n1838_), .A2(new_n1828_), .A3(new_n1798_), .ZN(new_n1839_));
  INV_X1     g1788(.I(new_n1798_), .ZN(new_n1840_));
  NOR3_X1    g1789(.A1(new_n1837_), .A2(new_n1836_), .A3(new_n1835_), .ZN(new_n1841_));
  AOI21_X1   g1790(.A1(new_n1820_), .A2(new_n1827_), .B(new_n1806_), .ZN(new_n1842_));
  OAI21_X1   g1791(.A1(new_n1841_), .A2(new_n1842_), .B(new_n1840_), .ZN(new_n1843_));
  NAND3_X1   g1792(.A1(new_n1843_), .A2(new_n1839_), .A3(new_n1796_), .ZN(new_n1844_));
  INV_X1     g1793(.I(new_n1692_), .ZN(new_n1845_));
  AOI21_X1   g1794(.A1(new_n1723_), .A2(new_n1726_), .B(new_n1718_), .ZN(new_n1846_));
  OAI21_X1   g1795(.A1(new_n1846_), .A2(new_n1737_), .B(new_n1729_), .ZN(new_n1847_));
  NOR3_X1    g1796(.A1(new_n1712_), .A2(new_n1715_), .A3(new_n1718_), .ZN(new_n1848_));
  AOI21_X1   g1797(.A1(new_n1723_), .A2(new_n1726_), .B(new_n1719_), .ZN(new_n1849_));
  OAI21_X1   g1798(.A1(new_n1849_), .A2(new_n1848_), .B(new_n1695_), .ZN(new_n1850_));
  AOI21_X1   g1799(.A1(new_n1850_), .A2(new_n1847_), .B(new_n1845_), .ZN(new_n1851_));
  NAND3_X1   g1800(.A1(new_n1850_), .A2(new_n1847_), .A3(new_n1845_), .ZN(new_n1852_));
  AOI21_X1   g1801(.A1(new_n1674_), .A2(new_n1852_), .B(new_n1851_), .ZN(new_n1853_));
  INV_X1     g1802(.I(new_n1796_), .ZN(new_n1854_));
  NOR3_X1    g1803(.A1(new_n1841_), .A2(new_n1842_), .A3(new_n1840_), .ZN(new_n1855_));
  AOI21_X1   g1804(.A1(new_n1838_), .A2(new_n1828_), .B(new_n1798_), .ZN(new_n1856_));
  OAI21_X1   g1805(.A1(new_n1855_), .A2(new_n1856_), .B(new_n1854_), .ZN(new_n1857_));
  NAND2_X1   g1806(.A1(new_n1857_), .A2(new_n1853_), .ZN(new_n1858_));
  NAND4_X1   g1807(.A1(new_n1858_), .A2(new_n1736_), .A3(new_n1338_), .A4(new_n1844_), .ZN(new_n1859_));
  NOR3_X1    g1808(.A1(new_n1855_), .A2(new_n1856_), .A3(new_n1854_), .ZN(new_n1860_));
  AOI21_X1   g1809(.A1(new_n1853_), .A2(new_n1857_), .B(new_n1860_), .ZN(new_n1861_));
  AOI21_X1   g1810(.A1(new_n1861_), .A2(new_n1736_), .B(new_n1338_), .ZN(new_n1862_));
  AOI21_X1   g1811(.A1(new_n1838_), .A2(new_n1828_), .B(new_n1840_), .ZN(new_n1863_));
  INV_X1     g1812(.I(new_n1863_), .ZN(new_n1864_));
  NAND2_X1   g1813(.A1(new_n1835_), .A2(new_n1817_), .ZN(new_n1865_));
  NOR2_X1    g1814(.A1(new_n1772_), .A2(new_n1739_), .ZN(new_n1866_));
  OAI22_X1   g1815(.A1(new_n1835_), .A2(new_n1817_), .B1(new_n1764_), .B2(new_n1866_), .ZN(new_n1867_));
  NAND2_X1   g1816(.A1(new_n1867_), .A2(new_n1865_), .ZN(new_n1868_));
  INV_X1     g1817(.I(new_n1868_), .ZN(new_n1869_));
  NOR2_X1    g1818(.A1(new_n1864_), .A2(new_n1869_), .ZN(new_n1870_));
  INV_X1     g1819(.I(new_n1870_), .ZN(new_n1871_));
  OAI21_X1   g1820(.A1(new_n1862_), .A2(new_n1871_), .B(new_n1859_), .ZN(new_n1872_));
  NAND2_X1   g1821(.A1(new_n1327_), .A2(new_n1310_), .ZN(new_n1873_));
  NAND2_X1   g1822(.A1(new_n1873_), .A2(new_n1326_), .ZN(new_n1874_));
  INV_X1     g1823(.I(new_n1874_), .ZN(new_n1875_));
  OAI21_X1   g1824(.A1(new_n1207_), .A2(new_n1211_), .B(new_n1174_), .ZN(new_n1876_));
  NOR3_X1    g1825(.A1(new_n1174_), .A2(new_n1207_), .A3(new_n1211_), .ZN(new_n1877_));
  NOR2_X1    g1826(.A1(new_n1130_), .A2(new_n1213_), .ZN(new_n1878_));
  INV_X1     g1827(.I(new_n1878_), .ZN(new_n1879_));
  OAI21_X1   g1828(.A1(new_n1877_), .A2(new_n1879_), .B(new_n1876_), .ZN(new_n1880_));
  NOR4_X1    g1829(.A1(new_n690_), .A2(new_n271_), .A3(new_n694_), .A4(new_n559_), .ZN(new_n1881_));
  NOR2_X1    g1830(.A1(new_n1184_), .A2(new_n576_), .ZN(new_n1882_));
  AOI21_X1   g1831(.A1(new_n576_), .A2(new_n1183_), .B(new_n1882_), .ZN(new_n1883_));
  NOR3_X1    g1832(.A1(new_n1883_), .A2(new_n1182_), .A3(new_n721_), .ZN(new_n1884_));
  NOR3_X1    g1833(.A1(new_n1883_), .A2(new_n1181_), .A3(new_n702_), .ZN(new_n1885_));
  OAI21_X1   g1834(.A1(new_n1884_), .A2(new_n1885_), .B(new_n1180_), .ZN(new_n1886_));
  INV_X1     g1835(.I(new_n1886_), .ZN(new_n1887_));
  NOR2_X1    g1836(.A1(new_n1019_), .A2(new_n645_), .ZN(new_n1888_));
  AOI21_X1   g1837(.A1(new_n645_), .A2(new_n1197_), .B(new_n1888_), .ZN(new_n1889_));
  NOR2_X1    g1838(.A1(new_n1889_), .A2(new_n1017_), .ZN(new_n1890_));
  NOR2_X1    g1839(.A1(new_n1889_), .A2(new_n708_), .ZN(new_n1891_));
  XOR2_X1    g1840(.A1(new_n1890_), .A2(new_n1891_), .Z(new_n1892_));
  NAND2_X1   g1841(.A1(new_n1892_), .A2(new_n1016_), .ZN(new_n1893_));
  NOR2_X1    g1842(.A1(new_n1893_), .A2(new_n1887_), .ZN(new_n1894_));
  XNOR2_X1   g1843(.A1(new_n1890_), .A2(new_n1891_), .ZN(new_n1895_));
  NOR2_X1    g1844(.A1(new_n1895_), .A2(new_n1339_), .ZN(new_n1896_));
  NOR2_X1    g1845(.A1(new_n1896_), .A2(new_n1886_), .ZN(new_n1897_));
  OAI21_X1   g1846(.A1(new_n1897_), .A2(new_n1894_), .B(new_n1881_), .ZN(new_n1898_));
  INV_X1     g1847(.I(new_n1881_), .ZN(new_n1899_));
  NOR2_X1    g1848(.A1(new_n1893_), .A2(new_n1886_), .ZN(new_n1900_));
  NOR2_X1    g1849(.A1(new_n1896_), .A2(new_n1887_), .ZN(new_n1901_));
  OAI21_X1   g1850(.A1(new_n1901_), .A2(new_n1900_), .B(new_n1899_), .ZN(new_n1902_));
  XOR2_X1    g1851(.A1(new_n266_), .A2(new_n1050_), .Z(new_n1903_));
  NAND3_X1   g1852(.A1(new_n1902_), .A2(new_n1898_), .A3(new_n1903_), .ZN(new_n1904_));
  NAND2_X1   g1853(.A1(new_n1896_), .A2(new_n1886_), .ZN(new_n1905_));
  NAND2_X1   g1854(.A1(new_n1893_), .A2(new_n1887_), .ZN(new_n1906_));
  AOI21_X1   g1855(.A1(new_n1905_), .A2(new_n1906_), .B(new_n1899_), .ZN(new_n1907_));
  NAND2_X1   g1856(.A1(new_n1896_), .A2(new_n1887_), .ZN(new_n1908_));
  NAND2_X1   g1857(.A1(new_n1893_), .A2(new_n1886_), .ZN(new_n1909_));
  AOI21_X1   g1858(.A1(new_n1908_), .A2(new_n1909_), .B(new_n1881_), .ZN(new_n1910_));
  INV_X1     g1859(.I(new_n1903_), .ZN(new_n1911_));
  OAI21_X1   g1860(.A1(new_n1910_), .A2(new_n1907_), .B(new_n1911_), .ZN(new_n1912_));
  OAI21_X1   g1861(.A1(new_n1189_), .A2(new_n1202_), .B(new_n1176_), .ZN(new_n1913_));
  NAND2_X1   g1862(.A1(new_n1913_), .A2(new_n1210_), .ZN(new_n1914_));
  INV_X1     g1863(.I(new_n1914_), .ZN(new_n1915_));
  NOR2_X1    g1864(.A1(new_n1056_), .A2(new_n1151_), .ZN(new_n1916_));
  AOI21_X1   g1865(.A1(new_n571_), .A2(new_n1151_), .B(new_n1916_), .ZN(new_n1917_));
  NOR3_X1    g1866(.A1(new_n1917_), .A2(new_n580_), .A3(new_n808_), .ZN(new_n1918_));
  NOR3_X1    g1867(.A1(new_n1917_), .A2(new_n565_), .A3(new_n809_), .ZN(new_n1919_));
  OAI21_X1   g1868(.A1(new_n1919_), .A2(new_n1918_), .B(new_n562_), .ZN(new_n1920_));
  NAND2_X1   g1869(.A1(new_n1253_), .A2(new_n438_), .ZN(new_n1921_));
  OAI21_X1   g1870(.A1(new_n438_), .A2(new_n1252_), .B(new_n1921_), .ZN(new_n1922_));
  NAND3_X1   g1871(.A1(new_n1922_), .A2(new_n875_), .A3(new_n1223_), .ZN(new_n1923_));
  NAND3_X1   g1872(.A1(new_n1922_), .A2(new_n645_), .A3(new_n1257_), .ZN(new_n1924_));
  AOI21_X1   g1873(.A1(new_n1923_), .A2(new_n1924_), .B(new_n925_), .ZN(new_n1925_));
  NAND3_X1   g1874(.A1(new_n1925_), .A2(new_n266_), .A3(new_n1061_), .ZN(new_n1926_));
  XOR2_X1    g1875(.A1(new_n1920_), .A2(new_n1926_), .Z(new_n1927_));
  INV_X1     g1876(.I(new_n1926_), .ZN(new_n1928_));
  NAND2_X1   g1877(.A1(new_n1920_), .A2(new_n1928_), .ZN(new_n1929_));
  NAND2_X1   g1878(.A1(new_n567_), .A2(new_n1149_), .ZN(new_n1930_));
  OAI21_X1   g1879(.A1(new_n572_), .A2(new_n1149_), .B(new_n1930_), .ZN(new_n1931_));
  NAND3_X1   g1880(.A1(new_n1931_), .A2(new_n565_), .A3(new_n809_), .ZN(new_n1932_));
  NAND3_X1   g1881(.A1(new_n1931_), .A2(new_n580_), .A3(new_n808_), .ZN(new_n1933_));
  NAND2_X1   g1882(.A1(new_n1933_), .A2(new_n1932_), .ZN(new_n1934_));
  NAND3_X1   g1883(.A1(new_n1934_), .A2(new_n562_), .A3(new_n1926_), .ZN(new_n1935_));
  NAND2_X1   g1884(.A1(new_n1935_), .A2(new_n1929_), .ZN(new_n1936_));
  NAND3_X1   g1885(.A1(new_n1936_), .A2(new_n1913_), .A3(new_n1210_), .ZN(new_n1937_));
  OAI21_X1   g1886(.A1(new_n1915_), .A2(new_n1927_), .B(new_n1937_), .ZN(new_n1938_));
  NAND3_X1   g1887(.A1(new_n1912_), .A2(new_n1938_), .A3(new_n1904_), .ZN(new_n1939_));
  NOR3_X1    g1888(.A1(new_n1910_), .A2(new_n1907_), .A3(new_n1911_), .ZN(new_n1940_));
  AOI21_X1   g1889(.A1(new_n1902_), .A2(new_n1898_), .B(new_n1903_), .ZN(new_n1941_));
  NOR2_X1    g1890(.A1(new_n1915_), .A2(new_n1927_), .ZN(new_n1942_));
  AOI21_X1   g1891(.A1(new_n1929_), .A2(new_n1935_), .B(new_n1914_), .ZN(new_n1943_));
  NOR2_X1    g1892(.A1(new_n1942_), .A2(new_n1943_), .ZN(new_n1944_));
  OAI21_X1   g1893(.A1(new_n1940_), .A2(new_n1941_), .B(new_n1944_), .ZN(new_n1945_));
  AOI21_X1   g1894(.A1(new_n1945_), .A2(new_n1939_), .B(new_n1880_), .ZN(new_n1946_));
  NOR2_X1    g1895(.A1(new_n1215_), .A2(new_n1212_), .ZN(new_n1947_));
  NOR2_X1    g1896(.A1(new_n1877_), .A2(new_n1879_), .ZN(new_n1948_));
  NOR2_X1    g1897(.A1(new_n1948_), .A2(new_n1947_), .ZN(new_n1949_));
  NOR3_X1    g1898(.A1(new_n1944_), .A2(new_n1941_), .A3(new_n1940_), .ZN(new_n1950_));
  AOI21_X1   g1899(.A1(new_n1904_), .A2(new_n1912_), .B(new_n1938_), .ZN(new_n1951_));
  NOR3_X1    g1900(.A1(new_n1949_), .A2(new_n1950_), .A3(new_n1951_), .ZN(new_n1952_));
  OAI21_X1   g1901(.A1(new_n1952_), .A2(new_n1946_), .B(new_n1875_), .ZN(new_n1953_));
  OAI21_X1   g1902(.A1(new_n1950_), .A2(new_n1951_), .B(new_n1949_), .ZN(new_n1954_));
  NAND3_X1   g1903(.A1(new_n1880_), .A2(new_n1945_), .A3(new_n1939_), .ZN(new_n1955_));
  NAND3_X1   g1904(.A1(new_n1954_), .A2(new_n1955_), .A3(new_n1874_), .ZN(new_n1956_));
  NAND2_X1   g1905(.A1(new_n1956_), .A2(new_n1953_), .ZN(new_n1957_));
  NAND2_X1   g1906(.A1(new_n1874_), .A2(new_n1911_), .ZN(new_n1958_));
  OAI22_X1   g1907(.A1(new_n1874_), .A2(new_n1911_), .B1(new_n1907_), .B2(new_n1910_), .ZN(new_n1959_));
  NAND2_X1   g1908(.A1(new_n1959_), .A2(new_n1958_), .ZN(new_n1960_));
  NOR2_X1    g1909(.A1(new_n1184_), .A2(new_n721_), .ZN(new_n1961_));
  AOI21_X1   g1910(.A1(new_n1183_), .A2(new_n721_), .B(new_n1961_), .ZN(new_n1962_));
  NOR3_X1    g1911(.A1(new_n1962_), .A2(new_n1182_), .A3(new_n708_), .ZN(new_n1963_));
  NOR3_X1    g1912(.A1(new_n1962_), .A2(new_n1181_), .A3(new_n711_), .ZN(new_n1964_));
  OAI21_X1   g1913(.A1(new_n1963_), .A2(new_n1964_), .B(new_n1180_), .ZN(new_n1965_));
  XOR2_X1    g1914(.A1(new_n266_), .A2(new_n1149_), .Z(new_n1966_));
  NOR2_X1    g1915(.A1(new_n566_), .A2(new_n1050_), .ZN(new_n1967_));
  NAND4_X1   g1916(.A1(new_n1967_), .A2(new_n437_), .A3(new_n1014_), .A4(new_n1251_), .ZN(new_n1968_));
  NOR2_X1    g1917(.A1(new_n1968_), .A2(new_n1966_), .ZN(new_n1969_));
  NAND2_X1   g1918(.A1(new_n1968_), .A2(new_n1966_), .ZN(new_n1970_));
  INV_X1     g1919(.I(new_n1970_), .ZN(new_n1971_));
  NOR2_X1    g1920(.A1(new_n1971_), .A2(new_n1969_), .ZN(new_n1972_));
  NOR2_X1    g1921(.A1(new_n1965_), .A2(new_n1972_), .ZN(new_n1973_));
  XNOR2_X1   g1922(.A1(new_n1968_), .A2(new_n1966_), .ZN(new_n1974_));
  INV_X1     g1923(.I(new_n1974_), .ZN(new_n1975_));
  AOI21_X1   g1924(.A1(new_n1965_), .A2(new_n1975_), .B(new_n1973_), .ZN(new_n1976_));
  XOR2_X1    g1925(.A1(new_n1960_), .A2(new_n1976_), .Z(new_n1977_));
  NAND2_X1   g1926(.A1(new_n1914_), .A2(new_n1935_), .ZN(new_n1978_));
  NAND2_X1   g1927(.A1(new_n1978_), .A2(new_n1929_), .ZN(new_n1979_));
  AOI21_X1   g1928(.A1(new_n1899_), .A2(new_n1908_), .B(new_n1901_), .ZN(new_n1980_));
  INV_X1     g1929(.I(new_n1032_), .ZN(new_n1981_));
  NAND2_X1   g1930(.A1(new_n1026_), .A2(new_n1035_), .ZN(new_n1982_));
  NAND2_X1   g1931(.A1(new_n1982_), .A2(new_n1981_), .ZN(new_n1983_));
  NOR2_X1    g1932(.A1(new_n1033_), .A2(new_n1025_), .ZN(new_n1984_));
  NOR2_X1    g1933(.A1(new_n983_), .A2(new_n1034_), .ZN(new_n1985_));
  OAI21_X1   g1934(.A1(new_n1985_), .A2(new_n1984_), .B(new_n1032_), .ZN(new_n1986_));
  AOI21_X1   g1935(.A1(new_n1983_), .A2(new_n1986_), .B(new_n1980_), .ZN(new_n1987_));
  OAI21_X1   g1936(.A1(new_n1881_), .A2(new_n1900_), .B(new_n1909_), .ZN(new_n1988_));
  AOI21_X1   g1937(.A1(new_n1026_), .A2(new_n1035_), .B(new_n1032_), .ZN(new_n1989_));
  INV_X1     g1938(.I(new_n1986_), .ZN(new_n1990_));
  NOR3_X1    g1939(.A1(new_n1990_), .A2(new_n1988_), .A3(new_n1989_), .ZN(new_n1991_));
  OAI21_X1   g1940(.A1(new_n1987_), .A2(new_n1991_), .B(new_n1979_), .ZN(new_n1992_));
  INV_X1     g1941(.I(new_n1979_), .ZN(new_n1993_));
  AOI21_X1   g1942(.A1(new_n1983_), .A2(new_n1986_), .B(new_n1988_), .ZN(new_n1994_));
  NOR3_X1    g1943(.A1(new_n1990_), .A2(new_n1980_), .A3(new_n1989_), .ZN(new_n1995_));
  OAI21_X1   g1944(.A1(new_n1995_), .A2(new_n1994_), .B(new_n1993_), .ZN(new_n1996_));
  NAND2_X1   g1945(.A1(new_n1992_), .A2(new_n1996_), .ZN(new_n1997_));
  NAND2_X1   g1946(.A1(new_n1880_), .A2(new_n1938_), .ZN(new_n1998_));
  NOR3_X1    g1947(.A1(new_n1941_), .A2(new_n1940_), .A3(new_n1875_), .ZN(new_n1999_));
  AOI21_X1   g1948(.A1(new_n1912_), .A2(new_n1904_), .B(new_n1874_), .ZN(new_n2000_));
  OAI22_X1   g1949(.A1(new_n1999_), .A2(new_n2000_), .B1(new_n1880_), .B2(new_n1938_), .ZN(new_n2001_));
  AOI21_X1   g1950(.A1(new_n2001_), .A2(new_n1998_), .B(new_n1997_), .ZN(new_n2002_));
  OAI21_X1   g1951(.A1(new_n1990_), .A2(new_n1989_), .B(new_n1988_), .ZN(new_n2003_));
  NAND3_X1   g1952(.A1(new_n1983_), .A2(new_n1980_), .A3(new_n1986_), .ZN(new_n2004_));
  AOI21_X1   g1953(.A1(new_n2003_), .A2(new_n2004_), .B(new_n1993_), .ZN(new_n2005_));
  OAI21_X1   g1954(.A1(new_n1990_), .A2(new_n1989_), .B(new_n1980_), .ZN(new_n2006_));
  NAND3_X1   g1955(.A1(new_n1983_), .A2(new_n1986_), .A3(new_n1988_), .ZN(new_n2007_));
  AOI21_X1   g1956(.A1(new_n2006_), .A2(new_n2007_), .B(new_n1979_), .ZN(new_n2008_));
  NOR2_X1    g1957(.A1(new_n2008_), .A2(new_n2005_), .ZN(new_n2009_));
  NOR2_X1    g1958(.A1(new_n1949_), .A2(new_n1944_), .ZN(new_n2010_));
  NAND3_X1   g1959(.A1(new_n1912_), .A2(new_n1904_), .A3(new_n1874_), .ZN(new_n2011_));
  OAI21_X1   g1960(.A1(new_n1941_), .A2(new_n1940_), .B(new_n1875_), .ZN(new_n2012_));
  AOI22_X1   g1961(.A1(new_n1949_), .A2(new_n1944_), .B1(new_n2012_), .B2(new_n2011_), .ZN(new_n2013_));
  NOR3_X1    g1962(.A1(new_n2013_), .A2(new_n2009_), .A3(new_n2010_), .ZN(new_n2014_));
  OAI21_X1   g1963(.A1(new_n2014_), .A2(new_n2002_), .B(new_n1977_), .ZN(new_n2015_));
  INV_X1     g1964(.I(new_n1976_), .ZN(new_n2016_));
  XOR2_X1    g1965(.A1(new_n1960_), .A2(new_n2016_), .Z(new_n2017_));
  AOI21_X1   g1966(.A1(new_n2001_), .A2(new_n1998_), .B(new_n2009_), .ZN(new_n2018_));
  NOR3_X1    g1967(.A1(new_n2013_), .A2(new_n1997_), .A3(new_n2010_), .ZN(new_n2019_));
  OAI21_X1   g1968(.A1(new_n2019_), .A2(new_n2018_), .B(new_n2017_), .ZN(new_n2020_));
  NAND2_X1   g1969(.A1(new_n2015_), .A2(new_n2020_), .ZN(new_n2021_));
  NOR2_X1    g1970(.A1(new_n2021_), .A2(new_n1957_), .ZN(new_n2022_));
  INV_X1     g1971(.I(new_n1332_), .ZN(new_n2023_));
  AOI21_X1   g1972(.A1(new_n1220_), .A2(new_n1221_), .B(new_n1129_), .ZN(new_n2024_));
  NOR3_X1    g1973(.A1(new_n1218_), .A2(new_n1130_), .A3(new_n1214_), .ZN(new_n2025_));
  NOR3_X1    g1974(.A1(new_n2025_), .A2(new_n2024_), .A3(new_n1330_), .ZN(new_n2026_));
  NOR2_X1    g1975(.A1(new_n2026_), .A2(new_n2023_), .ZN(new_n2027_));
  NAND2_X1   g1976(.A1(new_n2021_), .A2(new_n1957_), .ZN(new_n2028_));
  AOI21_X1   g1977(.A1(new_n2027_), .A2(new_n2028_), .B(new_n2022_), .ZN(new_n2029_));
  NAND2_X1   g1978(.A1(new_n1872_), .A2(new_n2029_), .ZN(new_n2030_));
  AOI21_X1   g1979(.A1(new_n1979_), .A2(new_n2006_), .B(new_n1995_), .ZN(new_n2031_));
  INV_X1     g1980(.I(new_n977_), .ZN(new_n2032_));
  AOI21_X1   g1981(.A1(new_n2032_), .A2(new_n1038_), .B(new_n1036_), .ZN(new_n2033_));
  INV_X1     g1982(.I(new_n976_), .ZN(new_n2034_));
  NOR2_X1    g1983(.A1(new_n973_), .A2(new_n2034_), .ZN(new_n2035_));
  INV_X1     g1984(.I(new_n2035_), .ZN(new_n2036_));
  NAND2_X1   g1985(.A1(new_n973_), .A2(new_n2034_), .ZN(new_n2037_));
  AOI21_X1   g1986(.A1(new_n2036_), .A2(new_n2037_), .B(new_n1037_), .ZN(new_n2038_));
  AOI21_X1   g1987(.A1(new_n1965_), .A2(new_n1970_), .B(new_n1969_), .ZN(new_n2039_));
  INV_X1     g1988(.I(new_n2039_), .ZN(new_n2040_));
  OAI21_X1   g1989(.A1(new_n2033_), .A2(new_n2038_), .B(new_n2040_), .ZN(new_n2041_));
  INV_X1     g1990(.I(new_n1038_), .ZN(new_n2042_));
  OAI21_X1   g1991(.A1(new_n2042_), .A2(new_n977_), .B(new_n1037_), .ZN(new_n2043_));
  INV_X1     g1992(.I(new_n2037_), .ZN(new_n2044_));
  OAI21_X1   g1993(.A1(new_n2044_), .A2(new_n2035_), .B(new_n1036_), .ZN(new_n2045_));
  NAND3_X1   g1994(.A1(new_n2043_), .A2(new_n2045_), .A3(new_n2039_), .ZN(new_n2046_));
  AOI21_X1   g1995(.A1(new_n2041_), .A2(new_n2046_), .B(new_n2031_), .ZN(new_n2047_));
  INV_X1     g1996(.I(new_n2031_), .ZN(new_n2048_));
  NAND3_X1   g1997(.A1(new_n2043_), .A2(new_n2045_), .A3(new_n2040_), .ZN(new_n2049_));
  OAI21_X1   g1998(.A1(new_n2033_), .A2(new_n2038_), .B(new_n2039_), .ZN(new_n2050_));
  AOI21_X1   g1999(.A1(new_n2050_), .A2(new_n2049_), .B(new_n2048_), .ZN(new_n2051_));
  NOR2_X1    g2000(.A1(new_n2047_), .A2(new_n2051_), .ZN(new_n2052_));
  NOR2_X1    g2001(.A1(new_n2030_), .A2(new_n2052_), .ZN(new_n2053_));
  NOR2_X1    g2002(.A1(new_n2013_), .A2(new_n2010_), .ZN(new_n2054_));
  XOR2_X1    g2003(.A1(new_n2017_), .A2(new_n2009_), .Z(new_n2055_));
  NAND2_X1   g2004(.A1(new_n2055_), .A2(new_n2054_), .ZN(new_n2056_));
  INV_X1     g2005(.I(new_n1960_), .ZN(new_n2057_));
  NOR2_X1    g2006(.A1(new_n2057_), .A2(new_n2016_), .ZN(new_n2058_));
  AOI21_X1   g2007(.A1(new_n2057_), .A2(new_n2016_), .B(new_n1997_), .ZN(new_n2059_));
  NOR2_X1    g2008(.A1(new_n2059_), .A2(new_n2058_), .ZN(new_n2060_));
  NOR2_X1    g2009(.A1(new_n2056_), .A2(new_n2060_), .ZN(new_n2061_));
  INV_X1     g2010(.I(new_n2061_), .ZN(new_n2062_));
  AOI21_X1   g2011(.A1(new_n2030_), .A2(new_n2052_), .B(new_n2062_), .ZN(new_n2063_));
  NOR2_X1    g2012(.A1(new_n2063_), .A2(new_n2053_), .ZN(new_n2064_));
  INV_X1     g2013(.I(new_n968_), .ZN(new_n2065_));
  AOI21_X1   g2014(.A1(new_n2065_), .A2(new_n1041_), .B(new_n1039_), .ZN(new_n2066_));
  NAND2_X1   g2015(.A1(new_n961_), .A2(new_n966_), .ZN(new_n2067_));
  OAI21_X1   g2016(.A1(new_n960_), .A2(new_n958_), .B(new_n967_), .ZN(new_n2068_));
  AOI21_X1   g2017(.A1(new_n2068_), .A2(new_n2067_), .B(new_n1040_), .ZN(new_n2069_));
  NOR2_X1    g2018(.A1(new_n2066_), .A2(new_n2069_), .ZN(new_n2070_));
  OAI21_X1   g2019(.A1(new_n955_), .A2(new_n956_), .B(new_n495_), .ZN(new_n2071_));
  NAND3_X1   g2020(.A1(new_n950_), .A2(new_n953_), .A3(new_n496_), .ZN(new_n2072_));
  AOI21_X1   g2021(.A1(new_n2071_), .A2(new_n2072_), .B(new_n1042_), .ZN(new_n2073_));
  NOR2_X1    g2022(.A1(new_n1044_), .A2(new_n2073_), .ZN(new_n2074_));
  NAND2_X1   g2023(.A1(new_n2074_), .A2(new_n2070_), .ZN(new_n2075_));
  AOI21_X1   g2024(.A1(new_n2043_), .A2(new_n2045_), .B(new_n2039_), .ZN(new_n2076_));
  AOI21_X1   g2025(.A1(new_n2048_), .A2(new_n2046_), .B(new_n2076_), .ZN(new_n2077_));
  INV_X1     g2026(.I(new_n2077_), .ZN(new_n2078_));
  NOR2_X1    g2027(.A1(new_n2074_), .A2(new_n2070_), .ZN(new_n2079_));
  OAI21_X1   g2028(.A1(new_n2078_), .A2(new_n2079_), .B(new_n2075_), .ZN(new_n2080_));
  INV_X1     g2029(.I(new_n944_), .ZN(new_n2081_));
  XOR2_X1    g2030(.A1(new_n495_), .A2(new_n945_), .Z(new_n2082_));
  AOI21_X1   g2031(.A1(new_n2081_), .A2(new_n818_), .B(new_n2082_), .ZN(new_n2083_));
  AOI21_X1   g2032(.A1(new_n951_), .A2(new_n944_), .B(new_n2083_), .ZN(new_n2084_));
  OAI21_X1   g2033(.A1(new_n717_), .A2(new_n813_), .B(new_n812_), .ZN(new_n2085_));
  NAND2_X1   g2034(.A1(new_n494_), .A2(new_n272_), .ZN(new_n2086_));
  OAI21_X1   g2035(.A1(new_n494_), .A2(new_n272_), .B(new_n946_), .ZN(new_n2087_));
  NAND2_X1   g2036(.A1(new_n2087_), .A2(new_n2086_), .ZN(new_n2088_));
  INV_X1     g2037(.I(new_n2088_), .ZN(new_n2089_));
  NOR2_X1    g2038(.A1(new_n703_), .A2(new_n875_), .ZN(new_n2090_));
  AOI21_X1   g2039(.A1(new_n697_), .A2(new_n875_), .B(new_n2090_), .ZN(new_n2091_));
  NOR3_X1    g2040(.A1(new_n2091_), .A2(new_n437_), .A3(new_n693_), .ZN(new_n2092_));
  NOR3_X1    g2041(.A1(new_n2091_), .A2(new_n438_), .A3(new_n710_), .ZN(new_n2093_));
  OAI21_X1   g2042(.A1(new_n2093_), .A2(new_n2092_), .B(new_n692_), .ZN(new_n2094_));
  NOR2_X1    g2043(.A1(new_n1056_), .A2(new_n702_), .ZN(new_n2095_));
  AOI21_X1   g2044(.A1(new_n571_), .A2(new_n702_), .B(new_n2095_), .ZN(new_n2096_));
  NOR3_X1    g2045(.A1(new_n2096_), .A2(new_n580_), .A3(new_n708_), .ZN(new_n2097_));
  NOR3_X1    g2046(.A1(new_n2096_), .A2(new_n565_), .A3(new_n711_), .ZN(new_n2098_));
  OAI21_X1   g2047(.A1(new_n2097_), .A2(new_n2098_), .B(new_n562_), .ZN(new_n2099_));
  XNOR2_X1   g2048(.A1(new_n2094_), .A2(new_n2099_), .ZN(new_n2100_));
  NOR2_X1    g2049(.A1(new_n2094_), .A2(new_n2099_), .ZN(new_n2101_));
  NAND2_X1   g2050(.A1(new_n2094_), .A2(new_n2099_), .ZN(new_n2102_));
  INV_X1     g2051(.I(new_n2102_), .ZN(new_n2103_));
  OAI21_X1   g2052(.A1(new_n2103_), .A2(new_n2101_), .B(new_n2089_), .ZN(new_n2104_));
  OAI21_X1   g2053(.A1(new_n2089_), .A2(new_n2100_), .B(new_n2104_), .ZN(new_n2105_));
  XOR2_X1    g2054(.A1(new_n1178_), .A2(new_n270_), .Z(new_n2106_));
  NAND2_X1   g2055(.A1(new_n2106_), .A2(new_n577_), .ZN(new_n2107_));
  XOR2_X1    g2056(.A1(new_n2107_), .A2(new_n266_), .Z(new_n2108_));
  XOR2_X1    g2057(.A1(new_n2105_), .A2(new_n2108_), .Z(new_n2109_));
  INV_X1     g2058(.I(new_n2109_), .ZN(new_n2110_));
  INV_X1     g2059(.I(new_n2108_), .ZN(new_n2111_));
  NAND2_X1   g2060(.A1(new_n2105_), .A2(new_n2111_), .ZN(new_n2112_));
  NOR2_X1    g2061(.A1(new_n2105_), .A2(new_n2111_), .ZN(new_n2113_));
  INV_X1     g2062(.I(new_n2113_), .ZN(new_n2114_));
  AOI21_X1   g2063(.A1(new_n2114_), .A2(new_n2112_), .B(new_n2085_), .ZN(new_n2115_));
  AOI21_X1   g2064(.A1(new_n2110_), .A2(new_n2085_), .B(new_n2115_), .ZN(new_n2116_));
  NOR2_X1    g2065(.A1(new_n2084_), .A2(new_n2116_), .ZN(new_n2117_));
  OAI21_X1   g2066(.A1(new_n2064_), .A2(new_n2080_), .B(new_n2117_), .ZN(new_n2118_));
  NAND2_X1   g2067(.A1(new_n1423_), .A2(new_n1417_), .ZN(new_n2119_));
  NAND2_X1   g2068(.A1(new_n2119_), .A2(new_n1582_), .ZN(new_n2120_));
  NAND2_X1   g2069(.A1(new_n1429_), .A2(new_n1430_), .ZN(new_n2121_));
  NAND2_X1   g2070(.A1(new_n2121_), .A2(new_n1407_), .ZN(new_n2122_));
  NAND2_X1   g2071(.A1(new_n2120_), .A2(new_n2122_), .ZN(new_n2123_));
  AOI21_X1   g2072(.A1(new_n1493_), .A2(new_n1492_), .B(new_n1459_), .ZN(new_n2124_));
  NOR3_X1    g2073(.A1(new_n1470_), .A2(new_n1490_), .A3(new_n1443_), .ZN(new_n2125_));
  NOR2_X1    g2074(.A1(new_n2125_), .A2(new_n2124_), .ZN(new_n2126_));
  NOR2_X1    g2075(.A1(new_n2126_), .A2(new_n2123_), .ZN(new_n2127_));
  NOR3_X1    g2076(.A1(new_n1455_), .A2(new_n1460_), .A3(new_n1478_), .ZN(new_n2128_));
  OAI21_X1   g2077(.A1(new_n1497_), .A2(new_n2128_), .B(new_n1487_), .ZN(new_n2129_));
  OAI21_X1   g2078(.A1(new_n1461_), .A2(new_n1488_), .B(new_n1467_), .ZN(new_n2130_));
  AOI21_X1   g2079(.A1(new_n2130_), .A2(new_n2129_), .B(new_n1515_), .ZN(new_n2131_));
  NOR4_X1    g2080(.A1(new_n1440_), .A2(new_n1051_), .A3(new_n1060_), .A4(new_n1075_), .ZN(new_n2132_));
  AOI21_X1   g2081(.A1(new_n1092_), .A2(new_n1061_), .B(new_n1050_), .ZN(new_n2133_));
  OAI21_X1   g2082(.A1(new_n2133_), .A2(new_n2132_), .B(new_n1061_), .ZN(new_n2134_));
  INV_X1     g2083(.I(new_n1524_), .ZN(new_n2135_));
  NAND2_X1   g2084(.A1(new_n2134_), .A2(new_n2135_), .ZN(new_n2136_));
  NAND3_X1   g2085(.A1(new_n925_), .A2(new_n1014_), .A3(new_n1122_), .ZN(new_n2137_));
  NAND3_X1   g2086(.A1(new_n925_), .A2(new_n798_), .A3(new_n1121_), .ZN(new_n2138_));
  NAND2_X1   g2087(.A1(new_n2138_), .A2(new_n2137_), .ZN(new_n2139_));
  AOI21_X1   g2088(.A1(new_n2136_), .A2(new_n2139_), .B(new_n1518_), .ZN(new_n2140_));
  INV_X1     g2089(.I(new_n1531_), .ZN(new_n2141_));
  NOR2_X1    g2090(.A1(new_n2140_), .A2(new_n2141_), .ZN(new_n2142_));
  AOI22_X1   g2091(.A1(new_n2140_), .A2(new_n2141_), .B1(new_n1537_), .B2(new_n1539_), .ZN(new_n2143_));
  INV_X1     g2092(.I(new_n1542_), .ZN(new_n2144_));
  OAI21_X1   g2093(.A1(new_n2143_), .A2(new_n2142_), .B(new_n2144_), .ZN(new_n2145_));
  NOR3_X1    g2094(.A1(new_n2143_), .A2(new_n2142_), .A3(new_n2144_), .ZN(new_n2146_));
  INV_X1     g2095(.I(new_n1552_), .ZN(new_n2147_));
  OAI21_X1   g2096(.A1(new_n2147_), .A2(new_n2146_), .B(new_n2145_), .ZN(new_n2148_));
  NAND3_X1   g2097(.A1(new_n2130_), .A2(new_n2129_), .A3(new_n1515_), .ZN(new_n2149_));
  AOI21_X1   g2098(.A1(new_n2148_), .A2(new_n2149_), .B(new_n2131_), .ZN(new_n2150_));
  AOI21_X1   g2099(.A1(new_n2126_), .A2(new_n2123_), .B(new_n2150_), .ZN(new_n2151_));
  INV_X1     g2100(.I(new_n1560_), .ZN(new_n2152_));
  OAI21_X1   g2101(.A1(new_n2151_), .A2(new_n2127_), .B(new_n2152_), .ZN(new_n2153_));
  NOR3_X1    g2102(.A1(new_n2151_), .A2(new_n2127_), .A3(new_n2152_), .ZN(new_n2154_));
  NOR2_X1    g2103(.A1(new_n1588_), .A2(new_n1591_), .ZN(new_n2155_));
  NAND2_X1   g2104(.A1(new_n1572_), .A2(new_n1375_), .ZN(new_n2156_));
  NAND2_X1   g2105(.A1(new_n1370_), .A2(new_n1567_), .ZN(new_n2157_));
  AOI21_X1   g2106(.A1(new_n2157_), .A2(new_n2156_), .B(new_n1378_), .ZN(new_n2158_));
  AOI21_X1   g2107(.A1(new_n1379_), .A2(new_n1602_), .B(new_n1377_), .ZN(new_n2159_));
  NOR2_X1    g2108(.A1(new_n2158_), .A2(new_n2159_), .ZN(new_n2160_));
  NOR2_X1    g2109(.A1(new_n2160_), .A2(new_n1586_), .ZN(new_n2161_));
  NOR2_X1    g2110(.A1(new_n2161_), .A2(new_n2155_), .ZN(new_n2162_));
  OAI21_X1   g2111(.A1(new_n2162_), .A2(new_n2154_), .B(new_n2153_), .ZN(new_n2163_));
  INV_X1     g2112(.I(new_n1598_), .ZN(new_n2164_));
  NAND2_X1   g2113(.A1(new_n2163_), .A2(new_n2164_), .ZN(new_n2165_));
  OAI21_X1   g2114(.A1(new_n1381_), .A2(new_n1607_), .B(new_n1400_), .ZN(new_n2166_));
  NAND3_X1   g2115(.A1(new_n1401_), .A2(new_n1605_), .A3(new_n1604_), .ZN(new_n2167_));
  NAND2_X1   g2116(.A1(new_n2166_), .A2(new_n2167_), .ZN(new_n2168_));
  OAI21_X1   g2117(.A1(new_n2163_), .A2(new_n2164_), .B(new_n2168_), .ZN(new_n2169_));
  NAND3_X1   g2118(.A1(new_n2169_), .A2(new_n2165_), .A3(new_n1402_), .ZN(new_n2170_));
  INV_X1     g2119(.I(new_n1659_), .ZN(new_n2171_));
  OAI21_X1   g2120(.A1(new_n2171_), .A2(new_n1660_), .B(new_n1647_), .ZN(new_n2172_));
  XOR2_X1    g2121(.A1(new_n1663_), .A2(new_n1658_), .Z(new_n2173_));
  OAI21_X1   g2122(.A1(new_n2173_), .A2(new_n1647_), .B(new_n2172_), .ZN(new_n2174_));
  NAND3_X1   g2123(.A1(new_n2174_), .A2(new_n1642_), .A3(new_n1645_), .ZN(new_n2175_));
  NAND2_X1   g2124(.A1(new_n1665_), .A2(new_n1646_), .ZN(new_n2176_));
  NAND2_X1   g2125(.A1(new_n2176_), .A2(new_n2175_), .ZN(new_n2177_));
  NAND2_X1   g2126(.A1(new_n2170_), .A2(new_n2177_), .ZN(new_n2178_));
  AOI21_X1   g2127(.A1(new_n2178_), .A2(new_n1611_), .B(new_n1670_), .ZN(new_n2179_));
  NAND3_X1   g2128(.A1(new_n2178_), .A2(new_n1611_), .A3(new_n1670_), .ZN(new_n2180_));
  AOI21_X1   g2129(.A1(new_n2180_), .A2(new_n1734_), .B(new_n2179_), .ZN(new_n2181_));
  INV_X1     g2130(.I(new_n1674_), .ZN(new_n2182_));
  OAI21_X1   g2131(.A1(new_n1728_), .A2(new_n1732_), .B(new_n1692_), .ZN(new_n2183_));
  NOR3_X1    g2132(.A1(new_n1728_), .A2(new_n1732_), .A3(new_n1692_), .ZN(new_n2184_));
  OAI21_X1   g2133(.A1(new_n2182_), .A2(new_n2184_), .B(new_n2183_), .ZN(new_n2185_));
  AOI21_X1   g2134(.A1(new_n1843_), .A2(new_n1839_), .B(new_n1796_), .ZN(new_n2186_));
  OAI21_X1   g2135(.A1(new_n2185_), .A2(new_n2186_), .B(new_n1844_), .ZN(new_n2187_));
  NOR3_X1    g2136(.A1(new_n2187_), .A2(new_n1337_), .A3(new_n2181_), .ZN(new_n2188_));
  OAI21_X1   g2137(.A1(new_n2187_), .A2(new_n2181_), .B(new_n1337_), .ZN(new_n2189_));
  AOI21_X1   g2138(.A1(new_n2189_), .A2(new_n1870_), .B(new_n2188_), .ZN(new_n2190_));
  AOI21_X1   g2139(.A1(new_n1954_), .A2(new_n1955_), .B(new_n1874_), .ZN(new_n2191_));
  NOR3_X1    g2140(.A1(new_n1952_), .A2(new_n1946_), .A3(new_n1875_), .ZN(new_n2192_));
  NOR2_X1    g2141(.A1(new_n2191_), .A2(new_n2192_), .ZN(new_n2193_));
  OAI21_X1   g2142(.A1(new_n2013_), .A2(new_n2010_), .B(new_n2009_), .ZN(new_n2194_));
  NAND3_X1   g2143(.A1(new_n2001_), .A2(new_n1997_), .A3(new_n1998_), .ZN(new_n2195_));
  AOI21_X1   g2144(.A1(new_n2194_), .A2(new_n2195_), .B(new_n2017_), .ZN(new_n2196_));
  OAI21_X1   g2145(.A1(new_n2013_), .A2(new_n2010_), .B(new_n1997_), .ZN(new_n2197_));
  NAND3_X1   g2146(.A1(new_n2001_), .A2(new_n2009_), .A3(new_n1998_), .ZN(new_n2198_));
  AOI21_X1   g2147(.A1(new_n2197_), .A2(new_n2198_), .B(new_n1977_), .ZN(new_n2199_));
  NOR2_X1    g2148(.A1(new_n2196_), .A2(new_n2199_), .ZN(new_n2200_));
  NAND2_X1   g2149(.A1(new_n2200_), .A2(new_n2193_), .ZN(new_n2201_));
  OAI21_X1   g2150(.A1(new_n1334_), .A2(new_n1330_), .B(new_n1332_), .ZN(new_n2202_));
  NOR2_X1    g2151(.A1(new_n2200_), .A2(new_n2193_), .ZN(new_n2203_));
  OAI21_X1   g2152(.A1(new_n2202_), .A2(new_n2203_), .B(new_n2201_), .ZN(new_n2204_));
  NOR2_X1    g2153(.A1(new_n2190_), .A2(new_n2204_), .ZN(new_n2205_));
  INV_X1     g2154(.I(new_n2052_), .ZN(new_n2206_));
  NAND2_X1   g2155(.A1(new_n2205_), .A2(new_n2206_), .ZN(new_n2207_));
  OAI21_X1   g2156(.A1(new_n2205_), .A2(new_n2206_), .B(new_n2061_), .ZN(new_n2208_));
  NAND2_X1   g2157(.A1(new_n2208_), .A2(new_n2207_), .ZN(new_n2209_));
  INV_X1     g2158(.I(new_n2075_), .ZN(new_n2210_));
  NOR2_X1    g2159(.A1(new_n2079_), .A2(new_n2078_), .ZN(new_n2211_));
  NOR2_X1    g2160(.A1(new_n2211_), .A2(new_n2210_), .ZN(new_n2212_));
  INV_X1     g2161(.I(new_n2117_), .ZN(new_n2213_));
  NAND3_X1   g2162(.A1(new_n2209_), .A2(new_n2212_), .A3(new_n2213_), .ZN(new_n2214_));
  AOI21_X1   g2163(.A1(new_n2214_), .A2(new_n2118_), .B(new_n1044_), .ZN(new_n2215_));
  INV_X1     g2164(.I(new_n1044_), .ZN(new_n2216_));
  AOI21_X1   g2165(.A1(new_n2209_), .A2(new_n2212_), .B(new_n2213_), .ZN(new_n2217_));
  NOR3_X1    g2166(.A1(new_n2064_), .A2(new_n2080_), .A3(new_n2117_), .ZN(new_n2218_));
  NOR3_X1    g2167(.A1(new_n2217_), .A2(new_n2218_), .A3(new_n2216_), .ZN(new_n2219_));
  INV_X1     g2168(.I(new_n484_), .ZN(new_n2220_));
  NOR3_X1    g2169(.A1(new_n548_), .A2(new_n374_), .A3(new_n212_), .ZN(new_n2221_));
  INV_X1     g2170(.I(new_n2221_), .ZN(new_n2222_));
  NOR3_X1    g2171(.A1(new_n218_), .A2(new_n228_), .A3(new_n522_), .ZN(new_n2223_));
  INV_X1     g2172(.I(new_n2223_), .ZN(new_n2224_));
  NOR3_X1    g2173(.A1(new_n2224_), .A2(new_n2222_), .A3(new_n312_), .ZN(new_n2225_));
  INV_X1     g2174(.I(new_n2225_), .ZN(new_n2226_));
  NOR2_X1    g2175(.A1(new_n205_), .A2(new_n156_), .ZN(new_n2227_));
  NAND3_X1   g2176(.A1(new_n2227_), .A2(new_n465_), .A3(new_n675_), .ZN(new_n2228_));
  NOR2_X1    g2177(.A1(new_n151_), .A2(new_n245_), .ZN(new_n2229_));
  NOR4_X1    g2178(.A1(new_n733_), .A2(new_n64_), .A3(new_n171_), .A4(new_n322_), .ZN(new_n2230_));
  NOR2_X1    g2179(.A1(new_n821_), .A2(new_n156_), .ZN(new_n2231_));
  NAND4_X1   g2180(.A1(new_n672_), .A2(new_n2230_), .A3(new_n2231_), .A4(new_n2229_), .ZN(new_n2232_));
  NOR4_X1    g2181(.A1(new_n2226_), .A2(new_n2232_), .A3(new_n2220_), .A4(new_n2228_), .ZN(new_n2233_));
  INV_X1     g2182(.I(new_n2233_), .ZN(new_n2234_));
  NAND2_X1   g2183(.A1(new_n401_), .A2(new_n230_), .ZN(new_n2235_));
  NOR3_X1    g2184(.A1(new_n2234_), .A2(new_n399_), .A3(new_n2235_), .ZN(new_n2236_));
  INV_X1     g2185(.I(new_n786_), .ZN(new_n2237_));
  NOR2_X1    g2186(.A1(new_n1073_), .A2(new_n332_), .ZN(new_n2238_));
  INV_X1     g2187(.I(new_n2238_), .ZN(new_n2239_));
  NOR2_X1    g2188(.A1(new_n735_), .A2(new_n734_), .ZN(new_n2240_));
  NOR2_X1    g2189(.A1(new_n366_), .A2(new_n243_), .ZN(new_n2241_));
  NAND4_X1   g2190(.A1(new_n2241_), .A2(new_n325_), .A3(new_n413_), .A4(new_n2240_), .ZN(new_n2242_));
  NOR3_X1    g2191(.A1(new_n820_), .A2(new_n384_), .A3(new_n232_), .ZN(new_n2243_));
  INV_X1     g2192(.I(new_n2243_), .ZN(new_n2244_));
  NOR4_X1    g2193(.A1(new_n2239_), .A2(new_n2242_), .A3(new_n2244_), .A4(new_n2237_), .ZN(new_n2245_));
  NOR3_X1    g2194(.A1(new_n635_), .A2(new_n314_), .A3(new_n299_), .ZN(new_n2246_));
  NAND4_X1   g2195(.A1(new_n342_), .A2(new_n2246_), .A3(new_n192_), .A4(new_n277_), .ZN(new_n2247_));
  NOR2_X1    g2196(.A1(new_n256_), .A2(new_n251_), .ZN(new_n2248_));
  NAND4_X1   g2197(.A1(new_n231_), .A2(new_n2248_), .A3(new_n649_), .A4(new_n1246_), .ZN(new_n2249_));
  NOR3_X1    g2198(.A1(new_n539_), .A2(new_n219_), .A3(new_n375_), .ZN(new_n2250_));
  INV_X1     g2199(.I(new_n2250_), .ZN(new_n2251_));
  NAND4_X1   g2200(.A1(new_n401_), .A2(new_n220_), .A3(new_n375_), .A4(new_n420_), .ZN(new_n2252_));
  NOR4_X1    g2201(.A1(new_n2247_), .A2(new_n2249_), .A3(new_n2251_), .A4(new_n2252_), .ZN(new_n2253_));
  NAND3_X1   g2202(.A1(new_n2236_), .A2(new_n2245_), .A3(new_n2253_), .ZN(new_n2254_));
  NOR3_X1    g2203(.A1(new_n2215_), .A2(new_n2219_), .A3(new_n2254_), .ZN(new_n2255_));
  OAI21_X1   g2204(.A1(new_n2217_), .A2(new_n2218_), .B(new_n2216_), .ZN(new_n2256_));
  NAND3_X1   g2205(.A1(new_n2214_), .A2(new_n2118_), .A3(new_n1044_), .ZN(new_n2257_));
  INV_X1     g2206(.I(new_n2254_), .ZN(new_n2258_));
  AOI21_X1   g2207(.A1(new_n2256_), .A2(new_n2257_), .B(new_n2258_), .ZN(new_n2259_));
  NOR2_X1    g2208(.A1(new_n2255_), .A2(new_n2259_), .ZN(new_n2260_));
  OR2_X2     g2209(.A1(new_n1044_), .A2(new_n2073_), .Z(new_n2261_));
  NOR2_X1    g2210(.A1(new_n2070_), .A2(new_n2077_), .ZN(new_n2262_));
  INV_X1     g2211(.I(new_n2262_), .ZN(new_n2263_));
  XOR2_X1    g2212(.A1(new_n2070_), .A2(new_n2077_), .Z(new_n2264_));
  NAND3_X1   g2213(.A1(new_n2261_), .A2(new_n2263_), .A3(new_n2264_), .ZN(new_n2265_));
  XNOR2_X1   g2214(.A1(new_n2070_), .A2(new_n2077_), .ZN(new_n2266_));
  OAI21_X1   g2215(.A1(new_n2074_), .A2(new_n2266_), .B(new_n2262_), .ZN(new_n2267_));
  NAND2_X1   g2216(.A1(new_n2265_), .A2(new_n2267_), .ZN(new_n2268_));
  NAND2_X1   g2217(.A1(new_n2064_), .A2(new_n2268_), .ZN(new_n2269_));
  INV_X1     g2218(.I(new_n2268_), .ZN(new_n2270_));
  NAND2_X1   g2219(.A1(new_n2270_), .A2(new_n2209_), .ZN(new_n2271_));
  NOR3_X1    g2220(.A1(new_n994_), .A2(new_n307_), .A3(new_n347_), .ZN(new_n2272_));
  INV_X1     g2221(.I(new_n2272_), .ZN(new_n2273_));
  NOR2_X1    g2222(.A1(new_n205_), .A2(new_n331_), .ZN(new_n2274_));
  NAND3_X1   g2223(.A1(new_n679_), .A2(new_n2274_), .A3(new_n1235_), .ZN(new_n2275_));
  NOR2_X1    g2224(.A1(new_n339_), .A2(new_n221_), .ZN(new_n2276_));
  NAND4_X1   g2225(.A1(new_n2276_), .A2(new_n654_), .A3(new_n319_), .A4(new_n384_), .ZN(new_n2277_));
  NOR3_X1    g2226(.A1(new_n2275_), .A2(new_n793_), .A3(new_n2277_), .ZN(new_n2278_));
  INV_X1     g2227(.I(new_n2278_), .ZN(new_n2279_));
  NAND4_X1   g2228(.A1(new_n514_), .A2(new_n821_), .A3(new_n292_), .A4(new_n363_), .ZN(new_n2280_));
  NAND4_X1   g2229(.A1(new_n380_), .A2(new_n197_), .A3(new_n313_), .A4(new_n447_), .ZN(new_n2281_));
  NOR2_X1    g2230(.A1(new_n2281_), .A2(new_n2280_), .ZN(new_n2282_));
  NOR2_X1    g2231(.A1(new_n510_), .A2(new_n1101_), .ZN(new_n2283_));
  NAND4_X1   g2232(.A1(new_n2283_), .A2(new_n201_), .A3(new_n222_), .A4(new_n317_), .ZN(new_n2284_));
  INV_X1     g2233(.I(new_n2284_), .ZN(new_n2285_));
  NAND2_X1   g2234(.A1(new_n310_), .A2(new_n847_), .ZN(new_n2286_));
  NAND4_X1   g2235(.A1(new_n228_), .A2(new_n363_), .A3(new_n374_), .A4(new_n921_), .ZN(new_n2287_));
  NOR4_X1    g2236(.A1(new_n2287_), .A2(new_n207_), .A3(new_n2286_), .A4(new_n892_), .ZN(new_n2288_));
  NAND3_X1   g2237(.A1(new_n2285_), .A2(new_n2282_), .A3(new_n2288_), .ZN(new_n2289_));
  NOR3_X1    g2238(.A1(new_n2273_), .A2(new_n2279_), .A3(new_n2289_), .ZN(new_n2290_));
  INV_X1     g2239(.I(new_n2290_), .ZN(new_n2291_));
  NAND3_X1   g2240(.A1(new_n2271_), .A2(new_n2269_), .A3(new_n2291_), .ZN(new_n2292_));
  NOR2_X1    g2241(.A1(new_n2193_), .A2(new_n2027_), .ZN(new_n2293_));
  AOI21_X1   g2242(.A1(new_n1953_), .A2(new_n1956_), .B(new_n2202_), .ZN(new_n2294_));
  NOR3_X1    g2243(.A1(new_n2027_), .A2(new_n2191_), .A3(new_n2192_), .ZN(new_n2295_));
  NOR2_X1    g2244(.A1(new_n2294_), .A2(new_n2295_), .ZN(new_n2296_));
  NOR3_X1    g2245(.A1(new_n2296_), .A2(new_n2200_), .A3(new_n2293_), .ZN(new_n2297_));
  NAND2_X1   g2246(.A1(new_n1957_), .A2(new_n2202_), .ZN(new_n2298_));
  OAI21_X1   g2247(.A1(new_n2191_), .A2(new_n2192_), .B(new_n2027_), .ZN(new_n2299_));
  NAND3_X1   g2248(.A1(new_n2202_), .A2(new_n1956_), .A3(new_n1953_), .ZN(new_n2300_));
  NAND2_X1   g2249(.A1(new_n2299_), .A2(new_n2300_), .ZN(new_n2301_));
  AOI21_X1   g2250(.A1(new_n2301_), .A2(new_n2021_), .B(new_n2298_), .ZN(new_n2302_));
  NOR2_X1    g2251(.A1(new_n2302_), .A2(new_n2297_), .ZN(new_n2303_));
  NOR2_X1    g2252(.A1(new_n1872_), .A2(new_n2303_), .ZN(new_n2304_));
  NAND3_X1   g2253(.A1(new_n2301_), .A2(new_n2021_), .A3(new_n2298_), .ZN(new_n2305_));
  OAI21_X1   g2254(.A1(new_n2296_), .A2(new_n2200_), .B(new_n2293_), .ZN(new_n2306_));
  NAND2_X1   g2255(.A1(new_n2306_), .A2(new_n2305_), .ZN(new_n2307_));
  NOR2_X1    g2256(.A1(new_n2190_), .A2(new_n2307_), .ZN(new_n2308_));
  NOR2_X1    g2257(.A1(new_n2308_), .A2(new_n2304_), .ZN(new_n2309_));
  NAND3_X1   g2258(.A1(new_n388_), .A2(new_n292_), .A3(new_n376_), .ZN(new_n2310_));
  NOR3_X1    g2259(.A1(new_n207_), .A2(new_n391_), .A3(new_n243_), .ZN(new_n2311_));
  INV_X1     g2260(.I(new_n2311_), .ZN(new_n2312_));
  NOR4_X1    g2261(.A1(new_n198_), .A2(new_n2312_), .A3(new_n448_), .A4(new_n2310_), .ZN(new_n2313_));
  AND4_X2    g2262(.A1(new_n413_), .A2(new_n2313_), .A3(new_n307_), .A4(new_n546_), .Z(new_n2314_));
  NOR4_X1    g2263(.A1(new_n366_), .A2(new_n132_), .A3(new_n222_), .A4(new_n456_), .ZN(new_n2315_));
  NAND3_X1   g2264(.A1(new_n2315_), .A2(new_n313_), .A3(new_n254_), .ZN(new_n2316_));
  NAND3_X1   g2265(.A1(new_n739_), .A2(new_n388_), .A3(new_n649_), .ZN(new_n2317_));
  INV_X1     g2266(.I(new_n359_), .ZN(new_n2318_));
  NOR2_X1    g2267(.A1(new_n2318_), .A2(new_n398_), .ZN(new_n2319_));
  NAND4_X1   g2268(.A1(new_n2319_), .A2(new_n1094_), .A3(new_n523_), .A4(new_n218_), .ZN(new_n2320_));
  NAND3_X1   g2269(.A1(new_n1226_), .A2(new_n1137_), .A3(new_n791_), .ZN(new_n2321_));
  NOR4_X1    g2270(.A1(new_n2320_), .A2(new_n2316_), .A3(new_n2321_), .A4(new_n2317_), .ZN(new_n2322_));
  NAND3_X1   g2271(.A1(new_n2314_), .A2(new_n613_), .A3(new_n2322_), .ZN(new_n2323_));
  INV_X1     g2272(.I(new_n2056_), .ZN(new_n2324_));
  NOR3_X1    g2273(.A1(new_n2033_), .A2(new_n2038_), .A3(new_n2040_), .ZN(new_n2325_));
  OAI21_X1   g2274(.A1(new_n2076_), .A2(new_n2325_), .B(new_n2048_), .ZN(new_n2326_));
  NOR3_X1    g2275(.A1(new_n2033_), .A2(new_n2038_), .A3(new_n2039_), .ZN(new_n2327_));
  AOI21_X1   g2276(.A1(new_n2043_), .A2(new_n2045_), .B(new_n2040_), .ZN(new_n2328_));
  OAI21_X1   g2277(.A1(new_n2328_), .A2(new_n2327_), .B(new_n2031_), .ZN(new_n2329_));
  NAND3_X1   g2278(.A1(new_n2326_), .A2(new_n2329_), .A3(new_n2060_), .ZN(new_n2330_));
  INV_X1     g2279(.I(new_n2060_), .ZN(new_n2331_));
  OAI21_X1   g2280(.A1(new_n2047_), .A2(new_n2051_), .B(new_n2331_), .ZN(new_n2332_));
  NOR4_X1    g2281(.A1(new_n653_), .A2(new_n317_), .A3(new_n1069_), .A4(new_n341_), .ZN(new_n2333_));
  INV_X1     g2282(.I(new_n2274_), .ZN(new_n2334_));
  NOR3_X1    g2283(.A1(new_n2334_), .A2(new_n671_), .A3(new_n332_), .ZN(new_n2335_));
  NAND4_X1   g2284(.A1(new_n2335_), .A2(new_n484_), .A3(new_n919_), .A4(new_n2333_), .ZN(new_n2336_));
  NOR3_X1    g2285(.A1(new_n2336_), .A2(new_n461_), .A3(new_n332_), .ZN(new_n2337_));
  INV_X1     g2286(.I(new_n2337_), .ZN(new_n2338_));
  NOR2_X1    g2287(.A1(new_n992_), .A2(new_n990_), .ZN(new_n2339_));
  NOR2_X1    g2288(.A1(new_n820_), .A2(new_n891_), .ZN(new_n2340_));
  NAND2_X1   g2289(.A1(new_n1224_), .A2(new_n424_), .ZN(new_n2341_));
  NOR4_X1    g2290(.A1(new_n2341_), .A2(new_n401_), .A3(new_n608_), .A4(new_n282_), .ZN(new_n2342_));
  NOR3_X1    g2291(.A1(new_n218_), .A2(new_n649_), .A3(new_n847_), .ZN(new_n2343_));
  NAND4_X1   g2292(.A1(new_n2342_), .A2(new_n2339_), .A3(new_n2340_), .A4(new_n2343_), .ZN(new_n2344_));
  INV_X1     g2293(.I(new_n540_), .ZN(new_n2345_));
  NOR2_X1    g2294(.A1(new_n160_), .A2(new_n243_), .ZN(new_n2346_));
  INV_X1     g2295(.I(new_n2346_), .ZN(new_n2347_));
  NOR4_X1    g2296(.A1(new_n2347_), .A2(new_n2345_), .A3(new_n449_), .A4(new_n655_), .ZN(new_n2348_));
  NOR4_X1    g2297(.A1(new_n385_), .A2(new_n151_), .A3(new_n227_), .A4(new_n245_), .ZN(new_n2349_));
  NOR4_X1    g2298(.A1(new_n400_), .A2(new_n733_), .A3(new_n668_), .A4(new_n339_), .ZN(new_n2350_));
  NAND3_X1   g2299(.A1(new_n2348_), .A2(new_n2349_), .A3(new_n2350_), .ZN(new_n2351_));
  NOR3_X1    g2300(.A1(new_n2338_), .A2(new_n2344_), .A3(new_n2351_), .ZN(new_n2352_));
  INV_X1     g2301(.I(new_n2352_), .ZN(new_n2353_));
  AOI21_X1   g2302(.A1(new_n2332_), .A2(new_n2330_), .B(new_n2353_), .ZN(new_n2354_));
  OAI21_X1   g2303(.A1(new_n2190_), .A2(new_n2204_), .B(new_n2354_), .ZN(new_n2355_));
  NOR3_X1    g2304(.A1(new_n2047_), .A2(new_n2051_), .A3(new_n2331_), .ZN(new_n2356_));
  AOI21_X1   g2305(.A1(new_n2326_), .A2(new_n2329_), .B(new_n2060_), .ZN(new_n2357_));
  OAI21_X1   g2306(.A1(new_n2357_), .A2(new_n2356_), .B(new_n2352_), .ZN(new_n2358_));
  NAND3_X1   g2307(.A1(new_n1872_), .A2(new_n2029_), .A3(new_n2358_), .ZN(new_n2359_));
  AOI21_X1   g2308(.A1(new_n2355_), .A2(new_n2359_), .B(new_n2324_), .ZN(new_n2360_));
  AOI21_X1   g2309(.A1(new_n1872_), .A2(new_n2029_), .B(new_n2358_), .ZN(new_n2361_));
  NOR3_X1    g2310(.A1(new_n2190_), .A2(new_n2204_), .A3(new_n2354_), .ZN(new_n2362_));
  NOR3_X1    g2311(.A1(new_n2362_), .A2(new_n2361_), .A3(new_n2056_), .ZN(new_n2363_));
  NOR2_X1    g2312(.A1(new_n2363_), .A2(new_n2360_), .ZN(new_n2364_));
  OAI21_X1   g2313(.A1(new_n2364_), .A2(new_n2323_), .B(new_n2309_), .ZN(new_n2365_));
  NOR2_X1    g2314(.A1(new_n1796_), .A2(new_n1853_), .ZN(new_n2366_));
  NOR3_X1    g2315(.A1(new_n1788_), .A2(new_n1785_), .A3(new_n1789_), .ZN(new_n2367_));
  AOI21_X1   g2316(.A1(new_n1773_), .A2(new_n1776_), .B(new_n1781_), .ZN(new_n2368_));
  OAI21_X1   g2317(.A1(new_n2368_), .A2(new_n2367_), .B(new_n1792_), .ZN(new_n2369_));
  NOR3_X1    g2318(.A1(new_n1788_), .A2(new_n1785_), .A3(new_n1781_), .ZN(new_n2370_));
  OAI21_X1   g2319(.A1(new_n1797_), .A2(new_n2370_), .B(new_n1738_), .ZN(new_n2371_));
  NAND3_X1   g2320(.A1(new_n2185_), .A2(new_n2371_), .A3(new_n2369_), .ZN(new_n2372_));
  OAI21_X1   g2321(.A1(new_n1791_), .A2(new_n1795_), .B(new_n1853_), .ZN(new_n2373_));
  NAND2_X1   g2322(.A1(new_n2373_), .A2(new_n2372_), .ZN(new_n2374_));
  OAI21_X1   g2323(.A1(new_n1855_), .A2(new_n1856_), .B(new_n2374_), .ZN(new_n2375_));
  NOR2_X1    g2324(.A1(new_n2375_), .A2(new_n2366_), .ZN(new_n2376_));
  NAND2_X1   g2325(.A1(new_n1843_), .A2(new_n1839_), .ZN(new_n2377_));
  INV_X1     g2326(.I(new_n2366_), .ZN(new_n2378_));
  AOI21_X1   g2327(.A1(new_n2377_), .A2(new_n2374_), .B(new_n2378_), .ZN(new_n2379_));
  OAI21_X1   g2328(.A1(new_n2376_), .A2(new_n2379_), .B(new_n2181_), .ZN(new_n2380_));
  NAND3_X1   g2329(.A1(new_n2377_), .A2(new_n2378_), .A3(new_n2374_), .ZN(new_n2381_));
  NAND2_X1   g2330(.A1(new_n2375_), .A2(new_n2366_), .ZN(new_n2382_));
  NAND3_X1   g2331(.A1(new_n2381_), .A2(new_n2382_), .A3(new_n1736_), .ZN(new_n2383_));
  INV_X1     g2332(.I(new_n2228_), .ZN(new_n2384_));
  NOR3_X1    g2333(.A1(new_n233_), .A2(new_n421_), .A3(new_n420_), .ZN(new_n2385_));
  INV_X1     g2334(.I(new_n2385_), .ZN(new_n2386_));
  NOR3_X1    g2335(.A1(new_n2386_), .A2(new_n400_), .A3(new_n848_), .ZN(new_n2387_));
  NOR3_X1    g2336(.A1(new_n453_), .A2(new_n425_), .A3(new_n619_), .ZN(new_n2388_));
  NAND2_X1   g2337(.A1(new_n221_), .A2(new_n222_), .ZN(new_n2389_));
  NOR4_X1    g2338(.A1(new_n2389_), .A2(new_n240_), .A3(new_n310_), .A4(new_n292_), .ZN(new_n2390_));
  NAND4_X1   g2339(.A1(new_n2384_), .A2(new_n2387_), .A3(new_n2388_), .A4(new_n2390_), .ZN(new_n2391_));
  INV_X1     g2340(.I(new_n2391_), .ZN(new_n2392_));
  NOR2_X1    g2341(.A1(new_n151_), .A2(new_n608_), .ZN(new_n2393_));
  INV_X1     g2342(.I(new_n2393_), .ZN(new_n2394_));
  NOR2_X1    g2343(.A1(new_n2394_), .A2(new_n444_), .ZN(new_n2395_));
  NAND3_X1   g2344(.A1(new_n2395_), .A2(new_n596_), .A3(new_n652_), .ZN(new_n2396_));
  INV_X1     g2345(.I(new_n414_), .ZN(new_n2397_));
  NOR4_X1    g2346(.A1(new_n110_), .A2(new_n201_), .A3(new_n292_), .A4(new_n345_), .ZN(new_n2398_));
  NAND3_X1   g2347(.A1(new_n2397_), .A2(new_n452_), .A3(new_n2398_), .ZN(new_n2399_));
  NOR4_X1    g2348(.A1(new_n2396_), .A2(new_n840_), .A3(new_n989_), .A4(new_n2399_), .ZN(new_n2400_));
  AND3_X2    g2349(.A1(new_n2314_), .A2(new_n2392_), .A3(new_n2400_), .Z(new_n2401_));
  NAND3_X1   g2350(.A1(new_n2380_), .A2(new_n2383_), .A3(new_n2401_), .ZN(new_n2402_));
  NAND2_X1   g2351(.A1(new_n256_), .A2(new_n209_), .ZN(new_n2403_));
  NOR4_X1    g2352(.A1(new_n2403_), .A2(new_n602_), .A3(new_n332_), .A4(new_n515_), .ZN(new_n2404_));
  NAND3_X1   g2353(.A1(new_n401_), .A2(new_n201_), .A3(new_n475_), .ZN(new_n2405_));
  NOR4_X1    g2354(.A1(new_n2405_), .A2(new_n921_), .A3(new_n257_), .A4(new_n452_), .ZN(new_n2406_));
  NAND2_X1   g2355(.A1(new_n230_), .A2(new_n243_), .ZN(new_n2407_));
  NOR4_X1    g2356(.A1(new_n2407_), .A2(new_n285_), .A3(new_n375_), .A4(new_n319_), .ZN(new_n2408_));
  NAND3_X1   g2357(.A1(new_n2406_), .A2(new_n2408_), .A3(new_n2404_), .ZN(new_n2409_));
  INV_X1     g2358(.I(new_n2409_), .ZN(new_n2410_));
  INV_X1     g2359(.I(new_n765_), .ZN(new_n2411_));
  NOR3_X1    g2360(.A1(new_n201_), .A2(new_n338_), .A3(new_n367_), .ZN(new_n2412_));
  INV_X1     g2361(.I(new_n2412_), .ZN(new_n2413_));
  NOR2_X1    g2362(.A1(new_n997_), .A2(new_n625_), .ZN(new_n2414_));
  INV_X1     g2363(.I(new_n2414_), .ZN(new_n2415_));
  NOR4_X1    g2364(.A1(new_n2415_), .A2(new_n405_), .A3(new_n2411_), .A4(new_n2413_), .ZN(new_n2416_));
  INV_X1     g2365(.I(new_n665_), .ZN(new_n2417_));
  NOR2_X1    g2366(.A1(new_n241_), .A2(new_n221_), .ZN(new_n2418_));
  NOR2_X1    g2367(.A1(new_n230_), .A2(new_n847_), .ZN(new_n2419_));
  NAND4_X1   g2368(.A1(new_n535_), .A2(new_n2418_), .A3(new_n2419_), .A4(new_n313_), .ZN(new_n2420_));
  NAND4_X1   g2369(.A1(new_n514_), .A2(new_n388_), .A3(new_n363_), .A4(new_n212_), .ZN(new_n2421_));
  NOR4_X1    g2370(.A1(new_n2420_), .A2(new_n2421_), .A3(new_n2417_), .A4(new_n355_), .ZN(new_n2422_));
  NAND3_X1   g2371(.A1(new_n2410_), .A2(new_n2416_), .A3(new_n2422_), .ZN(new_n2423_));
  NOR2_X1    g2372(.A1(new_n2402_), .A2(new_n2423_), .ZN(new_n2424_));
  OAI21_X1   g2373(.A1(new_n1336_), .A2(new_n1333_), .B(new_n1868_), .ZN(new_n2425_));
  AOI21_X1   g2374(.A1(new_n1861_), .A2(new_n1736_), .B(new_n2425_), .ZN(new_n2426_));
  NOR2_X1    g2375(.A1(new_n2186_), .A2(new_n2185_), .ZN(new_n2427_));
  INV_X1     g2376(.I(new_n2425_), .ZN(new_n2428_));
  NOR4_X1    g2377(.A1(new_n2181_), .A2(new_n2427_), .A3(new_n1860_), .A4(new_n2428_), .ZN(new_n2429_));
  OAI21_X1   g2378(.A1(new_n2426_), .A2(new_n2429_), .B(new_n1864_), .ZN(new_n2430_));
  OAI21_X1   g2379(.A1(new_n2187_), .A2(new_n2181_), .B(new_n2428_), .ZN(new_n2431_));
  NAND4_X1   g2380(.A1(new_n1858_), .A2(new_n1736_), .A3(new_n1844_), .A4(new_n2425_), .ZN(new_n2432_));
  NAND3_X1   g2381(.A1(new_n2431_), .A2(new_n2432_), .A3(new_n1863_), .ZN(new_n2433_));
  AOI22_X1   g2382(.A1(new_n2430_), .A2(new_n2433_), .B1(new_n2402_), .B2(new_n2423_), .ZN(new_n2434_));
  NAND3_X1   g2383(.A1(new_n462_), .A2(new_n467_), .A3(new_n464_), .ZN(new_n2435_));
  INV_X1     g2384(.I(new_n2435_), .ZN(new_n2436_));
  NOR2_X1    g2385(.A1(new_n277_), .A2(new_n649_), .ZN(new_n2437_));
  INV_X1     g2386(.I(new_n2437_), .ZN(new_n2438_));
  NOR3_X1    g2387(.A1(new_n2438_), .A2(new_n465_), .A3(new_n2394_), .ZN(new_n2439_));
  INV_X1     g2388(.I(new_n2419_), .ZN(new_n2440_));
  NOR3_X1    g2389(.A1(new_n151_), .A2(new_n589_), .A3(new_n367_), .ZN(new_n2441_));
  INV_X1     g2390(.I(new_n2441_), .ZN(new_n2442_));
  NOR4_X1    g2391(.A1(new_n2442_), .A2(new_n2440_), .A3(new_n341_), .A4(new_n774_), .ZN(new_n2443_));
  NOR4_X1    g2392(.A1(new_n516_), .A2(new_n205_), .A3(new_n319_), .A4(new_n548_), .ZN(new_n2444_));
  NOR3_X1    g2393(.A1(new_n2244_), .A2(new_n653_), .A3(new_n857_), .ZN(new_n2445_));
  NAND4_X1   g2394(.A1(new_n2443_), .A2(new_n2445_), .A3(new_n2439_), .A4(new_n2444_), .ZN(new_n2446_));
  INV_X1     g2395(.I(new_n2446_), .ZN(new_n2447_));
  NAND2_X1   g2396(.A1(new_n736_), .A2(new_n732_), .ZN(new_n2448_));
  INV_X1     g2397(.I(new_n2448_), .ZN(new_n2449_));
  NOR3_X1    g2398(.A1(new_n388_), .A2(new_n468_), .A3(new_n221_), .ZN(new_n2450_));
  NOR2_X1    g2399(.A1(new_n277_), .A2(new_n304_), .ZN(new_n2451_));
  NAND4_X1   g2400(.A1(new_n2449_), .A2(new_n786_), .A3(new_n2450_), .A4(new_n2451_), .ZN(new_n2452_));
  NAND4_X1   g2401(.A1(new_n357_), .A2(new_n231_), .A3(new_n205_), .A4(new_n413_), .ZN(new_n2453_));
  NOR4_X1    g2402(.A1(new_n2452_), .A2(new_n762_), .A3(new_n2320_), .A4(new_n2453_), .ZN(new_n2454_));
  NAND3_X1   g2403(.A1(new_n2447_), .A2(new_n2436_), .A3(new_n2454_), .ZN(new_n2455_));
  INV_X1     g2404(.I(new_n2455_), .ZN(new_n2456_));
  OAI21_X1   g2405(.A1(new_n2434_), .A2(new_n2424_), .B(new_n2456_), .ZN(new_n2457_));
  NAND2_X1   g2406(.A1(new_n2193_), .A2(new_n2027_), .ZN(new_n2458_));
  NAND2_X1   g2407(.A1(new_n2458_), .A2(new_n2298_), .ZN(new_n2459_));
  NAND2_X1   g2408(.A1(new_n1872_), .A2(new_n2459_), .ZN(new_n2460_));
  OAI21_X1   g2409(.A1(new_n1872_), .A2(new_n2296_), .B(new_n2460_), .ZN(new_n2461_));
  AOI21_X1   g2410(.A1(new_n2382_), .A2(new_n2381_), .B(new_n1736_), .ZN(new_n2462_));
  NOR3_X1    g2411(.A1(new_n2181_), .A2(new_n2376_), .A3(new_n2379_), .ZN(new_n2463_));
  INV_X1     g2412(.I(new_n2401_), .ZN(new_n2464_));
  NOR3_X1    g2413(.A1(new_n2463_), .A2(new_n2462_), .A3(new_n2464_), .ZN(new_n2465_));
  INV_X1     g2414(.I(new_n2423_), .ZN(new_n2466_));
  NAND2_X1   g2415(.A1(new_n2465_), .A2(new_n2466_), .ZN(new_n2467_));
  AOI21_X1   g2416(.A1(new_n2431_), .A2(new_n2432_), .B(new_n1863_), .ZN(new_n2468_));
  NOR3_X1    g2417(.A1(new_n2426_), .A2(new_n2429_), .A3(new_n1864_), .ZN(new_n2469_));
  OAI22_X1   g2418(.A1(new_n2469_), .A2(new_n2468_), .B1(new_n2465_), .B2(new_n2466_), .ZN(new_n2470_));
  NAND3_X1   g2419(.A1(new_n2470_), .A2(new_n2467_), .A3(new_n2455_), .ZN(new_n2471_));
  NAND2_X1   g2420(.A1(new_n2471_), .A2(new_n2461_), .ZN(new_n2472_));
  NAND2_X1   g2421(.A1(new_n2472_), .A2(new_n2457_), .ZN(new_n2473_));
  OAI21_X1   g2422(.A1(new_n2362_), .A2(new_n2361_), .B(new_n2056_), .ZN(new_n2474_));
  NAND3_X1   g2423(.A1(new_n2355_), .A2(new_n2359_), .A3(new_n2324_), .ZN(new_n2475_));
  NAND3_X1   g2424(.A1(new_n2474_), .A2(new_n2475_), .A3(new_n2323_), .ZN(new_n2476_));
  OAI21_X1   g2425(.A1(new_n2063_), .A2(new_n2053_), .B(new_n2264_), .ZN(new_n2477_));
  NAND2_X1   g2426(.A1(new_n2070_), .A2(new_n2077_), .ZN(new_n2478_));
  NAND2_X1   g2427(.A1(new_n2263_), .A2(new_n2478_), .ZN(new_n2479_));
  NAND3_X1   g2428(.A1(new_n2208_), .A2(new_n2207_), .A3(new_n2479_), .ZN(new_n2480_));
  NAND2_X1   g2429(.A1(new_n2480_), .A2(new_n2477_), .ZN(new_n2481_));
  NAND4_X1   g2430(.A1(new_n2365_), .A2(new_n2473_), .A3(new_n2481_), .A4(new_n2476_), .ZN(new_n2482_));
  NAND2_X1   g2431(.A1(new_n2190_), .A2(new_n2307_), .ZN(new_n2483_));
  NAND2_X1   g2432(.A1(new_n1872_), .A2(new_n2303_), .ZN(new_n2484_));
  NAND2_X1   g2433(.A1(new_n2483_), .A2(new_n2484_), .ZN(new_n2485_));
  INV_X1     g2434(.I(new_n2323_), .ZN(new_n2486_));
  NAND2_X1   g2435(.A1(new_n2474_), .A2(new_n2475_), .ZN(new_n2487_));
  AOI21_X1   g2436(.A1(new_n2487_), .A2(new_n2486_), .B(new_n2485_), .ZN(new_n2488_));
  AOI21_X1   g2437(.A1(new_n2470_), .A2(new_n2467_), .B(new_n2455_), .ZN(new_n2489_));
  AOI21_X1   g2438(.A1(new_n2461_), .A2(new_n2471_), .B(new_n2489_), .ZN(new_n2490_));
  INV_X1     g2439(.I(new_n2476_), .ZN(new_n2491_));
  NOR3_X1    g2440(.A1(new_n2488_), .A2(new_n2491_), .A3(new_n2490_), .ZN(new_n2492_));
  XOR2_X1    g2441(.A1(new_n2358_), .A2(new_n2324_), .Z(new_n2493_));
  NOR2_X1    g2442(.A1(new_n2493_), .A2(new_n2030_), .ZN(new_n2494_));
  INV_X1     g2443(.I(new_n2494_), .ZN(new_n2495_));
  INV_X1     g2444(.I(new_n2416_), .ZN(new_n2496_));
  NAND4_X1   g2445(.A1(new_n2444_), .A2(new_n842_), .A3(new_n846_), .A4(new_n731_), .ZN(new_n2497_));
  NAND2_X1   g2446(.A1(new_n2318_), .A2(new_n421_), .ZN(new_n2498_));
  NOR4_X1    g2447(.A1(new_n2498_), .A2(new_n660_), .A3(new_n168_), .A4(new_n826_), .ZN(new_n2499_));
  NOR3_X1    g2448(.A1(new_n347_), .A2(new_n388_), .A3(new_n233_), .ZN(new_n2500_));
  NAND2_X1   g2449(.A1(new_n2500_), .A2(new_n739_), .ZN(new_n2501_));
  INV_X1     g2450(.I(new_n2501_), .ZN(new_n2502_));
  NAND2_X1   g2451(.A1(new_n622_), .A2(new_n160_), .ZN(new_n2503_));
  NOR2_X1    g2452(.A1(new_n310_), .A2(new_n197_), .ZN(new_n2504_));
  INV_X1     g2453(.I(new_n2504_), .ZN(new_n2505_));
  NOR4_X1    g2454(.A1(new_n2505_), .A2(new_n246_), .A3(new_n2503_), .A4(new_n301_), .ZN(new_n2506_));
  NAND4_X1   g2455(.A1(new_n2506_), .A2(new_n2502_), .A3(new_n2499_), .A4(new_n1002_), .ZN(new_n2507_));
  NOR3_X1    g2456(.A1(new_n2496_), .A2(new_n2507_), .A3(new_n2497_), .ZN(new_n2508_));
  INV_X1     g2457(.I(new_n2508_), .ZN(new_n2509_));
  NOR2_X1    g2458(.A1(new_n2495_), .A2(new_n2509_), .ZN(new_n2510_));
  OAI21_X1   g2459(.A1(new_n2492_), .A2(new_n2481_), .B(new_n2510_), .ZN(new_n2511_));
  NOR2_X1    g2460(.A1(new_n2270_), .A2(new_n2209_), .ZN(new_n2512_));
  NOR2_X1    g2461(.A1(new_n2064_), .A2(new_n2268_), .ZN(new_n2513_));
  NOR3_X1    g2462(.A1(new_n2512_), .A2(new_n2513_), .A3(new_n2290_), .ZN(new_n2514_));
  AOI21_X1   g2463(.A1(new_n2271_), .A2(new_n2269_), .B(new_n2291_), .ZN(new_n2515_));
  NOR2_X1    g2464(.A1(new_n2514_), .A2(new_n2515_), .ZN(new_n2516_));
  NAND3_X1   g2465(.A1(new_n2511_), .A2(new_n2516_), .A3(new_n2482_), .ZN(new_n2517_));
  AOI21_X1   g2466(.A1(new_n2517_), .A2(new_n2292_), .B(new_n2260_), .ZN(new_n2518_));
  NAND2_X1   g2467(.A1(new_n2209_), .A2(new_n2212_), .ZN(new_n2519_));
  AOI21_X1   g2468(.A1(new_n2084_), .A2(new_n2116_), .B(new_n2216_), .ZN(new_n2520_));
  INV_X1     g2469(.I(new_n2520_), .ZN(new_n2521_));
  OAI21_X1   g2470(.A1(new_n2519_), .A2(new_n2521_), .B(new_n2213_), .ZN(new_n2522_));
  NAND2_X1   g2471(.A1(new_n2112_), .A2(new_n2085_), .ZN(new_n2523_));
  NAND2_X1   g2472(.A1(new_n2523_), .A2(new_n2114_), .ZN(new_n2524_));
  INV_X1     g2473(.I(new_n2524_), .ZN(new_n2525_));
  OAI21_X1   g2474(.A1(new_n2089_), .A2(new_n2101_), .B(new_n2102_), .ZN(new_n2526_));
  NAND2_X1   g2475(.A1(new_n567_), .A2(new_n708_), .ZN(new_n2527_));
  OAI21_X1   g2476(.A1(new_n572_), .A2(new_n708_), .B(new_n2527_), .ZN(new_n2528_));
  NAND3_X1   g2477(.A1(new_n2528_), .A2(new_n565_), .A3(new_n875_), .ZN(new_n2529_));
  NAND3_X1   g2478(.A1(new_n2528_), .A2(new_n580_), .A3(new_n645_), .ZN(new_n2530_));
  NAND2_X1   g2479(.A1(new_n2529_), .A2(new_n2530_), .ZN(new_n2531_));
  NAND2_X1   g2480(.A1(new_n2531_), .A2(new_n562_), .ZN(new_n2532_));
  INV_X1     g2481(.I(new_n2532_), .ZN(new_n2533_));
  XOR2_X1    g2482(.A1(new_n687_), .A2(new_n587_), .Z(new_n2534_));
  OR2_X2     g2483(.A1(new_n2534_), .A2(new_n550_), .Z(new_n2535_));
  NAND2_X1   g2484(.A1(new_n2535_), .A2(new_n438_), .ZN(new_n2536_));
  NOR2_X1    g2485(.A1(new_n2535_), .A2(new_n438_), .ZN(new_n2537_));
  NAND2_X1   g2486(.A1(new_n2534_), .A2(new_n1745_), .ZN(new_n2538_));
  NOR2_X1    g2487(.A1(new_n2537_), .A2(new_n2538_), .ZN(new_n2539_));
  NAND2_X1   g2488(.A1(new_n2539_), .A2(new_n2536_), .ZN(new_n2540_));
  NOR2_X1    g2489(.A1(new_n266_), .A2(new_n702_), .ZN(new_n2541_));
  AND2_X2    g2490(.A1(new_n2540_), .A2(new_n2541_), .Z(new_n2542_));
  NOR2_X1    g2491(.A1(new_n2540_), .A2(new_n2541_), .ZN(new_n2543_));
  OAI21_X1   g2492(.A1(new_n2542_), .A2(new_n2543_), .B(new_n2533_), .ZN(new_n2544_));
  XNOR2_X1   g2493(.A1(new_n2540_), .A2(new_n2541_), .ZN(new_n2545_));
  OAI21_X1   g2494(.A1(new_n2533_), .A2(new_n2545_), .B(new_n2544_), .ZN(new_n2546_));
  AOI21_X1   g2495(.A1(new_n266_), .A2(new_n271_), .B(new_n577_), .ZN(new_n2547_));
  NOR3_X1    g2496(.A1(new_n1178_), .A2(new_n2547_), .A3(new_n272_), .ZN(new_n2548_));
  INV_X1     g2497(.I(new_n2548_), .ZN(new_n2549_));
  NOR2_X1    g2498(.A1(new_n2546_), .A2(new_n2549_), .ZN(new_n2550_));
  NAND2_X1   g2499(.A1(new_n2546_), .A2(new_n2549_), .ZN(new_n2551_));
  INV_X1     g2500(.I(new_n2551_), .ZN(new_n2552_));
  OAI21_X1   g2501(.A1(new_n2552_), .A2(new_n2550_), .B(new_n2526_), .ZN(new_n2553_));
  INV_X1     g2502(.I(new_n2526_), .ZN(new_n2554_));
  XOR2_X1    g2503(.A1(new_n2546_), .A2(new_n2549_), .Z(new_n2555_));
  NAND2_X1   g2504(.A1(new_n2555_), .A2(new_n2554_), .ZN(new_n2556_));
  NAND2_X1   g2505(.A1(new_n2556_), .A2(new_n2553_), .ZN(new_n2557_));
  XOR2_X1    g2506(.A1(new_n2557_), .A2(new_n2525_), .Z(new_n2558_));
  INV_X1     g2507(.I(new_n2558_), .ZN(new_n2559_));
  NAND2_X1   g2508(.A1(new_n2522_), .A2(new_n2559_), .ZN(new_n2560_));
  XOR2_X1    g2509(.A1(new_n2557_), .A2(new_n2524_), .Z(new_n2561_));
  OAI21_X1   g2510(.A1(new_n2522_), .A2(new_n2561_), .B(new_n2560_), .ZN(new_n2562_));
  NAND2_X1   g2511(.A1(new_n2518_), .A2(new_n2562_), .ZN(new_n2563_));
  NOR2_X1    g2512(.A1(new_n2215_), .A2(new_n2219_), .ZN(new_n2564_));
  NAND2_X1   g2513(.A1(new_n2564_), .A2(new_n2254_), .ZN(new_n2565_));
  NOR2_X1    g2514(.A1(new_n257_), .A2(new_n151_), .ZN(new_n2566_));
  NAND3_X1   g2515(.A1(new_n2566_), .A2(new_n313_), .A3(new_n319_), .ZN(new_n2567_));
  NAND3_X1   g2516(.A1(new_n384_), .A2(new_n326_), .A3(new_n376_), .ZN(new_n2568_));
  NOR4_X1    g2517(.A1(new_n2568_), .A2(new_n201_), .A3(new_n314_), .A4(new_n505_), .ZN(new_n2569_));
  INV_X1     g2518(.I(new_n2569_), .ZN(new_n2570_));
  NOR4_X1    g2519(.A1(new_n2570_), .A2(new_n2567_), .A3(new_n471_), .A4(new_n659_), .ZN(new_n2571_));
  INV_X1     g2520(.I(new_n2571_), .ZN(new_n2572_));
  NOR4_X1    g2521(.A1(new_n2251_), .A2(new_n2312_), .A3(new_n201_), .A4(new_n452_), .ZN(new_n2573_));
  INV_X1     g2522(.I(new_n679_), .ZN(new_n2574_));
  NOR4_X1    g2523(.A1(new_n2574_), .A2(new_n222_), .A3(new_n461_), .A4(new_n538_), .ZN(new_n2575_));
  NAND3_X1   g2524(.A1(new_n2573_), .A2(new_n487_), .A3(new_n2575_), .ZN(new_n2576_));
  NOR3_X1    g2525(.A1(new_n2234_), .A2(new_n2576_), .A3(new_n2572_), .ZN(new_n2577_));
  INV_X1     g2526(.I(new_n2577_), .ZN(new_n2578_));
  NOR2_X1    g2527(.A1(new_n2565_), .A2(new_n2578_), .ZN(new_n2579_));
  OAI21_X1   g2528(.A1(new_n2518_), .A2(new_n2562_), .B(new_n2579_), .ZN(new_n2580_));
  NAND2_X1   g2529(.A1(new_n2580_), .A2(new_n2563_), .ZN(new_n2581_));
  NOR2_X1    g2530(.A1(new_n2064_), .A2(new_n2080_), .ZN(new_n2582_));
  AOI21_X1   g2531(.A1(new_n2582_), .A2(new_n2520_), .B(new_n2117_), .ZN(new_n2583_));
  NAND2_X1   g2532(.A1(new_n2557_), .A2(new_n2524_), .ZN(new_n2584_));
  NOR2_X1    g2533(.A1(new_n2552_), .A2(new_n2554_), .ZN(new_n2585_));
  NOR2_X1    g2534(.A1(new_n2585_), .A2(new_n2550_), .ZN(new_n2586_));
  NOR2_X1    g2535(.A1(new_n2533_), .A2(new_n2543_), .ZN(new_n2587_));
  NOR2_X1    g2536(.A1(new_n2587_), .A2(new_n2542_), .ZN(new_n2588_));
  NOR2_X1    g2537(.A1(new_n1056_), .A2(new_n875_), .ZN(new_n2589_));
  AOI21_X1   g2538(.A1(new_n571_), .A2(new_n875_), .B(new_n2589_), .ZN(new_n2590_));
  NOR3_X1    g2539(.A1(new_n2590_), .A2(new_n437_), .A3(new_n580_), .ZN(new_n2591_));
  NOR3_X1    g2540(.A1(new_n2590_), .A2(new_n438_), .A3(new_n565_), .ZN(new_n2592_));
  OAI21_X1   g2541(.A1(new_n2592_), .A2(new_n2591_), .B(new_n562_), .ZN(new_n2593_));
  XOR2_X1    g2542(.A1(new_n691_), .A2(new_n711_), .Z(new_n2594_));
  NAND2_X1   g2543(.A1(new_n2594_), .A2(new_n702_), .ZN(new_n2595_));
  XOR2_X1    g2544(.A1(new_n2595_), .A2(new_n266_), .Z(new_n2596_));
  XNOR2_X1   g2545(.A1(new_n2596_), .A2(new_n2593_), .ZN(new_n2597_));
  NOR2_X1    g2546(.A1(new_n2597_), .A2(new_n2588_), .ZN(new_n2598_));
  NOR2_X1    g2547(.A1(new_n2596_), .A2(new_n2593_), .ZN(new_n2599_));
  INV_X1     g2548(.I(new_n2599_), .ZN(new_n2600_));
  NAND2_X1   g2549(.A1(new_n2596_), .A2(new_n2593_), .ZN(new_n2601_));
  NAND2_X1   g2550(.A1(new_n2600_), .A2(new_n2601_), .ZN(new_n2602_));
  AOI21_X1   g2551(.A1(new_n2588_), .A2(new_n2602_), .B(new_n2598_), .ZN(new_n2603_));
  XOR2_X1    g2552(.A1(new_n2586_), .A2(new_n2603_), .Z(new_n2604_));
  INV_X1     g2553(.I(new_n2604_), .ZN(new_n2605_));
  NAND2_X1   g2554(.A1(new_n2559_), .A2(new_n2605_), .ZN(new_n2606_));
  XNOR2_X1   g2555(.A1(new_n2606_), .A2(new_n2584_), .ZN(new_n2607_));
  INV_X1     g2556(.I(new_n2607_), .ZN(new_n2608_));
  NAND2_X1   g2557(.A1(new_n2583_), .A2(new_n2608_), .ZN(new_n2609_));
  NAND2_X1   g2558(.A1(new_n2522_), .A2(new_n2607_), .ZN(new_n2610_));
  NAND2_X1   g2559(.A1(new_n2610_), .A2(new_n2609_), .ZN(new_n2611_));
  INV_X1     g2560(.I(new_n656_), .ZN(new_n2612_));
  NOR2_X1    g2561(.A1(new_n756_), .A2(new_n754_), .ZN(new_n2613_));
  INV_X1     g2562(.I(new_n2613_), .ZN(new_n2614_));
  INV_X1     g2563(.I(new_n482_), .ZN(new_n2615_));
  NOR2_X1    g2564(.A1(new_n2448_), .A2(new_n2386_), .ZN(new_n2616_));
  NAND4_X1   g2565(.A1(new_n318_), .A2(new_n360_), .A3(new_n329_), .A4(new_n750_), .ZN(new_n2617_));
  INV_X1     g2566(.I(new_n2617_), .ZN(new_n2618_));
  NAND4_X1   g2567(.A1(new_n2618_), .A2(new_n2616_), .A3(new_n2615_), .A4(new_n2395_), .ZN(new_n2619_));
  NAND3_X1   g2568(.A1(new_n350_), .A2(new_n214_), .A3(new_n465_), .ZN(new_n2620_));
  NOR4_X1    g2569(.A1(new_n2620_), .A2(new_n317_), .A3(new_n367_), .A4(new_n635_), .ZN(new_n2621_));
  NAND3_X1   g2570(.A1(new_n672_), .A2(new_n442_), .A3(new_n535_), .ZN(new_n2622_));
  NOR2_X1    g2571(.A1(new_n2622_), .A2(new_n414_), .ZN(new_n2623_));
  NAND4_X1   g2572(.A1(new_n2623_), .A2(new_n2621_), .A3(new_n327_), .A4(new_n760_), .ZN(new_n2624_));
  NOR4_X1    g2573(.A1(new_n2624_), .A2(new_n2612_), .A3(new_n2619_), .A4(new_n2614_), .ZN(new_n2625_));
  NAND2_X1   g2574(.A1(new_n2611_), .A2(new_n2625_), .ZN(new_n2626_));
  NAND3_X1   g2575(.A1(new_n2610_), .A2(new_n2609_), .A3(new_n2625_), .ZN(new_n2627_));
  NOR2_X1    g2576(.A1(new_n2522_), .A2(new_n2607_), .ZN(new_n2628_));
  NOR2_X1    g2577(.A1(new_n2583_), .A2(new_n2608_), .ZN(new_n2629_));
  INV_X1     g2578(.I(new_n2625_), .ZN(new_n2630_));
  OAI21_X1   g2579(.A1(new_n2628_), .A2(new_n2629_), .B(new_n2630_), .ZN(new_n2631_));
  NAND2_X1   g2580(.A1(new_n2631_), .A2(new_n2627_), .ZN(new_n2632_));
  NOR3_X1    g2581(.A1(new_n2585_), .A2(new_n2550_), .A3(new_n2603_), .ZN(new_n2633_));
  INV_X1     g2582(.I(new_n2633_), .ZN(new_n2634_));
  NOR2_X1    g2583(.A1(new_n2605_), .A2(new_n2557_), .ZN(new_n2635_));
  AOI21_X1   g2584(.A1(new_n2605_), .A2(new_n2557_), .B(new_n2524_), .ZN(new_n2636_));
  NOR2_X1    g2585(.A1(new_n2636_), .A2(new_n2635_), .ZN(new_n2637_));
  OAI21_X1   g2586(.A1(new_n2588_), .A2(new_n2599_), .B(new_n2601_), .ZN(new_n2638_));
  NOR2_X1    g2587(.A1(new_n266_), .A2(new_n711_), .ZN(new_n2639_));
  AOI21_X1   g2588(.A1(new_n266_), .A2(new_n711_), .B(new_n702_), .ZN(new_n2640_));
  NOR3_X1    g2589(.A1(new_n929_), .A2(new_n2639_), .A3(new_n2640_), .ZN(new_n2641_));
  AOI21_X1   g2590(.A1(new_n1053_), .A2(new_n566_), .B(new_n437_), .ZN(new_n2642_));
  AND3_X2    g2591(.A1(new_n1053_), .A2(new_n566_), .A3(new_n437_), .Z(new_n2643_));
  XOR2_X1    g2592(.A1(new_n559_), .A2(new_n266_), .Z(new_n2644_));
  NOR4_X1    g2593(.A1(new_n2643_), .A2(new_n1053_), .A3(new_n2642_), .A4(new_n2644_), .ZN(new_n2645_));
  NAND2_X1   g2594(.A1(new_n2645_), .A2(new_n2641_), .ZN(new_n2646_));
  XOR2_X1    g2595(.A1(new_n2646_), .A2(new_n266_), .Z(new_n2647_));
  XOR2_X1    g2596(.A1(new_n2647_), .A2(new_n875_), .Z(new_n2648_));
  XNOR2_X1   g2597(.A1(new_n2638_), .A2(new_n2648_), .ZN(new_n2649_));
  INV_X1     g2598(.I(new_n2247_), .ZN(new_n2650_));
  NOR2_X1    g2599(.A1(new_n292_), .A2(new_n522_), .ZN(new_n2651_));
  NAND4_X1   g2600(.A1(new_n2651_), .A2(new_n505_), .A3(new_n625_), .A4(new_n537_), .ZN(new_n2652_));
  NAND3_X1   g2601(.A1(new_n635_), .A2(new_n323_), .A3(new_n383_), .ZN(new_n2653_));
  NOR2_X1    g2602(.A1(new_n230_), .A2(new_n160_), .ZN(new_n2654_));
  NAND4_X1   g2603(.A1(new_n2654_), .A2(new_n600_), .A3(new_n413_), .A4(new_n253_), .ZN(new_n2655_));
  NOR3_X1    g2604(.A1(new_n2655_), .A2(new_n2652_), .A3(new_n2653_), .ZN(new_n2656_));
  NOR2_X1    g2605(.A1(new_n168_), .A2(new_n281_), .ZN(new_n2657_));
  NAND4_X1   g2606(.A1(new_n2657_), .A2(new_n234_), .A3(new_n223_), .A4(new_n304_), .ZN(new_n2658_));
  NOR4_X1    g2607(.A1(new_n1065_), .A2(new_n388_), .A3(new_n859_), .A4(new_n399_), .ZN(new_n2659_));
  INV_X1     g2608(.I(new_n2659_), .ZN(new_n2660_));
  NOR4_X1    g2609(.A1(new_n2660_), .A2(new_n2222_), .A3(new_n2658_), .A4(new_n595_), .ZN(new_n2661_));
  NAND4_X1   g2610(.A1(new_n2392_), .A2(new_n2661_), .A3(new_n2656_), .A4(new_n2650_), .ZN(new_n2662_));
  NOR2_X1    g2611(.A1(new_n2649_), .A2(new_n2662_), .ZN(new_n2663_));
  INV_X1     g2612(.I(new_n2663_), .ZN(new_n2664_));
  AOI21_X1   g2613(.A1(new_n2522_), .A2(new_n2637_), .B(new_n2664_), .ZN(new_n2665_));
  INV_X1     g2614(.I(new_n2637_), .ZN(new_n2666_));
  NOR3_X1    g2615(.A1(new_n2583_), .A2(new_n2666_), .A3(new_n2663_), .ZN(new_n2667_));
  OAI21_X1   g2616(.A1(new_n2665_), .A2(new_n2667_), .B(new_n2634_), .ZN(new_n2668_));
  OAI21_X1   g2617(.A1(new_n2583_), .A2(new_n2666_), .B(new_n2663_), .ZN(new_n2669_));
  NAND3_X1   g2618(.A1(new_n2522_), .A2(new_n2637_), .A3(new_n2664_), .ZN(new_n2670_));
  NAND3_X1   g2619(.A1(new_n2670_), .A2(new_n2669_), .A3(new_n2633_), .ZN(new_n2671_));
  NAND2_X1   g2620(.A1(new_n2668_), .A2(new_n2671_), .ZN(new_n2672_));
  NAND3_X1   g2621(.A1(new_n2672_), .A2(new_n2632_), .A3(new_n2626_), .ZN(new_n2673_));
  INV_X1     g2622(.I(new_n2611_), .ZN(new_n2674_));
  NOR2_X1    g2623(.A1(new_n2674_), .A2(new_n2630_), .ZN(new_n2676_));
  INV_X1     g2624(.I(new_n2676_), .ZN(new_n2677_));
  AND2_X2    g2625(.A1(new_n2673_), .A2(new_n2677_), .Z(new_n2678_));
  NOR2_X1    g2626(.A1(new_n2678_), .A2(new_n2581_), .ZN(new_n2679_));
  NAND2_X1   g2627(.A1(new_n2673_), .A2(new_n2677_), .ZN(new_n2680_));
  AOI21_X1   g2628(.A1(new_n2563_), .A2(new_n2580_), .B(new_n2680_), .ZN(new_n2681_));
  NOR2_X1    g2629(.A1(new_n2679_), .A2(new_n2681_), .ZN(new_n2682_));
  OR2_X2     g2630(.A1(new_n2255_), .A2(new_n2259_), .Z(new_n2683_));
  AOI22_X1   g2631(.A1(new_n2364_), .A2(new_n2323_), .B1(new_n2472_), .B2(new_n2457_), .ZN(new_n2684_));
  AOI21_X1   g2632(.A1(new_n2684_), .A2(new_n2365_), .B(new_n2481_), .ZN(new_n2685_));
  INV_X1     g2633(.I(new_n2510_), .ZN(new_n2686_));
  OAI21_X1   g2634(.A1(new_n2685_), .A2(new_n2686_), .B(new_n2482_), .ZN(new_n2687_));
  OAI21_X1   g2635(.A1(new_n2512_), .A2(new_n2513_), .B(new_n2290_), .ZN(new_n2688_));
  NAND2_X1   g2636(.A1(new_n2688_), .A2(new_n2292_), .ZN(new_n2689_));
  OAI21_X1   g2637(.A1(new_n2687_), .A2(new_n2689_), .B(new_n2292_), .ZN(new_n2690_));
  NAND2_X1   g2638(.A1(new_n2690_), .A2(new_n2683_), .ZN(new_n2691_));
  NOR2_X1    g2639(.A1(new_n2522_), .A2(new_n2561_), .ZN(new_n2692_));
  AOI21_X1   g2640(.A1(new_n2522_), .A2(new_n2559_), .B(new_n2692_), .ZN(new_n2693_));
  NOR2_X1    g2641(.A1(new_n2691_), .A2(new_n2693_), .ZN(new_n2694_));
  INV_X1     g2642(.I(new_n2579_), .ZN(new_n2695_));
  AOI21_X1   g2643(.A1(new_n2691_), .A2(new_n2693_), .B(new_n2695_), .ZN(new_n2696_));
  NAND2_X1   g2644(.A1(new_n2674_), .A2(new_n2630_), .ZN(new_n2697_));
  NAND2_X1   g2645(.A1(new_n2697_), .A2(new_n2626_), .ZN(new_n2698_));
  OAI21_X1   g2646(.A1(new_n2696_), .A2(new_n2694_), .B(new_n2698_), .ZN(new_n2699_));
  NAND3_X1   g2647(.A1(new_n2580_), .A2(new_n2563_), .A3(new_n2632_), .ZN(new_n2700_));
  NAND2_X1   g2648(.A1(new_n2699_), .A2(new_n2700_), .ZN(new_n2701_));
  NAND2_X1   g2649(.A1(new_n2562_), .A2(new_n2577_), .ZN(new_n2702_));
  AOI21_X1   g2650(.A1(new_n2683_), .A2(new_n2690_), .B(new_n2702_), .ZN(new_n2703_));
  AOI21_X1   g2651(.A1(new_n2208_), .A2(new_n2207_), .B(new_n2266_), .ZN(new_n2704_));
  INV_X1     g2652(.I(new_n2479_), .ZN(new_n2705_));
  NOR3_X1    g2653(.A1(new_n2063_), .A2(new_n2053_), .A3(new_n2705_), .ZN(new_n2706_));
  NOR2_X1    g2654(.A1(new_n2704_), .A2(new_n2706_), .ZN(new_n2707_));
  NOR4_X1    g2655(.A1(new_n2488_), .A2(new_n2491_), .A3(new_n2707_), .A4(new_n2490_), .ZN(new_n2708_));
  NAND2_X1   g2656(.A1(new_n2473_), .A2(new_n2476_), .ZN(new_n2709_));
  OAI21_X1   g2657(.A1(new_n2709_), .A2(new_n2488_), .B(new_n2707_), .ZN(new_n2710_));
  AOI21_X1   g2658(.A1(new_n2710_), .A2(new_n2510_), .B(new_n2708_), .ZN(new_n2711_));
  AOI21_X1   g2659(.A1(new_n2711_), .A2(new_n2516_), .B(new_n2514_), .ZN(new_n2712_));
  NOR2_X1    g2660(.A1(new_n2693_), .A2(new_n2578_), .ZN(new_n2713_));
  NOR3_X1    g2661(.A1(new_n2712_), .A2(new_n2713_), .A3(new_n2260_), .ZN(new_n2714_));
  OAI21_X1   g2662(.A1(new_n2714_), .A2(new_n2703_), .B(new_n2565_), .ZN(new_n2715_));
  INV_X1     g2663(.I(new_n2565_), .ZN(new_n2716_));
  OAI21_X1   g2664(.A1(new_n2712_), .A2(new_n2260_), .B(new_n2713_), .ZN(new_n2717_));
  NAND3_X1   g2665(.A1(new_n2690_), .A2(new_n2702_), .A3(new_n2683_), .ZN(new_n2718_));
  NAND3_X1   g2666(.A1(new_n2717_), .A2(new_n2718_), .A3(new_n2716_), .ZN(new_n2719_));
  NAND2_X1   g2667(.A1(new_n2715_), .A2(new_n2719_), .ZN(new_n2720_));
  AOI21_X1   g2668(.A1(new_n2717_), .A2(new_n2718_), .B(new_n2716_), .ZN(new_n2721_));
  NOR3_X1    g2669(.A1(new_n2714_), .A2(new_n2703_), .A3(new_n2565_), .ZN(new_n2722_));
  OAI21_X1   g2670(.A1(new_n2215_), .A2(new_n2219_), .B(new_n2258_), .ZN(new_n2723_));
  AOI21_X1   g2671(.A1(new_n2711_), .A2(new_n2516_), .B(new_n2723_), .ZN(new_n2724_));
  AOI21_X1   g2672(.A1(new_n2256_), .A2(new_n2257_), .B(new_n2254_), .ZN(new_n2725_));
  NOR3_X1    g2673(.A1(new_n2687_), .A2(new_n2689_), .A3(new_n2725_), .ZN(new_n2726_));
  OAI21_X1   g2674(.A1(new_n2724_), .A2(new_n2726_), .B(new_n2292_), .ZN(new_n2727_));
  OAI21_X1   g2675(.A1(new_n2564_), .A2(new_n2254_), .B(new_n2514_), .ZN(new_n2728_));
  NAND2_X1   g2676(.A1(new_n2727_), .A2(new_n2728_), .ZN(new_n2729_));
  NAND3_X1   g2677(.A1(new_n2365_), .A2(new_n2473_), .A3(new_n2476_), .ZN(new_n2730_));
  AOI21_X1   g2678(.A1(new_n2730_), .A2(new_n2707_), .B(new_n2686_), .ZN(new_n2731_));
  NOR3_X1    g2679(.A1(new_n2731_), .A2(new_n2708_), .A3(new_n2689_), .ZN(new_n2732_));
  AOI21_X1   g2680(.A1(new_n2511_), .A2(new_n2482_), .B(new_n2516_), .ZN(new_n2733_));
  NOR2_X1    g2681(.A1(new_n2733_), .A2(new_n2732_), .ZN(new_n2734_));
  OAI21_X1   g2682(.A1(new_n2704_), .A2(new_n2706_), .B(new_n2508_), .ZN(new_n2735_));
  AOI21_X1   g2683(.A1(new_n2684_), .A2(new_n2365_), .B(new_n2735_), .ZN(new_n2736_));
  AOI21_X1   g2684(.A1(new_n2480_), .A2(new_n2477_), .B(new_n2509_), .ZN(new_n2737_));
  NOR4_X1    g2685(.A1(new_n2488_), .A2(new_n2737_), .A3(new_n2491_), .A4(new_n2490_), .ZN(new_n2738_));
  OAI21_X1   g2686(.A1(new_n2736_), .A2(new_n2738_), .B(new_n2495_), .ZN(new_n2739_));
  OAI21_X1   g2687(.A1(new_n2709_), .A2(new_n2488_), .B(new_n2737_), .ZN(new_n2740_));
  NAND3_X1   g2688(.A1(new_n2684_), .A2(new_n2365_), .A3(new_n2735_), .ZN(new_n2741_));
  NAND3_X1   g2689(.A1(new_n2740_), .A2(new_n2494_), .A3(new_n2741_), .ZN(new_n2742_));
  NAND2_X1   g2690(.A1(new_n2742_), .A2(new_n2739_), .ZN(new_n2743_));
  NOR2_X1    g2691(.A1(new_n2309_), .A2(new_n2323_), .ZN(new_n2744_));
  NOR3_X1    g2692(.A1(new_n2308_), .A2(new_n2304_), .A3(new_n2323_), .ZN(new_n2745_));
  AOI21_X1   g2693(.A1(new_n2483_), .A2(new_n2484_), .B(new_n2486_), .ZN(new_n2746_));
  NOR2_X1    g2694(.A1(new_n2746_), .A2(new_n2745_), .ZN(new_n2747_));
  NOR3_X1    g2695(.A1(new_n2364_), .A2(new_n2747_), .A3(new_n2744_), .ZN(new_n2748_));
  NOR2_X1    g2696(.A1(new_n2309_), .A2(new_n2323_), .ZN(new_n2749_));
  OAI21_X1   g2697(.A1(new_n2748_), .A2(new_n2749_), .B(new_n2490_), .ZN(new_n2750_));
  NAND2_X1   g2698(.A1(new_n2485_), .A2(new_n2486_), .ZN(new_n2751_));
  NAND3_X1   g2699(.A1(new_n2483_), .A2(new_n2484_), .A3(new_n2486_), .ZN(new_n2752_));
  OAI21_X1   g2700(.A1(new_n2308_), .A2(new_n2304_), .B(new_n2323_), .ZN(new_n2753_));
  NAND2_X1   g2701(.A1(new_n2753_), .A2(new_n2752_), .ZN(new_n2754_));
  NAND3_X1   g2702(.A1(new_n2487_), .A2(new_n2754_), .A3(new_n2751_), .ZN(new_n2755_));
  INV_X1     g2703(.I(new_n2749_), .ZN(new_n2756_));
  NAND3_X1   g2704(.A1(new_n2755_), .A2(new_n2473_), .A3(new_n2756_), .ZN(new_n2757_));
  NAND2_X1   g2705(.A1(new_n2750_), .A2(new_n2757_), .ZN(new_n2758_));
  NOR2_X1    g2706(.A1(new_n1872_), .A2(new_n2296_), .ZN(new_n2759_));
  AOI21_X1   g2707(.A1(new_n1872_), .A2(new_n2459_), .B(new_n2759_), .ZN(new_n2760_));
  NOR3_X1    g2708(.A1(new_n2434_), .A2(new_n2424_), .A3(new_n2456_), .ZN(new_n2761_));
  NOR2_X1    g2709(.A1(new_n2761_), .A2(new_n2760_), .ZN(new_n2762_));
  NOR3_X1    g2710(.A1(new_n2762_), .A2(new_n2754_), .A3(new_n2489_), .ZN(new_n2763_));
  NOR2_X1    g2711(.A1(new_n2490_), .A2(new_n2747_), .ZN(new_n2764_));
  NOR2_X1    g2712(.A1(new_n2764_), .A2(new_n2763_), .ZN(new_n2765_));
  AOI21_X1   g2713(.A1(new_n2471_), .A2(new_n2457_), .B(new_n2760_), .ZN(new_n2766_));
  NAND3_X1   g2714(.A1(new_n2470_), .A2(new_n2467_), .A3(new_n2456_), .ZN(new_n2767_));
  OAI21_X1   g2715(.A1(new_n2434_), .A2(new_n2424_), .B(new_n2455_), .ZN(new_n2768_));
  AOI21_X1   g2716(.A1(new_n2767_), .A2(new_n2768_), .B(new_n2461_), .ZN(new_n2769_));
  NOR2_X1    g2717(.A1(new_n2766_), .A2(new_n2769_), .ZN(new_n2770_));
  OAI21_X1   g2718(.A1(new_n2489_), .A2(new_n2761_), .B(new_n2461_), .ZN(new_n2771_));
  NOR3_X1    g2719(.A1(new_n2434_), .A2(new_n2424_), .A3(new_n2455_), .ZN(new_n2772_));
  AOI21_X1   g2720(.A1(new_n2470_), .A2(new_n2467_), .B(new_n2456_), .ZN(new_n2773_));
  OAI21_X1   g2721(.A1(new_n2773_), .A2(new_n2772_), .B(new_n2760_), .ZN(new_n2774_));
  NAND2_X1   g2722(.A1(new_n2771_), .A2(new_n2774_), .ZN(new_n2775_));
  NOR2_X1    g2723(.A1(new_n2469_), .A2(new_n2468_), .ZN(new_n2776_));
  NAND2_X1   g2724(.A1(new_n2402_), .A2(new_n2423_), .ZN(new_n2777_));
  AOI21_X1   g2725(.A1(new_n2467_), .A2(new_n2777_), .B(new_n2776_), .ZN(new_n2778_));
  NAND2_X1   g2726(.A1(new_n2430_), .A2(new_n2433_), .ZN(new_n2779_));
  NAND2_X1   g2727(.A1(new_n2402_), .A2(new_n2466_), .ZN(new_n2780_));
  NAND2_X1   g2728(.A1(new_n2465_), .A2(new_n2423_), .ZN(new_n2781_));
  AOI21_X1   g2729(.A1(new_n2780_), .A2(new_n2781_), .B(new_n2779_), .ZN(new_n2782_));
  OR2_X2     g2730(.A1(new_n2778_), .A2(new_n2782_), .Z(new_n2783_));
  NAND3_X1   g2731(.A1(new_n2380_), .A2(new_n2383_), .A3(new_n2464_), .ZN(new_n2784_));
  OAI21_X1   g2732(.A1(new_n2463_), .A2(new_n2462_), .B(new_n2401_), .ZN(new_n2785_));
  NAND2_X1   g2733(.A1(new_n2785_), .A2(new_n2784_), .ZN(new_n2786_));
  AOI21_X1   g2734(.A1(new_n2775_), .A2(new_n2786_), .B(new_n2783_), .ZN(new_n2787_));
  NOR4_X1    g2735(.A1(new_n2758_), .A2(new_n2765_), .A3(new_n2770_), .A4(new_n2787_), .ZN(new_n2788_));
  NAND3_X1   g2736(.A1(new_n2472_), .A2(new_n2747_), .A3(new_n2457_), .ZN(new_n2789_));
  OAI21_X1   g2737(.A1(new_n2762_), .A2(new_n2489_), .B(new_n2754_), .ZN(new_n2790_));
  NAND2_X1   g2738(.A1(new_n2790_), .A2(new_n2789_), .ZN(new_n2791_));
  NOR2_X1    g2739(.A1(new_n2778_), .A2(new_n2782_), .ZN(new_n2792_));
  NOR3_X1    g2740(.A1(new_n2463_), .A2(new_n2462_), .A3(new_n2401_), .ZN(new_n2793_));
  AOI21_X1   g2741(.A1(new_n2380_), .A2(new_n2383_), .B(new_n2464_), .ZN(new_n2794_));
  NOR2_X1    g2742(.A1(new_n2794_), .A2(new_n2793_), .ZN(new_n2795_));
  NAND2_X1   g2743(.A1(new_n2770_), .A2(new_n2792_), .ZN(new_n2796_));
  NOR2_X1    g2744(.A1(new_n2796_), .A2(new_n2791_), .ZN(new_n2797_));
  OAI21_X1   g2745(.A1(new_n2770_), .A2(new_n2795_), .B(new_n2792_), .ZN(new_n2798_));
  NAND3_X1   g2746(.A1(new_n2798_), .A2(new_n2791_), .A3(new_n2775_), .ZN(new_n2799_));
  NAND3_X1   g2747(.A1(new_n2799_), .A2(new_n2797_), .A3(new_n2758_), .ZN(new_n2800_));
  OAI21_X1   g2748(.A1(new_n2788_), .A2(new_n2800_), .B(new_n2743_), .ZN(new_n2801_));
  AOI21_X1   g2749(.A1(new_n2755_), .A2(new_n2756_), .B(new_n2473_), .ZN(new_n2802_));
  NOR3_X1    g2750(.A1(new_n2748_), .A2(new_n2490_), .A3(new_n2749_), .ZN(new_n2803_));
  NOR2_X1    g2751(.A1(new_n2803_), .A2(new_n2802_), .ZN(new_n2804_));
  NOR2_X1    g2752(.A1(new_n2775_), .A2(new_n2783_), .ZN(new_n2805_));
  NAND2_X1   g2753(.A1(new_n2765_), .A2(new_n2805_), .ZN(new_n2806_));
  NOR3_X1    g2754(.A1(new_n2787_), .A2(new_n2765_), .A3(new_n2770_), .ZN(new_n2807_));
  NOR3_X1    g2755(.A1(new_n2807_), .A2(new_n2806_), .A3(new_n2804_), .ZN(new_n2808_));
  NOR2_X1    g2756(.A1(new_n2743_), .A2(new_n2788_), .ZN(new_n2809_));
  NAND2_X1   g2757(.A1(new_n2801_), .A2(new_n2734_), .ZN(new_n2810_));
  OAI22_X1   g2758(.A1(new_n2722_), .A2(new_n2721_), .B1(new_n2729_), .B2(new_n2810_), .ZN(new_n2811_));
  NAND2_X1   g2759(.A1(new_n2687_), .A2(new_n2689_), .ZN(new_n2812_));
  NAND2_X1   g2760(.A1(new_n2812_), .A2(new_n2517_), .ZN(new_n2813_));
  OAI22_X1   g2761(.A1(new_n2743_), .A2(new_n2788_), .B1(new_n2732_), .B2(new_n2733_), .ZN(new_n2814_));
  NAND2_X1   g2762(.A1(new_n2801_), .A2(new_n2814_), .ZN(new_n2815_));
  NAND3_X1   g2763(.A1(new_n2815_), .A2(new_n2729_), .A3(new_n2813_), .ZN(new_n2816_));
  NAND2_X1   g2764(.A1(new_n2811_), .A2(new_n2816_), .ZN(new_n2817_));
  NAND4_X1   g2765(.A1(new_n2817_), .A2(new_n2682_), .A3(new_n2701_), .A4(new_n2720_), .ZN(new_n2818_));
  INV_X1     g2766(.I(new_n2818_), .ZN(new_n2819_));
  XNOR2_X1   g2767(.A1(new_n2633_), .A2(new_n2663_), .ZN(new_n2820_));
  NOR3_X1    g2768(.A1(new_n2583_), .A2(new_n2666_), .A3(new_n2820_), .ZN(new_n2821_));
  INV_X1     g2769(.I(new_n2821_), .ZN(new_n2822_));
  AOI21_X1   g2770(.A1(new_n2670_), .A2(new_n2669_), .B(new_n2633_), .ZN(new_n2823_));
  NOR3_X1    g2771(.A1(new_n2665_), .A2(new_n2667_), .A3(new_n2634_), .ZN(new_n2824_));
  NOR2_X1    g2772(.A1(new_n2823_), .A2(new_n2824_), .ZN(new_n2825_));
  NAND2_X1   g2773(.A1(new_n2825_), .A2(new_n2630_), .ZN(new_n2826_));
  NOR2_X1    g2774(.A1(new_n2825_), .A2(new_n2630_), .ZN(new_n2827_));
  OAI21_X1   g2775(.A1(new_n2611_), .A2(new_n2827_), .B(new_n2826_), .ZN(new_n2828_));
  AOI21_X1   g2776(.A1(new_n2563_), .A2(new_n2580_), .B(new_n2828_), .ZN(new_n2829_));
  NAND2_X1   g2777(.A1(new_n2633_), .A2(new_n2638_), .ZN(new_n2830_));
  NOR2_X1    g2778(.A1(new_n2633_), .A2(new_n2638_), .ZN(new_n2831_));
  NOR2_X1    g2779(.A1(new_n2831_), .A2(new_n2648_), .ZN(new_n2832_));
  NAND3_X1   g2780(.A1(new_n2522_), .A2(new_n2637_), .A3(new_n2832_), .ZN(new_n2833_));
  NAND2_X1   g2781(.A1(new_n2833_), .A2(new_n2830_), .ZN(new_n2834_));
  NOR2_X1    g2782(.A1(new_n566_), .A2(new_n645_), .ZN(new_n2835_));
  OAI21_X1   g2783(.A1(new_n2645_), .A2(new_n2641_), .B(new_n2835_), .ZN(new_n2836_));
  NAND2_X1   g2784(.A1(new_n2836_), .A2(new_n2646_), .ZN(new_n2837_));
  XOR2_X1    g2785(.A1(new_n645_), .A2(new_n437_), .Z(new_n2838_));
  INV_X1     g2786(.I(new_n2838_), .ZN(new_n2839_));
  NAND2_X1   g2787(.A1(new_n266_), .A2(new_n2839_), .ZN(new_n2840_));
  XOR2_X1    g2788(.A1(new_n2840_), .A2(new_n552_), .Z(new_n2841_));
  NOR2_X1    g2789(.A1(new_n2841_), .A2(new_n559_), .ZN(new_n2842_));
  XNOR2_X1   g2790(.A1(new_n2837_), .A2(new_n2842_), .ZN(new_n2843_));
  INV_X1     g2791(.I(new_n2843_), .ZN(new_n2844_));
  XOR2_X1    g2792(.A1(new_n2837_), .A2(new_n2842_), .Z(new_n2845_));
  NOR2_X1    g2793(.A1(new_n2834_), .A2(new_n2845_), .ZN(new_n2846_));
  AOI21_X1   g2794(.A1(new_n2834_), .A2(new_n2844_), .B(new_n2846_), .ZN(new_n2847_));
  NOR4_X1    g2795(.A1(new_n450_), .A2(new_n203_), .A3(new_n366_), .A4(new_n424_), .ZN(new_n2848_));
  NOR4_X1    g2796(.A1(new_n312_), .A2(new_n191_), .A3(new_n398_), .A4(new_n317_), .ZN(new_n2849_));
  AND3_X2    g2797(.A1(new_n2849_), .A2(new_n2848_), .A3(new_n765_), .Z(new_n2850_));
  INV_X1     g2798(.I(new_n2850_), .ZN(new_n2851_));
  NOR2_X1    g2799(.A1(new_n548_), .A2(new_n228_), .ZN(new_n2852_));
  NOR2_X1    g2800(.A1(new_n205_), .A2(new_n313_), .ZN(new_n2853_));
  INV_X1     g2801(.I(new_n2853_), .ZN(new_n2854_));
  NOR2_X1    g2802(.A1(new_n2854_), .A2(new_n2237_), .ZN(new_n2855_));
  NOR2_X1    g2803(.A1(new_n388_), .A2(new_n420_), .ZN(new_n2856_));
  NAND4_X1   g2804(.A1(new_n2856_), .A2(new_n168_), .A3(new_n221_), .A4(new_n250_), .ZN(new_n2857_));
  INV_X1     g2805(.I(new_n2857_), .ZN(new_n2858_));
  INV_X1     g2806(.I(new_n500_), .ZN(new_n2859_));
  NOR4_X1    g2807(.A1(new_n2859_), .A2(new_n213_), .A3(new_n241_), .A4(new_n660_), .ZN(new_n2860_));
  NAND4_X1   g2808(.A1(new_n2858_), .A2(new_n2855_), .A3(new_n2852_), .A4(new_n2860_), .ZN(new_n2861_));
  NOR4_X1    g2809(.A1(new_n2224_), .A2(new_n243_), .A3(new_n442_), .A4(new_n625_), .ZN(new_n2862_));
  INV_X1     g2810(.I(new_n2862_), .ZN(new_n2863_));
  NOR4_X1    g2811(.A1(new_n2851_), .A2(new_n762_), .A3(new_n2861_), .A4(new_n2863_), .ZN(new_n2864_));
  AND2_X2    g2812(.A1(new_n2864_), .A2(new_n2337_), .Z(new_n2865_));
  INV_X1     g2813(.I(new_n2865_), .ZN(new_n2866_));
  NOR2_X1    g2814(.A1(new_n2847_), .A2(new_n2866_), .ZN(new_n2867_));
  INV_X1     g2815(.I(new_n2867_), .ZN(new_n2868_));
  NOR2_X1    g2816(.A1(new_n2829_), .A2(new_n2868_), .ZN(new_n2869_));
  NOR2_X1    g2817(.A1(new_n2672_), .A2(new_n2625_), .ZN(new_n2870_));
  NAND2_X1   g2818(.A1(new_n2672_), .A2(new_n2625_), .ZN(new_n2871_));
  AOI21_X1   g2819(.A1(new_n2674_), .A2(new_n2871_), .B(new_n2870_), .ZN(new_n2872_));
  NAND2_X1   g2820(.A1(new_n2581_), .A2(new_n2872_), .ZN(new_n2873_));
  NOR2_X1    g2821(.A1(new_n2873_), .A2(new_n2867_), .ZN(new_n2874_));
  OAI21_X1   g2822(.A1(new_n2869_), .A2(new_n2874_), .B(new_n2822_), .ZN(new_n2875_));
  NAND2_X1   g2823(.A1(new_n2873_), .A2(new_n2867_), .ZN(new_n2876_));
  NAND3_X1   g2824(.A1(new_n2868_), .A2(new_n2581_), .A3(new_n2872_), .ZN(new_n2877_));
  NAND3_X1   g2825(.A1(new_n2876_), .A2(new_n2821_), .A3(new_n2877_), .ZN(new_n2878_));
  NAND2_X1   g2826(.A1(new_n2875_), .A2(new_n2878_), .ZN(new_n2879_));
  NOR4_X1    g2827(.A1(new_n2817_), .A2(new_n2682_), .A3(new_n2701_), .A4(new_n2720_), .ZN(new_n2880_));
  INV_X1     g2828(.I(new_n2880_), .ZN(new_n2881_));
  AOI21_X1   g2829(.A1(new_n2879_), .A2(new_n2881_), .B(new_n2819_), .ZN(new_n2882_));
  NOR2_X1    g2830(.A1(new_n2873_), .A2(new_n2847_), .ZN(new_n2883_));
  NOR2_X1    g2831(.A1(new_n2822_), .A2(new_n2866_), .ZN(new_n2884_));
  INV_X1     g2832(.I(new_n2884_), .ZN(new_n2885_));
  AOI21_X1   g2833(.A1(new_n2873_), .A2(new_n2847_), .B(new_n2885_), .ZN(new_n2886_));
  NOR2_X1    g2834(.A1(new_n2886_), .A2(new_n2883_), .ZN(new_n2887_));
  NAND3_X1   g2835(.A1(new_n1137_), .A2(new_n649_), .A3(new_n546_), .ZN(new_n2888_));
  NAND4_X1   g2836(.A1(new_n232_), .A2(new_n356_), .A3(new_n273_), .A4(new_n383_), .ZN(new_n2889_));
  NOR4_X1    g2837(.A1(new_n2888_), .A2(new_n2386_), .A3(new_n538_), .A4(new_n2889_), .ZN(new_n2890_));
  NOR4_X1    g2838(.A1(new_n2235_), .A2(new_n921_), .A3(new_n205_), .A4(new_n447_), .ZN(new_n2891_));
  NAND2_X1   g2839(.A1(new_n2891_), .A2(new_n330_), .ZN(new_n2892_));
  NOR2_X1    g2840(.A1(new_n2892_), .A2(new_n666_), .ZN(new_n2893_));
  NAND4_X1   g2841(.A1(new_n2893_), .A2(new_n1100_), .A3(new_n2416_), .A4(new_n2890_), .ZN(new_n2894_));
  INV_X1     g2842(.I(new_n2894_), .ZN(new_n2895_));
  NAND2_X1   g2843(.A1(new_n2887_), .A2(new_n2895_), .ZN(new_n2896_));
  OAI21_X1   g2844(.A1(new_n2886_), .A2(new_n2883_), .B(new_n2894_), .ZN(new_n2897_));
  NAND2_X1   g2845(.A1(new_n2896_), .A2(new_n2897_), .ZN(new_n2898_));
  XOR2_X1    g2846(.A1(new_n2898_), .A2(new_n2879_), .Z(new_n2899_));
  NOR3_X1    g2847(.A1(new_n2886_), .A2(new_n2883_), .A3(new_n2894_), .ZN(new_n2900_));
  INV_X1     g2848(.I(new_n2897_), .ZN(new_n2901_));
  NOR2_X1    g2849(.A1(new_n2901_), .A2(new_n2900_), .ZN(new_n2902_));
  INV_X1     g2850(.I(new_n2847_), .ZN(new_n2903_));
  NAND2_X1   g2851(.A1(new_n2829_), .A2(new_n2903_), .ZN(new_n2904_));
  OAI21_X1   g2852(.A1(new_n2829_), .A2(new_n2903_), .B(new_n2884_), .ZN(new_n2905_));
  NAND2_X1   g2853(.A1(new_n2905_), .A2(new_n2904_), .ZN(new_n2906_));
  NAND4_X1   g2854(.A1(new_n228_), .A2(new_n384_), .A3(new_n292_), .A4(new_n420_), .ZN(new_n2907_));
  NOR4_X1    g2855(.A1(new_n2222_), .A2(new_n2907_), .A3(new_n372_), .A4(new_n253_), .ZN(new_n2908_));
  NAND2_X1   g2856(.A1(new_n347_), .A2(new_n332_), .ZN(new_n2909_));
  NOR3_X1    g2857(.A1(new_n307_), .A2(new_n388_), .A3(new_n859_), .ZN(new_n2910_));
  INV_X1     g2858(.I(new_n2910_), .ZN(new_n2911_));
  NOR2_X1    g2859(.A1(new_n891_), .A2(new_n383_), .ZN(new_n2912_));
  NAND4_X1   g2860(.A1(new_n2912_), .A2(new_n201_), .A3(new_n668_), .A4(new_n424_), .ZN(new_n2913_));
  NOR4_X1    g2861(.A1(new_n2911_), .A2(new_n2909_), .A3(new_n2913_), .A4(new_n537_), .ZN(new_n2914_));
  AND2_X2    g2862(.A1(new_n2908_), .A2(new_n2914_), .Z(new_n2915_));
  INV_X1     g2863(.I(new_n2343_), .ZN(new_n2916_));
  NOR4_X1    g2864(.A1(new_n675_), .A2(new_n160_), .A3(new_n201_), .A4(new_n209_), .ZN(new_n2917_));
  INV_X1     g2865(.I(new_n2566_), .ZN(new_n2918_));
  NOR2_X1    g2866(.A1(new_n2918_), .A2(new_n841_), .ZN(new_n2919_));
  NOR3_X1    g2867(.A1(new_n323_), .A2(new_n233_), .A3(new_n240_), .ZN(new_n2920_));
  NAND4_X1   g2868(.A1(new_n2919_), .A2(new_n1136_), .A3(new_n2917_), .A4(new_n2920_), .ZN(new_n2921_));
  NOR4_X1    g2869(.A1(new_n2921_), .A2(new_n422_), .A3(new_n423_), .A4(new_n2916_), .ZN(new_n2922_));
  NAND3_X1   g2870(.A1(new_n2915_), .A2(new_n2922_), .A3(new_n607_), .ZN(new_n2923_));
  OAI21_X1   g2871(.A1(new_n2886_), .A2(new_n2883_), .B(new_n2895_), .ZN(new_n2924_));
  NOR2_X1    g2872(.A1(new_n2923_), .A2(new_n2894_), .ZN(new_n2925_));
  AOI22_X1   g2873(.A1(new_n2923_), .A2(new_n2924_), .B1(new_n2906_), .B2(new_n2925_), .ZN(new_n2926_));
  XOR2_X1    g2874(.A1(new_n2902_), .A2(new_n2926_), .Z(new_n2927_));
  NAND3_X1   g2875(.A1(new_n2927_), .A2(new_n2899_), .A3(new_n2882_), .ZN(new_n2928_));
  AOI21_X1   g2876(.A1(new_n2876_), .A2(new_n2877_), .B(new_n2821_), .ZN(new_n2929_));
  NOR3_X1    g2877(.A1(new_n2869_), .A2(new_n2874_), .A3(new_n2822_), .ZN(new_n2930_));
  NOR2_X1    g2878(.A1(new_n2930_), .A2(new_n2929_), .ZN(new_n2931_));
  OAI21_X1   g2879(.A1(new_n2931_), .A2(new_n2880_), .B(new_n2818_), .ZN(new_n2932_));
  NAND2_X1   g2880(.A1(new_n2927_), .A2(new_n2899_), .ZN(new_n2933_));
  NAND2_X1   g2881(.A1(new_n2933_), .A2(new_n2932_), .ZN(new_n2934_));
  NAND2_X1   g2882(.A1(new_n2934_), .A2(new_n2928_), .ZN(new_n2935_));
  INV_X1     g2883(.I(\a[2] ), .ZN(new_n2936_));
  NOR2_X1    g2884(.A1(new_n2936_), .A2(\a[1] ), .ZN(new_n2937_));
  NOR2_X1    g2885(.A1(new_n1118_), .A2(\a[2] ), .ZN(new_n2938_));
  OAI21_X1   g2886(.A1(new_n2937_), .A2(new_n2938_), .B(\a[22] ), .ZN(new_n2939_));
  INV_X1     g2887(.I(new_n2939_), .ZN(new_n2940_));
  OAI21_X1   g2888(.A1(\a[2] ), .A2(\a[22] ), .B(\a[1] ), .ZN(new_n2941_));
  XOR2_X1    g2889(.A1(new_n2941_), .A2(\a[0] ), .Z(new_n2942_));
  INV_X1     g2890(.I(new_n2942_), .ZN(new_n2943_));
  NAND2_X1   g2891(.A1(new_n2924_), .A2(new_n2923_), .ZN(new_n2944_));
  NAND2_X1   g2892(.A1(new_n2906_), .A2(new_n2925_), .ZN(new_n2945_));
  NAND2_X1   g2893(.A1(new_n2944_), .A2(new_n2945_), .ZN(new_n2946_));
  NOR2_X1    g2894(.A1(new_n92_), .A2(new_n2936_), .ZN(new_n2947_));
  NAND2_X1   g2895(.A1(new_n2898_), .A2(new_n2947_), .ZN(new_n2948_));
  NOR2_X1    g2896(.A1(new_n1118_), .A2(\a[0] ), .ZN(new_n2949_));
  NAND2_X1   g2897(.A1(new_n2879_), .A2(new_n2949_), .ZN(new_n2950_));
  AOI22_X1   g2898(.A1(new_n2948_), .A2(new_n2950_), .B1(new_n2946_), .B2(new_n2940_), .ZN(new_n2951_));
  OAI21_X1   g2899(.A1(new_n2951_), .A2(new_n2943_), .B(new_n2940_), .ZN(new_n2952_));
  XOR2_X1    g2900(.A1(new_n2935_), .A2(new_n2952_), .Z(new_n2953_));
  AOI21_X1   g2901(.A1(new_n2740_), .A2(new_n2741_), .B(new_n2494_), .ZN(new_n2954_));
  NOR3_X1    g2902(.A1(new_n2736_), .A2(new_n2738_), .A3(new_n2495_), .ZN(new_n2955_));
  NOR2_X1    g2903(.A1(new_n2954_), .A2(new_n2955_), .ZN(new_n2956_));
  OAI21_X1   g2904(.A1(new_n2807_), .A2(new_n2806_), .B(new_n2758_), .ZN(new_n2957_));
  NAND2_X1   g2905(.A1(new_n2806_), .A2(new_n2758_), .ZN(new_n2958_));
  NAND3_X1   g2906(.A1(new_n2958_), .A2(new_n2804_), .A3(new_n2799_), .ZN(new_n2959_));
  AOI21_X1   g2907(.A1(new_n2959_), .A2(new_n2957_), .B(new_n2956_), .ZN(new_n2960_));
  AOI22_X1   g2908(.A1(new_n2765_), .A2(new_n2805_), .B1(new_n2750_), .B2(new_n2757_), .ZN(new_n2961_));
  OAI21_X1   g2909(.A1(new_n2961_), .A2(new_n2807_), .B(new_n2804_), .ZN(new_n2962_));
  AOI21_X1   g2910(.A1(new_n2962_), .A2(new_n2800_), .B(new_n2743_), .ZN(new_n2963_));
  NOR2_X1    g2911(.A1(new_n2960_), .A2(new_n2963_), .ZN(new_n2964_));
  NOR2_X1    g2912(.A1(new_n803_), .A2(new_n1149_), .ZN(new_n2965_));
  NOR2_X1    g2913(.A1(new_n1151_), .A2(new_n802_), .ZN(new_n2966_));
  XNOR2_X1   g2914(.A1(new_n808_), .A2(new_n1050_), .ZN(new_n2967_));
  INV_X1     g2915(.I(new_n2967_), .ZN(new_n2968_));
  OAI21_X1   g2916(.A1(new_n2965_), .A2(new_n2966_), .B(new_n2968_), .ZN(new_n2969_));
  NOR3_X1    g2917(.A1(new_n1051_), .A2(new_n808_), .A3(new_n1151_), .ZN(new_n2970_));
  NOR3_X1    g2918(.A1(new_n809_), .A2(new_n1050_), .A3(new_n1149_), .ZN(new_n2971_));
  NOR2_X1    g2919(.A1(new_n2971_), .A2(new_n2970_), .ZN(new_n2972_));
  XOR2_X1    g2920(.A1(new_n1050_), .A2(new_n1149_), .Z(new_n2973_));
  XOR2_X1    g2921(.A1(new_n1050_), .A2(new_n802_), .Z(new_n2974_));
  NAND3_X1   g2922(.A1(new_n2968_), .A2(new_n2973_), .A3(new_n2974_), .ZN(new_n2975_));
  OAI22_X1   g2923(.A1(new_n2804_), .A2(new_n2975_), .B1(new_n2765_), .B2(new_n2972_), .ZN(new_n2976_));
  INV_X1     g2924(.I(new_n2969_), .ZN(new_n2977_));
  NAND2_X1   g2925(.A1(new_n2956_), .A2(new_n2977_), .ZN(new_n2978_));
  AOI21_X1   g2926(.A1(new_n2978_), .A2(new_n2976_), .B(new_n803_), .ZN(new_n2979_));
  NOR2_X1    g2927(.A1(new_n2979_), .A2(new_n2969_), .ZN(new_n2980_));
  NAND2_X1   g2928(.A1(new_n2980_), .A2(new_n2964_), .ZN(new_n2981_));
  INV_X1     g2929(.I(new_n2981_), .ZN(new_n2982_));
  NOR2_X1    g2930(.A1(new_n2980_), .A2(new_n2964_), .ZN(new_n2983_));
  NAND2_X1   g2931(.A1(new_n2792_), .A2(new_n2795_), .ZN(new_n2984_));
  OAI21_X1   g2932(.A1(new_n2778_), .A2(new_n2782_), .B(new_n2786_), .ZN(new_n2985_));
  NAND2_X1   g2933(.A1(new_n2984_), .A2(new_n2985_), .ZN(new_n2986_));
  NOR2_X1    g2934(.A1(new_n576_), .A2(new_n803_), .ZN(new_n2987_));
  NOR2_X1    g2935(.A1(new_n577_), .A2(new_n802_), .ZN(new_n2988_));
  XOR2_X1    g2936(.A1(new_n702_), .A2(new_n270_), .Z(new_n2989_));
  INV_X1     g2937(.I(new_n2989_), .ZN(new_n2990_));
  OAI21_X1   g2938(.A1(new_n2987_), .A2(new_n2988_), .B(new_n2990_), .ZN(new_n2991_));
  INV_X1     g2939(.I(new_n2991_), .ZN(new_n2992_));
  NOR3_X1    g2940(.A1(new_n271_), .A2(new_n576_), .A3(new_n803_), .ZN(new_n2993_));
  AOI21_X1   g2941(.A1(new_n271_), .A2(new_n2988_), .B(new_n2993_), .ZN(new_n2994_));
  NOR2_X1    g2942(.A1(new_n2792_), .A2(new_n2994_), .ZN(new_n2995_));
  XOR2_X1    g2943(.A1(new_n270_), .A2(new_n803_), .Z(new_n2996_));
  XOR2_X1    g2944(.A1(new_n702_), .A2(new_n576_), .Z(new_n2997_));
  NOR2_X1    g2945(.A1(new_n2997_), .A2(new_n2996_), .ZN(new_n2998_));
  AOI21_X1   g2946(.A1(new_n2786_), .A2(new_n2998_), .B(new_n702_), .ZN(new_n2999_));
  INV_X1     g2947(.I(new_n2999_), .ZN(new_n3000_));
  OAI21_X1   g2948(.A1(new_n2995_), .A2(new_n3000_), .B(new_n2992_), .ZN(new_n3001_));
  OR2_X2     g2949(.A1(new_n3001_), .A2(new_n2986_), .Z(new_n3002_));
  NAND2_X1   g2950(.A1(new_n3001_), .A2(new_n2986_), .ZN(new_n3003_));
  NOR2_X1    g2951(.A1(new_n2786_), .A2(new_n2996_), .ZN(new_n3004_));
  NOR2_X1    g2952(.A1(new_n3004_), .A2(new_n702_), .ZN(new_n3005_));
  INV_X1     g2953(.I(new_n3005_), .ZN(new_n3006_));
  AOI21_X1   g2954(.A1(new_n3002_), .A2(new_n3003_), .B(new_n3006_), .ZN(new_n3007_));
  NOR2_X1    g2955(.A1(new_n2434_), .A2(new_n2424_), .ZN(new_n3008_));
  INV_X1     g2956(.I(new_n3008_), .ZN(new_n3009_));
  NOR2_X1    g2957(.A1(new_n2465_), .A2(new_n2423_), .ZN(new_n3010_));
  NOR2_X1    g2958(.A1(new_n2402_), .A2(new_n2466_), .ZN(new_n3011_));
  OAI21_X1   g2959(.A1(new_n3010_), .A2(new_n3011_), .B(new_n2795_), .ZN(new_n3012_));
  NAND3_X1   g2960(.A1(new_n2786_), .A2(new_n2781_), .A3(new_n2780_), .ZN(new_n3013_));
  AOI21_X1   g2961(.A1(new_n3012_), .A2(new_n3013_), .B(new_n2776_), .ZN(new_n3014_));
  NAND2_X1   g2962(.A1(new_n3014_), .A2(new_n2760_), .ZN(new_n3015_));
  AOI21_X1   g2963(.A1(new_n2780_), .A2(new_n2781_), .B(new_n2786_), .ZN(new_n3016_));
  NOR3_X1    g2964(.A1(new_n2795_), .A2(new_n3010_), .A3(new_n3011_), .ZN(new_n3017_));
  OAI21_X1   g2965(.A1(new_n3016_), .A2(new_n3017_), .B(new_n2779_), .ZN(new_n3018_));
  NAND2_X1   g2966(.A1(new_n3018_), .A2(new_n2461_), .ZN(new_n3019_));
  AOI21_X1   g2967(.A1(new_n3015_), .A2(new_n3019_), .B(new_n3009_), .ZN(new_n3020_));
  NOR2_X1    g2968(.A1(new_n3018_), .A2(new_n2461_), .ZN(new_n3021_));
  NOR2_X1    g2969(.A1(new_n3014_), .A2(new_n2760_), .ZN(new_n3022_));
  NOR3_X1    g2970(.A1(new_n3022_), .A2(new_n3021_), .A3(new_n3008_), .ZN(new_n3023_));
  OAI21_X1   g2971(.A1(new_n3020_), .A2(new_n3023_), .B(new_n2455_), .ZN(new_n3024_));
  OAI21_X1   g2972(.A1(new_n3022_), .A2(new_n3021_), .B(new_n3008_), .ZN(new_n3025_));
  NAND3_X1   g2973(.A1(new_n3015_), .A2(new_n3019_), .A3(new_n3009_), .ZN(new_n3026_));
  NAND3_X1   g2974(.A1(new_n3025_), .A2(new_n3026_), .A3(new_n2456_), .ZN(new_n3027_));
  INV_X1     g2975(.I(new_n2998_), .ZN(new_n3028_));
  XOR2_X1    g2976(.A1(new_n702_), .A2(new_n802_), .Z(new_n3029_));
  NOR3_X1    g2977(.A1(new_n2989_), .A2(new_n2997_), .A3(new_n3029_), .ZN(new_n3030_));
  INV_X1     g2978(.I(new_n3030_), .ZN(new_n3031_));
  OAI22_X1   g2979(.A1(new_n2792_), .A2(new_n3031_), .B1(new_n2795_), .B2(new_n2994_), .ZN(new_n3032_));
  OAI21_X1   g2980(.A1(new_n2775_), .A2(new_n3028_), .B(new_n3032_), .ZN(new_n3033_));
  AOI21_X1   g2981(.A1(new_n3033_), .A2(new_n721_), .B(new_n2991_), .ZN(new_n3034_));
  NAND3_X1   g2982(.A1(new_n3034_), .A2(new_n3024_), .A3(new_n3027_), .ZN(new_n3035_));
  AOI21_X1   g2983(.A1(new_n3025_), .A2(new_n3026_), .B(new_n2456_), .ZN(new_n3036_));
  NOR3_X1    g2984(.A1(new_n3020_), .A2(new_n3023_), .A3(new_n2455_), .ZN(new_n3037_));
  INV_X1     g2985(.I(new_n2994_), .ZN(new_n3038_));
  AOI22_X1   g2986(.A1(new_n2783_), .A2(new_n3030_), .B1(new_n2786_), .B2(new_n3038_), .ZN(new_n3039_));
  NOR3_X1    g2987(.A1(new_n2766_), .A2(new_n2769_), .A3(new_n3028_), .ZN(new_n3040_));
  OAI21_X1   g2988(.A1(new_n3039_), .A2(new_n3040_), .B(new_n721_), .ZN(new_n3041_));
  NAND2_X1   g2989(.A1(new_n3041_), .A2(new_n2992_), .ZN(new_n3042_));
  OAI21_X1   g2990(.A1(new_n3036_), .A2(new_n3037_), .B(new_n3042_), .ZN(new_n3043_));
  NAND2_X1   g2991(.A1(new_n3043_), .A2(new_n3035_), .ZN(new_n3044_));
  XNOR2_X1   g2992(.A1(new_n3044_), .A2(new_n3007_), .ZN(new_n3045_));
  OAI21_X1   g2993(.A1(new_n2982_), .A2(new_n2983_), .B(new_n3045_), .ZN(new_n3046_));
  NAND3_X1   g2994(.A1(new_n2775_), .A2(new_n2792_), .A3(new_n2795_), .ZN(new_n3047_));
  NAND2_X1   g2995(.A1(new_n2770_), .A2(new_n2783_), .ZN(new_n3048_));
  NAND2_X1   g2996(.A1(new_n3047_), .A2(new_n3048_), .ZN(new_n3049_));
  OAI21_X1   g2997(.A1(new_n2802_), .A2(new_n2803_), .B(new_n2787_), .ZN(new_n3050_));
  NAND3_X1   g2998(.A1(new_n2798_), .A2(new_n2750_), .A3(new_n2757_), .ZN(new_n3051_));
  NAND2_X1   g2999(.A1(new_n3050_), .A2(new_n3051_), .ZN(new_n3052_));
  NAND3_X1   g3000(.A1(new_n3052_), .A2(new_n2765_), .A3(new_n3049_), .ZN(new_n3053_));
  AOI21_X1   g3001(.A1(new_n2750_), .A2(new_n2757_), .B(new_n2798_), .ZN(new_n3054_));
  NOR3_X1    g3002(.A1(new_n2787_), .A2(new_n2803_), .A3(new_n2802_), .ZN(new_n3055_));
  OAI21_X1   g3003(.A1(new_n3054_), .A2(new_n3055_), .B(new_n3049_), .ZN(new_n3056_));
  NAND2_X1   g3004(.A1(new_n3056_), .A2(new_n2791_), .ZN(new_n3057_));
  NAND2_X1   g3005(.A1(new_n3057_), .A2(new_n3053_), .ZN(new_n3058_));
  OAI22_X1   g3006(.A1(new_n2765_), .A2(new_n2975_), .B1(new_n2770_), .B2(new_n2972_), .ZN(new_n3059_));
  OAI21_X1   g3007(.A1(new_n2804_), .A2(new_n2969_), .B(new_n3059_), .ZN(new_n3060_));
  AOI21_X1   g3008(.A1(new_n3060_), .A2(new_n802_), .B(new_n2969_), .ZN(new_n3061_));
  INV_X1     g3009(.I(new_n3061_), .ZN(new_n3062_));
  NOR2_X1    g3010(.A1(new_n3058_), .A2(new_n3062_), .ZN(new_n3063_));
  NOR2_X1    g3011(.A1(new_n3056_), .A2(new_n2791_), .ZN(new_n3064_));
  AOI21_X1   g3012(.A1(new_n3052_), .A2(new_n3049_), .B(new_n2765_), .ZN(new_n3065_));
  NOR2_X1    g3013(.A1(new_n3064_), .A2(new_n3065_), .ZN(new_n3066_));
  NOR2_X1    g3014(.A1(new_n3066_), .A2(new_n3061_), .ZN(new_n3067_));
  NOR2_X1    g3015(.A1(new_n3063_), .A2(new_n3067_), .ZN(new_n3068_));
  NAND2_X1   g3016(.A1(new_n3002_), .A2(new_n3003_), .ZN(new_n3069_));
  XOR2_X1    g3017(.A1(new_n3069_), .A2(new_n3006_), .Z(new_n3070_));
  NAND2_X1   g3018(.A1(new_n3068_), .A2(new_n3070_), .ZN(new_n3071_));
  INV_X1     g3019(.I(new_n3071_), .ZN(new_n3072_));
  AOI21_X1   g3020(.A1(new_n3047_), .A2(new_n3048_), .B(new_n2765_), .ZN(new_n3073_));
  OAI22_X1   g3021(.A1(new_n2783_), .A2(new_n2786_), .B1(new_n2766_), .B2(new_n2769_), .ZN(new_n3074_));
  AOI21_X1   g3022(.A1(new_n2796_), .A2(new_n3074_), .B(new_n2791_), .ZN(new_n3075_));
  INV_X1     g3023(.I(new_n2972_), .ZN(new_n3076_));
  NAND2_X1   g3024(.A1(new_n2783_), .A2(new_n3076_), .ZN(new_n3077_));
  OAI21_X1   g3025(.A1(new_n2770_), .A2(new_n2975_), .B(new_n3077_), .ZN(new_n3078_));
  NAND2_X1   g3026(.A1(new_n2791_), .A2(new_n2977_), .ZN(new_n3079_));
  AOI21_X1   g3027(.A1(new_n3079_), .A2(new_n3078_), .B(new_n803_), .ZN(new_n3080_));
  NOR4_X1    g3028(.A1(new_n3080_), .A2(new_n2969_), .A3(new_n3073_), .A4(new_n3075_), .ZN(new_n3081_));
  INV_X1     g3029(.I(new_n3081_), .ZN(new_n3082_));
  OAI22_X1   g3030(.A1(new_n3080_), .A2(new_n2969_), .B1(new_n3073_), .B2(new_n3075_), .ZN(new_n3083_));
  NAND2_X1   g3031(.A1(new_n3082_), .A2(new_n3083_), .ZN(new_n3084_));
  NOR2_X1    g3032(.A1(new_n3037_), .A2(new_n3036_), .ZN(new_n3085_));
  INV_X1     g3033(.I(new_n2975_), .ZN(new_n3086_));
  AOI22_X1   g3034(.A1(new_n2783_), .A2(new_n3086_), .B1(new_n2786_), .B2(new_n3076_), .ZN(new_n3087_));
  NOR2_X1    g3035(.A1(new_n2775_), .A2(new_n2969_), .ZN(new_n3088_));
  OAI21_X1   g3036(.A1(new_n3088_), .A2(new_n3087_), .B(new_n802_), .ZN(new_n3089_));
  NAND2_X1   g3037(.A1(new_n3089_), .A2(new_n2977_), .ZN(new_n3090_));
  INV_X1     g3038(.I(new_n3090_), .ZN(new_n3091_));
  NAND2_X1   g3039(.A1(new_n3091_), .A2(new_n3085_), .ZN(new_n3092_));
  INV_X1     g3040(.I(new_n3092_), .ZN(new_n3093_));
  NOR2_X1    g3041(.A1(new_n3091_), .A2(new_n3085_), .ZN(new_n3094_));
  AND2_X2    g3042(.A1(new_n2984_), .A2(new_n2985_), .Z(new_n3095_));
  AOI21_X1   g3043(.A1(new_n2786_), .A2(new_n2977_), .B(new_n803_), .ZN(new_n3096_));
  NAND2_X1   g3044(.A1(new_n3077_), .A2(new_n3096_), .ZN(new_n3097_));
  AND3_X2    g3045(.A1(new_n3095_), .A2(new_n2977_), .A3(new_n3097_), .Z(new_n3098_));
  AOI21_X1   g3046(.A1(new_n2977_), .A2(new_n3097_), .B(new_n3095_), .ZN(new_n3099_));
  NAND2_X1   g3047(.A1(new_n2795_), .A2(new_n2973_), .ZN(new_n3100_));
  INV_X1     g3048(.I(new_n3100_), .ZN(new_n3101_));
  NOR2_X1    g3049(.A1(new_n3101_), .A2(new_n803_), .ZN(new_n3102_));
  INV_X1     g3050(.I(new_n3102_), .ZN(new_n3103_));
  NOR3_X1    g3051(.A1(new_n3098_), .A2(new_n3099_), .A3(new_n3103_), .ZN(new_n3104_));
  OAI21_X1   g3052(.A1(new_n3093_), .A2(new_n3094_), .B(new_n3104_), .ZN(new_n3105_));
  NAND2_X1   g3053(.A1(new_n3105_), .A2(new_n3004_), .ZN(new_n3106_));
  INV_X1     g3054(.I(new_n3004_), .ZN(new_n3107_));
  INV_X1     g3055(.I(new_n3085_), .ZN(new_n3108_));
  NAND2_X1   g3056(.A1(new_n3108_), .A2(new_n3090_), .ZN(new_n3109_));
  INV_X1     g3057(.I(new_n3104_), .ZN(new_n3110_));
  AOI21_X1   g3058(.A1(new_n3109_), .A2(new_n3092_), .B(new_n3110_), .ZN(new_n3111_));
  NAND2_X1   g3059(.A1(new_n3111_), .A2(new_n3107_), .ZN(new_n3112_));
  AOI21_X1   g3060(.A1(new_n3106_), .A2(new_n3112_), .B(new_n3084_), .ZN(new_n3113_));
  NOR2_X1    g3061(.A1(new_n3105_), .A2(new_n3107_), .ZN(new_n3114_));
  INV_X1     g3062(.I(new_n3070_), .ZN(new_n3115_));
  OAI21_X1   g3063(.A1(new_n3063_), .A2(new_n3067_), .B(new_n3115_), .ZN(new_n3116_));
  INV_X1     g3064(.I(new_n3116_), .ZN(new_n3117_));
  NOR3_X1    g3065(.A1(new_n3117_), .A2(new_n3113_), .A3(new_n3114_), .ZN(new_n3118_));
  INV_X1     g3066(.I(new_n2983_), .ZN(new_n3119_));
  INV_X1     g3067(.I(new_n3045_), .ZN(new_n3120_));
  NAND3_X1   g3068(.A1(new_n3119_), .A2(new_n3120_), .A3(new_n2981_), .ZN(new_n3121_));
  OAI21_X1   g3069(.A1(new_n3118_), .A2(new_n3072_), .B(new_n3121_), .ZN(new_n3122_));
  NAND3_X1   g3070(.A1(new_n2962_), .A2(new_n2743_), .A3(new_n2808_), .ZN(new_n3123_));
  NAND2_X1   g3071(.A1(new_n2956_), .A2(new_n2788_), .ZN(new_n3124_));
  AOI21_X1   g3072(.A1(new_n3123_), .A2(new_n3124_), .B(new_n2734_), .ZN(new_n3125_));
  NAND2_X1   g3073(.A1(new_n2962_), .A2(new_n2956_), .ZN(new_n3126_));
  AOI21_X1   g3074(.A1(new_n2801_), .A2(new_n3126_), .B(new_n2813_), .ZN(new_n3127_));
  NOR2_X1    g3075(.A1(new_n3127_), .A2(new_n3125_), .ZN(new_n3128_));
  OAI22_X1   g3076(.A1(new_n2956_), .A2(new_n2975_), .B1(new_n2804_), .B2(new_n2972_), .ZN(new_n3129_));
  NAND2_X1   g3077(.A1(new_n2734_), .A2(new_n2977_), .ZN(new_n3130_));
  AOI21_X1   g3078(.A1(new_n3130_), .A2(new_n3129_), .B(new_n803_), .ZN(new_n3131_));
  NOR2_X1    g3079(.A1(new_n3131_), .A2(new_n2969_), .ZN(new_n3132_));
  NAND2_X1   g3080(.A1(new_n3132_), .A2(new_n3128_), .ZN(new_n3133_));
  NOR2_X1    g3081(.A1(new_n3132_), .A2(new_n3128_), .ZN(new_n3134_));
  INV_X1     g3082(.I(new_n3134_), .ZN(new_n3135_));
  NOR3_X1    g3083(.A1(new_n3042_), .A2(new_n3037_), .A3(new_n3036_), .ZN(new_n3136_));
  AOI21_X1   g3084(.A1(new_n3024_), .A2(new_n3027_), .B(new_n3034_), .ZN(new_n3137_));
  OAI21_X1   g3085(.A1(new_n3137_), .A2(new_n3136_), .B(new_n3007_), .ZN(new_n3138_));
  NOR3_X1    g3086(.A1(new_n2770_), .A2(new_n2783_), .A3(new_n2786_), .ZN(new_n3139_));
  NOR2_X1    g3087(.A1(new_n2775_), .A2(new_n2792_), .ZN(new_n3140_));
  OAI21_X1   g3088(.A1(new_n3139_), .A2(new_n3140_), .B(new_n2791_), .ZN(new_n3141_));
  INV_X1     g3089(.I(new_n3074_), .ZN(new_n3142_));
  OAI21_X1   g3090(.A1(new_n3142_), .A2(new_n2805_), .B(new_n2765_), .ZN(new_n3143_));
  AOI21_X1   g3091(.A1(new_n2775_), .A2(new_n3030_), .B(new_n2995_), .ZN(new_n3144_));
  NOR2_X1    g3092(.A1(new_n2765_), .A2(new_n3028_), .ZN(new_n3145_));
  OAI21_X1   g3093(.A1(new_n3145_), .A2(new_n3144_), .B(new_n721_), .ZN(new_n3146_));
  NAND4_X1   g3094(.A1(new_n3146_), .A2(new_n2992_), .A3(new_n3141_), .A4(new_n3143_), .ZN(new_n3147_));
  OAI22_X1   g3095(.A1(new_n2770_), .A2(new_n3031_), .B1(new_n2792_), .B2(new_n2994_), .ZN(new_n3148_));
  NAND2_X1   g3096(.A1(new_n2791_), .A2(new_n2998_), .ZN(new_n3149_));
  AOI21_X1   g3097(.A1(new_n3149_), .A2(new_n3148_), .B(new_n702_), .ZN(new_n3150_));
  OAI22_X1   g3098(.A1(new_n3150_), .A2(new_n2991_), .B1(new_n3073_), .B2(new_n3075_), .ZN(new_n3151_));
  NAND2_X1   g3099(.A1(new_n3147_), .A2(new_n3151_), .ZN(new_n3152_));
  XOR2_X1    g3100(.A1(new_n702_), .A2(new_n708_), .Z(new_n3153_));
  NOR2_X1    g3101(.A1(new_n2786_), .A2(new_n3153_), .ZN(new_n3154_));
  INV_X1     g3102(.I(new_n3154_), .ZN(new_n3155_));
  NOR2_X1    g3103(.A1(new_n3152_), .A2(new_n3155_), .ZN(new_n3156_));
  NOR4_X1    g3104(.A1(new_n3150_), .A2(new_n2991_), .A3(new_n3073_), .A4(new_n3075_), .ZN(new_n3157_));
  AOI22_X1   g3105(.A1(new_n3146_), .A2(new_n2992_), .B1(new_n3141_), .B2(new_n3143_), .ZN(new_n3158_));
  NOR2_X1    g3106(.A1(new_n3158_), .A2(new_n3157_), .ZN(new_n3159_));
  NOR2_X1    g3107(.A1(new_n3159_), .A2(new_n3154_), .ZN(new_n3160_));
  NOR2_X1    g3108(.A1(new_n3160_), .A2(new_n3156_), .ZN(new_n3161_));
  NOR2_X1    g3109(.A1(new_n3159_), .A2(new_n3155_), .ZN(new_n3162_));
  NOR2_X1    g3110(.A1(new_n3152_), .A2(new_n3154_), .ZN(new_n3163_));
  OAI21_X1   g3111(.A1(new_n3162_), .A2(new_n3163_), .B(new_n3138_), .ZN(new_n3164_));
  OAI21_X1   g3112(.A1(new_n3138_), .A2(new_n3161_), .B(new_n3164_), .ZN(new_n3165_));
  NAND3_X1   g3113(.A1(new_n3165_), .A2(new_n3135_), .A3(new_n3133_), .ZN(new_n3166_));
  AOI21_X1   g3114(.A1(new_n3133_), .A2(new_n3135_), .B(new_n3165_), .ZN(new_n3167_));
  INV_X1     g3115(.I(new_n3167_), .ZN(new_n3168_));
  AOI22_X1   g3116(.A1(new_n3168_), .A2(new_n3166_), .B1(new_n3122_), .B2(new_n3046_), .ZN(new_n3169_));
  NAND2_X1   g3117(.A1(new_n3122_), .A2(new_n3046_), .ZN(new_n3170_));
  INV_X1     g3118(.I(new_n3138_), .ZN(new_n3171_));
  OAI21_X1   g3119(.A1(new_n3160_), .A2(new_n3156_), .B(new_n3171_), .ZN(new_n3172_));
  AND2_X2    g3120(.A1(new_n3172_), .A2(new_n3164_), .Z(new_n3173_));
  AOI21_X1   g3121(.A1(new_n3133_), .A2(new_n3135_), .B(new_n3173_), .ZN(new_n3174_));
  INV_X1     g3122(.I(new_n3133_), .ZN(new_n3175_));
  NOR3_X1    g3123(.A1(new_n3165_), .A2(new_n3175_), .A3(new_n3134_), .ZN(new_n3176_));
  NOR2_X1    g3124(.A1(new_n3174_), .A2(new_n3176_), .ZN(new_n3177_));
  NOR2_X1    g3125(.A1(new_n3170_), .A2(new_n3177_), .ZN(new_n3178_));
  NOR2_X1    g3126(.A1(new_n3178_), .A2(new_n3169_), .ZN(new_n3179_));
  AOI22_X1   g3127(.A1(new_n2580_), .A2(new_n2563_), .B1(new_n2626_), .B2(new_n2697_), .ZN(new_n3180_));
  AND3_X2    g3128(.A1(new_n2580_), .A2(new_n2563_), .A3(new_n2632_), .Z(new_n3181_));
  NOR2_X1    g3129(.A1(new_n3181_), .A2(new_n3180_), .ZN(new_n3182_));
  NOR2_X1    g3130(.A1(new_n2722_), .A2(new_n2721_), .ZN(new_n3183_));
  NAND3_X1   g3131(.A1(new_n2811_), .A2(new_n3183_), .A3(new_n2816_), .ZN(new_n3184_));
  OAI21_X1   g3132(.A1(new_n2687_), .A2(new_n2689_), .B(new_n2725_), .ZN(new_n3185_));
  NAND3_X1   g3133(.A1(new_n2711_), .A2(new_n2516_), .A3(new_n2723_), .ZN(new_n3186_));
  AOI21_X1   g3134(.A1(new_n3186_), .A2(new_n3185_), .B(new_n2514_), .ZN(new_n3187_));
  INV_X1     g3135(.I(new_n2728_), .ZN(new_n3188_));
  NOR2_X1    g3136(.A1(new_n3187_), .A2(new_n3188_), .ZN(new_n3189_));
  AOI22_X1   g3137(.A1(new_n2962_), .A2(new_n2808_), .B1(new_n2739_), .B2(new_n2742_), .ZN(new_n3190_));
  NOR2_X1    g3138(.A1(new_n3190_), .A2(new_n2813_), .ZN(new_n3191_));
  NAND2_X1   g3139(.A1(new_n3191_), .A2(new_n3189_), .ZN(new_n3192_));
  AOI22_X1   g3140(.A1(new_n2962_), .A2(new_n2956_), .B1(new_n2517_), .B2(new_n2812_), .ZN(new_n3193_));
  NOR2_X1    g3141(.A1(new_n3193_), .A2(new_n3190_), .ZN(new_n3194_));
  NOR3_X1    g3142(.A1(new_n3194_), .A2(new_n3189_), .A3(new_n2734_), .ZN(new_n3195_));
  OAI21_X1   g3143(.A1(new_n3192_), .A2(new_n3195_), .B(new_n2720_), .ZN(new_n3196_));
  AOI21_X1   g3144(.A1(new_n3184_), .A2(new_n3196_), .B(new_n3182_), .ZN(new_n3197_));
  NOR2_X1    g3145(.A1(new_n2810_), .A2(new_n2729_), .ZN(new_n3198_));
  NAND3_X1   g3146(.A1(new_n2720_), .A2(new_n2816_), .A3(new_n3198_), .ZN(new_n3199_));
  NAND4_X1   g3147(.A1(new_n3183_), .A2(new_n2729_), .A3(new_n2813_), .A4(new_n2815_), .ZN(new_n3200_));
  AOI21_X1   g3148(.A1(new_n3200_), .A2(new_n3199_), .B(new_n2701_), .ZN(new_n3201_));
  NOR2_X1    g3149(.A1(new_n3197_), .A2(new_n3201_), .ZN(new_n3202_));
  NOR2_X1    g3150(.A1(new_n2943_), .A2(new_n1060_), .ZN(new_n3203_));
  NOR2_X1    g3151(.A1(new_n1061_), .A2(new_n2942_), .ZN(new_n3204_));
  XOR2_X1    g3152(.A1(new_n1050_), .A2(new_n1122_), .Z(new_n3205_));
  INV_X1     g3153(.I(new_n3205_), .ZN(new_n3206_));
  OAI21_X1   g3154(.A1(new_n3203_), .A2(new_n3204_), .B(new_n3206_), .ZN(new_n3207_));
  XOR2_X1    g3155(.A1(new_n1050_), .A2(new_n1061_), .Z(new_n3208_));
  XOR2_X1    g3156(.A1(new_n1050_), .A2(new_n2943_), .Z(new_n3209_));
  NOR3_X1    g3157(.A1(new_n3205_), .A2(new_n3208_), .A3(new_n3209_), .ZN(new_n3210_));
  INV_X1     g3158(.I(new_n3210_), .ZN(new_n3211_));
  NOR3_X1    g3159(.A1(new_n1061_), .A2(new_n1121_), .A3(new_n2942_), .ZN(new_n3212_));
  AOI21_X1   g3160(.A1(new_n1121_), .A2(new_n3203_), .B(new_n3212_), .ZN(new_n3213_));
  OAI22_X1   g3161(.A1(new_n3183_), .A2(new_n3211_), .B1(new_n3189_), .B2(new_n3213_), .ZN(new_n3214_));
  XOR2_X1    g3162(.A1(new_n1121_), .A2(new_n2943_), .Z(new_n3215_));
  NOR2_X1    g3163(.A1(new_n3208_), .A2(new_n3215_), .ZN(new_n3216_));
  NAND2_X1   g3164(.A1(new_n3182_), .A2(new_n3216_), .ZN(new_n3217_));
  AOI21_X1   g3165(.A1(new_n3217_), .A2(new_n3214_), .B(new_n1051_), .ZN(new_n3218_));
  NOR2_X1    g3166(.A1(new_n3218_), .A2(new_n3207_), .ZN(new_n3219_));
  NAND2_X1   g3167(.A1(new_n3219_), .A2(new_n3202_), .ZN(new_n3220_));
  OAI22_X1   g3168(.A1(new_n3218_), .A2(new_n3207_), .B1(new_n3197_), .B2(new_n3201_), .ZN(new_n3221_));
  NAND2_X1   g3169(.A1(new_n3220_), .A2(new_n3221_), .ZN(new_n3222_));
  NAND2_X1   g3170(.A1(new_n3179_), .A2(new_n3222_), .ZN(new_n3223_));
  NAND3_X1   g3171(.A1(new_n2813_), .A2(new_n2956_), .A3(new_n2962_), .ZN(new_n3224_));
  NAND2_X1   g3172(.A1(new_n3190_), .A2(new_n2734_), .ZN(new_n3225_));
  NAND2_X1   g3173(.A1(new_n3225_), .A2(new_n3224_), .ZN(new_n3226_));
  OAI21_X1   g3174(.A1(new_n2722_), .A2(new_n2721_), .B(new_n3194_), .ZN(new_n3227_));
  NAND3_X1   g3175(.A1(new_n2715_), .A2(new_n2719_), .A3(new_n2815_), .ZN(new_n3228_));
  NAND2_X1   g3176(.A1(new_n3227_), .A2(new_n3228_), .ZN(new_n3229_));
  NAND3_X1   g3177(.A1(new_n3229_), .A2(new_n3189_), .A3(new_n3226_), .ZN(new_n3230_));
  AOI21_X1   g3178(.A1(new_n2715_), .A2(new_n2719_), .B(new_n2815_), .ZN(new_n3231_));
  NOR3_X1    g3179(.A1(new_n2722_), .A2(new_n2721_), .A3(new_n3194_), .ZN(new_n3232_));
  OAI21_X1   g3180(.A1(new_n3232_), .A2(new_n3231_), .B(new_n3226_), .ZN(new_n3233_));
  NAND2_X1   g3181(.A1(new_n3233_), .A2(new_n2729_), .ZN(new_n3234_));
  NAND2_X1   g3182(.A1(new_n3234_), .A2(new_n3230_), .ZN(new_n3235_));
  INV_X1     g3183(.I(new_n3235_), .ZN(new_n3236_));
  INV_X1     g3184(.I(new_n3216_), .ZN(new_n3237_));
  OAI22_X1   g3185(.A1(new_n3183_), .A2(new_n3211_), .B1(new_n2734_), .B2(new_n3237_), .ZN(new_n3238_));
  OAI21_X1   g3186(.A1(new_n2729_), .A2(new_n3213_), .B(new_n3238_), .ZN(new_n3239_));
  AOI21_X1   g3187(.A1(new_n3239_), .A2(new_n1050_), .B(new_n3207_), .ZN(new_n3240_));
  NAND2_X1   g3188(.A1(new_n3236_), .A2(new_n3240_), .ZN(new_n3241_));
  NOR2_X1    g3189(.A1(new_n3236_), .A2(new_n3240_), .ZN(new_n3242_));
  INV_X1     g3190(.I(new_n3242_), .ZN(new_n3243_));
  NOR2_X1    g3191(.A1(new_n3118_), .A2(new_n3072_), .ZN(new_n3244_));
  INV_X1     g3192(.I(new_n3046_), .ZN(new_n3245_));
  NOR3_X1    g3193(.A1(new_n2982_), .A2(new_n2983_), .A3(new_n3045_), .ZN(new_n3246_));
  NOR2_X1    g3194(.A1(new_n3245_), .A2(new_n3246_), .ZN(new_n3247_));
  OAI21_X1   g3195(.A1(new_n2982_), .A2(new_n2983_), .B(new_n3120_), .ZN(new_n3248_));
  NAND3_X1   g3196(.A1(new_n3119_), .A2(new_n2981_), .A3(new_n3045_), .ZN(new_n3249_));
  NAND2_X1   g3197(.A1(new_n3248_), .A2(new_n3249_), .ZN(new_n3250_));
  NAND2_X1   g3198(.A1(new_n3244_), .A2(new_n3250_), .ZN(new_n3251_));
  OAI21_X1   g3199(.A1(new_n3244_), .A2(new_n3247_), .B(new_n3251_), .ZN(new_n3252_));
  NAND3_X1   g3200(.A1(new_n3252_), .A2(new_n3243_), .A3(new_n3241_), .ZN(new_n3253_));
  INV_X1     g3201(.I(new_n3241_), .ZN(new_n3254_));
  INV_X1     g3202(.I(new_n3083_), .ZN(new_n3255_));
  NOR2_X1    g3203(.A1(new_n3255_), .A2(new_n3081_), .ZN(new_n3256_));
  NOR2_X1    g3204(.A1(new_n3111_), .A2(new_n3107_), .ZN(new_n3257_));
  NOR2_X1    g3205(.A1(new_n3105_), .A2(new_n3004_), .ZN(new_n3258_));
  OAI21_X1   g3206(.A1(new_n3258_), .A2(new_n3257_), .B(new_n3256_), .ZN(new_n3259_));
  INV_X1     g3207(.I(new_n3114_), .ZN(new_n3260_));
  NAND3_X1   g3208(.A1(new_n3259_), .A2(new_n3260_), .A3(new_n3116_), .ZN(new_n3261_));
  AOI22_X1   g3209(.A1(new_n3261_), .A2(new_n3071_), .B1(new_n3046_), .B2(new_n3121_), .ZN(new_n3262_));
  AOI21_X1   g3210(.A1(new_n3244_), .A2(new_n3250_), .B(new_n3262_), .ZN(new_n3263_));
  OAI21_X1   g3211(.A1(new_n3254_), .A2(new_n3242_), .B(new_n3263_), .ZN(new_n3264_));
  NAND2_X1   g3212(.A1(new_n3253_), .A2(new_n3264_), .ZN(new_n3265_));
  AOI21_X1   g3213(.A1(new_n3225_), .A2(new_n3224_), .B(new_n3189_), .ZN(new_n3266_));
  AOI21_X1   g3214(.A1(new_n2956_), .A2(new_n2962_), .B(new_n2734_), .ZN(new_n3267_));
  OAI21_X1   g3215(.A1(new_n3191_), .A2(new_n3267_), .B(new_n3189_), .ZN(new_n3268_));
  INV_X1     g3216(.I(new_n3268_), .ZN(new_n3269_));
  NOR2_X1    g3217(.A1(new_n3269_), .A2(new_n3266_), .ZN(new_n3270_));
  OAI22_X1   g3218(.A1(new_n2734_), .A2(new_n3211_), .B1(new_n2956_), .B2(new_n3213_), .ZN(new_n3271_));
  OAI21_X1   g3219(.A1(new_n2729_), .A2(new_n3237_), .B(new_n3271_), .ZN(new_n3272_));
  AOI21_X1   g3220(.A1(new_n3272_), .A2(new_n1050_), .B(new_n3207_), .ZN(new_n3273_));
  XOR2_X1    g3221(.A1(new_n3270_), .A2(new_n3273_), .Z(new_n3274_));
  NOR3_X1    g3222(.A1(new_n2956_), .A2(new_n2788_), .A3(new_n2800_), .ZN(new_n3275_));
  NOR2_X1    g3223(.A1(new_n2962_), .A2(new_n2743_), .ZN(new_n3276_));
  OAI21_X1   g3224(.A1(new_n3275_), .A2(new_n3276_), .B(new_n2813_), .ZN(new_n3277_));
  OAI21_X1   g3225(.A1(new_n3190_), .A2(new_n2809_), .B(new_n2734_), .ZN(new_n3278_));
  NAND2_X1   g3226(.A1(new_n3278_), .A2(new_n3277_), .ZN(new_n3279_));
  INV_X1     g3227(.I(new_n3207_), .ZN(new_n3280_));
  NOR2_X1    g3228(.A1(new_n2956_), .A2(new_n2804_), .ZN(new_n3281_));
  NOR2_X1    g3229(.A1(new_n3211_), .A2(new_n3213_), .ZN(new_n3282_));
  OAI22_X1   g3230(.A1(new_n3281_), .A2(new_n3282_), .B1(new_n2813_), .B2(new_n3237_), .ZN(new_n3283_));
  NAND2_X1   g3231(.A1(new_n3283_), .A2(new_n1050_), .ZN(new_n3284_));
  NAND2_X1   g3232(.A1(new_n3284_), .A2(new_n3280_), .ZN(new_n3285_));
  NOR2_X1    g3233(.A1(new_n3285_), .A2(new_n3279_), .ZN(new_n3286_));
  NAND2_X1   g3234(.A1(new_n3285_), .A2(new_n3279_), .ZN(new_n3287_));
  INV_X1     g3235(.I(new_n3287_), .ZN(new_n3288_));
  NOR2_X1    g3236(.A1(new_n3288_), .A2(new_n3286_), .ZN(new_n3289_));
  NAND2_X1   g3237(.A1(new_n3084_), .A2(new_n3004_), .ZN(new_n3290_));
  NAND2_X1   g3238(.A1(new_n3256_), .A2(new_n3107_), .ZN(new_n3291_));
  AOI21_X1   g3239(.A1(new_n3291_), .A2(new_n3290_), .B(new_n3105_), .ZN(new_n3292_));
  NAND2_X1   g3240(.A1(new_n3256_), .A2(new_n3004_), .ZN(new_n3293_));
  NAND2_X1   g3241(.A1(new_n3084_), .A2(new_n3107_), .ZN(new_n3294_));
  AOI21_X1   g3242(.A1(new_n3293_), .A2(new_n3294_), .B(new_n3111_), .ZN(new_n3295_));
  NOR2_X1    g3243(.A1(new_n3295_), .A2(new_n3292_), .ZN(new_n3296_));
  INV_X1     g3244(.I(new_n3296_), .ZN(new_n3297_));
  NAND2_X1   g3245(.A1(new_n3289_), .A2(new_n3297_), .ZN(new_n3298_));
  NAND2_X1   g3246(.A1(new_n2758_), .A2(new_n2791_), .ZN(new_n3299_));
  OAI21_X1   g3247(.A1(new_n3211_), .A2(new_n3213_), .B(new_n3299_), .ZN(new_n3300_));
  NAND2_X1   g3248(.A1(new_n2956_), .A2(new_n3216_), .ZN(new_n3301_));
  NAND2_X1   g3249(.A1(new_n3301_), .A2(new_n3300_), .ZN(new_n3302_));
  AOI21_X1   g3250(.A1(new_n3302_), .A2(new_n1050_), .B(new_n3207_), .ZN(new_n3303_));
  XOR2_X1    g3251(.A1(new_n3303_), .A2(new_n2964_), .Z(new_n3304_));
  NOR2_X1    g3252(.A1(new_n3098_), .A2(new_n3099_), .ZN(new_n3305_));
  XOR2_X1    g3253(.A1(new_n3305_), .A2(new_n3103_), .Z(new_n3306_));
  INV_X1     g3254(.I(new_n3306_), .ZN(new_n3307_));
  INV_X1     g3255(.I(new_n3213_), .ZN(new_n3308_));
  OAI21_X1   g3256(.A1(new_n2778_), .A2(new_n2782_), .B(new_n3308_), .ZN(new_n3309_));
  AOI21_X1   g3257(.A1(new_n2786_), .A2(new_n3216_), .B(new_n1051_), .ZN(new_n3310_));
  AOI21_X1   g3258(.A1(new_n3309_), .A2(new_n3310_), .B(new_n3207_), .ZN(new_n3311_));
  INV_X1     g3259(.I(new_n3311_), .ZN(new_n3312_));
  NOR2_X1    g3260(.A1(new_n3312_), .A2(new_n2986_), .ZN(new_n3313_));
  NOR2_X1    g3261(.A1(new_n3095_), .A2(new_n3311_), .ZN(new_n3314_));
  NOR2_X1    g3262(.A1(new_n2786_), .A2(new_n3215_), .ZN(new_n3315_));
  NOR2_X1    g3263(.A1(new_n3315_), .A2(new_n1051_), .ZN(new_n3316_));
  OAI21_X1   g3264(.A1(new_n3314_), .A2(new_n3313_), .B(new_n3316_), .ZN(new_n3317_));
  AOI22_X1   g3265(.A1(new_n2783_), .A2(new_n3210_), .B1(new_n2786_), .B2(new_n3308_), .ZN(new_n3318_));
  NOR2_X1    g3266(.A1(new_n2775_), .A2(new_n3237_), .ZN(new_n3319_));
  OAI21_X1   g3267(.A1(new_n3319_), .A2(new_n3318_), .B(new_n1050_), .ZN(new_n3320_));
  NAND3_X1   g3268(.A1(new_n3085_), .A2(new_n3280_), .A3(new_n3320_), .ZN(new_n3321_));
  AOI22_X1   g3269(.A1(new_n3280_), .A2(new_n3320_), .B1(new_n3024_), .B2(new_n3027_), .ZN(new_n3322_));
  INV_X1     g3270(.I(new_n3322_), .ZN(new_n3323_));
  AOI21_X1   g3271(.A1(new_n3323_), .A2(new_n3321_), .B(new_n3317_), .ZN(new_n3324_));
  NAND2_X1   g3272(.A1(new_n3320_), .A2(new_n3280_), .ZN(new_n3325_));
  NOR3_X1    g3273(.A1(new_n3325_), .A2(new_n3036_), .A3(new_n3037_), .ZN(new_n3326_));
  NOR2_X1    g3274(.A1(new_n3317_), .A2(new_n3100_), .ZN(new_n3327_));
  OAI21_X1   g3275(.A1(new_n3326_), .A2(new_n3322_), .B(new_n3327_), .ZN(new_n3328_));
  OAI21_X1   g3276(.A1(new_n3324_), .A2(new_n3101_), .B(new_n3328_), .ZN(new_n3329_));
  OAI21_X1   g3277(.A1(new_n2770_), .A2(new_n3211_), .B(new_n3309_), .ZN(new_n3330_));
  NAND2_X1   g3278(.A1(new_n2791_), .A2(new_n3216_), .ZN(new_n3331_));
  AOI21_X1   g3279(.A1(new_n3331_), .A2(new_n3330_), .B(new_n1051_), .ZN(new_n3332_));
  NOR4_X1    g3280(.A1(new_n3332_), .A2(new_n3073_), .A3(new_n3075_), .A4(new_n3207_), .ZN(new_n3333_));
  INV_X1     g3281(.I(new_n3332_), .ZN(new_n3334_));
  AOI22_X1   g3282(.A1(new_n3334_), .A2(new_n3280_), .B1(new_n3141_), .B2(new_n3143_), .ZN(new_n3335_));
  NOR2_X1    g3283(.A1(new_n3335_), .A2(new_n3333_), .ZN(new_n3336_));
  NAND2_X1   g3284(.A1(new_n3324_), .A2(new_n3101_), .ZN(new_n3337_));
  OAI21_X1   g3285(.A1(new_n3329_), .A2(new_n3336_), .B(new_n3337_), .ZN(new_n3338_));
  NOR2_X1    g3286(.A1(new_n3338_), .A2(new_n3307_), .ZN(new_n3339_));
  OAI22_X1   g3287(.A1(new_n2765_), .A2(new_n3211_), .B1(new_n2770_), .B2(new_n3213_), .ZN(new_n3340_));
  OAI21_X1   g3288(.A1(new_n2804_), .A2(new_n3237_), .B(new_n3340_), .ZN(new_n3341_));
  AOI21_X1   g3289(.A1(new_n3341_), .A2(new_n1050_), .B(new_n3207_), .ZN(new_n3342_));
  NAND2_X1   g3290(.A1(new_n3066_), .A2(new_n3342_), .ZN(new_n3343_));
  INV_X1     g3291(.I(new_n3342_), .ZN(new_n3344_));
  NAND2_X1   g3292(.A1(new_n3058_), .A2(new_n3344_), .ZN(new_n3345_));
  NAND2_X1   g3293(.A1(new_n3345_), .A2(new_n3343_), .ZN(new_n3346_));
  AOI21_X1   g3294(.A1(new_n3338_), .A2(new_n3307_), .B(new_n3346_), .ZN(new_n3347_));
  NOR2_X1    g3295(.A1(new_n3347_), .A2(new_n3339_), .ZN(new_n3348_));
  NOR2_X1    g3296(.A1(new_n3348_), .A2(new_n3304_), .ZN(new_n3349_));
  NAND2_X1   g3297(.A1(new_n3109_), .A2(new_n3092_), .ZN(new_n3350_));
  XOR2_X1    g3298(.A1(new_n3350_), .A2(new_n3110_), .Z(new_n3351_));
  AOI21_X1   g3299(.A1(new_n3348_), .A2(new_n3304_), .B(new_n3351_), .ZN(new_n3352_));
  OAI22_X1   g3300(.A1(new_n3352_), .A2(new_n3349_), .B1(new_n3289_), .B2(new_n3297_), .ZN(new_n3353_));
  AOI21_X1   g3301(.A1(new_n3353_), .A2(new_n3298_), .B(new_n3274_), .ZN(new_n3354_));
  INV_X1     g3302(.I(new_n3354_), .ZN(new_n3355_));
  NAND3_X1   g3303(.A1(new_n3353_), .A2(new_n3274_), .A3(new_n3298_), .ZN(new_n3356_));
  NOR2_X1    g3304(.A1(new_n3113_), .A2(new_n3114_), .ZN(new_n3357_));
  NAND2_X1   g3305(.A1(new_n3068_), .A2(new_n3115_), .ZN(new_n3358_));
  OAI21_X1   g3306(.A1(new_n3063_), .A2(new_n3067_), .B(new_n3070_), .ZN(new_n3359_));
  NAND2_X1   g3307(.A1(new_n3358_), .A2(new_n3359_), .ZN(new_n3360_));
  XOR2_X1    g3308(.A1(new_n3360_), .A2(new_n3357_), .Z(new_n3361_));
  NAND2_X1   g3309(.A1(new_n3356_), .A2(new_n3361_), .ZN(new_n3362_));
  NAND2_X1   g3310(.A1(new_n3362_), .A2(new_n3355_), .ZN(new_n3363_));
  AOI21_X1   g3311(.A1(new_n3261_), .A2(new_n3071_), .B(new_n3246_), .ZN(new_n3364_));
  NOR3_X1    g3312(.A1(new_n3173_), .A2(new_n3134_), .A3(new_n3175_), .ZN(new_n3365_));
  OAI22_X1   g3313(.A1(new_n3364_), .A2(new_n3245_), .B1(new_n3167_), .B2(new_n3365_), .ZN(new_n3366_));
  OAI21_X1   g3314(.A1(new_n3170_), .A2(new_n3177_), .B(new_n3366_), .ZN(new_n3367_));
  NAND3_X1   g3315(.A1(new_n3367_), .A2(new_n3220_), .A3(new_n3221_), .ZN(new_n3368_));
  AOI21_X1   g3316(.A1(new_n3223_), .A2(new_n3368_), .B(new_n3264_), .ZN(new_n3369_));
  OAI21_X1   g3317(.A1(new_n3369_), .A2(new_n3363_), .B(new_n3265_), .ZN(new_n3370_));
  AOI21_X1   g3318(.A1(new_n3170_), .A2(new_n3168_), .B(new_n3365_), .ZN(new_n3371_));
  INV_X1     g3319(.I(new_n3266_), .ZN(new_n3372_));
  NAND2_X1   g3320(.A1(new_n3372_), .A2(new_n3268_), .ZN(new_n3373_));
  AOI22_X1   g3321(.A1(new_n2813_), .A2(new_n3086_), .B1(new_n2743_), .B2(new_n3076_), .ZN(new_n3374_));
  NOR2_X1    g3322(.A1(new_n2729_), .A2(new_n2969_), .ZN(new_n3375_));
  OAI21_X1   g3323(.A1(new_n3375_), .A2(new_n3374_), .B(new_n802_), .ZN(new_n3376_));
  NAND2_X1   g3324(.A1(new_n3376_), .A2(new_n2977_), .ZN(new_n3377_));
  XOR2_X1    g3325(.A1(new_n3373_), .A2(new_n3377_), .Z(new_n3378_));
  AOI21_X1   g3326(.A1(new_n3044_), .A2(new_n3007_), .B(new_n3155_), .ZN(new_n3379_));
  NOR2_X1    g3327(.A1(new_n3138_), .A2(new_n3154_), .ZN(new_n3380_));
  OAI21_X1   g3328(.A1(new_n3379_), .A2(new_n3380_), .B(new_n3152_), .ZN(new_n3381_));
  NOR2_X1    g3329(.A1(new_n3138_), .A2(new_n3155_), .ZN(new_n3382_));
  INV_X1     g3330(.I(new_n3382_), .ZN(new_n3383_));
  NOR2_X1    g3331(.A1(new_n2770_), .A2(new_n2994_), .ZN(new_n3384_));
  AOI21_X1   g3332(.A1(new_n2791_), .A2(new_n3030_), .B(new_n3384_), .ZN(new_n3385_));
  AOI21_X1   g3333(.A1(new_n2758_), .A2(new_n2998_), .B(new_n3385_), .ZN(new_n3386_));
  OAI21_X1   g3334(.A1(new_n3386_), .A2(new_n702_), .B(new_n2992_), .ZN(new_n3387_));
  NOR3_X1    g3335(.A1(new_n3387_), .A2(new_n3064_), .A3(new_n3065_), .ZN(new_n3388_));
  NOR2_X1    g3336(.A1(new_n2765_), .A2(new_n3031_), .ZN(new_n3389_));
  OAI22_X1   g3337(.A1(new_n2804_), .A2(new_n3028_), .B1(new_n3389_), .B2(new_n3384_), .ZN(new_n3390_));
  AOI21_X1   g3338(.A1(new_n3390_), .A2(new_n721_), .B(new_n2991_), .ZN(new_n3391_));
  AOI21_X1   g3339(.A1(new_n3053_), .A2(new_n3057_), .B(new_n3391_), .ZN(new_n3392_));
  NOR2_X1    g3340(.A1(new_n3153_), .A2(new_n2839_), .ZN(new_n3393_));
  NOR3_X1    g3341(.A1(new_n711_), .A2(new_n645_), .A3(new_n702_), .ZN(new_n3394_));
  NOR3_X1    g3342(.A1(new_n721_), .A2(new_n875_), .A3(new_n708_), .ZN(new_n3395_));
  NOR2_X1    g3343(.A1(new_n3395_), .A2(new_n3394_), .ZN(new_n3396_));
  NOR2_X1    g3344(.A1(new_n2792_), .A2(new_n3396_), .ZN(new_n3397_));
  NOR2_X1    g3345(.A1(new_n3153_), .A2(new_n2838_), .ZN(new_n3398_));
  AOI21_X1   g3346(.A1(new_n2786_), .A2(new_n3398_), .B(new_n438_), .ZN(new_n3399_));
  INV_X1     g3347(.I(new_n3399_), .ZN(new_n3400_));
  OAI21_X1   g3348(.A1(new_n3397_), .A2(new_n3400_), .B(new_n3393_), .ZN(new_n3401_));
  NOR2_X1    g3349(.A1(new_n3401_), .A2(new_n2986_), .ZN(new_n3402_));
  NAND2_X1   g3350(.A1(new_n3401_), .A2(new_n2986_), .ZN(new_n3403_));
  INV_X1     g3351(.I(new_n3403_), .ZN(new_n3404_));
  NOR2_X1    g3352(.A1(new_n3404_), .A2(new_n3402_), .ZN(new_n3405_));
  NOR2_X1    g3353(.A1(new_n3154_), .A2(new_n438_), .ZN(new_n3406_));
  XOR2_X1    g3354(.A1(new_n3405_), .A2(new_n3406_), .Z(new_n3407_));
  OAI21_X1   g3355(.A1(new_n3392_), .A2(new_n3388_), .B(new_n3407_), .ZN(new_n3408_));
  XOR2_X1    g3356(.A1(new_n3408_), .A2(new_n3383_), .Z(new_n3409_));
  NAND2_X1   g3357(.A1(new_n3409_), .A2(new_n3381_), .ZN(new_n3410_));
  NAND2_X1   g3358(.A1(new_n3138_), .A2(new_n3154_), .ZN(new_n3411_));
  NAND3_X1   g3359(.A1(new_n3044_), .A2(new_n3007_), .A3(new_n3155_), .ZN(new_n3412_));
  AOI21_X1   g3360(.A1(new_n3412_), .A2(new_n3411_), .B(new_n3159_), .ZN(new_n3413_));
  XOR2_X1    g3361(.A1(new_n3408_), .A2(new_n3382_), .Z(new_n3414_));
  NAND2_X1   g3362(.A1(new_n3414_), .A2(new_n3413_), .ZN(new_n3415_));
  NAND2_X1   g3363(.A1(new_n3410_), .A2(new_n3415_), .ZN(new_n3416_));
  NAND2_X1   g3364(.A1(new_n3416_), .A2(new_n3378_), .ZN(new_n3417_));
  XOR2_X1    g3365(.A1(new_n3270_), .A2(new_n3377_), .Z(new_n3418_));
  NOR2_X1    g3366(.A1(new_n3414_), .A2(new_n3413_), .ZN(new_n3419_));
  NOR2_X1    g3367(.A1(new_n3409_), .A2(new_n3381_), .ZN(new_n3420_));
  NOR2_X1    g3368(.A1(new_n3419_), .A2(new_n3420_), .ZN(new_n3421_));
  NAND2_X1   g3369(.A1(new_n3421_), .A2(new_n3418_), .ZN(new_n3422_));
  AOI21_X1   g3370(.A1(new_n3417_), .A2(new_n3422_), .B(new_n3371_), .ZN(new_n3423_));
  NAND2_X1   g3371(.A1(new_n3416_), .A2(new_n3418_), .ZN(new_n3424_));
  NAND2_X1   g3372(.A1(new_n3421_), .A2(new_n3378_), .ZN(new_n3425_));
  NAND2_X1   g3373(.A1(new_n3425_), .A2(new_n3424_), .ZN(new_n3426_));
  AOI21_X1   g3374(.A1(new_n3371_), .A2(new_n3426_), .B(new_n3423_), .ZN(new_n3427_));
  NOR3_X1    g3375(.A1(new_n3183_), .A2(new_n3195_), .A3(new_n3192_), .ZN(new_n3428_));
  NOR4_X1    g3376(.A1(new_n2720_), .A2(new_n3189_), .A3(new_n2734_), .A4(new_n3194_), .ZN(new_n3429_));
  NOR2_X1    g3377(.A1(new_n3429_), .A2(new_n3428_), .ZN(new_n3430_));
  XOR2_X1    g3378(.A1(new_n2817_), .A2(new_n2682_), .Z(new_n3431_));
  NOR3_X1    g3379(.A1(new_n3431_), .A2(new_n2701_), .A3(new_n3430_), .ZN(new_n3432_));
  INV_X1     g3380(.I(new_n3430_), .ZN(new_n3433_));
  NAND3_X1   g3381(.A1(new_n2680_), .A2(new_n2580_), .A3(new_n2563_), .ZN(new_n3434_));
  NAND2_X1   g3382(.A1(new_n2678_), .A2(new_n2581_), .ZN(new_n3435_));
  NAND2_X1   g3383(.A1(new_n3435_), .A2(new_n3434_), .ZN(new_n3436_));
  NAND3_X1   g3384(.A1(new_n3436_), .A2(new_n2811_), .A3(new_n2816_), .ZN(new_n3437_));
  NAND2_X1   g3385(.A1(new_n2817_), .A2(new_n2682_), .ZN(new_n3438_));
  NAND2_X1   g3386(.A1(new_n3438_), .A2(new_n3437_), .ZN(new_n3439_));
  AOI21_X1   g3387(.A1(new_n3439_), .A2(new_n3433_), .B(new_n3182_), .ZN(new_n3440_));
  NOR2_X1    g3388(.A1(new_n3432_), .A2(new_n3440_), .ZN(new_n3441_));
  OAI22_X1   g3389(.A1(new_n2682_), .A2(new_n3211_), .B1(new_n3183_), .B2(new_n3237_), .ZN(new_n3442_));
  OAI21_X1   g3390(.A1(new_n2701_), .A2(new_n3213_), .B(new_n3442_), .ZN(new_n3443_));
  AOI21_X1   g3391(.A1(new_n3443_), .A2(new_n1050_), .B(new_n3207_), .ZN(new_n3444_));
  XOR2_X1    g3392(.A1(new_n3441_), .A2(new_n3444_), .Z(new_n3445_));
  NOR2_X1    g3393(.A1(new_n3427_), .A2(new_n3445_), .ZN(new_n3446_));
  NAND2_X1   g3394(.A1(new_n3370_), .A2(new_n3446_), .ZN(new_n3447_));
  AND2_X2    g3395(.A1(new_n3253_), .A2(new_n3264_), .Z(new_n3448_));
  AOI21_X1   g3396(.A1(new_n3361_), .A2(new_n3356_), .B(new_n3354_), .ZN(new_n3449_));
  AOI21_X1   g3397(.A1(new_n3220_), .A2(new_n3221_), .B(new_n3367_), .ZN(new_n3450_));
  AOI21_X1   g3398(.A1(new_n3241_), .A2(new_n3243_), .B(new_n3252_), .ZN(new_n3451_));
  NOR2_X1    g3399(.A1(new_n3179_), .A2(new_n3222_), .ZN(new_n3452_));
  OAI21_X1   g3400(.A1(new_n3450_), .A2(new_n3452_), .B(new_n3451_), .ZN(new_n3453_));
  AOI21_X1   g3401(.A1(new_n3453_), .A2(new_n3449_), .B(new_n3448_), .ZN(new_n3454_));
  NOR2_X1    g3402(.A1(new_n3364_), .A2(new_n3245_), .ZN(new_n3455_));
  OAI21_X1   g3403(.A1(new_n3455_), .A2(new_n3167_), .B(new_n3166_), .ZN(new_n3456_));
  NOR2_X1    g3404(.A1(new_n3421_), .A2(new_n3418_), .ZN(new_n3457_));
  NOR2_X1    g3405(.A1(new_n3416_), .A2(new_n3378_), .ZN(new_n3458_));
  OAI21_X1   g3406(.A1(new_n3457_), .A2(new_n3458_), .B(new_n3456_), .ZN(new_n3459_));
  NAND2_X1   g3407(.A1(new_n3426_), .A2(new_n3371_), .ZN(new_n3460_));
  NAND2_X1   g3408(.A1(new_n3460_), .A2(new_n3459_), .ZN(new_n3461_));
  NAND3_X1   g3409(.A1(new_n3439_), .A2(new_n3433_), .A3(new_n3182_), .ZN(new_n3462_));
  OAI21_X1   g3410(.A1(new_n3431_), .A2(new_n3430_), .B(new_n2701_), .ZN(new_n3463_));
  NAND2_X1   g3411(.A1(new_n3463_), .A2(new_n3462_), .ZN(new_n3464_));
  XOR2_X1    g3412(.A1(new_n3464_), .A2(new_n3444_), .Z(new_n3465_));
  NAND2_X1   g3413(.A1(new_n3461_), .A2(new_n3465_), .ZN(new_n3466_));
  NAND2_X1   g3414(.A1(new_n3454_), .A2(new_n3466_), .ZN(new_n3467_));
  NAND2_X1   g3415(.A1(new_n3467_), .A2(new_n3447_), .ZN(new_n3468_));
  NAND2_X1   g3416(.A1(new_n3468_), .A2(new_n3223_), .ZN(new_n3469_));
  NAND3_X1   g3417(.A1(new_n3467_), .A2(new_n3447_), .A3(new_n3450_), .ZN(new_n3470_));
  NAND2_X1   g3418(.A1(new_n3469_), .A2(new_n3470_), .ZN(new_n3471_));
  INV_X1     g3419(.I(new_n3471_), .ZN(new_n3472_));
  AOI21_X1   g3420(.A1(new_n3427_), .A2(new_n3445_), .B(new_n3223_), .ZN(new_n3473_));
  AOI21_X1   g3421(.A1(new_n3454_), .A2(new_n3473_), .B(new_n3446_), .ZN(new_n3474_));
  OAI21_X1   g3422(.A1(new_n3371_), .A2(new_n3457_), .B(new_n3422_), .ZN(new_n3475_));
  NOR2_X1    g3423(.A1(new_n3233_), .A2(new_n2729_), .ZN(new_n3476_));
  AOI21_X1   g3424(.A1(new_n3229_), .A2(new_n3226_), .B(new_n3189_), .ZN(new_n3477_));
  NOR2_X1    g3425(.A1(new_n2734_), .A2(new_n2969_), .ZN(new_n3478_));
  INV_X1     g3426(.I(new_n3478_), .ZN(new_n3479_));
  OAI21_X1   g3427(.A1(new_n2722_), .A2(new_n2721_), .B(new_n3086_), .ZN(new_n3480_));
  NOR2_X1    g3428(.A1(new_n2729_), .A2(new_n2972_), .ZN(new_n3481_));
  AOI21_X1   g3429(.A1(new_n3480_), .A2(new_n3479_), .B(new_n3481_), .ZN(new_n3482_));
  OAI21_X1   g3430(.A1(new_n3482_), .A2(new_n803_), .B(new_n2977_), .ZN(new_n3483_));
  NOR3_X1    g3431(.A1(new_n3476_), .A2(new_n3483_), .A3(new_n3477_), .ZN(new_n3484_));
  AOI21_X1   g3432(.A1(new_n2720_), .A2(new_n3086_), .B(new_n3478_), .ZN(new_n3485_));
  OAI21_X1   g3433(.A1(new_n3485_), .A2(new_n3481_), .B(new_n802_), .ZN(new_n3486_));
  AOI22_X1   g3434(.A1(new_n3234_), .A2(new_n3230_), .B1(new_n3486_), .B2(new_n2977_), .ZN(new_n3487_));
  NOR2_X1    g3435(.A1(new_n3487_), .A2(new_n3484_), .ZN(new_n3488_));
  NOR2_X1    g3436(.A1(new_n2795_), .A2(new_n3396_), .ZN(new_n3489_));
  INV_X1     g3437(.I(new_n3153_), .ZN(new_n3490_));
  XOR2_X1    g3438(.A1(new_n702_), .A2(new_n875_), .Z(new_n3491_));
  XOR2_X1    g3439(.A1(new_n702_), .A2(new_n438_), .Z(new_n3492_));
  NAND3_X1   g3440(.A1(new_n3490_), .A2(new_n3492_), .A3(new_n3491_), .ZN(new_n3493_));
  INV_X1     g3441(.I(new_n3493_), .ZN(new_n3494_));
  AOI21_X1   g3442(.A1(new_n2783_), .A2(new_n3494_), .B(new_n3489_), .ZN(new_n3495_));
  INV_X1     g3443(.I(new_n3398_), .ZN(new_n3496_));
  NOR3_X1    g3444(.A1(new_n2766_), .A2(new_n2769_), .A3(new_n3496_), .ZN(new_n3497_));
  OAI21_X1   g3445(.A1(new_n3495_), .A2(new_n3497_), .B(new_n437_), .ZN(new_n3498_));
  NAND2_X1   g3446(.A1(new_n3498_), .A2(new_n3393_), .ZN(new_n3499_));
  NOR3_X1    g3447(.A1(new_n3499_), .A2(new_n3036_), .A3(new_n3037_), .ZN(new_n3500_));
  INV_X1     g3448(.I(new_n3393_), .ZN(new_n3501_));
  NOR2_X1    g3449(.A1(new_n2792_), .A2(new_n3493_), .ZN(new_n3502_));
  OAI22_X1   g3450(.A1(new_n2775_), .A2(new_n3496_), .B1(new_n3489_), .B2(new_n3502_), .ZN(new_n3503_));
  AOI21_X1   g3451(.A1(new_n3503_), .A2(new_n437_), .B(new_n3501_), .ZN(new_n3504_));
  AOI21_X1   g3452(.A1(new_n3024_), .A2(new_n3027_), .B(new_n3504_), .ZN(new_n3505_));
  NOR2_X1    g3453(.A1(new_n3505_), .A2(new_n3500_), .ZN(new_n3506_));
  AOI21_X1   g3454(.A1(new_n2799_), .A2(new_n2797_), .B(new_n2804_), .ZN(new_n3507_));
  NOR3_X1    g3455(.A1(new_n2961_), .A2(new_n2807_), .A3(new_n2758_), .ZN(new_n3508_));
  OAI21_X1   g3456(.A1(new_n3508_), .A2(new_n3507_), .B(new_n2743_), .ZN(new_n3509_));
  OAI21_X1   g3457(.A1(new_n2808_), .A2(new_n2788_), .B(new_n2956_), .ZN(new_n3510_));
  NAND2_X1   g3458(.A1(new_n3510_), .A2(new_n3509_), .ZN(new_n3511_));
  NOR2_X1    g3459(.A1(new_n3031_), .A2(new_n2994_), .ZN(new_n3512_));
  INV_X1     g3460(.I(new_n3512_), .ZN(new_n3513_));
  NAND2_X1   g3461(.A1(new_n3299_), .A2(new_n3513_), .ZN(new_n3514_));
  NAND2_X1   g3462(.A1(new_n2956_), .A2(new_n2998_), .ZN(new_n3515_));
  AOI21_X1   g3463(.A1(new_n3515_), .A2(new_n3514_), .B(new_n702_), .ZN(new_n3516_));
  NOR3_X1    g3464(.A1(new_n3511_), .A2(new_n2991_), .A3(new_n3516_), .ZN(new_n3517_));
  NOR2_X1    g3465(.A1(new_n3516_), .A2(new_n2991_), .ZN(new_n3518_));
  NOR2_X1    g3466(.A1(new_n3518_), .A2(new_n2964_), .ZN(new_n3519_));
  NOR2_X1    g3467(.A1(new_n3519_), .A2(new_n3517_), .ZN(new_n3520_));
  INV_X1     g3468(.I(new_n3520_), .ZN(new_n3521_));
  NAND3_X1   g3469(.A1(new_n3391_), .A2(new_n3057_), .A3(new_n3053_), .ZN(new_n3522_));
  OAI21_X1   g3470(.A1(new_n3064_), .A2(new_n3065_), .B(new_n3387_), .ZN(new_n3523_));
  INV_X1     g3471(.I(new_n3406_), .ZN(new_n3524_));
  XOR2_X1    g3472(.A1(new_n3405_), .A2(new_n3524_), .Z(new_n3525_));
  NAND3_X1   g3473(.A1(new_n3523_), .A2(new_n3522_), .A3(new_n3525_), .ZN(new_n3526_));
  NAND3_X1   g3474(.A1(new_n3526_), .A2(new_n3413_), .A3(new_n3382_), .ZN(new_n3527_));
  NOR3_X1    g3475(.A1(new_n3404_), .A2(new_n3402_), .A3(new_n3524_), .ZN(new_n3528_));
  NAND3_X1   g3476(.A1(new_n3527_), .A2(new_n3408_), .A3(new_n3528_), .ZN(new_n3529_));
  INV_X1     g3477(.I(new_n3408_), .ZN(new_n3530_));
  NOR3_X1    g3478(.A1(new_n3392_), .A2(new_n3388_), .A3(new_n3407_), .ZN(new_n3531_));
  NOR3_X1    g3479(.A1(new_n3531_), .A2(new_n3381_), .A3(new_n3383_), .ZN(new_n3532_));
  INV_X1     g3480(.I(new_n3402_), .ZN(new_n3533_));
  NAND3_X1   g3481(.A1(new_n3533_), .A2(new_n3403_), .A3(new_n3406_), .ZN(new_n3534_));
  OAI21_X1   g3482(.A1(new_n3532_), .A2(new_n3530_), .B(new_n3534_), .ZN(new_n3535_));
  AOI21_X1   g3483(.A1(new_n3535_), .A2(new_n3529_), .B(new_n3521_), .ZN(new_n3536_));
  NOR3_X1    g3484(.A1(new_n3532_), .A2(new_n3530_), .A3(new_n3534_), .ZN(new_n3537_));
  AOI21_X1   g3485(.A1(new_n3527_), .A2(new_n3408_), .B(new_n3528_), .ZN(new_n3538_));
  NOR3_X1    g3486(.A1(new_n3537_), .A2(new_n3538_), .A3(new_n3520_), .ZN(new_n3539_));
  OAI21_X1   g3487(.A1(new_n3539_), .A2(new_n3536_), .B(new_n3506_), .ZN(new_n3540_));
  INV_X1     g3488(.I(new_n3506_), .ZN(new_n3541_));
  OAI21_X1   g3489(.A1(new_n3537_), .A2(new_n3538_), .B(new_n3520_), .ZN(new_n3542_));
  NAND3_X1   g3490(.A1(new_n3535_), .A2(new_n3529_), .A3(new_n3521_), .ZN(new_n3543_));
  NAND3_X1   g3491(.A1(new_n3542_), .A2(new_n3543_), .A3(new_n3541_), .ZN(new_n3544_));
  NAND3_X1   g3492(.A1(new_n3488_), .A2(new_n3540_), .A3(new_n3544_), .ZN(new_n3545_));
  NAND4_X1   g3493(.A1(new_n3234_), .A2(new_n3230_), .A3(new_n3486_), .A4(new_n2977_), .ZN(new_n3546_));
  OAI21_X1   g3494(.A1(new_n3476_), .A2(new_n3477_), .B(new_n3483_), .ZN(new_n3547_));
  NAND2_X1   g3495(.A1(new_n3547_), .A2(new_n3546_), .ZN(new_n3548_));
  AOI21_X1   g3496(.A1(new_n3542_), .A2(new_n3543_), .B(new_n3541_), .ZN(new_n3549_));
  NOR3_X1    g3497(.A1(new_n3539_), .A2(new_n3536_), .A3(new_n3506_), .ZN(new_n3550_));
  OAI21_X1   g3498(.A1(new_n3550_), .A2(new_n3549_), .B(new_n3548_), .ZN(new_n3551_));
  NAND2_X1   g3499(.A1(new_n3551_), .A2(new_n3545_), .ZN(new_n3552_));
  NOR2_X1    g3500(.A1(new_n3552_), .A2(new_n3475_), .ZN(new_n3553_));
  AOI21_X1   g3501(.A1(new_n3456_), .A2(new_n3417_), .B(new_n3458_), .ZN(new_n3554_));
  NOR3_X1    g3502(.A1(new_n3549_), .A2(new_n3550_), .A3(new_n3548_), .ZN(new_n3555_));
  AOI21_X1   g3503(.A1(new_n3540_), .A2(new_n3544_), .B(new_n3488_), .ZN(new_n3556_));
  NOR2_X1    g3504(.A1(new_n3556_), .A2(new_n3555_), .ZN(new_n3557_));
  NOR2_X1    g3505(.A1(new_n3557_), .A2(new_n3554_), .ZN(new_n3558_));
  AOI22_X1   g3506(.A1(new_n2715_), .A2(new_n2719_), .B1(new_n3191_), .B2(new_n3189_), .ZN(new_n3559_));
  NOR3_X1    g3507(.A1(new_n3559_), .A2(new_n2720_), .A3(new_n3195_), .ZN(new_n3560_));
  AOI21_X1   g3508(.A1(new_n3560_), .A2(new_n3182_), .B(new_n2682_), .ZN(new_n3561_));
  INV_X1     g3509(.I(new_n3561_), .ZN(new_n3562_));
  NAND3_X1   g3510(.A1(new_n2817_), .A2(new_n2701_), .A3(new_n2720_), .ZN(new_n3563_));
  NAND3_X1   g3511(.A1(new_n2875_), .A2(new_n2878_), .A3(new_n2682_), .ZN(new_n3564_));
  OAI21_X1   g3512(.A1(new_n2930_), .A2(new_n2929_), .B(new_n3436_), .ZN(new_n3565_));
  NAND4_X1   g3513(.A1(new_n3562_), .A2(new_n3565_), .A3(new_n3564_), .A4(new_n3563_), .ZN(new_n3566_));
  INV_X1     g3514(.I(new_n3563_), .ZN(new_n3567_));
  NOR3_X1    g3515(.A1(new_n2930_), .A2(new_n2929_), .A3(new_n3436_), .ZN(new_n3568_));
  AOI21_X1   g3516(.A1(new_n2875_), .A2(new_n2878_), .B(new_n2682_), .ZN(new_n3569_));
  OAI22_X1   g3517(.A1(new_n3568_), .A2(new_n3569_), .B1(new_n3561_), .B2(new_n3567_), .ZN(new_n3570_));
  NAND2_X1   g3518(.A1(new_n3570_), .A2(new_n3566_), .ZN(new_n3571_));
  AOI22_X1   g3519(.A1(new_n3436_), .A2(new_n3210_), .B1(new_n2701_), .B2(new_n3308_), .ZN(new_n3572_));
  NOR2_X1    g3520(.A1(new_n2879_), .A2(new_n3237_), .ZN(new_n3573_));
  OAI21_X1   g3521(.A1(new_n3573_), .A2(new_n3572_), .B(new_n1050_), .ZN(new_n3574_));
  NAND2_X1   g3522(.A1(new_n3574_), .A2(new_n3280_), .ZN(new_n3575_));
  XOR2_X1    g3523(.A1(new_n3575_), .A2(new_n3571_), .Z(new_n3576_));
  NOR3_X1    g3524(.A1(new_n3576_), .A2(new_n3558_), .A3(new_n3553_), .ZN(new_n3577_));
  NAND2_X1   g3525(.A1(new_n3557_), .A2(new_n3554_), .ZN(new_n3578_));
  NAND2_X1   g3526(.A1(new_n3552_), .A2(new_n3475_), .ZN(new_n3579_));
  NOR4_X1    g3527(.A1(new_n3568_), .A2(new_n3569_), .A3(new_n3567_), .A4(new_n3561_), .ZN(new_n3580_));
  AOI22_X1   g3528(.A1(new_n3565_), .A2(new_n3564_), .B1(new_n3562_), .B2(new_n3563_), .ZN(new_n3581_));
  NOR2_X1    g3529(.A1(new_n3581_), .A2(new_n3580_), .ZN(new_n3582_));
  NAND3_X1   g3530(.A1(new_n3582_), .A2(new_n3280_), .A3(new_n3574_), .ZN(new_n3583_));
  NAND2_X1   g3531(.A1(new_n3575_), .A2(new_n3571_), .ZN(new_n3584_));
  NAND2_X1   g3532(.A1(new_n3584_), .A2(new_n3583_), .ZN(new_n3585_));
  AOI21_X1   g3533(.A1(new_n3578_), .A2(new_n3579_), .B(new_n3585_), .ZN(new_n3586_));
  NOR3_X1    g3534(.A1(new_n2879_), .A2(new_n2901_), .A3(new_n2900_), .ZN(new_n3587_));
  AOI21_X1   g3535(.A1(new_n2882_), .A2(new_n3587_), .B(new_n2926_), .ZN(new_n3588_));
  NOR3_X1    g3536(.A1(new_n2882_), .A2(new_n2931_), .A3(new_n2902_), .ZN(new_n3589_));
  NOR4_X1    g3537(.A1(new_n834_), .A2(new_n317_), .A3(new_n329_), .A4(new_n519_), .ZN(new_n3590_));
  NOR4_X1    g3538(.A1(new_n2570_), .A2(new_n820_), .A3(new_n1088_), .A4(new_n852_), .ZN(new_n3591_));
  NAND4_X1   g3539(.A1(new_n3591_), .A2(new_n2437_), .A3(new_n2444_), .A4(new_n3590_), .ZN(new_n3592_));
  NOR3_X1    g3540(.A1(new_n3592_), .A2(new_n226_), .A3(new_n556_), .ZN(new_n3593_));
  NAND2_X1   g3541(.A1(new_n2925_), .A2(new_n3593_), .ZN(new_n3594_));
  NOR3_X1    g3542(.A1(new_n2886_), .A2(new_n2883_), .A3(new_n3594_), .ZN(new_n3595_));
  AOI22_X1   g3543(.A1(new_n2905_), .A2(new_n2904_), .B1(new_n2925_), .B2(new_n3593_), .ZN(new_n3596_));
  NOR2_X1    g3544(.A1(new_n3596_), .A2(new_n3595_), .ZN(new_n3597_));
  NOR2_X1    g3545(.A1(new_n2926_), .A2(new_n3597_), .ZN(new_n3598_));
  NAND2_X1   g3546(.A1(new_n2926_), .A2(new_n3597_), .ZN(new_n3599_));
  INV_X1     g3547(.I(new_n3599_), .ZN(new_n3600_));
  OAI22_X1   g3548(.A1(new_n3589_), .A2(new_n3588_), .B1(new_n3598_), .B2(new_n3600_), .ZN(new_n3601_));
  NAND3_X1   g3549(.A1(new_n2931_), .A2(new_n2896_), .A3(new_n2897_), .ZN(new_n3602_));
  OAI21_X1   g3550(.A1(new_n2932_), .A2(new_n3602_), .B(new_n2946_), .ZN(new_n3603_));
  NAND3_X1   g3551(.A1(new_n2932_), .A2(new_n2898_), .A3(new_n2879_), .ZN(new_n3604_));
  XOR2_X1    g3552(.A1(new_n2926_), .A2(new_n3597_), .Z(new_n3605_));
  NAND3_X1   g3553(.A1(new_n3605_), .A2(new_n3603_), .A3(new_n3604_), .ZN(new_n3606_));
  NAND2_X1   g3554(.A1(new_n3601_), .A2(new_n3606_), .ZN(new_n3607_));
  NAND2_X1   g3555(.A1(new_n2946_), .A2(new_n2947_), .ZN(new_n3608_));
  NAND2_X1   g3556(.A1(new_n2898_), .A2(new_n2949_), .ZN(new_n3609_));
  AOI22_X1   g3557(.A1(new_n3608_), .A2(new_n3609_), .B1(new_n2940_), .B2(new_n3597_), .ZN(new_n3610_));
  INV_X1     g3558(.I(new_n3610_), .ZN(new_n3611_));
  AOI21_X1   g3559(.A1(new_n3607_), .A2(new_n2940_), .B(new_n3611_), .ZN(new_n3612_));
  NOR3_X1    g3560(.A1(new_n3577_), .A2(new_n3586_), .A3(new_n3612_), .ZN(new_n3613_));
  NAND3_X1   g3561(.A1(new_n3585_), .A2(new_n3578_), .A3(new_n3579_), .ZN(new_n3614_));
  OAI21_X1   g3562(.A1(new_n3553_), .A2(new_n3558_), .B(new_n3576_), .ZN(new_n3615_));
  INV_X1     g3563(.I(new_n3598_), .ZN(new_n3616_));
  AOI22_X1   g3564(.A1(new_n3603_), .A2(new_n3604_), .B1(new_n3616_), .B2(new_n3599_), .ZN(new_n3617_));
  NAND2_X1   g3565(.A1(new_n3603_), .A2(new_n3604_), .ZN(new_n3618_));
  XNOR2_X1   g3566(.A1(new_n2926_), .A2(new_n3597_), .ZN(new_n3619_));
  NOR2_X1    g3567(.A1(new_n3618_), .A2(new_n3619_), .ZN(new_n3620_));
  OAI21_X1   g3568(.A1(new_n3620_), .A2(new_n3617_), .B(new_n2940_), .ZN(new_n3621_));
  NAND2_X1   g3569(.A1(new_n3621_), .A2(new_n3610_), .ZN(new_n3622_));
  AOI21_X1   g3570(.A1(new_n3615_), .A2(new_n3614_), .B(new_n3622_), .ZN(new_n3623_));
  OAI21_X1   g3571(.A1(new_n3613_), .A2(new_n3623_), .B(new_n3474_), .ZN(new_n3624_));
  OAI21_X1   g3572(.A1(new_n3461_), .A2(new_n3465_), .B(new_n3450_), .ZN(new_n3625_));
  OAI21_X1   g3573(.A1(new_n3370_), .A2(new_n3625_), .B(new_n3466_), .ZN(new_n3626_));
  NAND3_X1   g3574(.A1(new_n3615_), .A2(new_n3622_), .A3(new_n3614_), .ZN(new_n3627_));
  OAI21_X1   g3575(.A1(new_n3577_), .A2(new_n3586_), .B(new_n3612_), .ZN(new_n3628_));
  NAND3_X1   g3576(.A1(new_n3626_), .A2(new_n3627_), .A3(new_n3628_), .ZN(new_n3629_));
  AOI21_X1   g3577(.A1(new_n3624_), .A2(new_n3629_), .B(new_n2943_), .ZN(new_n3630_));
  AOI21_X1   g3578(.A1(new_n3627_), .A2(new_n3628_), .B(new_n3626_), .ZN(new_n3631_));
  NOR3_X1    g3579(.A1(new_n3474_), .A2(new_n3623_), .A3(new_n3613_), .ZN(new_n3632_));
  NOR3_X1    g3580(.A1(new_n3632_), .A2(new_n3631_), .A3(new_n2942_), .ZN(new_n3633_));
  NOR2_X1    g3581(.A1(new_n3630_), .A2(new_n3633_), .ZN(new_n3634_));
  OAI21_X1   g3582(.A1(new_n3634_), .A2(new_n3472_), .B(new_n2953_), .ZN(new_n3635_));
  INV_X1     g3583(.I(new_n2949_), .ZN(new_n3636_));
  NAND2_X1   g3584(.A1(new_n2720_), .A2(new_n2940_), .ZN(new_n3637_));
  INV_X1     g3585(.I(new_n3637_), .ZN(new_n3638_));
  INV_X1     g3586(.I(new_n2947_), .ZN(new_n3639_));
  NOR2_X1    g3587(.A1(new_n2682_), .A2(new_n3639_), .ZN(new_n3640_));
  OAI22_X1   g3588(.A1(new_n3640_), .A2(new_n3638_), .B1(new_n2701_), .B2(new_n3636_), .ZN(new_n3641_));
  AOI21_X1   g3589(.A1(new_n3641_), .A2(new_n2942_), .B(new_n2939_), .ZN(new_n3642_));
  INV_X1     g3590(.I(new_n3642_), .ZN(new_n3643_));
  NOR2_X1    g3591(.A1(new_n3464_), .A2(new_n3643_), .ZN(new_n3644_));
  NOR2_X1    g3592(.A1(new_n3441_), .A2(new_n3642_), .ZN(new_n3645_));
  NOR2_X1    g3593(.A1(new_n3645_), .A2(new_n3644_), .ZN(new_n3646_));
  INV_X1     g3594(.I(new_n3646_), .ZN(new_n3647_));
  INV_X1     g3595(.I(new_n3357_), .ZN(new_n3648_));
  INV_X1     g3596(.I(new_n3298_), .ZN(new_n3649_));
  INV_X1     g3597(.I(new_n3304_), .ZN(new_n3650_));
  NAND2_X1   g3598(.A1(new_n3323_), .A2(new_n3321_), .ZN(new_n3651_));
  INV_X1     g3599(.I(new_n3317_), .ZN(new_n3652_));
  OAI21_X1   g3600(.A1(new_n3326_), .A2(new_n3322_), .B(new_n3652_), .ZN(new_n3653_));
  AOI22_X1   g3601(.A1(new_n3100_), .A2(new_n3653_), .B1(new_n3651_), .B2(new_n3327_), .ZN(new_n3654_));
  INV_X1     g3602(.I(new_n3336_), .ZN(new_n3655_));
  NOR2_X1    g3603(.A1(new_n3653_), .A2(new_n3100_), .ZN(new_n3656_));
  AOI21_X1   g3604(.A1(new_n3654_), .A2(new_n3655_), .B(new_n3656_), .ZN(new_n3657_));
  NAND2_X1   g3605(.A1(new_n3657_), .A2(new_n3306_), .ZN(new_n3658_));
  NOR2_X1    g3606(.A1(new_n3058_), .A2(new_n3344_), .ZN(new_n3659_));
  NOR2_X1    g3607(.A1(new_n3066_), .A2(new_n3342_), .ZN(new_n3660_));
  NOR2_X1    g3608(.A1(new_n3659_), .A2(new_n3660_), .ZN(new_n3661_));
  OAI21_X1   g3609(.A1(new_n3657_), .A2(new_n3306_), .B(new_n3661_), .ZN(new_n3662_));
  NAND2_X1   g3610(.A1(new_n3662_), .A2(new_n3658_), .ZN(new_n3663_));
  NAND2_X1   g3611(.A1(new_n3663_), .A2(new_n3650_), .ZN(new_n3664_));
  INV_X1     g3612(.I(new_n3351_), .ZN(new_n3665_));
  OAI21_X1   g3613(.A1(new_n3663_), .A2(new_n3650_), .B(new_n3665_), .ZN(new_n3666_));
  NOR2_X1    g3614(.A1(new_n3289_), .A2(new_n3297_), .ZN(new_n3667_));
  AOI21_X1   g3615(.A1(new_n3666_), .A2(new_n3664_), .B(new_n3667_), .ZN(new_n3668_));
  NOR3_X1    g3616(.A1(new_n3668_), .A2(new_n3648_), .A3(new_n3649_), .ZN(new_n3669_));
  AOI21_X1   g3617(.A1(new_n3353_), .A2(new_n3298_), .B(new_n3357_), .ZN(new_n3670_));
  OAI21_X1   g3618(.A1(new_n3669_), .A2(new_n3670_), .B(new_n3274_), .ZN(new_n3671_));
  INV_X1     g3619(.I(new_n3274_), .ZN(new_n3672_));
  NAND3_X1   g3620(.A1(new_n3353_), .A2(new_n3357_), .A3(new_n3298_), .ZN(new_n3673_));
  OAI21_X1   g3621(.A1(new_n3668_), .A2(new_n3649_), .B(new_n3648_), .ZN(new_n3674_));
  NAND3_X1   g3622(.A1(new_n3674_), .A2(new_n3673_), .A3(new_n3672_), .ZN(new_n3675_));
  AOI21_X1   g3623(.A1(new_n3671_), .A2(new_n3675_), .B(new_n3360_), .ZN(new_n3676_));
  INV_X1     g3624(.I(new_n3360_), .ZN(new_n3677_));
  AOI21_X1   g3625(.A1(new_n3674_), .A2(new_n3673_), .B(new_n3672_), .ZN(new_n3678_));
  NOR3_X1    g3626(.A1(new_n3669_), .A2(new_n3670_), .A3(new_n3274_), .ZN(new_n3679_));
  NOR3_X1    g3627(.A1(new_n3679_), .A2(new_n3678_), .A3(new_n3677_), .ZN(new_n3680_));
  NOR3_X1    g3628(.A1(new_n3680_), .A2(new_n3676_), .A3(new_n3647_), .ZN(new_n3681_));
  OAI22_X1   g3629(.A1(new_n2729_), .A2(new_n3636_), .B1(new_n2813_), .B2(new_n3639_), .ZN(new_n3682_));
  NAND3_X1   g3630(.A1(new_n2720_), .A2(new_n3682_), .A3(new_n2940_), .ZN(new_n3683_));
  AOI21_X1   g3631(.A1(new_n3683_), .A2(new_n2942_), .B(new_n2939_), .ZN(new_n3684_));
  NAND3_X1   g3632(.A1(new_n3234_), .A2(new_n3230_), .A3(new_n3684_), .ZN(new_n3685_));
  AOI21_X1   g3633(.A1(new_n3234_), .A2(new_n3230_), .B(new_n3684_), .ZN(new_n3686_));
  INV_X1     g3634(.I(new_n3686_), .ZN(new_n3687_));
  NAND2_X1   g3635(.A1(new_n3687_), .A2(new_n3685_), .ZN(new_n3688_));
  NAND4_X1   g3636(.A1(new_n3338_), .A2(new_n3305_), .A3(new_n3346_), .A4(new_n3102_), .ZN(new_n3689_));
  INV_X1     g3637(.I(new_n3689_), .ZN(new_n3690_));
  AOI21_X1   g3638(.A1(new_n3662_), .A2(new_n3658_), .B(new_n3104_), .ZN(new_n3691_));
  OAI21_X1   g3639(.A1(new_n3691_), .A2(new_n3690_), .B(new_n3304_), .ZN(new_n3692_));
  OAI21_X1   g3640(.A1(new_n3347_), .A2(new_n3339_), .B(new_n3110_), .ZN(new_n3693_));
  NAND3_X1   g3641(.A1(new_n3693_), .A2(new_n3650_), .A3(new_n3689_), .ZN(new_n3694_));
  AOI21_X1   g3642(.A1(new_n3692_), .A2(new_n3694_), .B(new_n3350_), .ZN(new_n3695_));
  INV_X1     g3643(.I(new_n3350_), .ZN(new_n3696_));
  AOI21_X1   g3644(.A1(new_n3693_), .A2(new_n3689_), .B(new_n3650_), .ZN(new_n3697_));
  NOR3_X1    g3645(.A1(new_n3691_), .A2(new_n3690_), .A3(new_n3304_), .ZN(new_n3698_));
  NOR3_X1    g3646(.A1(new_n3698_), .A2(new_n3697_), .A3(new_n3696_), .ZN(new_n3699_));
  NOR3_X1    g3647(.A1(new_n3699_), .A2(new_n3695_), .A3(new_n3688_), .ZN(new_n3700_));
  NAND2_X1   g3648(.A1(new_n2758_), .A2(new_n2940_), .ZN(new_n3701_));
  OAI21_X1   g3649(.A1(new_n2773_), .A2(new_n2772_), .B(new_n3639_), .ZN(new_n3702_));
  NAND3_X1   g3650(.A1(new_n2767_), .A2(new_n2768_), .A3(new_n2947_), .ZN(new_n3703_));
  AOI21_X1   g3651(.A1(new_n3702_), .A2(new_n3703_), .B(new_n2760_), .ZN(new_n3704_));
  AOI21_X1   g3652(.A1(new_n3704_), .A2(new_n2747_), .B(new_n2473_), .ZN(new_n3705_));
  OAI21_X1   g3653(.A1(new_n2747_), .A2(new_n3704_), .B(new_n3705_), .ZN(new_n3706_));
  NAND3_X1   g3654(.A1(new_n3701_), .A2(new_n3706_), .A3(new_n2949_), .ZN(new_n3707_));
  AOI21_X1   g3655(.A1(new_n3707_), .A2(new_n2942_), .B(new_n2939_), .ZN(new_n3708_));
  NAND2_X1   g3656(.A1(new_n3066_), .A2(new_n3708_), .ZN(new_n3709_));
  INV_X1     g3657(.I(new_n3708_), .ZN(new_n3710_));
  NAND2_X1   g3658(.A1(new_n3710_), .A2(new_n3058_), .ZN(new_n3711_));
  NOR2_X1    g3659(.A1(new_n3314_), .A2(new_n3313_), .ZN(new_n3712_));
  XOR2_X1    g3660(.A1(new_n3712_), .A2(new_n3316_), .Z(new_n3713_));
  AOI21_X1   g3661(.A1(new_n3711_), .A2(new_n3709_), .B(new_n3713_), .ZN(new_n3714_));
  NAND3_X1   g3662(.A1(new_n3711_), .A2(new_n3709_), .A3(new_n3713_), .ZN(new_n3715_));
  NOR2_X1    g3663(.A1(new_n2792_), .A2(new_n3636_), .ZN(new_n3716_));
  NOR2_X1    g3664(.A1(new_n2770_), .A2(new_n3639_), .ZN(new_n3717_));
  OAI22_X1   g3665(.A1(new_n2765_), .A2(new_n2939_), .B1(new_n3717_), .B2(new_n3716_), .ZN(new_n3718_));
  AOI22_X1   g3666(.A1(new_n2783_), .A2(new_n2947_), .B1(new_n2786_), .B2(new_n2949_), .ZN(new_n3719_));
  OAI21_X1   g3667(.A1(new_n3719_), .A2(new_n2942_), .B(new_n2939_), .ZN(new_n3720_));
  AOI21_X1   g3668(.A1(new_n2786_), .A2(new_n2943_), .B(\a[0] ), .ZN(new_n3721_));
  NOR4_X1    g3669(.A1(new_n3721_), .A2(new_n2939_), .A3(new_n2943_), .A4(new_n3636_), .ZN(new_n3722_));
  OAI21_X1   g3670(.A1(new_n2783_), .A2(new_n2939_), .B(new_n3722_), .ZN(new_n3723_));
  AOI22_X1   g3671(.A1(new_n3720_), .A2(new_n2775_), .B1(new_n3095_), .B2(new_n3723_), .ZN(new_n3724_));
  NAND2_X1   g3672(.A1(new_n3108_), .A2(new_n3724_), .ZN(new_n3725_));
  NOR2_X1    g3673(.A1(new_n3315_), .A2(new_n2942_), .ZN(new_n3726_));
  NAND3_X1   g3674(.A1(new_n3725_), .A2(new_n3718_), .A3(new_n3726_), .ZN(new_n3727_));
  INV_X1     g3675(.I(new_n3718_), .ZN(new_n3728_));
  INV_X1     g3676(.I(new_n3724_), .ZN(new_n3729_));
  NOR2_X1    g3677(.A1(new_n3729_), .A2(new_n3085_), .ZN(new_n3730_));
  INV_X1     g3678(.I(new_n3726_), .ZN(new_n3731_));
  OAI21_X1   g3679(.A1(new_n3730_), .A2(new_n3731_), .B(new_n3728_), .ZN(new_n3732_));
  XOR2_X1    g3680(.A1(new_n3049_), .A2(new_n2939_), .Z(new_n3733_));
  NAND2_X1   g3681(.A1(new_n2791_), .A2(new_n3315_), .ZN(new_n3734_));
  NOR3_X1    g3682(.A1(new_n3725_), .A2(new_n3733_), .A3(new_n3734_), .ZN(new_n3735_));
  INV_X1     g3683(.I(new_n3735_), .ZN(new_n3736_));
  AOI21_X1   g3684(.A1(new_n3727_), .A2(new_n3732_), .B(new_n3736_), .ZN(new_n3737_));
  AOI21_X1   g3685(.A1(new_n3737_), .A2(new_n3715_), .B(new_n3714_), .ZN(new_n3738_));
  NOR2_X1    g3686(.A1(new_n3639_), .A2(new_n3636_), .ZN(new_n3739_));
  INV_X1     g3687(.I(new_n3739_), .ZN(new_n3740_));
  AOI22_X1   g3688(.A1(new_n2956_), .A2(new_n2940_), .B1(new_n3299_), .B2(new_n3740_), .ZN(new_n3741_));
  NOR2_X1    g3689(.A1(new_n3741_), .A2(new_n2943_), .ZN(new_n3742_));
  NOR2_X1    g3690(.A1(new_n3742_), .A2(new_n2939_), .ZN(new_n3743_));
  XOR2_X1    g3691(.A1(new_n3743_), .A2(new_n2964_), .Z(new_n3744_));
  NOR2_X1    g3692(.A1(new_n3738_), .A2(new_n3744_), .ZN(new_n3745_));
  XOR2_X1    g3693(.A1(new_n3651_), .A2(new_n3317_), .Z(new_n3746_));
  AOI21_X1   g3694(.A1(new_n3738_), .A2(new_n3744_), .B(new_n3746_), .ZN(new_n3747_));
  NOR2_X1    g3695(.A1(new_n3281_), .A2(new_n3739_), .ZN(new_n3748_));
  NOR2_X1    g3696(.A1(new_n2813_), .A2(new_n2939_), .ZN(new_n3749_));
  OAI21_X1   g3697(.A1(new_n3748_), .A2(new_n3749_), .B(new_n2942_), .ZN(new_n3750_));
  NAND2_X1   g3698(.A1(new_n3750_), .A2(new_n2940_), .ZN(new_n3751_));
  NOR2_X1    g3699(.A1(new_n3751_), .A2(new_n3279_), .ZN(new_n3752_));
  AOI21_X1   g3700(.A1(new_n2940_), .A2(new_n3750_), .B(new_n3128_), .ZN(new_n3753_));
  NOR2_X1    g3701(.A1(new_n3752_), .A2(new_n3753_), .ZN(new_n3754_));
  INV_X1     g3702(.I(new_n3754_), .ZN(new_n3755_));
  OAI21_X1   g3703(.A1(new_n3747_), .A2(new_n3745_), .B(new_n3755_), .ZN(new_n3756_));
  NOR3_X1    g3704(.A1(new_n3747_), .A2(new_n3745_), .A3(new_n3755_), .ZN(new_n3757_));
  XOR2_X1    g3705(.A1(new_n3654_), .A2(new_n3655_), .Z(new_n3758_));
  OAI21_X1   g3706(.A1(new_n3757_), .A2(new_n3758_), .B(new_n3756_), .ZN(new_n3759_));
  OAI22_X1   g3707(.A1(new_n2734_), .A2(new_n3639_), .B1(new_n2956_), .B2(new_n3636_), .ZN(new_n3760_));
  OAI21_X1   g3708(.A1(new_n2729_), .A2(new_n2939_), .B(new_n3760_), .ZN(new_n3761_));
  AOI21_X1   g3709(.A1(new_n3761_), .A2(new_n2942_), .B(new_n2939_), .ZN(new_n3762_));
  XOR2_X1    g3710(.A1(new_n3270_), .A2(new_n3762_), .Z(new_n3763_));
  INV_X1     g3711(.I(new_n3763_), .ZN(new_n3764_));
  NAND2_X1   g3712(.A1(new_n3759_), .A2(new_n3764_), .ZN(new_n3765_));
  XOR2_X1    g3713(.A1(new_n3346_), .A2(new_n3306_), .Z(new_n3766_));
  XOR2_X1    g3714(.A1(new_n3766_), .A2(new_n3338_), .Z(new_n3767_));
  OAI21_X1   g3715(.A1(new_n3759_), .A2(new_n3764_), .B(new_n3767_), .ZN(new_n3768_));
  INV_X1     g3716(.I(new_n3684_), .ZN(new_n3769_));
  NOR2_X1    g3717(.A1(new_n3235_), .A2(new_n3769_), .ZN(new_n3770_));
  NOR2_X1    g3718(.A1(new_n3770_), .A2(new_n3686_), .ZN(new_n3771_));
  OAI21_X1   g3719(.A1(new_n3698_), .A2(new_n3697_), .B(new_n3696_), .ZN(new_n3772_));
  NAND3_X1   g3720(.A1(new_n3692_), .A2(new_n3694_), .A3(new_n3350_), .ZN(new_n3773_));
  AOI21_X1   g3721(.A1(new_n3772_), .A2(new_n3773_), .B(new_n3771_), .ZN(new_n3774_));
  AOI21_X1   g3722(.A1(new_n3768_), .A2(new_n3765_), .B(new_n3774_), .ZN(new_n3775_));
  AOI22_X1   g3723(.A1(new_n2720_), .A2(new_n2947_), .B1(new_n2729_), .B2(new_n2949_), .ZN(new_n3776_));
  NOR2_X1    g3724(.A1(new_n2701_), .A2(new_n2939_), .ZN(new_n3777_));
  OAI21_X1   g3725(.A1(new_n3777_), .A2(new_n3776_), .B(new_n2942_), .ZN(new_n3778_));
  NAND2_X1   g3726(.A1(new_n3778_), .A2(new_n2940_), .ZN(new_n3779_));
  XNOR2_X1   g3727(.A1(new_n3202_), .A2(new_n3779_), .ZN(new_n3780_));
  INV_X1     g3728(.I(new_n3780_), .ZN(new_n3781_));
  OAI21_X1   g3729(.A1(new_n3775_), .A2(new_n3700_), .B(new_n3781_), .ZN(new_n3782_));
  NOR3_X1    g3730(.A1(new_n3775_), .A2(new_n3700_), .A3(new_n3781_), .ZN(new_n3783_));
  NOR2_X1    g3731(.A1(new_n3352_), .A2(new_n3349_), .ZN(new_n3784_));
  NOR2_X1    g3732(.A1(new_n3649_), .A2(new_n3667_), .ZN(new_n3785_));
  XNOR2_X1   g3733(.A1(new_n3785_), .A2(new_n3784_), .ZN(new_n3786_));
  OAI21_X1   g3734(.A1(new_n3783_), .A2(new_n3786_), .B(new_n3782_), .ZN(new_n3787_));
  OAI21_X1   g3735(.A1(new_n3680_), .A2(new_n3676_), .B(new_n3647_), .ZN(new_n3788_));
  AOI21_X1   g3736(.A1(new_n3787_), .A2(new_n3788_), .B(new_n3681_), .ZN(new_n3789_));
  XOR2_X1    g3737(.A1(new_n3265_), .A2(new_n3449_), .Z(new_n3790_));
  NOR2_X1    g3738(.A1(new_n3789_), .A2(new_n3790_), .ZN(new_n3791_));
  NOR2_X1    g3739(.A1(new_n3582_), .A2(new_n2939_), .ZN(new_n3792_));
  NOR2_X1    g3740(.A1(new_n3182_), .A2(new_n3636_), .ZN(new_n3793_));
  OAI22_X1   g3741(.A1(new_n2879_), .A2(new_n2939_), .B1(new_n3640_), .B2(new_n3793_), .ZN(new_n3794_));
  NOR2_X1    g3742(.A1(new_n3792_), .A2(new_n3794_), .ZN(new_n3795_));
  NOR2_X1    g3743(.A1(new_n3795_), .A2(new_n2942_), .ZN(new_n3796_));
  NOR3_X1    g3744(.A1(new_n3792_), .A2(new_n2943_), .A3(new_n3794_), .ZN(new_n3797_));
  NOR2_X1    g3745(.A1(new_n3796_), .A2(new_n3797_), .ZN(new_n3798_));
  AOI21_X1   g3746(.A1(new_n3789_), .A2(new_n3790_), .B(new_n3798_), .ZN(new_n3799_));
  NAND3_X1   g3747(.A1(new_n3223_), .A2(new_n3368_), .A3(new_n3264_), .ZN(new_n3800_));
  AND3_X2    g3748(.A1(new_n3800_), .A2(new_n3448_), .A3(new_n3363_), .Z(new_n3801_));
  AOI21_X1   g3749(.A1(new_n3800_), .A2(new_n3363_), .B(new_n3448_), .ZN(new_n3802_));
  OAI22_X1   g3750(.A1(new_n3799_), .A2(new_n3791_), .B1(new_n3801_), .B2(new_n3802_), .ZN(new_n3803_));
  OAI21_X1   g3751(.A1(new_n3679_), .A2(new_n3678_), .B(new_n3677_), .ZN(new_n3804_));
  NAND3_X1   g3752(.A1(new_n3671_), .A2(new_n3675_), .A3(new_n3360_), .ZN(new_n3805_));
  NAND3_X1   g3753(.A1(new_n3804_), .A2(new_n3805_), .A3(new_n3646_), .ZN(new_n3806_));
  INV_X1     g3754(.I(new_n3700_), .ZN(new_n3807_));
  NOR2_X1    g3755(.A1(new_n3710_), .A2(new_n3058_), .ZN(new_n3808_));
  NOR2_X1    g3756(.A1(new_n3066_), .A2(new_n3708_), .ZN(new_n3809_));
  INV_X1     g3757(.I(new_n3713_), .ZN(new_n3810_));
  OAI21_X1   g3758(.A1(new_n3808_), .A2(new_n3809_), .B(new_n3810_), .ZN(new_n3811_));
  NOR3_X1    g3759(.A1(new_n3808_), .A2(new_n3809_), .A3(new_n3810_), .ZN(new_n3812_));
  NAND2_X1   g3760(.A1(new_n3727_), .A2(new_n3732_), .ZN(new_n3813_));
  NAND2_X1   g3761(.A1(new_n3813_), .A2(new_n3735_), .ZN(new_n3814_));
  OAI21_X1   g3762(.A1(new_n3812_), .A2(new_n3814_), .B(new_n3811_), .ZN(new_n3815_));
  XOR2_X1    g3763(.A1(new_n3743_), .A2(new_n3511_), .Z(new_n3816_));
  NAND2_X1   g3764(.A1(new_n3815_), .A2(new_n3816_), .ZN(new_n3817_));
  INV_X1     g3765(.I(new_n3746_), .ZN(new_n3818_));
  OAI21_X1   g3766(.A1(new_n3815_), .A2(new_n3816_), .B(new_n3818_), .ZN(new_n3819_));
  AOI21_X1   g3767(.A1(new_n3819_), .A2(new_n3817_), .B(new_n3754_), .ZN(new_n3820_));
  NAND3_X1   g3768(.A1(new_n3819_), .A2(new_n3817_), .A3(new_n3754_), .ZN(new_n3821_));
  INV_X1     g3769(.I(new_n3758_), .ZN(new_n3822_));
  AOI21_X1   g3770(.A1(new_n3821_), .A2(new_n3822_), .B(new_n3820_), .ZN(new_n3823_));
  NOR2_X1    g3771(.A1(new_n3823_), .A2(new_n3763_), .ZN(new_n3824_));
  XOR2_X1    g3772(.A1(new_n3766_), .A2(new_n3657_), .Z(new_n3825_));
  AOI21_X1   g3773(.A1(new_n3823_), .A2(new_n3763_), .B(new_n3825_), .ZN(new_n3826_));
  OAI21_X1   g3774(.A1(new_n3699_), .A2(new_n3695_), .B(new_n3688_), .ZN(new_n3827_));
  OAI21_X1   g3775(.A1(new_n3826_), .A2(new_n3824_), .B(new_n3827_), .ZN(new_n3828_));
  AOI21_X1   g3776(.A1(new_n3828_), .A2(new_n3807_), .B(new_n3780_), .ZN(new_n3829_));
  NAND3_X1   g3777(.A1(new_n3828_), .A2(new_n3807_), .A3(new_n3780_), .ZN(new_n3830_));
  INV_X1     g3778(.I(new_n3786_), .ZN(new_n3831_));
  AOI21_X1   g3779(.A1(new_n3830_), .A2(new_n3831_), .B(new_n3829_), .ZN(new_n3832_));
  AOI21_X1   g3780(.A1(new_n3804_), .A2(new_n3805_), .B(new_n3646_), .ZN(new_n3833_));
  OAI21_X1   g3781(.A1(new_n3832_), .A2(new_n3833_), .B(new_n3806_), .ZN(new_n3834_));
  INV_X1     g3782(.I(new_n3790_), .ZN(new_n3835_));
  NAND2_X1   g3783(.A1(new_n3834_), .A2(new_n3835_), .ZN(new_n3836_));
  INV_X1     g3784(.I(new_n3798_), .ZN(new_n3837_));
  OAI21_X1   g3785(.A1(new_n3834_), .A2(new_n3835_), .B(new_n3837_), .ZN(new_n3838_));
  NOR2_X1    g3786(.A1(new_n3801_), .A2(new_n3802_), .ZN(new_n3839_));
  NAND3_X1   g3787(.A1(new_n3838_), .A2(new_n3836_), .A3(new_n3839_), .ZN(new_n3840_));
  XOR2_X1    g3788(.A1(new_n2898_), .A2(new_n2931_), .Z(new_n3841_));
  NAND2_X1   g3789(.A1(new_n3841_), .A2(new_n2882_), .ZN(new_n3842_));
  NAND2_X1   g3790(.A1(new_n2899_), .A2(new_n2932_), .ZN(new_n3843_));
  NAND2_X1   g3791(.A1(new_n3842_), .A2(new_n3843_), .ZN(new_n3844_));
  AOI22_X1   g3792(.A1(new_n2931_), .A2(new_n2949_), .B1(new_n3436_), .B2(new_n2940_), .ZN(new_n3845_));
  AOI21_X1   g3793(.A1(new_n2948_), .A2(new_n3845_), .B(new_n2939_), .ZN(new_n3846_));
  NAND2_X1   g3794(.A1(new_n3844_), .A2(new_n3846_), .ZN(new_n3847_));
  XOR2_X1    g3795(.A1(new_n3847_), .A2(new_n2943_), .Z(new_n3848_));
  INV_X1     g3796(.I(new_n3848_), .ZN(new_n3849_));
  NAND2_X1   g3797(.A1(new_n3840_), .A2(new_n3849_), .ZN(new_n3850_));
  NAND2_X1   g3798(.A1(new_n3850_), .A2(new_n3803_), .ZN(new_n3851_));
  NAND2_X1   g3799(.A1(new_n3634_), .A2(new_n3472_), .ZN(new_n3852_));
  NAND3_X1   g3800(.A1(new_n3635_), .A2(new_n3851_), .A3(new_n3852_), .ZN(new_n3853_));
  NOR2_X1    g3801(.A1(new_n3577_), .A2(new_n3586_), .ZN(new_n3854_));
  XOR2_X1    g3802(.A1(new_n3626_), .A2(new_n3854_), .Z(new_n3855_));
  XOR2_X1    g3803(.A1(new_n3612_), .A2(new_n2942_), .Z(new_n3856_));
  NOR2_X1    g3804(.A1(new_n3855_), .A2(new_n3856_), .ZN(new_n3857_));
  NOR2_X1    g3805(.A1(new_n2682_), .A2(new_n3237_), .ZN(new_n3858_));
  NAND2_X1   g3806(.A1(new_n2898_), .A2(new_n3210_), .ZN(new_n3859_));
  INV_X1     g3807(.I(new_n3859_), .ZN(new_n3860_));
  OAI22_X1   g3808(.A1(new_n3860_), .A2(new_n3858_), .B1(new_n2879_), .B2(new_n3213_), .ZN(new_n3861_));
  AOI21_X1   g3809(.A1(new_n3842_), .A2(new_n3843_), .B(new_n3207_), .ZN(new_n3862_));
  OAI21_X1   g3810(.A1(new_n3189_), .A2(new_n2972_), .B(new_n3480_), .ZN(new_n3863_));
  NAND3_X1   g3811(.A1(new_n2699_), .A2(new_n2700_), .A3(new_n2977_), .ZN(new_n3864_));
  AOI21_X1   g3812(.A1(new_n3863_), .A2(new_n3864_), .B(new_n803_), .ZN(new_n3865_));
  NOR4_X1    g3813(.A1(new_n3865_), .A2(new_n3197_), .A3(new_n3201_), .A4(new_n2969_), .ZN(new_n3866_));
  AOI22_X1   g3814(.A1(new_n2816_), .A2(new_n3198_), .B1(new_n2715_), .B2(new_n2719_), .ZN(new_n3867_));
  OAI21_X1   g3815(.A1(new_n3560_), .A2(new_n3867_), .B(new_n2701_), .ZN(new_n3868_));
  OAI21_X1   g3816(.A1(new_n3429_), .A2(new_n3428_), .B(new_n3182_), .ZN(new_n3869_));
  AOI22_X1   g3817(.A1(new_n2720_), .A2(new_n3086_), .B1(new_n2729_), .B2(new_n3076_), .ZN(new_n3870_));
  INV_X1     g3818(.I(new_n3864_), .ZN(new_n3871_));
  OAI21_X1   g3819(.A1(new_n3871_), .A2(new_n3870_), .B(new_n802_), .ZN(new_n3872_));
  AOI22_X1   g3820(.A1(new_n3868_), .A2(new_n3869_), .B1(new_n3872_), .B2(new_n2977_), .ZN(new_n3873_));
  NAND2_X1   g3821(.A1(new_n3527_), .A2(new_n3408_), .ZN(new_n3874_));
  NAND2_X1   g3822(.A1(new_n3874_), .A2(new_n3521_), .ZN(new_n3875_));
  NOR2_X1    g3823(.A1(new_n3506_), .A2(new_n3528_), .ZN(new_n3876_));
  NOR2_X1    g3824(.A1(new_n3541_), .A2(new_n3534_), .ZN(new_n3877_));
  NOR2_X1    g3825(.A1(new_n3877_), .A2(new_n3876_), .ZN(new_n3878_));
  INV_X1     g3826(.I(new_n3878_), .ZN(new_n3879_));
  OAI21_X1   g3827(.A1(new_n3874_), .A2(new_n3521_), .B(new_n3879_), .ZN(new_n3880_));
  AOI21_X1   g3828(.A1(new_n2743_), .A2(new_n2758_), .B(new_n3512_), .ZN(new_n3881_));
  NOR3_X1    g3829(.A1(new_n2733_), .A2(new_n2732_), .A3(new_n3028_), .ZN(new_n3882_));
  OAI21_X1   g3830(.A1(new_n3881_), .A2(new_n3882_), .B(new_n721_), .ZN(new_n3883_));
  NAND4_X1   g3831(.A1(new_n3278_), .A2(new_n3277_), .A3(new_n3883_), .A4(new_n2992_), .ZN(new_n3884_));
  OAI21_X1   g3832(.A1(new_n2956_), .A2(new_n2804_), .B(new_n3513_), .ZN(new_n3885_));
  NAND3_X1   g3833(.A1(new_n2812_), .A2(new_n2517_), .A3(new_n2998_), .ZN(new_n3886_));
  AOI21_X1   g3834(.A1(new_n3885_), .A2(new_n3886_), .B(new_n702_), .ZN(new_n3887_));
  OAI22_X1   g3835(.A1(new_n3127_), .A2(new_n3125_), .B1(new_n3887_), .B2(new_n2991_), .ZN(new_n3888_));
  NAND2_X1   g3836(.A1(new_n3888_), .A2(new_n3884_), .ZN(new_n3889_));
  OAI21_X1   g3837(.A1(new_n3505_), .A2(new_n3500_), .B(new_n3528_), .ZN(new_n3890_));
  OAI22_X1   g3838(.A1(new_n2770_), .A2(new_n3493_), .B1(new_n2792_), .B2(new_n3396_), .ZN(new_n3891_));
  OAI21_X1   g3839(.A1(new_n2764_), .A2(new_n2763_), .B(new_n3398_), .ZN(new_n3892_));
  AOI21_X1   g3840(.A1(new_n3891_), .A2(new_n3892_), .B(new_n438_), .ZN(new_n3893_));
  NOR4_X1    g3841(.A1(new_n3893_), .A2(new_n3073_), .A3(new_n3075_), .A4(new_n3501_), .ZN(new_n3894_));
  AOI21_X1   g3842(.A1(new_n2775_), .A2(new_n3494_), .B(new_n3397_), .ZN(new_n3895_));
  AOI21_X1   g3843(.A1(new_n2790_), .A2(new_n2789_), .B(new_n3496_), .ZN(new_n3896_));
  OAI21_X1   g3844(.A1(new_n3895_), .A2(new_n3896_), .B(new_n437_), .ZN(new_n3897_));
  AOI22_X1   g3845(.A1(new_n3143_), .A2(new_n3141_), .B1(new_n3897_), .B2(new_n3393_), .ZN(new_n3898_));
  NOR2_X1    g3846(.A1(new_n3898_), .A2(new_n3894_), .ZN(new_n3899_));
  NOR3_X1    g3847(.A1(new_n3890_), .A2(new_n3899_), .A3(new_n2786_), .ZN(new_n3900_));
  NAND3_X1   g3848(.A1(new_n3504_), .A2(new_n3024_), .A3(new_n3027_), .ZN(new_n3901_));
  OAI21_X1   g3849(.A1(new_n3036_), .A2(new_n3037_), .B(new_n3499_), .ZN(new_n3902_));
  AOI21_X1   g3850(.A1(new_n3902_), .A2(new_n3901_), .B(new_n3534_), .ZN(new_n3903_));
  NAND4_X1   g3851(.A1(new_n3143_), .A2(new_n3897_), .A3(new_n3141_), .A4(new_n3393_), .ZN(new_n3904_));
  OAI22_X1   g3852(.A1(new_n3893_), .A2(new_n3501_), .B1(new_n3073_), .B2(new_n3075_), .ZN(new_n3905_));
  NAND2_X1   g3853(.A1(new_n3905_), .A2(new_n3904_), .ZN(new_n3906_));
  AOI21_X1   g3854(.A1(new_n3903_), .A2(new_n3906_), .B(new_n2795_), .ZN(new_n3907_));
  OAI21_X1   g3855(.A1(new_n3900_), .A2(new_n3907_), .B(new_n437_), .ZN(new_n3908_));
  NAND3_X1   g3856(.A1(new_n3903_), .A2(new_n3906_), .A3(new_n2795_), .ZN(new_n3909_));
  OAI21_X1   g3857(.A1(new_n3890_), .A2(new_n3899_), .B(new_n2786_), .ZN(new_n3910_));
  NAND3_X1   g3858(.A1(new_n3910_), .A2(new_n3909_), .A3(new_n438_), .ZN(new_n3911_));
  NAND2_X1   g3859(.A1(new_n3908_), .A2(new_n3911_), .ZN(new_n3912_));
  NAND2_X1   g3860(.A1(new_n3889_), .A2(new_n3912_), .ZN(new_n3913_));
  NAND4_X1   g3861(.A1(new_n3884_), .A2(new_n3908_), .A3(new_n3888_), .A4(new_n3911_), .ZN(new_n3914_));
  AOI22_X1   g3862(.A1(new_n3880_), .A2(new_n3875_), .B1(new_n3913_), .B2(new_n3914_), .ZN(new_n3915_));
  NOR2_X1    g3863(.A1(new_n3532_), .A2(new_n3530_), .ZN(new_n3916_));
  NOR2_X1    g3864(.A1(new_n3916_), .A2(new_n3520_), .ZN(new_n3917_));
  AOI21_X1   g3865(.A1(new_n3916_), .A2(new_n3520_), .B(new_n3878_), .ZN(new_n3918_));
  AOI21_X1   g3866(.A1(new_n3910_), .A2(new_n3909_), .B(new_n438_), .ZN(new_n3919_));
  NOR3_X1    g3867(.A1(new_n3900_), .A2(new_n3907_), .A3(new_n437_), .ZN(new_n3920_));
  NOR2_X1    g3868(.A1(new_n3920_), .A2(new_n3919_), .ZN(new_n3921_));
  NOR2_X1    g3869(.A1(new_n3921_), .A2(new_n3889_), .ZN(new_n3922_));
  NOR4_X1    g3870(.A1(new_n3127_), .A2(new_n3125_), .A3(new_n3887_), .A4(new_n2991_), .ZN(new_n3923_));
  AOI22_X1   g3871(.A1(new_n3278_), .A2(new_n3277_), .B1(new_n3883_), .B2(new_n2992_), .ZN(new_n3924_));
  NOR2_X1    g3872(.A1(new_n3924_), .A2(new_n3923_), .ZN(new_n3925_));
  NOR2_X1    g3873(.A1(new_n3925_), .A2(new_n3912_), .ZN(new_n3926_));
  NOR2_X1    g3874(.A1(new_n3922_), .A2(new_n3926_), .ZN(new_n3927_));
  NOR3_X1    g3875(.A1(new_n3927_), .A2(new_n3918_), .A3(new_n3917_), .ZN(new_n3928_));
  NOR4_X1    g3876(.A1(new_n3915_), .A2(new_n3928_), .A3(new_n3866_), .A4(new_n3873_), .ZN(new_n3929_));
  NAND4_X1   g3877(.A1(new_n3868_), .A2(new_n3872_), .A3(new_n3869_), .A4(new_n2977_), .ZN(new_n3930_));
  OAI22_X1   g3878(.A1(new_n2969_), .A2(new_n3865_), .B1(new_n3197_), .B2(new_n3201_), .ZN(new_n3931_));
  NAND2_X1   g3879(.A1(new_n3913_), .A2(new_n3914_), .ZN(new_n3932_));
  OAI21_X1   g3880(.A1(new_n3918_), .A2(new_n3917_), .B(new_n3932_), .ZN(new_n3933_));
  NAND2_X1   g3881(.A1(new_n3925_), .A2(new_n3912_), .ZN(new_n3934_));
  NAND2_X1   g3882(.A1(new_n3921_), .A2(new_n3889_), .ZN(new_n3935_));
  NAND2_X1   g3883(.A1(new_n3935_), .A2(new_n3934_), .ZN(new_n3936_));
  NAND3_X1   g3884(.A1(new_n3936_), .A2(new_n3880_), .A3(new_n3875_), .ZN(new_n3937_));
  AOI22_X1   g3885(.A1(new_n3933_), .A2(new_n3937_), .B1(new_n3930_), .B2(new_n3931_), .ZN(new_n3938_));
  NOR3_X1    g3886(.A1(new_n3556_), .A2(new_n3929_), .A3(new_n3938_), .ZN(new_n3939_));
  NOR3_X1    g3887(.A1(new_n3939_), .A2(new_n3557_), .A3(new_n3475_), .ZN(new_n3940_));
  NAND4_X1   g3888(.A1(new_n3933_), .A2(new_n3937_), .A3(new_n3930_), .A4(new_n3931_), .ZN(new_n3941_));
  OAI22_X1   g3889(.A1(new_n3915_), .A2(new_n3928_), .B1(new_n3866_), .B2(new_n3873_), .ZN(new_n3942_));
  NAND3_X1   g3890(.A1(new_n3551_), .A2(new_n3942_), .A3(new_n3941_), .ZN(new_n3943_));
  AOI21_X1   g3891(.A1(new_n3943_), .A2(new_n3552_), .B(new_n3554_), .ZN(new_n3944_));
  OAI21_X1   g3892(.A1(new_n3940_), .A2(new_n3944_), .B(new_n1051_), .ZN(new_n3945_));
  NOR2_X1    g3893(.A1(new_n3945_), .A2(new_n3862_), .ZN(new_n3946_));
  NAND2_X1   g3894(.A1(new_n3844_), .A2(new_n3280_), .ZN(new_n3947_));
  NAND3_X1   g3895(.A1(new_n3943_), .A2(new_n3552_), .A3(new_n3554_), .ZN(new_n3948_));
  OAI21_X1   g3896(.A1(new_n3939_), .A2(new_n3557_), .B(new_n3475_), .ZN(new_n3949_));
  NAND2_X1   g3897(.A1(new_n3949_), .A2(new_n3948_), .ZN(new_n3950_));
  AOI21_X1   g3898(.A1(new_n3950_), .A2(new_n1051_), .B(new_n3947_), .ZN(new_n3951_));
  OAI21_X1   g3899(.A1(new_n3946_), .A2(new_n3951_), .B(new_n3861_), .ZN(new_n3952_));
  INV_X1     g3900(.I(new_n3861_), .ZN(new_n3953_));
  NAND3_X1   g3901(.A1(new_n3950_), .A2(new_n1051_), .A3(new_n3947_), .ZN(new_n3954_));
  NAND2_X1   g3902(.A1(new_n3945_), .A2(new_n3862_), .ZN(new_n3955_));
  NAND3_X1   g3903(.A1(new_n3955_), .A2(new_n3954_), .A3(new_n3953_), .ZN(new_n3956_));
  NAND3_X1   g3904(.A1(new_n3952_), .A2(new_n3956_), .A3(new_n3614_), .ZN(new_n3957_));
  NAND3_X1   g3905(.A1(new_n3957_), .A2(new_n3626_), .A3(new_n3854_), .ZN(new_n3958_));
  INV_X1     g3906(.I(new_n3958_), .ZN(new_n3959_));
  AOI21_X1   g3907(.A1(new_n3957_), .A2(new_n3626_), .B(new_n3854_), .ZN(new_n3960_));
  NOR2_X1    g3908(.A1(new_n3589_), .A2(new_n3588_), .ZN(new_n3961_));
  INV_X1     g3909(.I(new_n2924_), .ZN(new_n3962_));
  NOR4_X1    g3910(.A1(new_n2923_), .A2(new_n226_), .A3(new_n556_), .A4(new_n3592_), .ZN(new_n3963_));
  NAND2_X1   g3911(.A1(new_n3962_), .A2(new_n3963_), .ZN(new_n3964_));
  INV_X1     g3912(.I(new_n504_), .ZN(new_n3965_));
  INV_X1     g3913(.I(new_n234_), .ZN(new_n3966_));
  NOR2_X1    g3914(.A1(new_n200_), .A2(new_n212_), .ZN(new_n3967_));
  INV_X1     g3915(.I(new_n3967_), .ZN(new_n3968_));
  NOR3_X1    g3916(.A1(new_n3966_), .A2(new_n2859_), .A3(new_n3968_), .ZN(new_n3969_));
  NOR3_X1    g3917(.A1(new_n922_), .A2(new_n246_), .A3(new_n187_), .ZN(new_n3970_));
  NAND2_X1   g3918(.A1(new_n3969_), .A2(new_n3970_), .ZN(new_n3971_));
  NOR3_X1    g3919(.A1(new_n3971_), .A2(new_n259_), .A3(new_n3965_), .ZN(new_n3972_));
  NAND4_X1   g3920(.A1(new_n3972_), .A2(new_n176_), .A3(new_n531_), .A4(new_n542_), .ZN(new_n3973_));
  NAND2_X1   g3921(.A1(new_n3964_), .A2(new_n3973_), .ZN(new_n3974_));
  INV_X1     g3922(.I(new_n3973_), .ZN(new_n3975_));
  NAND3_X1   g3923(.A1(new_n3962_), .A2(new_n3963_), .A3(new_n3975_), .ZN(new_n3976_));
  NAND2_X1   g3924(.A1(new_n3974_), .A2(new_n3976_), .ZN(new_n3977_));
  XOR2_X1    g3925(.A1(new_n3977_), .A2(new_n2946_), .Z(new_n3978_));
  NAND3_X1   g3926(.A1(new_n3978_), .A2(new_n3961_), .A3(new_n3605_), .ZN(new_n3979_));
  NAND2_X1   g3927(.A1(new_n3978_), .A2(new_n3605_), .ZN(new_n3980_));
  NAND2_X1   g3928(.A1(new_n3980_), .A2(new_n3618_), .ZN(new_n3981_));
  NAND2_X1   g3929(.A1(new_n3981_), .A2(new_n3979_), .ZN(new_n3982_));
  INV_X1     g3930(.I(new_n3595_), .ZN(new_n3983_));
  NAND2_X1   g3931(.A1(new_n2906_), .A2(new_n3594_), .ZN(new_n3984_));
  NAND2_X1   g3932(.A1(new_n3984_), .A2(new_n3983_), .ZN(new_n3985_));
  AOI22_X1   g3933(.A1(new_n2946_), .A2(new_n2949_), .B1(new_n3985_), .B2(new_n2947_), .ZN(new_n3986_));
  INV_X1     g3934(.I(new_n3977_), .ZN(new_n3987_));
  NOR2_X1    g3935(.A1(new_n3987_), .A2(new_n2939_), .ZN(new_n3988_));
  OAI21_X1   g3936(.A1(new_n3988_), .A2(new_n3986_), .B(new_n2942_), .ZN(new_n3989_));
  NAND2_X1   g3937(.A1(new_n3989_), .A2(new_n2940_), .ZN(new_n3990_));
  XNOR2_X1   g3938(.A1(new_n3982_), .A2(new_n3990_), .ZN(new_n3991_));
  OAI21_X1   g3939(.A1(new_n3959_), .A2(new_n3960_), .B(new_n3991_), .ZN(new_n3992_));
  NOR2_X1    g3940(.A1(new_n3992_), .A2(new_n3857_), .ZN(new_n3993_));
  INV_X1     g3941(.I(new_n3857_), .ZN(new_n3994_));
  INV_X1     g3942(.I(new_n3960_), .ZN(new_n3995_));
  NAND2_X1   g3943(.A1(new_n3995_), .A2(new_n3958_), .ZN(new_n3996_));
  AOI21_X1   g3944(.A1(new_n3996_), .A2(new_n3991_), .B(new_n3994_), .ZN(new_n3997_));
  OAI21_X1   g3945(.A1(new_n3993_), .A2(new_n3997_), .B(new_n3853_), .ZN(new_n3998_));
  INV_X1     g3946(.I(new_n2953_), .ZN(new_n3999_));
  OAI21_X1   g3947(.A1(new_n3632_), .A2(new_n3631_), .B(new_n2942_), .ZN(new_n4000_));
  NAND3_X1   g3948(.A1(new_n3624_), .A2(new_n3629_), .A3(new_n2943_), .ZN(new_n4001_));
  NAND2_X1   g3949(.A1(new_n4001_), .A2(new_n4000_), .ZN(new_n4002_));
  AOI21_X1   g3950(.A1(new_n4002_), .A2(new_n3471_), .B(new_n3999_), .ZN(new_n4003_));
  NOR2_X1    g3951(.A1(new_n3799_), .A2(new_n3791_), .ZN(new_n4004_));
  NOR2_X1    g3952(.A1(new_n4004_), .A2(new_n3839_), .ZN(new_n4005_));
  AOI21_X1   g3953(.A1(new_n4004_), .A2(new_n3839_), .B(new_n3848_), .ZN(new_n4006_));
  NOR2_X1    g3954(.A1(new_n4006_), .A2(new_n4005_), .ZN(new_n4007_));
  NOR2_X1    g3955(.A1(new_n4002_), .A2(new_n3471_), .ZN(new_n4008_));
  NOR3_X1    g3956(.A1(new_n4007_), .A2(new_n4003_), .A3(new_n4008_), .ZN(new_n4009_));
  NAND3_X1   g3957(.A1(new_n3996_), .A2(new_n3994_), .A3(new_n3991_), .ZN(new_n4010_));
  NAND2_X1   g3958(.A1(new_n3992_), .A2(new_n3857_), .ZN(new_n4011_));
  NAND3_X1   g3959(.A1(new_n4009_), .A2(new_n4010_), .A3(new_n4011_), .ZN(new_n4012_));
  NAND2_X1   g3960(.A1(new_n3998_), .A2(new_n4012_), .ZN(new_n4013_));
  NOR2_X1    g3961(.A1(new_n3471_), .A2(new_n2953_), .ZN(new_n4014_));
  AOI22_X1   g3962(.A1(new_n3850_), .A2(new_n3803_), .B1(new_n2953_), .B2(new_n3471_), .ZN(new_n4015_));
  NOR3_X1    g3963(.A1(new_n4015_), .A2(new_n3855_), .A3(new_n4014_), .ZN(new_n4016_));
  INV_X1     g3964(.I(new_n3855_), .ZN(new_n4017_));
  INV_X1     g3965(.I(new_n4014_), .ZN(new_n4018_));
  NAND2_X1   g3966(.A1(new_n3471_), .A2(new_n2953_), .ZN(new_n4019_));
  OAI21_X1   g3967(.A1(new_n4006_), .A2(new_n4005_), .B(new_n4019_), .ZN(new_n4020_));
  AOI21_X1   g3968(.A1(new_n4020_), .A2(new_n4018_), .B(new_n4017_), .ZN(new_n4021_));
  OAI21_X1   g3969(.A1(new_n4016_), .A2(new_n4021_), .B(new_n3856_), .ZN(new_n4022_));
  INV_X1     g3970(.I(new_n3856_), .ZN(new_n4023_));
  NAND3_X1   g3971(.A1(new_n4020_), .A2(new_n4017_), .A3(new_n4018_), .ZN(new_n4024_));
  OAI21_X1   g3972(.A1(new_n4015_), .A2(new_n4014_), .B(new_n3855_), .ZN(new_n4025_));
  NAND3_X1   g3973(.A1(new_n4025_), .A2(new_n4024_), .A3(new_n4023_), .ZN(new_n4026_));
  NOR4_X1    g3974(.A1(new_n2440_), .A2(new_n413_), .A3(new_n1069_), .A4(new_n332_), .ZN(new_n4027_));
  NAND3_X1   g3975(.A1(new_n223_), .A2(new_n374_), .A3(new_n517_), .ZN(new_n4028_));
  NOR2_X1    g3976(.A1(new_n4028_), .A2(new_n660_), .ZN(new_n4029_));
  NAND4_X1   g3977(.A1(new_n2348_), .A2(new_n4027_), .A3(new_n4029_), .A4(new_n2451_), .ZN(new_n4030_));
  NOR3_X1    g3978(.A1(new_n2394_), .A2(new_n214_), .A3(new_n367_), .ZN(new_n4031_));
  NAND4_X1   g3979(.A1(new_n2282_), .A2(new_n4031_), .A3(new_n234_), .A4(new_n2243_), .ZN(new_n4032_));
  NOR2_X1    g3980(.A1(new_n321_), .A2(new_n312_), .ZN(new_n4033_));
  NAND4_X1   g3981(.A1(new_n4033_), .A2(new_n463_), .A3(new_n364_), .A4(new_n2858_), .ZN(new_n4034_));
  NOR3_X1    g3982(.A1(new_n4034_), .A2(new_n4030_), .A3(new_n4032_), .ZN(new_n4035_));
  INV_X1     g3983(.I(new_n4035_), .ZN(new_n4036_));
  AOI21_X1   g3984(.A1(new_n4022_), .A2(new_n4026_), .B(new_n4036_), .ZN(new_n4037_));
  NAND2_X1   g3985(.A1(new_n4037_), .A2(new_n4013_), .ZN(new_n4038_));
  NAND4_X1   g3986(.A1(new_n305_), .A2(new_n539_), .A3(new_n602_), .A4(new_n510_), .ZN(new_n4039_));
  NOR4_X1    g3987(.A1(new_n4039_), .A2(new_n217_), .A3(new_n609_), .A4(new_n834_), .ZN(new_n4040_));
  NAND3_X1   g3988(.A1(new_n4040_), .A2(new_n905_), .A3(new_n2335_), .ZN(new_n4041_));
  NOR4_X1    g3989(.A1(new_n4041_), .A2(new_n151_), .A3(new_n398_), .A4(new_n355_), .ZN(new_n4042_));
  NOR4_X1    g3990(.A1(new_n1088_), .A2(new_n619_), .A3(new_n375_), .A4(new_n292_), .ZN(new_n4043_));
  INV_X1     g3991(.I(new_n4043_), .ZN(new_n4044_));
  NAND4_X1   g3992(.A1(new_n228_), .A2(new_n220_), .A3(new_n326_), .A4(new_n375_), .ZN(new_n4045_));
  NAND2_X1   g3993(.A1(new_n2346_), .A2(new_n347_), .ZN(new_n4046_));
  NOR4_X1    g3994(.A1(new_n4044_), .A2(new_n358_), .A3(new_n4045_), .A4(new_n4046_), .ZN(new_n4047_));
  NAND3_X1   g3995(.A1(new_n2240_), .A2(new_n310_), .A3(new_n608_), .ZN(new_n4048_));
  NAND3_X1   g3996(.A1(new_n781_), .A2(new_n160_), .A3(new_n232_), .ZN(new_n4049_));
  NOR4_X1    g3997(.A1(new_n4049_), .A2(new_n4048_), .A3(new_n505_), .A4(new_n791_), .ZN(new_n4050_));
  NAND4_X1   g3998(.A1(new_n4042_), .A2(new_n2406_), .A3(new_n4047_), .A4(new_n4050_), .ZN(new_n4051_));
  INV_X1     g3999(.I(new_n4051_), .ZN(new_n4052_));
  OAI21_X1   g4000(.A1(new_n4037_), .A2(new_n4013_), .B(new_n4052_), .ZN(new_n4053_));
  NAND2_X1   g4001(.A1(new_n254_), .A2(new_n341_), .ZN(new_n4054_));
  NOR4_X1    g4002(.A1(new_n2918_), .A2(new_n4054_), .A3(new_n222_), .A4(new_n363_), .ZN(new_n4055_));
  NOR2_X1    g4003(.A1(new_n160_), .A2(new_n245_), .ZN(new_n4056_));
  NAND4_X1   g4004(.A1(new_n2231_), .A2(new_n4056_), .A3(new_n602_), .A4(new_n510_), .ZN(new_n4057_));
  NOR2_X1    g4005(.A1(new_n820_), .A2(new_n388_), .ZN(new_n4058_));
  NOR4_X1    g4006(.A1(new_n132_), .A2(new_n367_), .A3(new_n485_), .A4(new_n416_), .ZN(new_n4059_));
  NAND2_X1   g4007(.A1(new_n4059_), .A2(new_n4058_), .ZN(new_n4060_));
  NOR2_X1    g4008(.A1(new_n4057_), .A2(new_n4060_), .ZN(new_n4061_));
  NOR4_X1    g4009(.A1(new_n205_), .A2(new_n468_), .A3(new_n395_), .A4(new_n311_), .ZN(new_n4062_));
  AND3_X2    g4010(.A1(new_n4061_), .A2(new_n4055_), .A3(new_n4062_), .Z(new_n4063_));
  INV_X1     g4011(.I(new_n4063_), .ZN(new_n4064_));
  OR4_X2     g4012(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .A4(new_n444_), .Z(new_n4065_));
  NOR4_X1    g4013(.A1(new_n227_), .A2(new_n401_), .A3(new_n156_), .A4(new_n353_), .ZN(new_n4066_));
  INV_X1     g4014(.I(new_n4066_), .ZN(new_n4067_));
  NOR3_X1    g4015(.A1(new_n4065_), .A2(new_n2913_), .A3(new_n4067_), .ZN(new_n4068_));
  INV_X1     g4016(.I(new_n4068_), .ZN(new_n4069_));
  NOR4_X1    g4017(.A1(new_n207_), .A2(new_n417_), .A3(new_n141_), .A4(new_n251_), .ZN(new_n4070_));
  NOR4_X1    g4018(.A1(new_n2417_), .A2(new_n465_), .A3(new_n2318_), .A4(new_n367_), .ZN(new_n4071_));
  NAND4_X1   g4019(.A1(new_n4071_), .A2(new_n2853_), .A3(new_n2920_), .A4(new_n4070_), .ZN(new_n4072_));
  NOR4_X1    g4020(.A1(new_n4064_), .A2(new_n2435_), .A3(new_n4069_), .A4(new_n4072_), .ZN(new_n4073_));
  INV_X1     g4021(.I(new_n4073_), .ZN(new_n4074_));
  AOI21_X1   g4022(.A1(new_n4053_), .A2(new_n4038_), .B(new_n4074_), .ZN(new_n4075_));
  NAND3_X1   g4023(.A1(new_n4053_), .A2(new_n4038_), .A3(new_n4074_), .ZN(new_n4076_));
  OAI21_X1   g4024(.A1(new_n3996_), .A2(new_n3991_), .B(new_n3857_), .ZN(new_n4077_));
  OAI21_X1   g4025(.A1(new_n3853_), .A2(new_n4077_), .B(new_n3992_), .ZN(new_n4078_));
  NOR2_X1    g4026(.A1(new_n3945_), .A2(new_n3953_), .ZN(new_n4079_));
  AOI21_X1   g4027(.A1(new_n3950_), .A2(new_n1051_), .B(new_n3861_), .ZN(new_n4080_));
  OAI21_X1   g4028(.A1(new_n4079_), .A2(new_n4080_), .B(new_n3862_), .ZN(new_n4081_));
  INV_X1     g4029(.I(new_n4081_), .ZN(new_n4082_));
  INV_X1     g4030(.I(new_n3854_), .ZN(new_n4083_));
  AOI21_X1   g4031(.A1(new_n3952_), .A2(new_n3956_), .B(new_n3614_), .ZN(new_n4084_));
  OAI21_X1   g4032(.A1(new_n4084_), .A2(new_n3626_), .B(new_n4083_), .ZN(new_n4085_));
  NOR2_X1    g4033(.A1(new_n2931_), .A2(new_n3213_), .ZN(new_n4086_));
  OAI22_X1   g4034(.A1(new_n3860_), .A2(new_n4086_), .B1(new_n2926_), .B2(new_n3237_), .ZN(new_n4087_));
  AOI21_X1   g4035(.A1(new_n4087_), .A2(new_n1050_), .B(new_n3207_), .ZN(new_n4088_));
  NAND3_X1   g4036(.A1(new_n2934_), .A2(new_n4088_), .A3(new_n2928_), .ZN(new_n4089_));
  AOI21_X1   g4037(.A1(new_n2934_), .A2(new_n2928_), .B(new_n4088_), .ZN(new_n4090_));
  INV_X1     g4038(.I(new_n4090_), .ZN(new_n4091_));
  NAND2_X1   g4039(.A1(new_n4091_), .A2(new_n4089_), .ZN(new_n4092_));
  NOR2_X1    g4040(.A1(new_n3183_), .A2(new_n2969_), .ZN(new_n4093_));
  INV_X1     g4041(.I(new_n4093_), .ZN(new_n4094_));
  NAND2_X1   g4042(.A1(new_n3436_), .A2(new_n3086_), .ZN(new_n4095_));
  AOI22_X1   g4043(.A1(new_n4095_), .A2(new_n4094_), .B1(new_n3182_), .B2(new_n3076_), .ZN(new_n4096_));
  OAI21_X1   g4044(.A1(new_n4096_), .A2(new_n803_), .B(new_n2977_), .ZN(new_n4097_));
  NOR3_X1    g4045(.A1(new_n3432_), .A2(new_n3440_), .A3(new_n4097_), .ZN(new_n4098_));
  NOR2_X1    g4046(.A1(new_n2682_), .A2(new_n2975_), .ZN(new_n4099_));
  OAI22_X1   g4047(.A1(new_n4099_), .A2(new_n4093_), .B1(new_n2701_), .B2(new_n2972_), .ZN(new_n4100_));
  AOI21_X1   g4048(.A1(new_n4100_), .A2(new_n802_), .B(new_n2969_), .ZN(new_n4101_));
  AOI21_X1   g4049(.A1(new_n3463_), .A2(new_n3462_), .B(new_n4101_), .ZN(new_n4102_));
  NOR2_X1    g4050(.A1(new_n4098_), .A2(new_n4102_), .ZN(new_n4103_));
  OAI21_X1   g4051(.A1(new_n3918_), .A2(new_n3917_), .B(new_n3935_), .ZN(new_n4104_));
  NAND2_X1   g4052(.A1(new_n4104_), .A2(new_n3934_), .ZN(new_n4105_));
  AOI22_X1   g4053(.A1(new_n2813_), .A2(new_n3030_), .B1(new_n2743_), .B2(new_n3038_), .ZN(new_n4106_));
  NOR2_X1    g4054(.A1(new_n2729_), .A2(new_n3028_), .ZN(new_n4107_));
  OAI21_X1   g4055(.A1(new_n4107_), .A2(new_n4106_), .B(new_n721_), .ZN(new_n4108_));
  NAND4_X1   g4056(.A1(new_n3372_), .A2(new_n4108_), .A3(new_n2992_), .A4(new_n3268_), .ZN(new_n4109_));
  INV_X1     g4057(.I(new_n4106_), .ZN(new_n4110_));
  NAND2_X1   g4058(.A1(new_n3189_), .A2(new_n2998_), .ZN(new_n4111_));
  AOI21_X1   g4059(.A1(new_n4111_), .A2(new_n4110_), .B(new_n702_), .ZN(new_n4112_));
  OAI22_X1   g4060(.A1(new_n3266_), .A2(new_n3269_), .B1(new_n4112_), .B2(new_n2991_), .ZN(new_n4113_));
  NAND2_X1   g4061(.A1(new_n4113_), .A2(new_n4109_), .ZN(new_n4114_));
  NAND2_X1   g4062(.A1(new_n3903_), .A2(new_n3906_), .ZN(new_n4115_));
  NOR2_X1    g4063(.A1(new_n2795_), .A2(new_n437_), .ZN(new_n4116_));
  OAI21_X1   g4064(.A1(new_n3903_), .A2(new_n3906_), .B(new_n4116_), .ZN(new_n4117_));
  NAND2_X1   g4065(.A1(new_n4117_), .A2(new_n4115_), .ZN(new_n4118_));
  NAND3_X1   g4066(.A1(new_n3057_), .A2(new_n3053_), .A3(new_n3393_), .ZN(new_n4119_));
  OAI22_X1   g4067(.A1(new_n2765_), .A2(new_n3493_), .B1(new_n2770_), .B2(new_n3396_), .ZN(new_n4120_));
  NAND2_X1   g4068(.A1(new_n2758_), .A2(new_n3398_), .ZN(new_n4121_));
  NAND2_X1   g4069(.A1(new_n4121_), .A2(new_n4120_), .ZN(new_n4122_));
  INV_X1     g4070(.I(new_n4122_), .ZN(new_n4123_));
  NAND3_X1   g4071(.A1(new_n4118_), .A2(new_n4119_), .A3(new_n4123_), .ZN(new_n4124_));
  NOR2_X1    g4072(.A1(new_n4124_), .A2(new_n438_), .ZN(new_n4125_));
  NAND2_X1   g4073(.A1(new_n4124_), .A2(new_n438_), .ZN(new_n4126_));
  INV_X1     g4074(.I(new_n4126_), .ZN(new_n4127_));
  OAI21_X1   g4075(.A1(new_n4127_), .A2(new_n4125_), .B(new_n2792_), .ZN(new_n4128_));
  NOR2_X1    g4076(.A1(new_n3890_), .A2(new_n3899_), .ZN(new_n4129_));
  INV_X1     g4077(.I(new_n4116_), .ZN(new_n4130_));
  AOI21_X1   g4078(.A1(new_n3890_), .A2(new_n3899_), .B(new_n4130_), .ZN(new_n4131_));
  NOR2_X1    g4079(.A1(new_n4131_), .A2(new_n4129_), .ZN(new_n4132_));
  NOR3_X1    g4080(.A1(new_n3064_), .A2(new_n3065_), .A3(new_n3501_), .ZN(new_n4133_));
  NOR3_X1    g4081(.A1(new_n4132_), .A2(new_n4133_), .A3(new_n4122_), .ZN(new_n4134_));
  NAND2_X1   g4082(.A1(new_n4134_), .A2(new_n437_), .ZN(new_n4135_));
  NAND3_X1   g4083(.A1(new_n4135_), .A2(new_n4126_), .A3(new_n2783_), .ZN(new_n4136_));
  AOI21_X1   g4084(.A1(new_n4128_), .A2(new_n4136_), .B(new_n4114_), .ZN(new_n4137_));
  INV_X1     g4085(.I(new_n4114_), .ZN(new_n4138_));
  AOI21_X1   g4086(.A1(new_n4135_), .A2(new_n4126_), .B(new_n2783_), .ZN(new_n4139_));
  NOR3_X1    g4087(.A1(new_n4127_), .A2(new_n4125_), .A3(new_n2792_), .ZN(new_n4140_));
  NOR3_X1    g4088(.A1(new_n4138_), .A2(new_n4140_), .A3(new_n4139_), .ZN(new_n4141_));
  OAI21_X1   g4089(.A1(new_n4137_), .A2(new_n4141_), .B(new_n4105_), .ZN(new_n4142_));
  OAI21_X1   g4090(.A1(new_n4140_), .A2(new_n4139_), .B(new_n4114_), .ZN(new_n4143_));
  NAND3_X1   g4091(.A1(new_n4138_), .A2(new_n4128_), .A3(new_n4136_), .ZN(new_n4144_));
  NAND2_X1   g4092(.A1(new_n4144_), .A2(new_n4143_), .ZN(new_n4145_));
  NAND3_X1   g4093(.A1(new_n4145_), .A2(new_n3934_), .A3(new_n4104_), .ZN(new_n4146_));
  NAND3_X1   g4094(.A1(new_n4103_), .A2(new_n4146_), .A3(new_n4142_), .ZN(new_n4147_));
  NAND3_X1   g4095(.A1(new_n3463_), .A2(new_n4101_), .A3(new_n3462_), .ZN(new_n4148_));
  OAI21_X1   g4096(.A1(new_n3432_), .A2(new_n3440_), .B(new_n4097_), .ZN(new_n4149_));
  NAND2_X1   g4097(.A1(new_n4149_), .A2(new_n4148_), .ZN(new_n4150_));
  OAI21_X1   g4098(.A1(new_n4139_), .A2(new_n4140_), .B(new_n4138_), .ZN(new_n4151_));
  NAND3_X1   g4099(.A1(new_n4128_), .A2(new_n4136_), .A3(new_n4114_), .ZN(new_n4152_));
  AOI22_X1   g4100(.A1(new_n4151_), .A2(new_n4152_), .B1(new_n3934_), .B2(new_n4104_), .ZN(new_n4153_));
  AOI21_X1   g4101(.A1(new_n4143_), .A2(new_n4144_), .B(new_n4105_), .ZN(new_n4154_));
  OAI21_X1   g4102(.A1(new_n4153_), .A2(new_n4154_), .B(new_n4150_), .ZN(new_n4155_));
  NAND2_X1   g4103(.A1(new_n4155_), .A2(new_n4147_), .ZN(new_n4156_));
  OAI21_X1   g4104(.A1(new_n3555_), .A2(new_n3556_), .B(new_n3475_), .ZN(new_n4158_));
  AOI21_X1   g4105(.A1(new_n3942_), .A2(new_n4158_), .B(new_n4156_), .ZN(new_n4159_));
  NAND3_X1   g4106(.A1(new_n4156_), .A2(new_n3942_), .A3(new_n4158_), .ZN(new_n4160_));
  INV_X1     g4107(.I(new_n4160_), .ZN(new_n4161_));
  OAI21_X1   g4108(.A1(new_n4161_), .A2(new_n4159_), .B(new_n4092_), .ZN(new_n4162_));
  INV_X1     g4109(.I(new_n4162_), .ZN(new_n4163_));
  NAND2_X1   g4110(.A1(new_n4085_), .A2(new_n4163_), .ZN(new_n4164_));
  AOI21_X1   g4111(.A1(new_n3955_), .A2(new_n3954_), .B(new_n3953_), .ZN(new_n4165_));
  NOR3_X1    g4112(.A1(new_n3946_), .A2(new_n3951_), .A3(new_n3861_), .ZN(new_n4166_));
  OAI21_X1   g4113(.A1(new_n4166_), .A2(new_n4165_), .B(new_n3577_), .ZN(new_n4167_));
  NAND2_X1   g4114(.A1(new_n4167_), .A2(new_n3474_), .ZN(new_n4168_));
  NAND3_X1   g4115(.A1(new_n4168_), .A2(new_n4083_), .A3(new_n4162_), .ZN(new_n4169_));
  AOI21_X1   g4116(.A1(new_n4169_), .A2(new_n4164_), .B(new_n4082_), .ZN(new_n4170_));
  AOI21_X1   g4117(.A1(new_n4168_), .A2(new_n4083_), .B(new_n4162_), .ZN(new_n4171_));
  NOR2_X1    g4118(.A1(new_n4085_), .A2(new_n4163_), .ZN(new_n4172_));
  NOR3_X1    g4119(.A1(new_n4171_), .A2(new_n4172_), .A3(new_n4081_), .ZN(new_n4173_));
  NAND3_X1   g4120(.A1(new_n248_), .A2(new_n363_), .A3(new_n1248_), .ZN(new_n4174_));
  NAND2_X1   g4121(.A1(new_n208_), .A2(new_n521_), .ZN(new_n4175_));
  INV_X1     g4122(.I(new_n531_), .ZN(new_n4176_));
  NOR3_X1    g4123(.A1(new_n4176_), .A2(new_n233_), .A3(new_n407_), .ZN(new_n4177_));
  INV_X1     g4124(.I(new_n4177_), .ZN(new_n4178_));
  NOR4_X1    g4125(.A1(new_n4178_), .A2(new_n556_), .A3(new_n4174_), .A4(new_n4175_), .ZN(new_n4179_));
  AND2_X2    g4126(.A1(new_n3976_), .A2(new_n4179_), .Z(new_n4180_));
  NOR2_X1    g4127(.A1(new_n3976_), .A2(new_n4179_), .ZN(new_n4181_));
  NOR2_X1    g4128(.A1(new_n4180_), .A2(new_n4181_), .ZN(new_n4182_));
  OAI21_X1   g4129(.A1(new_n3618_), .A2(new_n3599_), .B(new_n3977_), .ZN(new_n4183_));
  NAND2_X1   g4130(.A1(new_n3618_), .A2(new_n3598_), .ZN(new_n4184_));
  NAND2_X1   g4131(.A1(new_n4183_), .A2(new_n4184_), .ZN(new_n4185_));
  NAND2_X1   g4132(.A1(new_n4185_), .A2(new_n3977_), .ZN(new_n4186_));
  AOI21_X1   g4133(.A1(new_n3961_), .A2(new_n3600_), .B(new_n3987_), .ZN(new_n4187_));
  NOR2_X1    g4134(.A1(new_n3961_), .A2(new_n3616_), .ZN(new_n4188_));
  NOR2_X1    g4135(.A1(new_n4187_), .A2(new_n4188_), .ZN(new_n4189_));
  NAND2_X1   g4136(.A1(new_n4189_), .A2(new_n3987_), .ZN(new_n4190_));
  AOI21_X1   g4137(.A1(new_n4190_), .A2(new_n4186_), .B(new_n4182_), .ZN(new_n4191_));
  INV_X1     g4138(.I(new_n4182_), .ZN(new_n4192_));
  NOR4_X1    g4139(.A1(new_n3618_), .A2(new_n3987_), .A3(new_n2946_), .A4(new_n3985_), .ZN(new_n4193_));
  NAND4_X1   g4140(.A1(new_n3618_), .A2(new_n3987_), .A3(new_n2946_), .A4(new_n3985_), .ZN(new_n4194_));
  INV_X1     g4141(.I(new_n4194_), .ZN(new_n4195_));
  NOR2_X1    g4142(.A1(new_n4195_), .A2(new_n4193_), .ZN(new_n4196_));
  NOR2_X1    g4143(.A1(new_n4196_), .A2(new_n4192_), .ZN(new_n4197_));
  NOR2_X1    g4144(.A1(new_n4191_), .A2(new_n4197_), .ZN(new_n4198_));
  OAI22_X1   g4145(.A1(new_n3987_), .A2(new_n3639_), .B1(new_n3636_), .B2(new_n3597_), .ZN(new_n4199_));
  OAI21_X1   g4146(.A1(new_n2939_), .A2(new_n4192_), .B(new_n4199_), .ZN(new_n4200_));
  AOI21_X1   g4147(.A1(new_n4200_), .A2(new_n2942_), .B(new_n2939_), .ZN(new_n4201_));
  XOR2_X1    g4148(.A1(new_n4198_), .A2(new_n4201_), .Z(new_n4202_));
  NOR3_X1    g4149(.A1(new_n4170_), .A2(new_n4173_), .A3(new_n4202_), .ZN(new_n4203_));
  OAI21_X1   g4150(.A1(new_n4171_), .A2(new_n4172_), .B(new_n4081_), .ZN(new_n4204_));
  NAND3_X1   g4151(.A1(new_n4169_), .A2(new_n4164_), .A3(new_n4082_), .ZN(new_n4205_));
  INV_X1     g4152(.I(new_n4202_), .ZN(new_n4206_));
  AOI21_X1   g4153(.A1(new_n4204_), .A2(new_n4205_), .B(new_n4206_), .ZN(new_n4207_));
  NOR2_X1    g4154(.A1(new_n4203_), .A2(new_n4207_), .ZN(new_n4208_));
  XOR2_X1    g4155(.A1(new_n4208_), .A2(new_n4078_), .Z(new_n4209_));
  INV_X1     g4156(.I(new_n4209_), .ZN(new_n4210_));
  AOI21_X1   g4157(.A1(new_n4076_), .A2(new_n4210_), .B(new_n4075_), .ZN(new_n4211_));
  NAND3_X1   g4158(.A1(new_n4204_), .A2(new_n4205_), .A3(new_n4206_), .ZN(new_n4212_));
  OAI21_X1   g4159(.A1(new_n4170_), .A2(new_n4173_), .B(new_n4202_), .ZN(new_n4213_));
  NAND2_X1   g4160(.A1(new_n4213_), .A2(new_n4212_), .ZN(new_n4214_));
  NAND2_X1   g4161(.A1(new_n4204_), .A2(new_n4205_), .ZN(new_n4215_));
  NAND2_X1   g4162(.A1(new_n4215_), .A2(new_n4206_), .ZN(new_n4216_));
  NOR3_X1    g4163(.A1(new_n4161_), .A2(new_n4092_), .A3(new_n4159_), .ZN(new_n4217_));
  NOR2_X1    g4164(.A1(new_n4217_), .A2(new_n4081_), .ZN(new_n4218_));
  INV_X1     g4165(.I(new_n4218_), .ZN(new_n4219_));
  OAI21_X1   g4166(.A1(new_n4085_), .A2(new_n4219_), .B(new_n4162_), .ZN(new_n4220_));
  INV_X1     g4167(.I(new_n4179_), .ZN(new_n4221_));
  NOR2_X1    g4168(.A1(new_n3976_), .A2(new_n4221_), .ZN(new_n4222_));
  NAND3_X1   g4169(.A1(new_n409_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n4223_));
  NOR4_X1    g4170(.A1(new_n4223_), .A2(new_n277_), .A3(new_n649_), .A4(new_n399_), .ZN(new_n4224_));
  NOR4_X1    g4171(.A1(new_n482_), .A2(new_n311_), .A3(new_n341_), .A4(new_n548_), .ZN(new_n4225_));
  AND2_X2    g4172(.A1(new_n4224_), .A2(new_n4225_), .Z(new_n4226_));
  NAND4_X1   g4173(.A1(new_n1226_), .A2(new_n313_), .A3(new_n820_), .A4(new_n332_), .ZN(new_n4227_));
  NOR4_X1    g4174(.A1(new_n4227_), .A2(new_n201_), .A3(new_n243_), .A4(new_n281_), .ZN(new_n4228_));
  NAND4_X1   g4175(.A1(new_n4226_), .A2(new_n1234_), .A3(new_n2862_), .A4(new_n4228_), .ZN(new_n4229_));
  XNOR2_X1   g4176(.A1(new_n4222_), .A2(new_n4229_), .ZN(new_n4230_));
  NOR3_X1    g4177(.A1(new_n4187_), .A2(new_n4188_), .A3(new_n4230_), .ZN(new_n4231_));
  XOR2_X1    g4178(.A1(new_n4222_), .A2(new_n4229_), .Z(new_n4232_));
  AOI21_X1   g4179(.A1(new_n4183_), .A2(new_n4184_), .B(new_n4232_), .ZN(new_n4233_));
  NOR2_X1    g4180(.A1(new_n4231_), .A2(new_n4233_), .ZN(new_n4234_));
  NOR3_X1    g4181(.A1(new_n4234_), .A2(new_n4192_), .A3(new_n4196_), .ZN(new_n4235_));
  INV_X1     g4182(.I(new_n4193_), .ZN(new_n4236_));
  NAND2_X1   g4183(.A1(new_n4236_), .A2(new_n4194_), .ZN(new_n4237_));
  NAND3_X1   g4184(.A1(new_n4183_), .A2(new_n4184_), .A3(new_n4232_), .ZN(new_n4238_));
  OAI21_X1   g4185(.A1(new_n4187_), .A2(new_n4188_), .B(new_n4230_), .ZN(new_n4239_));
  NAND2_X1   g4186(.A1(new_n4239_), .A2(new_n4238_), .ZN(new_n4240_));
  AOI21_X1   g4187(.A1(new_n4240_), .A2(new_n4237_), .B(new_n4182_), .ZN(new_n4241_));
  OAI21_X1   g4188(.A1(new_n4235_), .A2(new_n4241_), .B(new_n2940_), .ZN(new_n4242_));
  NOR2_X1    g4189(.A1(new_n4182_), .A2(new_n3987_), .ZN(new_n4243_));
  OAI22_X1   g4190(.A1(new_n4243_), .A2(new_n3739_), .B1(new_n4230_), .B2(new_n2939_), .ZN(new_n4244_));
  INV_X1     g4191(.I(new_n4244_), .ZN(new_n4245_));
  OAI21_X1   g4192(.A1(new_n3182_), .A2(new_n2972_), .B(new_n4095_), .ZN(new_n4246_));
  NAND3_X1   g4193(.A1(new_n2875_), .A2(new_n2878_), .A3(new_n2977_), .ZN(new_n4247_));
  AOI21_X1   g4194(.A1(new_n4246_), .A2(new_n4247_), .B(new_n803_), .ZN(new_n4248_));
  NOR4_X1    g4195(.A1(new_n3581_), .A2(new_n3580_), .A3(new_n4248_), .A4(new_n2969_), .ZN(new_n4249_));
  AOI21_X1   g4196(.A1(new_n2701_), .A2(new_n3076_), .B(new_n4099_), .ZN(new_n4250_));
  NOR3_X1    g4197(.A1(new_n2930_), .A2(new_n2929_), .A3(new_n2969_), .ZN(new_n4251_));
  OAI21_X1   g4198(.A1(new_n4250_), .A2(new_n4251_), .B(new_n802_), .ZN(new_n4252_));
  AOI22_X1   g4199(.A1(new_n3570_), .A2(new_n3566_), .B1(new_n4252_), .B2(new_n2977_), .ZN(new_n4253_));
  NOR2_X1    g4200(.A1(new_n4253_), .A2(new_n4249_), .ZN(new_n4254_));
  NOR2_X1    g4201(.A1(new_n2734_), .A2(new_n3028_), .ZN(new_n4255_));
  INV_X1     g4202(.I(new_n4255_), .ZN(new_n4256_));
  NAND2_X1   g4203(.A1(new_n2720_), .A2(new_n3030_), .ZN(new_n4257_));
  AOI22_X1   g4204(.A1(new_n4257_), .A2(new_n4256_), .B1(new_n3189_), .B2(new_n3038_), .ZN(new_n4258_));
  OAI21_X1   g4205(.A1(new_n4258_), .A2(new_n702_), .B(new_n2992_), .ZN(new_n4259_));
  NOR2_X1    g4206(.A1(new_n3235_), .A2(new_n4259_), .ZN(new_n4260_));
  AND2_X2    g4207(.A1(new_n3235_), .A2(new_n4259_), .Z(new_n4261_));
  NOR2_X1    g4208(.A1(new_n2792_), .A2(new_n438_), .ZN(new_n4262_));
  OAI21_X1   g4209(.A1(new_n4133_), .A2(new_n4122_), .B(new_n4262_), .ZN(new_n4263_));
  INV_X1     g4210(.I(new_n4262_), .ZN(new_n4264_));
  NAND3_X1   g4211(.A1(new_n4119_), .A2(new_n4123_), .A3(new_n4264_), .ZN(new_n4265_));
  NAND2_X1   g4212(.A1(new_n4263_), .A2(new_n4265_), .ZN(new_n4266_));
  NAND4_X1   g4213(.A1(new_n4119_), .A2(new_n437_), .A3(new_n2783_), .A4(new_n4123_), .ZN(new_n4267_));
  OAI21_X1   g4214(.A1(new_n4266_), .A2(new_n4118_), .B(new_n4267_), .ZN(new_n4268_));
  AOI21_X1   g4215(.A1(new_n3510_), .A2(new_n3509_), .B(new_n3501_), .ZN(new_n4269_));
  INV_X1     g4216(.I(new_n3396_), .ZN(new_n4270_));
  AOI22_X1   g4217(.A1(new_n2758_), .A2(new_n3494_), .B1(new_n2791_), .B2(new_n4270_), .ZN(new_n4271_));
  NOR2_X1    g4218(.A1(new_n2743_), .A2(new_n3496_), .ZN(new_n4272_));
  OR2_X2     g4219(.A1(new_n4272_), .A2(new_n4271_), .Z(new_n4273_));
  OAI22_X1   g4220(.A1(new_n4269_), .A2(new_n4273_), .B1(new_n438_), .B2(new_n2770_), .ZN(new_n4274_));
  OAI21_X1   g4221(.A1(new_n2960_), .A2(new_n2963_), .B(new_n3393_), .ZN(new_n4275_));
  NOR2_X1    g4222(.A1(new_n4272_), .A2(new_n4271_), .ZN(new_n4276_));
  NOR2_X1    g4223(.A1(new_n2770_), .A2(new_n438_), .ZN(new_n4277_));
  NAND3_X1   g4224(.A1(new_n4275_), .A2(new_n4276_), .A3(new_n4277_), .ZN(new_n4278_));
  NAND2_X1   g4225(.A1(new_n4274_), .A2(new_n4278_), .ZN(new_n4279_));
  XOR2_X1    g4226(.A1(new_n4268_), .A2(new_n4279_), .Z(new_n4280_));
  OAI21_X1   g4227(.A1(new_n4261_), .A2(new_n4260_), .B(new_n4280_), .ZN(new_n4281_));
  INV_X1     g4228(.I(new_n4260_), .ZN(new_n4282_));
  NAND2_X1   g4229(.A1(new_n3235_), .A2(new_n4259_), .ZN(new_n4283_));
  INV_X1     g4230(.I(new_n4267_), .ZN(new_n4284_));
  AOI21_X1   g4231(.A1(new_n4119_), .A2(new_n4123_), .B(new_n4264_), .ZN(new_n4285_));
  NOR3_X1    g4232(.A1(new_n4133_), .A2(new_n4122_), .A3(new_n4262_), .ZN(new_n4286_));
  NOR3_X1    g4233(.A1(new_n4118_), .A2(new_n4286_), .A3(new_n4285_), .ZN(new_n4287_));
  OAI21_X1   g4234(.A1(new_n4284_), .A2(new_n4287_), .B(new_n4279_), .ZN(new_n4288_));
  NOR2_X1    g4235(.A1(new_n4287_), .A2(new_n4284_), .ZN(new_n4289_));
  AOI21_X1   g4236(.A1(new_n4275_), .A2(new_n4276_), .B(new_n4277_), .ZN(new_n4290_));
  NOR4_X1    g4237(.A1(new_n4269_), .A2(new_n4273_), .A3(new_n438_), .A4(new_n2770_), .ZN(new_n4291_));
  NOR2_X1    g4238(.A1(new_n4291_), .A2(new_n4290_), .ZN(new_n4292_));
  NAND2_X1   g4239(.A1(new_n4289_), .A2(new_n4292_), .ZN(new_n4293_));
  NAND2_X1   g4240(.A1(new_n4293_), .A2(new_n4288_), .ZN(new_n4294_));
  NAND3_X1   g4241(.A1(new_n4282_), .A2(new_n4294_), .A3(new_n4283_), .ZN(new_n4295_));
  AOI21_X1   g4242(.A1(new_n4105_), .A2(new_n4152_), .B(new_n4137_), .ZN(new_n4296_));
  NAND3_X1   g4243(.A1(new_n4296_), .A2(new_n4295_), .A3(new_n4281_), .ZN(new_n4297_));
  INV_X1     g4244(.I(new_n4280_), .ZN(new_n4298_));
  AOI21_X1   g4245(.A1(new_n4282_), .A2(new_n4283_), .B(new_n4298_), .ZN(new_n4299_));
  INV_X1     g4246(.I(new_n4294_), .ZN(new_n4300_));
  NOR3_X1    g4247(.A1(new_n4261_), .A2(new_n4260_), .A3(new_n4300_), .ZN(new_n4301_));
  AOI21_X1   g4248(.A1(new_n3934_), .A2(new_n4104_), .B(new_n4141_), .ZN(new_n4302_));
  OAI22_X1   g4249(.A1(new_n4302_), .A2(new_n4137_), .B1(new_n4299_), .B2(new_n4301_), .ZN(new_n4303_));
  NAND3_X1   g4250(.A1(new_n4303_), .A2(new_n4254_), .A3(new_n4297_), .ZN(new_n4304_));
  NAND4_X1   g4251(.A1(new_n3570_), .A2(new_n3566_), .A3(new_n4252_), .A4(new_n2977_), .ZN(new_n4305_));
  OAI22_X1   g4252(.A1(new_n3581_), .A2(new_n3580_), .B1(new_n4248_), .B2(new_n2969_), .ZN(new_n4306_));
  NAND2_X1   g4253(.A1(new_n4306_), .A2(new_n4305_), .ZN(new_n4307_));
  NOR4_X1    g4254(.A1(new_n4302_), .A2(new_n4299_), .A3(new_n4301_), .A4(new_n4137_), .ZN(new_n4308_));
  AOI21_X1   g4255(.A1(new_n4281_), .A2(new_n4295_), .B(new_n4296_), .ZN(new_n4309_));
  OAI21_X1   g4256(.A1(new_n4309_), .A2(new_n4308_), .B(new_n4307_), .ZN(new_n4310_));
  OAI22_X1   g4257(.A1(new_n4150_), .A2(new_n3938_), .B1(new_n4154_), .B2(new_n4153_), .ZN(new_n4311_));
  OAI22_X1   g4258(.A1(new_n4311_), .A2(new_n4158_), .B1(new_n3942_), .B2(new_n4103_), .ZN(new_n4312_));
  NAND3_X1   g4259(.A1(new_n4312_), .A2(new_n4304_), .A3(new_n4310_), .ZN(new_n4313_));
  NAND2_X1   g4260(.A1(new_n4310_), .A2(new_n4304_), .ZN(new_n4314_));
  AOI21_X1   g4261(.A1(new_n3545_), .A2(new_n3551_), .B(new_n3554_), .ZN(new_n4315_));
  AOI22_X1   g4262(.A1(new_n3942_), .A2(new_n4103_), .B1(new_n4146_), .B2(new_n4142_), .ZN(new_n4316_));
  AOI22_X1   g4263(.A1(new_n4316_), .A2(new_n4315_), .B1(new_n3938_), .B2(new_n4150_), .ZN(new_n4317_));
  NAND2_X1   g4264(.A1(new_n4314_), .A2(new_n4317_), .ZN(new_n4318_));
  NAND2_X1   g4265(.A1(new_n2946_), .A2(new_n3210_), .ZN(new_n4319_));
  NAND2_X1   g4266(.A1(new_n2898_), .A2(new_n3308_), .ZN(new_n4320_));
  AOI22_X1   g4267(.A1(new_n4319_), .A2(new_n4320_), .B1(new_n3216_), .B2(new_n3597_), .ZN(new_n4321_));
  OAI21_X1   g4268(.A1(new_n4321_), .A2(new_n1051_), .B(new_n3280_), .ZN(new_n4322_));
  XOR2_X1    g4269(.A1(new_n3607_), .A2(new_n4322_), .Z(new_n4323_));
  NAND3_X1   g4270(.A1(new_n4318_), .A2(new_n4313_), .A3(new_n4323_), .ZN(new_n4324_));
  NOR2_X1    g4271(.A1(new_n4314_), .A2(new_n4317_), .ZN(new_n4325_));
  NOR3_X1    g4272(.A1(new_n4309_), .A2(new_n4308_), .A3(new_n4307_), .ZN(new_n4326_));
  AOI21_X1   g4273(.A1(new_n4303_), .A2(new_n4297_), .B(new_n4254_), .ZN(new_n4327_));
  NOR2_X1    g4274(.A1(new_n4326_), .A2(new_n4327_), .ZN(new_n4328_));
  NOR2_X1    g4275(.A1(new_n4328_), .A2(new_n4312_), .ZN(new_n4329_));
  XNOR2_X1   g4276(.A1(new_n3607_), .A2(new_n4322_), .ZN(new_n4330_));
  OAI21_X1   g4277(.A1(new_n4325_), .A2(new_n4329_), .B(new_n4330_), .ZN(new_n4331_));
  AOI22_X1   g4278(.A1(new_n4242_), .A2(new_n4245_), .B1(new_n4331_), .B2(new_n4324_), .ZN(new_n4332_));
  NAND3_X1   g4279(.A1(new_n4240_), .A2(new_n4182_), .A3(new_n4237_), .ZN(new_n4333_));
  OAI21_X1   g4280(.A1(new_n4234_), .A2(new_n4196_), .B(new_n4192_), .ZN(new_n4334_));
  AOI21_X1   g4281(.A1(new_n4334_), .A2(new_n4333_), .B(new_n2939_), .ZN(new_n4335_));
  NOR3_X1    g4282(.A1(new_n4325_), .A2(new_n4329_), .A3(new_n4330_), .ZN(new_n4336_));
  AOI21_X1   g4283(.A1(new_n4318_), .A2(new_n4313_), .B(new_n4323_), .ZN(new_n4337_));
  NOR4_X1    g4284(.A1(new_n4335_), .A2(new_n4336_), .A3(new_n4337_), .A4(new_n4244_), .ZN(new_n4338_));
  NOR2_X1    g4285(.A1(new_n4332_), .A2(new_n4338_), .ZN(new_n4339_));
  NOR2_X1    g4286(.A1(new_n4220_), .A2(new_n4339_), .ZN(new_n4340_));
  NAND3_X1   g4287(.A1(new_n4168_), .A2(new_n4083_), .A3(new_n4218_), .ZN(new_n4341_));
  OAI22_X1   g4288(.A1(new_n4335_), .A2(new_n4244_), .B1(new_n4336_), .B2(new_n4337_), .ZN(new_n4342_));
  NAND4_X1   g4289(.A1(new_n4242_), .A2(new_n4331_), .A3(new_n4324_), .A4(new_n4245_), .ZN(new_n4343_));
  NAND2_X1   g4290(.A1(new_n4342_), .A2(new_n4343_), .ZN(new_n4344_));
  AOI21_X1   g4291(.A1(new_n4341_), .A2(new_n4162_), .B(new_n4344_), .ZN(new_n4345_));
  OAI21_X1   g4292(.A1(new_n4345_), .A2(new_n4340_), .B(new_n2942_), .ZN(new_n4346_));
  NAND3_X1   g4293(.A1(new_n4341_), .A2(new_n4162_), .A3(new_n4344_), .ZN(new_n4347_));
  NAND2_X1   g4294(.A1(new_n4220_), .A2(new_n4339_), .ZN(new_n4348_));
  NAND3_X1   g4295(.A1(new_n4348_), .A2(new_n4347_), .A3(new_n2943_), .ZN(new_n4349_));
  NAND2_X1   g4296(.A1(new_n4346_), .A2(new_n4349_), .ZN(new_n4350_));
  NAND3_X1   g4297(.A1(new_n4214_), .A2(new_n4350_), .A3(new_n4216_), .ZN(new_n4351_));
  NOR2_X1    g4298(.A1(new_n4170_), .A2(new_n4173_), .ZN(new_n4352_));
  AOI21_X1   g4299(.A1(new_n4348_), .A2(new_n4347_), .B(new_n2943_), .ZN(new_n4353_));
  NOR3_X1    g4300(.A1(new_n4345_), .A2(new_n4340_), .A3(new_n2942_), .ZN(new_n4354_));
  NOR2_X1    g4301(.A1(new_n4354_), .A2(new_n4353_), .ZN(new_n4355_));
  NOR2_X1    g4302(.A1(new_n4352_), .A2(new_n4202_), .ZN(new_n4356_));
  INV_X1     g4303(.I(new_n4356_), .ZN(new_n4357_));
  AOI21_X1   g4304(.A1(new_n4351_), .A2(new_n4357_), .B(new_n4078_), .ZN(new_n4358_));
  INV_X1     g4305(.I(new_n4078_), .ZN(new_n4359_));
  NOR2_X1    g4306(.A1(new_n4352_), .A2(new_n4202_), .ZN(new_n4360_));
  NOR3_X1    g4307(.A1(new_n4208_), .A2(new_n4355_), .A3(new_n4360_), .ZN(new_n4361_));
  NOR3_X1    g4308(.A1(new_n4361_), .A2(new_n4359_), .A3(new_n4356_), .ZN(new_n4362_));
  NOR2_X1    g4309(.A1(new_n4362_), .A2(new_n4358_), .ZN(new_n4363_));
  NOR2_X1    g4310(.A1(new_n308_), .A2(new_n294_), .ZN(new_n4364_));
  NAND3_X1   g4311(.A1(new_n2238_), .A2(new_n2920_), .A3(new_n4058_), .ZN(new_n4365_));
  NAND4_X1   g4312(.A1(new_n357_), .A2(new_n218_), .A3(new_n407_), .A4(new_n548_), .ZN(new_n4366_));
  NOR4_X1    g4313(.A1(new_n4366_), .A2(new_n482_), .A3(new_n674_), .A4(new_n4365_), .ZN(new_n4367_));
  AND3_X2    g4314(.A1(new_n4367_), .A2(new_n4364_), .A3(new_n2278_), .Z(new_n4368_));
  INV_X1     g4315(.I(new_n4368_), .ZN(new_n4369_));
  NAND2_X1   g4316(.A1(new_n4363_), .A2(new_n4369_), .ZN(new_n4370_));
  OAI21_X1   g4317(.A1(new_n4362_), .A2(new_n4358_), .B(new_n4368_), .ZN(new_n4371_));
  NAND2_X1   g4318(.A1(new_n4370_), .A2(new_n4371_), .ZN(new_n4372_));
  NAND3_X1   g4319(.A1(new_n4053_), .A2(new_n4038_), .A3(new_n4214_), .ZN(new_n4373_));
  AOI21_X1   g4320(.A1(new_n4011_), .A2(new_n4010_), .B(new_n4009_), .ZN(new_n4374_));
  NOR3_X1    g4321(.A1(new_n3853_), .A2(new_n3997_), .A3(new_n3993_), .ZN(new_n4375_));
  NOR2_X1    g4322(.A1(new_n4374_), .A2(new_n4375_), .ZN(new_n4376_));
  AOI21_X1   g4323(.A1(new_n4025_), .A2(new_n4024_), .B(new_n4023_), .ZN(new_n4377_));
  NOR3_X1    g4324(.A1(new_n4016_), .A2(new_n4021_), .A3(new_n3856_), .ZN(new_n4378_));
  OAI21_X1   g4325(.A1(new_n4378_), .A2(new_n4377_), .B(new_n4035_), .ZN(new_n4379_));
  NOR2_X1    g4326(.A1(new_n4379_), .A2(new_n4376_), .ZN(new_n4380_));
  AOI21_X1   g4327(.A1(new_n4379_), .A2(new_n4376_), .B(new_n4051_), .ZN(new_n4381_));
  OAI21_X1   g4328(.A1(new_n4381_), .A2(new_n4380_), .B(new_n4208_), .ZN(new_n4382_));
  AOI21_X1   g4329(.A1(new_n4382_), .A2(new_n4373_), .B(new_n4078_), .ZN(new_n4383_));
  NOR3_X1    g4330(.A1(new_n4381_), .A2(new_n4380_), .A3(new_n4208_), .ZN(new_n4384_));
  AOI21_X1   g4331(.A1(new_n4053_), .A2(new_n4038_), .B(new_n4214_), .ZN(new_n4385_));
  NOR3_X1    g4332(.A1(new_n4384_), .A2(new_n4385_), .A3(new_n4359_), .ZN(new_n4386_));
  OAI21_X1   g4333(.A1(new_n4386_), .A2(new_n4383_), .B(new_n4074_), .ZN(new_n4387_));
  OAI21_X1   g4334(.A1(new_n4384_), .A2(new_n4385_), .B(new_n4359_), .ZN(new_n4388_));
  NAND3_X1   g4335(.A1(new_n4382_), .A2(new_n4373_), .A3(new_n4078_), .ZN(new_n4389_));
  NAND3_X1   g4336(.A1(new_n4388_), .A2(new_n4389_), .A3(new_n4073_), .ZN(new_n4390_));
  NAND2_X1   g4337(.A1(new_n4387_), .A2(new_n4390_), .ZN(new_n4391_));
  NAND2_X1   g4338(.A1(new_n4391_), .A2(new_n4372_), .ZN(new_n4392_));
  INV_X1     g4339(.I(new_n4372_), .ZN(new_n4393_));
  NAND3_X1   g4340(.A1(new_n4393_), .A2(new_n4387_), .A3(new_n4390_), .ZN(new_n4394_));
  AOI21_X1   g4341(.A1(new_n4392_), .A2(new_n4394_), .B(new_n4211_), .ZN(new_n4395_));
  OAI21_X1   g4342(.A1(new_n4381_), .A2(new_n4380_), .B(new_n4073_), .ZN(new_n4396_));
  NOR3_X1    g4343(.A1(new_n4381_), .A2(new_n4380_), .A3(new_n4073_), .ZN(new_n4397_));
  OAI21_X1   g4344(.A1(new_n4397_), .A2(new_n4209_), .B(new_n4396_), .ZN(new_n4398_));
  NAND2_X1   g4345(.A1(new_n4391_), .A2(new_n4393_), .ZN(new_n4399_));
  NAND3_X1   g4346(.A1(new_n4387_), .A2(new_n4390_), .A3(new_n4372_), .ZN(new_n4400_));
  AOI21_X1   g4347(.A1(new_n4399_), .A2(new_n4400_), .B(new_n4398_), .ZN(new_n4401_));
  NOR2_X1    g4348(.A1(new_n4395_), .A2(new_n4401_), .ZN(new_n4402_));
  INV_X1     g4349(.I(new_n4402_), .ZN(\sin[0] ));
  XOR2_X1    g4350(.A1(\a[22] ), .A2(\a[23] ), .Z(new_n4404_));
  NAND2_X1   g4351(.A1(new_n4372_), .A2(new_n4398_), .ZN(new_n4405_));
  NAND3_X1   g4352(.A1(new_n4211_), .A2(new_n4370_), .A3(new_n4371_), .ZN(new_n4406_));
  NAND2_X1   g4353(.A1(new_n4405_), .A2(new_n4406_), .ZN(new_n4407_));
  NAND3_X1   g4354(.A1(new_n4407_), .A2(new_n4387_), .A3(new_n4390_), .ZN(new_n4408_));
  NAND2_X1   g4355(.A1(new_n4331_), .A2(new_n4324_), .ZN(new_n4409_));
  XOR2_X1    g4356(.A1(new_n4409_), .A2(new_n2943_), .Z(new_n4410_));
  INV_X1     g4357(.I(new_n4220_), .ZN(new_n4411_));
  NOR2_X1    g4358(.A1(new_n4335_), .A2(new_n4244_), .ZN(new_n4412_));
  NOR2_X1    g4359(.A1(new_n4411_), .A2(new_n4412_), .ZN(new_n4413_));
  NOR3_X1    g4360(.A1(new_n4220_), .A2(new_n4335_), .A3(new_n4244_), .ZN(new_n4414_));
  OAI21_X1   g4361(.A1(new_n4413_), .A2(new_n4414_), .B(new_n4410_), .ZN(new_n4415_));
  OAI21_X1   g4362(.A1(new_n4355_), .A2(new_n4202_), .B(new_n4352_), .ZN(new_n4416_));
  NOR3_X1    g4363(.A1(new_n4354_), .A2(new_n4353_), .A3(new_n4206_), .ZN(new_n4417_));
  NOR2_X1    g4364(.A1(new_n4359_), .A2(new_n4417_), .ZN(new_n4418_));
  NAND3_X1   g4365(.A1(new_n4418_), .A2(new_n4416_), .A3(new_n4415_), .ZN(new_n4419_));
  INV_X1     g4366(.I(new_n4415_), .ZN(new_n4420_));
  AOI21_X1   g4367(.A1(new_n4350_), .A2(new_n4206_), .B(new_n4215_), .ZN(new_n4421_));
  OAI21_X1   g4368(.A1(new_n4350_), .A2(new_n4206_), .B(new_n4078_), .ZN(new_n4422_));
  OAI21_X1   g4369(.A1(new_n4421_), .A2(new_n4422_), .B(new_n4420_), .ZN(new_n4423_));
  NAND2_X1   g4370(.A1(new_n4419_), .A2(new_n4423_), .ZN(new_n4424_));
  OAI21_X1   g4371(.A1(new_n4362_), .A2(new_n4358_), .B(new_n4369_), .ZN(new_n4425_));
  OAI21_X1   g4372(.A1(new_n4361_), .A2(new_n4356_), .B(new_n4359_), .ZN(new_n4426_));
  NAND3_X1   g4373(.A1(new_n4351_), .A2(new_n4078_), .A3(new_n4357_), .ZN(new_n4427_));
  NAND3_X1   g4374(.A1(new_n4426_), .A2(new_n4427_), .A3(new_n4368_), .ZN(new_n4428_));
  NAND2_X1   g4375(.A1(new_n4425_), .A2(new_n4428_), .ZN(new_n4429_));
  NAND3_X1   g4376(.A1(new_n4429_), .A2(new_n4371_), .A3(new_n4424_), .ZN(new_n4430_));
  NOR2_X1    g4377(.A1(new_n4421_), .A2(new_n4422_), .ZN(new_n4431_));
  NOR2_X1    g4378(.A1(new_n4363_), .A2(new_n4369_), .ZN(new_n4432_));
  INV_X1     g4379(.I(new_n4432_), .ZN(new_n4433_));
  AOI21_X1   g4380(.A1(new_n4430_), .A2(new_n4433_), .B(new_n4398_), .ZN(new_n4434_));
  INV_X1     g4381(.I(new_n4371_), .ZN(new_n4435_));
  AOI21_X1   g4382(.A1(new_n4426_), .A2(new_n4427_), .B(new_n4368_), .ZN(new_n4436_));
  NOR3_X1    g4383(.A1(new_n4362_), .A2(new_n4358_), .A3(new_n4369_), .ZN(new_n4437_));
  OAI21_X1   g4384(.A1(new_n4437_), .A2(new_n4436_), .B(new_n4424_), .ZN(new_n4438_));
  NOR2_X1    g4385(.A1(new_n4438_), .A2(new_n4435_), .ZN(new_n4439_));
  NOR3_X1    g4386(.A1(new_n4439_), .A2(new_n4211_), .A3(new_n4432_), .ZN(new_n4440_));
  NOR2_X1    g4387(.A1(new_n4440_), .A2(new_n4434_), .ZN(new_n4441_));
  NOR2_X1    g4388(.A1(new_n4408_), .A2(new_n4441_), .ZN(new_n4442_));
  XOR2_X1    g4389(.A1(new_n4442_), .A2(new_n4404_), .Z(new_n4443_));
  XOR2_X1    g4390(.A1(new_n4443_), .A2(new_n4402_), .Z(\sin[1] ));
  INV_X1     g4391(.I(new_n4404_), .ZN(new_n4445_));
  INV_X1     g4392(.I(new_n4442_), .ZN(new_n4446_));
  NAND2_X1   g4393(.A1(new_n4408_), .A2(new_n4441_), .ZN(new_n4447_));
  NAND2_X1   g4394(.A1(new_n4446_), .A2(new_n4447_), .ZN(new_n4448_));
  NAND2_X1   g4395(.A1(new_n4448_), .A2(new_n4402_), .ZN(new_n4449_));
  NAND2_X1   g4396(.A1(new_n4418_), .A2(new_n4416_), .ZN(new_n4450_));
  NOR2_X1    g4397(.A1(new_n4450_), .A2(new_n4415_), .ZN(new_n4451_));
  NOR3_X1    g4398(.A1(new_n4421_), .A2(new_n4422_), .A3(new_n4420_), .ZN(new_n4452_));
  AOI21_X1   g4399(.A1(new_n4418_), .A2(new_n4416_), .B(new_n4415_), .ZN(new_n4453_));
  NOR2_X1    g4400(.A1(new_n4453_), .A2(new_n4452_), .ZN(new_n4454_));
  OAI21_X1   g4401(.A1(new_n4454_), .A2(new_n4363_), .B(new_n4369_), .ZN(new_n4455_));
  NAND2_X1   g4402(.A1(new_n4454_), .A2(new_n4363_), .ZN(new_n4456_));
  NAND3_X1   g4403(.A1(new_n4455_), .A2(new_n4398_), .A3(new_n4456_), .ZN(new_n4457_));
  NOR2_X1    g4404(.A1(new_n4185_), .A2(new_n3977_), .ZN(new_n4458_));
  AOI21_X1   g4405(.A1(new_n4458_), .A2(new_n4182_), .B(new_n4230_), .ZN(new_n4459_));
  NOR3_X1    g4406(.A1(new_n4189_), .A2(new_n3987_), .A3(new_n4182_), .ZN(new_n4460_));
  NOR2_X1    g4407(.A1(new_n4459_), .A2(new_n4460_), .ZN(new_n4461_));
  NAND2_X1   g4408(.A1(new_n4222_), .A2(new_n2447_), .ZN(new_n4462_));
  NAND3_X1   g4409(.A1(new_n359_), .A2(new_n439_), .A3(new_n376_), .ZN(new_n4463_));
  NAND2_X1   g4410(.A1(new_n2231_), .A2(new_n380_), .ZN(new_n4464_));
  NAND2_X1   g4411(.A1(new_n2451_), .A2(new_n603_), .ZN(new_n4465_));
  NOR4_X1    g4412(.A1(new_n4464_), .A2(new_n4465_), .A3(new_n507_), .A4(new_n4463_), .ZN(new_n4466_));
  INV_X1     g4413(.I(new_n4466_), .ZN(new_n4467_));
  NOR4_X1    g4414(.A1(new_n625_), .A2(new_n292_), .A3(new_n383_), .A4(new_n517_), .ZN(new_n4468_));
  NOR4_X1    g4415(.A1(new_n453_), .A2(new_n160_), .A3(new_n256_), .A4(new_n609_), .ZN(new_n4469_));
  NAND4_X1   g4416(.A1(new_n324_), .A2(new_n1436_), .A3(new_n4468_), .A4(new_n4469_), .ZN(new_n4470_));
  NOR3_X1    g4417(.A1(new_n4229_), .A2(new_n4467_), .A3(new_n4470_), .ZN(new_n4471_));
  AND2_X2    g4418(.A1(new_n4462_), .A2(new_n4471_), .Z(new_n4472_));
  NOR2_X1    g4419(.A1(new_n4462_), .A2(new_n4471_), .ZN(new_n4473_));
  NOR2_X1    g4420(.A1(new_n4472_), .A2(new_n4473_), .ZN(new_n4474_));
  INV_X1     g4421(.I(new_n4474_), .ZN(new_n4475_));
  NAND2_X1   g4422(.A1(new_n4475_), .A2(new_n4230_), .ZN(new_n4476_));
  NAND2_X1   g4423(.A1(new_n4474_), .A2(new_n4232_), .ZN(new_n4477_));
  AOI21_X1   g4424(.A1(new_n4476_), .A2(new_n4477_), .B(new_n4461_), .ZN(new_n4478_));
  INV_X1     g4425(.I(new_n4461_), .ZN(new_n4479_));
  NOR2_X1    g4426(.A1(new_n4474_), .A2(new_n4230_), .ZN(new_n4480_));
  NOR2_X1    g4427(.A1(new_n4475_), .A2(new_n4232_), .ZN(new_n4481_));
  NOR2_X1    g4428(.A1(new_n4481_), .A2(new_n4480_), .ZN(new_n4482_));
  NOR2_X1    g4429(.A1(new_n4479_), .A2(new_n4482_), .ZN(new_n4483_));
  NOR2_X1    g4430(.A1(new_n4483_), .A2(new_n4478_), .ZN(new_n4484_));
  OAI22_X1   g4431(.A1(new_n4230_), .A2(new_n3639_), .B1(new_n4182_), .B2(new_n3636_), .ZN(new_n4485_));
  NOR2_X1    g4432(.A1(new_n4474_), .A2(new_n2939_), .ZN(new_n4486_));
  INV_X1     g4433(.I(new_n4486_), .ZN(new_n4487_));
  NAND2_X1   g4434(.A1(new_n4487_), .A2(new_n4485_), .ZN(new_n4488_));
  AOI21_X1   g4435(.A1(new_n4488_), .A2(new_n2942_), .B(new_n2939_), .ZN(new_n4489_));
  XOR2_X1    g4436(.A1(new_n4484_), .A2(new_n4489_), .Z(new_n4490_));
  NOR2_X1    g4437(.A1(new_n4415_), .A2(new_n4490_), .ZN(new_n4491_));
  INV_X1     g4438(.I(new_n4491_), .ZN(new_n4492_));
  INV_X1     g4439(.I(new_n4490_), .ZN(new_n4493_));
  NOR2_X1    g4440(.A1(new_n2682_), .A2(new_n2969_), .ZN(new_n4494_));
  INV_X1     g4441(.I(new_n4494_), .ZN(new_n4495_));
  NAND2_X1   g4442(.A1(new_n2898_), .A2(new_n3086_), .ZN(new_n4496_));
  AOI22_X1   g4443(.A1(new_n4496_), .A2(new_n4495_), .B1(new_n2931_), .B2(new_n3076_), .ZN(new_n4497_));
  INV_X1     g4444(.I(new_n4497_), .ZN(new_n4498_));
  AOI21_X1   g4445(.A1(new_n3842_), .A2(new_n3843_), .B(new_n2969_), .ZN(new_n4499_));
  NAND2_X1   g4446(.A1(new_n4295_), .A2(new_n4281_), .ZN(new_n4500_));
  AOI22_X1   g4447(.A1(new_n2720_), .A2(new_n3030_), .B1(new_n2729_), .B2(new_n3038_), .ZN(new_n4501_));
  NOR3_X1    g4448(.A1(new_n3181_), .A2(new_n3180_), .A3(new_n3028_), .ZN(new_n4502_));
  OAI21_X1   g4449(.A1(new_n4501_), .A2(new_n4502_), .B(new_n721_), .ZN(new_n4503_));
  NAND4_X1   g4450(.A1(new_n3868_), .A2(new_n3869_), .A3(new_n4503_), .A4(new_n2992_), .ZN(new_n4504_));
  NAND2_X1   g4451(.A1(new_n2729_), .A2(new_n3038_), .ZN(new_n4505_));
  OAI21_X1   g4452(.A1(new_n3183_), .A2(new_n3031_), .B(new_n4505_), .ZN(new_n4506_));
  NAND3_X1   g4453(.A1(new_n2699_), .A2(new_n2700_), .A3(new_n2998_), .ZN(new_n4507_));
  AOI21_X1   g4454(.A1(new_n4506_), .A2(new_n4507_), .B(new_n702_), .ZN(new_n4508_));
  OAI22_X1   g4455(.A1(new_n3197_), .A2(new_n3201_), .B1(new_n4508_), .B2(new_n2991_), .ZN(new_n4509_));
  NAND2_X1   g4456(.A1(new_n4509_), .A2(new_n4504_), .ZN(new_n4510_));
  NAND3_X1   g4457(.A1(new_n4132_), .A2(new_n4263_), .A3(new_n4265_), .ZN(new_n4511_));
  AOI22_X1   g4458(.A1(new_n4511_), .A2(new_n4267_), .B1(new_n4274_), .B2(new_n4278_), .ZN(new_n4512_));
  NOR4_X1    g4459(.A1(new_n4269_), .A2(new_n4273_), .A3(new_n438_), .A4(new_n2775_), .ZN(new_n4513_));
  AOI22_X1   g4460(.A1(new_n2743_), .A2(new_n3494_), .B1(new_n2758_), .B2(new_n4270_), .ZN(new_n4514_));
  NOR2_X1    g4461(.A1(new_n2813_), .A2(new_n3496_), .ZN(new_n4515_));
  NOR2_X1    g4462(.A1(new_n4515_), .A2(new_n4514_), .ZN(new_n4516_));
  OAI21_X1   g4463(.A1(new_n3128_), .A2(new_n3501_), .B(new_n4516_), .ZN(new_n4517_));
  NOR4_X1    g4464(.A1(new_n4512_), .A2(new_n2791_), .A3(new_n4513_), .A4(new_n4517_), .ZN(new_n4518_));
  AOI21_X1   g4465(.A1(new_n4268_), .A2(new_n4279_), .B(new_n4513_), .ZN(new_n4519_));
  INV_X1     g4466(.I(new_n4517_), .ZN(new_n4520_));
  AOI21_X1   g4467(.A1(new_n4519_), .A2(new_n4520_), .B(new_n2765_), .ZN(new_n4521_));
  OAI21_X1   g4468(.A1(new_n4521_), .A2(new_n4518_), .B(new_n437_), .ZN(new_n4522_));
  INV_X1     g4469(.I(new_n4513_), .ZN(new_n4523_));
  NAND4_X1   g4470(.A1(new_n4288_), .A2(new_n2765_), .A3(new_n4523_), .A4(new_n4520_), .ZN(new_n4524_));
  OAI21_X1   g4471(.A1(new_n4289_), .A2(new_n4292_), .B(new_n4523_), .ZN(new_n4525_));
  OAI21_X1   g4472(.A1(new_n4525_), .A2(new_n4517_), .B(new_n2791_), .ZN(new_n4526_));
  NAND3_X1   g4473(.A1(new_n4526_), .A2(new_n438_), .A3(new_n4524_), .ZN(new_n4527_));
  AOI21_X1   g4474(.A1(new_n4527_), .A2(new_n4522_), .B(new_n4510_), .ZN(new_n4528_));
  NOR4_X1    g4475(.A1(new_n3197_), .A2(new_n3201_), .A3(new_n4508_), .A4(new_n2991_), .ZN(new_n4529_));
  AOI22_X1   g4476(.A1(new_n3868_), .A2(new_n3869_), .B1(new_n4503_), .B2(new_n2992_), .ZN(new_n4530_));
  NOR2_X1    g4477(.A1(new_n4530_), .A2(new_n4529_), .ZN(new_n4531_));
  AOI21_X1   g4478(.A1(new_n4526_), .A2(new_n4524_), .B(new_n438_), .ZN(new_n4532_));
  NOR3_X1    g4479(.A1(new_n4521_), .A2(new_n437_), .A3(new_n4518_), .ZN(new_n4533_));
  NOR3_X1    g4480(.A1(new_n4532_), .A2(new_n4533_), .A3(new_n4531_), .ZN(new_n4534_));
  NOR3_X1    g4481(.A1(new_n4528_), .A2(new_n4534_), .A3(new_n4299_), .ZN(new_n4535_));
  NOR3_X1    g4482(.A1(new_n4535_), .A2(new_n4500_), .A3(new_n4296_), .ZN(new_n4536_));
  NOR2_X1    g4483(.A1(new_n4299_), .A2(new_n4301_), .ZN(new_n4537_));
  INV_X1     g4484(.I(new_n4296_), .ZN(new_n4538_));
  OAI21_X1   g4485(.A1(new_n4532_), .A2(new_n4533_), .B(new_n4531_), .ZN(new_n4539_));
  NAND3_X1   g4486(.A1(new_n4527_), .A2(new_n4522_), .A3(new_n4510_), .ZN(new_n4540_));
  NAND3_X1   g4487(.A1(new_n4539_), .A2(new_n4540_), .A3(new_n4281_), .ZN(new_n4541_));
  AOI21_X1   g4488(.A1(new_n4541_), .A2(new_n4538_), .B(new_n4537_), .ZN(new_n4542_));
  OAI21_X1   g4489(.A1(new_n4536_), .A2(new_n4542_), .B(new_n803_), .ZN(new_n4543_));
  NOR2_X1    g4490(.A1(new_n4543_), .A2(new_n4499_), .ZN(new_n4544_));
  INV_X1     g4491(.I(new_n4499_), .ZN(new_n4545_));
  NAND3_X1   g4492(.A1(new_n4541_), .A2(new_n4537_), .A3(new_n4538_), .ZN(new_n4546_));
  OAI21_X1   g4493(.A1(new_n4535_), .A2(new_n4296_), .B(new_n4500_), .ZN(new_n4547_));
  NAND2_X1   g4494(.A1(new_n4547_), .A2(new_n4546_), .ZN(new_n4548_));
  AOI21_X1   g4495(.A1(new_n4548_), .A2(new_n803_), .B(new_n4545_), .ZN(new_n4549_));
  OAI21_X1   g4496(.A1(new_n4544_), .A2(new_n4549_), .B(new_n4498_), .ZN(new_n4550_));
  NAND3_X1   g4497(.A1(new_n4548_), .A2(new_n803_), .A3(new_n4545_), .ZN(new_n4551_));
  NAND2_X1   g4498(.A1(new_n4543_), .A2(new_n4499_), .ZN(new_n4552_));
  NAND3_X1   g4499(.A1(new_n4552_), .A2(new_n4551_), .A3(new_n4497_), .ZN(new_n4553_));
  NAND3_X1   g4500(.A1(new_n4550_), .A2(new_n4553_), .A3(new_n4304_), .ZN(new_n4554_));
  NAND3_X1   g4501(.A1(new_n4554_), .A2(new_n4328_), .A3(new_n4312_), .ZN(new_n4555_));
  AOI21_X1   g4502(.A1(new_n4552_), .A2(new_n4551_), .B(new_n4497_), .ZN(new_n4556_));
  NOR3_X1    g4503(.A1(new_n4544_), .A2(new_n4549_), .A3(new_n4498_), .ZN(new_n4557_));
  NOR3_X1    g4504(.A1(new_n4557_), .A2(new_n4556_), .A3(new_n4326_), .ZN(new_n4558_));
  OAI21_X1   g4505(.A1(new_n4558_), .A2(new_n4317_), .B(new_n4314_), .ZN(new_n4559_));
  AOI22_X1   g4506(.A1(new_n2946_), .A2(new_n3308_), .B1(new_n3985_), .B2(new_n3210_), .ZN(new_n4560_));
  NOR2_X1    g4507(.A1(new_n3987_), .A2(new_n3237_), .ZN(new_n4561_));
  OAI21_X1   g4508(.A1(new_n4561_), .A2(new_n4560_), .B(new_n1050_), .ZN(new_n4562_));
  NAND2_X1   g4509(.A1(new_n4562_), .A2(new_n3280_), .ZN(new_n4563_));
  XOR2_X1    g4510(.A1(new_n3982_), .A2(new_n4563_), .Z(new_n4564_));
  NAND3_X1   g4511(.A1(new_n4559_), .A2(new_n4555_), .A3(new_n4564_), .ZN(new_n4565_));
  NOR3_X1    g4512(.A1(new_n4558_), .A2(new_n4314_), .A3(new_n4317_), .ZN(new_n4566_));
  AOI21_X1   g4513(.A1(new_n4554_), .A2(new_n4312_), .B(new_n4328_), .ZN(new_n4567_));
  INV_X1     g4514(.I(new_n4564_), .ZN(new_n4568_));
  OAI21_X1   g4515(.A1(new_n4566_), .A2(new_n4567_), .B(new_n4568_), .ZN(new_n4569_));
  NAND2_X1   g4516(.A1(new_n4569_), .A2(new_n4565_), .ZN(new_n4570_));
  NOR2_X1    g4517(.A1(new_n4325_), .A2(new_n4329_), .ZN(new_n4571_));
  XOR2_X1    g4518(.A1(new_n4571_), .A2(new_n4323_), .Z(new_n4572_));
  NAND3_X1   g4519(.A1(new_n4570_), .A2(new_n4331_), .A3(new_n4572_), .ZN(new_n4573_));
  NOR2_X1    g4520(.A1(new_n4571_), .A2(new_n4323_), .ZN(new_n4575_));
  INV_X1     g4521(.I(new_n4575_), .ZN(new_n4576_));
  AOI21_X1   g4522(.A1(new_n4573_), .A2(new_n4576_), .B(new_n4220_), .ZN(new_n4577_));
  NOR3_X1    g4523(.A1(new_n4566_), .A2(new_n4567_), .A3(new_n4568_), .ZN(new_n4578_));
  AOI21_X1   g4524(.A1(new_n4559_), .A2(new_n4555_), .B(new_n4564_), .ZN(new_n4579_));
  OAI21_X1   g4525(.A1(new_n4578_), .A2(new_n4579_), .B(new_n4572_), .ZN(new_n4580_));
  NOR2_X1    g4526(.A1(new_n4580_), .A2(new_n4337_), .ZN(new_n4581_));
  NOR3_X1    g4527(.A1(new_n4581_), .A2(new_n4411_), .A3(new_n4575_), .ZN(new_n4582_));
  OAI22_X1   g4528(.A1(new_n4420_), .A2(new_n4493_), .B1(new_n4582_), .B2(new_n4577_), .ZN(new_n4583_));
  OAI21_X1   g4529(.A1(new_n4450_), .A2(new_n4583_), .B(new_n4492_), .ZN(new_n4584_));
  NAND3_X1   g4530(.A1(new_n4548_), .A2(new_n803_), .A3(new_n4498_), .ZN(new_n4585_));
  NAND2_X1   g4531(.A1(new_n4543_), .A2(new_n4497_), .ZN(new_n4586_));
  AOI21_X1   g4532(.A1(new_n4586_), .A2(new_n4585_), .B(new_n4545_), .ZN(new_n4587_));
  INV_X1     g4533(.I(new_n4587_), .ZN(new_n4588_));
  OAI21_X1   g4534(.A1(new_n4557_), .A2(new_n4556_), .B(new_n4326_), .ZN(new_n4589_));
  NAND2_X1   g4535(.A1(new_n4589_), .A2(new_n4317_), .ZN(new_n4590_));
  NAND2_X1   g4536(.A1(new_n2879_), .A2(new_n3076_), .ZN(new_n4591_));
  AOI22_X1   g4537(.A1(new_n4496_), .A2(new_n4591_), .B1(new_n2946_), .B2(new_n2977_), .ZN(new_n4592_));
  OAI21_X1   g4538(.A1(new_n4592_), .A2(new_n803_), .B(new_n2977_), .ZN(new_n4593_));
  XOR2_X1    g4539(.A1(new_n2935_), .A2(new_n4593_), .Z(new_n4594_));
  INV_X1     g4540(.I(new_n4594_), .ZN(new_n4595_));
  NOR2_X1    g4541(.A1(new_n4308_), .A2(new_n4299_), .ZN(new_n4596_));
  INV_X1     g4542(.I(new_n4596_), .ZN(new_n4597_));
  NAND2_X1   g4543(.A1(new_n4527_), .A2(new_n4522_), .ZN(new_n4598_));
  NAND2_X1   g4544(.A1(new_n4598_), .A2(new_n4510_), .ZN(new_n4599_));
  INV_X1     g4545(.I(new_n4599_), .ZN(new_n4600_));
  NAND2_X1   g4546(.A1(new_n4539_), .A2(new_n4540_), .ZN(new_n4601_));
  NOR2_X1    g4547(.A1(new_n3183_), .A2(new_n3028_), .ZN(new_n4602_));
  NOR2_X1    g4548(.A1(new_n2682_), .A2(new_n3031_), .ZN(new_n4603_));
  OAI22_X1   g4549(.A1(new_n4603_), .A2(new_n4602_), .B1(new_n2701_), .B2(new_n2994_), .ZN(new_n4604_));
  AOI21_X1   g4550(.A1(new_n4604_), .A2(new_n721_), .B(new_n2991_), .ZN(new_n4605_));
  NAND3_X1   g4551(.A1(new_n3463_), .A2(new_n4605_), .A3(new_n3462_), .ZN(new_n4606_));
  INV_X1     g4552(.I(new_n4602_), .ZN(new_n4607_));
  NAND2_X1   g4553(.A1(new_n3436_), .A2(new_n3030_), .ZN(new_n4608_));
  AOI22_X1   g4554(.A1(new_n4608_), .A2(new_n4607_), .B1(new_n3182_), .B2(new_n3038_), .ZN(new_n4609_));
  OAI21_X1   g4555(.A1(new_n4609_), .A2(new_n702_), .B(new_n2992_), .ZN(new_n4610_));
  OAI21_X1   g4556(.A1(new_n3432_), .A2(new_n3440_), .B(new_n4610_), .ZN(new_n4611_));
  NAND2_X1   g4557(.A1(new_n4611_), .A2(new_n4606_), .ZN(new_n4612_));
  NOR2_X1    g4558(.A1(new_n2791_), .A2(new_n437_), .ZN(new_n4613_));
  NAND2_X1   g4559(.A1(new_n4517_), .A2(new_n4613_), .ZN(new_n4614_));
  NAND2_X1   g4560(.A1(new_n3279_), .A2(new_n3393_), .ZN(new_n4615_));
  INV_X1     g4561(.I(new_n4613_), .ZN(new_n4616_));
  NAND3_X1   g4562(.A1(new_n4615_), .A2(new_n4516_), .A3(new_n4616_), .ZN(new_n4617_));
  NAND2_X1   g4563(.A1(new_n4614_), .A2(new_n4617_), .ZN(new_n4618_));
  NOR3_X1    g4564(.A1(new_n4517_), .A2(new_n437_), .A3(new_n2791_), .ZN(new_n4619_));
  INV_X1     g4565(.I(new_n4619_), .ZN(new_n4620_));
  OAI21_X1   g4566(.A1(new_n4519_), .A2(new_n4618_), .B(new_n4620_), .ZN(new_n4621_));
  NOR2_X1    g4567(.A1(new_n3270_), .A2(new_n3501_), .ZN(new_n4622_));
  OAI22_X1   g4568(.A1(new_n2734_), .A2(new_n3493_), .B1(new_n2956_), .B2(new_n3396_), .ZN(new_n4623_));
  OAI21_X1   g4569(.A1(new_n2729_), .A2(new_n3496_), .B(new_n4623_), .ZN(new_n4624_));
  NOR2_X1    g4570(.A1(new_n4622_), .A2(new_n4624_), .ZN(new_n4625_));
  INV_X1     g4571(.I(new_n4625_), .ZN(new_n4626_));
  NOR3_X1    g4572(.A1(new_n4626_), .A2(new_n4621_), .A3(new_n2758_), .ZN(new_n4627_));
  INV_X1     g4573(.I(new_n4621_), .ZN(new_n4628_));
  AOI21_X1   g4574(.A1(new_n4628_), .A2(new_n4625_), .B(new_n2804_), .ZN(new_n4629_));
  OAI21_X1   g4575(.A1(new_n4629_), .A2(new_n4627_), .B(new_n437_), .ZN(new_n4630_));
  NAND3_X1   g4576(.A1(new_n4525_), .A2(new_n4614_), .A3(new_n4617_), .ZN(new_n4631_));
  NAND4_X1   g4577(.A1(new_n4631_), .A2(new_n2804_), .A3(new_n4620_), .A4(new_n4625_), .ZN(new_n4632_));
  OAI21_X1   g4578(.A1(new_n4626_), .A2(new_n4621_), .B(new_n2758_), .ZN(new_n4633_));
  NAND3_X1   g4579(.A1(new_n4633_), .A2(new_n4632_), .A3(new_n438_), .ZN(new_n4634_));
  AOI21_X1   g4580(.A1(new_n4630_), .A2(new_n4634_), .B(new_n4612_), .ZN(new_n4635_));
  NOR3_X1    g4581(.A1(new_n3432_), .A2(new_n3440_), .A3(new_n4610_), .ZN(new_n4636_));
  AOI21_X1   g4582(.A1(new_n3463_), .A2(new_n3462_), .B(new_n4605_), .ZN(new_n4637_));
  NOR2_X1    g4583(.A1(new_n4636_), .A2(new_n4637_), .ZN(new_n4638_));
  AOI21_X1   g4584(.A1(new_n4633_), .A2(new_n4632_), .B(new_n438_), .ZN(new_n4639_));
  NOR3_X1    g4585(.A1(new_n4629_), .A2(new_n437_), .A3(new_n4627_), .ZN(new_n4640_));
  NOR3_X1    g4586(.A1(new_n4640_), .A2(new_n4638_), .A3(new_n4639_), .ZN(new_n4641_));
  OAI21_X1   g4587(.A1(new_n4635_), .A2(new_n4641_), .B(new_n4601_), .ZN(new_n4642_));
  NOR2_X1    g4588(.A1(new_n4642_), .A2(new_n4600_), .ZN(new_n4643_));
  OAI21_X1   g4589(.A1(new_n4640_), .A2(new_n4639_), .B(new_n4638_), .ZN(new_n4644_));
  NAND3_X1   g4590(.A1(new_n4630_), .A2(new_n4612_), .A3(new_n4634_), .ZN(new_n4645_));
  NAND2_X1   g4591(.A1(new_n4644_), .A2(new_n4645_), .ZN(new_n4646_));
  NAND2_X1   g4592(.A1(new_n4598_), .A2(new_n4510_), .ZN(new_n4648_));
  INV_X1     g4593(.I(new_n4648_), .ZN(new_n4649_));
  OAI21_X1   g4594(.A1(new_n4643_), .A2(new_n4649_), .B(new_n4597_), .ZN(new_n4650_));
  NAND3_X1   g4595(.A1(new_n4646_), .A2(new_n4601_), .A3(new_n4599_), .ZN(new_n4651_));
  NAND3_X1   g4596(.A1(new_n4651_), .A2(new_n4596_), .A3(new_n4648_), .ZN(new_n4652_));
  NAND2_X1   g4597(.A1(new_n4650_), .A2(new_n4652_), .ZN(new_n4653_));
  NAND2_X1   g4598(.A1(new_n4653_), .A2(new_n4595_), .ZN(new_n4654_));
  AOI21_X1   g4599(.A1(new_n4590_), .A2(new_n4314_), .B(new_n4654_), .ZN(new_n4655_));
  AOI21_X1   g4600(.A1(new_n4550_), .A2(new_n4553_), .B(new_n4304_), .ZN(new_n4656_));
  OAI21_X1   g4601(.A1(new_n4656_), .A2(new_n4312_), .B(new_n4314_), .ZN(new_n4657_));
  INV_X1     g4602(.I(new_n4654_), .ZN(new_n4658_));
  NOR2_X1    g4603(.A1(new_n4657_), .A2(new_n4658_), .ZN(new_n4659_));
  OAI21_X1   g4604(.A1(new_n4655_), .A2(new_n4659_), .B(new_n4588_), .ZN(new_n4660_));
  NAND2_X1   g4605(.A1(new_n4657_), .A2(new_n4658_), .ZN(new_n4661_));
  NAND3_X1   g4606(.A1(new_n4590_), .A2(new_n4314_), .A3(new_n4654_), .ZN(new_n4662_));
  NAND3_X1   g4607(.A1(new_n4662_), .A2(new_n4661_), .A3(new_n4587_), .ZN(new_n4663_));
  OAI22_X1   g4608(.A1(new_n3987_), .A2(new_n3211_), .B1(new_n3213_), .B2(new_n3597_), .ZN(new_n4664_));
  OAI21_X1   g4609(.A1(new_n3237_), .A2(new_n4192_), .B(new_n4664_), .ZN(new_n4665_));
  AOI21_X1   g4610(.A1(new_n4665_), .A2(new_n1050_), .B(new_n3207_), .ZN(new_n4666_));
  XOR2_X1    g4611(.A1(new_n4198_), .A2(new_n4666_), .Z(new_n4667_));
  NAND3_X1   g4612(.A1(new_n4660_), .A2(new_n4663_), .A3(new_n4667_), .ZN(new_n4668_));
  AOI21_X1   g4613(.A1(new_n4662_), .A2(new_n4661_), .B(new_n4587_), .ZN(new_n4669_));
  NOR3_X1    g4614(.A1(new_n4655_), .A2(new_n4659_), .A3(new_n4588_), .ZN(new_n4670_));
  INV_X1     g4615(.I(new_n4667_), .ZN(new_n4671_));
  OAI21_X1   g4616(.A1(new_n4669_), .A2(new_n4670_), .B(new_n4671_), .ZN(new_n4672_));
  NAND2_X1   g4617(.A1(new_n4672_), .A2(new_n4668_), .ZN(new_n4673_));
  INV_X1     g4618(.I(new_n4673_), .ZN(new_n4674_));
  INV_X1     g4619(.I(new_n4571_), .ZN(new_n4675_));
  AOI21_X1   g4620(.A1(new_n4570_), .A2(new_n4330_), .B(new_n4675_), .ZN(new_n4676_));
  NAND3_X1   g4621(.A1(new_n4569_), .A2(new_n4565_), .A3(new_n4323_), .ZN(new_n4677_));
  NAND2_X1   g4622(.A1(new_n4677_), .A2(new_n4220_), .ZN(new_n4678_));
  OAI21_X1   g4623(.A1(new_n4676_), .A2(new_n4678_), .B(new_n4569_), .ZN(new_n4679_));
  NAND2_X1   g4624(.A1(new_n4674_), .A2(new_n4679_), .ZN(new_n4680_));
  OAI21_X1   g4625(.A1(new_n4578_), .A2(new_n4579_), .B(new_n4330_), .ZN(new_n4681_));
  NAND2_X1   g4626(.A1(new_n4681_), .A2(new_n4571_), .ZN(new_n4682_));
  NOR3_X1    g4627(.A1(new_n4578_), .A2(new_n4579_), .A3(new_n4330_), .ZN(new_n4683_));
  NOR2_X1    g4628(.A1(new_n4683_), .A2(new_n4411_), .ZN(new_n4684_));
  AOI21_X1   g4629(.A1(new_n4684_), .A2(new_n4682_), .B(new_n4579_), .ZN(new_n4685_));
  NAND2_X1   g4630(.A1(new_n4685_), .A2(new_n4673_), .ZN(new_n4686_));
  NAND3_X1   g4631(.A1(new_n4461_), .A2(new_n4232_), .A3(new_n4474_), .ZN(new_n4687_));
  OAI21_X1   g4632(.A1(new_n4461_), .A2(new_n4476_), .B(new_n4687_), .ZN(new_n4688_));
  NOR2_X1    g4633(.A1(new_n4474_), .A2(new_n3639_), .ZN(new_n4689_));
  OAI21_X1   g4634(.A1(new_n4230_), .A2(new_n3636_), .B(new_n2942_), .ZN(new_n4690_));
  OAI21_X1   g4635(.A1(new_n4689_), .A2(new_n4690_), .B(new_n2940_), .ZN(new_n4691_));
  XOR2_X1    g4636(.A1(new_n4688_), .A2(new_n4691_), .Z(new_n4692_));
  AOI21_X1   g4637(.A1(new_n4680_), .A2(new_n4686_), .B(new_n4692_), .ZN(new_n4693_));
  NOR2_X1    g4638(.A1(new_n4685_), .A2(new_n4673_), .ZN(new_n4694_));
  NOR2_X1    g4639(.A1(new_n4674_), .A2(new_n4679_), .ZN(new_n4695_));
  INV_X1     g4640(.I(new_n4692_), .ZN(new_n4696_));
  NOR3_X1    g4641(.A1(new_n4695_), .A2(new_n4694_), .A3(new_n4696_), .ZN(new_n4697_));
  OAI21_X1   g4642(.A1(new_n4693_), .A2(new_n4697_), .B(new_n4584_), .ZN(new_n4698_));
  OAI21_X1   g4643(.A1(new_n4581_), .A2(new_n4575_), .B(new_n4411_), .ZN(new_n4699_));
  NAND3_X1   g4644(.A1(new_n4573_), .A2(new_n4220_), .A3(new_n4576_), .ZN(new_n4700_));
  AOI22_X1   g4645(.A1(new_n4699_), .A2(new_n4700_), .B1(new_n4415_), .B2(new_n4490_), .ZN(new_n4701_));
  AOI21_X1   g4646(.A1(new_n4431_), .A2(new_n4701_), .B(new_n4491_), .ZN(new_n4702_));
  NOR3_X1    g4647(.A1(new_n4695_), .A2(new_n4694_), .A3(new_n4692_), .ZN(new_n4703_));
  AOI21_X1   g4648(.A1(new_n4680_), .A2(new_n4686_), .B(new_n4696_), .ZN(new_n4704_));
  OAI21_X1   g4649(.A1(new_n4703_), .A2(new_n4704_), .B(new_n4702_), .ZN(new_n4705_));
  INV_X1     g4650(.I(new_n2852_), .ZN(new_n4706_));
  NAND4_X1   g4651(.A1(new_n187_), .A2(new_n219_), .A3(new_n465_), .A4(new_n222_), .ZN(new_n4707_));
  NOR3_X1    g4652(.A1(new_n4706_), .A2(new_n399_), .A3(new_n4707_), .ZN(new_n4708_));
  NAND3_X1   g4653(.A1(new_n650_), .A2(new_n228_), .A3(new_n232_), .ZN(new_n4709_));
  NOR3_X1    g4654(.A1(new_n4709_), .A2(new_n217_), .A3(new_n625_), .ZN(new_n4710_));
  NOR4_X1    g4655(.A1(new_n658_), .A2(new_n317_), .A3(new_n519_), .A4(new_n635_), .ZN(new_n4711_));
  NAND3_X1   g4656(.A1(new_n4708_), .A2(new_n4710_), .A3(new_n4711_), .ZN(new_n4712_));
  NOR3_X1    g4657(.A1(new_n4712_), .A2(new_n633_), .A3(new_n4032_), .ZN(new_n4713_));
  INV_X1     g4658(.I(new_n4713_), .ZN(new_n4714_));
  AOI21_X1   g4659(.A1(new_n4698_), .A2(new_n4705_), .B(new_n4714_), .ZN(new_n4715_));
  NAND2_X1   g4660(.A1(new_n4715_), .A2(new_n4457_), .ZN(new_n4716_));
  NAND2_X1   g4661(.A1(new_n4426_), .A2(new_n4427_), .ZN(new_n4717_));
  AOI21_X1   g4662(.A1(new_n4424_), .A2(new_n4717_), .B(new_n4368_), .ZN(new_n4718_));
  NOR2_X1    g4663(.A1(new_n4424_), .A2(new_n4717_), .ZN(new_n4719_));
  NOR3_X1    g4664(.A1(new_n4211_), .A2(new_n4718_), .A3(new_n4719_), .ZN(new_n4720_));
  NAND3_X1   g4665(.A1(new_n4701_), .A2(new_n4416_), .A3(new_n4418_), .ZN(new_n4721_));
  OAI21_X1   g4666(.A1(new_n4695_), .A2(new_n4694_), .B(new_n4696_), .ZN(new_n4722_));
  NAND3_X1   g4667(.A1(new_n4680_), .A2(new_n4686_), .A3(new_n4692_), .ZN(new_n4723_));
  AOI22_X1   g4668(.A1(new_n4722_), .A2(new_n4723_), .B1(new_n4721_), .B2(new_n4492_), .ZN(new_n4724_));
  NAND3_X1   g4669(.A1(new_n4680_), .A2(new_n4686_), .A3(new_n4696_), .ZN(new_n4725_));
  OAI21_X1   g4670(.A1(new_n4695_), .A2(new_n4694_), .B(new_n4692_), .ZN(new_n4726_));
  AOI21_X1   g4671(.A1(new_n4725_), .A2(new_n4726_), .B(new_n4584_), .ZN(new_n4727_));
  NOR2_X1    g4672(.A1(new_n4727_), .A2(new_n4724_), .ZN(new_n4728_));
  OAI21_X1   g4673(.A1(new_n4728_), .A2(new_n4714_), .B(new_n4720_), .ZN(new_n4729_));
  AOI21_X1   g4674(.A1(new_n4729_), .A2(new_n4716_), .B(new_n4451_), .ZN(new_n4730_));
  INV_X1     g4675(.I(new_n4451_), .ZN(new_n4731_));
  NOR3_X1    g4676(.A1(new_n4720_), .A2(new_n4728_), .A3(new_n4714_), .ZN(new_n4732_));
  NOR2_X1    g4677(.A1(new_n4715_), .A2(new_n4457_), .ZN(new_n4733_));
  NOR3_X1    g4678(.A1(new_n4732_), .A2(new_n4733_), .A3(new_n4731_), .ZN(new_n4734_));
  NOR2_X1    g4679(.A1(new_n4730_), .A2(new_n4734_), .ZN(new_n4735_));
  INV_X1     g4680(.I(new_n4735_), .ZN(new_n4736_));
  NAND2_X1   g4681(.A1(new_n4736_), .A2(new_n4442_), .ZN(new_n4737_));
  XOR2_X1    g4682(.A1(new_n4449_), .A2(new_n4737_), .Z(new_n4738_));
  XOR2_X1    g4683(.A1(new_n4738_), .A2(new_n4445_), .Z(\sin[2] ));
  NAND2_X1   g4684(.A1(new_n4698_), .A2(new_n4705_), .ZN(new_n4740_));
  NAND2_X1   g4685(.A1(new_n4720_), .A2(new_n4740_), .ZN(new_n4741_));
  NAND2_X1   g4686(.A1(new_n4451_), .A2(new_n4713_), .ZN(new_n4742_));
  INV_X1     g4687(.I(new_n4742_), .ZN(new_n4743_));
  OAI21_X1   g4688(.A1(new_n4720_), .A2(new_n4740_), .B(new_n4743_), .ZN(new_n4744_));
  NAND2_X1   g4689(.A1(new_n4744_), .A2(new_n4741_), .ZN(new_n4745_));
  NOR2_X1    g4690(.A1(new_n4703_), .A2(new_n4704_), .ZN(new_n4746_));
  AOI21_X1   g4691(.A1(new_n4479_), .A2(new_n4230_), .B(new_n4474_), .ZN(new_n4747_));
  AOI21_X1   g4692(.A1(new_n4747_), .A2(new_n2947_), .B(new_n4486_), .ZN(new_n4748_));
  AOI21_X1   g4693(.A1(new_n4646_), .A2(new_n4510_), .B(new_n4598_), .ZN(new_n4749_));
  OAI21_X1   g4694(.A1(new_n4646_), .A2(new_n4510_), .B(new_n4596_), .ZN(new_n4750_));
  OAI21_X1   g4695(.A1(new_n3182_), .A2(new_n2994_), .B(new_n4608_), .ZN(new_n4751_));
  NAND2_X1   g4696(.A1(new_n2931_), .A2(new_n2998_), .ZN(new_n4752_));
  NAND2_X1   g4697(.A1(new_n4752_), .A2(new_n4751_), .ZN(new_n4753_));
  NAND2_X1   g4698(.A1(new_n4753_), .A2(new_n721_), .ZN(new_n4754_));
  NAND3_X1   g4699(.A1(new_n4754_), .A2(new_n3582_), .A3(new_n2992_), .ZN(new_n4755_));
  NAND2_X1   g4700(.A1(new_n4754_), .A2(new_n2992_), .ZN(new_n4756_));
  NAND2_X1   g4701(.A1(new_n4756_), .A2(new_n3571_), .ZN(new_n4757_));
  NAND2_X1   g4702(.A1(new_n2804_), .A2(new_n438_), .ZN(new_n4758_));
  XOR2_X1    g4703(.A1(new_n4625_), .A2(new_n4758_), .Z(new_n4759_));
  NOR2_X1    g4704(.A1(new_n4626_), .A2(new_n437_), .ZN(new_n4760_));
  OAI21_X1   g4705(.A1(new_n4621_), .A2(new_n4760_), .B(new_n4759_), .ZN(new_n4761_));
  NOR2_X1    g4706(.A1(new_n2734_), .A2(new_n3496_), .ZN(new_n4762_));
  INV_X1     g4707(.I(new_n4762_), .ZN(new_n4763_));
  NAND2_X1   g4708(.A1(new_n2720_), .A2(new_n3494_), .ZN(new_n4764_));
  AOI22_X1   g4709(.A1(new_n4764_), .A2(new_n4763_), .B1(new_n3189_), .B2(new_n4270_), .ZN(new_n4765_));
  INV_X1     g4710(.I(new_n4765_), .ZN(new_n4766_));
  AOI21_X1   g4711(.A1(new_n3235_), .A2(new_n3393_), .B(new_n4766_), .ZN(new_n4767_));
  NAND3_X1   g4712(.A1(new_n4761_), .A2(new_n437_), .A3(new_n4767_), .ZN(new_n4768_));
  INV_X1     g4713(.I(new_n4768_), .ZN(new_n4769_));
  AOI21_X1   g4714(.A1(new_n4761_), .A2(new_n4767_), .B(new_n437_), .ZN(new_n4770_));
  OAI21_X1   g4715(.A1(new_n4769_), .A2(new_n4770_), .B(new_n2956_), .ZN(new_n4771_));
  INV_X1     g4716(.I(new_n4770_), .ZN(new_n4772_));
  NAND3_X1   g4717(.A1(new_n4772_), .A2(new_n4768_), .A3(new_n2743_), .ZN(new_n4773_));
  AOI22_X1   g4718(.A1(new_n4773_), .A2(new_n4771_), .B1(new_n4755_), .B2(new_n4757_), .ZN(new_n4774_));
  OAI21_X1   g4719(.A1(new_n4749_), .A2(new_n4750_), .B(new_n4774_), .ZN(new_n4775_));
  NOR2_X1    g4720(.A1(new_n4749_), .A2(new_n4750_), .ZN(new_n4776_));
  NAND2_X1   g4721(.A1(new_n4757_), .A2(new_n4755_), .ZN(new_n4777_));
  AOI21_X1   g4722(.A1(new_n4772_), .A2(new_n4768_), .B(new_n2743_), .ZN(new_n4778_));
  NOR3_X1    g4723(.A1(new_n4769_), .A2(new_n4770_), .A3(new_n2956_), .ZN(new_n4779_));
  OAI21_X1   g4724(.A1(new_n4778_), .A2(new_n4779_), .B(new_n4777_), .ZN(new_n4780_));
  NAND2_X1   g4725(.A1(new_n4776_), .A2(new_n4780_), .ZN(new_n4781_));
  AOI21_X1   g4726(.A1(new_n4775_), .A2(new_n4781_), .B(new_n4641_), .ZN(new_n4782_));
  NOR2_X1    g4727(.A1(new_n4776_), .A2(new_n4780_), .ZN(new_n4783_));
  NOR3_X1    g4728(.A1(new_n4774_), .A2(new_n4749_), .A3(new_n4750_), .ZN(new_n4784_));
  NOR3_X1    g4729(.A1(new_n4784_), .A2(new_n4783_), .A3(new_n4645_), .ZN(new_n4785_));
  NAND2_X1   g4730(.A1(new_n3086_), .A2(new_n3076_), .ZN(new_n4786_));
  NAND2_X1   g4731(.A1(new_n2946_), .A2(new_n2898_), .ZN(new_n4787_));
  AOI22_X1   g4732(.A1(new_n4787_), .A2(new_n4786_), .B1(new_n2977_), .B2(new_n3597_), .ZN(new_n4788_));
  OAI21_X1   g4733(.A1(new_n4788_), .A2(new_n803_), .B(new_n2977_), .ZN(new_n4789_));
  XOR2_X1    g4734(.A1(new_n3607_), .A2(new_n4789_), .Z(new_n4790_));
  NOR3_X1    g4735(.A1(new_n4782_), .A2(new_n4785_), .A3(new_n4790_), .ZN(new_n4791_));
  OAI21_X1   g4736(.A1(new_n4784_), .A2(new_n4783_), .B(new_n4645_), .ZN(new_n4792_));
  NAND3_X1   g4737(.A1(new_n4775_), .A2(new_n4781_), .A3(new_n4641_), .ZN(new_n4793_));
  INV_X1     g4738(.I(new_n4790_), .ZN(new_n4794_));
  AOI21_X1   g4739(.A1(new_n4793_), .A2(new_n4792_), .B(new_n4794_), .ZN(new_n4795_));
  NOR2_X1    g4740(.A1(new_n4791_), .A2(new_n4795_), .ZN(new_n4796_));
  NAND2_X1   g4741(.A1(new_n4595_), .A2(new_n4587_), .ZN(new_n4797_));
  OAI21_X1   g4742(.A1(new_n4587_), .A2(new_n4595_), .B(new_n4653_), .ZN(new_n4798_));
  OAI21_X1   g4743(.A1(new_n4657_), .A2(new_n4798_), .B(new_n4797_), .ZN(new_n4799_));
  NAND2_X1   g4744(.A1(new_n4334_), .A2(new_n4333_), .ZN(new_n4800_));
  OAI22_X1   g4745(.A1(new_n4243_), .A2(new_n3282_), .B1(new_n4230_), .B2(new_n3237_), .ZN(new_n4801_));
  AOI21_X1   g4746(.A1(new_n4801_), .A2(new_n1050_), .B(new_n3207_), .ZN(new_n4802_));
  XOR2_X1    g4747(.A1(new_n4800_), .A2(new_n4802_), .Z(new_n4803_));
  NAND2_X1   g4748(.A1(new_n4799_), .A2(new_n4803_), .ZN(new_n4804_));
  AOI22_X1   g4749(.A1(new_n4588_), .A2(new_n4594_), .B1(new_n4650_), .B2(new_n4652_), .ZN(new_n4805_));
  NAND3_X1   g4750(.A1(new_n4590_), .A2(new_n4805_), .A3(new_n4314_), .ZN(new_n4806_));
  XNOR2_X1   g4751(.A1(new_n4800_), .A2(new_n4802_), .ZN(new_n4807_));
  NAND3_X1   g4752(.A1(new_n4806_), .A2(new_n4797_), .A3(new_n4807_), .ZN(new_n4808_));
  AOI21_X1   g4753(.A1(new_n4808_), .A2(new_n4804_), .B(new_n4796_), .ZN(new_n4809_));
  NAND3_X1   g4754(.A1(new_n4793_), .A2(new_n4792_), .A3(new_n4794_), .ZN(new_n4810_));
  OAI21_X1   g4755(.A1(new_n4782_), .A2(new_n4785_), .B(new_n4790_), .ZN(new_n4811_));
  NAND2_X1   g4756(.A1(new_n4811_), .A2(new_n4810_), .ZN(new_n4812_));
  NAND3_X1   g4757(.A1(new_n4806_), .A2(new_n4797_), .A3(new_n4803_), .ZN(new_n4813_));
  NAND2_X1   g4758(.A1(new_n4799_), .A2(new_n4807_), .ZN(new_n4814_));
  AOI21_X1   g4759(.A1(new_n4813_), .A2(new_n4814_), .B(new_n4812_), .ZN(new_n4815_));
  OAI21_X1   g4760(.A1(new_n4809_), .A2(new_n4815_), .B(new_n2943_), .ZN(new_n4816_));
  AOI21_X1   g4761(.A1(new_n4806_), .A2(new_n4797_), .B(new_n4807_), .ZN(new_n4817_));
  NOR2_X1    g4762(.A1(new_n4799_), .A2(new_n4803_), .ZN(new_n4818_));
  OAI21_X1   g4763(.A1(new_n4817_), .A2(new_n4818_), .B(new_n4812_), .ZN(new_n4819_));
  INV_X1     g4764(.I(new_n4797_), .ZN(new_n4820_));
  NAND2_X1   g4765(.A1(new_n4550_), .A2(new_n4553_), .ZN(new_n4821_));
  AOI21_X1   g4766(.A1(new_n4821_), .A2(new_n4326_), .B(new_n4312_), .ZN(new_n4822_));
  NOR3_X1    g4767(.A1(new_n4822_), .A2(new_n4328_), .A3(new_n4798_), .ZN(new_n4823_));
  NOR3_X1    g4768(.A1(new_n4823_), .A2(new_n4820_), .A3(new_n4807_), .ZN(new_n4824_));
  AOI21_X1   g4769(.A1(new_n4806_), .A2(new_n4797_), .B(new_n4803_), .ZN(new_n4825_));
  OAI21_X1   g4770(.A1(new_n4825_), .A2(new_n4824_), .B(new_n4796_), .ZN(new_n4826_));
  NAND3_X1   g4771(.A1(new_n4819_), .A2(new_n4826_), .A3(new_n2942_), .ZN(new_n4827_));
  AOI21_X1   g4772(.A1(new_n4816_), .A2(new_n4827_), .B(new_n4748_), .ZN(new_n4828_));
  INV_X1     g4773(.I(new_n4748_), .ZN(new_n4829_));
  NAND3_X1   g4774(.A1(new_n4819_), .A2(new_n4826_), .A3(new_n2943_), .ZN(new_n4830_));
  OAI21_X1   g4775(.A1(new_n4809_), .A2(new_n4815_), .B(new_n2942_), .ZN(new_n4831_));
  AOI21_X1   g4776(.A1(new_n4831_), .A2(new_n4830_), .B(new_n4829_), .ZN(new_n4832_));
  INV_X1     g4777(.I(new_n4672_), .ZN(new_n4833_));
  AOI21_X1   g4778(.A1(new_n4679_), .A2(new_n4668_), .B(new_n4833_), .ZN(new_n4834_));
  NOR3_X1    g4779(.A1(new_n4828_), .A2(new_n4832_), .A3(new_n4834_), .ZN(new_n4835_));
  AOI21_X1   g4780(.A1(new_n4819_), .A2(new_n4826_), .B(new_n2942_), .ZN(new_n4836_));
  NOR3_X1    g4781(.A1(new_n4809_), .A2(new_n4815_), .A3(new_n2943_), .ZN(new_n4837_));
  OAI21_X1   g4782(.A1(new_n4836_), .A2(new_n4837_), .B(new_n4829_), .ZN(new_n4838_));
  NOR3_X1    g4783(.A1(new_n4809_), .A2(new_n4815_), .A3(new_n2942_), .ZN(new_n4839_));
  AOI21_X1   g4784(.A1(new_n4819_), .A2(new_n4826_), .B(new_n2943_), .ZN(new_n4840_));
  OAI21_X1   g4785(.A1(new_n4840_), .A2(new_n4839_), .B(new_n4748_), .ZN(new_n4841_));
  OAI21_X1   g4786(.A1(new_n4685_), .A2(new_n4673_), .B(new_n4672_), .ZN(new_n4842_));
  AOI21_X1   g4787(.A1(new_n4838_), .A2(new_n4841_), .B(new_n4842_), .ZN(new_n4843_));
  NOR2_X1    g4788(.A1(new_n4843_), .A2(new_n4835_), .ZN(new_n4844_));
  NOR3_X1    g4789(.A1(new_n4746_), .A2(new_n4844_), .A3(new_n4693_), .ZN(new_n4845_));
  NOR2_X1    g4790(.A1(new_n4695_), .A2(new_n4694_), .ZN(new_n4846_));
  NOR2_X1    g4791(.A1(new_n4846_), .A2(new_n4692_), .ZN(new_n4848_));
  OAI21_X1   g4792(.A1(new_n4845_), .A2(new_n4848_), .B(new_n4702_), .ZN(new_n4849_));
  NAND2_X1   g4793(.A1(new_n4726_), .A2(new_n4725_), .ZN(new_n4850_));
  NAND3_X1   g4794(.A1(new_n4838_), .A2(new_n4841_), .A3(new_n4842_), .ZN(new_n4851_));
  OAI21_X1   g4795(.A1(new_n4828_), .A2(new_n4832_), .B(new_n4834_), .ZN(new_n4852_));
  NAND2_X1   g4796(.A1(new_n4851_), .A2(new_n4852_), .ZN(new_n4853_));
  NAND3_X1   g4797(.A1(new_n4850_), .A2(new_n4853_), .A3(new_n4722_), .ZN(new_n4854_));
  INV_X1     g4798(.I(new_n4848_), .ZN(new_n4855_));
  NAND3_X1   g4799(.A1(new_n4854_), .A2(new_n4584_), .A3(new_n4855_), .ZN(new_n4856_));
  NOR2_X1    g4800(.A1(new_n2220_), .A2(new_n591_), .ZN(new_n4857_));
  NAND4_X1   g4801(.A1(new_n234_), .A2(new_n2504_), .A3(new_n313_), .A4(new_n332_), .ZN(new_n4858_));
  NAND4_X1   g4802(.A1(new_n788_), .A2(new_n673_), .A3(new_n468_), .A4(new_n326_), .ZN(new_n4859_));
  NOR3_X1    g4803(.A1(new_n4044_), .A2(new_n4858_), .A3(new_n4859_), .ZN(new_n4860_));
  NAND4_X1   g4804(.A1(new_n4857_), .A2(new_n4860_), .A3(new_n1100_), .A4(new_n2650_), .ZN(new_n4861_));
  INV_X1     g4805(.I(new_n4861_), .ZN(new_n4862_));
  NAND3_X1   g4806(.A1(new_n4849_), .A2(new_n4856_), .A3(new_n4862_), .ZN(new_n4863_));
  AOI21_X1   g4807(.A1(new_n4854_), .A2(new_n4855_), .B(new_n4584_), .ZN(new_n4864_));
  NOR3_X1    g4808(.A1(new_n4845_), .A2(new_n4702_), .A3(new_n4848_), .ZN(new_n4865_));
  OAI21_X1   g4809(.A1(new_n4865_), .A2(new_n4864_), .B(new_n4861_), .ZN(new_n4866_));
  NAND2_X1   g4810(.A1(new_n4866_), .A2(new_n4863_), .ZN(new_n4867_));
  NAND3_X1   g4811(.A1(new_n4735_), .A2(new_n4745_), .A3(new_n4867_), .ZN(new_n4868_));
  NOR2_X1    g4812(.A1(new_n4457_), .A2(new_n4728_), .ZN(new_n4869_));
  AOI21_X1   g4813(.A1(new_n4457_), .A2(new_n4728_), .B(new_n4742_), .ZN(new_n4870_));
  NOR2_X1    g4814(.A1(new_n4870_), .A2(new_n4869_), .ZN(new_n4871_));
  NOR3_X1    g4815(.A1(new_n4865_), .A2(new_n4864_), .A3(new_n4861_), .ZN(new_n4872_));
  AOI21_X1   g4816(.A1(new_n4849_), .A2(new_n4856_), .B(new_n4862_), .ZN(new_n4873_));
  NOR2_X1    g4817(.A1(new_n4872_), .A2(new_n4873_), .ZN(new_n4874_));
  OAI22_X1   g4818(.A1(new_n4874_), .A2(new_n4871_), .B1(new_n4730_), .B2(new_n4734_), .ZN(new_n4875_));
  AOI21_X1   g4819(.A1(new_n4868_), .A2(new_n4875_), .B(new_n4442_), .ZN(new_n4876_));
  AND3_X2    g4820(.A1(new_n4868_), .A2(new_n4442_), .A3(new_n4875_), .Z(new_n4877_));
  NOR2_X1    g4821(.A1(new_n4877_), .A2(new_n4876_), .ZN(new_n4878_));
  NAND2_X1   g4822(.A1(new_n4736_), .A2(new_n4446_), .ZN(new_n4879_));
  NAND2_X1   g4823(.A1(new_n4735_), .A2(new_n4442_), .ZN(new_n4880_));
  NAND2_X1   g4824(.A1(new_n4879_), .A2(new_n4880_), .ZN(new_n4881_));
  NAND3_X1   g4825(.A1(new_n4881_), .A2(new_n4402_), .A3(new_n4448_), .ZN(new_n4882_));
  NAND2_X1   g4826(.A1(new_n4882_), .A2(new_n4404_), .ZN(new_n4883_));
  XNOR2_X1   g4827(.A1(new_n4883_), .A2(new_n4878_), .ZN(\sin[3] ));
  NAND2_X1   g4828(.A1(new_n4210_), .A2(new_n4076_), .ZN(new_n4885_));
  AOI22_X1   g4829(.A1(new_n4396_), .A2(new_n4885_), .B1(new_n4370_), .B2(new_n4371_), .ZN(new_n4886_));
  NOR2_X1    g4830(.A1(new_n4372_), .A2(new_n4398_), .ZN(new_n4887_));
  NOR2_X1    g4831(.A1(new_n4887_), .A2(new_n4886_), .ZN(new_n4888_));
  NOR2_X1    g4832(.A1(new_n4888_), .A2(new_n4391_), .ZN(new_n4889_));
  OAI21_X1   g4833(.A1(new_n4439_), .A2(new_n4432_), .B(new_n4211_), .ZN(new_n4890_));
  NAND3_X1   g4834(.A1(new_n4430_), .A2(new_n4398_), .A3(new_n4433_), .ZN(new_n4891_));
  NAND2_X1   g4835(.A1(new_n4890_), .A2(new_n4891_), .ZN(new_n4892_));
  NAND4_X1   g4836(.A1(new_n4889_), .A2(new_n4892_), .A3(new_n4866_), .A4(new_n4863_), .ZN(new_n4893_));
  OAI22_X1   g4837(.A1(new_n4408_), .A2(new_n4441_), .B1(new_n4872_), .B2(new_n4873_), .ZN(new_n4894_));
  OAI21_X1   g4838(.A1(new_n4730_), .A2(new_n4734_), .B(new_n4745_), .ZN(new_n4895_));
  AOI21_X1   g4839(.A1(new_n4893_), .A2(new_n4894_), .B(new_n4895_), .ZN(new_n4896_));
  INV_X1     g4840(.I(new_n4896_), .ZN(new_n4897_));
  OAI21_X1   g4841(.A1(new_n4828_), .A2(new_n4832_), .B(new_n4842_), .ZN(new_n4898_));
  OAI21_X1   g4842(.A1(new_n4843_), .A2(new_n4835_), .B(new_n4696_), .ZN(new_n4899_));
  NAND2_X1   g4843(.A1(new_n4899_), .A2(new_n4846_), .ZN(new_n4900_));
  AOI21_X1   g4844(.A1(new_n4844_), .A2(new_n4692_), .B(new_n4702_), .ZN(new_n4901_));
  XOR2_X1    g4845(.A1(new_n4748_), .A2(new_n2943_), .Z(new_n4902_));
  NAND2_X1   g4846(.A1(new_n4902_), .A2(new_n4803_), .ZN(new_n4903_));
  INV_X1     g4847(.I(new_n4903_), .ZN(new_n4904_));
  NOR2_X1    g4848(.A1(new_n4902_), .A2(new_n4803_), .ZN(new_n4905_));
  INV_X1     g4849(.I(new_n4799_), .ZN(new_n4906_));
  NAND2_X1   g4850(.A1(new_n4906_), .A2(new_n4812_), .ZN(new_n4907_));
  NAND2_X1   g4851(.A1(new_n4796_), .A2(new_n4799_), .ZN(new_n4908_));
  AOI21_X1   g4852(.A1(new_n4908_), .A2(new_n4907_), .B(new_n4905_), .ZN(new_n4909_));
  NAND2_X1   g4853(.A1(new_n4799_), .A2(new_n4811_), .ZN(new_n4910_));
  NAND2_X1   g4854(.A1(new_n4910_), .A2(new_n4810_), .ZN(new_n4911_));
  INV_X1     g4855(.I(new_n4911_), .ZN(new_n4912_));
  OAI22_X1   g4856(.A1(new_n4230_), .A2(new_n3211_), .B1(new_n3213_), .B2(new_n4182_), .ZN(new_n4913_));
  OAI21_X1   g4857(.A1(new_n3237_), .A2(new_n4474_), .B(new_n4913_), .ZN(new_n4914_));
  AOI21_X1   g4858(.A1(new_n4914_), .A2(new_n1050_), .B(new_n3207_), .ZN(new_n4915_));
  INV_X1     g4859(.I(new_n4915_), .ZN(new_n4916_));
  NOR3_X1    g4860(.A1(new_n4483_), .A2(new_n4478_), .A3(new_n4916_), .ZN(new_n4917_));
  NOR2_X1    g4861(.A1(new_n4484_), .A2(new_n4915_), .ZN(new_n4918_));
  NOR2_X1    g4862(.A1(new_n4918_), .A2(new_n4917_), .ZN(new_n4919_));
  NAND2_X1   g4863(.A1(new_n4777_), .A2(new_n4641_), .ZN(new_n4920_));
  INV_X1     g4864(.I(new_n4920_), .ZN(new_n4921_));
  NOR2_X1    g4865(.A1(new_n4778_), .A2(new_n4779_), .ZN(new_n4922_));
  NOR2_X1    g4866(.A1(new_n4777_), .A2(new_n4641_), .ZN(new_n4923_));
  NOR4_X1    g4867(.A1(new_n4922_), .A2(new_n4749_), .A3(new_n4750_), .A4(new_n4923_), .ZN(new_n4924_));
  NOR2_X1    g4868(.A1(new_n4924_), .A2(new_n4921_), .ZN(new_n4925_));
  NAND2_X1   g4869(.A1(new_n3436_), .A2(new_n2998_), .ZN(new_n4926_));
  NAND2_X1   g4870(.A1(new_n2898_), .A2(new_n3030_), .ZN(new_n4927_));
  AOI22_X1   g4871(.A1(new_n4927_), .A2(new_n4926_), .B1(new_n2931_), .B2(new_n3038_), .ZN(new_n4928_));
  OAI21_X1   g4872(.A1(new_n4928_), .A2(new_n702_), .B(new_n2992_), .ZN(new_n4929_));
  XOR2_X1    g4873(.A1(new_n3844_), .A2(new_n4929_), .Z(new_n4930_));
  INV_X1     g4874(.I(new_n4764_), .ZN(new_n4931_));
  NOR2_X1    g4875(.A1(new_n3189_), .A2(new_n3396_), .ZN(new_n4932_));
  OAI22_X1   g4876(.A1(new_n4931_), .A2(new_n4932_), .B1(new_n2701_), .B2(new_n3496_), .ZN(new_n4933_));
  AOI21_X1   g4877(.A1(new_n4933_), .A2(new_n437_), .B(new_n3501_), .ZN(new_n4934_));
  XNOR2_X1   g4878(.A1(new_n4934_), .A2(new_n3202_), .ZN(new_n4935_));
  NAND2_X1   g4879(.A1(new_n4935_), .A2(new_n2943_), .ZN(new_n4936_));
  NOR2_X1    g4880(.A1(new_n4936_), .A2(new_n2813_), .ZN(new_n4937_));
  NAND2_X1   g4881(.A1(new_n4936_), .A2(new_n2813_), .ZN(new_n4938_));
  INV_X1     g4882(.I(new_n4938_), .ZN(new_n4939_));
  OAI21_X1   g4883(.A1(new_n4939_), .A2(new_n4937_), .B(new_n437_), .ZN(new_n4940_));
  INV_X1     g4884(.I(new_n4937_), .ZN(new_n4941_));
  NAND3_X1   g4885(.A1(new_n4941_), .A2(new_n438_), .A3(new_n4938_), .ZN(new_n4942_));
  NAND3_X1   g4886(.A1(new_n4767_), .A2(new_n437_), .A3(new_n2743_), .ZN(new_n4943_));
  INV_X1     g4887(.I(new_n4761_), .ZN(new_n4944_));
  NOR2_X1    g4888(.A1(new_n2956_), .A2(new_n438_), .ZN(new_n4945_));
  INV_X1     g4889(.I(new_n4945_), .ZN(new_n4946_));
  XOR2_X1    g4890(.A1(new_n4767_), .A2(new_n4946_), .Z(new_n4947_));
  NAND2_X1   g4891(.A1(new_n4944_), .A2(new_n4947_), .ZN(new_n4948_));
  NAND2_X1   g4892(.A1(new_n4948_), .A2(new_n4943_), .ZN(new_n4949_));
  INV_X1     g4893(.I(new_n4949_), .ZN(new_n4950_));
  NAND3_X1   g4894(.A1(new_n4950_), .A2(new_n4940_), .A3(new_n4942_), .ZN(new_n4951_));
  AOI21_X1   g4895(.A1(new_n4941_), .A2(new_n4938_), .B(new_n438_), .ZN(new_n4952_));
  NOR3_X1    g4896(.A1(new_n4939_), .A2(new_n437_), .A3(new_n4937_), .ZN(new_n4953_));
  OAI21_X1   g4897(.A1(new_n4952_), .A2(new_n4953_), .B(new_n4949_), .ZN(new_n4954_));
  AOI21_X1   g4898(.A1(new_n4951_), .A2(new_n4954_), .B(new_n4930_), .ZN(new_n4955_));
  INV_X1     g4899(.I(new_n4955_), .ZN(new_n4956_));
  AOI21_X1   g4900(.A1(new_n4940_), .A2(new_n4942_), .B(new_n4949_), .ZN(new_n4957_));
  NOR3_X1    g4901(.A1(new_n4950_), .A2(new_n4952_), .A3(new_n4953_), .ZN(new_n4958_));
  OAI21_X1   g4902(.A1(new_n4958_), .A2(new_n4957_), .B(new_n4930_), .ZN(new_n4959_));
  OAI22_X1   g4903(.A1(new_n2926_), .A2(new_n2972_), .B1(new_n3597_), .B2(new_n2975_), .ZN(new_n4960_));
  OAI21_X1   g4904(.A1(new_n3987_), .A2(new_n2969_), .B(new_n4960_), .ZN(new_n4961_));
  AOI21_X1   g4905(.A1(new_n4961_), .A2(new_n802_), .B(new_n2969_), .ZN(new_n4962_));
  XOR2_X1    g4906(.A1(new_n3982_), .A2(new_n4962_), .Z(new_n4963_));
  NAND3_X1   g4907(.A1(new_n4956_), .A2(new_n4959_), .A3(new_n4963_), .ZN(new_n4964_));
  INV_X1     g4908(.I(new_n4959_), .ZN(new_n4965_));
  XNOR2_X1   g4909(.A1(new_n3982_), .A2(new_n4962_), .ZN(new_n4966_));
  OAI21_X1   g4910(.A1(new_n4965_), .A2(new_n4955_), .B(new_n4966_), .ZN(new_n4967_));
  AOI21_X1   g4911(.A1(new_n4967_), .A2(new_n4964_), .B(new_n4925_), .ZN(new_n4968_));
  AOI21_X1   g4912(.A1(new_n4956_), .A2(new_n4959_), .B(new_n4966_), .ZN(new_n4969_));
  NOR3_X1    g4913(.A1(new_n4965_), .A2(new_n4963_), .A3(new_n4955_), .ZN(new_n4970_));
  OAI21_X1   g4914(.A1(new_n4969_), .A2(new_n4970_), .B(new_n4925_), .ZN(new_n4971_));
  INV_X1     g4915(.I(new_n4971_), .ZN(new_n4972_));
  OAI21_X1   g4916(.A1(new_n4972_), .A2(new_n4968_), .B(new_n4919_), .ZN(new_n4973_));
  INV_X1     g4917(.I(new_n4919_), .ZN(new_n4974_));
  INV_X1     g4918(.I(new_n4968_), .ZN(new_n4975_));
  NAND3_X1   g4919(.A1(new_n4974_), .A2(new_n4975_), .A3(new_n4971_), .ZN(new_n4976_));
  AOI21_X1   g4920(.A1(new_n4973_), .A2(new_n4976_), .B(new_n4912_), .ZN(new_n4977_));
  AOI21_X1   g4921(.A1(new_n4975_), .A2(new_n4971_), .B(new_n4919_), .ZN(new_n4978_));
  INV_X1     g4922(.I(new_n4978_), .ZN(new_n4979_));
  NOR3_X1    g4923(.A1(new_n4974_), .A2(new_n4972_), .A3(new_n4968_), .ZN(new_n4980_));
  INV_X1     g4924(.I(new_n4980_), .ZN(new_n4981_));
  AOI21_X1   g4925(.A1(new_n4981_), .A2(new_n4979_), .B(new_n4911_), .ZN(new_n4982_));
  NOR4_X1    g4926(.A1(new_n4982_), .A2(new_n4904_), .A3(new_n4977_), .A4(new_n4909_), .ZN(new_n4983_));
  NAND2_X1   g4927(.A1(new_n4907_), .A2(new_n4908_), .ZN(new_n4984_));
  OAI21_X1   g4928(.A1(new_n4803_), .A2(new_n4902_), .B(new_n4984_), .ZN(new_n4985_));
  NAND2_X1   g4929(.A1(new_n4976_), .A2(new_n4973_), .ZN(new_n4986_));
  NAND2_X1   g4930(.A1(new_n4986_), .A2(new_n4911_), .ZN(new_n4987_));
  OAI21_X1   g4931(.A1(new_n4978_), .A2(new_n4980_), .B(new_n4912_), .ZN(new_n4988_));
  AOI22_X1   g4932(.A1(new_n4987_), .A2(new_n4988_), .B1(new_n4985_), .B2(new_n4903_), .ZN(new_n4989_));
  NOR2_X1    g4933(.A1(new_n753_), .A2(new_n749_), .ZN(new_n4990_));
  NAND4_X1   g4934(.A1(new_n526_), .A2(new_n251_), .A3(new_n366_), .A4(new_n892_), .ZN(new_n4991_));
  NAND2_X1   g4935(.A1(new_n2852_), .A2(new_n2437_), .ZN(new_n4992_));
  NOR4_X1    g4936(.A1(new_n4992_), .A2(new_n4991_), .A3(new_n2574_), .A4(new_n312_), .ZN(new_n4993_));
  NAND4_X1   g4937(.A1(new_n2410_), .A2(new_n613_), .A3(new_n4990_), .A4(new_n4993_), .ZN(new_n4994_));
  INV_X1     g4938(.I(new_n4994_), .ZN(new_n4995_));
  OAI21_X1   g4939(.A1(new_n4989_), .A2(new_n4983_), .B(new_n4995_), .ZN(new_n4996_));
  AOI21_X1   g4940(.A1(new_n4901_), .A2(new_n4900_), .B(new_n4996_), .ZN(new_n4997_));
  INV_X1     g4941(.I(new_n4846_), .ZN(new_n4998_));
  AOI21_X1   g4942(.A1(new_n4853_), .A2(new_n4696_), .B(new_n4998_), .ZN(new_n4999_));
  OAI21_X1   g4943(.A1(new_n4853_), .A2(new_n4696_), .B(new_n4584_), .ZN(new_n5000_));
  INV_X1     g4944(.I(new_n4996_), .ZN(new_n5001_));
  NOR3_X1    g4945(.A1(new_n4999_), .A2(new_n5000_), .A3(new_n5001_), .ZN(new_n5002_));
  OAI21_X1   g4946(.A1(new_n4997_), .A2(new_n5002_), .B(new_n4898_), .ZN(new_n5003_));
  INV_X1     g4947(.I(new_n4898_), .ZN(new_n5004_));
  OAI21_X1   g4948(.A1(new_n4999_), .A2(new_n5000_), .B(new_n5001_), .ZN(new_n5005_));
  NAND3_X1   g4949(.A1(new_n4901_), .A2(new_n4900_), .A3(new_n4996_), .ZN(new_n5006_));
  NAND3_X1   g4950(.A1(new_n5005_), .A2(new_n5006_), .A3(new_n5004_), .ZN(new_n5007_));
  NAND3_X1   g4951(.A1(new_n4866_), .A2(new_n5003_), .A3(new_n5007_), .ZN(new_n5008_));
  NAND3_X1   g4952(.A1(new_n5008_), .A2(new_n4867_), .A3(new_n4871_), .ZN(new_n5009_));
  AOI21_X1   g4953(.A1(new_n5005_), .A2(new_n5006_), .B(new_n5004_), .ZN(new_n5010_));
  NOR3_X1    g4954(.A1(new_n4997_), .A2(new_n5002_), .A3(new_n4898_), .ZN(new_n5011_));
  NOR3_X1    g4955(.A1(new_n5010_), .A2(new_n5011_), .A3(new_n4873_), .ZN(new_n5012_));
  OAI21_X1   g4956(.A1(new_n5012_), .A2(new_n4874_), .B(new_n4745_), .ZN(new_n5013_));
  NAND2_X1   g4957(.A1(new_n5013_), .A2(new_n5009_), .ZN(new_n5014_));
  NAND2_X1   g4958(.A1(new_n4897_), .A2(new_n5014_), .ZN(new_n5015_));
  NAND3_X1   g4959(.A1(new_n4896_), .A2(new_n5009_), .A3(new_n5013_), .ZN(new_n5016_));
  NAND2_X1   g4960(.A1(new_n5015_), .A2(new_n5016_), .ZN(new_n5017_));
  NOR2_X1    g4961(.A1(new_n4878_), .A2(new_n4882_), .ZN(new_n5018_));
  NOR2_X1    g4962(.A1(new_n5018_), .A2(new_n4445_), .ZN(new_n5019_));
  XOR2_X1    g4963(.A1(new_n5019_), .A2(new_n5017_), .Z(\sin[4] ));
  NOR3_X1    g4964(.A1(new_n5017_), .A2(new_n4878_), .A3(new_n4882_), .ZN(new_n5021_));
  NAND2_X1   g4965(.A1(new_n4894_), .A2(new_n4893_), .ZN(new_n5022_));
  NAND2_X1   g4966(.A1(new_n5008_), .A2(new_n4867_), .ZN(new_n5023_));
  NAND4_X1   g4967(.A1(new_n5022_), .A2(new_n4736_), .A3(new_n5023_), .A4(new_n4745_), .ZN(new_n5024_));
  NOR2_X1    g4968(.A1(new_n4898_), .A2(new_n4983_), .ZN(new_n5025_));
  INV_X1     g4969(.I(new_n5025_), .ZN(new_n5026_));
  NOR3_X1    g4970(.A1(new_n4999_), .A2(new_n5000_), .A3(new_n5026_), .ZN(new_n5027_));
  NOR2_X1    g4971(.A1(new_n5027_), .A2(new_n4989_), .ZN(new_n5028_));
  AOI21_X1   g4972(.A1(new_n4979_), .A2(new_n4911_), .B(new_n4980_), .ZN(new_n5029_));
  NOR2_X1    g4973(.A1(new_n4474_), .A2(new_n3211_), .ZN(new_n5030_));
  OAI21_X1   g4974(.A1(new_n4230_), .A2(new_n3213_), .B(new_n1050_), .ZN(new_n5031_));
  OAI21_X1   g4975(.A1(new_n5030_), .A2(new_n5031_), .B(new_n3280_), .ZN(new_n5032_));
  XOR2_X1    g4976(.A1(new_n4688_), .A2(new_n5032_), .Z(new_n5033_));
  NOR2_X1    g4977(.A1(new_n4970_), .A2(new_n4925_), .ZN(new_n5034_));
  NOR2_X1    g4978(.A1(new_n5034_), .A2(new_n4969_), .ZN(new_n5035_));
  INV_X1     g4979(.I(new_n4958_), .ZN(new_n5036_));
  AOI21_X1   g4980(.A1(new_n5036_), .A2(new_n4930_), .B(new_n4957_), .ZN(new_n5037_));
  OAI21_X1   g4981(.A1(new_n4191_), .A2(new_n4197_), .B(new_n2977_), .ZN(new_n5038_));
  NOR2_X1    g4982(.A1(new_n3597_), .A2(new_n2972_), .ZN(new_n5039_));
  NOR2_X1    g4983(.A1(new_n3987_), .A2(new_n2975_), .ZN(new_n5040_));
  OAI22_X1   g4984(.A1(new_n5039_), .A2(new_n5040_), .B1(new_n4192_), .B2(new_n2969_), .ZN(new_n5041_));
  INV_X1     g4985(.I(new_n5041_), .ZN(new_n5042_));
  NAND2_X1   g4986(.A1(new_n5038_), .A2(new_n5042_), .ZN(new_n5043_));
  INV_X1     g4987(.I(new_n5043_), .ZN(new_n5044_));
  NOR2_X1    g4988(.A1(new_n2729_), .A2(new_n438_), .ZN(new_n5045_));
  INV_X1     g4989(.I(new_n5045_), .ZN(new_n5046_));
  NOR2_X1    g4990(.A1(new_n438_), .A2(new_n2943_), .ZN(new_n5047_));
  AOI22_X1   g4991(.A1(new_n5046_), .A2(new_n2943_), .B1(new_n3189_), .B2(new_n5047_), .ZN(new_n5048_));
  NOR2_X1    g4992(.A1(new_n2734_), .A2(new_n437_), .ZN(new_n5049_));
  OAI21_X1   g4993(.A1(new_n4935_), .A2(new_n2943_), .B(new_n5049_), .ZN(new_n5050_));
  NAND2_X1   g4994(.A1(new_n5050_), .A2(new_n4936_), .ZN(new_n5051_));
  OAI22_X1   g4995(.A1(new_n2902_), .A2(new_n3031_), .B1(new_n2931_), .B2(new_n2994_), .ZN(new_n5052_));
  OAI21_X1   g4996(.A1(new_n2926_), .A2(new_n3028_), .B(new_n5052_), .ZN(new_n5053_));
  AOI21_X1   g4997(.A1(new_n5053_), .A2(new_n721_), .B(new_n2991_), .ZN(new_n5054_));
  NAND3_X1   g4998(.A1(new_n2934_), .A2(new_n2928_), .A3(new_n5054_), .ZN(new_n5055_));
  AOI21_X1   g4999(.A1(new_n2934_), .A2(new_n2928_), .B(new_n5054_), .ZN(new_n5056_));
  INV_X1     g5000(.I(new_n5056_), .ZN(new_n5057_));
  NAND2_X1   g5001(.A1(new_n2720_), .A2(new_n3398_), .ZN(new_n5058_));
  NAND2_X1   g5002(.A1(new_n3436_), .A2(new_n3494_), .ZN(new_n5059_));
  AOI22_X1   g5003(.A1(new_n5059_), .A2(new_n5058_), .B1(new_n3182_), .B2(new_n4270_), .ZN(new_n5060_));
  OAI21_X1   g5004(.A1(new_n5060_), .A2(new_n438_), .B(new_n3393_), .ZN(new_n5061_));
  XOR2_X1    g5005(.A1(new_n3464_), .A2(new_n5061_), .Z(new_n5062_));
  INV_X1     g5006(.I(new_n5062_), .ZN(new_n5063_));
  NAND3_X1   g5007(.A1(new_n5057_), .A2(new_n5055_), .A3(new_n5063_), .ZN(new_n5064_));
  INV_X1     g5008(.I(new_n5055_), .ZN(new_n5065_));
  OAI21_X1   g5009(.A1(new_n5065_), .A2(new_n5056_), .B(new_n5062_), .ZN(new_n5066_));
  AOI21_X1   g5010(.A1(new_n5064_), .A2(new_n5066_), .B(new_n5051_), .ZN(new_n5067_));
  INV_X1     g5011(.I(new_n5051_), .ZN(new_n5068_));
  NOR3_X1    g5012(.A1(new_n5065_), .A2(new_n5056_), .A3(new_n5062_), .ZN(new_n5069_));
  AOI21_X1   g5013(.A1(new_n5057_), .A2(new_n5055_), .B(new_n5063_), .ZN(new_n5070_));
  NOR3_X1    g5014(.A1(new_n5070_), .A2(new_n5069_), .A3(new_n5068_), .ZN(new_n5071_));
  OAI21_X1   g5015(.A1(new_n5067_), .A2(new_n5071_), .B(new_n5048_), .ZN(new_n5072_));
  INV_X1     g5016(.I(new_n5048_), .ZN(new_n5073_));
  OAI21_X1   g5017(.A1(new_n5070_), .A2(new_n5069_), .B(new_n5068_), .ZN(new_n5074_));
  NAND3_X1   g5018(.A1(new_n5064_), .A2(new_n5066_), .A3(new_n5051_), .ZN(new_n5075_));
  NAND3_X1   g5019(.A1(new_n5074_), .A2(new_n5075_), .A3(new_n5073_), .ZN(new_n5076_));
  AOI21_X1   g5020(.A1(new_n5072_), .A2(new_n5076_), .B(new_n5044_), .ZN(new_n5077_));
  AOI21_X1   g5021(.A1(new_n5074_), .A2(new_n5075_), .B(new_n5073_), .ZN(new_n5078_));
  NOR3_X1    g5022(.A1(new_n5067_), .A2(new_n5071_), .A3(new_n5048_), .ZN(new_n5079_));
  NOR3_X1    g5023(.A1(new_n5079_), .A2(new_n5078_), .A3(new_n5043_), .ZN(new_n5080_));
  OAI21_X1   g5024(.A1(new_n5077_), .A2(new_n5080_), .B(new_n5037_), .ZN(new_n5081_));
  INV_X1     g5025(.I(new_n5037_), .ZN(new_n5082_));
  OAI21_X1   g5026(.A1(new_n5079_), .A2(new_n5078_), .B(new_n5043_), .ZN(new_n5083_));
  NAND3_X1   g5027(.A1(new_n5044_), .A2(new_n5072_), .A3(new_n5076_), .ZN(new_n5084_));
  NAND3_X1   g5028(.A1(new_n5084_), .A2(new_n5083_), .A3(new_n5082_), .ZN(new_n5085_));
  AOI21_X1   g5029(.A1(new_n5081_), .A2(new_n5085_), .B(new_n803_), .ZN(new_n5086_));
  AOI21_X1   g5030(.A1(new_n5084_), .A2(new_n5083_), .B(new_n5082_), .ZN(new_n5087_));
  NOR3_X1    g5031(.A1(new_n5077_), .A2(new_n5080_), .A3(new_n5037_), .ZN(new_n5088_));
  NOR3_X1    g5032(.A1(new_n5088_), .A2(new_n5087_), .A3(new_n802_), .ZN(new_n5089_));
  OAI21_X1   g5033(.A1(new_n5089_), .A2(new_n5086_), .B(new_n5035_), .ZN(new_n5090_));
  INV_X1     g5034(.I(new_n5035_), .ZN(new_n5091_));
  OAI21_X1   g5035(.A1(new_n5088_), .A2(new_n5087_), .B(new_n802_), .ZN(new_n5092_));
  NAND3_X1   g5036(.A1(new_n5081_), .A2(new_n5085_), .A3(new_n803_), .ZN(new_n5093_));
  NAND3_X1   g5037(.A1(new_n5092_), .A2(new_n5093_), .A3(new_n5091_), .ZN(new_n5094_));
  AOI21_X1   g5038(.A1(new_n5090_), .A2(new_n5094_), .B(new_n5033_), .ZN(new_n5095_));
  INV_X1     g5039(.I(new_n5033_), .ZN(new_n5096_));
  OAI21_X1   g5040(.A1(new_n5089_), .A2(new_n5086_), .B(new_n5091_), .ZN(new_n5097_));
  NAND3_X1   g5041(.A1(new_n5092_), .A2(new_n5093_), .A3(new_n5035_), .ZN(new_n5098_));
  AOI21_X1   g5042(.A1(new_n5097_), .A2(new_n5098_), .B(new_n5096_), .ZN(new_n5099_));
  NOR2_X1    g5043(.A1(new_n5095_), .A2(new_n5099_), .ZN(new_n5100_));
  NAND2_X1   g5044(.A1(new_n5100_), .A2(new_n5029_), .ZN(new_n5101_));
  INV_X1     g5045(.I(new_n5029_), .ZN(new_n5102_));
  AOI21_X1   g5046(.A1(new_n5092_), .A2(new_n5093_), .B(new_n5091_), .ZN(new_n5103_));
  INV_X1     g5047(.I(new_n5094_), .ZN(new_n5104_));
  OAI21_X1   g5048(.A1(new_n5104_), .A2(new_n5103_), .B(new_n5096_), .ZN(new_n5105_));
  AOI21_X1   g5049(.A1(new_n5092_), .A2(new_n5093_), .B(new_n5035_), .ZN(new_n5106_));
  NOR3_X1    g5050(.A1(new_n5089_), .A2(new_n5086_), .A3(new_n5091_), .ZN(new_n5107_));
  OAI21_X1   g5051(.A1(new_n5107_), .A2(new_n5106_), .B(new_n5033_), .ZN(new_n5108_));
  NAND2_X1   g5052(.A1(new_n5105_), .A2(new_n5108_), .ZN(new_n5109_));
  NAND2_X1   g5053(.A1(new_n5109_), .A2(new_n5102_), .ZN(new_n5110_));
  NAND2_X1   g5054(.A1(new_n5110_), .A2(new_n5101_), .ZN(new_n5111_));
  NOR4_X1    g5055(.A1(new_n636_), .A2(new_n151_), .A3(new_n191_), .A4(new_n251_), .ZN(new_n5112_));
  NOR3_X1    g5056(.A1(new_n110_), .A2(new_n468_), .A3(new_n375_), .ZN(new_n5113_));
  AND3_X2    g5057(.A1(new_n5112_), .A2(new_n2274_), .A3(new_n5113_), .Z(new_n5114_));
  NOR4_X1    g5058(.A1(new_n207_), .A2(new_n187_), .A3(new_n390_), .A4(new_n675_), .ZN(new_n5115_));
  INV_X1     g5059(.I(new_n5115_), .ZN(new_n5116_));
  NOR2_X1    g5060(.A1(new_n401_), .A2(new_n156_), .ZN(new_n5117_));
  NAND2_X1   g5061(.A1(new_n5117_), .A2(new_n1240_), .ZN(new_n5118_));
  NOR4_X1    g5062(.A1(new_n5116_), .A2(new_n2284_), .A3(new_n350_), .A4(new_n5118_), .ZN(new_n5119_));
  NAND4_X1   g5063(.A1(new_n2915_), .A2(new_n4466_), .A3(new_n5114_), .A4(new_n5119_), .ZN(new_n5120_));
  INV_X1     g5064(.I(new_n5120_), .ZN(new_n5121_));
  NAND2_X1   g5065(.A1(new_n5111_), .A2(new_n5121_), .ZN(new_n5122_));
  INV_X1     g5066(.I(new_n5101_), .ZN(new_n5123_));
  NOR2_X1    g5067(.A1(new_n5100_), .A2(new_n5029_), .ZN(new_n5124_));
  NOR2_X1    g5068(.A1(new_n5123_), .A2(new_n5124_), .ZN(new_n5125_));
  NAND2_X1   g5069(.A1(new_n5125_), .A2(new_n5120_), .ZN(new_n5126_));
  AND2_X2    g5070(.A1(new_n5126_), .A2(new_n5122_), .Z(new_n5127_));
  INV_X1     g5071(.I(new_n4989_), .ZN(new_n5128_));
  NAND3_X1   g5072(.A1(new_n4901_), .A2(new_n4900_), .A3(new_n5025_), .ZN(new_n5129_));
  NAND3_X1   g5073(.A1(new_n5110_), .A2(new_n5101_), .A3(new_n5121_), .ZN(new_n5130_));
  AOI21_X1   g5074(.A1(new_n5110_), .A2(new_n5101_), .B(new_n5121_), .ZN(new_n5131_));
  INV_X1     g5075(.I(new_n5131_), .ZN(new_n5132_));
  NAND2_X1   g5076(.A1(new_n5132_), .A2(new_n5130_), .ZN(new_n5133_));
  NAND3_X1   g5077(.A1(new_n5133_), .A2(new_n5129_), .A3(new_n5128_), .ZN(new_n5134_));
  OAI21_X1   g5078(.A1(new_n5028_), .A2(new_n5127_), .B(new_n5134_), .ZN(new_n5135_));
  OAI21_X1   g5079(.A1(new_n4872_), .A2(new_n4873_), .B(new_n4745_), .ZN(new_n5137_));
  XOR2_X1    g5080(.A1(new_n4996_), .A2(new_n4898_), .Z(new_n5138_));
  NAND3_X1   g5081(.A1(new_n5138_), .A2(new_n4900_), .A3(new_n4901_), .ZN(new_n5139_));
  AOI21_X1   g5082(.A1(new_n5137_), .A2(new_n5139_), .B(new_n5135_), .ZN(new_n5140_));
  AOI21_X1   g5083(.A1(new_n4863_), .A2(new_n4866_), .B(new_n4871_), .ZN(new_n5141_));
  AOI22_X1   g5084(.A1(new_n5129_), .A2(new_n5128_), .B1(new_n5122_), .B2(new_n5126_), .ZN(new_n5142_));
  INV_X1     g5085(.I(new_n5130_), .ZN(new_n5143_));
  NOR2_X1    g5086(.A1(new_n5143_), .A2(new_n5131_), .ZN(new_n5144_));
  NOR3_X1    g5087(.A1(new_n5144_), .A2(new_n5027_), .A3(new_n4989_), .ZN(new_n5145_));
  OAI21_X1   g5088(.A1(new_n5145_), .A2(new_n5142_), .B(new_n5139_), .ZN(new_n5146_));
  NOR2_X1    g5089(.A1(new_n5141_), .A2(new_n5146_), .ZN(new_n5147_));
  NOR2_X1    g5090(.A1(new_n5140_), .A2(new_n5147_), .ZN(new_n5148_));
  NOR2_X1    g5091(.A1(new_n5024_), .A2(new_n5148_), .ZN(new_n5149_));
  XOR2_X1    g5092(.A1(new_n5021_), .A2(new_n5149_), .Z(new_n5150_));
  XOR2_X1    g5093(.A1(new_n5150_), .A2(new_n4445_), .Z(\sin[5] ));
  INV_X1     g5094(.I(new_n5149_), .ZN(new_n5152_));
  NAND3_X1   g5095(.A1(new_n5129_), .A2(new_n5128_), .A3(new_n5125_), .ZN(new_n5153_));
  INV_X1     g5096(.I(new_n5153_), .ZN(new_n5154_));
  NOR2_X1    g5097(.A1(new_n5028_), .A2(new_n5125_), .ZN(new_n5155_));
  NOR2_X1    g5098(.A1(new_n5155_), .A2(new_n5154_), .ZN(new_n5156_));
  NOR2_X1    g5099(.A1(new_n5156_), .A2(new_n5137_), .ZN(new_n5157_));
  NOR2_X1    g5100(.A1(new_n5139_), .A2(new_n5120_), .ZN(new_n5158_));
  INV_X1     g5101(.I(new_n5158_), .ZN(new_n5159_));
  AOI21_X1   g5102(.A1(new_n5156_), .A2(new_n5137_), .B(new_n5159_), .ZN(new_n5160_));
  NOR2_X1    g5103(.A1(new_n5160_), .A2(new_n5157_), .ZN(new_n5161_));
  OAI21_X1   g5104(.A1(new_n5096_), .A2(new_n5103_), .B(new_n5094_), .ZN(new_n5162_));
  INV_X1     g5105(.I(new_n5162_), .ZN(new_n5163_));
  OAI22_X1   g5106(.A1(new_n4182_), .A2(new_n2975_), .B1(new_n3987_), .B2(new_n2972_), .ZN(new_n5164_));
  OAI21_X1   g5107(.A1(new_n2969_), .A2(new_n4230_), .B(new_n5164_), .ZN(new_n5165_));
  AOI21_X1   g5108(.A1(new_n5165_), .A2(new_n802_), .B(new_n2969_), .ZN(new_n5166_));
  XNOR2_X1   g5109(.A1(new_n4800_), .A2(new_n5166_), .ZN(new_n5167_));
  NAND2_X1   g5110(.A1(new_n2946_), .A2(new_n3030_), .ZN(new_n5168_));
  AOI22_X1   g5111(.A1(new_n2898_), .A2(new_n3038_), .B1(new_n3597_), .B2(new_n2998_), .ZN(new_n5169_));
  AOI21_X1   g5112(.A1(new_n5169_), .A2(new_n5168_), .B(new_n2991_), .ZN(new_n5170_));
  NAND2_X1   g5113(.A1(new_n3607_), .A2(new_n5170_), .ZN(new_n5171_));
  XOR2_X1    g5114(.A1(new_n5171_), .A2(new_n702_), .Z(new_n5172_));
  OAI21_X1   g5115(.A1(new_n4935_), .A2(new_n5049_), .B(new_n2943_), .ZN(new_n5173_));
  AOI21_X1   g5116(.A1(new_n4935_), .A2(new_n5049_), .B(new_n2943_), .ZN(new_n5174_));
  NOR2_X1    g5117(.A1(new_n3189_), .A2(new_n437_), .ZN(new_n5175_));
  INV_X1     g5118(.I(new_n5175_), .ZN(new_n5176_));
  OAI21_X1   g5119(.A1(new_n5174_), .A2(new_n5176_), .B(new_n5173_), .ZN(new_n5177_));
  NAND2_X1   g5120(.A1(new_n5177_), .A2(new_n2943_), .ZN(new_n5178_));
  NOR2_X1    g5121(.A1(new_n5178_), .A2(new_n438_), .ZN(new_n5179_));
  NAND2_X1   g5122(.A1(new_n5178_), .A2(new_n438_), .ZN(new_n5180_));
  INV_X1     g5123(.I(new_n5180_), .ZN(new_n5181_));
  OAI21_X1   g5124(.A1(new_n5181_), .A2(new_n5179_), .B(new_n3183_), .ZN(new_n5182_));
  INV_X1     g5125(.I(new_n5179_), .ZN(new_n5183_));
  NAND3_X1   g5126(.A1(new_n5183_), .A2(new_n2720_), .A3(new_n5180_), .ZN(new_n5184_));
  OAI21_X1   g5127(.A1(new_n3182_), .A2(new_n3396_), .B(new_n5059_), .ZN(new_n5185_));
  OAI21_X1   g5128(.A1(new_n2879_), .A2(new_n3496_), .B(new_n5185_), .ZN(new_n5186_));
  AOI21_X1   g5129(.A1(new_n5186_), .A2(new_n437_), .B(new_n3501_), .ZN(new_n5187_));
  XOR2_X1    g5130(.A1(new_n3582_), .A2(new_n5187_), .Z(new_n5188_));
  INV_X1     g5131(.I(new_n5188_), .ZN(new_n5189_));
  NAND3_X1   g5132(.A1(new_n5182_), .A2(new_n5184_), .A3(new_n5189_), .ZN(new_n5190_));
  AOI21_X1   g5133(.A1(new_n5182_), .A2(new_n5184_), .B(new_n5189_), .ZN(new_n5191_));
  INV_X1     g5134(.I(new_n5191_), .ZN(new_n5192_));
  AOI21_X1   g5135(.A1(new_n5192_), .A2(new_n5190_), .B(new_n5172_), .ZN(new_n5193_));
  INV_X1     g5136(.I(new_n5172_), .ZN(new_n5194_));
  AOI21_X1   g5137(.A1(new_n5183_), .A2(new_n5180_), .B(new_n2720_), .ZN(new_n5195_));
  INV_X1     g5138(.I(new_n5184_), .ZN(new_n5196_));
  OAI21_X1   g5139(.A1(new_n5196_), .A2(new_n5195_), .B(new_n5189_), .ZN(new_n5197_));
  NAND3_X1   g5140(.A1(new_n5182_), .A2(new_n5184_), .A3(new_n5188_), .ZN(new_n5198_));
  AOI21_X1   g5141(.A1(new_n5197_), .A2(new_n5198_), .B(new_n5194_), .ZN(new_n5199_));
  NOR2_X1    g5142(.A1(new_n5065_), .A2(new_n5056_), .ZN(new_n5200_));
  NOR2_X1    g5143(.A1(new_n5200_), .A2(new_n5062_), .ZN(new_n5201_));
  NAND2_X1   g5144(.A1(new_n5200_), .A2(new_n5062_), .ZN(new_n5202_));
  XOR2_X1    g5145(.A1(new_n5051_), .A2(new_n5048_), .Z(new_n5203_));
  INV_X1     g5146(.I(new_n5203_), .ZN(new_n5204_));
  AOI21_X1   g5147(.A1(new_n5204_), .A2(new_n5202_), .B(new_n5201_), .ZN(new_n5205_));
  INV_X1     g5148(.I(new_n5205_), .ZN(new_n5206_));
  OAI21_X1   g5149(.A1(new_n5193_), .A2(new_n5199_), .B(new_n5206_), .ZN(new_n5207_));
  INV_X1     g5150(.I(new_n5190_), .ZN(new_n5208_));
  OAI21_X1   g5151(.A1(new_n5208_), .A2(new_n5191_), .B(new_n5194_), .ZN(new_n5209_));
  AOI21_X1   g5152(.A1(new_n5182_), .A2(new_n5184_), .B(new_n5188_), .ZN(new_n5210_));
  INV_X1     g5153(.I(new_n5198_), .ZN(new_n5211_));
  OAI21_X1   g5154(.A1(new_n5211_), .A2(new_n5210_), .B(new_n5172_), .ZN(new_n5212_));
  NAND3_X1   g5155(.A1(new_n5209_), .A2(new_n5212_), .A3(new_n5205_), .ZN(new_n5213_));
  AOI21_X1   g5156(.A1(new_n5213_), .A2(new_n5207_), .B(new_n5167_), .ZN(new_n5214_));
  INV_X1     g5157(.I(new_n5167_), .ZN(new_n5215_));
  NAND3_X1   g5158(.A1(new_n5209_), .A2(new_n5212_), .A3(new_n5206_), .ZN(new_n5216_));
  OAI21_X1   g5159(.A1(new_n5193_), .A2(new_n5199_), .B(new_n5205_), .ZN(new_n5217_));
  AOI21_X1   g5160(.A1(new_n5216_), .A2(new_n5217_), .B(new_n5215_), .ZN(new_n5218_));
  AOI22_X1   g5161(.A1(new_n4747_), .A2(new_n3210_), .B1(new_n3280_), .B2(new_n4475_), .ZN(new_n5219_));
  INV_X1     g5162(.I(new_n5219_), .ZN(new_n5220_));
  OAI21_X1   g5163(.A1(new_n5079_), .A2(new_n5078_), .B(new_n5082_), .ZN(new_n5221_));
  NAND3_X1   g5164(.A1(new_n5072_), .A2(new_n5076_), .A3(new_n5037_), .ZN(new_n5222_));
  NAND2_X1   g5165(.A1(new_n5043_), .A2(new_n803_), .ZN(new_n5223_));
  NAND3_X1   g5166(.A1(new_n5038_), .A2(new_n802_), .A3(new_n5042_), .ZN(new_n5224_));
  NAND2_X1   g5167(.A1(new_n5223_), .A2(new_n5224_), .ZN(new_n5225_));
  NAND2_X1   g5168(.A1(new_n5222_), .A2(new_n5225_), .ZN(new_n5226_));
  AOI21_X1   g5169(.A1(new_n5226_), .A2(new_n5221_), .B(new_n5220_), .ZN(new_n5227_));
  NOR2_X1    g5170(.A1(new_n5079_), .A2(new_n5078_), .ZN(new_n5228_));
  NOR2_X1    g5171(.A1(new_n5228_), .A2(new_n5037_), .ZN(new_n5229_));
  AOI22_X1   g5172(.A1(new_n5228_), .A2(new_n5037_), .B1(new_n5223_), .B2(new_n5224_), .ZN(new_n5230_));
  NOR3_X1    g5173(.A1(new_n5230_), .A2(new_n5219_), .A3(new_n5229_), .ZN(new_n5231_));
  NOR2_X1    g5174(.A1(new_n5231_), .A2(new_n5227_), .ZN(new_n5232_));
  NOR3_X1    g5175(.A1(new_n5214_), .A2(new_n5218_), .A3(new_n5232_), .ZN(new_n5233_));
  AOI21_X1   g5176(.A1(new_n5209_), .A2(new_n5212_), .B(new_n5205_), .ZN(new_n5234_));
  NOR3_X1    g5177(.A1(new_n5193_), .A2(new_n5199_), .A3(new_n5206_), .ZN(new_n5235_));
  OAI21_X1   g5178(.A1(new_n5234_), .A2(new_n5235_), .B(new_n5215_), .ZN(new_n5236_));
  NOR3_X1    g5179(.A1(new_n5193_), .A2(new_n5199_), .A3(new_n5205_), .ZN(new_n5237_));
  AOI21_X1   g5180(.A1(new_n5209_), .A2(new_n5212_), .B(new_n5206_), .ZN(new_n5238_));
  OAI21_X1   g5181(.A1(new_n5238_), .A2(new_n5237_), .B(new_n5167_), .ZN(new_n5239_));
  OAI21_X1   g5182(.A1(new_n5230_), .A2(new_n5229_), .B(new_n5219_), .ZN(new_n5240_));
  NAND3_X1   g5183(.A1(new_n5226_), .A2(new_n5220_), .A3(new_n5221_), .ZN(new_n5241_));
  NAND2_X1   g5184(.A1(new_n5240_), .A2(new_n5241_), .ZN(new_n5242_));
  AOI21_X1   g5185(.A1(new_n5236_), .A2(new_n5239_), .B(new_n5242_), .ZN(new_n5243_));
  OAI21_X1   g5186(.A1(new_n5233_), .A2(new_n5243_), .B(new_n1050_), .ZN(new_n5244_));
  NAND3_X1   g5187(.A1(new_n5236_), .A2(new_n5239_), .A3(new_n5242_), .ZN(new_n5245_));
  OAI21_X1   g5188(.A1(new_n5214_), .A2(new_n5218_), .B(new_n5232_), .ZN(new_n5246_));
  NAND3_X1   g5189(.A1(new_n5246_), .A2(new_n5245_), .A3(new_n1051_), .ZN(new_n5247_));
  NAND3_X1   g5190(.A1(new_n5244_), .A2(new_n5247_), .A3(new_n5163_), .ZN(new_n5248_));
  AOI21_X1   g5191(.A1(new_n5246_), .A2(new_n5245_), .B(new_n1051_), .ZN(new_n5249_));
  NOR3_X1    g5192(.A1(new_n5233_), .A2(new_n5243_), .A3(new_n1050_), .ZN(new_n5250_));
  OAI21_X1   g5193(.A1(new_n5249_), .A2(new_n5250_), .B(new_n5162_), .ZN(new_n5251_));
  NAND2_X1   g5194(.A1(new_n5251_), .A2(new_n5248_), .ZN(new_n5252_));
  XOR2_X1    g5195(.A1(new_n5100_), .A2(new_n5029_), .Z(new_n5253_));
  NAND3_X1   g5196(.A1(new_n5253_), .A2(new_n5252_), .A3(new_n5110_), .ZN(new_n5254_));
  NOR3_X1    g5197(.A1(new_n5249_), .A2(new_n5250_), .A3(new_n5162_), .ZN(new_n5255_));
  AOI21_X1   g5198(.A1(new_n5244_), .A2(new_n5247_), .B(new_n5163_), .ZN(new_n5256_));
  NOR2_X1    g5199(.A1(new_n5256_), .A2(new_n5255_), .ZN(new_n5257_));
  NOR2_X1    g5200(.A1(new_n5100_), .A2(new_n5029_), .ZN(new_n5258_));
  INV_X1     g5201(.I(new_n5258_), .ZN(new_n5259_));
  NAND2_X1   g5202(.A1(new_n5254_), .A2(new_n5259_), .ZN(new_n5260_));
  NAND3_X1   g5203(.A1(new_n5260_), .A2(new_n5129_), .A3(new_n5128_), .ZN(new_n5261_));
  NAND2_X1   g5204(.A1(new_n5129_), .A2(new_n5128_), .ZN(new_n5262_));
  XOR2_X1    g5205(.A1(new_n5100_), .A2(new_n5102_), .Z(new_n5263_));
  NOR3_X1    g5206(.A1(new_n5263_), .A2(new_n5257_), .A3(new_n5124_), .ZN(new_n5264_));
  NOR2_X1    g5207(.A1(new_n5264_), .A2(new_n5258_), .ZN(new_n5265_));
  NAND2_X1   g5208(.A1(new_n5262_), .A2(new_n5265_), .ZN(new_n5266_));
  NAND2_X1   g5209(.A1(new_n5266_), .A2(new_n5261_), .ZN(new_n5267_));
  NAND4_X1   g5210(.A1(new_n476_), .A2(new_n921_), .A3(new_n388_), .A4(new_n514_), .ZN(new_n5268_));
  NOR4_X1    g5211(.A1(new_n2505_), .A2(new_n292_), .A3(new_n383_), .A4(new_n517_), .ZN(new_n5269_));
  NAND2_X1   g5212(.A1(new_n5269_), .A2(new_n2439_), .ZN(new_n5270_));
  NOR4_X1    g5213(.A1(new_n5270_), .A2(new_n461_), .A3(new_n2334_), .A4(new_n5268_), .ZN(new_n5271_));
  NAND2_X1   g5214(.A1(new_n363_), .A2(new_n407_), .ZN(new_n5272_));
  NAND2_X1   g5215(.A1(new_n3967_), .A2(new_n1238_), .ZN(new_n5273_));
  NOR4_X1    g5216(.A1(new_n5273_), .A2(new_n593_), .A3(new_n857_), .A4(new_n5272_), .ZN(new_n5274_));
  NAND4_X1   g5217(.A1(new_n5271_), .A2(new_n4063_), .A3(new_n2404_), .A4(new_n5274_), .ZN(new_n5275_));
  INV_X1     g5218(.I(new_n5275_), .ZN(new_n5276_));
  NOR2_X1    g5219(.A1(new_n5267_), .A2(new_n5276_), .ZN(new_n5277_));
  NOR2_X1    g5220(.A1(new_n5262_), .A2(new_n5265_), .ZN(new_n5278_));
  AOI21_X1   g5221(.A1(new_n5128_), .A2(new_n5129_), .B(new_n5260_), .ZN(new_n5279_));
  NOR2_X1    g5222(.A1(new_n5278_), .A2(new_n5279_), .ZN(new_n5280_));
  NOR2_X1    g5223(.A1(new_n5280_), .A2(new_n5275_), .ZN(new_n5281_));
  NOR2_X1    g5224(.A1(new_n5281_), .A2(new_n5277_), .ZN(new_n5282_));
  NAND2_X1   g5225(.A1(new_n5161_), .A2(new_n5282_), .ZN(new_n5283_));
  OAI22_X1   g5226(.A1(new_n5160_), .A2(new_n5157_), .B1(new_n5281_), .B2(new_n5277_), .ZN(new_n5284_));
  NAND2_X1   g5227(.A1(new_n5283_), .A2(new_n5284_), .ZN(new_n5285_));
  XOR2_X1    g5228(.A1(new_n5285_), .A2(new_n5152_), .Z(new_n5286_));
  NOR2_X1    g5229(.A1(new_n5145_), .A2(new_n5142_), .ZN(new_n5287_));
  INV_X1     g5230(.I(new_n5139_), .ZN(new_n5288_));
  OAI21_X1   g5231(.A1(new_n5141_), .A2(new_n5288_), .B(new_n5287_), .ZN(new_n5289_));
  NAND3_X1   g5232(.A1(new_n5137_), .A2(new_n5135_), .A3(new_n5139_), .ZN(new_n5290_));
  NAND2_X1   g5233(.A1(new_n5289_), .A2(new_n5290_), .ZN(new_n5291_));
  NOR3_X1    g5234(.A1(new_n4878_), .A2(new_n4882_), .A3(new_n5291_), .ZN(new_n5292_));
  NOR2_X1    g5235(.A1(new_n5018_), .A2(new_n5148_), .ZN(new_n5293_));
  AOI21_X1   g5236(.A1(new_n5015_), .A2(new_n5016_), .B(new_n5024_), .ZN(new_n5294_));
  OAI21_X1   g5237(.A1(new_n5293_), .A2(new_n5292_), .B(new_n5294_), .ZN(new_n5295_));
  NAND2_X1   g5238(.A1(new_n5295_), .A2(new_n4404_), .ZN(new_n5296_));
  XOR2_X1    g5239(.A1(new_n5296_), .A2(new_n5286_), .Z(\sin[6] ));
  INV_X1     g5240(.I(new_n5295_), .ZN(new_n5298_));
  AOI21_X1   g5241(.A1(new_n5298_), .A2(new_n5286_), .B(new_n4445_), .ZN(new_n5299_));
  NAND2_X1   g5242(.A1(new_n5024_), .A2(new_n5291_), .ZN(new_n5300_));
  NAND3_X1   g5243(.A1(new_n5148_), .A2(new_n5014_), .A3(new_n4896_), .ZN(new_n5301_));
  AOI21_X1   g5244(.A1(new_n5300_), .A2(new_n5301_), .B(new_n5284_), .ZN(new_n5302_));
  NAND2_X1   g5245(.A1(new_n5244_), .A2(new_n5247_), .ZN(new_n5303_));
  NAND2_X1   g5246(.A1(new_n5303_), .A2(new_n5163_), .ZN(new_n5304_));
  INV_X1     g5247(.I(new_n5304_), .ZN(new_n5305_));
  NOR3_X1    g5248(.A1(new_n5256_), .A2(new_n5255_), .A3(new_n5109_), .ZN(new_n5306_));
  OAI21_X1   g5249(.A1(new_n5256_), .A2(new_n5255_), .B(new_n5109_), .ZN(new_n5307_));
  AOI21_X1   g5250(.A1(new_n5029_), .A2(new_n5307_), .B(new_n5306_), .ZN(new_n5308_));
  OAI21_X1   g5251(.A1(new_n5027_), .A2(new_n4989_), .B(new_n5308_), .ZN(new_n5309_));
  NOR2_X1    g5252(.A1(new_n5230_), .A2(new_n5229_), .ZN(new_n5310_));
  AOI21_X1   g5253(.A1(new_n5236_), .A2(new_n5239_), .B(new_n5310_), .ZN(new_n5311_));
  NOR4_X1    g5254(.A1(new_n5214_), .A2(new_n5218_), .A3(new_n5229_), .A4(new_n5230_), .ZN(new_n5312_));
  XOR2_X1    g5255(.A1(new_n5219_), .A2(new_n1051_), .Z(new_n5313_));
  NOR2_X1    g5256(.A1(new_n5312_), .A2(new_n5313_), .ZN(new_n5314_));
  NOR2_X1    g5257(.A1(new_n5314_), .A2(new_n5311_), .ZN(new_n5315_));
  AOI21_X1   g5258(.A1(new_n5215_), .A2(new_n5217_), .B(new_n5237_), .ZN(new_n5316_));
  INV_X1     g5259(.I(new_n5316_), .ZN(new_n5317_));
  OAI22_X1   g5260(.A1(new_n4230_), .A2(new_n2975_), .B1(new_n4182_), .B2(new_n2972_), .ZN(new_n5318_));
  OAI21_X1   g5261(.A1(new_n2969_), .A2(new_n4474_), .B(new_n5318_), .ZN(new_n5319_));
  AOI21_X1   g5262(.A1(new_n5319_), .A2(new_n802_), .B(new_n2969_), .ZN(new_n5320_));
  XOR2_X1    g5263(.A1(new_n4484_), .A2(new_n5320_), .Z(new_n5321_));
  INV_X1     g5264(.I(new_n5321_), .ZN(new_n5322_));
  AOI21_X1   g5265(.A1(new_n5172_), .A2(new_n5190_), .B(new_n5191_), .ZN(new_n5323_));
  NOR2_X1    g5266(.A1(new_n5177_), .A2(new_n2943_), .ZN(new_n5324_));
  NAND2_X1   g5267(.A1(new_n2720_), .A2(new_n438_), .ZN(new_n5325_));
  OAI21_X1   g5268(.A1(new_n5324_), .A2(new_n5325_), .B(new_n5178_), .ZN(new_n5326_));
  AOI22_X1   g5269(.A1(new_n2898_), .A2(new_n3494_), .B1(new_n3436_), .B2(new_n3398_), .ZN(new_n5327_));
  NOR2_X1    g5270(.A1(new_n2879_), .A2(new_n3396_), .ZN(new_n5328_));
  OAI21_X1   g5271(.A1(new_n5327_), .A2(new_n5328_), .B(new_n437_), .ZN(new_n5329_));
  NAND2_X1   g5272(.A1(new_n5329_), .A2(new_n3393_), .ZN(new_n5330_));
  XOR2_X1    g5273(.A1(new_n3844_), .A2(new_n5330_), .Z(new_n5331_));
  NAND2_X1   g5274(.A1(new_n3182_), .A2(new_n437_), .ZN(new_n5332_));
  NAND2_X1   g5275(.A1(new_n1051_), .A2(new_n2943_), .ZN(new_n5333_));
  NAND2_X1   g5276(.A1(new_n1050_), .A2(new_n2942_), .ZN(new_n5334_));
  AOI21_X1   g5277(.A1(new_n5333_), .A2(new_n5334_), .B(new_n5332_), .ZN(new_n5335_));
  AOI21_X1   g5278(.A1(new_n3182_), .A2(new_n437_), .B(new_n3209_), .ZN(new_n5336_));
  NOR2_X1    g5279(.A1(new_n5335_), .A2(new_n5336_), .ZN(new_n5337_));
  INV_X1     g5280(.I(new_n5337_), .ZN(new_n5338_));
  NAND2_X1   g5281(.A1(new_n5331_), .A2(new_n5338_), .ZN(new_n5339_));
  NOR2_X1    g5282(.A1(new_n5331_), .A2(new_n5338_), .ZN(new_n5340_));
  INV_X1     g5283(.I(new_n5340_), .ZN(new_n5341_));
  NAND2_X1   g5284(.A1(new_n5341_), .A2(new_n5339_), .ZN(new_n5342_));
  AND2_X2    g5285(.A1(new_n5342_), .A2(new_n5326_), .Z(new_n5343_));
  XOR2_X1    g5286(.A1(new_n5331_), .A2(new_n5337_), .Z(new_n5344_));
  NOR2_X1    g5287(.A1(new_n5344_), .A2(new_n5326_), .ZN(new_n5345_));
  NOR2_X1    g5288(.A1(new_n5343_), .A2(new_n5345_), .ZN(new_n5346_));
  AOI22_X1   g5289(.A1(new_n2946_), .A2(new_n3038_), .B1(new_n3985_), .B2(new_n3030_), .ZN(new_n5347_));
  NOR2_X1    g5290(.A1(new_n3987_), .A2(new_n3028_), .ZN(new_n5348_));
  OAI21_X1   g5291(.A1(new_n5348_), .A2(new_n5347_), .B(new_n721_), .ZN(new_n5349_));
  NAND2_X1   g5292(.A1(new_n5349_), .A2(new_n2992_), .ZN(new_n5350_));
  XOR2_X1    g5293(.A1(new_n3982_), .A2(new_n5350_), .Z(new_n5351_));
  INV_X1     g5294(.I(new_n5351_), .ZN(new_n5352_));
  NAND2_X1   g5295(.A1(new_n5346_), .A2(new_n5352_), .ZN(new_n5353_));
  OAI21_X1   g5296(.A1(new_n5343_), .A2(new_n5345_), .B(new_n5351_), .ZN(new_n5354_));
  AOI21_X1   g5297(.A1(new_n5353_), .A2(new_n5354_), .B(new_n5323_), .ZN(new_n5355_));
  INV_X1     g5298(.I(new_n5323_), .ZN(new_n5356_));
  XOR2_X1    g5299(.A1(new_n5346_), .A2(new_n5351_), .Z(new_n5357_));
  NOR2_X1    g5300(.A1(new_n5357_), .A2(new_n5356_), .ZN(new_n5358_));
  NOR2_X1    g5301(.A1(new_n5358_), .A2(new_n5355_), .ZN(new_n5359_));
  NOR2_X1    g5302(.A1(new_n5359_), .A2(new_n5322_), .ZN(new_n5360_));
  INV_X1     g5303(.I(new_n5355_), .ZN(new_n5361_));
  XOR2_X1    g5304(.A1(new_n5346_), .A2(new_n5352_), .Z(new_n5362_));
  NAND2_X1   g5305(.A1(new_n5362_), .A2(new_n5323_), .ZN(new_n5363_));
  NAND2_X1   g5306(.A1(new_n5363_), .A2(new_n5361_), .ZN(new_n5364_));
  NOR2_X1    g5307(.A1(new_n5364_), .A2(new_n5321_), .ZN(new_n5365_));
  OAI21_X1   g5308(.A1(new_n5360_), .A2(new_n5365_), .B(new_n5317_), .ZN(new_n5366_));
  NOR2_X1    g5309(.A1(new_n5359_), .A2(new_n5321_), .ZN(new_n5367_));
  NOR2_X1    g5310(.A1(new_n5364_), .A2(new_n5322_), .ZN(new_n5368_));
  OAI21_X1   g5311(.A1(new_n5367_), .A2(new_n5368_), .B(new_n5316_), .ZN(new_n5369_));
  NAND3_X1   g5312(.A1(new_n5366_), .A2(new_n5369_), .A3(new_n5315_), .ZN(new_n5370_));
  INV_X1     g5313(.I(new_n5370_), .ZN(new_n5371_));
  AOI21_X1   g5314(.A1(new_n5369_), .A2(new_n5366_), .B(new_n5315_), .ZN(new_n5372_));
  INV_X1     g5315(.I(new_n5271_), .ZN(new_n5373_));
  NOR2_X1    g5316(.A1(new_n233_), .A2(new_n251_), .ZN(new_n5374_));
  NAND4_X1   g5317(.A1(new_n320_), .A2(new_n5374_), .A3(new_n777_), .A4(new_n313_), .ZN(new_n5375_));
  NOR3_X1    g5318(.A1(new_n892_), .A2(new_n203_), .A3(new_n421_), .ZN(new_n5376_));
  NAND4_X1   g5319(.A1(new_n5376_), .A2(new_n156_), .A3(new_n5113_), .A4(new_n380_), .ZN(new_n5377_));
  NOR3_X1    g5320(.A1(new_n5373_), .A2(new_n5375_), .A3(new_n5377_), .ZN(new_n5378_));
  AND2_X2    g5321(.A1(new_n2236_), .A2(new_n5378_), .Z(new_n5379_));
  OAI21_X1   g5322(.A1(new_n5371_), .A2(new_n5372_), .B(new_n5379_), .ZN(new_n5380_));
  INV_X1     g5323(.I(new_n5380_), .ZN(new_n5381_));
  NAND2_X1   g5324(.A1(new_n5309_), .A2(new_n5381_), .ZN(new_n5382_));
  NAND3_X1   g5325(.A1(new_n5262_), .A2(new_n5308_), .A3(new_n5380_), .ZN(new_n5383_));
  AOI21_X1   g5326(.A1(new_n5382_), .A2(new_n5383_), .B(new_n5305_), .ZN(new_n5384_));
  NAND3_X1   g5327(.A1(new_n5251_), .A2(new_n5248_), .A3(new_n5100_), .ZN(new_n5385_));
  AOI21_X1   g5328(.A1(new_n5251_), .A2(new_n5248_), .B(new_n5100_), .ZN(new_n5386_));
  OAI21_X1   g5329(.A1(new_n5102_), .A2(new_n5386_), .B(new_n5385_), .ZN(new_n5387_));
  AOI21_X1   g5330(.A1(new_n5129_), .A2(new_n5128_), .B(new_n5387_), .ZN(new_n5388_));
  NOR2_X1    g5331(.A1(new_n5388_), .A2(new_n5380_), .ZN(new_n5389_));
  NOR2_X1    g5332(.A1(new_n5309_), .A2(new_n5381_), .ZN(new_n5390_));
  NOR3_X1    g5333(.A1(new_n5390_), .A2(new_n5389_), .A3(new_n5304_), .ZN(new_n5391_));
  NOR2_X1    g5334(.A1(new_n5391_), .A2(new_n5384_), .ZN(new_n5392_));
  AOI21_X1   g5335(.A1(new_n5266_), .A2(new_n5261_), .B(new_n5276_), .ZN(new_n5393_));
  NOR3_X1    g5336(.A1(new_n5278_), .A2(new_n5279_), .A3(new_n5275_), .ZN(new_n5394_));
  NOR2_X1    g5337(.A1(new_n5394_), .A2(new_n5393_), .ZN(new_n5395_));
  NOR3_X1    g5338(.A1(new_n5392_), .A2(new_n5281_), .A3(new_n5395_), .ZN(new_n5396_));
  NOR2_X1    g5339(.A1(new_n5280_), .A2(new_n5275_), .ZN(new_n5397_));
  OAI21_X1   g5340(.A1(new_n5396_), .A2(new_n5397_), .B(new_n5161_), .ZN(new_n5398_));
  NAND2_X1   g5341(.A1(new_n5262_), .A2(new_n5111_), .ZN(new_n5399_));
  NAND2_X1   g5342(.A1(new_n5399_), .A2(new_n5153_), .ZN(new_n5400_));
  NAND2_X1   g5343(.A1(new_n5141_), .A2(new_n5400_), .ZN(new_n5401_));
  OAI21_X1   g5344(.A1(new_n5141_), .A2(new_n5400_), .B(new_n5158_), .ZN(new_n5402_));
  NAND2_X1   g5345(.A1(new_n5402_), .A2(new_n5401_), .ZN(new_n5403_));
  NAND2_X1   g5346(.A1(new_n5267_), .A2(new_n5276_), .ZN(new_n5404_));
  OAI21_X1   g5347(.A1(new_n5390_), .A2(new_n5389_), .B(new_n5304_), .ZN(new_n5405_));
  NAND3_X1   g5348(.A1(new_n5382_), .A2(new_n5383_), .A3(new_n5305_), .ZN(new_n5406_));
  NAND2_X1   g5349(.A1(new_n5405_), .A2(new_n5406_), .ZN(new_n5407_));
  OAI21_X1   g5350(.A1(new_n5278_), .A2(new_n5279_), .B(new_n5275_), .ZN(new_n5408_));
  NAND3_X1   g5351(.A1(new_n5266_), .A2(new_n5261_), .A3(new_n5276_), .ZN(new_n5409_));
  NAND2_X1   g5352(.A1(new_n5408_), .A2(new_n5409_), .ZN(new_n5410_));
  NAND3_X1   g5353(.A1(new_n5407_), .A2(new_n5404_), .A3(new_n5410_), .ZN(new_n5411_));
  INV_X1     g5354(.I(new_n5397_), .ZN(new_n5412_));
  NAND3_X1   g5355(.A1(new_n5411_), .A2(new_n5412_), .A3(new_n5403_), .ZN(new_n5413_));
  NAND2_X1   g5356(.A1(new_n5398_), .A2(new_n5413_), .ZN(new_n5414_));
  NAND2_X1   g5357(.A1(new_n5414_), .A2(new_n5302_), .ZN(new_n5415_));
  NOR2_X1    g5358(.A1(new_n5161_), .A2(new_n5282_), .ZN(new_n5416_));
  AOI21_X1   g5359(.A1(new_n4896_), .A2(new_n5014_), .B(new_n5148_), .ZN(new_n5417_));
  NOR2_X1    g5360(.A1(new_n5024_), .A2(new_n5291_), .ZN(new_n5418_));
  OAI21_X1   g5361(.A1(new_n5417_), .A2(new_n5418_), .B(new_n5416_), .ZN(new_n5419_));
  AOI21_X1   g5362(.A1(new_n5411_), .A2(new_n5412_), .B(new_n5403_), .ZN(new_n5420_));
  NOR3_X1    g5363(.A1(new_n5396_), .A2(new_n5161_), .A3(new_n5397_), .ZN(new_n5421_));
  NOR2_X1    g5364(.A1(new_n5421_), .A2(new_n5420_), .ZN(new_n5422_));
  NAND2_X1   g5365(.A1(new_n5422_), .A2(new_n5419_), .ZN(new_n5423_));
  NAND2_X1   g5366(.A1(new_n5423_), .A2(new_n5415_), .ZN(new_n5424_));
  NAND2_X1   g5367(.A1(new_n5299_), .A2(new_n5424_), .ZN(new_n5425_));
  XOR2_X1    g5368(.A1(new_n5422_), .A2(new_n5302_), .Z(new_n5426_));
  OAI21_X1   g5369(.A1(new_n5299_), .A2(new_n5426_), .B(new_n5425_), .ZN(\sin[7] ));
  INV_X1     g5370(.I(new_n5285_), .ZN(new_n5428_));
  XOR2_X1    g5371(.A1(new_n5018_), .A2(new_n5291_), .Z(new_n5429_));
  NAND3_X1   g5372(.A1(new_n5429_), .A2(new_n5428_), .A3(new_n5294_), .ZN(new_n5430_));
  NAND2_X1   g5373(.A1(new_n5295_), .A2(new_n5285_), .ZN(new_n5431_));
  NOR2_X1    g5374(.A1(new_n5422_), .A2(new_n5285_), .ZN(new_n5432_));
  NOR2_X1    g5375(.A1(new_n5428_), .A2(new_n5414_), .ZN(new_n5433_));
  OAI21_X1   g5376(.A1(new_n5433_), .A2(new_n5432_), .B(new_n5149_), .ZN(new_n5434_));
  AOI21_X1   g5377(.A1(new_n5430_), .A2(new_n5431_), .B(new_n5434_), .ZN(new_n5435_));
  INV_X1     g5378(.I(new_n5315_), .ZN(new_n5436_));
  NAND2_X1   g5379(.A1(new_n5305_), .A2(new_n5436_), .ZN(new_n5437_));
  AOI22_X1   g5380(.A1(new_n5304_), .A2(new_n5315_), .B1(new_n5366_), .B2(new_n5369_), .ZN(new_n5438_));
  INV_X1     g5381(.I(new_n5438_), .ZN(new_n5439_));
  OAI21_X1   g5382(.A1(new_n5309_), .A2(new_n5439_), .B(new_n5437_), .ZN(new_n5440_));
  INV_X1     g5383(.I(new_n5360_), .ZN(new_n5441_));
  OAI21_X1   g5384(.A1(new_n5316_), .A2(new_n5365_), .B(new_n5441_), .ZN(new_n5442_));
  NAND2_X1   g5385(.A1(new_n4786_), .A2(new_n802_), .ZN(new_n5443_));
  OAI21_X1   g5386(.A1(new_n4480_), .A2(new_n5443_), .B(new_n2977_), .ZN(new_n5444_));
  XOR2_X1    g5387(.A1(new_n4688_), .A2(new_n5444_), .Z(new_n5445_));
  INV_X1     g5388(.I(new_n5445_), .ZN(new_n5446_));
  AOI22_X1   g5389(.A1(new_n2898_), .A2(new_n3494_), .B1(new_n2879_), .B2(new_n4270_), .ZN(new_n5447_));
  AOI21_X1   g5390(.A1(new_n2946_), .A2(new_n3398_), .B(new_n5447_), .ZN(new_n5448_));
  OAI21_X1   g5391(.A1(new_n5448_), .A2(new_n438_), .B(new_n3393_), .ZN(new_n5449_));
  XNOR2_X1   g5392(.A1(new_n2935_), .A2(new_n5449_), .ZN(new_n5450_));
  NAND2_X1   g5393(.A1(new_n5332_), .A2(new_n5333_), .ZN(new_n5451_));
  NAND2_X1   g5394(.A1(new_n5451_), .A2(new_n5334_), .ZN(new_n5452_));
  INV_X1     g5395(.I(new_n5452_), .ZN(new_n5453_));
  NOR2_X1    g5396(.A1(new_n2682_), .A2(new_n438_), .ZN(new_n5454_));
  INV_X1     g5397(.I(new_n5454_), .ZN(new_n5455_));
  NOR2_X1    g5398(.A1(new_n5453_), .A2(new_n5455_), .ZN(new_n5456_));
  NOR2_X1    g5399(.A1(new_n5452_), .A2(new_n5454_), .ZN(new_n5457_));
  OAI21_X1   g5400(.A1(new_n5456_), .A2(new_n5457_), .B(new_n5450_), .ZN(new_n5458_));
  XOR2_X1    g5401(.A1(new_n5452_), .A2(new_n5455_), .Z(new_n5459_));
  OR2_X2     g5402(.A1(new_n5450_), .A2(new_n5459_), .Z(new_n5460_));
  NAND2_X1   g5403(.A1(new_n5460_), .A2(new_n5458_), .ZN(new_n5461_));
  INV_X1     g5404(.I(new_n5461_), .ZN(new_n5462_));
  AND2_X2    g5405(.A1(new_n5339_), .A2(new_n5326_), .Z(new_n5463_));
  NOR2_X1    g5406(.A1(new_n5463_), .A2(new_n5340_), .ZN(new_n5464_));
  NOR2_X1    g5407(.A1(new_n4198_), .A2(new_n2991_), .ZN(new_n5465_));
  OAI22_X1   g5408(.A1(new_n3987_), .A2(new_n3031_), .B1(new_n2994_), .B2(new_n3597_), .ZN(new_n5466_));
  OAI21_X1   g5409(.A1(new_n3028_), .A2(new_n4192_), .B(new_n5466_), .ZN(new_n5467_));
  NOR2_X1    g5410(.A1(new_n5465_), .A2(new_n5467_), .ZN(new_n5468_));
  NAND2_X1   g5411(.A1(new_n5464_), .A2(new_n5468_), .ZN(new_n5469_));
  INV_X1     g5412(.I(new_n5469_), .ZN(new_n5470_));
  NOR2_X1    g5413(.A1(new_n5464_), .A2(new_n5468_), .ZN(new_n5471_));
  OAI21_X1   g5414(.A1(new_n5470_), .A2(new_n5471_), .B(new_n5462_), .ZN(new_n5472_));
  INV_X1     g5415(.I(new_n5471_), .ZN(new_n5473_));
  NAND3_X1   g5416(.A1(new_n5473_), .A2(new_n5461_), .A3(new_n5469_), .ZN(new_n5474_));
  AOI21_X1   g5417(.A1(new_n5472_), .A2(new_n5474_), .B(new_n702_), .ZN(new_n5475_));
  NAND3_X1   g5418(.A1(new_n5472_), .A2(new_n5474_), .A3(new_n702_), .ZN(new_n5476_));
  INV_X1     g5419(.I(new_n5476_), .ZN(new_n5477_));
  OAI21_X1   g5420(.A1(new_n5477_), .A2(new_n5475_), .B(new_n5446_), .ZN(new_n5478_));
  NOR2_X1    g5421(.A1(new_n5478_), .A2(new_n5358_), .ZN(new_n5479_));
  AOI21_X1   g5422(.A1(new_n5473_), .A2(new_n5469_), .B(new_n5461_), .ZN(new_n5480_));
  INV_X1     g5423(.I(new_n5474_), .ZN(new_n5481_));
  OAI21_X1   g5424(.A1(new_n5481_), .A2(new_n5480_), .B(new_n721_), .ZN(new_n5482_));
  AOI21_X1   g5425(.A1(new_n5482_), .A2(new_n5476_), .B(new_n5445_), .ZN(new_n5483_));
  NOR2_X1    g5426(.A1(new_n5483_), .A2(new_n5363_), .ZN(new_n5484_));
  OAI21_X1   g5427(.A1(new_n5479_), .A2(new_n5484_), .B(new_n5353_), .ZN(new_n5485_));
  NAND2_X1   g5428(.A1(new_n5483_), .A2(new_n5363_), .ZN(new_n5486_));
  NAND2_X1   g5429(.A1(new_n5478_), .A2(new_n5358_), .ZN(new_n5487_));
  NAND4_X1   g5430(.A1(new_n5487_), .A2(new_n5486_), .A3(new_n5346_), .A4(new_n5352_), .ZN(new_n5488_));
  NAND2_X1   g5431(.A1(new_n5488_), .A2(new_n5485_), .ZN(new_n5489_));
  NOR2_X1    g5432(.A1(new_n5489_), .A2(new_n5442_), .ZN(new_n5490_));
  NAND2_X1   g5433(.A1(new_n5489_), .A2(new_n5442_), .ZN(new_n5491_));
  INV_X1     g5434(.I(new_n5491_), .ZN(new_n5492_));
  NOR2_X1    g5435(.A1(new_n5492_), .A2(new_n5490_), .ZN(new_n5493_));
  INV_X1     g5436(.I(new_n5493_), .ZN(new_n5494_));
  INV_X1     g5437(.I(new_n4042_), .ZN(new_n5495_));
  NOR4_X1    g5438(.A1(new_n283_), .A2(new_n110_), .A3(new_n132_), .A4(new_n465_), .ZN(new_n5496_));
  NOR4_X1    g5439(.A1(new_n227_), .A2(new_n388_), .A3(new_n454_), .A4(new_n311_), .ZN(new_n5497_));
  NAND3_X1   g5440(.A1(new_n2390_), .A2(new_n5496_), .A3(new_n5497_), .ZN(new_n5498_));
  NOR2_X1    g5441(.A1(new_n2435_), .A2(new_n5498_), .ZN(new_n5499_));
  INV_X1     g5442(.I(new_n5499_), .ZN(new_n5500_));
  NOR4_X1    g5443(.A1(new_n754_), .A2(new_n281_), .A3(new_n398_), .A4(new_n675_), .ZN(new_n5501_));
  NOR4_X1    g5444(.A1(new_n372_), .A2(new_n187_), .A3(new_n201_), .A4(new_n625_), .ZN(new_n5502_));
  NAND4_X1   g5445(.A1(new_n5501_), .A2(new_n853_), .A3(new_n2500_), .A4(new_n5502_), .ZN(new_n5503_));
  NOR3_X1    g5446(.A1(new_n5495_), .A2(new_n5500_), .A3(new_n5503_), .ZN(new_n5504_));
  NAND2_X1   g5447(.A1(new_n5494_), .A2(new_n5504_), .ZN(new_n5505_));
  INV_X1     g5448(.I(new_n5504_), .ZN(new_n5506_));
  NAND2_X1   g5449(.A1(new_n5493_), .A2(new_n5506_), .ZN(new_n5507_));
  NAND2_X1   g5450(.A1(new_n5505_), .A2(new_n5507_), .ZN(new_n5508_));
  NAND2_X1   g5451(.A1(new_n5508_), .A2(new_n5440_), .ZN(new_n5509_));
  AOI22_X1   g5452(.A1(new_n5388_), .A2(new_n5438_), .B1(new_n5305_), .B2(new_n5436_), .ZN(new_n5510_));
  NOR2_X1    g5453(.A1(new_n5494_), .A2(new_n5506_), .ZN(new_n5511_));
  NOR2_X1    g5454(.A1(new_n5493_), .A2(new_n5504_), .ZN(new_n5512_));
  OAI21_X1   g5455(.A1(new_n5511_), .A2(new_n5512_), .B(new_n5510_), .ZN(new_n5513_));
  NAND2_X1   g5456(.A1(new_n5509_), .A2(new_n5513_), .ZN(new_n5514_));
  NAND3_X1   g5457(.A1(new_n5405_), .A2(new_n5406_), .A3(new_n5280_), .ZN(new_n5515_));
  OAI21_X1   g5458(.A1(new_n5391_), .A2(new_n5384_), .B(new_n5267_), .ZN(new_n5516_));
  NAND2_X1   g5459(.A1(new_n5516_), .A2(new_n5275_), .ZN(new_n5517_));
  NAND3_X1   g5460(.A1(new_n5517_), .A2(new_n5403_), .A3(new_n5515_), .ZN(new_n5518_));
  XOR2_X1    g5461(.A1(new_n5380_), .A2(new_n5305_), .Z(new_n5519_));
  NOR2_X1    g5462(.A1(new_n5519_), .A2(new_n5309_), .ZN(new_n5520_));
  INV_X1     g5463(.I(new_n5520_), .ZN(new_n5521_));
  AOI21_X1   g5464(.A1(new_n5518_), .A2(new_n5521_), .B(new_n5514_), .ZN(new_n5522_));
  NOR3_X1    g5465(.A1(new_n5391_), .A2(new_n5384_), .A3(new_n5267_), .ZN(new_n5523_));
  AOI21_X1   g5466(.A1(new_n5405_), .A2(new_n5406_), .B(new_n5280_), .ZN(new_n5524_));
  NOR2_X1    g5467(.A1(new_n5524_), .A2(new_n5276_), .ZN(new_n5525_));
  NOR3_X1    g5468(.A1(new_n5525_), .A2(new_n5161_), .A3(new_n5523_), .ZN(new_n5526_));
  AOI21_X1   g5469(.A1(new_n5509_), .A2(new_n5513_), .B(new_n5520_), .ZN(new_n5527_));
  INV_X1     g5470(.I(new_n5527_), .ZN(new_n5528_));
  NOR2_X1    g5471(.A1(new_n5526_), .A2(new_n5528_), .ZN(new_n5529_));
  NOR2_X1    g5472(.A1(new_n5522_), .A2(new_n5529_), .ZN(new_n5530_));
  NOR2_X1    g5473(.A1(new_n5530_), .A2(new_n5415_), .ZN(new_n5531_));
  INV_X1     g5474(.I(new_n5531_), .ZN(new_n5532_));
  XOR2_X1    g5475(.A1(new_n5435_), .A2(new_n5532_), .Z(new_n5533_));
  XOR2_X1    g5476(.A1(new_n5533_), .A2(new_n4404_), .Z(\sin[8] ));
  XOR2_X1    g5477(.A1(new_n5440_), .A2(new_n5493_), .Z(new_n5535_));
  NAND4_X1   g5478(.A1(new_n5517_), .A2(new_n5403_), .A3(new_n5515_), .A4(new_n5535_), .ZN(new_n5536_));
  NOR2_X1    g5479(.A1(new_n5521_), .A2(new_n5506_), .ZN(new_n5537_));
  OAI21_X1   g5480(.A1(new_n5526_), .A2(new_n5535_), .B(new_n5537_), .ZN(new_n5538_));
  NAND3_X1   g5481(.A1(new_n5482_), .A2(new_n5476_), .A3(new_n5445_), .ZN(new_n5539_));
  NOR2_X1    g5482(.A1(new_n5363_), .A2(new_n5353_), .ZN(new_n5540_));
  NAND2_X1   g5483(.A1(new_n5540_), .A2(new_n5539_), .ZN(new_n5541_));
  NAND2_X1   g5484(.A1(new_n5541_), .A2(new_n5478_), .ZN(new_n5542_));
  AOI22_X1   g5485(.A1(new_n4747_), .A2(new_n4475_), .B1(new_n2977_), .B2(new_n3086_), .ZN(new_n5543_));
  OAI22_X1   g5486(.A1(new_n4243_), .A2(new_n3512_), .B1(new_n4230_), .B2(new_n3028_), .ZN(new_n5544_));
  AOI21_X1   g5487(.A1(new_n5544_), .A2(new_n721_), .B(new_n2991_), .ZN(new_n5545_));
  XNOR2_X1   g5488(.A1(new_n4800_), .A2(new_n5545_), .ZN(new_n5546_));
  INV_X1     g5489(.I(new_n5546_), .ZN(new_n5547_));
  INV_X1     g5490(.I(new_n5456_), .ZN(new_n5548_));
  OAI21_X1   g5491(.A1(new_n5450_), .A2(new_n5457_), .B(new_n5548_), .ZN(new_n5549_));
  NAND2_X1   g5492(.A1(new_n3494_), .A2(new_n4270_), .ZN(new_n5550_));
  AOI22_X1   g5493(.A1(new_n4787_), .A2(new_n5550_), .B1(new_n3398_), .B2(new_n3597_), .ZN(new_n5551_));
  OAI21_X1   g5494(.A1(new_n5551_), .A2(new_n438_), .B(new_n3393_), .ZN(new_n5552_));
  XNOR2_X1   g5495(.A1(new_n3607_), .A2(new_n5552_), .ZN(new_n5553_));
  OAI21_X1   g5496(.A1(new_n3568_), .A2(new_n3569_), .B(new_n437_), .ZN(new_n5554_));
  XOR2_X1    g5497(.A1(new_n5553_), .A2(new_n5554_), .Z(new_n5555_));
  XOR2_X1    g5498(.A1(new_n5555_), .A2(new_n5549_), .Z(new_n5556_));
  NAND2_X1   g5499(.A1(new_n5556_), .A2(new_n5547_), .ZN(new_n5557_));
  INV_X1     g5500(.I(new_n5549_), .ZN(new_n5558_));
  INV_X1     g5501(.I(new_n5555_), .ZN(new_n5559_));
  NOR2_X1    g5502(.A1(new_n5559_), .A2(new_n5558_), .ZN(new_n5560_));
  NOR2_X1    g5503(.A1(new_n5555_), .A2(new_n5549_), .ZN(new_n5561_));
  OAI21_X1   g5504(.A1(new_n5560_), .A2(new_n5561_), .B(new_n5546_), .ZN(new_n5562_));
  NAND2_X1   g5505(.A1(new_n5557_), .A2(new_n5562_), .ZN(new_n5563_));
  NOR2_X1    g5506(.A1(new_n5462_), .A2(new_n5464_), .ZN(new_n5564_));
  NAND2_X1   g5507(.A1(new_n5462_), .A2(new_n5464_), .ZN(new_n5565_));
  XOR2_X1    g5508(.A1(new_n5468_), .A2(new_n702_), .Z(new_n5566_));
  AOI21_X1   g5509(.A1(new_n5566_), .A2(new_n5565_), .B(new_n5564_), .ZN(new_n5567_));
  NOR2_X1    g5510(.A1(new_n5563_), .A2(new_n5567_), .ZN(new_n5568_));
  NAND2_X1   g5511(.A1(new_n5563_), .A2(new_n5567_), .ZN(new_n5569_));
  INV_X1     g5512(.I(new_n5569_), .ZN(new_n5570_));
  OAI21_X1   g5513(.A1(new_n5570_), .A2(new_n5568_), .B(new_n5543_), .ZN(new_n5571_));
  INV_X1     g5514(.I(new_n5543_), .ZN(new_n5572_));
  INV_X1     g5515(.I(new_n5568_), .ZN(new_n5573_));
  NAND3_X1   g5516(.A1(new_n5573_), .A2(new_n5572_), .A3(new_n5569_), .ZN(new_n5574_));
  AOI21_X1   g5517(.A1(new_n5571_), .A2(new_n5574_), .B(new_n803_), .ZN(new_n5575_));
  AOI21_X1   g5518(.A1(new_n5573_), .A2(new_n5569_), .B(new_n5572_), .ZN(new_n5576_));
  NOR3_X1    g5519(.A1(new_n5570_), .A2(new_n5543_), .A3(new_n5568_), .ZN(new_n5577_));
  NOR3_X1    g5520(.A1(new_n5576_), .A2(new_n5577_), .A3(new_n802_), .ZN(new_n5578_));
  NOR3_X1    g5521(.A1(new_n5542_), .A2(new_n5575_), .A3(new_n5578_), .ZN(new_n5579_));
  OAI21_X1   g5522(.A1(new_n5576_), .A2(new_n5577_), .B(new_n802_), .ZN(new_n5580_));
  NAND3_X1   g5523(.A1(new_n5571_), .A2(new_n5574_), .A3(new_n803_), .ZN(new_n5581_));
  AOI22_X1   g5524(.A1(new_n5580_), .A2(new_n5581_), .B1(new_n5478_), .B2(new_n5541_), .ZN(new_n5582_));
  NOR2_X1    g5525(.A1(new_n5582_), .A2(new_n5579_), .ZN(new_n5583_));
  NOR2_X1    g5526(.A1(new_n5365_), .A2(new_n5316_), .ZN(new_n5584_));
  NOR2_X1    g5527(.A1(new_n5584_), .A2(new_n5360_), .ZN(new_n5585_));
  XOR2_X1    g5528(.A1(new_n5489_), .A2(new_n5585_), .Z(new_n5586_));
  NOR3_X1    g5529(.A1(new_n5586_), .A2(new_n5492_), .A3(new_n5583_), .ZN(new_n5587_));
  INV_X1     g5530(.I(new_n5489_), .ZN(new_n5588_));
  NOR2_X1    g5531(.A1(new_n5588_), .A2(new_n5585_), .ZN(new_n5589_));
  NOR2_X1    g5532(.A1(new_n5587_), .A2(new_n5589_), .ZN(new_n5590_));
  NOR2_X1    g5533(.A1(new_n5590_), .A2(new_n5440_), .ZN(new_n5591_));
  OR2_X2     g5534(.A1(new_n5582_), .A2(new_n5579_), .Z(new_n5592_));
  NAND3_X1   g5535(.A1(new_n5442_), .A2(new_n5485_), .A3(new_n5488_), .ZN(new_n5593_));
  NAND2_X1   g5536(.A1(new_n5489_), .A2(new_n5585_), .ZN(new_n5594_));
  NAND2_X1   g5537(.A1(new_n5593_), .A2(new_n5594_), .ZN(new_n5595_));
  NAND3_X1   g5538(.A1(new_n5595_), .A2(new_n5491_), .A3(new_n5592_), .ZN(new_n5596_));
  INV_X1     g5539(.I(new_n5589_), .ZN(new_n5597_));
  NAND2_X1   g5540(.A1(new_n5596_), .A2(new_n5597_), .ZN(new_n5598_));
  NOR2_X1    g5541(.A1(new_n5510_), .A2(new_n5598_), .ZN(new_n5599_));
  NOR2_X1    g5542(.A1(new_n5591_), .A2(new_n5599_), .ZN(new_n5600_));
  NOR4_X1    g5543(.A1(new_n151_), .A2(new_n367_), .A3(new_n221_), .A4(new_n456_), .ZN(new_n5601_));
  NOR3_X1    g5544(.A1(new_n2347_), .A2(new_n3968_), .A3(new_n1088_), .ZN(new_n5602_));
  NAND2_X1   g5545(.A1(new_n5602_), .A2(new_n5601_), .ZN(new_n5603_));
  NOR3_X1    g5546(.A1(new_n5603_), .A2(new_n606_), .A3(new_n2911_), .ZN(new_n5604_));
  NAND3_X1   g5547(.A1(new_n2447_), .A2(new_n4068_), .A3(new_n5604_), .ZN(new_n5605_));
  NAND2_X1   g5548(.A1(new_n5600_), .A2(new_n5605_), .ZN(new_n5606_));
  NAND2_X1   g5549(.A1(new_n5510_), .A2(new_n5598_), .ZN(new_n5607_));
  NAND2_X1   g5550(.A1(new_n5590_), .A2(new_n5440_), .ZN(new_n5608_));
  NAND2_X1   g5551(.A1(new_n5608_), .A2(new_n5607_), .ZN(new_n5609_));
  INV_X1     g5552(.I(new_n5605_), .ZN(new_n5610_));
  NAND2_X1   g5553(.A1(new_n5609_), .A2(new_n5610_), .ZN(new_n5611_));
  NAND2_X1   g5554(.A1(new_n5606_), .A2(new_n5611_), .ZN(new_n5612_));
  INV_X1     g5555(.I(new_n5612_), .ZN(new_n5613_));
  NAND3_X1   g5556(.A1(new_n5538_), .A2(new_n5536_), .A3(new_n5613_), .ZN(new_n5614_));
  INV_X1     g5557(.I(new_n5536_), .ZN(new_n5615_));
  INV_X1     g5558(.I(new_n5535_), .ZN(new_n5616_));
  INV_X1     g5559(.I(new_n5537_), .ZN(new_n5617_));
  AOI21_X1   g5560(.A1(new_n5518_), .A2(new_n5616_), .B(new_n5617_), .ZN(new_n5618_));
  OAI21_X1   g5561(.A1(new_n5618_), .A2(new_n5615_), .B(new_n5612_), .ZN(new_n5619_));
  NAND2_X1   g5562(.A1(new_n5619_), .A2(new_n5614_), .ZN(new_n5620_));
  XNOR2_X1   g5563(.A1(new_n5620_), .A2(new_n5531_), .ZN(new_n5621_));
  NAND2_X1   g5564(.A1(new_n5530_), .A2(new_n5415_), .ZN(new_n5622_));
  NAND2_X1   g5565(.A1(new_n5532_), .A2(new_n5622_), .ZN(new_n5623_));
  NAND2_X1   g5566(.A1(new_n5435_), .A2(new_n5623_), .ZN(new_n5624_));
  NAND2_X1   g5567(.A1(new_n5624_), .A2(new_n4404_), .ZN(new_n5625_));
  XOR2_X1    g5568(.A1(new_n5625_), .A2(new_n5621_), .Z(\sin[9] ));
  INV_X1     g5569(.I(new_n5621_), .ZN(new_n5627_));
  OAI21_X1   g5570(.A1(new_n5624_), .A2(new_n5627_), .B(new_n4404_), .ZN(new_n5628_));
  AOI21_X1   g5571(.A1(new_n5538_), .A2(new_n5536_), .B(new_n5613_), .ZN(new_n5629_));
  INV_X1     g5572(.I(new_n5514_), .ZN(new_n5630_));
  OAI21_X1   g5573(.A1(new_n5526_), .A2(new_n5520_), .B(new_n5630_), .ZN(new_n5631_));
  OAI21_X1   g5574(.A1(new_n5524_), .A2(new_n5276_), .B(new_n5515_), .ZN(new_n5632_));
  OAI21_X1   g5575(.A1(new_n5632_), .A2(new_n5161_), .B(new_n5527_), .ZN(new_n5633_));
  AOI22_X1   g5576(.A1(new_n5631_), .A2(new_n5633_), .B1(new_n5414_), .B2(new_n5302_), .ZN(new_n5634_));
  NOR4_X1    g5577(.A1(new_n5422_), .A2(new_n5522_), .A3(new_n5529_), .A4(new_n5419_), .ZN(new_n5635_));
  OAI21_X1   g5578(.A1(new_n5635_), .A2(new_n5634_), .B(new_n5629_), .ZN(new_n5636_));
  AOI21_X1   g5579(.A1(new_n5275_), .A2(new_n5516_), .B(new_n5523_), .ZN(new_n5637_));
  AOI21_X1   g5580(.A1(new_n5637_), .A2(new_n5403_), .B(new_n5535_), .ZN(new_n5638_));
  OAI21_X1   g5581(.A1(new_n5638_), .A2(new_n5617_), .B(new_n5536_), .ZN(new_n5639_));
  NOR2_X1    g5582(.A1(new_n5600_), .A2(new_n5605_), .ZN(new_n5640_));
  NOR2_X1    g5583(.A1(new_n5592_), .A2(new_n5489_), .ZN(new_n5641_));
  INV_X1     g5584(.I(new_n5641_), .ZN(new_n5642_));
  NAND2_X1   g5585(.A1(new_n5592_), .A2(new_n5489_), .ZN(new_n5643_));
  NAND2_X1   g5586(.A1(new_n5643_), .A2(new_n5585_), .ZN(new_n5644_));
  NAND2_X1   g5587(.A1(new_n5644_), .A2(new_n5642_), .ZN(new_n5645_));
  INV_X1     g5588(.I(new_n5563_), .ZN(new_n5646_));
  NOR2_X1    g5589(.A1(new_n5646_), .A2(new_n5567_), .ZN(new_n5647_));
  NAND2_X1   g5590(.A1(new_n5646_), .A2(new_n5567_), .ZN(new_n5648_));
  XOR2_X1    g5591(.A1(new_n5543_), .A2(new_n802_), .Z(new_n5649_));
  AOI21_X1   g5592(.A1(new_n5648_), .A2(new_n5649_), .B(new_n5647_), .ZN(new_n5650_));
  XOR2_X1    g5593(.A1(new_n2879_), .A2(new_n438_), .Z(new_n5651_));
  NAND2_X1   g5594(.A1(new_n5553_), .A2(new_n5651_), .ZN(new_n5652_));
  MUX2_X1    g5595(.I0(new_n3436_), .I1(new_n438_), .S(new_n5652_), .Z(new_n5653_));
  NOR2_X1    g5596(.A1(new_n2898_), .A2(new_n438_), .ZN(new_n5654_));
  INV_X1     g5597(.I(new_n5654_), .ZN(new_n5655_));
  XOR2_X1    g5598(.A1(new_n5454_), .A2(new_n802_), .Z(new_n5656_));
  NOR2_X1    g5599(.A1(new_n5455_), .A2(new_n802_), .ZN(new_n5657_));
  NOR2_X1    g5600(.A1(new_n5454_), .A2(new_n803_), .ZN(new_n5658_));
  OAI21_X1   g5601(.A1(new_n5657_), .A2(new_n5658_), .B(new_n5655_), .ZN(new_n5659_));
  OAI21_X1   g5602(.A1(new_n5655_), .A2(new_n5656_), .B(new_n5659_), .ZN(new_n5660_));
  NOR2_X1    g5603(.A1(new_n5653_), .A2(new_n5660_), .ZN(new_n5661_));
  INV_X1     g5604(.I(new_n5661_), .ZN(new_n5662_));
  NAND2_X1   g5605(.A1(new_n5653_), .A2(new_n5660_), .ZN(new_n5663_));
  NAND2_X1   g5606(.A1(new_n5662_), .A2(new_n5663_), .ZN(new_n5664_));
  AOI22_X1   g5607(.A1(new_n2946_), .A2(new_n4270_), .B1(new_n3985_), .B2(new_n3494_), .ZN(new_n5665_));
  NOR2_X1    g5608(.A1(new_n3987_), .A2(new_n3496_), .ZN(new_n5666_));
  OAI21_X1   g5609(.A1(new_n5666_), .A2(new_n5665_), .B(new_n437_), .ZN(new_n5667_));
  NAND2_X1   g5610(.A1(new_n5667_), .A2(new_n3393_), .ZN(new_n5668_));
  XOR2_X1    g5611(.A1(new_n3982_), .A2(new_n5668_), .Z(new_n5669_));
  XOR2_X1    g5612(.A1(new_n5664_), .A2(new_n5669_), .Z(new_n5670_));
  NAND2_X1   g5613(.A1(new_n5555_), .A2(new_n5549_), .ZN(new_n5671_));
  OAI21_X1   g5614(.A1(new_n5547_), .A2(new_n5561_), .B(new_n5671_), .ZN(new_n5672_));
  OAI22_X1   g5615(.A1(new_n4230_), .A2(new_n3031_), .B1(new_n4182_), .B2(new_n2994_), .ZN(new_n5673_));
  OAI21_X1   g5616(.A1(new_n3028_), .A2(new_n4474_), .B(new_n5673_), .ZN(new_n5674_));
  AOI21_X1   g5617(.A1(new_n5674_), .A2(new_n721_), .B(new_n2991_), .ZN(new_n5675_));
  XOR2_X1    g5618(.A1(new_n4484_), .A2(new_n5675_), .Z(new_n5676_));
  XOR2_X1    g5619(.A1(new_n5672_), .A2(new_n5676_), .Z(new_n5677_));
  OR2_X2     g5620(.A1(new_n5672_), .A2(new_n5676_), .Z(new_n5678_));
  NAND2_X1   g5621(.A1(new_n5672_), .A2(new_n5676_), .ZN(new_n5679_));
  AOI21_X1   g5622(.A1(new_n5678_), .A2(new_n5679_), .B(new_n5670_), .ZN(new_n5680_));
  AOI21_X1   g5623(.A1(new_n5670_), .A2(new_n5677_), .B(new_n5680_), .ZN(new_n5681_));
  NAND2_X1   g5624(.A1(new_n5681_), .A2(new_n5650_), .ZN(new_n5682_));
  OR2_X2     g5625(.A1(new_n5681_), .A2(new_n5650_), .Z(new_n5683_));
  NAND2_X1   g5626(.A1(new_n5683_), .A2(new_n5682_), .ZN(new_n5684_));
  INV_X1     g5627(.I(new_n2619_), .ZN(new_n5685_));
  NOR4_X1    g5628(.A1(new_n2854_), .A2(new_n201_), .A3(new_n345_), .A4(new_n1001_), .ZN(new_n5686_));
  NOR4_X1    g5629(.A1(new_n3968_), .A2(new_n425_), .A3(new_n624_), .A4(new_n852_), .ZN(new_n5687_));
  AND3_X2    g5630(.A1(new_n5686_), .A2(new_n2920_), .A3(new_n5687_), .Z(new_n5688_));
  AND4_X2    g5631(.A1(new_n667_), .A2(new_n5688_), .A3(new_n5685_), .A4(new_n4047_), .Z(new_n5689_));
  NAND2_X1   g5632(.A1(new_n5684_), .A2(new_n5689_), .ZN(new_n5690_));
  INV_X1     g5633(.I(new_n5690_), .ZN(new_n5691_));
  OAI21_X1   g5634(.A1(new_n5510_), .A2(new_n5645_), .B(new_n5691_), .ZN(new_n5692_));
  AOI21_X1   g5635(.A1(new_n5585_), .A2(new_n5643_), .B(new_n5641_), .ZN(new_n5693_));
  NAND3_X1   g5636(.A1(new_n5440_), .A2(new_n5693_), .A3(new_n5690_), .ZN(new_n5694_));
  AOI21_X1   g5637(.A1(new_n5692_), .A2(new_n5694_), .B(new_n5579_), .ZN(new_n5695_));
  INV_X1     g5638(.I(new_n5579_), .ZN(new_n5696_));
  AOI21_X1   g5639(.A1(new_n5440_), .A2(new_n5693_), .B(new_n5690_), .ZN(new_n5697_));
  NOR3_X1    g5640(.A1(new_n5510_), .A2(new_n5645_), .A3(new_n5691_), .ZN(new_n5698_));
  NOR3_X1    g5641(.A1(new_n5698_), .A2(new_n5697_), .A3(new_n5696_), .ZN(new_n5699_));
  NOR2_X1    g5642(.A1(new_n5695_), .A2(new_n5699_), .ZN(new_n5700_));
  AOI21_X1   g5643(.A1(new_n5608_), .A2(new_n5607_), .B(new_n5610_), .ZN(new_n5701_));
  NOR3_X1    g5644(.A1(new_n5591_), .A2(new_n5599_), .A3(new_n5605_), .ZN(new_n5702_));
  NOR2_X1    g5645(.A1(new_n5701_), .A2(new_n5702_), .ZN(new_n5703_));
  NOR3_X1    g5646(.A1(new_n5700_), .A2(new_n5703_), .A3(new_n5640_), .ZN(new_n5704_));
  NOR2_X1    g5647(.A1(new_n5600_), .A2(new_n5605_), .ZN(new_n5705_));
  NOR2_X1    g5648(.A1(new_n5704_), .A2(new_n5705_), .ZN(new_n5706_));
  NOR2_X1    g5649(.A1(new_n5639_), .A2(new_n5706_), .ZN(new_n5707_));
  OAI21_X1   g5650(.A1(new_n5698_), .A2(new_n5697_), .B(new_n5696_), .ZN(new_n5708_));
  NAND3_X1   g5651(.A1(new_n5692_), .A2(new_n5694_), .A3(new_n5579_), .ZN(new_n5709_));
  NAND2_X1   g5652(.A1(new_n5708_), .A2(new_n5709_), .ZN(new_n5710_));
  OAI21_X1   g5653(.A1(new_n5591_), .A2(new_n5599_), .B(new_n5605_), .ZN(new_n5711_));
  NAND3_X1   g5654(.A1(new_n5608_), .A2(new_n5607_), .A3(new_n5610_), .ZN(new_n5712_));
  NAND2_X1   g5655(.A1(new_n5711_), .A2(new_n5712_), .ZN(new_n5713_));
  NAND3_X1   g5656(.A1(new_n5710_), .A2(new_n5713_), .A3(new_n5611_), .ZN(new_n5714_));
  INV_X1     g5657(.I(new_n5705_), .ZN(new_n5715_));
  NAND2_X1   g5658(.A1(new_n5714_), .A2(new_n5715_), .ZN(new_n5716_));
  AOI21_X1   g5659(.A1(new_n5536_), .A2(new_n5538_), .B(new_n5716_), .ZN(new_n5717_));
  NOR2_X1    g5660(.A1(new_n5717_), .A2(new_n5707_), .ZN(new_n5718_));
  NOR2_X1    g5661(.A1(new_n5636_), .A2(new_n5718_), .ZN(new_n5719_));
  OAI22_X1   g5662(.A1(new_n5522_), .A2(new_n5529_), .B1(new_n5422_), .B2(new_n5419_), .ZN(new_n5720_));
  NAND4_X1   g5663(.A1(new_n5631_), .A2(new_n5414_), .A3(new_n5302_), .A4(new_n5633_), .ZN(new_n5721_));
  AOI21_X1   g5664(.A1(new_n5720_), .A2(new_n5721_), .B(new_n5619_), .ZN(new_n5722_));
  NAND3_X1   g5665(.A1(new_n5716_), .A2(new_n5538_), .A3(new_n5536_), .ZN(new_n5723_));
  NAND2_X1   g5666(.A1(new_n5639_), .A2(new_n5706_), .ZN(new_n5724_));
  NAND2_X1   g5667(.A1(new_n5724_), .A2(new_n5723_), .ZN(new_n5725_));
  NOR2_X1    g5668(.A1(new_n5722_), .A2(new_n5725_), .ZN(new_n5726_));
  NOR2_X1    g5669(.A1(new_n5719_), .A2(new_n5726_), .ZN(new_n5727_));
  XOR2_X1    g5670(.A1(new_n5722_), .A2(new_n5725_), .Z(new_n5728_));
  NAND2_X1   g5671(.A1(new_n5628_), .A2(new_n5728_), .ZN(new_n5729_));
  OAI21_X1   g5672(.A1(new_n5628_), .A2(new_n5727_), .B(new_n5729_), .ZN(\sin[10] ));
  INV_X1     g5673(.I(new_n5620_), .ZN(new_n5731_));
  NAND3_X1   g5674(.A1(new_n5435_), .A2(new_n5731_), .A3(new_n5623_), .ZN(new_n5732_));
  NOR2_X1    g5675(.A1(new_n5295_), .A2(new_n5285_), .ZN(new_n5733_));
  AOI21_X1   g5676(.A1(new_n5429_), .A2(new_n5294_), .B(new_n5428_), .ZN(new_n5734_));
  INV_X1     g5677(.I(new_n5434_), .ZN(new_n5735_));
  OAI21_X1   g5678(.A1(new_n5734_), .A2(new_n5733_), .B(new_n5735_), .ZN(new_n5736_));
  INV_X1     g5679(.I(new_n5623_), .ZN(new_n5737_));
  OAI21_X1   g5680(.A1(new_n5736_), .A2(new_n5737_), .B(new_n5620_), .ZN(new_n5738_));
  NOR2_X1    g5681(.A1(new_n5718_), .A2(new_n5620_), .ZN(new_n5739_));
  NAND2_X1   g5682(.A1(new_n5718_), .A2(new_n5620_), .ZN(new_n5740_));
  INV_X1     g5683(.I(new_n5740_), .ZN(new_n5741_));
  OAI21_X1   g5684(.A1(new_n5741_), .A2(new_n5739_), .B(new_n5531_), .ZN(new_n5742_));
  AOI21_X1   g5685(.A1(new_n5738_), .A2(new_n5732_), .B(new_n5742_), .ZN(new_n5743_));
  INV_X1     g5686(.I(new_n5683_), .ZN(new_n5744_));
  NAND2_X1   g5687(.A1(new_n5579_), .A2(new_n5682_), .ZN(new_n5745_));
  NOR3_X1    g5688(.A1(new_n5510_), .A2(new_n5645_), .A3(new_n5745_), .ZN(new_n5746_));
  NOR2_X1    g5689(.A1(new_n5746_), .A2(new_n5744_), .ZN(new_n5747_));
  NAND2_X1   g5690(.A1(new_n5670_), .A2(new_n5678_), .ZN(new_n5748_));
  NAND2_X1   g5691(.A1(new_n5748_), .A2(new_n5679_), .ZN(new_n5749_));
  INV_X1     g5692(.I(new_n5749_), .ZN(new_n5750_));
  INV_X1     g5693(.I(new_n5669_), .ZN(new_n5751_));
  NOR2_X1    g5694(.A1(new_n5664_), .A2(new_n5751_), .ZN(new_n5752_));
  NAND2_X1   g5695(.A1(new_n4475_), .A2(new_n3030_), .ZN(new_n5753_));
  AOI21_X1   g5696(.A1(new_n4232_), .A2(new_n3038_), .B(new_n702_), .ZN(new_n5754_));
  AOI21_X1   g5697(.A1(new_n5753_), .A2(new_n5754_), .B(new_n2991_), .ZN(new_n5755_));
  XNOR2_X1   g5698(.A1(new_n4688_), .A2(new_n5755_), .ZN(new_n5756_));
  INV_X1     g5699(.I(new_n5756_), .ZN(new_n5757_));
  OAI22_X1   g5700(.A1(new_n3987_), .A2(new_n3493_), .B1(new_n3396_), .B2(new_n3597_), .ZN(new_n5758_));
  OAI21_X1   g5701(.A1(new_n3496_), .A2(new_n4192_), .B(new_n5758_), .ZN(new_n5759_));
  AOI21_X1   g5702(.A1(new_n5759_), .A2(new_n437_), .B(new_n3501_), .ZN(new_n5760_));
  XNOR2_X1   g5703(.A1(new_n4198_), .A2(new_n5760_), .ZN(new_n5761_));
  NOR2_X1    g5704(.A1(new_n5654_), .A2(new_n5657_), .ZN(new_n5762_));
  NOR2_X1    g5705(.A1(new_n5762_), .A2(new_n5658_), .ZN(new_n5763_));
  NOR2_X1    g5706(.A1(new_n2926_), .A2(new_n438_), .ZN(new_n5764_));
  INV_X1     g5707(.I(new_n5764_), .ZN(new_n5765_));
  NOR2_X1    g5708(.A1(new_n5763_), .A2(new_n5765_), .ZN(new_n5766_));
  NOR3_X1    g5709(.A1(new_n5762_), .A2(new_n5658_), .A3(new_n5764_), .ZN(new_n5767_));
  OAI21_X1   g5710(.A1(new_n5766_), .A2(new_n5767_), .B(new_n5761_), .ZN(new_n5768_));
  XOR2_X1    g5711(.A1(new_n5763_), .A2(new_n5764_), .Z(new_n5769_));
  OAI21_X1   g5712(.A1(new_n5761_), .A2(new_n5769_), .B(new_n5768_), .ZN(new_n5770_));
  NAND2_X1   g5713(.A1(new_n5757_), .A2(new_n5770_), .ZN(new_n5771_));
  XOR2_X1    g5714(.A1(new_n5771_), .A2(new_n5752_), .Z(new_n5772_));
  XOR2_X1    g5715(.A1(new_n5772_), .A2(new_n5661_), .Z(new_n5773_));
  XOR2_X1    g5716(.A1(new_n5773_), .A2(new_n5750_), .Z(new_n5774_));
  NOR3_X1    g5717(.A1(new_n3965_), .A2(new_n201_), .A3(new_n479_), .ZN(new_n5775_));
  NOR2_X1    g5718(.A1(new_n527_), .A2(new_n749_), .ZN(new_n5776_));
  NAND4_X1   g5719(.A1(new_n663_), .A2(new_n4228_), .A3(new_n5775_), .A4(new_n5776_), .ZN(new_n5777_));
  XOR2_X1    g5720(.A1(new_n5774_), .A2(new_n5777_), .Z(new_n5778_));
  NOR2_X1    g5721(.A1(new_n5747_), .A2(new_n5778_), .ZN(new_n5779_));
  XNOR2_X1   g5722(.A1(new_n5774_), .A2(new_n5777_), .ZN(new_n5780_));
  INV_X1     g5723(.I(new_n5780_), .ZN(new_n5781_));
  AOI21_X1   g5724(.A1(new_n5747_), .A2(new_n5781_), .B(new_n5779_), .ZN(new_n5782_));
  NAND3_X1   g5725(.A1(new_n5708_), .A2(new_n5709_), .A3(new_n5600_), .ZN(new_n5783_));
  AOI21_X1   g5726(.A1(new_n5708_), .A2(new_n5709_), .B(new_n5600_), .ZN(new_n5784_));
  OAI21_X1   g5727(.A1(new_n5784_), .A2(new_n5610_), .B(new_n5783_), .ZN(new_n5785_));
  AOI21_X1   g5728(.A1(new_n5538_), .A2(new_n5536_), .B(new_n5785_), .ZN(new_n5786_));
  NOR2_X1    g5729(.A1(new_n5510_), .A2(new_n5645_), .ZN(new_n5787_));
  XOR2_X1    g5730(.A1(new_n5690_), .A2(new_n5696_), .Z(new_n5788_));
  NAND2_X1   g5731(.A1(new_n5787_), .A2(new_n5788_), .ZN(new_n5789_));
  INV_X1     g5732(.I(new_n5789_), .ZN(new_n5790_));
  OAI21_X1   g5733(.A1(new_n5786_), .A2(new_n5790_), .B(new_n5782_), .ZN(new_n5791_));
  INV_X1     g5734(.I(new_n5782_), .ZN(new_n5792_));
  NOR3_X1    g5735(.A1(new_n5695_), .A2(new_n5699_), .A3(new_n5609_), .ZN(new_n5793_));
  OAI21_X1   g5736(.A1(new_n5695_), .A2(new_n5699_), .B(new_n5609_), .ZN(new_n5794_));
  AOI21_X1   g5737(.A1(new_n5605_), .A2(new_n5794_), .B(new_n5793_), .ZN(new_n5795_));
  OAI21_X1   g5738(.A1(new_n5618_), .A2(new_n5615_), .B(new_n5795_), .ZN(new_n5796_));
  NAND3_X1   g5739(.A1(new_n5796_), .A2(new_n5792_), .A3(new_n5789_), .ZN(new_n5797_));
  NAND2_X1   g5740(.A1(new_n5791_), .A2(new_n5797_), .ZN(new_n5798_));
  NAND2_X1   g5741(.A1(new_n5719_), .A2(new_n5798_), .ZN(new_n5799_));
  XOR2_X1    g5742(.A1(new_n5743_), .A2(new_n5799_), .Z(new_n5800_));
  XOR2_X1    g5743(.A1(new_n5800_), .A2(new_n4404_), .Z(\sin[11] ));
  AOI21_X1   g5744(.A1(new_n5796_), .A2(new_n5789_), .B(new_n5792_), .ZN(new_n5802_));
  NOR3_X1    g5745(.A1(new_n5786_), .A2(new_n5782_), .A3(new_n5790_), .ZN(new_n5803_));
  NOR2_X1    g5746(.A1(new_n5802_), .A2(new_n5803_), .ZN(new_n5804_));
  XOR2_X1    g5747(.A1(new_n5747_), .A2(new_n5774_), .Z(new_n5805_));
  NOR2_X1    g5748(.A1(new_n5796_), .A2(new_n5805_), .ZN(new_n5806_));
  NAND2_X1   g5749(.A1(new_n5796_), .A2(new_n5805_), .ZN(new_n5807_));
  NOR2_X1    g5750(.A1(new_n5789_), .A2(new_n5777_), .ZN(new_n5808_));
  AOI21_X1   g5751(.A1(new_n5807_), .A2(new_n5808_), .B(new_n5806_), .ZN(new_n5809_));
  NOR2_X1    g5752(.A1(new_n5773_), .A2(new_n5750_), .ZN(new_n5810_));
  NOR3_X1    g5753(.A1(new_n5664_), .A2(new_n5662_), .A3(new_n5751_), .ZN(new_n5811_));
  OAI21_X1   g5754(.A1(new_n5757_), .A2(new_n5770_), .B(new_n5811_), .ZN(new_n5812_));
  NAND2_X1   g5755(.A1(new_n5812_), .A2(new_n5771_), .ZN(new_n5813_));
  NOR2_X1    g5756(.A1(new_n5761_), .A2(new_n5767_), .ZN(new_n5814_));
  NOR2_X1    g5757(.A1(new_n5814_), .A2(new_n5766_), .ZN(new_n5815_));
  NOR3_X1    g5758(.A1(new_n2946_), .A2(new_n3985_), .A3(new_n438_), .ZN(new_n5816_));
  INV_X1     g5759(.I(new_n5816_), .ZN(new_n5817_));
  NOR2_X1    g5760(.A1(new_n3985_), .A2(new_n438_), .ZN(new_n5818_));
  NOR2_X1    g5761(.A1(new_n5765_), .A2(new_n5818_), .ZN(new_n5819_));
  INV_X1     g5762(.I(new_n5819_), .ZN(new_n5820_));
  AOI21_X1   g5763(.A1(new_n5817_), .A2(new_n5820_), .B(new_n5815_), .ZN(new_n5821_));
  INV_X1     g5764(.I(new_n5815_), .ZN(new_n5822_));
  XOR2_X1    g5765(.A1(new_n5818_), .A2(new_n5764_), .Z(new_n5823_));
  NOR2_X1    g5766(.A1(new_n5822_), .A2(new_n5823_), .ZN(new_n5824_));
  NOR2_X1    g5767(.A1(new_n5824_), .A2(new_n5821_), .ZN(new_n5825_));
  INV_X1     g5768(.I(new_n4747_), .ZN(new_n5826_));
  OAI22_X1   g5769(.A1(new_n5826_), .A2(new_n3031_), .B1(new_n2991_), .B2(new_n4474_), .ZN(new_n5827_));
  OAI22_X1   g5770(.A1(new_n4182_), .A2(new_n3493_), .B1(new_n3987_), .B2(new_n3396_), .ZN(new_n5828_));
  OAI21_X1   g5771(.A1(new_n3496_), .A2(new_n4230_), .B(new_n5828_), .ZN(new_n5829_));
  AOI21_X1   g5772(.A1(new_n5829_), .A2(new_n437_), .B(new_n3501_), .ZN(new_n5830_));
  XOR2_X1    g5773(.A1(new_n4800_), .A2(new_n5830_), .Z(new_n5831_));
  XOR2_X1    g5774(.A1(new_n5827_), .A2(new_n5831_), .Z(new_n5832_));
  XOR2_X1    g5775(.A1(new_n5825_), .A2(new_n5832_), .Z(new_n5833_));
  XOR2_X1    g5776(.A1(new_n5833_), .A2(new_n702_), .Z(new_n5834_));
  XOR2_X1    g5777(.A1(new_n5834_), .A2(new_n5813_), .Z(new_n5835_));
  XOR2_X1    g5778(.A1(new_n5773_), .A2(new_n5749_), .Z(new_n5836_));
  NOR2_X1    g5779(.A1(new_n5835_), .A2(new_n5836_), .ZN(new_n5837_));
  XNOR2_X1   g5780(.A1(new_n5837_), .A2(new_n5810_), .ZN(new_n5838_));
  INV_X1     g5781(.I(new_n5838_), .ZN(new_n5839_));
  NAND2_X1   g5782(.A1(new_n5839_), .A2(new_n5747_), .ZN(new_n5840_));
  OAI21_X1   g5783(.A1(new_n5744_), .A2(new_n5746_), .B(new_n5838_), .ZN(new_n5841_));
  NAND2_X1   g5784(.A1(new_n5840_), .A2(new_n5841_), .ZN(new_n5842_));
  INV_X1     g5785(.I(new_n5842_), .ZN(new_n5843_));
  NOR4_X1    g5786(.A1(new_n821_), .A2(new_n156_), .A3(new_n233_), .A4(new_n420_), .ZN(new_n5844_));
  NOR4_X1    g5787(.A1(new_n1004_), .A2(new_n213_), .A3(new_n416_), .A4(new_n311_), .ZN(new_n5845_));
  NAND4_X1   g5788(.A1(new_n4708_), .A2(new_n2340_), .A3(new_n5844_), .A4(new_n5845_), .ZN(new_n5846_));
  NOR3_X1    g5789(.A1(new_n2572_), .A2(new_n2336_), .A3(new_n5846_), .ZN(new_n5847_));
  INV_X1     g5790(.I(new_n5847_), .ZN(new_n5848_));
  NAND2_X1   g5791(.A1(new_n5843_), .A2(new_n5848_), .ZN(new_n5849_));
  NAND2_X1   g5792(.A1(new_n5842_), .A2(new_n5847_), .ZN(new_n5850_));
  AND2_X2    g5793(.A1(new_n5849_), .A2(new_n5850_), .Z(new_n5851_));
  NOR3_X1    g5794(.A1(new_n5719_), .A2(new_n5809_), .A3(new_n5851_), .ZN(new_n5852_));
  NAND2_X1   g5795(.A1(new_n5722_), .A2(new_n5725_), .ZN(new_n5853_));
  INV_X1     g5796(.I(new_n5805_), .ZN(new_n5854_));
  NAND2_X1   g5797(.A1(new_n5786_), .A2(new_n5854_), .ZN(new_n5855_));
  OAI21_X1   g5798(.A1(new_n5786_), .A2(new_n5854_), .B(new_n5808_), .ZN(new_n5856_));
  AOI22_X1   g5799(.A1(new_n5856_), .A2(new_n5855_), .B1(new_n5849_), .B2(new_n5850_), .ZN(new_n5857_));
  NOR2_X1    g5800(.A1(new_n5857_), .A2(new_n5853_), .ZN(new_n5858_));
  OAI21_X1   g5801(.A1(new_n5852_), .A2(new_n5858_), .B(new_n5804_), .ZN(new_n5859_));
  INV_X1     g5802(.I(new_n5859_), .ZN(new_n5860_));
  NOR3_X1    g5803(.A1(new_n5852_), .A2(new_n5858_), .A3(new_n5804_), .ZN(new_n5861_));
  NOR2_X1    g5804(.A1(new_n5860_), .A2(new_n5861_), .ZN(new_n5862_));
  NOR3_X1    g5805(.A1(new_n5736_), .A2(new_n5620_), .A3(new_n5737_), .ZN(new_n5863_));
  AOI21_X1   g5806(.A1(new_n5435_), .A2(new_n5623_), .B(new_n5731_), .ZN(new_n5864_));
  INV_X1     g5807(.I(new_n5739_), .ZN(new_n5865_));
  AOI21_X1   g5808(.A1(new_n5865_), .A2(new_n5740_), .B(new_n5532_), .ZN(new_n5866_));
  OAI21_X1   g5809(.A1(new_n5863_), .A2(new_n5864_), .B(new_n5866_), .ZN(new_n5867_));
  NAND2_X1   g5810(.A1(new_n5853_), .A2(new_n5804_), .ZN(new_n5868_));
  NAND2_X1   g5811(.A1(new_n5799_), .A2(new_n5868_), .ZN(new_n5869_));
  INV_X1     g5812(.I(new_n5869_), .ZN(new_n5870_));
  OAI21_X1   g5813(.A1(new_n5867_), .A2(new_n5870_), .B(new_n4404_), .ZN(new_n5871_));
  XOR2_X1    g5814(.A1(new_n5871_), .A2(new_n5862_), .Z(\sin[12] ));
  INV_X1     g5815(.I(new_n2656_), .ZN(new_n5873_));
  NOR3_X1    g5816(.A1(new_n372_), .A2(new_n1069_), .A3(new_n449_), .ZN(new_n5874_));
  NAND2_X1   g5817(.A1(new_n2240_), .A2(new_n439_), .ZN(new_n5875_));
  NOR4_X1    g5818(.A1(new_n5875_), .A2(new_n461_), .A3(new_n465_), .A4(new_n668_), .ZN(new_n5876_));
  NAND2_X1   g5819(.A1(new_n227_), .A2(new_n217_), .ZN(new_n5877_));
  NOR4_X1    g5820(.A1(new_n5877_), .A2(new_n273_), .A3(new_n359_), .A4(new_n891_), .ZN(new_n5878_));
  NAND4_X1   g5821(.A1(new_n5876_), .A2(new_n5878_), .A3(new_n5115_), .A4(new_n5874_), .ZN(new_n5879_));
  NOR4_X1    g5822(.A1(new_n2851_), .A2(new_n5873_), .A3(new_n4032_), .A4(new_n5879_), .ZN(new_n5880_));
  INV_X1     g5823(.I(new_n5880_), .ZN(new_n5881_));
  NOR2_X1    g5824(.A1(new_n5842_), .A2(new_n5848_), .ZN(new_n5882_));
  INV_X1     g5825(.I(new_n5882_), .ZN(new_n5883_));
  NOR2_X1    g5826(.A1(new_n5843_), .A2(new_n5847_), .ZN(new_n5884_));
  OAI21_X1   g5827(.A1(new_n5809_), .A2(new_n5884_), .B(new_n5883_), .ZN(new_n5885_));
  AOI22_X1   g5828(.A1(new_n5722_), .A2(new_n5725_), .B1(new_n5791_), .B2(new_n5797_), .ZN(new_n5886_));
  NOR4_X1    g5829(.A1(new_n5636_), .A2(new_n5718_), .A3(new_n5802_), .A4(new_n5803_), .ZN(new_n5887_));
  OAI21_X1   g5830(.A1(new_n5887_), .A2(new_n5886_), .B(new_n5857_), .ZN(new_n5888_));
  NAND2_X1   g5831(.A1(new_n5822_), .A2(new_n5820_), .ZN(new_n5889_));
  NAND2_X1   g5832(.A1(new_n5889_), .A2(new_n5817_), .ZN(new_n5890_));
  OAI22_X1   g5833(.A1(new_n4230_), .A2(new_n3493_), .B1(new_n4182_), .B2(new_n3396_), .ZN(new_n5891_));
  OAI21_X1   g5834(.A1(new_n3496_), .A2(new_n4474_), .B(new_n5891_), .ZN(new_n5892_));
  AOI21_X1   g5835(.A1(new_n5892_), .A2(new_n437_), .B(new_n3501_), .ZN(new_n5893_));
  XOR2_X1    g5836(.A1(new_n4484_), .A2(new_n5893_), .Z(new_n5894_));
  XOR2_X1    g5837(.A1(new_n3597_), .A2(new_n721_), .Z(new_n5895_));
  NAND2_X1   g5838(.A1(new_n5895_), .A2(new_n3977_), .ZN(new_n5896_));
  XOR2_X1    g5839(.A1(new_n5896_), .A2(new_n438_), .Z(new_n5897_));
  INV_X1     g5840(.I(new_n5897_), .ZN(new_n5898_));
  AND2_X2    g5841(.A1(new_n5894_), .A2(new_n5898_), .Z(new_n5899_));
  NOR2_X1    g5842(.A1(new_n5894_), .A2(new_n5898_), .ZN(new_n5900_));
  OAI21_X1   g5843(.A1(new_n5899_), .A2(new_n5900_), .B(new_n5890_), .ZN(new_n5901_));
  INV_X1     g5844(.I(new_n5890_), .ZN(new_n5902_));
  XOR2_X1    g5845(.A1(new_n5894_), .A2(new_n5898_), .Z(new_n5903_));
  NAND2_X1   g5846(.A1(new_n5902_), .A2(new_n5903_), .ZN(new_n5904_));
  NAND2_X1   g5847(.A1(new_n5904_), .A2(new_n5901_), .ZN(new_n5905_));
  INV_X1     g5848(.I(new_n5825_), .ZN(new_n5906_));
  INV_X1     g5849(.I(new_n5831_), .ZN(new_n5907_));
  XOR2_X1    g5850(.A1(new_n5827_), .A2(new_n721_), .Z(new_n5908_));
  AOI21_X1   g5851(.A1(new_n5825_), .A2(new_n5907_), .B(new_n5908_), .ZN(new_n5909_));
  AOI21_X1   g5852(.A1(new_n5906_), .A2(new_n5831_), .B(new_n5909_), .ZN(new_n5910_));
  XOR2_X1    g5853(.A1(new_n5905_), .A2(new_n5910_), .Z(new_n5911_));
  AND2_X2    g5854(.A1(new_n5835_), .A2(new_n5773_), .Z(new_n5912_));
  NOR2_X1    g5855(.A1(new_n5835_), .A2(new_n5773_), .ZN(new_n5913_));
  NOR2_X1    g5856(.A1(new_n5913_), .A2(new_n5749_), .ZN(new_n5914_));
  NOR3_X1    g5857(.A1(new_n5747_), .A2(new_n5912_), .A3(new_n5914_), .ZN(new_n5915_));
  NAND3_X1   g5858(.A1(new_n5834_), .A2(new_n5771_), .A3(new_n5812_), .ZN(new_n5916_));
  INV_X1     g5859(.I(new_n5916_), .ZN(new_n5917_));
  OAI21_X1   g5860(.A1(new_n5915_), .A2(new_n5917_), .B(new_n5911_), .ZN(new_n5918_));
  OR3_X2     g5861(.A1(new_n5915_), .A2(new_n5911_), .A3(new_n5917_), .Z(new_n5919_));
  NAND2_X1   g5862(.A1(new_n5919_), .A2(new_n5918_), .ZN(new_n5920_));
  NAND2_X1   g5863(.A1(new_n5888_), .A2(new_n5920_), .ZN(new_n5921_));
  OAI22_X1   g5864(.A1(new_n5636_), .A2(new_n5718_), .B1(new_n5802_), .B2(new_n5803_), .ZN(new_n5922_));
  NAND4_X1   g5865(.A1(new_n5722_), .A2(new_n5725_), .A3(new_n5791_), .A4(new_n5797_), .ZN(new_n5923_));
  NAND2_X1   g5866(.A1(new_n5922_), .A2(new_n5923_), .ZN(new_n5924_));
  INV_X1     g5867(.I(new_n5920_), .ZN(new_n5925_));
  NAND3_X1   g5868(.A1(new_n5924_), .A2(new_n5857_), .A3(new_n5925_), .ZN(new_n5926_));
  AOI21_X1   g5869(.A1(new_n5921_), .A2(new_n5926_), .B(new_n5885_), .ZN(new_n5927_));
  INV_X1     g5870(.I(new_n5885_), .ZN(new_n5928_));
  AOI21_X1   g5871(.A1(new_n5924_), .A2(new_n5857_), .B(new_n5925_), .ZN(new_n5929_));
  NOR2_X1    g5872(.A1(new_n5888_), .A2(new_n5920_), .ZN(new_n5930_));
  NOR3_X1    g5873(.A1(new_n5930_), .A2(new_n5929_), .A3(new_n5928_), .ZN(new_n5931_));
  OAI21_X1   g5874(.A1(new_n5931_), .A2(new_n5927_), .B(new_n5881_), .ZN(new_n5932_));
  OAI21_X1   g5875(.A1(new_n5930_), .A2(new_n5929_), .B(new_n5928_), .ZN(new_n5933_));
  NAND3_X1   g5876(.A1(new_n5921_), .A2(new_n5926_), .A3(new_n5885_), .ZN(new_n5934_));
  NAND3_X1   g5877(.A1(new_n5933_), .A2(new_n5934_), .A3(new_n5880_), .ZN(new_n5935_));
  NAND2_X1   g5878(.A1(new_n5932_), .A2(new_n5935_), .ZN(new_n5936_));
  NOR4_X1    g5879(.A1(new_n5867_), .A2(new_n5860_), .A3(new_n5861_), .A4(new_n5870_), .ZN(new_n5937_));
  NOR2_X1    g5880(.A1(new_n5937_), .A2(new_n4445_), .ZN(new_n5938_));
  XOR2_X1    g5881(.A1(new_n5936_), .A2(new_n5938_), .Z(\sin[13] ));
  NAND2_X1   g5882(.A1(new_n5920_), .A2(new_n5881_), .ZN(new_n5940_));
  NOR2_X1    g5883(.A1(new_n5914_), .A2(new_n5912_), .ZN(new_n5941_));
  OAI21_X1   g5884(.A1(new_n5746_), .A2(new_n5744_), .B(new_n5941_), .ZN(new_n5942_));
  NOR2_X1    g5885(.A1(new_n5911_), .A2(new_n5881_), .ZN(new_n5943_));
  NAND2_X1   g5886(.A1(new_n5942_), .A2(new_n5943_), .ZN(new_n5944_));
  OAI21_X1   g5887(.A1(new_n5881_), .A2(new_n5911_), .B(new_n5915_), .ZN(new_n5945_));
  NAND2_X1   g5888(.A1(new_n5945_), .A2(new_n5944_), .ZN(new_n5946_));
  NAND2_X1   g5889(.A1(new_n5946_), .A2(new_n5916_), .ZN(new_n5947_));
  NAND3_X1   g5890(.A1(new_n5945_), .A2(new_n5917_), .A3(new_n5944_), .ZN(new_n5948_));
  NAND3_X1   g5891(.A1(new_n5947_), .A2(new_n5843_), .A3(new_n5948_), .ZN(new_n5949_));
  AOI21_X1   g5892(.A1(new_n5947_), .A2(new_n5948_), .B(new_n5843_), .ZN(new_n5950_));
  OAI21_X1   g5893(.A1(new_n5847_), .A2(new_n5950_), .B(new_n5949_), .ZN(new_n5951_));
  OAI21_X1   g5894(.A1(new_n5951_), .A2(new_n5809_), .B(new_n5940_), .ZN(new_n5952_));
  INV_X1     g5895(.I(new_n5952_), .ZN(new_n5953_));
  NAND2_X1   g5896(.A1(new_n5925_), .A2(new_n5880_), .ZN(new_n5954_));
  NAND2_X1   g5897(.A1(new_n5954_), .A2(new_n5940_), .ZN(new_n5955_));
  INV_X1     g5898(.I(new_n5955_), .ZN(new_n5956_));
  AOI21_X1   g5899(.A1(new_n5924_), .A2(new_n5857_), .B(new_n5956_), .ZN(new_n5957_));
  NOR2_X1    g5900(.A1(new_n5888_), .A2(new_n5955_), .ZN(new_n5958_));
  OAI21_X1   g5901(.A1(new_n5958_), .A2(new_n5957_), .B(new_n5885_), .ZN(new_n5959_));
  INV_X1     g5902(.I(new_n5905_), .ZN(new_n5960_));
  AOI21_X1   g5903(.A1(new_n5916_), .A2(new_n5960_), .B(new_n5910_), .ZN(new_n5961_));
  INV_X1     g5904(.I(new_n5961_), .ZN(new_n5962_));
  OAI22_X1   g5905(.A1(new_n5942_), .A2(new_n5962_), .B1(new_n5960_), .B2(new_n5916_), .ZN(new_n5963_));
  INV_X1     g5906(.I(new_n5963_), .ZN(new_n5964_));
  NOR2_X1    g5907(.A1(new_n5902_), .A2(new_n5899_), .ZN(new_n5965_));
  NOR2_X1    g5908(.A1(new_n5965_), .A2(new_n5900_), .ZN(new_n5966_));
  NAND2_X1   g5909(.A1(new_n5550_), .A2(new_n437_), .ZN(new_n5967_));
  OAI21_X1   g5910(.A1(new_n4480_), .A2(new_n5967_), .B(new_n3393_), .ZN(new_n5968_));
  XOR2_X1    g5911(.A1(new_n4688_), .A2(new_n5968_), .Z(new_n5969_));
  NOR2_X1    g5912(.A1(new_n4192_), .A2(new_n438_), .ZN(new_n5970_));
  INV_X1     g5913(.I(new_n5970_), .ZN(new_n5971_));
  NAND2_X1   g5914(.A1(new_n721_), .A2(new_n437_), .ZN(new_n5972_));
  OAI21_X1   g5915(.A1(new_n437_), .A2(new_n721_), .B(new_n3597_), .ZN(new_n5973_));
  NAND3_X1   g5916(.A1(new_n3977_), .A2(new_n5972_), .A3(new_n5973_), .ZN(new_n5974_));
  NOR2_X1    g5917(.A1(new_n5971_), .A2(new_n5974_), .ZN(new_n5975_));
  INV_X1     g5918(.I(new_n5975_), .ZN(new_n5976_));
  NAND2_X1   g5919(.A1(new_n5971_), .A2(new_n5974_), .ZN(new_n5977_));
  AOI21_X1   g5920(.A1(new_n5976_), .A2(new_n5977_), .B(new_n5969_), .ZN(new_n5978_));
  XOR2_X1    g5921(.A1(new_n5970_), .A2(new_n5974_), .Z(new_n5979_));
  INV_X1     g5922(.I(new_n5979_), .ZN(new_n5980_));
  AOI21_X1   g5923(.A1(new_n5969_), .A2(new_n5980_), .B(new_n5978_), .ZN(new_n5981_));
  NOR2_X1    g5924(.A1(new_n5966_), .A2(new_n5981_), .ZN(new_n5982_));
  INV_X1     g5925(.I(new_n5966_), .ZN(new_n5983_));
  INV_X1     g5926(.I(new_n5981_), .ZN(new_n5984_));
  NOR2_X1    g5927(.A1(new_n5983_), .A2(new_n5984_), .ZN(new_n5985_));
  NOR2_X1    g5928(.A1(new_n5985_), .A2(new_n5982_), .ZN(new_n5986_));
  NOR2_X1    g5929(.A1(new_n5964_), .A2(new_n5986_), .ZN(new_n5987_));
  XOR2_X1    g5930(.A1(new_n5966_), .A2(new_n5984_), .Z(new_n5988_));
  NOR2_X1    g5931(.A1(new_n5963_), .A2(new_n5988_), .ZN(new_n5989_));
  NOR2_X1    g5932(.A1(new_n5987_), .A2(new_n5989_), .ZN(new_n5990_));
  NAND2_X1   g5933(.A1(new_n523_), .A2(new_n3967_), .ZN(new_n5991_));
  NAND4_X1   g5934(.A1(new_n331_), .A2(new_n197_), .A3(new_n375_), .A4(new_n325_), .ZN(new_n5992_));
  NAND2_X1   g5935(.A1(new_n2340_), .A2(new_n2451_), .ZN(new_n5993_));
  OR3_X2     g5936(.A1(new_n5993_), .A2(new_n2448_), .A3(new_n5992_), .Z(new_n5994_));
  NOR4_X1    g5937(.A1(new_n5994_), .A2(new_n404_), .A3(new_n543_), .A4(new_n5991_), .ZN(new_n5995_));
  NAND4_X1   g5938(.A1(new_n5995_), .A2(new_n2392_), .A3(new_n2613_), .A4(new_n1439_), .ZN(new_n5996_));
  INV_X1     g5939(.I(new_n5996_), .ZN(new_n5997_));
  XOR2_X1    g5940(.A1(new_n5990_), .A2(new_n5997_), .Z(new_n5998_));
  NAND2_X1   g5941(.A1(new_n5959_), .A2(new_n5998_), .ZN(new_n5999_));
  INV_X1     g5942(.I(new_n5999_), .ZN(new_n6000_));
  NOR2_X1    g5943(.A1(new_n5959_), .A2(new_n5998_), .ZN(new_n6001_));
  OAI21_X1   g5944(.A1(new_n6000_), .A2(new_n6001_), .B(new_n5953_), .ZN(new_n6002_));
  INV_X1     g5945(.I(new_n5998_), .ZN(new_n6003_));
  NOR2_X1    g5946(.A1(new_n5959_), .A2(new_n6003_), .ZN(new_n6004_));
  OR2_X2     g5947(.A1(new_n5958_), .A2(new_n5957_), .Z(new_n6005_));
  AOI21_X1   g5948(.A1(new_n6005_), .A2(new_n5885_), .B(new_n5998_), .ZN(new_n6006_));
  OAI21_X1   g5949(.A1(new_n6006_), .A2(new_n6004_), .B(new_n5952_), .ZN(new_n6007_));
  NAND2_X1   g5950(.A1(new_n6002_), .A2(new_n6007_), .ZN(new_n6008_));
  AOI21_X1   g5951(.A1(new_n5933_), .A2(new_n5934_), .B(new_n5880_), .ZN(new_n6009_));
  NOR3_X1    g5952(.A1(new_n5931_), .A2(new_n5927_), .A3(new_n5881_), .ZN(new_n6010_));
  INV_X1     g5953(.I(new_n5861_), .ZN(new_n6011_));
  NAND4_X1   g5954(.A1(new_n5743_), .A2(new_n6011_), .A3(new_n5869_), .A4(new_n5859_), .ZN(new_n6012_));
  NOR3_X1    g5955(.A1(new_n6010_), .A2(new_n6009_), .A3(new_n6012_), .ZN(new_n6013_));
  NOR2_X1    g5956(.A1(new_n6013_), .A2(new_n4445_), .ZN(new_n6014_));
  XOR2_X1    g5957(.A1(new_n6008_), .A2(new_n6014_), .Z(\sin[14] ));
  NAND3_X1   g5958(.A1(new_n5932_), .A2(new_n5935_), .A3(new_n5937_), .ZN(new_n6016_));
  NOR2_X1    g5959(.A1(new_n6008_), .A2(new_n6016_), .ZN(new_n6017_));
  NOR2_X1    g5960(.A1(new_n6017_), .A2(new_n4445_), .ZN(new_n6018_));
  XOR2_X1    g5961(.A1(new_n5952_), .A2(new_n5998_), .Z(new_n6019_));
  AND3_X2    g5962(.A1(new_n6005_), .A2(new_n5885_), .A3(new_n6019_), .Z(new_n6020_));
  NOR2_X1    g5963(.A1(new_n5951_), .A2(new_n5809_), .ZN(new_n6021_));
  INV_X1     g5964(.I(new_n5990_), .ZN(new_n6022_));
  NAND2_X1   g5965(.A1(new_n6021_), .A2(new_n6022_), .ZN(new_n6023_));
  NOR2_X1    g5966(.A1(new_n5940_), .A2(new_n5996_), .ZN(new_n6024_));
  OAI21_X1   g5967(.A1(new_n6021_), .A2(new_n6022_), .B(new_n6024_), .ZN(new_n6025_));
  AOI22_X1   g5968(.A1(new_n4747_), .A2(new_n3494_), .B1(new_n3393_), .B2(new_n4475_), .ZN(new_n6026_));
  XOR2_X1    g5969(.A1(new_n6026_), .A2(new_n4182_), .Z(new_n6027_));
  NAND2_X1   g5970(.A1(new_n6027_), .A2(new_n4232_), .ZN(new_n6028_));
  XOR2_X1    g5971(.A1(new_n6028_), .A2(new_n438_), .Z(new_n6029_));
  AOI21_X1   g5972(.A1(new_n5969_), .A2(new_n5977_), .B(new_n5975_), .ZN(new_n6030_));
  INV_X1     g5973(.I(new_n6030_), .ZN(new_n6031_));
  XOR2_X1    g5974(.A1(new_n6029_), .A2(new_n6031_), .Z(new_n6032_));
  NOR2_X1    g5975(.A1(new_n5988_), .A2(new_n6032_), .ZN(new_n6033_));
  XNOR2_X1   g5976(.A1(new_n6033_), .A2(new_n5982_), .ZN(new_n6034_));
  XOR2_X1    g5977(.A1(new_n5963_), .A2(new_n6034_), .Z(new_n6035_));
  AOI21_X1   g5978(.A1(new_n6025_), .A2(new_n6023_), .B(new_n6035_), .ZN(new_n6036_));
  NAND2_X1   g5979(.A1(new_n6025_), .A2(new_n6023_), .ZN(new_n6037_));
  INV_X1     g5980(.I(new_n6035_), .ZN(new_n6038_));
  NOR2_X1    g5981(.A1(new_n6037_), .A2(new_n6038_), .ZN(new_n6039_));
  NOR2_X1    g5982(.A1(new_n6039_), .A2(new_n6036_), .ZN(new_n6040_));
  NOR2_X1    g5983(.A1(new_n6020_), .A2(new_n6040_), .ZN(new_n6041_));
  NAND3_X1   g5984(.A1(new_n6005_), .A2(new_n5885_), .A3(new_n6019_), .ZN(new_n6042_));
  OR2_X2     g5985(.A1(new_n6039_), .A2(new_n6036_), .Z(new_n6043_));
  NOR2_X1    g5986(.A1(new_n6043_), .A2(new_n6042_), .ZN(new_n6044_));
  OAI21_X1   g5987(.A1(new_n6041_), .A2(new_n6044_), .B(new_n6018_), .ZN(new_n6045_));
  XOR2_X1    g5988(.A1(new_n6042_), .A2(new_n6040_), .Z(new_n6046_));
  OAI21_X1   g5989(.A1(new_n6018_), .A2(new_n6046_), .B(new_n6045_), .ZN(\sin[15] ));
  AOI21_X1   g5990(.A1(new_n6025_), .A2(new_n6023_), .B(new_n6038_), .ZN(new_n6048_));
  INV_X1     g5991(.I(new_n6029_), .ZN(new_n6049_));
  NOR2_X1    g5992(.A1(new_n6032_), .A2(new_n5981_), .ZN(new_n6050_));
  NOR2_X1    g5993(.A1(new_n6050_), .A2(new_n5983_), .ZN(new_n6051_));
  AOI21_X1   g5994(.A1(new_n5981_), .A2(new_n6032_), .B(new_n6051_), .ZN(new_n6052_));
  XOR2_X1    g5995(.A1(new_n6026_), .A2(new_n4232_), .Z(new_n6053_));
  XOR2_X1    g5996(.A1(new_n6026_), .A2(new_n438_), .Z(new_n6054_));
  AOI21_X1   g5997(.A1(new_n6054_), .A2(new_n6053_), .B(new_n4182_), .ZN(new_n6055_));
  XOR2_X1    g5998(.A1(new_n6055_), .A2(new_n4230_), .Z(new_n6056_));
  INV_X1     g5999(.I(new_n6056_), .ZN(new_n6057_));
  AOI21_X1   g6000(.A1(new_n5963_), .A2(new_n6052_), .B(new_n6057_), .ZN(new_n6058_));
  NOR3_X1    g6001(.A1(new_n6058_), .A2(new_n6049_), .A3(new_n6030_), .ZN(new_n6059_));
  INV_X1     g6002(.I(new_n6059_), .ZN(new_n6060_));
  OAI21_X1   g6003(.A1(new_n6058_), .A2(new_n6030_), .B(new_n6049_), .ZN(new_n6061_));
  AOI21_X1   g6004(.A1(new_n6060_), .A2(new_n6061_), .B(new_n4192_), .ZN(new_n6062_));
  INV_X1     g6005(.I(new_n6061_), .ZN(new_n6063_));
  NOR3_X1    g6006(.A1(new_n6063_), .A2(new_n4182_), .A3(new_n6059_), .ZN(new_n6064_));
  OAI21_X1   g6007(.A1(new_n6062_), .A2(new_n6064_), .B(new_n4475_), .ZN(new_n6065_));
  NOR2_X1    g6008(.A1(new_n6065_), .A2(new_n438_), .ZN(new_n6066_));
  OAI21_X1   g6009(.A1(new_n6063_), .A2(new_n6059_), .B(new_n4182_), .ZN(new_n6067_));
  NAND3_X1   g6010(.A1(new_n6060_), .A2(new_n4192_), .A3(new_n6061_), .ZN(new_n6068_));
  NAND2_X1   g6011(.A1(new_n6067_), .A2(new_n6068_), .ZN(new_n6069_));
  AOI21_X1   g6012(.A1(new_n6069_), .A2(new_n4475_), .B(new_n437_), .ZN(new_n6070_));
  INV_X1     g6013(.I(new_n4034_), .ZN(new_n6071_));
  NOR2_X1    g6014(.A1(new_n209_), .A2(new_n608_), .ZN(new_n6072_));
  NAND4_X1   g6015(.A1(new_n6072_), .A2(new_n151_), .A3(new_n241_), .A4(new_n593_), .ZN(new_n6073_));
  NOR3_X1    g6016(.A1(new_n2251_), .A2(new_n6073_), .A3(new_n896_), .ZN(new_n6074_));
  NAND4_X1   g6017(.A1(new_n6071_), .A2(new_n4055_), .A3(new_n5878_), .A4(new_n6074_), .ZN(new_n6075_));
  NOR2_X1    g6018(.A1(new_n6075_), .A2(new_n2273_), .ZN(new_n6076_));
  OAI21_X1   g6019(.A1(new_n6066_), .A2(new_n6070_), .B(new_n6076_), .ZN(new_n6077_));
  NAND3_X1   g6020(.A1(new_n6069_), .A2(new_n437_), .A3(new_n4475_), .ZN(new_n6078_));
  NAND2_X1   g6021(.A1(new_n6065_), .A2(new_n438_), .ZN(new_n6079_));
  INV_X1     g6022(.I(new_n6076_), .ZN(new_n6080_));
  NAND3_X1   g6023(.A1(new_n6079_), .A2(new_n6078_), .A3(new_n6080_), .ZN(new_n6081_));
  NAND2_X1   g6024(.A1(new_n6077_), .A2(new_n6081_), .ZN(new_n6082_));
  NAND2_X1   g6025(.A1(new_n6082_), .A2(new_n6048_), .ZN(new_n6083_));
  NAND3_X1   g6026(.A1(new_n6079_), .A2(new_n6078_), .A3(new_n6076_), .ZN(new_n6084_));
  OAI21_X1   g6027(.A1(new_n6066_), .A2(new_n6070_), .B(new_n6080_), .ZN(new_n6085_));
  AOI21_X1   g6028(.A1(new_n6084_), .A2(new_n6085_), .B(new_n6048_), .ZN(new_n6086_));
  INV_X1     g6029(.I(new_n6086_), .ZN(new_n6087_));
  NAND2_X1   g6030(.A1(new_n6087_), .A2(new_n6083_), .ZN(new_n6088_));
  XOR2_X1    g6031(.A1(new_n6044_), .A2(new_n6088_), .Z(new_n6089_));
  NAND4_X1   g6032(.A1(new_n5932_), .A2(new_n6040_), .A3(new_n5935_), .A4(new_n5937_), .ZN(new_n6090_));
  NAND2_X1   g6033(.A1(new_n6016_), .A2(new_n6043_), .ZN(new_n6091_));
  NAND2_X1   g6034(.A1(new_n6091_), .A2(new_n6090_), .ZN(new_n6092_));
  AOI21_X1   g6035(.A1(new_n6002_), .A2(new_n6007_), .B(new_n6042_), .ZN(new_n6093_));
  NAND2_X1   g6036(.A1(new_n6092_), .A2(new_n6093_), .ZN(new_n6094_));
  INV_X1     g6037(.I(new_n6094_), .ZN(new_n6095_));
  NOR2_X1    g6038(.A1(new_n6095_), .A2(new_n4445_), .ZN(new_n6096_));
  NAND2_X1   g6039(.A1(new_n6089_), .A2(new_n4404_), .ZN(new_n6097_));
  OAI22_X1   g6040(.A1(new_n6096_), .A2(new_n6089_), .B1(new_n6095_), .B2(new_n6097_), .ZN(\sin[16] ));
  NAND2_X1   g6041(.A1(new_n6085_), .A2(new_n6084_), .ZN(new_n6099_));
  INV_X1     g6042(.I(new_n2915_), .ZN(new_n6100_));
  NAND4_X1   g6043(.A1(new_n2240_), .A2(new_n201_), .A3(new_n310_), .A4(new_n353_), .ZN(new_n6101_));
  NOR3_X1    g6044(.A1(new_n2854_), .A2(new_n6101_), .A3(new_n392_), .ZN(new_n6102_));
  NOR4_X1    g6045(.A1(new_n372_), .A2(new_n416_), .A3(new_n281_), .A4(new_n399_), .ZN(new_n6103_));
  NAND4_X1   g6046(.A1(new_n584_), .A2(new_n462_), .A3(new_n6102_), .A4(new_n6103_), .ZN(new_n6104_));
  NOR2_X1    g6047(.A1(new_n6100_), .A2(new_n6104_), .ZN(new_n6105_));
  NAND3_X1   g6048(.A1(new_n6099_), .A2(new_n6077_), .A3(new_n6105_), .ZN(new_n6106_));
  AOI21_X1   g6049(.A1(new_n6079_), .A2(new_n6078_), .B(new_n6080_), .ZN(new_n6107_));
  INV_X1     g6050(.I(new_n6107_), .ZN(new_n6108_));
  AOI21_X1   g6051(.A1(new_n6106_), .A2(new_n6108_), .B(new_n6048_), .ZN(new_n6109_));
  INV_X1     g6052(.I(new_n6048_), .ZN(new_n6110_));
  INV_X1     g6053(.I(new_n6077_), .ZN(new_n6111_));
  NOR3_X1    g6054(.A1(new_n6066_), .A2(new_n6070_), .A3(new_n6080_), .ZN(new_n6112_));
  AOI21_X1   g6055(.A1(new_n6079_), .A2(new_n6078_), .B(new_n6076_), .ZN(new_n6113_));
  OAI21_X1   g6056(.A1(new_n6112_), .A2(new_n6113_), .B(new_n6105_), .ZN(new_n6114_));
  NOR2_X1    g6057(.A1(new_n6114_), .A2(new_n6111_), .ZN(new_n6115_));
  NOR3_X1    g6058(.A1(new_n6115_), .A2(new_n6110_), .A3(new_n6107_), .ZN(new_n6116_));
  NOR2_X1    g6059(.A1(new_n6116_), .A2(new_n6109_), .ZN(new_n6117_));
  AOI21_X1   g6060(.A1(new_n6048_), .A2(new_n6082_), .B(new_n6086_), .ZN(new_n6118_));
  NAND2_X1   g6061(.A1(new_n6044_), .A2(new_n6118_), .ZN(new_n6119_));
  NOR2_X1    g6062(.A1(new_n6119_), .A2(new_n6117_), .ZN(new_n6120_));
  INV_X1     g6063(.I(new_n6120_), .ZN(new_n6121_));
  AOI21_X1   g6064(.A1(new_n6119_), .A2(new_n6117_), .B(new_n4445_), .ZN(new_n6122_));
  AOI21_X1   g6065(.A1(new_n6121_), .A2(new_n6122_), .B(new_n6094_), .ZN(new_n6123_));
  XNOR2_X1   g6066(.A1(new_n6123_), .A2(new_n6089_), .ZN(\sin[17] ));
  NOR2_X1    g6067(.A1(new_n1227_), .A2(new_n1225_), .ZN(new_n6125_));
  INV_X1     g6068(.I(new_n4041_), .ZN(new_n6126_));
  NOR2_X1    g6069(.A1(new_n388_), .A2(new_n325_), .ZN(new_n6127_));
  NAND4_X1   g6070(.A1(new_n6127_), .A2(new_n281_), .A3(new_n257_), .A4(new_n299_), .ZN(new_n6128_));
  NAND4_X1   g6071(.A1(new_n739_), .A2(new_n221_), .A3(new_n416_), .A4(new_n367_), .ZN(new_n6129_));
  NOR4_X1    g6072(.A1(new_n6128_), .A2(new_n6129_), .A3(new_n2652_), .A4(new_n911_), .ZN(new_n6130_));
  NAND4_X1   g6073(.A1(new_n6126_), .A2(new_n1142_), .A3(new_n6125_), .A4(new_n6130_), .ZN(new_n6131_));
  NAND2_X1   g6074(.A1(new_n6076_), .A2(new_n6105_), .ZN(new_n6132_));
  NAND3_X1   g6075(.A1(new_n6079_), .A2(new_n6078_), .A3(new_n6132_), .ZN(new_n6133_));
  OAI21_X1   g6076(.A1(new_n6076_), .A2(new_n6105_), .B(new_n6133_), .ZN(new_n6134_));
  NOR2_X1    g6077(.A1(new_n6134_), .A2(new_n6110_), .ZN(new_n6135_));
  NOR2_X1    g6078(.A1(new_n6135_), .A2(new_n6131_), .ZN(new_n6136_));
  INV_X1     g6079(.I(new_n6136_), .ZN(new_n6137_));
  INV_X1     g6080(.I(new_n6131_), .ZN(new_n6138_));
  INV_X1     g6081(.I(new_n6135_), .ZN(new_n6139_));
  NOR2_X1    g6082(.A1(new_n6139_), .A2(new_n6138_), .ZN(new_n6140_));
  OR3_X2     g6083(.A1(new_n6120_), .A2(new_n6136_), .A3(new_n6140_), .Z(new_n6141_));
  OAI21_X1   g6084(.A1(new_n6121_), .A2(new_n6137_), .B(new_n6141_), .ZN(new_n6142_));
  NAND3_X1   g6085(.A1(new_n6092_), .A2(new_n6093_), .A3(new_n6117_), .ZN(new_n6143_));
  NOR4_X1    g6086(.A1(new_n6043_), .A2(new_n6010_), .A3(new_n6009_), .A4(new_n6012_), .ZN(new_n6144_));
  NOR2_X1    g6087(.A1(new_n6013_), .A2(new_n6040_), .ZN(new_n6145_));
  NOR2_X1    g6088(.A1(new_n6145_), .A2(new_n6144_), .ZN(new_n6146_));
  INV_X1     g6089(.I(new_n6001_), .ZN(new_n6147_));
  AOI21_X1   g6090(.A1(new_n6147_), .A2(new_n5999_), .B(new_n5952_), .ZN(new_n6148_));
  INV_X1     g6091(.I(new_n6004_), .ZN(new_n6149_));
  NAND2_X1   g6092(.A1(new_n5959_), .A2(new_n6003_), .ZN(new_n6150_));
  AOI21_X1   g6093(.A1(new_n6149_), .A2(new_n6150_), .B(new_n5953_), .ZN(new_n6151_));
  OAI21_X1   g6094(.A1(new_n6148_), .A2(new_n6151_), .B(new_n6020_), .ZN(new_n6152_));
  OAI21_X1   g6095(.A1(new_n6115_), .A2(new_n6107_), .B(new_n6110_), .ZN(new_n6153_));
  NAND3_X1   g6096(.A1(new_n6106_), .A2(new_n6048_), .A3(new_n6108_), .ZN(new_n6154_));
  NAND2_X1   g6097(.A1(new_n6153_), .A2(new_n6154_), .ZN(new_n6155_));
  OAI21_X1   g6098(.A1(new_n6146_), .A2(new_n6152_), .B(new_n6155_), .ZN(new_n6156_));
  NOR2_X1    g6099(.A1(new_n6155_), .A2(new_n6118_), .ZN(new_n6157_));
  AOI21_X1   g6100(.A1(new_n6153_), .A2(new_n6154_), .B(new_n6088_), .ZN(new_n6158_));
  OAI21_X1   g6101(.A1(new_n6157_), .A2(new_n6158_), .B(new_n6044_), .ZN(new_n6159_));
  AOI21_X1   g6102(.A1(new_n6156_), .A2(new_n6143_), .B(new_n6159_), .ZN(new_n6160_));
  OAI21_X1   g6103(.A1(new_n4445_), .A2(new_n6160_), .B(new_n6142_), .ZN(new_n6161_));
  OR3_X2     g6104(.A1(new_n6142_), .A2(new_n4445_), .A3(new_n6160_), .Z(new_n6162_));
  NAND2_X1   g6105(.A1(new_n6162_), .A2(new_n6161_), .ZN(\sin[18] ));
  NOR2_X1    g6106(.A1(new_n505_), .A2(new_n221_), .ZN(new_n6164_));
  NAND3_X1   g6107(.A1(new_n323_), .A2(new_n859_), .A3(new_n363_), .ZN(new_n6165_));
  NAND4_X1   g6108(.A1(new_n401_), .A2(new_n388_), .A3(new_n921_), .A4(new_n240_), .ZN(new_n6166_));
  NAND2_X1   g6109(.A1(new_n652_), .A2(new_n5113_), .ZN(new_n6167_));
  NOR4_X1    g6110(.A1(new_n2892_), .A2(new_n6165_), .A3(new_n6166_), .A4(new_n6167_), .ZN(new_n6168_));
  NAND4_X1   g6111(.A1(new_n6168_), .A2(new_n785_), .A3(new_n1243_), .A4(new_n6164_), .ZN(new_n6169_));
  INV_X1     g6112(.I(new_n6169_), .ZN(new_n6170_));
  NAND2_X1   g6113(.A1(new_n6135_), .A2(new_n6170_), .ZN(new_n6171_));
  OAI22_X1   g6114(.A1(new_n6140_), .A2(new_n6170_), .B1(new_n6138_), .B2(new_n6171_), .ZN(new_n6172_));
  NAND2_X1   g6115(.A1(new_n6120_), .A2(new_n6137_), .ZN(new_n6173_));
  NOR2_X1    g6116(.A1(new_n6172_), .A2(new_n6136_), .ZN(new_n6174_));
  AOI22_X1   g6117(.A1(new_n6173_), .A2(new_n6172_), .B1(new_n6174_), .B2(new_n6120_), .ZN(new_n6175_));
  NOR4_X1    g6118(.A1(new_n6160_), .A2(new_n6121_), .A3(new_n6138_), .A4(new_n6139_), .ZN(new_n6176_));
  NOR2_X1    g6119(.A1(new_n6176_), .A2(new_n4445_), .ZN(new_n6177_));
  NAND2_X1   g6120(.A1(new_n6175_), .A2(new_n4404_), .ZN(new_n6178_));
  OAI22_X1   g6121(.A1(new_n6177_), .A2(new_n6175_), .B1(new_n6176_), .B2(new_n6178_), .ZN(\sin[19] ));
  NOR3_X1    g6122(.A1(new_n6146_), .A2(new_n6152_), .A3(new_n6155_), .ZN(new_n6180_));
  AOI21_X1   g6123(.A1(new_n6092_), .A2(new_n6093_), .B(new_n6117_), .ZN(new_n6181_));
  NAND2_X1   g6124(.A1(new_n6020_), .A2(new_n6040_), .ZN(new_n6182_));
  NAND3_X1   g6125(.A1(new_n6088_), .A2(new_n6153_), .A3(new_n6154_), .ZN(new_n6183_));
  OAI21_X1   g6126(.A1(new_n6109_), .A2(new_n6116_), .B(new_n6118_), .ZN(new_n6184_));
  AOI21_X1   g6127(.A1(new_n6184_), .A2(new_n6183_), .B(new_n6182_), .ZN(new_n6185_));
  OAI21_X1   g6128(.A1(new_n6180_), .A2(new_n6181_), .B(new_n6185_), .ZN(new_n6186_));
  NAND4_X1   g6129(.A1(new_n6186_), .A2(new_n6120_), .A3(new_n6131_), .A4(new_n6135_), .ZN(new_n6187_));
  NAND2_X1   g6130(.A1(new_n6175_), .A2(new_n4445_), .ZN(new_n6188_));
  NAND3_X1   g6131(.A1(new_n5117_), .A2(new_n499_), .A3(new_n649_), .ZN(new_n6189_));
  NOR3_X1    g6132(.A1(new_n892_), .A2(new_n160_), .A3(new_n395_), .ZN(new_n6190_));
  NAND4_X1   g6133(.A1(new_n6190_), .A2(new_n2274_), .A3(new_n258_), .A4(new_n205_), .ZN(new_n6191_));
  NOR3_X1    g6134(.A1(new_n4176_), .A2(new_n6189_), .A3(new_n6191_), .ZN(new_n6192_));
  NAND3_X1   g6135(.A1(new_n6192_), .A2(new_n5499_), .A3(new_n742_), .ZN(new_n6193_));
  NOR4_X1    g6136(.A1(new_n6135_), .A2(new_n6131_), .A3(new_n6170_), .A4(new_n6193_), .ZN(new_n6194_));
  INV_X1     g6137(.I(new_n6194_), .ZN(new_n6195_));
  NOR3_X1    g6138(.A1(new_n6121_), .A2(new_n6137_), .A3(new_n6195_), .ZN(new_n6200_));
  OAI21_X1   g6139(.A1(new_n6188_), .A2(new_n6187_), .B(new_n6200_), .ZN(new_n6201_));
  INV_X1     g6140(.I(new_n6200_), .ZN(new_n6202_));
  NAND4_X1   g6141(.A1(new_n6176_), .A2(new_n4445_), .A3(new_n6175_), .A4(new_n6202_), .ZN(new_n6203_));
  NAND2_X1   g6142(.A1(new_n6203_), .A2(new_n6201_), .ZN(\sin[20] ));
  NAND4_X1   g6143(.A1(new_n6155_), .A2(new_n6044_), .A3(new_n6118_), .A4(new_n6194_), .ZN(new_n6205_));
  NOR3_X1    g6144(.A1(new_n6131_), .A2(new_n6169_), .A3(new_n6193_), .ZN(new_n6206_));
  INV_X1     g6145(.I(new_n6206_), .ZN(new_n6207_));
  NOR3_X1    g6146(.A1(new_n6134_), .A2(new_n6110_), .A3(new_n6207_), .ZN(new_n6208_));
  INV_X1     g6147(.I(new_n6208_), .ZN(new_n6209_));
  NOR2_X1    g6148(.A1(new_n227_), .A2(new_n366_), .ZN(new_n6210_));
  NAND4_X1   g6149(.A1(new_n266_), .A2(new_n557_), .A3(new_n4177_), .A4(new_n6210_), .ZN(new_n6211_));
  NAND2_X1   g6150(.A1(new_n6209_), .A2(new_n6211_), .ZN(new_n6212_));
  INV_X1     g6151(.I(new_n6211_), .ZN(new_n6213_));
  NAND2_X1   g6152(.A1(new_n6208_), .A2(new_n6213_), .ZN(new_n6214_));
  NAND2_X1   g6153(.A1(new_n6212_), .A2(new_n6214_), .ZN(new_n6215_));
  XOR2_X1    g6154(.A1(new_n6205_), .A2(new_n6215_), .Z(new_n6216_));
  AOI21_X1   g6155(.A1(new_n6187_), .A2(new_n6175_), .B(new_n6202_), .ZN(new_n6217_));
  NOR2_X1    g6156(.A1(new_n6217_), .A2(new_n4445_), .ZN(new_n6218_));
  NAND2_X1   g6157(.A1(new_n6216_), .A2(new_n4404_), .ZN(new_n6219_));
  OAI22_X1   g6158(.A1(new_n6218_), .A2(new_n6216_), .B1(new_n6217_), .B2(new_n6219_), .ZN(\sin[21] ));
  INV_X1     g6159(.I(new_n6215_), .ZN(new_n6221_));
  NOR2_X1    g6160(.A1(new_n6221_), .A2(new_n6205_), .ZN(new_n6222_));
  NOR3_X1    g6161(.A1(new_n6119_), .A2(new_n6117_), .A3(new_n6195_), .ZN(new_n6223_));
  NAND2_X1   g6162(.A1(new_n6208_), .A2(new_n6211_), .ZN(new_n6224_));
  NAND2_X1   g6163(.A1(new_n266_), .A2(new_n525_), .ZN(new_n6225_));
  NAND2_X1   g6164(.A1(new_n6224_), .A2(new_n6225_), .ZN(new_n6226_));
  OAI21_X1   g6165(.A1(new_n6223_), .A2(new_n6215_), .B(new_n6226_), .ZN(new_n6227_));
  NOR2_X1    g6166(.A1(new_n6227_), .A2(new_n6222_), .ZN(new_n6228_));
  NOR3_X1    g6167(.A1(new_n6221_), .A2(new_n6205_), .A3(new_n6226_), .ZN(new_n6229_));
  NOR3_X1    g6168(.A1(new_n6228_), .A2(new_n4445_), .A3(new_n6229_), .ZN(new_n6230_));
  INV_X1     g6169(.I(new_n6230_), .ZN(new_n6231_));
  NAND3_X1   g6170(.A1(new_n6217_), .A2(new_n6231_), .A3(new_n6216_), .ZN(new_n6232_));
  INV_X1     g6171(.I(new_n6216_), .ZN(new_n6233_));
  INV_X1     g6172(.I(new_n6175_), .ZN(new_n6234_));
  OAI21_X1   g6173(.A1(new_n6176_), .A2(new_n6234_), .B(new_n6200_), .ZN(new_n6235_));
  OAI21_X1   g6174(.A1(new_n6235_), .A2(new_n6230_), .B(new_n6233_), .ZN(new_n6236_));
  NAND2_X1   g6175(.A1(new_n6236_), .A2(new_n6232_), .ZN(\sin[22] ));
  INV_X1     g6176(.I(new_n6228_), .ZN(new_n6238_));
  INV_X1     g6177(.I(new_n6229_), .ZN(new_n6239_));
  NAND2_X1   g6178(.A1(new_n6238_), .A2(new_n6239_), .ZN(new_n6240_));
  NOR2_X1    g6179(.A1(new_n6224_), .A2(new_n6225_), .ZN(new_n6241_));
  AOI22_X1   g6180(.A1(new_n6212_), .A2(new_n6214_), .B1(new_n6224_), .B2(new_n6225_), .ZN(new_n6242_));
  AOI21_X1   g6181(.A1(new_n6223_), .A2(new_n6242_), .B(new_n6241_), .ZN(new_n6243_));
  NOR3_X1    g6182(.A1(new_n84_), .A2(\a[21] ), .A3(\a[22] ), .ZN(new_n6244_));
  NAND3_X1   g6183(.A1(new_n6223_), .A2(new_n6215_), .A3(new_n6241_), .ZN(new_n6245_));
  NAND3_X1   g6184(.A1(new_n6243_), .A2(new_n6245_), .A3(new_n6244_), .ZN(new_n6246_));
  XOR2_X1    g6185(.A1(new_n6246_), .A2(new_n4445_), .Z(new_n6247_));
  NOR4_X1    g6186(.A1(new_n6247_), .A2(new_n6233_), .A3(new_n6235_), .A4(new_n6240_), .ZN(\sin[23] ));
  NAND2_X1   g6187(.A1(new_n6216_), .A2(new_n6245_), .ZN(new_n6249_));
  OAI21_X1   g6188(.A1(new_n6217_), .A2(new_n6249_), .B(new_n6240_), .ZN(new_n6250_));
  NOR2_X1    g6189(.A1(new_n6244_), .A2(new_n4445_), .ZN(new_n6251_));
  NAND2_X1   g6190(.A1(new_n6187_), .A2(new_n6175_), .ZN(new_n6252_));
  NOR4_X1    g6191(.A1(new_n6205_), .A2(new_n6209_), .A3(new_n6213_), .A4(new_n6225_), .ZN(new_n6253_));
  NAND3_X1   g6192(.A1(new_n6252_), .A2(new_n6200_), .A3(new_n6253_), .ZN(new_n6254_));
  AOI21_X1   g6193(.A1(new_n6250_), .A2(new_n6251_), .B(new_n6254_), .ZN(\sin[24] ));
endmodule


