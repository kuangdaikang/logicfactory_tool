// Benchmark "i2c" written by ABC on Fri Feb 25 15:09:05 2022

module i2c ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1136_, new_n1137_, new_n1138_, new_n1140_,
    new_n1141_, new_n1142_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1157_, new_n1158_, new_n1159_, new_n1162_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1236_, new_n1237_, new_n1238_, new_n1240_,
    new_n1241_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1276_,
    new_n1277_, new_n1278_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1300_, new_n1301_, new_n1302_, new_n1304_, new_n1305_, new_n1306_,
    new_n1308_, new_n1309_, new_n1310_, new_n1312_, new_n1313_, new_n1314_,
    new_n1316_, new_n1317_, new_n1318_, new_n1320_, new_n1321_, new_n1322_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1330_,
    new_n1331_, new_n1332_, new_n1334_, new_n1335_, new_n1336_, new_n1338_,
    new_n1339_, new_n1340_, new_n1342_, new_n1343_, new_n1344_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1365_,
    new_n1366_, new_n1367_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1377_, new_n1378_, new_n1379_,
    new_n1381_, new_n1382_, new_n1383_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1391_, new_n1392_, new_n1393_, new_n1395_,
    new_n1396_, new_n1397_, new_n1399_, new_n1400_, new_n1401_, new_n1403_,
    new_n1404_, new_n1405_, new_n1407_, new_n1408_, new_n1409_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1428_, new_n1429_, new_n1430_, new_n1432_,
    new_n1433_, new_n1434_, new_n1436_, new_n1437_, new_n1438_, new_n1440_,
    new_n1441_, new_n1442_, new_n1444_, new_n1445_, new_n1446_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1619_, new_n1620_, new_n1621_, new_n1623_,
    new_n1628_, new_n1629_, new_n1631_;
  assign new_n291_ = ~pi013 & ~pi014;
  assign new_n292_ = ~pi006 & ~pi007;
  assign new_n293_ = new_n291_ & new_n292_;
  assign new_n294_ = ~pi017 & ~pi021;
  assign new_n295_ = ~pi008 & new_n294_;
  assign new_n296_ = ~pi012 & new_n295_;
  assign new_n297_ = new_n293_ & new_n296_;
  assign new_n298_ = ~pi018 & ~pi019;
  assign new_n299_ = ~pi004 & ~pi016;
  assign new_n300_ = new_n298_ & new_n299_;
  assign new_n301_ = ~pi005 & ~pi022;
  assign new_n302_ = ~pi009 & ~pi011;
  assign new_n303_ = new_n301_ & new_n302_;
  assign new_n304_ = new_n300_ & new_n303_;
  assign new_n305_ = new_n297_ & new_n304_;
  assign new_n306_ = pi054 & ~new_n305_;
  assign new_n307_ = ~pi000 & ~new_n306_;
  assign new_n308_ = new_n301_ & ~new_n302_;
  assign new_n309_ = ~pi056 & new_n308_;
  assign new_n310_ = ~pi056 & ~new_n301_;
  assign new_n311_ = ~pi008 & ~pi021;
  assign new_n312_ = ~pi007 & pi013;
  assign new_n313_ = new_n311_ & new_n312_;
  assign new_n314_ = ~pi007 & new_n311_;
  assign new_n315_ = pi007 & ~new_n311_;
  assign new_n316_ = ~new_n314_ & ~new_n315_;
  assign new_n317_ = pi008 & pi021;
  assign new_n318_ = ~pi013 & ~new_n317_;
  assign new_n319_ = new_n316_ & new_n318_;
  assign new_n320_ = ~new_n313_ & ~new_n319_;
  assign new_n321_ = ~pi014 & ~new_n320_;
  assign new_n322_ = ~pi013 & pi014;
  assign new_n323_ = new_n314_ & new_n322_;
  assign new_n324_ = ~new_n321_ & ~new_n323_;
  assign new_n325_ = ~pi010 & ~new_n324_;
  assign new_n326_ = pi010 & new_n291_;
  assign new_n327_ = new_n314_ & new_n326_;
  assign new_n328_ = ~new_n325_ & ~new_n327_;
  assign new_n329_ = new_n301_ & ~new_n328_;
  assign new_n330_ = new_n300_ & new_n329_;
  assign new_n331_ = ~pi017 & new_n330_;
  assign new_n332_ = ~pi006 & ~pi012;
  assign new_n333_ = new_n331_ & new_n332_;
  assign new_n334_ = ~new_n310_ & ~new_n333_;
  assign new_n335_ = new_n302_ & ~new_n334_;
  assign new_n336_ = ~new_n309_ & ~new_n335_;
  assign new_n337_ = pi054 & ~new_n336_;
  assign new_n338_ = ~new_n307_ & ~new_n337_;
  assign new_n339_ = ~pi129 & ~new_n338_;
  assign po015 = pi003 | ~new_n339_;
  assign new_n341_ = ~pi011 & ~pi012;
  assign new_n342_ = new_n311_ & new_n341_;
  assign new_n343_ = new_n300_ & new_n342_;
  assign new_n344_ = ~pi010 & ~pi022;
  assign new_n345_ = ~pi007 & ~pi013;
  assign new_n346_ = ~pi005 & ~pi006;
  assign new_n347_ = new_n345_ & new_n346_;
  assign new_n348_ = ~pi014 & new_n347_;
  assign new_n349_ = new_n344_ & new_n348_;
  assign new_n350_ = new_n343_ & new_n349_;
  assign new_n351_ = ~pi017 & pi054;
  assign new_n352_ = ~new_n350_ & new_n351_;
  assign new_n353_ = ~pi001 & ~new_n352_;
  assign new_n354_ = ~pi014 & pi054;
  assign new_n355_ = ~pi008 & ~pi011;
  assign new_n356_ = new_n294_ & new_n355_;
  assign new_n357_ = ~pi005 & new_n332_;
  assign new_n358_ = pi005 & ~new_n332_;
  assign new_n359_ = ~new_n357_ & ~new_n358_;
  assign new_n360_ = pi006 & pi012;
  assign new_n361_ = ~pi007 & ~new_n360_;
  assign new_n362_ = new_n359_ & new_n361_;
  assign new_n363_ = pi007 & new_n357_;
  assign new_n364_ = ~new_n362_ & ~new_n363_;
  assign new_n365_ = ~pi013 & ~new_n364_;
  assign new_n366_ = new_n312_ & new_n357_;
  assign new_n367_ = ~new_n365_ & ~new_n366_;
  assign new_n368_ = ~pi009 & ~new_n367_;
  assign new_n369_ = new_n345_ & new_n357_;
  assign new_n370_ = pi009 & new_n369_;
  assign new_n371_ = ~new_n368_ & ~new_n370_;
  assign new_n372_ = new_n300_ & ~new_n371_;
  assign new_n373_ = new_n356_ & new_n372_;
  assign new_n374_ = new_n354_ & new_n373_;
  assign new_n375_ = new_n344_ & new_n374_;
  assign new_n376_ = ~new_n353_ & ~new_n375_;
  assign new_n377_ = ~pi129 & ~new_n376_;
  assign po016 = pi003 | ~new_n377_;
  assign new_n379_ = pi122 & pi127;
  assign new_n380_ = ~pi045 & ~pi048;
  assign new_n381_ = ~pi043 & ~pi047;
  assign new_n382_ = new_n380_ & new_n381_;
  assign new_n383_ = ~pi015 & ~pi020;
  assign new_n384_ = ~pi024 & ~pi049;
  assign new_n385_ = new_n383_ & new_n384_;
  assign new_n386_ = new_n382_ & new_n385_;
  assign new_n387_ = ~pi041 & ~pi046;
  assign new_n388_ = ~pi038 & ~pi050;
  assign new_n389_ = new_n387_ & new_n388_;
  assign new_n390_ = ~pi042 & ~pi044;
  assign new_n391_ = ~pi040 & new_n390_;
  assign new_n392_ = ~pi002 & new_n391_;
  assign new_n393_ = new_n389_ & new_n392_;
  assign new_n394_ = new_n386_ & new_n393_;
  assign new_n395_ = pi082 & ~new_n394_;
  assign new_n396_ = ~new_n379_ & ~new_n395_;
  assign new_n397_ = ~pi065 & new_n396_;
  assign new_n398_ = ~pi024 & ~pi045;
  assign new_n399_ = ~pi047 & ~pi048;
  assign new_n400_ = new_n398_ & new_n399_;
  assign new_n401_ = ~pi049 & new_n383_;
  assign new_n402_ = new_n400_ & new_n401_;
  assign new_n403_ = ~pi038 & ~pi040;
  assign new_n404_ = new_n390_ & new_n403_;
  assign new_n405_ = ~pi046 & ~pi050;
  assign new_n406_ = ~pi041 & new_n405_;
  assign new_n407_ = new_n404_ & new_n406_;
  assign new_n408_ = ~pi043 & new_n407_;
  assign new_n409_ = new_n402_ & new_n408_;
  assign new_n410_ = pi082 & ~new_n409_;
  assign new_n411_ = ~pi082 & new_n379_;
  assign new_n412_ = ~new_n410_ & ~new_n411_;
  assign new_n413_ = pi002 & ~new_n412_;
  assign new_n414_ = ~new_n397_ & ~new_n413_;
  assign po017 = ~pi129 & ~new_n414_;
  assign new_n416_ = ~pi009 & ~pi014;
  assign new_n417_ = new_n344_ & new_n416_;
  assign new_n418_ = new_n347_ & new_n417_;
  assign new_n419_ = ~pi008 & ~pi017;
  assign new_n420_ = new_n341_ & new_n419_;
  assign new_n421_ = ~pi021 & new_n300_;
  assign new_n422_ = new_n420_ & new_n421_;
  assign new_n423_ = new_n418_ & new_n422_;
  assign new_n424_ = ~pi061 & ~pi118;
  assign new_n425_ = ~new_n423_ & new_n424_;
  assign new_n426_ = pi000 & ~pi123;
  assign new_n427_ = ~pi113 & new_n426_;
  assign new_n428_ = ~new_n425_ & ~new_n427_;
  assign po018 = ~pi129 & ~new_n428_;
  assign new_n430_ = pi010 & ~pi022;
  assign new_n431_ = new_n416_ & new_n430_;
  assign new_n432_ = new_n369_ & new_n431_;
  assign new_n433_ = pi054 & new_n300_;
  assign new_n434_ = new_n356_ & new_n433_;
  assign new_n435_ = new_n432_ & new_n434_;
  assign new_n436_ = pi004 & ~pi054;
  assign new_n437_ = ~new_n435_ & ~new_n436_;
  assign new_n438_ = ~pi129 & ~new_n437_;
  assign po019 = ~pi003 & new_n438_;
  assign new_n440_ = pi005 & ~pi054;
  assign new_n441_ = ~pi007 & new_n332_;
  assign new_n442_ = ~pi025 & ~pi029;
  assign new_n443_ = pi028 & new_n442_;
  assign new_n444_ = new_n441_ & new_n443_;
  assign new_n445_ = ~pi013 & new_n417_;
  assign new_n446_ = new_n444_ & new_n445_;
  assign new_n447_ = ~pi059 & new_n356_;
  assign new_n448_ = ~pi016 & pi054;
  assign new_n449_ = ~pi004 & ~pi019;
  assign new_n450_ = ~pi018 & new_n449_;
  assign new_n451_ = ~pi005 & new_n450_;
  assign new_n452_ = new_n448_ & new_n451_;
  assign new_n453_ = new_n447_ & new_n452_;
  assign new_n454_ = new_n446_ & new_n453_;
  assign new_n455_ = ~new_n440_ & ~new_n454_;
  assign new_n456_ = ~pi129 & ~new_n455_;
  assign po020 = ~pi003 & new_n456_;
  assign new_n458_ = pi006 & ~pi054;
  assign new_n459_ = ~pi005 & ~pi007;
  assign new_n460_ = pi025 & ~pi029;
  assign new_n461_ = ~pi028 & new_n460_;
  assign new_n462_ = ~pi012 & new_n461_;
  assign new_n463_ = new_n459_ & new_n462_;
  assign new_n464_ = new_n445_ & new_n463_;
  assign new_n465_ = ~pi006 & new_n450_;
  assign new_n466_ = new_n448_ & new_n465_;
  assign new_n467_ = new_n447_ & new_n466_;
  assign new_n468_ = new_n464_ & new_n467_;
  assign new_n469_ = ~new_n458_ & ~new_n468_;
  assign new_n470_ = ~pi129 & ~new_n469_;
  assign po021 = ~pi003 & new_n470_;
  assign new_n472_ = pi007 & ~pi054;
  assign new_n473_ = ~pi018 & ~pi021;
  assign new_n474_ = pi008 & ~pi017;
  assign new_n475_ = new_n473_ & new_n474_;
  assign new_n476_ = ~pi007 & new_n449_;
  assign new_n477_ = new_n448_ & new_n476_;
  assign new_n478_ = new_n475_ & new_n477_;
  assign new_n479_ = ~pi006 & new_n341_;
  assign new_n480_ = ~pi005 & new_n479_;
  assign new_n481_ = new_n445_ & new_n480_;
  assign new_n482_ = new_n478_ & new_n481_;
  assign new_n483_ = ~new_n472_ & ~new_n482_;
  assign new_n484_ = ~pi129 & ~new_n483_;
  assign po022 = ~pi003 & new_n484_;
  assign new_n486_ = pi008 & ~pi054;
  assign new_n487_ = new_n369_ & new_n417_;
  assign new_n488_ = ~pi017 & ~pi018;
  assign new_n489_ = ~pi011 & pi021;
  assign new_n490_ = new_n488_ & new_n489_;
  assign new_n491_ = ~pi008 & new_n449_;
  assign new_n492_ = new_n448_ & new_n491_;
  assign new_n493_ = new_n490_ & new_n492_;
  assign new_n494_ = new_n487_ & new_n493_;
  assign new_n495_ = ~new_n486_ & ~new_n494_;
  assign new_n496_ = ~pi129 & ~new_n495_;
  assign po023 = ~pi003 & new_n496_;
  assign new_n498_ = pi009 & ~pi054;
  assign new_n499_ = new_n291_ & new_n344_;
  assign new_n500_ = pi011 & new_n459_;
  assign new_n501_ = new_n332_ & new_n500_;
  assign new_n502_ = new_n499_ & new_n501_;
  assign new_n503_ = new_n419_ & new_n473_;
  assign new_n504_ = ~pi009 & new_n449_;
  assign new_n505_ = new_n448_ & new_n504_;
  assign new_n506_ = new_n503_ & new_n505_;
  assign new_n507_ = new_n502_ & new_n506_;
  assign new_n508_ = ~new_n498_ & ~new_n507_;
  assign new_n509_ = ~pi129 & ~new_n508_;
  assign po024 = ~pi003 & new_n509_;
  assign new_n511_ = pi010 & ~pi054;
  assign new_n512_ = ~pi010 & new_n449_;
  assign new_n513_ = new_n448_ & new_n512_;
  assign new_n514_ = new_n503_ & new_n513_;
  assign new_n515_ = new_n459_ & new_n479_;
  assign new_n516_ = ~pi009 & ~pi022;
  assign new_n517_ = new_n322_ & new_n516_;
  assign new_n518_ = new_n515_ & new_n517_;
  assign new_n519_ = new_n514_ & new_n518_;
  assign new_n520_ = ~new_n511_ & ~new_n519_;
  assign new_n521_ = ~pi129 & ~new_n520_;
  assign po025 = ~pi003 & new_n521_;
  assign new_n523_ = pi011 & ~pi054;
  assign new_n524_ = ~pi011 & new_n449_;
  assign new_n525_ = new_n448_ & new_n524_;
  assign new_n526_ = new_n503_ & new_n525_;
  assign new_n527_ = ~pi010 & pi022;
  assign new_n528_ = new_n416_ & new_n527_;
  assign new_n529_ = new_n369_ & new_n528_;
  assign new_n530_ = new_n526_ & new_n529_;
  assign new_n531_ = ~new_n523_ & ~new_n530_;
  assign new_n532_ = ~pi129 & ~new_n531_;
  assign po026 = ~pi003 & new_n532_;
  assign new_n534_ = pi012 & ~pi054;
  assign new_n535_ = ~pi012 & new_n449_;
  assign new_n536_ = new_n448_ & new_n535_;
  assign new_n537_ = pi018 & new_n295_;
  assign new_n538_ = new_n536_ & new_n537_;
  assign new_n539_ = ~pi011 & new_n418_;
  assign new_n540_ = new_n538_ & new_n539_;
  assign new_n541_ = ~new_n534_ & ~new_n540_;
  assign new_n542_ = ~pi129 & ~new_n541_;
  assign po027 = ~pi003 & new_n542_;
  assign new_n544_ = pi013 & ~pi054;
  assign new_n545_ = ~pi013 & new_n450_;
  assign new_n546_ = new_n448_ & new_n545_;
  assign new_n547_ = new_n447_ & new_n546_;
  assign new_n548_ = ~pi025 & pi029;
  assign new_n549_ = ~pi028 & new_n548_;
  assign new_n550_ = new_n357_ & new_n549_;
  assign new_n551_ = ~pi007 & new_n417_;
  assign new_n552_ = new_n550_ & new_n551_;
  assign new_n553_ = new_n547_ & new_n552_;
  assign new_n554_ = ~new_n544_ & ~new_n553_;
  assign new_n555_ = ~pi129 & ~new_n554_;
  assign po028 = ~pi003 & new_n555_;
  assign new_n557_ = pi014 & ~pi054;
  assign new_n558_ = ~pi016 & new_n354_;
  assign new_n559_ = new_n449_ & new_n558_;
  assign new_n560_ = new_n503_ & new_n559_;
  assign new_n561_ = ~pi009 & pi013;
  assign new_n562_ = new_n344_ & new_n561_;
  assign new_n563_ = new_n515_ & new_n562_;
  assign new_n564_ = new_n560_ & new_n563_;
  assign new_n565_ = ~new_n557_ & ~new_n564_;
  assign new_n566_ = ~pi129 & ~new_n565_;
  assign po029 = ~pi003 & new_n566_;
  assign new_n568_ = ~pi041 & ~pi043;
  assign new_n569_ = new_n399_ & new_n568_;
  assign new_n570_ = ~pi045 & new_n384_;
  assign new_n571_ = new_n569_ & new_n570_;
  assign new_n572_ = ~pi046 & new_n388_;
  assign new_n573_ = new_n391_ & new_n572_;
  assign new_n574_ = ~pi015 & new_n573_;
  assign new_n575_ = new_n571_ & new_n574_;
  assign new_n576_ = pi082 & ~new_n575_;
  assign new_n577_ = ~new_n379_ & ~new_n576_;
  assign new_n578_ = ~pi070 & new_n577_;
  assign new_n579_ = ~pi048 & new_n381_;
  assign new_n580_ = new_n570_ & new_n579_;
  assign new_n581_ = new_n407_ & new_n580_;
  assign new_n582_ = pi015 & ~new_n581_;
  assign new_n583_ = ~pi045 & new_n399_;
  assign new_n584_ = ~pi002 & ~pi020;
  assign new_n585_ = ~pi015 & ~new_n584_;
  assign new_n586_ = new_n408_ & new_n585_;
  assign new_n587_ = new_n384_ & new_n586_;
  assign new_n588_ = new_n583_ & new_n587_;
  assign new_n589_ = ~new_n582_ & ~new_n588_;
  assign new_n590_ = pi082 & ~new_n589_;
  assign new_n591_ = pi015 & new_n411_;
  assign new_n592_ = ~new_n590_ & ~new_n591_;
  assign new_n593_ = ~new_n578_ & new_n592_;
  assign po030 = ~pi129 & ~new_n593_;
  assign new_n595_ = pi016 & ~pi054;
  assign new_n596_ = pi006 & ~pi012;
  assign new_n597_ = ~pi005 & new_n596_;
  assign new_n598_ = new_n345_ & new_n597_;
  assign new_n599_ = new_n417_ & new_n598_;
  assign new_n600_ = new_n434_ & new_n599_;
  assign new_n601_ = ~new_n595_ & ~new_n600_;
  assign new_n602_ = ~pi129 & ~new_n601_;
  assign po031 = ~pi003 & new_n602_;
  assign new_n604_ = pi017 & ~pi054;
  assign new_n605_ = ~pi007 & new_n346_;
  assign new_n606_ = ~pi025 & ~pi028;
  assign new_n607_ = ~pi012 & new_n606_;
  assign new_n608_ = new_n605_ & new_n607_;
  assign new_n609_ = new_n445_ & new_n608_;
  assign new_n610_ = ~pi016 & new_n351_;
  assign new_n611_ = new_n450_ & new_n610_;
  assign new_n612_ = ~pi011 & new_n311_;
  assign new_n613_ = ~pi029 & pi059;
  assign new_n614_ = new_n612_ & new_n613_;
  assign new_n615_ = new_n611_ & new_n614_;
  assign new_n616_ = new_n609_ & new_n615_;
  assign new_n617_ = ~new_n604_ & ~new_n616_;
  assign new_n618_ = ~pi129 & ~new_n617_;
  assign po032 = ~pi003 & new_n618_;
  assign new_n620_ = pi018 & ~pi054;
  assign new_n621_ = pi016 & pi054;
  assign new_n622_ = new_n450_ & new_n621_;
  assign new_n623_ = new_n356_ & new_n622_;
  assign new_n624_ = new_n487_ & new_n623_;
  assign new_n625_ = ~new_n620_ & ~new_n624_;
  assign new_n626_ = ~pi129 & ~new_n625_;
  assign po033 = ~pi003 & new_n626_;
  assign new_n628_ = pi019 & ~pi054;
  assign new_n629_ = pi017 & new_n612_;
  assign new_n630_ = ~pi004 & ~pi018;
  assign new_n631_ = ~pi019 & new_n630_;
  assign new_n632_ = new_n448_ & new_n631_;
  assign new_n633_ = new_n629_ & new_n632_;
  assign new_n634_ = new_n487_ & new_n633_;
  assign new_n635_ = ~new_n628_ & ~new_n634_;
  assign new_n636_ = ~pi129 & ~new_n635_;
  assign po034 = ~pi003 & new_n636_;
  assign new_n638_ = new_n381_ & new_n387_;
  assign new_n639_ = ~pi024 & new_n380_;
  assign new_n640_ = new_n638_ & new_n639_;
  assign new_n641_ = ~pi040 & ~pi042;
  assign new_n642_ = new_n388_ & new_n641_;
  assign new_n643_ = ~pi044 & new_n401_;
  assign new_n644_ = new_n642_ & new_n643_;
  assign new_n645_ = new_n640_ & new_n644_;
  assign new_n646_ = pi082 & ~new_n645_;
  assign new_n647_ = ~new_n379_ & ~new_n646_;
  assign new_n648_ = ~pi071 & new_n647_;
  assign new_n649_ = ~pi050 & new_n403_;
  assign new_n650_ = ~pi015 & ~pi049;
  assign new_n651_ = new_n390_ & new_n650_;
  assign new_n652_ = new_n649_ & new_n651_;
  assign new_n653_ = new_n640_ & new_n652_;
  assign new_n654_ = pi020 & ~new_n653_;
  assign new_n655_ = pi002 & new_n645_;
  assign new_n656_ = ~new_n654_ & ~new_n655_;
  assign new_n657_ = pi082 & ~new_n656_;
  assign new_n658_ = pi020 & new_n411_;
  assign new_n659_ = ~new_n657_ & ~new_n658_;
  assign new_n660_ = ~new_n648_ & new_n659_;
  assign po035 = ~pi129 & ~new_n660_;
  assign new_n662_ = pi021 & ~pi054;
  assign new_n663_ = new_n355_ & new_n488_;
  assign new_n664_ = ~pi021 & pi054;
  assign new_n665_ = pi019 & new_n664_;
  assign new_n666_ = new_n299_ & new_n665_;
  assign new_n667_ = new_n663_ & new_n666_;
  assign new_n668_ = new_n487_ & new_n667_;
  assign new_n669_ = ~new_n662_ & ~new_n668_;
  assign new_n670_ = ~pi129 & ~new_n669_;
  assign po036 = ~pi003 & new_n670_;
  assign new_n672_ = pi022 & ~pi054;
  assign new_n673_ = ~pi022 & new_n449_;
  assign new_n674_ = new_n448_ & new_n673_;
  assign new_n675_ = new_n503_ & new_n674_;
  assign new_n676_ = ~pi009 & ~pi010;
  assign new_n677_ = new_n291_ & new_n676_;
  assign new_n678_ = pi005 & ~pi007;
  assign new_n679_ = new_n479_ & new_n678_;
  assign new_n680_ = new_n677_ & new_n679_;
  assign new_n681_ = new_n675_ & new_n680_;
  assign new_n682_ = ~new_n672_ & ~new_n681_;
  assign new_n683_ = ~pi129 & ~new_n682_;
  assign po037 = ~pi003 & new_n683_;
  assign new_n685_ = ~pi023 & pi055;
  assign new_n686_ = ~pi129 & ~new_n685_;
  assign po038 = pi061 & new_n686_;
  assign new_n688_ = ~pi047 & new_n568_;
  assign new_n689_ = new_n380_ & new_n688_;
  assign new_n690_ = new_n573_ & new_n689_;
  assign new_n691_ = pi082 & ~new_n690_;
  assign new_n692_ = new_n584_ & new_n650_;
  assign new_n693_ = pi082 & ~new_n692_;
  assign new_n694_ = new_n379_ & ~new_n693_;
  assign new_n695_ = ~new_n691_ & ~new_n694_;
  assign new_n696_ = ~pi024 & ~new_n695_;
  assign new_n697_ = ~pi002 & ~pi045;
  assign new_n698_ = new_n399_ & new_n697_;
  assign new_n699_ = new_n401_ & new_n698_;
  assign new_n700_ = new_n408_ & new_n699_;
  assign new_n701_ = pi082 & ~new_n700_;
  assign new_n702_ = ~new_n379_ & ~new_n701_;
  assign new_n703_ = pi063 & new_n702_;
  assign new_n704_ = ~pi043 & new_n387_;
  assign new_n705_ = new_n583_ & new_n704_;
  assign new_n706_ = pi024 & pi082;
  assign new_n707_ = new_n390_ & new_n706_;
  assign new_n708_ = new_n649_ & new_n707_;
  assign new_n709_ = new_n705_ & new_n708_;
  assign new_n710_ = ~pi129 & ~new_n709_;
  assign new_n711_ = ~new_n703_ & new_n710_;
  assign po039 = ~new_n696_ & new_n711_;
  assign new_n713_ = pi085 & pi116;
  assign new_n714_ = ~pi085 & ~pi110;
  assign new_n715_ = ~pi096 & new_n714_;
  assign new_n716_ = ~new_n713_ & ~new_n715_;
  assign new_n717_ = pi100 & ~new_n716_;
  assign new_n718_ = pi025 & ~pi116;
  assign new_n719_ = pi085 & new_n718_;
  assign new_n720_ = ~new_n717_ & ~new_n719_;
  assign new_n721_ = ~pi026 & ~new_n720_;
  assign new_n722_ = ~pi051 & ~pi052;
  assign new_n723_ = ~pi039 & new_n722_;
  assign new_n724_ = ~pi095 & ~pi100;
  assign new_n725_ = ~pi097 & new_n724_;
  assign new_n726_ = ~pi110 & ~new_n725_;
  assign new_n727_ = pi025 & ~new_n726_;
  assign new_n728_ = pi026 & pi116;
  assign new_n729_ = ~new_n727_ & ~new_n728_;
  assign new_n730_ = ~new_n723_ & ~new_n729_;
  assign new_n731_ = pi026 & new_n718_;
  assign new_n732_ = ~new_n730_ & ~new_n731_;
  assign new_n733_ = ~pi085 & ~new_n732_;
  assign new_n734_ = ~new_n721_ & ~new_n733_;
  assign new_n735_ = ~pi027 & ~new_n734_;
  assign new_n736_ = ~pi039 & ~pi052;
  assign new_n737_ = ~pi051 & new_n736_;
  assign new_n738_ = pi116 & new_n737_;
  assign new_n739_ = ~new_n718_ & ~new_n738_;
  assign new_n740_ = pi027 & ~new_n739_;
  assign new_n741_ = new_n723_ & new_n727_;
  assign new_n742_ = ~new_n740_ & ~new_n741_;
  assign new_n743_ = ~pi026 & ~pi085;
  assign new_n744_ = ~new_n742_ & new_n743_;
  assign new_n745_ = ~new_n735_ & ~new_n744_;
  assign new_n746_ = ~pi053 & ~new_n745_;
  assign new_n747_ = pi025 & ~pi026;
  assign new_n748_ = ~pi116 & new_n747_;
  assign new_n749_ = pi053 & ~pi085;
  assign new_n750_ = ~pi027 & new_n749_;
  assign new_n751_ = new_n748_ & new_n750_;
  assign new_n752_ = ~new_n746_ & ~new_n751_;
  assign new_n753_ = ~pi058 & ~new_n752_;
  assign new_n754_ = ~pi027 & ~pi085;
  assign new_n755_ = ~pi053 & pi058;
  assign new_n756_ = new_n754_ & new_n755_;
  assign new_n757_ = new_n748_ & new_n756_;
  assign new_n758_ = ~new_n753_ & ~new_n757_;
  assign new_n759_ = ~pi129 & ~new_n758_;
  assign po040 = ~pi003 & new_n759_;
  assign new_n761_ = pi085 & ~pi116;
  assign new_n762_ = ~pi110 & ~new_n761_;
  assign new_n763_ = ~new_n728_ & new_n762_;
  assign new_n764_ = ~pi096 & new_n763_;
  assign new_n765_ = ~pi026 & new_n713_;
  assign new_n766_ = ~new_n764_ & ~new_n765_;
  assign new_n767_ = pi100 & ~new_n766_;
  assign new_n768_ = ~pi085 & ~new_n738_;
  assign new_n769_ = pi026 & new_n768_;
  assign new_n770_ = ~new_n767_ & ~new_n769_;
  assign new_n771_ = ~pi129 & ~new_n770_;
  assign new_n772_ = ~pi003 & new_n771_;
  assign new_n773_ = ~pi027 & ~pi053;
  assign new_n774_ = ~pi058 & new_n773_;
  assign po041 = new_n772_ & new_n774_;
  assign new_n776_ = pi095 & ~pi096;
  assign new_n777_ = pi027 & pi116;
  assign new_n778_ = new_n762_ & ~new_n777_;
  assign new_n779_ = new_n776_ & new_n778_;
  assign new_n780_ = ~pi027 & new_n713_;
  assign new_n781_ = ~new_n779_ & ~new_n780_;
  assign new_n782_ = ~pi100 & ~new_n781_;
  assign new_n783_ = pi027 & new_n768_;
  assign new_n784_ = ~new_n782_ & ~new_n783_;
  assign new_n785_ = ~pi129 & ~new_n784_;
  assign new_n786_ = ~pi003 & new_n785_;
  assign new_n787_ = ~pi053 & ~pi058;
  assign new_n788_ = ~pi026 & new_n787_;
  assign po042 = new_n786_ & new_n788_;
  assign new_n790_ = ~pi026 & ~new_n723_;
  assign new_n791_ = ~pi027 & new_n737_;
  assign new_n792_ = ~new_n790_ & ~new_n791_;
  assign new_n793_ = ~new_n726_ & ~new_n792_;
  assign new_n794_ = pi026 & ~pi027;
  assign new_n795_ = ~pi026 & pi027;
  assign new_n796_ = ~new_n794_ & ~new_n795_;
  assign new_n797_ = ~pi116 & ~new_n796_;
  assign new_n798_ = ~new_n793_ & ~new_n797_;
  assign new_n799_ = pi028 & ~new_n798_;
  assign new_n800_ = ~pi026 & ~pi100;
  assign new_n801_ = ~pi110 & new_n800_;
  assign new_n802_ = new_n776_ & new_n801_;
  assign new_n803_ = new_n728_ & new_n737_;
  assign new_n804_ = ~new_n802_ & ~new_n803_;
  assign new_n805_ = ~pi027 & ~new_n804_;
  assign new_n806_ = new_n777_ & new_n790_;
  assign new_n807_ = ~new_n805_ & ~new_n806_;
  assign new_n808_ = ~new_n799_ & new_n807_;
  assign new_n809_ = ~pi085 & ~new_n808_;
  assign new_n810_ = pi028 & ~pi116;
  assign new_n811_ = ~pi100 & pi116;
  assign new_n812_ = ~new_n810_ & ~new_n811_;
  assign new_n813_ = pi085 & ~new_n812_;
  assign new_n814_ = ~pi026 & ~pi027;
  assign new_n815_ = new_n813_ & new_n814_;
  assign new_n816_ = ~new_n809_ & ~new_n815_;
  assign new_n817_ = ~pi053 & ~new_n816_;
  assign new_n818_ = ~pi027 & pi028;
  assign new_n819_ = ~pi116 & new_n818_;
  assign new_n820_ = ~pi026 & new_n749_;
  assign new_n821_ = new_n819_ & new_n820_;
  assign new_n822_ = ~new_n817_ & ~new_n821_;
  assign new_n823_ = ~pi058 & ~new_n822_;
  assign new_n824_ = new_n743_ & new_n755_;
  assign new_n825_ = new_n819_ & new_n824_;
  assign new_n826_ = ~new_n823_ & ~new_n825_;
  assign new_n827_ = ~pi129 & ~new_n826_;
  assign po043 = ~pi003 & new_n827_;
  assign new_n829_ = pi029 & pi110;
  assign new_n830_ = pi097 & ~pi110;
  assign new_n831_ = ~pi096 & new_n830_;
  assign new_n832_ = pi029 & ~pi097;
  assign new_n833_ = ~new_n831_ & ~new_n832_;
  assign new_n834_ = new_n724_ & ~new_n833_;
  assign new_n835_ = ~new_n829_ & ~new_n834_;
  assign new_n836_ = ~pi058 & ~new_n835_;
  assign new_n837_ = pi097 & pi116;
  assign new_n838_ = pi029 & ~pi116;
  assign new_n839_ = ~new_n837_ & ~new_n838_;
  assign new_n840_ = pi058 & ~new_n839_;
  assign new_n841_ = ~new_n836_ & ~new_n840_;
  assign new_n842_ = ~pi053 & ~new_n841_;
  assign new_n843_ = pi053 & ~pi058;
  assign new_n844_ = new_n838_ & new_n843_;
  assign new_n845_ = ~new_n842_ & ~new_n844_;
  assign new_n846_ = ~pi027 & ~new_n845_;
  assign new_n847_ = pi027 & new_n838_;
  assign new_n848_ = new_n787_ & new_n847_;
  assign new_n849_ = ~new_n846_ & ~new_n848_;
  assign new_n850_ = ~pi085 & ~new_n849_;
  assign new_n851_ = pi085 & new_n774_;
  assign new_n852_ = new_n838_ & new_n851_;
  assign new_n853_ = ~new_n850_ & ~new_n852_;
  assign new_n854_ = ~pi026 & ~new_n853_;
  assign new_n855_ = new_n754_ & new_n787_;
  assign new_n856_ = pi026 & new_n855_;
  assign new_n857_ = new_n838_ & new_n856_;
  assign new_n858_ = ~new_n854_ & ~new_n857_;
  assign new_n859_ = ~pi129 & ~new_n858_;
  assign po044 = ~pi003 & new_n859_;
  assign new_n861_ = pi030 & ~pi109;
  assign new_n862_ = pi060 & pi109;
  assign new_n863_ = ~new_n861_ & ~new_n862_;
  assign new_n864_ = ~pi106 & ~new_n863_;
  assign new_n865_ = pi088 & pi106;
  assign new_n866_ = ~new_n864_ & ~new_n865_;
  assign po045 = ~pi129 & ~new_n866_;
  assign new_n868_ = pi089 & pi106;
  assign new_n869_ = pi030 & pi109;
  assign new_n870_ = pi031 & ~pi109;
  assign new_n871_ = ~new_n869_ & ~new_n870_;
  assign new_n872_ = ~pi106 & ~new_n871_;
  assign new_n873_ = ~new_n868_ & ~new_n872_;
  assign po046 = ~pi129 & ~new_n873_;
  assign new_n875_ = pi099 & pi106;
  assign new_n876_ = pi031 & pi109;
  assign new_n877_ = pi032 & ~pi109;
  assign new_n878_ = ~new_n876_ & ~new_n877_;
  assign new_n879_ = ~pi106 & ~new_n878_;
  assign new_n880_ = ~new_n875_ & ~new_n879_;
  assign po047 = ~pi129 & ~new_n880_;
  assign new_n882_ = pi090 & pi106;
  assign new_n883_ = pi032 & pi109;
  assign new_n884_ = pi033 & ~pi109;
  assign new_n885_ = ~new_n883_ & ~new_n884_;
  assign new_n886_ = ~pi106 & ~new_n885_;
  assign new_n887_ = ~new_n882_ & ~new_n886_;
  assign po048 = ~pi129 & ~new_n887_;
  assign new_n889_ = pi091 & pi106;
  assign new_n890_ = pi033 & pi109;
  assign new_n891_ = pi034 & ~pi109;
  assign new_n892_ = ~new_n890_ & ~new_n891_;
  assign new_n893_ = ~pi106 & ~new_n892_;
  assign new_n894_ = ~new_n889_ & ~new_n893_;
  assign po049 = ~pi129 & ~new_n894_;
  assign new_n896_ = pi092 & pi106;
  assign new_n897_ = pi034 & pi109;
  assign new_n898_ = pi035 & ~pi109;
  assign new_n899_ = ~new_n897_ & ~new_n898_;
  assign new_n900_ = ~pi106 & ~new_n899_;
  assign new_n901_ = ~new_n896_ & ~new_n900_;
  assign po050 = ~pi129 & ~new_n901_;
  assign new_n903_ = pi098 & pi106;
  assign new_n904_ = pi035 & pi109;
  assign new_n905_ = pi036 & ~pi109;
  assign new_n906_ = ~new_n904_ & ~new_n905_;
  assign new_n907_ = ~pi106 & ~new_n906_;
  assign new_n908_ = ~new_n903_ & ~new_n907_;
  assign po051 = ~pi129 & ~new_n908_;
  assign new_n910_ = pi093 & pi106;
  assign new_n911_ = pi036 & pi109;
  assign new_n912_ = pi037 & ~pi109;
  assign new_n913_ = ~new_n911_ & ~new_n912_;
  assign new_n914_ = ~pi106 & ~new_n913_;
  assign new_n915_ = ~new_n910_ & ~new_n914_;
  assign po052 = ~pi129 & ~new_n915_;
  assign new_n917_ = pi082 & ~new_n391_;
  assign new_n918_ = new_n406_ & new_n579_;
  assign new_n919_ = new_n385_ & new_n697_;
  assign new_n920_ = new_n918_ & new_n919_;
  assign new_n921_ = pi082 & ~new_n920_;
  assign new_n922_ = new_n379_ & ~new_n921_;
  assign new_n923_ = ~new_n917_ & ~new_n922_;
  assign new_n924_ = ~pi038 & ~new_n923_;
  assign new_n925_ = ~pi002 & ~pi048;
  assign new_n926_ = new_n398_ & new_n925_;
  assign new_n927_ = new_n401_ & new_n926_;
  assign new_n928_ = ~pi050 & new_n391_;
  assign new_n929_ = new_n638_ & new_n928_;
  assign new_n930_ = new_n927_ & new_n929_;
  assign new_n931_ = pi082 & ~new_n930_;
  assign new_n932_ = ~new_n379_ & ~new_n931_;
  assign new_n933_ = pi074 & new_n932_;
  assign new_n934_ = ~pi044 & pi082;
  assign new_n935_ = pi038 & new_n641_;
  assign new_n936_ = new_n934_ & new_n935_;
  assign new_n937_ = ~pi129 & ~new_n936_;
  assign new_n938_ = ~new_n933_ & new_n937_;
  assign po053 = ~new_n924_ & new_n938_;
  assign new_n940_ = ~pi051 & pi109;
  assign new_n941_ = new_n736_ & new_n940_;
  assign new_n942_ = ~pi106 & ~new_n941_;
  assign new_n943_ = pi109 & new_n722_;
  assign new_n944_ = pi039 & ~new_n943_;
  assign new_n945_ = new_n942_ & ~new_n944_;
  assign po054 = ~pi129 & ~new_n945_;
  assign new_n947_ = pi082 & ~new_n390_;
  assign new_n948_ = new_n579_ & new_n919_;
  assign new_n949_ = new_n389_ & new_n948_;
  assign new_n950_ = pi082 & ~new_n949_;
  assign new_n951_ = new_n379_ & ~new_n950_;
  assign new_n952_ = ~new_n947_ & ~new_n951_;
  assign new_n953_ = ~pi040 & ~new_n952_;
  assign new_n954_ = new_n388_ & new_n390_;
  assign new_n955_ = new_n638_ & new_n954_;
  assign new_n956_ = new_n927_ & new_n955_;
  assign new_n957_ = pi082 & ~new_n956_;
  assign new_n958_ = ~new_n379_ & ~new_n957_;
  assign new_n959_ = pi073 & new_n958_;
  assign new_n960_ = pi040 & pi082;
  assign new_n961_ = new_n390_ & new_n960_;
  assign new_n962_ = ~pi129 & ~new_n961_;
  assign new_n963_ = ~new_n959_ & new_n962_;
  assign po055 = ~new_n953_ & new_n963_;
  assign new_n965_ = pi082 & ~new_n573_;
  assign new_n966_ = pi082 & ~new_n948_;
  assign new_n967_ = new_n379_ & ~new_n966_;
  assign new_n968_ = ~new_n965_ & ~new_n967_;
  assign new_n969_ = ~pi041 & ~new_n968_;
  assign new_n970_ = new_n381_ & new_n405_;
  assign new_n971_ = new_n404_ & new_n970_;
  assign new_n972_ = new_n927_ & new_n971_;
  assign new_n973_ = pi082 & ~new_n972_;
  assign new_n974_ = ~new_n379_ & ~new_n973_;
  assign new_n975_ = pi076 & new_n974_;
  assign new_n976_ = new_n403_ & new_n405_;
  assign new_n977_ = pi041 & pi082;
  assign new_n978_ = new_n390_ & new_n977_;
  assign new_n979_ = new_n976_ & new_n978_;
  assign new_n980_ = ~pi129 & ~new_n979_;
  assign new_n981_ = ~new_n975_ & new_n980_;
  assign po056 = ~new_n969_ & new_n981_;
  assign new_n983_ = pi044 & pi082;
  assign new_n984_ = new_n688_ & new_n976_;
  assign new_n985_ = new_n927_ & new_n984_;
  assign new_n986_ = pi082 & ~new_n985_;
  assign new_n987_ = new_n379_ & ~new_n986_;
  assign new_n988_ = ~new_n983_ & ~new_n987_;
  assign new_n989_ = ~pi042 & ~new_n988_;
  assign new_n990_ = ~pi044 & new_n649_;
  assign new_n991_ = new_n638_ & new_n990_;
  assign new_n992_ = new_n927_ & new_n991_;
  assign new_n993_ = pi082 & ~new_n992_;
  assign new_n994_ = ~new_n379_ & ~new_n993_;
  assign new_n995_ = pi072 & new_n994_;
  assign new_n996_ = pi042 & new_n934_;
  assign new_n997_ = ~pi129 & ~new_n996_;
  assign new_n998_ = ~new_n995_ & new_n997_;
  assign po057 = ~new_n989_ & new_n998_;
  assign new_n1000_ = pi082 & ~new_n407_;
  assign new_n1001_ = new_n385_ & new_n698_;
  assign new_n1002_ = pi082 & ~new_n1001_;
  assign new_n1003_ = new_n379_ & ~new_n1002_;
  assign new_n1004_ = ~new_n1000_ & ~new_n1003_;
  assign new_n1005_ = ~pi043 & ~new_n1004_;
  assign new_n1006_ = ~pi047 & new_n407_;
  assign new_n1007_ = new_n927_ & new_n1006_;
  assign new_n1008_ = pi082 & ~new_n1007_;
  assign new_n1009_ = ~new_n379_ & ~new_n1008_;
  assign new_n1010_ = pi077 & new_n1009_;
  assign new_n1011_ = pi043 & new_n641_;
  assign new_n1012_ = new_n934_ & new_n1011_;
  assign new_n1013_ = new_n389_ & new_n1012_;
  assign new_n1014_ = ~pi129 & ~new_n1013_;
  assign new_n1015_ = ~new_n1010_ & new_n1014_;
  assign po058 = ~new_n1005_ & new_n1015_;
  assign new_n1017_ = new_n638_ & new_n642_;
  assign new_n1018_ = new_n927_ & new_n1017_;
  assign new_n1019_ = pi082 & ~new_n1018_;
  assign new_n1020_ = pi067 & ~new_n379_;
  assign new_n1021_ = ~pi044 & new_n379_;
  assign new_n1022_ = ~new_n1020_ & ~new_n1021_;
  assign new_n1023_ = ~new_n1019_ & ~new_n1022_;
  assign new_n1024_ = ~pi129 & ~new_n983_;
  assign po059 = ~new_n1023_ & new_n1024_;
  assign new_n1026_ = new_n399_ & new_n704_;
  assign new_n1027_ = new_n388_ & new_n391_;
  assign new_n1028_ = new_n1026_ & new_n1027_;
  assign new_n1029_ = pi082 & ~new_n1028_;
  assign new_n1030_ = ~pi024 & new_n692_;
  assign new_n1031_ = pi082 & ~new_n1030_;
  assign new_n1032_ = new_n379_ & ~new_n1031_;
  assign new_n1033_ = ~new_n1029_ & ~new_n1032_;
  assign new_n1034_ = ~pi045 & ~new_n1033_;
  assign new_n1035_ = ~pi002 & new_n399_;
  assign new_n1036_ = new_n385_ & new_n1035_;
  assign new_n1037_ = new_n408_ & new_n1036_;
  assign new_n1038_ = pi082 & ~new_n1037_;
  assign new_n1039_ = ~new_n379_ & ~new_n1038_;
  assign new_n1040_ = pi068 & new_n1039_;
  assign new_n1041_ = ~pi038 & new_n641_;
  assign new_n1042_ = pi045 & new_n1041_;
  assign new_n1043_ = new_n934_ & new_n1042_;
  assign new_n1044_ = new_n918_ & new_n1043_;
  assign new_n1045_ = ~pi129 & ~new_n1044_;
  assign new_n1046_ = ~new_n1040_ & new_n1045_;
  assign po060 = ~new_n1034_ & new_n1046_;
  assign new_n1048_ = pi082 & ~new_n1027_;
  assign new_n1049_ = new_n688_ & new_n927_;
  assign new_n1050_ = pi082 & ~new_n1049_;
  assign new_n1051_ = new_n379_ & ~new_n1050_;
  assign new_n1052_ = ~new_n1048_ & ~new_n1051_;
  assign new_n1053_ = ~pi046 & ~new_n1052_;
  assign new_n1054_ = ~pi050 & new_n404_;
  assign new_n1055_ = new_n1049_ & new_n1054_;
  assign new_n1056_ = pi082 & ~new_n1055_;
  assign new_n1057_ = ~new_n379_ & ~new_n1056_;
  assign new_n1058_ = pi075 & new_n1057_;
  assign new_n1059_ = pi046 & pi082;
  assign new_n1060_ = new_n1054_ & new_n1059_;
  assign new_n1061_ = ~pi129 & ~new_n1060_;
  assign new_n1062_ = ~new_n1058_ & new_n1061_;
  assign po061 = ~new_n1053_ & new_n1062_;
  assign new_n1064_ = pi082 & ~new_n408_;
  assign new_n1065_ = pi082 & ~new_n927_;
  assign new_n1066_ = new_n379_ & ~new_n1065_;
  assign new_n1067_ = ~new_n1064_ & ~new_n1066_;
  assign new_n1068_ = ~pi047 & ~new_n1067_;
  assign new_n1069_ = new_n408_ & new_n927_;
  assign new_n1070_ = pi082 & ~new_n1069_;
  assign new_n1071_ = ~new_n379_ & ~new_n1070_;
  assign new_n1072_ = pi064 & new_n1071_;
  assign new_n1073_ = new_n568_ & new_n572_;
  assign new_n1074_ = pi047 & new_n641_;
  assign new_n1075_ = new_n934_ & new_n1074_;
  assign new_n1076_ = new_n1073_ & new_n1075_;
  assign new_n1077_ = ~pi129 & ~new_n1076_;
  assign new_n1078_ = ~new_n1072_ & new_n1077_;
  assign po062 = ~new_n1068_ & new_n1078_;
  assign new_n1080_ = new_n638_ & new_n1027_;
  assign new_n1081_ = pi082 & ~new_n1080_;
  assign new_n1082_ = pi082 & ~new_n919_;
  assign new_n1083_ = new_n379_ & ~new_n1082_;
  assign new_n1084_ = ~new_n1081_ & ~new_n1083_;
  assign new_n1085_ = ~pi048 & ~new_n1084_;
  assign new_n1086_ = ~pi002 & ~pi047;
  assign new_n1087_ = new_n398_ & new_n401_;
  assign new_n1088_ = new_n1086_ & new_n1087_;
  assign new_n1089_ = new_n408_ & new_n1088_;
  assign new_n1090_ = pi082 & ~new_n1089_;
  assign new_n1091_ = ~new_n379_ & ~new_n1090_;
  assign new_n1092_ = pi062 & new_n1091_;
  assign new_n1093_ = new_n381_ & new_n406_;
  assign new_n1094_ = pi048 & new_n1041_;
  assign new_n1095_ = new_n934_ & new_n1094_;
  assign new_n1096_ = new_n1093_ & new_n1095_;
  assign new_n1097_ = ~pi129 & ~new_n1096_;
  assign new_n1098_ = ~new_n1092_ & new_n1097_;
  assign po063 = ~new_n1085_ & new_n1098_;
  assign new_n1100_ = new_n384_ & new_n1054_;
  assign new_n1101_ = new_n705_ & new_n1100_;
  assign new_n1102_ = pi082 & ~new_n1101_;
  assign new_n1103_ = ~new_n379_ & ~new_n1102_;
  assign new_n1104_ = ~pi069 & new_n1103_;
  assign new_n1105_ = ~pi024 & ~pi042;
  assign new_n1106_ = new_n990_ & new_n1105_;
  assign new_n1107_ = new_n705_ & new_n1106_;
  assign new_n1108_ = pi049 & ~new_n1107_;
  assign new_n1109_ = ~pi002 & new_n383_;
  assign new_n1110_ = new_n1100_ & ~new_n1109_;
  assign new_n1111_ = new_n638_ & new_n1110_;
  assign new_n1112_ = new_n380_ & new_n1111_;
  assign new_n1113_ = ~new_n1108_ & ~new_n1112_;
  assign new_n1114_ = pi082 & ~new_n1113_;
  assign new_n1115_ = pi049 & new_n411_;
  assign new_n1116_ = ~new_n1114_ & ~new_n1115_;
  assign new_n1117_ = ~new_n1104_ & new_n1116_;
  assign po064 = ~pi129 & ~new_n1117_;
  assign new_n1119_ = pi082 & ~new_n404_;
  assign new_n1120_ = new_n704_ & new_n1035_;
  assign new_n1121_ = new_n1087_ & new_n1120_;
  assign new_n1122_ = pi082 & ~new_n1121_;
  assign new_n1123_ = new_n379_ & ~new_n1122_;
  assign new_n1124_ = ~new_n1119_ & ~new_n1123_;
  assign new_n1125_ = ~pi050 & ~new_n1124_;
  assign new_n1126_ = new_n404_ & new_n638_;
  assign new_n1127_ = new_n927_ & new_n1126_;
  assign new_n1128_ = pi082 & ~new_n1127_;
  assign new_n1129_ = ~new_n379_ & ~new_n1128_;
  assign new_n1130_ = pi066 & new_n1129_;
  assign new_n1131_ = pi050 & new_n1041_;
  assign new_n1132_ = new_n934_ & new_n1131_;
  assign new_n1133_ = ~pi129 & ~new_n1132_;
  assign new_n1134_ = ~new_n1130_ & new_n1133_;
  assign po065 = ~new_n1125_ & new_n1134_;
  assign new_n1136_ = pi051 & ~pi109;
  assign new_n1137_ = ~new_n940_ & ~new_n1136_;
  assign new_n1138_ = ~pi106 & new_n1137_;
  assign po066 = ~pi129 & ~new_n1138_;
  assign new_n1140_ = pi052 & ~new_n940_;
  assign new_n1141_ = ~pi106 & ~new_n943_;
  assign new_n1142_ = ~new_n1140_ & new_n1141_;
  assign po067 = ~pi129 & ~new_n1142_;
  assign new_n1144_ = pi058 & pi116;
  assign new_n1145_ = ~pi058 & ~pi110;
  assign new_n1146_ = ~pi096 & new_n1145_;
  assign new_n1147_ = new_n724_ & new_n1146_;
  assign new_n1148_ = ~new_n1144_ & ~new_n1147_;
  assign new_n1149_ = ~pi053 & ~new_n1148_;
  assign new_n1150_ = pi097 & new_n1149_;
  assign new_n1151_ = ~pi116 & new_n843_;
  assign new_n1152_ = ~new_n1150_ & ~new_n1151_;
  assign new_n1153_ = ~pi129 & ~new_n1152_;
  assign new_n1154_ = ~pi003 & new_n1153_;
  assign new_n1155_ = new_n754_ & new_n1154_;
  assign po068 = ~pi026 & new_n1155_;
  assign new_n1157_ = new_n408_ & new_n1001_;
  assign new_n1158_ = pi082 & ~new_n1157_;
  assign new_n1159_ = ~new_n379_ & ~new_n1158_;
  assign po069 = pi129 | new_n1159_;
  assign po129 = pi123 | pi129;
  assign new_n1162_ = pi114 & ~pi122;
  assign po070 = ~po129 & new_n1162_;
  assign new_n1164_ = ~pi026 & pi058;
  assign new_n1165_ = pi026 & ~pi058;
  assign new_n1166_ = pi116 & new_n1165_;
  assign new_n1167_ = ~new_n1164_ & ~new_n1166_;
  assign new_n1168_ = pi094 & ~new_n1167_;
  assign new_n1169_ = pi058 & ~pi116;
  assign new_n1170_ = pi037 & ~pi116;
  assign new_n1171_ = ~new_n1164_ & ~new_n1170_;
  assign new_n1172_ = ~new_n1169_ & ~new_n1171_;
  assign new_n1173_ = ~new_n1168_ & ~new_n1172_;
  assign new_n1174_ = ~pi053 & ~new_n1173_;
  assign new_n1175_ = ~pi026 & pi037;
  assign new_n1176_ = ~pi058 & new_n1175_;
  assign new_n1177_ = ~new_n1174_ & ~new_n1176_;
  assign new_n1178_ = ~pi085 & ~new_n1177_;
  assign new_n1179_ = new_n787_ & new_n1175_;
  assign new_n1180_ = ~new_n1178_ & ~new_n1179_;
  assign new_n1181_ = ~pi027 & ~new_n1180_;
  assign new_n1182_ = ~pi085 & new_n787_;
  assign new_n1183_ = new_n1175_ & new_n1182_;
  assign new_n1184_ = ~new_n1181_ & ~new_n1183_;
  assign new_n1185_ = ~pi129 & ~new_n1184_;
  assign po071 = ~pi003 & new_n1185_;
  assign new_n1187_ = ~pi026 & ~pi053;
  assign new_n1188_ = pi026 & pi053;
  assign new_n1189_ = ~pi085 & ~new_n1188_;
  assign new_n1190_ = ~new_n1187_ & ~new_n1189_;
  assign new_n1191_ = ~pi058 & ~new_n1190_;
  assign new_n1192_ = ~pi085 & new_n1187_;
  assign new_n1193_ = ~pi116 & new_n1192_;
  assign new_n1194_ = ~new_n1191_ & ~new_n1193_;
  assign new_n1195_ = pi057 & ~new_n1194_;
  assign new_n1196_ = pi060 & new_n1144_;
  assign new_n1197_ = new_n1192_ & new_n1196_;
  assign new_n1198_ = ~new_n1195_ & ~new_n1197_;
  assign new_n1199_ = ~pi027 & ~new_n1198_;
  assign new_n1200_ = pi057 & ~pi058;
  assign new_n1201_ = new_n1192_ & new_n1200_;
  assign new_n1202_ = ~new_n1199_ & ~new_n1201_;
  assign new_n1203_ = ~pi129 & ~new_n1202_;
  assign po072 = ~pi003 & new_n1203_;
  assign new_n1205_ = new_n814_ & new_n1169_;
  assign new_n1206_ = pi116 & ~new_n796_;
  assign new_n1207_ = ~pi058 & new_n1206_;
  assign new_n1208_ = new_n737_ & new_n1207_;
  assign new_n1209_ = ~new_n1205_ & ~new_n1208_;
  assign new_n1210_ = ~pi129 & ~new_n1209_;
  assign new_n1211_ = ~pi003 & new_n1210_;
  assign new_n1212_ = ~pi053 & new_n1211_;
  assign po073 = ~pi085 & new_n1212_;
  assign new_n1214_ = ~new_n755_ & ~new_n843_;
  assign new_n1215_ = ~pi116 & ~new_n1214_;
  assign new_n1216_ = ~new_n726_ & new_n787_;
  assign new_n1217_ = ~new_n1215_ & ~new_n1216_;
  assign new_n1218_ = pi059 & ~new_n1217_;
  assign new_n1219_ = new_n726_ & new_n787_;
  assign new_n1220_ = pi096 & new_n1219_;
  assign new_n1221_ = ~new_n1218_ & ~new_n1220_;
  assign new_n1222_ = ~pi085 & ~new_n1221_;
  assign new_n1223_ = pi059 & ~pi116;
  assign new_n1224_ = pi085 & new_n787_;
  assign new_n1225_ = new_n1223_ & new_n1224_;
  assign new_n1226_ = ~new_n1222_ & ~new_n1225_;
  assign new_n1227_ = ~pi027 & ~new_n1226_;
  assign new_n1228_ = pi027 & new_n1182_;
  assign new_n1229_ = new_n1223_ & new_n1228_;
  assign new_n1230_ = ~new_n1227_ & ~new_n1229_;
  assign new_n1231_ = ~pi026 & ~new_n1230_;
  assign new_n1232_ = new_n856_ & new_n1223_;
  assign new_n1233_ = ~new_n1231_ & ~new_n1232_;
  assign new_n1234_ = ~pi129 & ~new_n1233_;
  assign po074 = ~pi003 & new_n1234_;
  assign new_n1236_ = ~pi117 & ~pi122;
  assign new_n1237_ = pi060 & ~new_n1236_;
  assign new_n1238_ = pi123 & new_n1236_;
  assign po075 = new_n1237_ | new_n1238_;
  assign new_n1240_ = ~pi114 & pi123;
  assign new_n1241_ = ~pi122 & new_n1240_;
  assign po076 = ~pi129 & new_n1241_;
  assign new_n1243_ = ~pi137 & ~pi138;
  assign new_n1244_ = pi136 & new_n1243_;
  assign new_n1245_ = pi132 & pi133;
  assign new_n1246_ = pi131 & new_n1245_;
  assign new_n1247_ = new_n1244_ & new_n1246_;
  assign new_n1248_ = pi062 & ~new_n1247_;
  assign new_n1249_ = pi136 & ~pi137;
  assign new_n1250_ = ~pi140 & new_n1249_;
  assign new_n1251_ = ~pi138 & new_n1246_;
  assign new_n1252_ = new_n1250_ & new_n1251_;
  assign new_n1253_ = ~new_n1248_ & ~new_n1252_;
  assign po077 = pi129 | new_n1253_;
  assign new_n1255_ = pi063 & ~new_n1247_;
  assign new_n1256_ = ~pi142 & new_n1249_;
  assign new_n1257_ = new_n1251_ & new_n1256_;
  assign new_n1258_ = ~new_n1255_ & ~new_n1257_;
  assign po078 = pi129 | new_n1258_;
  assign new_n1260_ = pi064 & ~new_n1247_;
  assign new_n1261_ = ~pi139 & new_n1249_;
  assign new_n1262_ = new_n1251_ & new_n1261_;
  assign new_n1263_ = ~new_n1260_ & ~new_n1262_;
  assign po079 = pi129 | new_n1263_;
  assign new_n1265_ = pi065 & ~new_n1247_;
  assign new_n1266_ = ~pi146 & new_n1249_;
  assign new_n1267_ = new_n1251_ & new_n1266_;
  assign new_n1268_ = ~new_n1265_ & ~new_n1267_;
  assign po080 = pi129 | new_n1268_;
  assign new_n1270_ = ~pi136 & ~pi137;
  assign new_n1271_ = new_n1251_ & new_n1270_;
  assign new_n1272_ = pi066 & ~new_n1271_;
  assign new_n1273_ = ~pi143 & new_n1271_;
  assign new_n1274_ = ~new_n1272_ & ~new_n1273_;
  assign po081 = pi129 | new_n1274_;
  assign new_n1276_ = pi067 & ~new_n1271_;
  assign new_n1277_ = ~pi139 & new_n1271_;
  assign new_n1278_ = ~new_n1276_ & ~new_n1277_;
  assign po082 = pi129 | new_n1278_;
  assign new_n1280_ = pi068 & ~new_n1247_;
  assign new_n1281_ = ~pi141 & new_n1249_;
  assign new_n1282_ = new_n1251_ & new_n1281_;
  assign new_n1283_ = ~new_n1280_ & ~new_n1282_;
  assign po083 = pi129 | new_n1283_;
  assign new_n1285_ = pi069 & ~new_n1247_;
  assign new_n1286_ = ~pi143 & new_n1249_;
  assign new_n1287_ = new_n1251_ & new_n1286_;
  assign new_n1288_ = ~new_n1285_ & ~new_n1287_;
  assign po084 = pi129 | new_n1288_;
  assign new_n1290_ = pi070 & ~new_n1247_;
  assign new_n1291_ = ~pi144 & new_n1249_;
  assign new_n1292_ = new_n1251_ & new_n1291_;
  assign new_n1293_ = ~new_n1290_ & ~new_n1292_;
  assign po085 = pi129 | new_n1293_;
  assign new_n1295_ = pi071 & ~new_n1247_;
  assign new_n1296_ = ~pi145 & new_n1249_;
  assign new_n1297_ = new_n1251_ & new_n1296_;
  assign new_n1298_ = ~new_n1295_ & ~new_n1297_;
  assign po086 = pi129 | new_n1298_;
  assign new_n1300_ = pi072 & ~new_n1271_;
  assign new_n1301_ = ~pi140 & new_n1271_;
  assign new_n1302_ = ~new_n1300_ & ~new_n1301_;
  assign po087 = pi129 | new_n1302_;
  assign new_n1304_ = pi073 & ~new_n1271_;
  assign new_n1305_ = ~pi141 & new_n1271_;
  assign new_n1306_ = ~new_n1304_ & ~new_n1305_;
  assign po088 = pi129 | new_n1306_;
  assign new_n1308_ = pi074 & ~new_n1271_;
  assign new_n1309_ = ~pi142 & new_n1271_;
  assign new_n1310_ = ~new_n1308_ & ~new_n1309_;
  assign po089 = pi129 | new_n1310_;
  assign new_n1312_ = pi075 & ~new_n1271_;
  assign new_n1313_ = ~pi144 & new_n1271_;
  assign new_n1314_ = ~new_n1312_ & ~new_n1313_;
  assign po090 = pi129 | new_n1314_;
  assign new_n1316_ = pi076 & ~new_n1271_;
  assign new_n1317_ = ~pi145 & new_n1271_;
  assign new_n1318_ = ~new_n1316_ & ~new_n1317_;
  assign po091 = pi129 | new_n1318_;
  assign new_n1320_ = pi077 & ~new_n1271_;
  assign new_n1321_ = ~pi146 & new_n1271_;
  assign new_n1322_ = ~new_n1320_ & ~new_n1321_;
  assign po092 = pi129 | new_n1322_;
  assign new_n1324_ = ~pi136 & pi137;
  assign new_n1325_ = new_n1251_ & new_n1324_;
  assign new_n1326_ = pi078 & ~new_n1325_;
  assign new_n1327_ = pi142 & new_n1325_;
  assign new_n1328_ = ~new_n1326_ & ~new_n1327_;
  assign po093 = ~pi129 & ~new_n1328_;
  assign new_n1330_ = pi079 & ~new_n1325_;
  assign new_n1331_ = pi143 & new_n1325_;
  assign new_n1332_ = ~new_n1330_ & ~new_n1331_;
  assign po094 = ~pi129 & ~new_n1332_;
  assign new_n1334_ = pi080 & ~new_n1325_;
  assign new_n1335_ = pi144 & new_n1325_;
  assign new_n1336_ = ~new_n1334_ & ~new_n1335_;
  assign po095 = ~pi129 & ~new_n1336_;
  assign new_n1338_ = pi081 & ~new_n1325_;
  assign new_n1339_ = pi145 & new_n1325_;
  assign new_n1340_ = ~new_n1338_ & ~new_n1339_;
  assign po096 = ~pi129 & ~new_n1340_;
  assign new_n1342_ = pi082 & ~new_n1325_;
  assign new_n1343_ = pi146 & new_n1325_;
  assign new_n1344_ = ~new_n1342_ & ~new_n1343_;
  assign po097 = ~pi129 & ~new_n1344_;
  assign new_n1346_ = pi089 & pi138;
  assign new_n1347_ = ~pi062 & ~pi138;
  assign new_n1348_ = ~new_n1346_ & ~new_n1347_;
  assign new_n1349_ = pi136 & ~new_n1348_;
  assign new_n1350_ = pi119 & pi138;
  assign new_n1351_ = ~pi072 & ~pi138;
  assign new_n1352_ = ~new_n1350_ & ~new_n1351_;
  assign new_n1353_ = ~pi136 & ~new_n1352_;
  assign new_n1354_ = ~new_n1349_ & ~new_n1353_;
  assign new_n1355_ = ~pi137 & ~new_n1354_;
  assign new_n1356_ = ~pi115 & pi138;
  assign new_n1357_ = pi087 & ~pi138;
  assign new_n1358_ = ~new_n1356_ & ~new_n1357_;
  assign new_n1359_ = ~pi136 & ~new_n1358_;
  assign new_n1360_ = pi136 & ~pi138;
  assign new_n1361_ = pi031 & new_n1360_;
  assign new_n1362_ = ~new_n1359_ & ~new_n1361_;
  assign new_n1363_ = pi137 & ~new_n1362_;
  assign po098 = new_n1355_ | new_n1363_;
  assign new_n1365_ = pi084 & ~new_n1325_;
  assign new_n1366_ = pi141 & new_n1325_;
  assign new_n1367_ = ~new_n1365_ & ~new_n1366_;
  assign po099 = ~pi129 & ~new_n1367_;
  assign new_n1369_ = ~pi085 & ~new_n725_;
  assign new_n1370_ = ~pi110 & new_n1369_;
  assign new_n1371_ = pi096 & new_n1370_;
  assign new_n1372_ = ~new_n761_ & ~new_n1371_;
  assign new_n1373_ = ~pi129 & ~new_n1372_;
  assign new_n1374_ = ~pi003 & new_n1373_;
  assign new_n1375_ = new_n774_ & new_n1374_;
  assign po100 = ~pi026 & new_n1375_;
  assign new_n1377_ = pi086 & ~new_n1325_;
  assign new_n1378_ = pi139 & new_n1325_;
  assign new_n1379_ = ~new_n1377_ & ~new_n1378_;
  assign po101 = ~pi129 & ~new_n1379_;
  assign new_n1381_ = pi087 & ~new_n1325_;
  assign new_n1382_ = pi140 & new_n1325_;
  assign new_n1383_ = ~new_n1381_ & ~new_n1382_;
  assign po102 = ~pi129 & ~new_n1383_;
  assign new_n1385_ = pi136 & pi137;
  assign new_n1386_ = new_n1251_ & new_n1385_;
  assign new_n1387_ = pi088 & ~new_n1386_;
  assign new_n1388_ = pi139 & new_n1386_;
  assign new_n1389_ = ~new_n1387_ & ~new_n1388_;
  assign po103 = ~pi129 & ~new_n1389_;
  assign new_n1391_ = pi089 & ~new_n1386_;
  assign new_n1392_ = pi140 & new_n1386_;
  assign new_n1393_ = ~new_n1391_ & ~new_n1392_;
  assign po104 = ~pi129 & ~new_n1393_;
  assign new_n1395_ = pi090 & ~new_n1386_;
  assign new_n1396_ = pi142 & new_n1386_;
  assign new_n1397_ = ~new_n1395_ & ~new_n1396_;
  assign po105 = ~pi129 & ~new_n1397_;
  assign new_n1399_ = pi091 & ~new_n1386_;
  assign new_n1400_ = pi143 & new_n1386_;
  assign new_n1401_ = ~new_n1399_ & ~new_n1400_;
  assign po106 = ~pi129 & ~new_n1401_;
  assign new_n1403_ = pi092 & ~new_n1386_;
  assign new_n1404_ = pi144 & new_n1386_;
  assign new_n1405_ = ~new_n1403_ & ~new_n1404_;
  assign po107 = ~pi129 & ~new_n1405_;
  assign new_n1407_ = pi093 & ~new_n1386_;
  assign new_n1408_ = pi146 & new_n1386_;
  assign new_n1409_ = ~new_n1407_ & ~new_n1408_;
  assign po108 = ~pi129 & ~new_n1409_;
  assign new_n1411_ = pi082 & ~pi137;
  assign new_n1412_ = ~pi136 & new_n1411_;
  assign new_n1413_ = pi138 & new_n1246_;
  assign new_n1414_ = new_n1412_ & new_n1413_;
  assign new_n1415_ = pi094 & ~new_n1414_;
  assign new_n1416_ = pi142 & new_n1414_;
  assign new_n1417_ = ~new_n1415_ & ~new_n1416_;
  assign po109 = ~pi129 & ~new_n1417_;
  assign new_n1419_ = ~pi003 & ~new_n1246_;
  assign new_n1420_ = ~pi110 & new_n1419_;
  assign new_n1421_ = pi138 & new_n1412_;
  assign new_n1422_ = new_n1246_ & ~new_n1421_;
  assign new_n1423_ = ~new_n1420_ & ~new_n1422_;
  assign new_n1424_ = pi095 & ~new_n1423_;
  assign new_n1425_ = pi143 & new_n1414_;
  assign new_n1426_ = ~new_n1424_ & ~new_n1425_;
  assign po110 = ~pi129 & ~new_n1426_;
  assign new_n1428_ = pi096 & ~new_n1423_;
  assign new_n1429_ = pi146 & new_n1414_;
  assign new_n1430_ = ~new_n1428_ & ~new_n1429_;
  assign po111 = ~pi129 & ~new_n1430_;
  assign new_n1432_ = pi097 & ~new_n1423_;
  assign new_n1433_ = pi145 & new_n1414_;
  assign new_n1434_ = ~new_n1432_ & ~new_n1433_;
  assign po112 = ~pi129 & ~new_n1434_;
  assign new_n1436_ = pi098 & ~new_n1386_;
  assign new_n1437_ = pi145 & new_n1386_;
  assign new_n1438_ = ~new_n1436_ & ~new_n1437_;
  assign po113 = ~pi129 & ~new_n1438_;
  assign new_n1440_ = pi099 & ~new_n1386_;
  assign new_n1441_ = pi141 & new_n1386_;
  assign new_n1442_ = ~new_n1440_ & ~new_n1441_;
  assign po114 = ~pi129 & ~new_n1442_;
  assign new_n1444_ = pi100 & ~new_n1423_;
  assign new_n1445_ = pi144 & new_n1414_;
  assign new_n1446_ = ~new_n1444_ & ~new_n1445_;
  assign po115 = ~pi129 & ~new_n1446_;
  assign new_n1448_ = pi124 & pi138;
  assign new_n1449_ = ~pi077 & ~pi138;
  assign new_n1450_ = ~new_n1448_ & ~new_n1449_;
  assign new_n1451_ = ~pi136 & ~new_n1450_;
  assign new_n1452_ = ~pi065 & ~pi138;
  assign new_n1453_ = pi093 & pi138;
  assign new_n1454_ = ~new_n1452_ & ~new_n1453_;
  assign new_n1455_ = pi136 & ~new_n1454_;
  assign new_n1456_ = ~new_n1451_ & ~new_n1455_;
  assign new_n1457_ = ~pi137 & ~new_n1456_;
  assign new_n1458_ = pi037 & new_n1360_;
  assign new_n1459_ = pi096 & pi138;
  assign new_n1460_ = pi082 & ~pi138;
  assign new_n1461_ = ~new_n1459_ & ~new_n1460_;
  assign new_n1462_ = ~pi136 & ~new_n1461_;
  assign new_n1463_ = ~new_n1458_ & ~new_n1462_;
  assign new_n1464_ = pi137 & ~new_n1463_;
  assign po116 = new_n1457_ | new_n1464_;
  assign new_n1466_ = pi091 & new_n1249_;
  assign new_n1467_ = pi095 & new_n1324_;
  assign new_n1468_ = ~new_n1466_ & ~new_n1467_;
  assign new_n1469_ = pi138 & ~new_n1468_;
  assign new_n1470_ = pi079 & ~pi136;
  assign new_n1471_ = pi034 & pi136;
  assign new_n1472_ = ~new_n1470_ & ~new_n1471_;
  assign new_n1473_ = pi137 & ~new_n1472_;
  assign new_n1474_ = ~pi069 & pi136;
  assign new_n1475_ = ~pi066 & ~pi136;
  assign new_n1476_ = ~new_n1474_ & ~new_n1475_;
  assign new_n1477_ = ~pi137 & ~new_n1476_;
  assign new_n1478_ = ~new_n1473_ & ~new_n1477_;
  assign new_n1479_ = ~pi138 & ~new_n1478_;
  assign po117 = new_n1469_ | new_n1479_;
  assign new_n1481_ = pi090 & new_n1249_;
  assign new_n1482_ = pi094 & new_n1324_;
  assign new_n1483_ = ~new_n1481_ & ~new_n1482_;
  assign new_n1484_ = pi138 & ~new_n1483_;
  assign new_n1485_ = pi078 & ~pi136;
  assign new_n1486_ = pi033 & pi136;
  assign new_n1487_ = ~new_n1485_ & ~new_n1486_;
  assign new_n1488_ = pi137 & ~new_n1487_;
  assign new_n1489_ = ~pi063 & pi136;
  assign new_n1490_ = ~pi074 & ~pi136;
  assign new_n1491_ = ~new_n1489_ & ~new_n1490_;
  assign new_n1492_ = ~pi137 & ~new_n1491_;
  assign new_n1493_ = ~new_n1488_ & ~new_n1492_;
  assign new_n1494_ = ~pi138 & ~new_n1493_;
  assign po118 = new_n1484_ | new_n1494_;
  assign new_n1496_ = pi099 & new_n1249_;
  assign new_n1497_ = ~pi112 & new_n1324_;
  assign new_n1498_ = ~new_n1496_ & ~new_n1497_;
  assign new_n1499_ = pi138 & ~new_n1498_;
  assign new_n1500_ = ~pi068 & pi136;
  assign new_n1501_ = ~pi073 & ~pi136;
  assign new_n1502_ = ~new_n1500_ & ~new_n1501_;
  assign new_n1503_ = ~pi137 & ~new_n1502_;
  assign new_n1504_ = pi084 & ~pi136;
  assign new_n1505_ = pi032 & pi136;
  assign new_n1506_ = ~new_n1504_ & ~new_n1505_;
  assign new_n1507_ = pi137 & ~new_n1506_;
  assign new_n1508_ = ~new_n1503_ & ~new_n1507_;
  assign new_n1509_ = ~pi138 & ~new_n1508_;
  assign po119 = new_n1499_ | new_n1509_;
  assign new_n1511_ = pi092 & pi138;
  assign new_n1512_ = ~pi070 & ~pi138;
  assign new_n1513_ = ~new_n1511_ & ~new_n1512_;
  assign new_n1514_ = pi136 & ~new_n1513_;
  assign new_n1515_ = pi125 & pi138;
  assign new_n1516_ = ~pi075 & ~pi138;
  assign new_n1517_ = ~new_n1515_ & ~new_n1516_;
  assign new_n1518_ = ~pi136 & ~new_n1517_;
  assign new_n1519_ = ~new_n1514_ & ~new_n1518_;
  assign new_n1520_ = ~pi137 & ~new_n1519_;
  assign new_n1521_ = pi080 & ~pi138;
  assign new_n1522_ = pi100 & pi138;
  assign new_n1523_ = ~new_n1521_ & ~new_n1522_;
  assign new_n1524_ = ~pi136 & ~new_n1523_;
  assign new_n1525_ = pi035 & new_n1360_;
  assign new_n1526_ = ~new_n1524_ & ~new_n1525_;
  assign new_n1527_ = pi137 & ~new_n1526_;
  assign po120 = new_n1520_ | new_n1527_;
  assign new_n1529_ = new_n788_ & new_n1370_;
  assign new_n1530_ = ~pi027 & new_n1529_;
  assign new_n1531_ = ~new_n713_ & ~new_n1530_;
  assign new_n1532_ = ~pi129 & ~new_n1531_;
  assign po121 = ~pi003 & new_n1532_;
  assign new_n1534_ = pi098 & pi138;
  assign new_n1535_ = ~pi071 & ~pi138;
  assign new_n1536_ = ~new_n1534_ & ~new_n1535_;
  assign new_n1537_ = pi136 & ~new_n1536_;
  assign new_n1538_ = ~pi076 & ~pi138;
  assign new_n1539_ = pi023 & pi138;
  assign new_n1540_ = ~new_n1538_ & ~new_n1539_;
  assign new_n1541_ = ~pi136 & ~new_n1540_;
  assign new_n1542_ = ~new_n1537_ & ~new_n1541_;
  assign new_n1543_ = ~pi137 & ~new_n1542_;
  assign new_n1544_ = pi036 & new_n1360_;
  assign new_n1545_ = pi081 & ~pi138;
  assign new_n1546_ = pi097 & pi138;
  assign new_n1547_ = ~new_n1545_ & ~new_n1546_;
  assign new_n1548_ = ~pi136 & ~new_n1547_;
  assign new_n1549_ = ~new_n1544_ & ~new_n1548_;
  assign new_n1550_ = pi137 & ~new_n1549_;
  assign po122 = new_n1543_ | new_n1550_;
  assign new_n1552_ = pi088 & pi138;
  assign new_n1553_ = ~pi064 & ~pi138;
  assign new_n1554_ = ~new_n1552_ & ~new_n1553_;
  assign new_n1555_ = pi136 & ~new_n1554_;
  assign new_n1556_ = pi120 & pi138;
  assign new_n1557_ = ~pi067 & ~pi138;
  assign new_n1558_ = ~new_n1556_ & ~new_n1557_;
  assign new_n1559_ = ~pi136 & ~new_n1558_;
  assign new_n1560_ = ~new_n1555_ & ~new_n1559_;
  assign new_n1561_ = ~pi137 & ~new_n1560_;
  assign new_n1562_ = pi086 & ~pi138;
  assign new_n1563_ = pi111 & pi138;
  assign new_n1564_ = ~new_n1562_ & ~new_n1563_;
  assign new_n1565_ = ~pi136 & ~new_n1564_;
  assign new_n1566_ = pi030 & new_n1360_;
  assign new_n1567_ = ~new_n1565_ & ~new_n1566_;
  assign new_n1568_ = pi137 & ~new_n1567_;
  assign po123 = new_n1561_ | new_n1568_;
  assign new_n1570_ = ~new_n737_ & new_n795_;
  assign new_n1571_ = ~new_n794_ & ~new_n1570_;
  assign new_n1572_ = ~pi129 & ~new_n1571_;
  assign new_n1573_ = ~pi003 & new_n1572_;
  assign po124 = pi116 & new_n1573_;
  assign new_n1575_ = ~pi097 & new_n755_;
  assign new_n1576_ = ~new_n843_ & ~new_n1575_;
  assign new_n1577_ = ~pi129 & ~new_n1576_;
  assign new_n1578_ = ~pi003 & new_n1577_;
  assign po125 = pi116 & new_n1578_;
  assign new_n1580_ = pi111 & ~new_n1421_;
  assign new_n1581_ = ~pi136 & pi139;
  assign new_n1582_ = ~pi137 & pi138;
  assign new_n1583_ = pi082 & new_n1582_;
  assign new_n1584_ = new_n1581_ & new_n1583_;
  assign new_n1585_ = ~new_n1580_ & ~new_n1584_;
  assign new_n1586_ = new_n1246_ & ~new_n1585_;
  assign po126 = ~pi129 & new_n1586_;
  assign new_n1588_ = ~pi136 & pi141;
  assign new_n1589_ = new_n1583_ & new_n1588_;
  assign new_n1590_ = ~pi112 & ~new_n1421_;
  assign new_n1591_ = ~new_n1589_ & ~new_n1590_;
  assign new_n1592_ = new_n1246_ & ~new_n1591_;
  assign po127 = ~pi129 & new_n1592_;
  assign new_n1594_ = ~pi054 & ~pi113;
  assign new_n1595_ = ~pi011 & ~pi022;
  assign new_n1596_ = pi054 & ~new_n1595_;
  assign new_n1597_ = ~new_n1594_ & ~new_n1596_;
  assign new_n1598_ = ~pi129 & ~new_n1597_;
  assign po128 = ~pi003 & new_n1598_;
  assign new_n1600_ = ~pi136 & pi140;
  assign new_n1601_ = new_n1583_ & new_n1600_;
  assign new_n1602_ = ~pi115 & ~new_n1421_;
  assign new_n1603_ = ~new_n1601_ & ~new_n1602_;
  assign new_n1604_ = new_n1246_ & ~new_n1603_;
  assign po130 = ~pi129 & new_n1604_;
  assign new_n1606_ = ~pi004 & ~pi012;
  assign new_n1607_ = ~pi007 & ~pi009;
  assign new_n1608_ = new_n1606_ & new_n1607_;
  assign new_n1609_ = ~pi129 & ~new_n1608_;
  assign new_n1610_ = ~pi003 & new_n1609_;
  assign po131 = pi054 & new_n1610_;
  assign po132 = ~pi122 | pi129;
  assign new_n1613_ = ~pi054 & pi118;
  assign new_n1614_ = pi054 & ~pi059;
  assign new_n1615_ = new_n549_ & new_n1614_;
  assign new_n1616_ = ~new_n1613_ & ~new_n1615_;
  assign po133 = ~pi129 & ~new_n1616_;
  assign po134 = ~pi129 & ~new_n724_;
  assign new_n1619_ = ~pi110 & ~pi120;
  assign new_n1620_ = ~pi003 & new_n1619_;
  assign new_n1621_ = ~pi129 & ~new_n1620_;
  assign po135 = ~pi111 & new_n1621_;
  assign new_n1623_ = pi081 & pi120;
  assign po136 = ~pi129 & new_n1623_;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi057 & ~pi129;
  assign new_n1628_ = ~pi096 & pi125;
  assign new_n1629_ = ~pi003 & ~new_n1628_;
  assign po140 = ~pi129 & ~new_n1629_;
  assign new_n1631_ = ~pi126 & pi132;
  assign po141 = pi133 & new_n1631_;
  assign po012 = 1'b1;
  assign po000 = pi108;
  assign po001 = pi083;
  assign po002 = pi104;
  assign po003 = pi103;
  assign po004 = pi102;
  assign po005 = pi105;
  assign po006 = pi107;
  assign po007 = pi101;
  assign po008 = pi126;
  assign po009 = pi121;
  assign po010 = pi001;
  assign po011 = pi000;
  assign po013 = pi130;
  assign po014 = pi128;
endmodule


