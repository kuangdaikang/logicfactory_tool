// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:30 2022

module b3  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
    v30, v31,
    \v32.0 , \v32.1 , \v32.2 , \v32.3 , \v32.4 , \v32.5 , \v32.6 , \v32.7 ,
    \v32.8 , \v32.9 , \v32.10 , \v32.11 , \v32.12 , \v32.13 , \v32.14 ,
    \v32.15 , \v32.16 , \v32.17 , \v32.18 , \v32.19   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28,
    v29, v30, v31;
  output \v32.0 , \v32.1 , \v32.2 , \v32.3 , \v32.4 , \v32.5 , \v32.6 ,
    \v32.7 , \v32.8 , \v32.9 , \v32.10 , \v32.11 , \v32.12 , \v32.13 ,
    \v32.14 , \v32.15 , \v32.16 , \v32.17 , \v32.18 , \v32.19 ;
  wire new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_,
    new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_,
    new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_,
    new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_,
    new_n82_, new_n83_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n345_, new_n346_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n479_, new_n480_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_;
  assign new_n54_ = v17 & v18;
  assign new_n55_ = ~v20 & ~v21;
  assign new_n56_ = ~v18 & new_n55_;
  assign new_n57_ = ~new_n54_ & ~new_n56_;
  assign new_n58_ = v3 & v9;
  assign new_n59_ = ~v4 & ~new_n58_;
  assign new_n60_ = ~new_n57_ & ~new_n59_;
  assign new_n61_ = v27 & new_n60_;
  assign new_n62_ = ~v19 & new_n61_;
  assign new_n63_ = ~v16 & new_n62_;
  assign new_n64_ = v0 & new_n63_;
  assign new_n65_ = ~v7 & v31;
  assign new_n66_ = ~v4 & ~v5;
  assign new_n67_ = ~v2 & new_n66_;
  assign new_n68_ = ~v5 & ~new_n67_;
  assign new_n69_ = ~new_n65_ & ~new_n68_;
  assign new_n70_ = ~v2 & ~v4;
  assign new_n71_ = ~v5 & ~v6;
  assign new_n72_ = new_n70_ & new_n71_;
  assign new_n73_ = ~new_n69_ & ~new_n72_;
  assign new_n74_ = ~v27 & ~new_n73_;
  assign new_n75_ = v3 & new_n74_;
  assign new_n76_ = ~new_n64_ & ~new_n75_;
  assign new_n77_ = ~v25 & ~new_n76_;
  assign new_n78_ = ~v28 & ~new_n73_;
  assign new_n79_ = ~v27 & new_n78_;
  assign new_n80_ = ~v26 & new_n79_;
  assign new_n81_ = v25 & new_n80_;
  assign new_n82_ = v3 & new_n81_;
  assign new_n83_ = ~new_n77_ & ~new_n82_;
  assign \v32.1  = ~v1 & ~new_n83_;
  assign new_n85_ = ~v26 & ~v28;
  assign new_n86_ = v25 & new_n85_;
  assign new_n87_ = v25 & ~new_n86_;
  assign new_n88_ = ~v7 & v23;
  assign new_n89_ = ~v5 & ~new_n88_;
  assign new_n90_ = ~v3 & v5;
  assign new_n91_ = ~new_n89_ & ~new_n90_;
  assign new_n92_ = ~new_n70_ & ~new_n91_;
  assign new_n93_ = v2 & ~v29;
  assign new_n94_ = v4 & ~v30;
  assign new_n95_ = ~new_n93_ & ~new_n94_;
  assign new_n96_ = ~v5 & ~new_n95_;
  assign new_n97_ = ~new_n92_ & ~new_n96_;
  assign new_n98_ = v0 & ~new_n97_;
  assign new_n99_ = v3 & ~new_n73_;
  assign new_n100_ = ~new_n98_ & ~new_n99_;
  assign new_n101_ = ~new_n87_ & ~new_n100_;
  assign new_n102_ = v9 & v29;
  assign new_n103_ = v2 & new_n102_;
  assign new_n104_ = v4 & v30;
  assign new_n105_ = ~new_n103_ & ~new_n104_;
  assign new_n106_ = v23 & ~new_n105_;
  assign new_n107_ = v0 & new_n106_;
  assign new_n108_ = v16 & ~v19;
  assign new_n109_ = v16 & ~new_n108_;
  assign new_n110_ = ~v17 & ~new_n109_;
  assign new_n111_ = ~v0 & new_n110_;
  assign new_n112_ = v17 & ~v19;
  assign new_n113_ = ~v16 & new_n112_;
  assign new_n114_ = ~new_n111_ & ~new_n113_;
  assign new_n115_ = v18 & ~new_n114_;
  assign new_n116_ = v15 & ~v16;
  assign new_n117_ = ~v0 & new_n116_;
  assign new_n118_ = ~v18 & v19;
  assign new_n119_ = ~v17 & new_n118_;
  assign new_n120_ = new_n117_ & new_n119_;
  assign new_n121_ = ~new_n115_ & ~new_n120_;
  assign new_n122_ = v31 & ~new_n121_;
  assign new_n123_ = v6 & new_n122_;
  assign new_n124_ = ~v4 & new_n123_;
  assign new_n125_ = v3 & new_n124_;
  assign new_n126_ = ~v2 & new_n125_;
  assign new_n127_ = ~new_n107_ & ~new_n126_;
  assign new_n128_ = ~v5 & ~new_n127_;
  assign new_n129_ = ~v4 & v6;
  assign new_n130_ = ~v2 & new_n129_;
  assign new_n131_ = ~v5 & ~new_n130_;
  assign new_n132_ = ~v21 & ~new_n131_;
  assign new_n133_ = ~v20 & new_n132_;
  assign new_n134_ = ~v15 & new_n133_;
  assign new_n135_ = v5 & v15;
  assign new_n136_ = ~new_n134_ & ~new_n135_;
  assign new_n137_ = v19 & ~new_n136_;
  assign new_n138_ = ~v18 & new_n137_;
  assign new_n139_ = v5 & v18;
  assign new_n140_ = ~new_n138_ & ~new_n139_;
  assign new_n141_ = ~v16 & ~new_n140_;
  assign new_n142_ = v5 & v16;
  assign new_n143_ = v18 & ~v19;
  assign new_n144_ = new_n142_ & new_n143_;
  assign new_n145_ = ~new_n141_ & ~new_n144_;
  assign new_n146_ = ~v17 & ~new_n145_;
  assign new_n147_ = v22 & ~new_n131_;
  assign new_n148_ = ~v21 & new_n147_;
  assign new_n149_ = ~v20 & new_n148_;
  assign new_n150_ = ~v19 & new_n149_;
  assign new_n151_ = ~v18 & new_n150_;
  assign new_n152_ = ~v16 & new_n151_;
  assign new_n153_ = ~new_n146_ & ~new_n152_;
  assign new_n154_ = ~v0 & ~new_n153_;
  assign new_n155_ = ~v18 & ~v20;
  assign new_n156_ = ~v21 & ~v22;
  assign new_n157_ = new_n155_ & new_n156_;
  assign new_n158_ = ~new_n54_ & ~new_n157_;
  assign new_n159_ = v5 & ~new_n158_;
  assign new_n160_ = new_n130_ & new_n157_;
  assign new_n161_ = ~new_n159_ & ~new_n160_;
  assign new_n162_ = ~v19 & ~new_n161_;
  assign new_n163_ = ~v16 & new_n162_;
  assign new_n164_ = ~new_n154_ & ~new_n163_;
  assign new_n165_ = v31 & ~new_n164_;
  assign new_n166_ = v3 & new_n165_;
  assign new_n167_ = ~new_n128_ & ~new_n166_;
  assign new_n168_ = ~v7 & ~new_n167_;
  assign new_n169_ = ~v3 & ~v4;
  assign new_n170_ = ~v2 & new_n169_;
  assign new_n171_ = ~new_n168_ & ~new_n170_;
  assign new_n172_ = ~v25 & ~new_n171_;
  assign new_n173_ = ~v0 & v24;
  assign new_n174_ = v0 & ~v24;
  assign new_n175_ = ~new_n173_ & ~new_n174_;
  assign new_n176_ = ~v26 & ~new_n175_;
  assign new_n177_ = v25 & new_n176_;
  assign new_n178_ = ~new_n172_ & ~new_n177_;
  assign new_n179_ = ~new_n101_ & new_n178_;
  assign new_n180_ = ~v27 & ~new_n179_;
  assign new_n181_ = v10 & ~v12;
  assign new_n182_ = ~v13 & ~v14;
  assign new_n183_ = new_n181_ & new_n182_;
  assign new_n184_ = ~v9 & ~new_n183_;
  assign new_n185_ = v2 & ~new_n184_;
  assign new_n186_ = ~v4 & ~new_n185_;
  assign new_n187_ = ~v8 & ~new_n186_;
  assign new_n188_ = ~v8 & ~new_n187_;
  assign new_n189_ = v27 & ~new_n188_;
  assign new_n190_ = ~v25 & new_n189_;
  assign new_n191_ = v0 & new_n190_;
  assign new_n192_ = ~new_n180_ & ~new_n191_;
  assign new_n193_ = ~v1 & ~new_n192_;
  assign \v32.2  = v1 | new_n193_;
  assign new_n195_ = ~v9 & ~v10;
  assign new_n196_ = v27 & ~new_n195_;
  assign new_n197_ = ~v25 & new_n196_;
  assign new_n198_ = ~v8 & new_n197_;
  assign new_n199_ = v2 & new_n198_;
  assign new_n200_ = ~v1 & new_n199_;
  assign new_n201_ = v0 & new_n200_;
  assign \v32.3  = v1 | new_n201_;
  assign new_n203_ = ~v17 & v19;
  assign new_n204_ = ~v15 & new_n203_;
  assign new_n205_ = ~v19 & v20;
  assign new_n206_ = ~new_n204_ & ~new_n205_;
  assign new_n207_ = ~v20 & v21;
  assign new_n208_ = ~v19 & new_n207_;
  assign new_n209_ = new_n206_ & ~new_n208_;
  assign new_n210_ = ~v19 & ~v20;
  assign new_n211_ = ~v21 & v22;
  assign new_n212_ = new_n210_ & new_n211_;
  assign new_n213_ = new_n209_ & ~new_n212_;
  assign new_n214_ = ~v0 & ~new_n213_;
  assign new_n215_ = new_n156_ & new_n210_;
  assign new_n216_ = ~new_n214_ & ~new_n215_;
  assign new_n217_ = ~v18 & ~new_n216_;
  assign new_n218_ = ~v16 & new_n217_;
  assign new_n219_ = v5 & ~new_n218_;
  assign new_n220_ = v6 & ~new_n219_;
  assign new_n221_ = ~v4 & new_n220_;
  assign new_n222_ = ~v2 & new_n221_;
  assign new_n223_ = ~v5 & ~new_n222_;
  assign new_n224_ = v31 & ~new_n223_;
  assign new_n225_ = ~v27 & new_n224_;
  assign new_n226_ = ~v25 & new_n225_;
  assign new_n227_ = ~v7 & new_n226_;
  assign new_n228_ = v3 & new_n227_;
  assign new_n229_ = ~v1 & new_n228_;
  assign \v32.4  = v1 | new_n229_;
  assign new_n231_ = ~v1 & v4;
  assign new_n232_ = v0 & new_n231_;
  assign new_n233_ = ~v25 & v27;
  assign new_n234_ = ~v8 & new_n233_;
  assign new_n235_ = new_n232_ & new_n234_;
  assign \v32.5  = v1 | new_n235_;
  assign new_n237_ = v8 & v27;
  assign new_n238_ = v27 & ~new_n237_;
  assign new_n239_ = ~v25 & ~new_n238_;
  assign new_n240_ = v25 & ~v26;
  assign new_n241_ = ~v27 & ~v28;
  assign new_n242_ = new_n240_ & new_n241_;
  assign new_n243_ = ~new_n239_ & ~new_n242_;
  assign new_n244_ = v23 & v29;
  assign new_n245_ = ~v7 & new_n244_;
  assign new_n246_ = ~v5 & ~new_n245_;
  assign new_n247_ = ~new_n90_ & ~new_n246_;
  assign new_n248_ = ~new_n243_ & ~new_n247_;
  assign new_n249_ = v2 & new_n248_;
  assign new_n250_ = ~v1 & new_n249_;
  assign \v32.6  = v0 & new_n250_;
  assign new_n252_ = v0 & ~v1;
  assign new_n253_ = v2 & new_n252_;
  assign new_n254_ = ~v5 & new_n253_;
  assign new_n255_ = ~v7 & new_n254_;
  assign new_n256_ = v23 & new_n255_;
  assign new_n257_ = ~v25 & new_n256_;
  assign new_n258_ = ~v27 & new_n257_;
  assign \v32.7  = v29 & new_n258_;
  assign new_n260_ = v23 & v30;
  assign new_n261_ = ~v7 & new_n260_;
  assign new_n262_ = ~v5 & ~new_n261_;
  assign new_n263_ = ~new_n90_ & ~new_n262_;
  assign new_n264_ = ~new_n243_ & ~new_n263_;
  assign new_n265_ = ~v11 & new_n264_;
  assign new_n266_ = v4 & new_n265_;
  assign new_n267_ = ~v27 & v28;
  assign new_n268_ = ~v26 & new_n267_;
  assign new_n269_ = ~v26 & v27;
  assign new_n270_ = ~v26 & ~new_n269_;
  assign new_n271_ = ~new_n268_ & new_n270_;
  assign new_n272_ = v25 & ~new_n271_;
  assign new_n273_ = ~v24 & new_n272_;
  assign new_n274_ = v10 & new_n233_;
  assign new_n275_ = ~v8 & new_n274_;
  assign new_n276_ = v2 & new_n275_;
  assign new_n277_ = ~new_n273_ & ~new_n276_;
  assign new_n278_ = ~new_n266_ & new_n277_;
  assign new_n279_ = ~v1 & ~new_n278_;
  assign \v32.8  = v0 & new_n279_;
  assign new_n281_ = v27 & ~new_n59_;
  assign new_n282_ = v0 & new_n281_;
  assign new_n283_ = v31 & ~new_n131_;
  assign new_n284_ = ~v27 & new_n283_;
  assign new_n285_ = v22 & new_n284_;
  assign new_n286_ = ~v7 & new_n285_;
  assign new_n287_ = v3 & new_n286_;
  assign new_n288_ = ~v0 & new_n287_;
  assign new_n289_ = ~new_n282_ & ~new_n288_;
  assign new_n290_ = ~v21 & ~new_n289_;
  assign new_n291_ = v21 & new_n284_;
  assign new_n292_ = ~v7 & new_n291_;
  assign new_n293_ = v3 & new_n292_;
  assign new_n294_ = ~v0 & new_n293_;
  assign new_n295_ = ~new_n290_ & ~new_n294_;
  assign new_n296_ = ~v20 & ~new_n295_;
  assign new_n297_ = v20 & new_n283_;
  assign new_n298_ = ~v7 & new_n297_;
  assign new_n299_ = ~v0 & new_n298_;
  assign new_n300_ = ~new_n72_ & ~new_n299_;
  assign new_n301_ = ~new_n69_ & new_n300_;
  assign new_n302_ = ~v27 & ~new_n301_;
  assign new_n303_ = v3 & new_n302_;
  assign new_n304_ = ~new_n296_ & ~new_n303_;
  assign new_n305_ = ~v19 & ~new_n304_;
  assign new_n306_ = ~v20 & ~new_n207_;
  assign new_n307_ = ~v20 & new_n211_;
  assign new_n308_ = new_n306_ & ~new_n307_;
  assign new_n309_ = ~new_n131_ & ~new_n308_;
  assign new_n310_ = v31 & new_n309_;
  assign new_n311_ = ~v7 & new_n310_;
  assign new_n312_ = ~new_n72_ & ~new_n311_;
  assign new_n313_ = ~new_n69_ & new_n312_;
  assign new_n314_ = ~v27 & ~new_n313_;
  assign new_n315_ = v19 & new_n314_;
  assign new_n316_ = ~v17 & new_n315_;
  assign new_n317_ = ~v15 & new_n316_;
  assign new_n318_ = v3 & new_n317_;
  assign new_n319_ = ~v0 & new_n318_;
  assign new_n320_ = ~new_n305_ & ~new_n319_;
  assign new_n321_ = ~v25 & ~new_n320_;
  assign new_n322_ = ~v0 & ~v15;
  assign new_n323_ = new_n203_ & new_n322_;
  assign new_n324_ = v19 & ~new_n323_;
  assign new_n325_ = ~new_n73_ & ~new_n324_;
  assign new_n326_ = ~v28 & new_n325_;
  assign new_n327_ = ~v27 & new_n326_;
  assign new_n328_ = ~v26 & new_n327_;
  assign new_n329_ = v25 & new_n328_;
  assign new_n330_ = v3 & new_n329_;
  assign new_n331_ = ~new_n321_ & ~new_n330_;
  assign new_n332_ = ~v18 & ~new_n331_;
  assign new_n333_ = ~v16 & new_n332_;
  assign new_n334_ = v26 & ~v27;
  assign new_n335_ = ~new_n269_ & ~new_n334_;
  assign new_n336_ = v27 & ~v28;
  assign new_n337_ = v26 & new_n336_;
  assign new_n338_ = ~new_n268_ & ~new_n337_;
  assign new_n339_ = new_n335_ & new_n338_;
  assign new_n340_ = v25 & ~new_n339_;
  assign new_n341_ = v24 & new_n340_;
  assign new_n342_ = ~v0 & new_n341_;
  assign new_n343_ = ~new_n333_ & ~new_n342_;
  assign \v32.9  = ~v1 & ~new_n343_;
  assign new_n345_ = v4 & new_n264_;
  assign new_n346_ = ~v1 & new_n345_;
  assign \v32.10  = v0 & new_n346_;
  assign new_n348_ = ~new_n73_ & ~new_n87_;
  assign new_n349_ = ~v27 & new_n348_;
  assign new_n350_ = v19 & new_n349_;
  assign new_n351_ = v18 & new_n350_;
  assign new_n352_ = ~v17 & new_n351_;
  assign new_n353_ = ~v16 & new_n352_;
  assign new_n354_ = v3 & new_n353_;
  assign new_n355_ = ~v1 & new_n354_;
  assign \v32.11  = ~v0 & new_n355_;
  assign new_n357_ = ~v18 & new_n350_;
  assign new_n358_ = ~v17 & new_n357_;
  assign new_n359_ = ~v16 & new_n358_;
  assign new_n360_ = v15 & new_n359_;
  assign new_n361_ = v3 & new_n360_;
  assign new_n362_ = ~v1 & new_n361_;
  assign \v32.12  = ~v0 & new_n362_;
  assign new_n364_ = v2 & v29;
  assign new_n365_ = ~new_n104_ & ~new_n364_;
  assign new_n366_ = v23 & ~new_n365_;
  assign new_n367_ = v0 & new_n366_;
  assign new_n368_ = ~v2 & v3;
  assign new_n369_ = v6 & v31;
  assign new_n370_ = ~v4 & new_n369_;
  assign new_n371_ = new_n368_ & new_n370_;
  assign new_n372_ = ~new_n367_ & ~new_n371_;
  assign new_n373_ = ~v5 & ~new_n372_;
  assign new_n374_ = v6 & new_n218_;
  assign new_n375_ = ~v4 & new_n374_;
  assign new_n376_ = ~v2 & new_n375_;
  assign new_n377_ = ~v5 & ~new_n376_;
  assign new_n378_ = v31 & ~new_n377_;
  assign new_n379_ = v3 & new_n378_;
  assign new_n380_ = ~new_n373_ & ~new_n379_;
  assign new_n381_ = ~v27 & ~new_n380_;
  assign new_n382_ = ~v7 & new_n381_;
  assign new_n383_ = ~v8 & new_n196_;
  assign new_n384_ = v2 & new_n383_;
  assign new_n385_ = v0 & new_n384_;
  assign new_n386_ = ~new_n382_ & ~new_n385_;
  assign new_n387_ = ~v25 & ~new_n386_;
  assign new_n388_ = v24 & ~v26;
  assign new_n389_ = ~v0 & new_n388_;
  assign new_n390_ = ~new_n174_ & ~new_n389_;
  assign new_n391_ = new_n173_ & new_n334_;
  assign new_n392_ = new_n390_ & ~new_n391_;
  assign new_n393_ = new_n173_ & new_n337_;
  assign new_n394_ = new_n392_ & ~new_n393_;
  assign new_n395_ = v25 & ~new_n394_;
  assign new_n396_ = ~new_n387_ & ~new_n395_;
  assign \v32.13  = ~v1 & ~new_n396_;
  assign new_n398_ = v19 & ~new_n204_;
  assign new_n399_ = ~new_n131_ & ~new_n398_;
  assign new_n400_ = v31 & new_n399_;
  assign new_n401_ = ~v22 & new_n400_;
  assign new_n402_ = v21 & new_n401_;
  assign new_n403_ = ~v7 & new_n402_;
  assign new_n404_ = ~v21 & ~new_n73_;
  assign new_n405_ = v19 & new_n404_;
  assign new_n406_ = ~v17 & new_n405_;
  assign new_n407_ = ~v15 & new_n406_;
  assign new_n408_ = ~new_n403_ & ~new_n407_;
  assign new_n409_ = ~v25 & ~new_n408_;
  assign new_n410_ = ~v26 & new_n78_;
  assign new_n411_ = v25 & new_n410_;
  assign new_n412_ = ~v21 & new_n411_;
  assign new_n413_ = v19 & new_n412_;
  assign new_n414_ = ~v17 & new_n413_;
  assign new_n415_ = ~v15 & new_n414_;
  assign new_n416_ = ~new_n409_ & ~new_n415_;
  assign new_n417_ = ~v20 & ~new_n416_;
  assign new_n418_ = v19 & new_n348_;
  assign new_n419_ = ~v17 & new_n418_;
  assign new_n420_ = v15 & new_n419_;
  assign new_n421_ = ~new_n417_ & ~new_n420_;
  assign new_n422_ = ~v18 & ~new_n421_;
  assign new_n423_ = v18 & new_n348_;
  assign new_n424_ = ~v17 & new_n423_;
  assign new_n425_ = ~new_n422_ & ~new_n424_;
  assign new_n426_ = ~v0 & ~new_n425_;
  assign new_n427_ = ~new_n57_ & ~new_n73_;
  assign new_n428_ = ~new_n87_ & new_n427_;
  assign new_n429_ = ~v19 & new_n428_;
  assign new_n430_ = ~new_n426_ & ~new_n429_;
  assign new_n431_ = ~v16 & ~new_n430_;
  assign new_n432_ = ~v19 & new_n348_;
  assign new_n433_ = v18 & new_n432_;
  assign new_n434_ = ~v17 & new_n433_;
  assign new_n435_ = v16 & new_n434_;
  assign new_n436_ = ~v0 & new_n435_;
  assign new_n437_ = ~new_n431_ & ~new_n436_;
  assign new_n438_ = v3 & ~new_n437_;
  assign new_n439_ = v2 & v9;
  assign new_n440_ = ~v4 & ~new_n439_;
  assign new_n441_ = ~new_n91_ & ~new_n440_;
  assign new_n442_ = v9 & ~v29;
  assign new_n443_ = v2 & new_n442_;
  assign new_n444_ = ~new_n94_ & ~new_n443_;
  assign new_n445_ = ~v5 & ~new_n444_;
  assign new_n446_ = ~new_n441_ & ~new_n445_;
  assign new_n447_ = ~new_n87_ & ~new_n446_;
  assign new_n448_ = v2 & ~v5;
  assign new_n449_ = ~v7 & new_n181_;
  assign new_n450_ = new_n448_ & new_n449_;
  assign new_n451_ = ~v25 & v29;
  assign new_n452_ = v23 & new_n451_;
  assign new_n453_ = new_n182_ & new_n452_;
  assign new_n454_ = new_n450_ & new_n453_;
  assign new_n455_ = ~new_n447_ & ~new_n454_;
  assign new_n456_ = v0 & ~new_n455_;
  assign new_n457_ = ~new_n438_ & ~new_n456_;
  assign new_n458_ = ~v27 & ~new_n457_;
  assign new_n459_ = ~v19 & new_n60_;
  assign new_n460_ = ~v16 & new_n459_;
  assign new_n461_ = v8 & ~new_n446_;
  assign new_n462_ = ~v8 & v10;
  assign new_n463_ = v2 & new_n462_;
  assign new_n464_ = ~v13 & v14;
  assign new_n465_ = ~v12 & new_n464_;
  assign new_n466_ = new_n463_ & new_n465_;
  assign new_n467_ = ~new_n461_ & ~new_n466_;
  assign new_n468_ = ~new_n460_ & new_n467_;
  assign new_n469_ = ~v25 & ~new_n468_;
  assign new_n470_ = ~v24 & v25;
  assign new_n471_ = new_n85_ & new_n470_;
  assign new_n472_ = ~new_n469_ & ~new_n471_;
  assign new_n473_ = v0 & ~new_n472_;
  assign new_n474_ = new_n86_ & new_n173_;
  assign new_n475_ = ~new_n473_ & ~new_n474_;
  assign new_n476_ = v27 & ~new_n475_;
  assign new_n477_ = ~new_n458_ & ~new_n476_;
  assign \v32.14  = ~v1 & ~new_n477_;
  assign new_n479_ = v23 & ~new_n234_;
  assign new_n480_ = ~v1 & new_n479_;
  assign \v32.15  = v0 & new_n480_;
  assign new_n482_ = v24 & new_n272_;
  assign new_n483_ = new_n309_ & ~new_n398_;
  assign new_n484_ = v31 & new_n483_;
  assign new_n485_ = ~v27 & new_n484_;
  assign new_n486_ = ~v25 & new_n485_;
  assign new_n487_ = ~v18 & new_n486_;
  assign new_n488_ = ~v16 & new_n487_;
  assign new_n489_ = ~v7 & new_n488_;
  assign new_n490_ = v3 & new_n489_;
  assign new_n491_ = ~new_n482_ & ~new_n490_;
  assign new_n492_ = ~v1 & ~new_n491_;
  assign \v32.16  = ~v0 & new_n492_;
  assign new_n494_ = v10 & v27;
  assign new_n495_ = ~v8 & new_n494_;
  assign new_n496_ = v2 & new_n495_;
  assign new_n497_ = v0 & new_n496_;
  assign new_n498_ = ~v18 & new_n485_;
  assign new_n499_ = ~v16 & new_n498_;
  assign new_n500_ = ~v7 & new_n499_;
  assign new_n501_ = v3 & new_n500_;
  assign new_n502_ = ~v0 & new_n501_;
  assign new_n503_ = ~new_n497_ & ~new_n502_;
  assign new_n504_ = ~v25 & ~new_n503_;
  assign new_n505_ = ~new_n175_ & ~new_n335_;
  assign new_n506_ = v26 & v27;
  assign new_n507_ = new_n174_ & new_n506_;
  assign new_n508_ = ~new_n505_ & ~new_n507_;
  assign new_n509_ = v24 & ~new_n338_;
  assign new_n510_ = ~v0 & new_n509_;
  assign new_n511_ = new_n174_ & new_n268_;
  assign new_n512_ = ~new_n510_ & ~new_n511_;
  assign new_n513_ = new_n508_ & new_n512_;
  assign new_n514_ = v25 & ~new_n513_;
  assign new_n515_ = ~new_n504_ & ~new_n514_;
  assign \v32.17  = ~v1 & ~new_n515_;
  assign new_n517_ = v12 & v27;
  assign new_n518_ = v10 & new_n517_;
  assign new_n519_ = ~v8 & new_n518_;
  assign new_n520_ = v2 & new_n519_;
  assign new_n521_ = v0 & new_n520_;
  assign new_n522_ = ~v21 & ~new_n211_;
  assign new_n523_ = ~new_n131_ & ~new_n522_;
  assign new_n524_ = ~new_n398_ & new_n523_;
  assign new_n525_ = v31 & new_n524_;
  assign new_n526_ = ~v27 & new_n525_;
  assign new_n527_ = v20 & new_n526_;
  assign new_n528_ = ~v18 & new_n527_;
  assign new_n529_ = ~v16 & new_n528_;
  assign new_n530_ = ~v7 & new_n529_;
  assign new_n531_ = v3 & new_n530_;
  assign new_n532_ = ~v0 & new_n531_;
  assign new_n533_ = ~new_n521_ & ~new_n532_;
  assign new_n534_ = ~v25 & ~new_n533_;
  assign new_n535_ = ~new_n267_ & ~new_n336_;
  assign new_n536_ = ~new_n175_ & ~new_n535_;
  assign new_n537_ = v27 & v28;
  assign new_n538_ = new_n174_ & new_n537_;
  assign new_n539_ = ~new_n536_ & ~new_n538_;
  assign new_n540_ = v26 & ~new_n539_;
  assign new_n541_ = v25 & new_n540_;
  assign new_n542_ = ~new_n534_ & ~new_n541_;
  assign \v32.18  = ~v1 & ~new_n542_;
  assign new_n544_ = ~v5 & new_n366_;
  assign new_n545_ = v0 & new_n544_;
  assign new_n546_ = v21 & v22;
  assign new_n547_ = ~new_n156_ & ~new_n546_;
  assign new_n548_ = v20 & ~new_n547_;
  assign new_n549_ = ~v20 & new_n546_;
  assign new_n550_ = ~new_n548_ & ~new_n549_;
  assign new_n551_ = ~new_n131_ & ~new_n550_;
  assign new_n552_ = ~new_n398_ & new_n551_;
  assign new_n553_ = v31 & new_n552_;
  assign new_n554_ = ~v18 & new_n553_;
  assign new_n555_ = ~v16 & new_n554_;
  assign new_n556_ = v3 & new_n555_;
  assign new_n557_ = ~v0 & new_n556_;
  assign new_n558_ = ~new_n545_ & ~new_n557_;
  assign new_n559_ = ~v27 & ~new_n558_;
  assign new_n560_ = ~v7 & new_n559_;
  assign new_n561_ = v13 & v27;
  assign new_n562_ = v10 & new_n561_;
  assign new_n563_ = ~v8 & new_n562_;
  assign new_n564_ = v2 & new_n563_;
  assign new_n565_ = v0 & new_n564_;
  assign new_n566_ = ~new_n560_ & ~new_n565_;
  assign new_n567_ = ~v25 & ~new_n566_;
  assign new_n568_ = ~v26 & new_n537_;
  assign new_n569_ = v26 & new_n241_;
  assign new_n570_ = ~new_n568_ & ~new_n569_;
  assign new_n571_ = ~new_n175_ & ~new_n570_;
  assign new_n572_ = v26 & new_n537_;
  assign new_n573_ = new_n174_ & new_n572_;
  assign new_n574_ = ~new_n571_ & ~new_n573_;
  assign new_n575_ = v25 & ~new_n574_;
  assign new_n576_ = ~new_n567_ & ~new_n575_;
  assign \v32.19  = ~v1 & ~new_n576_;
  assign \v32.0  = 1'b0;
endmodule


