// Benchmark "c1908.blif" written by ABC on Fri Feb 25 15:12:56 2022

module c1908  ( 
    G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
    G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237,
    G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_;
  assign new_n59_ = ~G237 & ~G902;
  assign new_n60_ = G214 & ~new_n59_;
  assign new_n61_ = G143 & ~G146;
  assign new_n62_ = ~G143 & G146;
  assign new_n63_ = ~new_n61_ & ~new_n62_;
  assign new_n64_ = G128 & ~new_n63_;
  assign new_n65_ = ~G128 & new_n63_;
  assign new_n66_ = ~new_n64_ & ~new_n65_;
  assign new_n67_ = G125 & ~new_n66_;
  assign new_n68_ = ~G125 & new_n66_;
  assign new_n69_ = ~new_n67_ & ~new_n68_;
  assign new_n70_ = G224 & ~G953;
  assign new_n71_ = ~new_n69_ & ~new_n70_;
  assign new_n72_ = new_n69_ & new_n70_;
  assign new_n73_ = ~new_n71_ & ~new_n72_;
  assign new_n74_ = G104 & ~G107;
  assign new_n75_ = ~G104 & G107;
  assign new_n76_ = ~new_n74_ & ~new_n75_;
  assign new_n77_ = G101 & ~new_n76_;
  assign new_n78_ = ~G101 & new_n76_;
  assign new_n79_ = ~new_n77_ & ~new_n78_;
  assign new_n80_ = G116 & ~G119;
  assign new_n81_ = ~G116 & G119;
  assign new_n82_ = ~new_n80_ & ~new_n81_;
  assign new_n83_ = G113 & ~new_n82_;
  assign new_n84_ = ~G113 & new_n82_;
  assign new_n85_ = ~new_n83_ & ~new_n84_;
  assign new_n86_ = new_n79_ & new_n85_;
  assign new_n87_ = ~new_n79_ & ~new_n85_;
  assign new_n88_ = ~new_n86_ & ~new_n87_;
  assign new_n89_ = G110 & ~G122;
  assign new_n90_ = ~G110 & G122;
  assign new_n91_ = ~new_n89_ & ~new_n90_;
  assign new_n92_ = ~new_n88_ & ~new_n91_;
  assign new_n93_ = new_n88_ & new_n91_;
  assign new_n94_ = ~new_n92_ & ~new_n93_;
  assign new_n95_ = new_n73_ & new_n94_;
  assign new_n96_ = ~new_n73_ & ~new_n94_;
  assign new_n97_ = ~new_n95_ & ~new_n96_;
  assign new_n98_ = ~G902 & new_n97_;
  assign new_n99_ = G210 & ~new_n59_;
  assign new_n100_ = ~new_n98_ & new_n99_;
  assign new_n101_ = new_n98_ & ~new_n99_;
  assign new_n102_ = ~new_n100_ & ~new_n101_;
  assign new_n103_ = ~new_n60_ & ~new_n102_;
  assign new_n104_ = G234 & ~G902;
  assign new_n105_ = G221 & ~new_n104_;
  assign new_n106_ = ~G110 & G140;
  assign new_n107_ = G110 & ~G140;
  assign new_n108_ = ~new_n106_ & ~new_n107_;
  assign new_n109_ = G227 & ~G953;
  assign new_n110_ = ~new_n108_ & ~new_n109_;
  assign new_n111_ = new_n108_ & new_n109_;
  assign new_n112_ = ~new_n110_ & ~new_n111_;
  assign new_n113_ = ~new_n66_ & ~new_n79_;
  assign new_n114_ = new_n66_ & new_n79_;
  assign new_n115_ = ~new_n113_ & ~new_n114_;
  assign new_n116_ = G134 & ~G137;
  assign new_n117_ = ~G134 & G137;
  assign new_n118_ = ~new_n116_ & ~new_n117_;
  assign new_n119_ = G131 & ~new_n118_;
  assign new_n120_ = ~G131 & new_n118_;
  assign new_n121_ = ~new_n119_ & ~new_n120_;
  assign new_n122_ = ~new_n115_ & ~new_n121_;
  assign new_n123_ = new_n115_ & new_n121_;
  assign new_n124_ = ~new_n122_ & ~new_n123_;
  assign new_n125_ = ~new_n112_ & ~new_n124_;
  assign new_n126_ = new_n112_ & new_n124_;
  assign new_n127_ = ~new_n125_ & ~new_n126_;
  assign new_n128_ = ~G902 & ~new_n127_;
  assign new_n129_ = G469 & ~new_n128_;
  assign new_n130_ = ~G469 & new_n128_;
  assign new_n131_ = ~new_n129_ & ~new_n130_;
  assign new_n132_ = ~new_n105_ & ~new_n131_;
  assign new_n133_ = ~G125 & G140;
  assign new_n134_ = G125 & ~G140;
  assign new_n135_ = ~new_n133_ & ~new_n134_;
  assign new_n136_ = G146 & ~new_n135_;
  assign new_n137_ = ~G146 & new_n135_;
  assign new_n138_ = ~new_n136_ & ~new_n137_;
  assign new_n139_ = G119 & ~G128;
  assign new_n140_ = ~G119 & G128;
  assign new_n141_ = ~new_n139_ & ~new_n140_;
  assign new_n142_ = G110 & ~new_n141_;
  assign new_n143_ = ~G110 & new_n141_;
  assign new_n144_ = ~new_n142_ & ~new_n143_;
  assign new_n145_ = new_n138_ & ~new_n144_;
  assign new_n146_ = ~new_n138_ & new_n144_;
  assign new_n147_ = ~new_n145_ & ~new_n146_;
  assign new_n148_ = G221 & G234;
  assign new_n149_ = ~G953 & new_n148_;
  assign new_n150_ = G137 & new_n149_;
  assign new_n151_ = ~G137 & ~new_n149_;
  assign new_n152_ = ~new_n150_ & ~new_n151_;
  assign new_n153_ = ~new_n147_ & ~new_n152_;
  assign new_n154_ = new_n147_ & new_n152_;
  assign new_n155_ = ~new_n153_ & ~new_n154_;
  assign new_n156_ = ~G902 & ~new_n155_;
  assign new_n157_ = G217 & ~new_n104_;
  assign new_n158_ = ~new_n156_ & new_n157_;
  assign new_n159_ = new_n156_ & ~new_n157_;
  assign new_n160_ = ~new_n158_ & ~new_n159_;
  assign new_n161_ = G210 & ~G237;
  assign new_n162_ = ~G953 & new_n161_;
  assign new_n163_ = ~G101 & ~new_n162_;
  assign new_n164_ = G101 & new_n162_;
  assign new_n165_ = ~new_n163_ & ~new_n164_;
  assign new_n166_ = new_n66_ & new_n121_;
  assign new_n167_ = ~new_n66_ & ~new_n121_;
  assign new_n168_ = ~new_n166_ & ~new_n167_;
  assign new_n169_ = ~new_n85_ & ~new_n168_;
  assign new_n170_ = new_n85_ & new_n168_;
  assign new_n171_ = ~new_n169_ & ~new_n170_;
  assign new_n172_ = new_n165_ & ~new_n171_;
  assign new_n173_ = ~new_n165_ & new_n171_;
  assign new_n174_ = ~new_n172_ & ~new_n173_;
  assign new_n175_ = ~G902 & ~new_n174_;
  assign new_n176_ = G472 & ~new_n175_;
  assign new_n177_ = ~G472 & new_n175_;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign new_n179_ = new_n160_ & ~new_n178_;
  assign new_n180_ = G116 & ~G122;
  assign new_n181_ = ~G116 & G122;
  assign new_n182_ = ~new_n180_ & ~new_n181_;
  assign new_n183_ = G107 & ~new_n182_;
  assign new_n184_ = ~G107 & new_n182_;
  assign new_n185_ = ~new_n183_ & ~new_n184_;
  assign new_n186_ = G128 & ~G143;
  assign new_n187_ = ~G128 & G143;
  assign new_n188_ = ~new_n186_ & ~new_n187_;
  assign new_n189_ = G134 & ~new_n188_;
  assign new_n190_ = ~G134 & new_n188_;
  assign new_n191_ = ~new_n189_ & ~new_n190_;
  assign new_n192_ = ~new_n185_ & new_n191_;
  assign new_n193_ = new_n185_ & ~new_n191_;
  assign new_n194_ = ~new_n192_ & ~new_n193_;
  assign new_n195_ = G217 & G234;
  assign new_n196_ = ~G953 & new_n195_;
  assign new_n197_ = ~new_n194_ & ~new_n196_;
  assign new_n198_ = new_n194_ & new_n196_;
  assign new_n199_ = ~new_n197_ & ~new_n198_;
  assign new_n200_ = ~G902 & ~new_n199_;
  assign new_n201_ = G478 & ~new_n200_;
  assign new_n202_ = ~G478 & new_n200_;
  assign new_n203_ = ~new_n201_ & ~new_n202_;
  assign new_n204_ = G214 & ~G237;
  assign new_n205_ = ~G953 & new_n204_;
  assign new_n206_ = ~G143 & ~new_n205_;
  assign new_n207_ = G143 & new_n205_;
  assign new_n208_ = ~new_n206_ & ~new_n207_;
  assign new_n209_ = G131 & ~new_n208_;
  assign new_n210_ = ~G131 & new_n208_;
  assign new_n211_ = ~new_n209_ & ~new_n210_;
  assign new_n212_ = ~new_n138_ & new_n211_;
  assign new_n213_ = new_n138_ & ~new_n211_;
  assign new_n214_ = ~new_n212_ & ~new_n213_;
  assign new_n215_ = G113 & ~G122;
  assign new_n216_ = ~G113 & G122;
  assign new_n217_ = ~new_n215_ & ~new_n216_;
  assign new_n218_ = G104 & ~new_n217_;
  assign new_n219_ = ~G104 & new_n217_;
  assign new_n220_ = ~new_n218_ & ~new_n219_;
  assign new_n221_ = ~new_n214_ & new_n220_;
  assign new_n222_ = new_n214_ & ~new_n220_;
  assign new_n223_ = ~new_n221_ & ~new_n222_;
  assign new_n224_ = ~G902 & ~new_n223_;
  assign new_n225_ = G475 & ~new_n224_;
  assign new_n226_ = ~G475 & new_n224_;
  assign new_n227_ = ~new_n225_ & ~new_n226_;
  assign new_n228_ = new_n203_ & new_n227_;
  assign new_n229_ = G234 & G237;
  assign new_n230_ = ~G898 & G902;
  assign new_n231_ = G953 & ~new_n229_;
  assign new_n232_ = new_n230_ & new_n231_;
  assign new_n233_ = G952 & ~G953;
  assign new_n234_ = ~new_n229_ & new_n233_;
  assign new_n235_ = ~new_n232_ & ~new_n234_;
  assign new_n236_ = new_n103_ & new_n132_;
  assign new_n237_ = new_n179_ & new_n236_;
  assign new_n238_ = new_n228_ & new_n237_;
  assign new_n239_ = ~new_n235_ & new_n238_;
  assign new_n240_ = ~G101 & new_n239_;
  assign new_n241_ = G101 & ~new_n239_;
  assign G3 = new_n240_ | new_n241_;
  assign new_n243_ = new_n160_ & new_n178_;
  assign new_n244_ = new_n203_ & ~new_n227_;
  assign new_n245_ = new_n236_ & new_n243_;
  assign new_n246_ = new_n244_ & new_n245_;
  assign new_n247_ = ~new_n235_ & new_n246_;
  assign new_n248_ = ~G104 & new_n247_;
  assign new_n249_ = G104 & ~new_n247_;
  assign G6 = new_n248_ | new_n249_;
  assign new_n251_ = ~new_n203_ & new_n227_;
  assign new_n252_ = new_n245_ & new_n251_;
  assign new_n253_ = ~new_n235_ & new_n252_;
  assign new_n254_ = ~G107 & new_n253_;
  assign new_n255_ = G107 & ~new_n253_;
  assign G9 = new_n254_ | new_n255_;
  assign new_n257_ = ~new_n160_ & new_n178_;
  assign new_n258_ = new_n236_ & new_n257_;
  assign new_n259_ = new_n228_ & new_n258_;
  assign new_n260_ = ~new_n235_ & new_n259_;
  assign new_n261_ = ~G110 & new_n260_;
  assign new_n262_ = G110 & ~new_n260_;
  assign G12 = new_n261_ | new_n262_;
  assign new_n264_ = ~new_n160_ & ~new_n178_;
  assign new_n265_ = ~G900 & G902;
  assign new_n266_ = new_n231_ & new_n265_;
  assign new_n267_ = ~new_n234_ & ~new_n266_;
  assign new_n268_ = new_n236_ & new_n264_;
  assign new_n269_ = new_n251_ & new_n268_;
  assign new_n270_ = ~new_n267_ & new_n269_;
  assign new_n271_ = ~G128 & new_n270_;
  assign new_n272_ = G128 & ~new_n270_;
  assign G30 = new_n271_ | new_n272_;
  assign new_n274_ = ~new_n203_ & ~new_n227_;
  assign new_n275_ = new_n237_ & new_n274_;
  assign new_n276_ = ~new_n267_ & new_n275_;
  assign new_n277_ = ~G143 & new_n276_;
  assign new_n278_ = G143 & ~new_n276_;
  assign G45 = new_n277_ | new_n278_;
  assign new_n280_ = new_n244_ & new_n268_;
  assign new_n281_ = ~new_n267_ & new_n280_;
  assign new_n282_ = ~G146 & new_n281_;
  assign new_n283_ = G146 & ~new_n281_;
  assign G48 = new_n282_ | new_n283_;
  assign new_n285_ = ~new_n105_ & new_n131_;
  assign new_n286_ = new_n103_ & new_n285_;
  assign new_n287_ = new_n179_ & new_n286_;
  assign new_n288_ = new_n244_ & new_n287_;
  assign new_n289_ = ~new_n235_ & new_n288_;
  assign new_n290_ = ~G113 & new_n289_;
  assign new_n291_ = G113 & ~new_n289_;
  assign G15 = new_n290_ | new_n291_;
  assign new_n293_ = new_n251_ & new_n287_;
  assign new_n294_ = ~new_n235_ & new_n293_;
  assign new_n295_ = ~G116 & new_n294_;
  assign new_n296_ = G116 & ~new_n294_;
  assign G18 = new_n295_ | new_n296_;
  assign new_n298_ = new_n264_ & new_n286_;
  assign new_n299_ = new_n228_ & new_n298_;
  assign new_n300_ = ~new_n235_ & new_n299_;
  assign new_n301_ = ~G119 & new_n300_;
  assign new_n302_ = G119 & ~new_n300_;
  assign G21 = new_n301_ | new_n302_;
  assign new_n304_ = new_n243_ & new_n286_;
  assign new_n305_ = new_n274_ & new_n304_;
  assign new_n306_ = ~new_n235_ & new_n305_;
  assign new_n307_ = ~G122 & new_n306_;
  assign new_n308_ = G122 & ~new_n306_;
  assign G24 = new_n307_ | new_n308_;
  assign new_n310_ = new_n257_ & new_n286_;
  assign new_n311_ = new_n244_ & new_n310_;
  assign new_n312_ = ~new_n267_ & new_n311_;
  assign new_n313_ = ~G125 & new_n312_;
  assign new_n314_ = G125 & ~new_n312_;
  assign G27 = new_n313_ | new_n314_;
  assign new_n316_ = ~new_n60_ & new_n102_;
  assign new_n317_ = new_n132_ & new_n316_;
  assign new_n318_ = new_n179_ & new_n317_;
  assign new_n319_ = new_n244_ & new_n318_;
  assign new_n320_ = ~new_n267_ & new_n319_;
  assign new_n321_ = ~G131 & new_n320_;
  assign new_n322_ = G131 & ~new_n320_;
  assign G33 = new_n321_ | new_n322_;
  assign new_n324_ = new_n251_ & new_n318_;
  assign new_n325_ = ~new_n267_ & new_n324_;
  assign new_n326_ = ~G134 & new_n325_;
  assign new_n327_ = G134 & ~new_n325_;
  assign G36 = new_n326_ | new_n327_;
  assign new_n329_ = new_n264_ & new_n317_;
  assign new_n330_ = new_n228_ & new_n329_;
  assign new_n331_ = ~new_n267_ & new_n330_;
  assign new_n332_ = ~G137 & new_n331_;
  assign new_n333_ = G137 & ~new_n331_;
  assign G39 = new_n332_ | new_n333_;
  assign new_n335_ = new_n257_ & new_n317_;
  assign new_n336_ = new_n244_ & new_n335_;
  assign new_n337_ = ~new_n267_ & new_n336_;
  assign new_n338_ = ~G140 & new_n337_;
  assign new_n339_ = G140 & ~new_n337_;
  assign G42 = new_n338_ | new_n339_;
  assign new_n341_ = new_n160_ & new_n203_;
  assign new_n342_ = new_n178_ & new_n227_;
  assign new_n343_ = new_n341_ & new_n342_;
  assign new_n344_ = new_n102_ & ~new_n105_;
  assign new_n345_ = ~new_n60_ & new_n131_;
  assign new_n346_ = new_n344_ & new_n345_;
  assign new_n347_ = new_n343_ & new_n346_;
  assign new_n348_ = ~G952 & ~G953;
  assign new_n349_ = ~new_n347_ & new_n348_;
  assign new_n350_ = new_n228_ & ~new_n235_;
  assign new_n351_ = new_n237_ & new_n350_;
  assign new_n352_ = ~new_n235_ & new_n244_;
  assign new_n353_ = new_n245_ & new_n352_;
  assign new_n354_ = ~new_n235_ & new_n251_;
  assign new_n355_ = new_n245_ & new_n354_;
  assign new_n356_ = new_n258_ & new_n350_;
  assign new_n357_ = new_n287_ & new_n352_;
  assign new_n358_ = new_n287_ & new_n354_;
  assign new_n359_ = new_n298_ & new_n350_;
  assign new_n360_ = ~new_n235_ & new_n274_;
  assign new_n361_ = new_n304_ & new_n360_;
  assign new_n362_ = ~new_n351_ & ~new_n353_;
  assign new_n363_ = ~new_n355_ & new_n362_;
  assign new_n364_ = ~new_n356_ & new_n363_;
  assign new_n365_ = ~new_n357_ & new_n364_;
  assign new_n366_ = ~new_n358_ & new_n365_;
  assign new_n367_ = ~new_n359_ & new_n366_;
  assign new_n368_ = ~new_n361_ & new_n367_;
  assign new_n369_ = new_n244_ & ~new_n267_;
  assign new_n370_ = new_n310_ & new_n369_;
  assign new_n371_ = new_n251_ & ~new_n267_;
  assign new_n372_ = new_n268_ & new_n371_;
  assign new_n373_ = new_n318_ & new_n369_;
  assign new_n374_ = new_n318_ & new_n371_;
  assign new_n375_ = new_n228_ & ~new_n267_;
  assign new_n376_ = new_n329_ & new_n375_;
  assign new_n377_ = new_n335_ & new_n369_;
  assign new_n378_ = ~new_n267_ & new_n274_;
  assign new_n379_ = new_n237_ & new_n378_;
  assign new_n380_ = new_n268_ & new_n369_;
  assign new_n381_ = ~new_n370_ & ~new_n372_;
  assign new_n382_ = ~new_n373_ & new_n381_;
  assign new_n383_ = ~new_n374_ & new_n382_;
  assign new_n384_ = ~new_n376_ & new_n383_;
  assign new_n385_ = ~new_n377_ & new_n384_;
  assign new_n386_ = ~new_n379_ & new_n385_;
  assign new_n387_ = ~new_n380_ & new_n386_;
  assign new_n388_ = new_n228_ & new_n234_;
  assign new_n389_ = new_n304_ & new_n388_;
  assign new_n390_ = new_n243_ & new_n317_;
  assign new_n391_ = new_n388_ & new_n390_;
  assign new_n392_ = new_n285_ & new_n316_;
  assign new_n393_ = new_n179_ & new_n392_;
  assign new_n394_ = new_n388_ & new_n393_;
  assign new_n395_ = new_n243_ & new_n392_;
  assign new_n396_ = new_n234_ & new_n244_;
  assign new_n397_ = new_n395_ & new_n396_;
  assign new_n398_ = new_n234_ & new_n251_;
  assign new_n399_ = new_n395_ & new_n398_;
  assign new_n400_ = new_n257_ & new_n392_;
  assign new_n401_ = new_n388_ & new_n400_;
  assign new_n402_ = new_n105_ & new_n131_;
  assign new_n403_ = new_n316_ & new_n402_;
  assign new_n404_ = new_n243_ & new_n403_;
  assign new_n405_ = new_n388_ & new_n404_;
  assign new_n406_ = new_n60_ & new_n102_;
  assign new_n407_ = new_n285_ & new_n406_;
  assign new_n408_ = new_n243_ & new_n407_;
  assign new_n409_ = new_n388_ & new_n408_;
  assign new_n410_ = ~new_n389_ & ~new_n391_;
  assign new_n411_ = ~new_n394_ & new_n410_;
  assign new_n412_ = ~new_n397_ & new_n411_;
  assign new_n413_ = ~new_n399_ & new_n412_;
  assign new_n414_ = ~new_n401_ & new_n413_;
  assign new_n415_ = ~new_n405_ & new_n414_;
  assign new_n416_ = ~new_n409_ & new_n415_;
  assign new_n417_ = new_n368_ & new_n387_;
  assign new_n418_ = new_n416_ & new_n417_;
  assign new_n419_ = ~G953 & ~new_n347_;
  assign new_n420_ = G952 & new_n419_;
  assign new_n421_ = new_n418_ & new_n420_;
  assign G75 = ~new_n349_ & ~new_n421_;
  assign new_n423_ = ~new_n73_ & new_n94_;
  assign new_n424_ = new_n73_ & ~new_n94_;
  assign new_n425_ = ~new_n423_ & ~new_n424_;
  assign new_n426_ = G902 & new_n99_;
  assign new_n427_ = ~new_n417_ & new_n426_;
  assign new_n428_ = ~new_n425_ & ~new_n427_;
  assign new_n429_ = new_n425_ & new_n427_;
  assign new_n430_ = ~new_n428_ & ~new_n429_;
  assign new_n431_ = ~G952 & G953;
  assign G51 = ~new_n430_ & ~new_n431_;
  assign new_n433_ = G469 & G902;
  assign new_n434_ = ~new_n417_ & new_n433_;
  assign new_n435_ = ~new_n127_ & ~new_n434_;
  assign new_n436_ = new_n127_ & new_n434_;
  assign new_n437_ = ~new_n435_ & ~new_n436_;
  assign G54 = ~new_n431_ & ~new_n437_;
  assign new_n439_ = G475 & G902;
  assign new_n440_ = ~new_n417_ & new_n439_;
  assign new_n441_ = ~new_n223_ & ~new_n440_;
  assign new_n442_ = new_n223_ & new_n440_;
  assign new_n443_ = ~new_n441_ & ~new_n442_;
  assign G60 = ~new_n431_ & ~new_n443_;
  assign new_n445_ = G478 & G902;
  assign new_n446_ = ~new_n417_ & new_n445_;
  assign new_n447_ = ~new_n199_ & ~new_n446_;
  assign new_n448_ = new_n199_ & new_n446_;
  assign new_n449_ = ~new_n447_ & ~new_n448_;
  assign G63 = ~new_n431_ & ~new_n449_;
  assign new_n451_ = G902 & new_n157_;
  assign new_n452_ = ~new_n417_ & new_n451_;
  assign new_n453_ = ~new_n155_ & ~new_n452_;
  assign new_n454_ = new_n155_ & new_n452_;
  assign new_n455_ = ~new_n453_ & ~new_n454_;
  assign G66 = ~new_n431_ & ~new_n455_;
  assign new_n457_ = ~new_n355_ & ~new_n356_;
  assign new_n458_ = new_n362_ & new_n457_;
  assign new_n459_ = ~new_n359_ & ~new_n361_;
  assign new_n460_ = ~new_n357_ & ~new_n358_;
  assign new_n461_ = new_n459_ & new_n460_;
  assign new_n462_ = new_n458_ & new_n461_;
  assign new_n463_ = ~G953 & ~new_n462_;
  assign new_n464_ = ~G898 & G953;
  assign new_n465_ = new_n94_ & ~new_n464_;
  assign new_n466_ = new_n463_ & ~new_n465_;
  assign new_n467_ = ~new_n463_ & new_n465_;
  assign new_n468_ = ~new_n466_ & ~new_n467_;
  assign new_n469_ = G224 & G898;
  assign new_n470_ = G953 & ~new_n469_;
  assign new_n471_ = ~new_n468_ & ~new_n470_;
  assign new_n472_ = new_n468_ & new_n470_;
  assign G69 = new_n471_ | new_n472_;
  assign new_n474_ = ~new_n373_ & ~new_n374_;
  assign new_n475_ = new_n381_ & new_n474_;
  assign new_n476_ = ~new_n379_ & ~new_n380_;
  assign new_n477_ = ~new_n376_ & ~new_n377_;
  assign new_n478_ = new_n476_ & new_n477_;
  assign new_n479_ = new_n475_ & new_n478_;
  assign new_n480_ = ~G953 & ~new_n479_;
  assign new_n481_ = ~G900 & G953;
  assign new_n482_ = ~new_n135_ & ~new_n168_;
  assign new_n483_ = new_n135_ & new_n168_;
  assign new_n484_ = ~new_n482_ & ~new_n483_;
  assign new_n485_ = ~new_n481_ & new_n484_;
  assign new_n486_ = new_n480_ & ~new_n485_;
  assign new_n487_ = ~new_n480_ & new_n485_;
  assign new_n488_ = ~new_n486_ & ~new_n487_;
  assign new_n489_ = G227 & G900;
  assign new_n490_ = G953 & ~new_n489_;
  assign new_n491_ = ~new_n488_ & ~new_n490_;
  assign new_n492_ = new_n488_ & new_n490_;
  assign G72 = new_n491_ | new_n492_;
  assign new_n494_ = G472 & G902;
  assign new_n495_ = ~new_n417_ & new_n494_;
  assign new_n496_ = ~new_n171_ & ~new_n495_;
  assign new_n497_ = new_n171_ & new_n495_;
  assign new_n498_ = ~new_n496_ & ~new_n497_;
  assign new_n499_ = new_n165_ & ~new_n498_;
  assign new_n500_ = ~new_n165_ & new_n498_;
  assign new_n501_ = ~new_n499_ & ~new_n500_;
  assign G57 = ~new_n431_ & ~new_n501_;
endmodule


