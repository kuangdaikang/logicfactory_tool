// Benchmark "priority" written by ABC on Mon Sep 11 23:42:39 2023

module priority ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] ,
    \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] ;
  output \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F;
  wire new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n914_, new_n915_, new_n916_, new_n917_;
  INV_X1     g000(.I(\A[9] ), .ZN(new_n137_));
  INV_X1     g001(.I(\A[11] ), .ZN(new_n138_));
  INV_X1     g002(.I(\A[17] ), .ZN(new_n139_));
  INV_X1     g003(.I(\A[19] ), .ZN(new_n140_));
  INV_X1     g004(.I(\A[21] ), .ZN(new_n141_));
  INV_X1     g005(.I(\A[23] ), .ZN(new_n142_));
  INV_X1     g006(.I(\A[25] ), .ZN(new_n143_));
  INV_X1     g007(.I(\A[27] ), .ZN(new_n144_));
  INV_X1     g008(.I(\A[29] ), .ZN(new_n145_));
  INV_X1     g009(.I(\A[31] ), .ZN(new_n146_));
  INV_X1     g010(.I(\A[33] ), .ZN(new_n147_));
  INV_X1     g011(.I(\A[35] ), .ZN(new_n148_));
  INV_X1     g012(.I(\A[37] ), .ZN(new_n149_));
  INV_X1     g013(.I(\A[39] ), .ZN(new_n150_));
  INV_X1     g014(.I(\A[41] ), .ZN(new_n151_));
  INV_X1     g015(.I(\A[43] ), .ZN(new_n152_));
  INV_X1     g016(.I(\A[45] ), .ZN(new_n153_));
  INV_X1     g017(.I(\A[47] ), .ZN(new_n154_));
  INV_X1     g018(.I(\A[49] ), .ZN(new_n155_));
  INV_X1     g019(.I(\A[51] ), .ZN(new_n156_));
  INV_X1     g020(.I(\A[53] ), .ZN(new_n157_));
  INV_X1     g021(.I(\A[55] ), .ZN(new_n158_));
  INV_X1     g022(.I(\A[57] ), .ZN(new_n159_));
  INV_X1     g023(.I(\A[59] ), .ZN(new_n160_));
  INV_X1     g024(.I(\A[61] ), .ZN(new_n161_));
  INV_X1     g025(.I(\A[63] ), .ZN(new_n162_));
  INV_X1     g026(.I(\A[65] ), .ZN(new_n163_));
  INV_X1     g027(.I(\A[67] ), .ZN(new_n164_));
  INV_X1     g028(.I(\A[69] ), .ZN(new_n165_));
  INV_X1     g029(.I(\A[71] ), .ZN(new_n166_));
  INV_X1     g030(.I(\A[73] ), .ZN(new_n167_));
  INV_X1     g031(.I(\A[75] ), .ZN(new_n168_));
  INV_X1     g032(.I(\A[77] ), .ZN(new_n169_));
  INV_X1     g033(.I(\A[79] ), .ZN(new_n170_));
  INV_X1     g034(.I(\A[81] ), .ZN(new_n171_));
  INV_X1     g035(.I(\A[83] ), .ZN(new_n172_));
  INV_X1     g036(.I(\A[85] ), .ZN(new_n173_));
  INV_X1     g037(.I(\A[87] ), .ZN(new_n174_));
  INV_X1     g038(.I(\A[89] ), .ZN(new_n175_));
  INV_X1     g039(.I(\A[91] ), .ZN(new_n176_));
  INV_X1     g040(.I(\A[93] ), .ZN(new_n177_));
  INV_X1     g041(.I(\A[95] ), .ZN(new_n178_));
  INV_X1     g042(.I(\A[97] ), .ZN(new_n179_));
  INV_X1     g043(.I(\A[101] ), .ZN(new_n180_));
  INV_X1     g044(.I(\A[105] ), .ZN(new_n181_));
  INV_X1     g045(.I(\A[109] ), .ZN(new_n182_));
  INV_X1     g046(.I(\A[113] ), .ZN(new_n183_));
  INV_X1     g047(.I(\A[117] ), .ZN(new_n184_));
  INV_X1     g048(.I(\A[121] ), .ZN(new_n185_));
  INV_X1     g049(.I(\A[123] ), .ZN(new_n186_));
  INV_X1     g050(.I(\A[126] ), .ZN(new_n187_));
  AOI21_X1   g051(.A1(new_n187_), .A2(\A[125] ), .B(\A[127] ), .ZN(new_n188_));
  NAND2_X1   g052(.A1(new_n188_), .A2(new_n186_), .ZN(new_n189_));
  INV_X1     g053(.I(\A[127] ), .ZN(new_n190_));
  INV_X1     g054(.I(\A[124] ), .ZN(new_n191_));
  NOR2_X1    g055(.A1(new_n191_), .A2(\A[125] ), .ZN(new_n192_));
  OAI21_X1   g056(.A1(new_n192_), .A2(\A[126] ), .B(new_n190_), .ZN(new_n193_));
  OAI21_X1   g057(.A1(new_n186_), .A2(new_n193_), .B(new_n189_), .ZN(new_n194_));
  NAND2_X1   g058(.A1(new_n194_), .A2(new_n185_), .ZN(new_n195_));
  NAND2_X1   g059(.A1(new_n186_), .A2(\A[122] ), .ZN(new_n196_));
  MUX2_X1    g060(.I0(new_n193_), .I1(new_n188_), .S(new_n196_), .Z(new_n197_));
  NAND2_X1   g061(.A1(new_n197_), .A2(\A[121] ), .ZN(new_n198_));
  AOI21_X1   g062(.A1(new_n198_), .A2(new_n195_), .B(\A[119] ), .ZN(new_n199_));
  INV_X1     g063(.I(\A[119] ), .ZN(new_n200_));
  INV_X1     g064(.I(\A[125] ), .ZN(new_n201_));
  OAI21_X1   g065(.A1(new_n201_), .A2(\A[126] ), .B(new_n190_), .ZN(new_n202_));
  NOR2_X1    g066(.A1(new_n202_), .A2(\A[123] ), .ZN(new_n203_));
  NAND2_X1   g067(.A1(new_n201_), .A2(\A[124] ), .ZN(new_n204_));
  AOI21_X1   g068(.A1(new_n204_), .A2(new_n187_), .B(\A[127] ), .ZN(new_n205_));
  AOI21_X1   g069(.A1(\A[123] ), .A2(new_n205_), .B(new_n203_), .ZN(new_n206_));
  NAND2_X1   g070(.A1(new_n185_), .A2(\A[120] ), .ZN(new_n207_));
  MUX2_X1    g071(.I0(new_n197_), .I1(new_n206_), .S(new_n207_), .Z(new_n208_));
  NOR2_X1    g072(.A1(new_n208_), .A2(new_n200_), .ZN(new_n209_));
  OAI21_X1   g073(.A1(new_n209_), .A2(new_n199_), .B(new_n184_), .ZN(new_n210_));
  NAND2_X1   g074(.A1(new_n198_), .A2(new_n195_), .ZN(new_n211_));
  NAND2_X1   g075(.A1(new_n200_), .A2(\A[118] ), .ZN(new_n212_));
  MUX2_X1    g076(.I0(new_n208_), .I1(new_n211_), .S(new_n212_), .Z(new_n213_));
  NAND2_X1   g077(.A1(new_n213_), .A2(\A[117] ), .ZN(new_n214_));
  AOI21_X1   g078(.A1(new_n214_), .A2(new_n210_), .B(\A[115] ), .ZN(new_n215_));
  INV_X1     g079(.I(\A[115] ), .ZN(new_n216_));
  MUX2_X1    g080(.I0(new_n205_), .I1(new_n202_), .S(new_n196_), .Z(new_n217_));
  MUX2_X1    g081(.I0(new_n217_), .I1(new_n194_), .S(new_n207_), .Z(new_n218_));
  AOI21_X1   g082(.A1(\A[119] ), .A2(new_n218_), .B(new_n199_), .ZN(new_n219_));
  NAND2_X1   g083(.A1(new_n184_), .A2(\A[116] ), .ZN(new_n220_));
  MUX2_X1    g084(.I0(new_n213_), .I1(new_n219_), .S(new_n220_), .Z(new_n221_));
  NOR2_X1    g085(.A1(new_n221_), .A2(new_n216_), .ZN(new_n222_));
  OAI21_X1   g086(.A1(new_n222_), .A2(new_n215_), .B(new_n183_), .ZN(new_n223_));
  NAND2_X1   g087(.A1(new_n214_), .A2(new_n210_), .ZN(new_n224_));
  NAND2_X1   g088(.A1(new_n216_), .A2(\A[114] ), .ZN(new_n225_));
  MUX2_X1    g089(.I0(new_n221_), .I1(new_n224_), .S(new_n225_), .Z(new_n226_));
  NAND2_X1   g090(.A1(new_n226_), .A2(\A[113] ), .ZN(new_n227_));
  AOI21_X1   g091(.A1(new_n227_), .A2(new_n223_), .B(\A[111] ), .ZN(new_n228_));
  INV_X1     g092(.I(\A[111] ), .ZN(new_n229_));
  MUX2_X1    g093(.I0(new_n218_), .I1(new_n211_), .S(new_n200_), .Z(new_n230_));
  MUX2_X1    g094(.I0(new_n217_), .I1(new_n206_), .S(new_n185_), .Z(new_n231_));
  MUX2_X1    g095(.I0(new_n218_), .I1(new_n231_), .S(new_n212_), .Z(new_n232_));
  MUX2_X1    g096(.I0(new_n232_), .I1(new_n230_), .S(new_n220_), .Z(new_n233_));
  AOI21_X1   g097(.A1(\A[115] ), .A2(new_n233_), .B(new_n215_), .ZN(new_n234_));
  NAND2_X1   g098(.A1(new_n183_), .A2(\A[112] ), .ZN(new_n235_));
  MUX2_X1    g099(.I0(new_n226_), .I1(new_n234_), .S(new_n235_), .Z(new_n236_));
  NOR2_X1    g100(.A1(new_n236_), .A2(new_n229_), .ZN(new_n237_));
  OAI21_X1   g101(.A1(new_n237_), .A2(new_n228_), .B(new_n182_), .ZN(new_n238_));
  NAND2_X1   g102(.A1(new_n227_), .A2(new_n223_), .ZN(new_n239_));
  NAND2_X1   g103(.A1(new_n229_), .A2(\A[110] ), .ZN(new_n240_));
  MUX2_X1    g104(.I0(new_n236_), .I1(new_n239_), .S(new_n240_), .Z(new_n241_));
  NAND2_X1   g105(.A1(new_n241_), .A2(\A[109] ), .ZN(new_n242_));
  AOI21_X1   g106(.A1(new_n242_), .A2(new_n238_), .B(\A[107] ), .ZN(new_n243_));
  INV_X1     g107(.I(\A[107] ), .ZN(new_n244_));
  MUX2_X1    g108(.I0(new_n233_), .I1(new_n224_), .S(new_n216_), .Z(new_n245_));
  MUX2_X1    g109(.I0(new_n232_), .I1(new_n219_), .S(new_n184_), .Z(new_n246_));
  MUX2_X1    g110(.I0(new_n233_), .I1(new_n246_), .S(new_n225_), .Z(new_n247_));
  MUX2_X1    g111(.I0(new_n247_), .I1(new_n245_), .S(new_n235_), .Z(new_n248_));
  AOI21_X1   g112(.A1(\A[111] ), .A2(new_n248_), .B(new_n228_), .ZN(new_n249_));
  NAND2_X1   g113(.A1(new_n182_), .A2(\A[108] ), .ZN(new_n250_));
  MUX2_X1    g114(.I0(new_n241_), .I1(new_n249_), .S(new_n250_), .Z(new_n251_));
  NOR2_X1    g115(.A1(new_n251_), .A2(new_n244_), .ZN(new_n252_));
  OAI21_X1   g116(.A1(new_n252_), .A2(new_n243_), .B(new_n181_), .ZN(new_n253_));
  NAND2_X1   g117(.A1(new_n242_), .A2(new_n238_), .ZN(new_n254_));
  NAND2_X1   g118(.A1(new_n244_), .A2(\A[106] ), .ZN(new_n255_));
  MUX2_X1    g119(.I0(new_n251_), .I1(new_n254_), .S(new_n255_), .Z(new_n256_));
  NAND2_X1   g120(.A1(new_n256_), .A2(\A[105] ), .ZN(new_n257_));
  AOI21_X1   g121(.A1(new_n257_), .A2(new_n253_), .B(\A[103] ), .ZN(new_n258_));
  INV_X1     g122(.I(\A[103] ), .ZN(new_n259_));
  MUX2_X1    g123(.I0(new_n248_), .I1(new_n239_), .S(new_n229_), .Z(new_n260_));
  MUX2_X1    g124(.I0(new_n247_), .I1(new_n234_), .S(new_n183_), .Z(new_n261_));
  MUX2_X1    g125(.I0(new_n248_), .I1(new_n261_), .S(new_n240_), .Z(new_n262_));
  MUX2_X1    g126(.I0(new_n262_), .I1(new_n260_), .S(new_n250_), .Z(new_n263_));
  AOI21_X1   g127(.A1(\A[107] ), .A2(new_n263_), .B(new_n243_), .ZN(new_n264_));
  NAND2_X1   g128(.A1(new_n181_), .A2(\A[104] ), .ZN(new_n265_));
  MUX2_X1    g129(.I0(new_n256_), .I1(new_n264_), .S(new_n265_), .Z(new_n266_));
  NOR2_X1    g130(.A1(new_n266_), .A2(new_n259_), .ZN(new_n267_));
  OAI21_X1   g131(.A1(new_n267_), .A2(new_n258_), .B(new_n180_), .ZN(new_n268_));
  NAND2_X1   g132(.A1(new_n257_), .A2(new_n253_), .ZN(new_n269_));
  NAND2_X1   g133(.A1(new_n259_), .A2(\A[102] ), .ZN(new_n270_));
  MUX2_X1    g134(.I0(new_n266_), .I1(new_n269_), .S(new_n270_), .Z(new_n271_));
  NAND2_X1   g135(.A1(new_n271_), .A2(\A[101] ), .ZN(new_n272_));
  AOI21_X1   g136(.A1(new_n272_), .A2(new_n268_), .B(\A[99] ), .ZN(new_n273_));
  INV_X1     g137(.I(\A[99] ), .ZN(new_n274_));
  MUX2_X1    g138(.I0(new_n263_), .I1(new_n254_), .S(new_n244_), .Z(new_n275_));
  MUX2_X1    g139(.I0(new_n262_), .I1(new_n249_), .S(new_n182_), .Z(new_n276_));
  MUX2_X1    g140(.I0(new_n263_), .I1(new_n276_), .S(new_n255_), .Z(new_n277_));
  MUX2_X1    g141(.I0(new_n277_), .I1(new_n275_), .S(new_n265_), .Z(new_n278_));
  AOI21_X1   g142(.A1(\A[103] ), .A2(new_n278_), .B(new_n258_), .ZN(new_n279_));
  NAND2_X1   g143(.A1(new_n180_), .A2(\A[100] ), .ZN(new_n280_));
  MUX2_X1    g144(.I0(new_n271_), .I1(new_n279_), .S(new_n280_), .Z(new_n281_));
  NOR2_X1    g145(.A1(new_n281_), .A2(new_n274_), .ZN(new_n282_));
  OAI21_X1   g146(.A1(new_n282_), .A2(new_n273_), .B(new_n179_), .ZN(new_n283_));
  NAND2_X1   g147(.A1(new_n272_), .A2(new_n268_), .ZN(new_n284_));
  NAND2_X1   g148(.A1(new_n274_), .A2(\A[98] ), .ZN(new_n285_));
  MUX2_X1    g149(.I0(new_n281_), .I1(new_n284_), .S(new_n285_), .Z(new_n286_));
  NAND2_X1   g150(.A1(new_n286_), .A2(\A[97] ), .ZN(new_n287_));
  NAND2_X1   g151(.A1(new_n287_), .A2(new_n283_), .ZN(new_n288_));
  MUX2_X1    g152(.I0(new_n278_), .I1(new_n269_), .S(new_n259_), .Z(new_n289_));
  MUX2_X1    g153(.I0(new_n277_), .I1(new_n264_), .S(new_n181_), .Z(new_n290_));
  MUX2_X1    g154(.I0(new_n278_), .I1(new_n290_), .S(new_n270_), .Z(new_n291_));
  MUX2_X1    g155(.I0(new_n291_), .I1(new_n289_), .S(new_n280_), .Z(new_n292_));
  MUX2_X1    g156(.I0(new_n292_), .I1(new_n284_), .S(new_n274_), .Z(new_n293_));
  MUX2_X1    g157(.I0(new_n291_), .I1(new_n279_), .S(new_n180_), .Z(new_n294_));
  MUX2_X1    g158(.I0(new_n292_), .I1(new_n294_), .S(new_n285_), .Z(new_n295_));
  NAND2_X1   g159(.A1(new_n179_), .A2(\A[96] ), .ZN(new_n296_));
  MUX2_X1    g160(.I0(new_n295_), .I1(new_n293_), .S(new_n296_), .Z(new_n297_));
  MUX2_X1    g161(.I0(new_n297_), .I1(new_n288_), .S(new_n178_), .Z(new_n298_));
  AOI21_X1   g162(.A1(\A[99] ), .A2(new_n292_), .B(new_n273_), .ZN(new_n299_));
  MUX2_X1    g163(.I0(new_n286_), .I1(new_n299_), .S(new_n296_), .Z(new_n300_));
  NAND2_X1   g164(.A1(new_n178_), .A2(\A[94] ), .ZN(new_n301_));
  MUX2_X1    g165(.I0(new_n300_), .I1(new_n288_), .S(new_n301_), .Z(new_n302_));
  MUX2_X1    g166(.I0(new_n302_), .I1(new_n298_), .S(new_n177_), .Z(new_n303_));
  MUX2_X1    g167(.I0(new_n295_), .I1(new_n299_), .S(new_n179_), .Z(new_n304_));
  MUX2_X1    g168(.I0(new_n297_), .I1(new_n304_), .S(new_n301_), .Z(new_n305_));
  NAND2_X1   g169(.A1(new_n177_), .A2(\A[92] ), .ZN(new_n306_));
  MUX2_X1    g170(.I0(new_n305_), .I1(new_n298_), .S(new_n306_), .Z(new_n307_));
  MUX2_X1    g171(.I0(new_n307_), .I1(new_n303_), .S(new_n176_), .Z(new_n308_));
  AOI21_X1   g172(.A1(new_n287_), .A2(new_n283_), .B(\A[95] ), .ZN(new_n309_));
  AOI21_X1   g173(.A1(\A[95] ), .A2(new_n297_), .B(new_n309_), .ZN(new_n310_));
  MUX2_X1    g174(.I0(new_n302_), .I1(new_n310_), .S(new_n306_), .Z(new_n311_));
  NAND2_X1   g175(.A1(new_n176_), .A2(\A[90] ), .ZN(new_n312_));
  MUX2_X1    g176(.I0(new_n311_), .I1(new_n303_), .S(new_n312_), .Z(new_n313_));
  MUX2_X1    g177(.I0(new_n313_), .I1(new_n308_), .S(new_n175_), .Z(new_n314_));
  NOR2_X1    g178(.A1(new_n310_), .A2(\A[93] ), .ZN(new_n315_));
  NOR2_X1    g179(.A1(new_n305_), .A2(new_n177_), .ZN(new_n316_));
  NOR2_X1    g180(.A1(new_n316_), .A2(new_n315_), .ZN(new_n317_));
  MUX2_X1    g181(.I0(new_n307_), .I1(new_n317_), .S(new_n312_), .Z(new_n318_));
  NAND2_X1   g182(.A1(new_n175_), .A2(\A[88] ), .ZN(new_n319_));
  MUX2_X1    g183(.I0(new_n318_), .I1(new_n308_), .S(new_n319_), .Z(new_n320_));
  MUX2_X1    g184(.I0(new_n320_), .I1(new_n314_), .S(new_n174_), .Z(new_n321_));
  MUX2_X1    g185(.I0(new_n311_), .I1(new_n317_), .S(new_n176_), .Z(new_n322_));
  MUX2_X1    g186(.I0(new_n313_), .I1(new_n322_), .S(new_n319_), .Z(new_n323_));
  NAND2_X1   g187(.A1(new_n174_), .A2(\A[86] ), .ZN(new_n324_));
  MUX2_X1    g188(.I0(new_n323_), .I1(new_n314_), .S(new_n324_), .Z(new_n325_));
  MUX2_X1    g189(.I0(new_n325_), .I1(new_n321_), .S(new_n173_), .Z(new_n326_));
  MUX2_X1    g190(.I0(new_n318_), .I1(new_n322_), .S(new_n175_), .Z(new_n327_));
  MUX2_X1    g191(.I0(new_n320_), .I1(new_n327_), .S(new_n324_), .Z(new_n328_));
  NAND2_X1   g192(.A1(new_n173_), .A2(\A[84] ), .ZN(new_n329_));
  MUX2_X1    g193(.I0(new_n328_), .I1(new_n321_), .S(new_n329_), .Z(new_n330_));
  MUX2_X1    g194(.I0(new_n330_), .I1(new_n326_), .S(new_n172_), .Z(new_n331_));
  MUX2_X1    g195(.I0(new_n323_), .I1(new_n327_), .S(new_n174_), .Z(new_n332_));
  MUX2_X1    g196(.I0(new_n325_), .I1(new_n332_), .S(new_n329_), .Z(new_n333_));
  NAND2_X1   g197(.A1(new_n172_), .A2(\A[82] ), .ZN(new_n334_));
  MUX2_X1    g198(.I0(new_n333_), .I1(new_n326_), .S(new_n334_), .Z(new_n335_));
  MUX2_X1    g199(.I0(new_n335_), .I1(new_n331_), .S(new_n171_), .Z(new_n336_));
  MUX2_X1    g200(.I0(new_n328_), .I1(new_n332_), .S(new_n173_), .Z(new_n337_));
  MUX2_X1    g201(.I0(new_n330_), .I1(new_n337_), .S(new_n334_), .Z(new_n338_));
  NAND2_X1   g202(.A1(new_n171_), .A2(\A[80] ), .ZN(new_n339_));
  MUX2_X1    g203(.I0(new_n338_), .I1(new_n331_), .S(new_n339_), .Z(new_n340_));
  MUX2_X1    g204(.I0(new_n340_), .I1(new_n336_), .S(new_n170_), .Z(new_n341_));
  MUX2_X1    g205(.I0(new_n333_), .I1(new_n337_), .S(new_n172_), .Z(new_n342_));
  MUX2_X1    g206(.I0(new_n335_), .I1(new_n342_), .S(new_n339_), .Z(new_n343_));
  NAND2_X1   g207(.A1(new_n170_), .A2(\A[78] ), .ZN(new_n344_));
  MUX2_X1    g208(.I0(new_n343_), .I1(new_n336_), .S(new_n344_), .Z(new_n345_));
  MUX2_X1    g209(.I0(new_n345_), .I1(new_n341_), .S(new_n169_), .Z(new_n346_));
  MUX2_X1    g210(.I0(new_n338_), .I1(new_n342_), .S(new_n171_), .Z(new_n347_));
  MUX2_X1    g211(.I0(new_n340_), .I1(new_n347_), .S(new_n344_), .Z(new_n348_));
  NAND2_X1   g212(.A1(new_n169_), .A2(\A[76] ), .ZN(new_n349_));
  MUX2_X1    g213(.I0(new_n348_), .I1(new_n341_), .S(new_n349_), .Z(new_n350_));
  MUX2_X1    g214(.I0(new_n350_), .I1(new_n346_), .S(new_n168_), .Z(new_n351_));
  MUX2_X1    g215(.I0(new_n343_), .I1(new_n347_), .S(new_n170_), .Z(new_n352_));
  MUX2_X1    g216(.I0(new_n345_), .I1(new_n352_), .S(new_n349_), .Z(new_n353_));
  NAND2_X1   g217(.A1(new_n168_), .A2(\A[74] ), .ZN(new_n354_));
  MUX2_X1    g218(.I0(new_n353_), .I1(new_n346_), .S(new_n354_), .Z(new_n355_));
  MUX2_X1    g219(.I0(new_n355_), .I1(new_n351_), .S(new_n167_), .Z(new_n356_));
  MUX2_X1    g220(.I0(new_n348_), .I1(new_n352_), .S(new_n169_), .Z(new_n357_));
  MUX2_X1    g221(.I0(new_n350_), .I1(new_n357_), .S(new_n354_), .Z(new_n358_));
  NAND2_X1   g222(.A1(new_n167_), .A2(\A[72] ), .ZN(new_n359_));
  MUX2_X1    g223(.I0(new_n358_), .I1(new_n351_), .S(new_n359_), .Z(new_n360_));
  MUX2_X1    g224(.I0(new_n360_), .I1(new_n356_), .S(new_n166_), .Z(new_n361_));
  MUX2_X1    g225(.I0(new_n353_), .I1(new_n357_), .S(new_n168_), .Z(new_n362_));
  MUX2_X1    g226(.I0(new_n355_), .I1(new_n362_), .S(new_n359_), .Z(new_n363_));
  NAND2_X1   g227(.A1(new_n166_), .A2(\A[70] ), .ZN(new_n364_));
  MUX2_X1    g228(.I0(new_n363_), .I1(new_n356_), .S(new_n364_), .Z(new_n365_));
  MUX2_X1    g229(.I0(new_n365_), .I1(new_n361_), .S(new_n165_), .Z(new_n366_));
  MUX2_X1    g230(.I0(new_n358_), .I1(new_n362_), .S(new_n167_), .Z(new_n367_));
  MUX2_X1    g231(.I0(new_n360_), .I1(new_n367_), .S(new_n364_), .Z(new_n368_));
  NAND2_X1   g232(.A1(new_n165_), .A2(\A[68] ), .ZN(new_n369_));
  MUX2_X1    g233(.I0(new_n368_), .I1(new_n361_), .S(new_n369_), .Z(new_n370_));
  MUX2_X1    g234(.I0(new_n370_), .I1(new_n366_), .S(new_n164_), .Z(new_n371_));
  MUX2_X1    g235(.I0(new_n363_), .I1(new_n367_), .S(new_n166_), .Z(new_n372_));
  MUX2_X1    g236(.I0(new_n365_), .I1(new_n372_), .S(new_n369_), .Z(new_n373_));
  NAND2_X1   g237(.A1(new_n164_), .A2(\A[66] ), .ZN(new_n374_));
  MUX2_X1    g238(.I0(new_n373_), .I1(new_n366_), .S(new_n374_), .Z(new_n375_));
  MUX2_X1    g239(.I0(new_n375_), .I1(new_n371_), .S(new_n163_), .Z(new_n376_));
  MUX2_X1    g240(.I0(new_n368_), .I1(new_n372_), .S(new_n165_), .Z(new_n377_));
  MUX2_X1    g241(.I0(new_n370_), .I1(new_n377_), .S(new_n374_), .Z(new_n378_));
  NAND2_X1   g242(.A1(new_n163_), .A2(\A[64] ), .ZN(new_n379_));
  MUX2_X1    g243(.I0(new_n378_), .I1(new_n371_), .S(new_n379_), .Z(new_n380_));
  MUX2_X1    g244(.I0(new_n380_), .I1(new_n376_), .S(new_n162_), .Z(new_n381_));
  MUX2_X1    g245(.I0(new_n373_), .I1(new_n377_), .S(new_n164_), .Z(new_n382_));
  MUX2_X1    g246(.I0(new_n375_), .I1(new_n382_), .S(new_n379_), .Z(new_n383_));
  NAND2_X1   g247(.A1(new_n162_), .A2(\A[62] ), .ZN(new_n384_));
  MUX2_X1    g248(.I0(new_n383_), .I1(new_n376_), .S(new_n384_), .Z(new_n385_));
  MUX2_X1    g249(.I0(new_n385_), .I1(new_n381_), .S(new_n161_), .Z(new_n386_));
  MUX2_X1    g250(.I0(new_n378_), .I1(new_n382_), .S(new_n163_), .Z(new_n387_));
  MUX2_X1    g251(.I0(new_n380_), .I1(new_n387_), .S(new_n384_), .Z(new_n388_));
  NAND2_X1   g252(.A1(new_n161_), .A2(\A[60] ), .ZN(new_n389_));
  MUX2_X1    g253(.I0(new_n388_), .I1(new_n381_), .S(new_n389_), .Z(new_n390_));
  MUX2_X1    g254(.I0(new_n390_), .I1(new_n386_), .S(new_n160_), .Z(new_n391_));
  MUX2_X1    g255(.I0(new_n383_), .I1(new_n387_), .S(new_n162_), .Z(new_n392_));
  MUX2_X1    g256(.I0(new_n385_), .I1(new_n392_), .S(new_n389_), .Z(new_n393_));
  NAND2_X1   g257(.A1(new_n160_), .A2(\A[58] ), .ZN(new_n394_));
  MUX2_X1    g258(.I0(new_n393_), .I1(new_n386_), .S(new_n394_), .Z(new_n395_));
  MUX2_X1    g259(.I0(new_n395_), .I1(new_n391_), .S(new_n159_), .Z(new_n396_));
  MUX2_X1    g260(.I0(new_n388_), .I1(new_n392_), .S(new_n161_), .Z(new_n397_));
  MUX2_X1    g261(.I0(new_n390_), .I1(new_n397_), .S(new_n394_), .Z(new_n398_));
  NAND2_X1   g262(.A1(new_n159_), .A2(\A[56] ), .ZN(new_n399_));
  MUX2_X1    g263(.I0(new_n398_), .I1(new_n391_), .S(new_n399_), .Z(new_n400_));
  MUX2_X1    g264(.I0(new_n400_), .I1(new_n396_), .S(new_n158_), .Z(new_n401_));
  MUX2_X1    g265(.I0(new_n393_), .I1(new_n397_), .S(new_n160_), .Z(new_n402_));
  MUX2_X1    g266(.I0(new_n395_), .I1(new_n402_), .S(new_n399_), .Z(new_n403_));
  NAND2_X1   g267(.A1(new_n158_), .A2(\A[54] ), .ZN(new_n404_));
  MUX2_X1    g268(.I0(new_n403_), .I1(new_n396_), .S(new_n404_), .Z(new_n405_));
  MUX2_X1    g269(.I0(new_n405_), .I1(new_n401_), .S(new_n157_), .Z(new_n406_));
  MUX2_X1    g270(.I0(new_n398_), .I1(new_n402_), .S(new_n159_), .Z(new_n407_));
  MUX2_X1    g271(.I0(new_n400_), .I1(new_n407_), .S(new_n404_), .Z(new_n408_));
  NAND2_X1   g272(.A1(new_n157_), .A2(\A[52] ), .ZN(new_n409_));
  MUX2_X1    g273(.I0(new_n408_), .I1(new_n401_), .S(new_n409_), .Z(new_n410_));
  MUX2_X1    g274(.I0(new_n410_), .I1(new_n406_), .S(new_n156_), .Z(new_n411_));
  MUX2_X1    g275(.I0(new_n403_), .I1(new_n407_), .S(new_n158_), .Z(new_n412_));
  MUX2_X1    g276(.I0(new_n405_), .I1(new_n412_), .S(new_n409_), .Z(new_n413_));
  NAND2_X1   g277(.A1(new_n156_), .A2(\A[50] ), .ZN(new_n414_));
  MUX2_X1    g278(.I0(new_n413_), .I1(new_n406_), .S(new_n414_), .Z(new_n415_));
  MUX2_X1    g279(.I0(new_n415_), .I1(new_n411_), .S(new_n155_), .Z(new_n416_));
  MUX2_X1    g280(.I0(new_n408_), .I1(new_n412_), .S(new_n157_), .Z(new_n417_));
  MUX2_X1    g281(.I0(new_n410_), .I1(new_n417_), .S(new_n414_), .Z(new_n418_));
  NAND2_X1   g282(.A1(new_n155_), .A2(\A[48] ), .ZN(new_n419_));
  MUX2_X1    g283(.I0(new_n418_), .I1(new_n411_), .S(new_n419_), .Z(new_n420_));
  MUX2_X1    g284(.I0(new_n420_), .I1(new_n416_), .S(new_n154_), .Z(new_n421_));
  MUX2_X1    g285(.I0(new_n413_), .I1(new_n417_), .S(new_n156_), .Z(new_n422_));
  MUX2_X1    g286(.I0(new_n415_), .I1(new_n422_), .S(new_n419_), .Z(new_n423_));
  NAND2_X1   g287(.A1(new_n154_), .A2(\A[46] ), .ZN(new_n424_));
  MUX2_X1    g288(.I0(new_n423_), .I1(new_n416_), .S(new_n424_), .Z(new_n425_));
  MUX2_X1    g289(.I0(new_n425_), .I1(new_n421_), .S(new_n153_), .Z(new_n426_));
  MUX2_X1    g290(.I0(new_n418_), .I1(new_n422_), .S(new_n155_), .Z(new_n427_));
  MUX2_X1    g291(.I0(new_n420_), .I1(new_n427_), .S(new_n424_), .Z(new_n428_));
  NAND2_X1   g292(.A1(new_n153_), .A2(\A[44] ), .ZN(new_n429_));
  MUX2_X1    g293(.I0(new_n428_), .I1(new_n421_), .S(new_n429_), .Z(new_n430_));
  MUX2_X1    g294(.I0(new_n430_), .I1(new_n426_), .S(new_n152_), .Z(new_n431_));
  MUX2_X1    g295(.I0(new_n423_), .I1(new_n427_), .S(new_n154_), .Z(new_n432_));
  MUX2_X1    g296(.I0(new_n425_), .I1(new_n432_), .S(new_n429_), .Z(new_n433_));
  NAND2_X1   g297(.A1(new_n152_), .A2(\A[42] ), .ZN(new_n434_));
  MUX2_X1    g298(.I0(new_n433_), .I1(new_n426_), .S(new_n434_), .Z(new_n435_));
  MUX2_X1    g299(.I0(new_n435_), .I1(new_n431_), .S(new_n151_), .Z(new_n436_));
  MUX2_X1    g300(.I0(new_n428_), .I1(new_n432_), .S(new_n153_), .Z(new_n437_));
  MUX2_X1    g301(.I0(new_n430_), .I1(new_n437_), .S(new_n434_), .Z(new_n438_));
  NAND2_X1   g302(.A1(new_n151_), .A2(\A[40] ), .ZN(new_n439_));
  MUX2_X1    g303(.I0(new_n438_), .I1(new_n431_), .S(new_n439_), .Z(new_n440_));
  MUX2_X1    g304(.I0(new_n440_), .I1(new_n436_), .S(new_n150_), .Z(new_n441_));
  MUX2_X1    g305(.I0(new_n433_), .I1(new_n437_), .S(new_n152_), .Z(new_n442_));
  MUX2_X1    g306(.I0(new_n435_), .I1(new_n442_), .S(new_n439_), .Z(new_n443_));
  NAND2_X1   g307(.A1(new_n150_), .A2(\A[38] ), .ZN(new_n444_));
  MUX2_X1    g308(.I0(new_n443_), .I1(new_n436_), .S(new_n444_), .Z(new_n445_));
  MUX2_X1    g309(.I0(new_n445_), .I1(new_n441_), .S(new_n149_), .Z(new_n446_));
  MUX2_X1    g310(.I0(new_n438_), .I1(new_n442_), .S(new_n151_), .Z(new_n447_));
  MUX2_X1    g311(.I0(new_n440_), .I1(new_n447_), .S(new_n444_), .Z(new_n448_));
  NAND2_X1   g312(.A1(new_n149_), .A2(\A[36] ), .ZN(new_n449_));
  MUX2_X1    g313(.I0(new_n448_), .I1(new_n441_), .S(new_n449_), .Z(new_n450_));
  MUX2_X1    g314(.I0(new_n450_), .I1(new_n446_), .S(new_n148_), .Z(new_n451_));
  MUX2_X1    g315(.I0(new_n443_), .I1(new_n447_), .S(new_n150_), .Z(new_n452_));
  MUX2_X1    g316(.I0(new_n445_), .I1(new_n452_), .S(new_n449_), .Z(new_n453_));
  NAND2_X1   g317(.A1(new_n148_), .A2(\A[34] ), .ZN(new_n454_));
  MUX2_X1    g318(.I0(new_n453_), .I1(new_n446_), .S(new_n454_), .Z(new_n455_));
  MUX2_X1    g319(.I0(new_n455_), .I1(new_n451_), .S(new_n147_), .Z(new_n456_));
  MUX2_X1    g320(.I0(new_n448_), .I1(new_n452_), .S(new_n149_), .Z(new_n457_));
  MUX2_X1    g321(.I0(new_n450_), .I1(new_n457_), .S(new_n454_), .Z(new_n458_));
  NAND2_X1   g322(.A1(new_n147_), .A2(\A[32] ), .ZN(new_n459_));
  MUX2_X1    g323(.I0(new_n458_), .I1(new_n451_), .S(new_n459_), .Z(new_n460_));
  MUX2_X1    g324(.I0(new_n460_), .I1(new_n456_), .S(new_n146_), .Z(new_n461_));
  MUX2_X1    g325(.I0(new_n453_), .I1(new_n457_), .S(new_n148_), .Z(new_n462_));
  MUX2_X1    g326(.I0(new_n455_), .I1(new_n462_), .S(new_n459_), .Z(new_n463_));
  NAND2_X1   g327(.A1(new_n146_), .A2(\A[30] ), .ZN(new_n464_));
  MUX2_X1    g328(.I0(new_n463_), .I1(new_n456_), .S(new_n464_), .Z(new_n465_));
  MUX2_X1    g329(.I0(new_n465_), .I1(new_n461_), .S(new_n145_), .Z(new_n466_));
  MUX2_X1    g330(.I0(new_n458_), .I1(new_n462_), .S(new_n147_), .Z(new_n467_));
  MUX2_X1    g331(.I0(new_n460_), .I1(new_n467_), .S(new_n464_), .Z(new_n468_));
  NAND2_X1   g332(.A1(new_n145_), .A2(\A[28] ), .ZN(new_n469_));
  MUX2_X1    g333(.I0(new_n468_), .I1(new_n461_), .S(new_n469_), .Z(new_n470_));
  MUX2_X1    g334(.I0(new_n470_), .I1(new_n466_), .S(new_n144_), .Z(new_n471_));
  MUX2_X1    g335(.I0(new_n463_), .I1(new_n467_), .S(new_n146_), .Z(new_n472_));
  MUX2_X1    g336(.I0(new_n465_), .I1(new_n472_), .S(new_n469_), .Z(new_n473_));
  NAND2_X1   g337(.A1(new_n144_), .A2(\A[26] ), .ZN(new_n474_));
  MUX2_X1    g338(.I0(new_n473_), .I1(new_n466_), .S(new_n474_), .Z(new_n475_));
  MUX2_X1    g339(.I0(new_n475_), .I1(new_n471_), .S(new_n143_), .Z(new_n476_));
  MUX2_X1    g340(.I0(new_n468_), .I1(new_n472_), .S(new_n145_), .Z(new_n477_));
  MUX2_X1    g341(.I0(new_n470_), .I1(new_n477_), .S(new_n474_), .Z(new_n478_));
  NAND2_X1   g342(.A1(new_n143_), .A2(\A[24] ), .ZN(new_n479_));
  MUX2_X1    g343(.I0(new_n478_), .I1(new_n471_), .S(new_n479_), .Z(new_n480_));
  MUX2_X1    g344(.I0(new_n480_), .I1(new_n476_), .S(new_n142_), .Z(new_n481_));
  MUX2_X1    g345(.I0(new_n473_), .I1(new_n477_), .S(new_n144_), .Z(new_n482_));
  MUX2_X1    g346(.I0(new_n475_), .I1(new_n482_), .S(new_n479_), .Z(new_n483_));
  NAND2_X1   g347(.A1(new_n142_), .A2(\A[22] ), .ZN(new_n484_));
  MUX2_X1    g348(.I0(new_n483_), .I1(new_n476_), .S(new_n484_), .Z(new_n485_));
  MUX2_X1    g349(.I0(new_n485_), .I1(new_n481_), .S(new_n141_), .Z(new_n486_));
  MUX2_X1    g350(.I0(new_n478_), .I1(new_n482_), .S(new_n143_), .Z(new_n487_));
  MUX2_X1    g351(.I0(new_n480_), .I1(new_n487_), .S(new_n484_), .Z(new_n488_));
  NAND2_X1   g352(.A1(new_n141_), .A2(\A[20] ), .ZN(new_n489_));
  MUX2_X1    g353(.I0(new_n488_), .I1(new_n481_), .S(new_n489_), .Z(new_n490_));
  MUX2_X1    g354(.I0(new_n490_), .I1(new_n486_), .S(new_n140_), .Z(new_n491_));
  NAND2_X1   g355(.A1(new_n491_), .A2(new_n139_), .ZN(new_n492_));
  MUX2_X1    g356(.I0(new_n483_), .I1(new_n487_), .S(new_n142_), .Z(new_n493_));
  MUX2_X1    g357(.I0(new_n485_), .I1(new_n493_), .S(new_n489_), .Z(new_n494_));
  NAND2_X1   g358(.A1(new_n140_), .A2(\A[18] ), .ZN(new_n495_));
  MUX2_X1    g359(.I0(new_n494_), .I1(new_n486_), .S(new_n495_), .Z(new_n496_));
  NAND2_X1   g360(.A1(new_n496_), .A2(\A[17] ), .ZN(new_n497_));
  AOI21_X1   g361(.A1(new_n497_), .A2(new_n492_), .B(\A[15] ), .ZN(new_n498_));
  MUX2_X1    g362(.I0(new_n488_), .I1(new_n493_), .S(new_n141_), .Z(new_n499_));
  MUX2_X1    g363(.I0(new_n490_), .I1(new_n499_), .S(new_n495_), .Z(new_n500_));
  NAND2_X1   g364(.A1(new_n139_), .A2(\A[16] ), .ZN(new_n501_));
  MUX2_X1    g365(.I0(new_n500_), .I1(new_n491_), .S(new_n501_), .Z(new_n502_));
  AOI21_X1   g366(.A1(\A[15] ), .A2(new_n502_), .B(new_n498_), .ZN(new_n503_));
  NOR2_X1    g367(.A1(new_n503_), .A2(\A[13] ), .ZN(new_n504_));
  INV_X1     g368(.I(\A[13] ), .ZN(new_n505_));
  MUX2_X1    g369(.I0(new_n494_), .I1(new_n499_), .S(new_n140_), .Z(new_n506_));
  MUX2_X1    g370(.I0(new_n500_), .I1(new_n506_), .S(new_n139_), .Z(new_n507_));
  INV_X1     g371(.I(\A[15] ), .ZN(new_n508_));
  NAND2_X1   g372(.A1(new_n508_), .A2(\A[14] ), .ZN(new_n509_));
  MUX2_X1    g373(.I0(new_n502_), .I1(new_n507_), .S(new_n509_), .Z(new_n510_));
  NOR2_X1    g374(.A1(new_n510_), .A2(new_n505_), .ZN(new_n511_));
  OAI21_X1   g375(.A1(new_n511_), .A2(new_n504_), .B(new_n138_), .ZN(new_n512_));
  MUX2_X1    g376(.I0(new_n496_), .I1(new_n491_), .S(new_n139_), .Z(new_n513_));
  MUX2_X1    g377(.I0(new_n496_), .I1(new_n506_), .S(new_n501_), .Z(new_n514_));
  MUX2_X1    g378(.I0(new_n514_), .I1(new_n513_), .S(new_n509_), .Z(new_n515_));
  NAND2_X1   g379(.A1(new_n505_), .A2(\A[12] ), .ZN(new_n516_));
  MUX2_X1    g380(.I0(new_n515_), .I1(new_n503_), .S(new_n516_), .Z(new_n517_));
  OAI21_X1   g381(.A1(new_n138_), .A2(new_n517_), .B(new_n512_), .ZN(new_n518_));
  NAND2_X1   g382(.A1(new_n518_), .A2(new_n137_), .ZN(new_n519_));
  NOR2_X1    g383(.A1(new_n514_), .A2(new_n508_), .ZN(new_n520_));
  OAI21_X1   g384(.A1(new_n520_), .A2(new_n498_), .B(new_n505_), .ZN(new_n521_));
  NAND2_X1   g385(.A1(new_n515_), .A2(\A[13] ), .ZN(new_n522_));
  NAND2_X1   g386(.A1(new_n522_), .A2(new_n521_), .ZN(new_n523_));
  INV_X1     g387(.I(\A[10] ), .ZN(new_n524_));
  NOR2_X1    g388(.A1(new_n524_), .A2(\A[11] ), .ZN(new_n525_));
  INV_X1     g389(.I(new_n525_), .ZN(new_n526_));
  MUX2_X1    g390(.I0(new_n517_), .I1(new_n523_), .S(new_n526_), .Z(new_n527_));
  NAND2_X1   g391(.A1(new_n527_), .A2(\A[9] ), .ZN(new_n528_));
  AOI21_X1   g392(.A1(new_n528_), .A2(new_n519_), .B(\A[7] ), .ZN(new_n529_));
  NOR2_X1    g393(.A1(new_n511_), .A2(new_n504_), .ZN(new_n530_));
  MUX2_X1    g394(.I0(new_n502_), .I1(new_n513_), .S(new_n508_), .Z(new_n531_));
  MUX2_X1    g395(.I0(new_n510_), .I1(new_n531_), .S(new_n516_), .Z(new_n532_));
  MUX2_X1    g396(.I0(new_n532_), .I1(new_n530_), .S(new_n526_), .Z(new_n533_));
  NAND2_X1   g397(.A1(new_n137_), .A2(\A[8] ), .ZN(new_n534_));
  MUX2_X1    g398(.I0(new_n533_), .I1(new_n518_), .S(new_n534_), .Z(new_n535_));
  AOI21_X1   g399(.A1(\A[7] ), .A2(new_n535_), .B(new_n529_), .ZN(new_n536_));
  INV_X1     g400(.I(\A[7] ), .ZN(new_n537_));
  AOI21_X1   g401(.A1(new_n522_), .A2(new_n521_), .B(\A[11] ), .ZN(new_n538_));
  AOI21_X1   g402(.A1(\A[11] ), .A2(new_n532_), .B(new_n538_), .ZN(new_n539_));
  NOR2_X1    g403(.A1(new_n539_), .A2(\A[9] ), .ZN(new_n540_));
  NOR2_X1    g404(.A1(new_n533_), .A2(new_n137_), .ZN(new_n541_));
  NOR2_X1    g405(.A1(new_n541_), .A2(new_n540_), .ZN(new_n542_));
  MUX2_X1    g406(.I0(new_n527_), .I1(new_n539_), .S(new_n534_), .Z(new_n543_));
  NAND4_X1   g407(.A1(new_n542_), .A2(new_n543_), .A3(\A[6] ), .A4(new_n537_), .ZN(new_n544_));
  NAND2_X1   g408(.A1(new_n528_), .A2(new_n519_), .ZN(new_n545_));
  NAND2_X1   g409(.A1(new_n537_), .A2(\A[6] ), .ZN(new_n546_));
  OAI21_X1   g410(.A1(new_n543_), .A2(new_n546_), .B(new_n545_), .ZN(new_n547_));
  INV_X1     g411(.I(\A[4] ), .ZN(new_n548_));
  NOR2_X1    g412(.A1(new_n548_), .A2(\A[5] ), .ZN(new_n549_));
  NAND4_X1   g413(.A1(new_n536_), .A2(new_n544_), .A3(new_n547_), .A4(new_n549_), .ZN(new_n550_));
  OAI21_X1   g414(.A1(new_n541_), .A2(new_n540_), .B(new_n537_), .ZN(new_n551_));
  NOR3_X1    g415(.A1(new_n532_), .A2(new_n523_), .A3(new_n526_), .ZN(new_n552_));
  AOI21_X1   g416(.A1(new_n532_), .A2(new_n525_), .B(new_n530_), .ZN(new_n553_));
  NOR4_X1    g417(.A1(new_n518_), .A2(new_n553_), .A3(new_n552_), .A4(new_n534_), .ZN(new_n554_));
  INV_X1     g418(.I(new_n534_), .ZN(new_n555_));
  AOI21_X1   g419(.A1(new_n527_), .A2(new_n555_), .B(new_n539_), .ZN(new_n556_));
  OAI21_X1   g420(.A1(new_n556_), .A2(new_n554_), .B(\A[7] ), .ZN(new_n557_));
  NAND2_X1   g421(.A1(new_n557_), .A2(new_n551_), .ZN(new_n558_));
  MUX2_X1    g422(.I0(new_n535_), .I1(new_n542_), .S(new_n546_), .Z(new_n559_));
  INV_X1     g423(.I(new_n549_), .ZN(new_n560_));
  OAI21_X1   g424(.A1(new_n559_), .A2(new_n560_), .B(new_n558_), .ZN(new_n561_));
  MUX2_X1    g425(.I0(new_n543_), .I1(new_n545_), .S(new_n546_), .Z(new_n562_));
  AOI21_X1   g426(.A1(new_n557_), .A2(new_n551_), .B(\A[5] ), .ZN(new_n563_));
  AOI21_X1   g427(.A1(new_n562_), .A2(\A[5] ), .B(new_n563_), .ZN(new_n564_));
  INV_X1     g428(.I(\A[2] ), .ZN(new_n565_));
  AOI21_X1   g429(.A1(new_n565_), .A2(\A[1] ), .B(\A[3] ), .ZN(new_n566_));
  INV_X1     g430(.I(new_n566_), .ZN(new_n567_));
  NAND4_X1   g431(.A1(new_n561_), .A2(new_n564_), .A3(new_n550_), .A4(new_n567_), .ZN(new_n568_));
  NOR3_X1    g432(.A1(new_n562_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n569_));
  AOI21_X1   g433(.A1(new_n562_), .A2(new_n549_), .B(new_n536_), .ZN(new_n570_));
  OAI22_X1   g434(.A1(new_n569_), .A2(new_n570_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n571_));
  NAND2_X1   g435(.A1(new_n571_), .A2(new_n568_), .ZN(\P[0] ));
  NOR2_X1    g436(.A1(\A[76] ), .A2(\A[77] ), .ZN(new_n573_));
  NOR2_X1    g437(.A1(\A[122] ), .A2(\A[123] ), .ZN(new_n574_));
  INV_X1     g438(.I(\A[120] ), .ZN(new_n575_));
  NOR2_X1    g439(.A1(\A[126] ), .A2(\A[127] ), .ZN(new_n576_));
  NAND4_X1   g440(.A1(new_n576_), .A2(new_n575_), .A3(new_n191_), .A4(new_n201_), .ZN(new_n577_));
  AOI21_X1   g441(.A1(\A[121] ), .A2(new_n574_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1   g442(.A1(new_n191_), .A2(new_n201_), .ZN(new_n579_));
  OAI21_X1   g443(.A1(new_n579_), .A2(new_n574_), .B(new_n576_), .ZN(new_n580_));
  NOR2_X1    g444(.A1(new_n580_), .A2(new_n575_), .ZN(new_n581_));
  XOR2_X1    g445(.A1(new_n581_), .A2(new_n578_), .Z(new_n582_));
  INV_X1     g446(.I(new_n582_), .ZN(new_n583_));
  NOR2_X1    g447(.A1(\A[116] ), .A2(\A[117] ), .ZN(new_n584_));
  NOR2_X1    g448(.A1(\A[118] ), .A2(\A[119] ), .ZN(new_n585_));
  MUX2_X1    g449(.I0(new_n580_), .I1(new_n582_), .S(new_n585_), .Z(new_n586_));
  MUX2_X1    g450(.I0(new_n586_), .I1(new_n583_), .S(new_n584_), .Z(new_n587_));
  NOR2_X1    g451(.A1(\A[112] ), .A2(\A[113] ), .ZN(new_n588_));
  NAND2_X1   g452(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR3_X1    g453(.A1(new_n586_), .A2(\A[114] ), .A3(\A[115] ), .ZN(new_n590_));
  NOR2_X1    g454(.A1(\A[114] ), .A2(\A[115] ), .ZN(new_n591_));
  NOR2_X1    g455(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1    g456(.A1(new_n592_), .A2(new_n590_), .Z(new_n593_));
  NOR2_X1    g457(.A1(new_n593_), .A2(new_n588_), .ZN(new_n594_));
  XNOR2_X1   g458(.A1(new_n594_), .A2(new_n589_), .ZN(new_n595_));
  NOR2_X1    g459(.A1(\A[108] ), .A2(\A[109] ), .ZN(new_n596_));
  INV_X1     g460(.I(new_n593_), .ZN(new_n597_));
  NOR2_X1    g461(.A1(\A[110] ), .A2(\A[111] ), .ZN(new_n598_));
  MUX2_X1    g462(.I0(new_n595_), .I1(new_n597_), .S(new_n598_), .Z(new_n599_));
  MUX2_X1    g463(.I0(new_n599_), .I1(new_n595_), .S(new_n596_), .Z(new_n600_));
  NOR2_X1    g464(.A1(\A[104] ), .A2(\A[105] ), .ZN(new_n601_));
  NOR2_X1    g465(.A1(\A[106] ), .A2(\A[107] ), .ZN(new_n602_));
  MUX2_X1    g466(.I0(new_n600_), .I1(new_n599_), .S(new_n602_), .Z(new_n603_));
  MUX2_X1    g467(.I0(new_n603_), .I1(new_n600_), .S(new_n601_), .Z(new_n604_));
  INV_X1     g468(.I(new_n604_), .ZN(new_n605_));
  NOR2_X1    g469(.A1(\A[100] ), .A2(\A[101] ), .ZN(new_n606_));
  NOR2_X1    g470(.A1(\A[102] ), .A2(\A[103] ), .ZN(new_n607_));
  INV_X1     g471(.I(new_n607_), .ZN(new_n608_));
  INV_X1     g472(.I(new_n603_), .ZN(new_n609_));
  NOR2_X1    g473(.A1(new_n609_), .A2(new_n608_), .ZN(new_n610_));
  AOI21_X1   g474(.A1(new_n604_), .A2(new_n608_), .B(new_n610_), .ZN(new_n611_));
  MUX2_X1    g475(.I0(new_n611_), .I1(new_n605_), .S(new_n606_), .Z(new_n612_));
  NOR2_X1    g476(.A1(\A[96] ), .A2(\A[97] ), .ZN(new_n613_));
  NOR2_X1    g477(.A1(\A[98] ), .A2(\A[99] ), .ZN(new_n614_));
  MUX2_X1    g478(.I0(new_n612_), .I1(new_n611_), .S(new_n614_), .Z(new_n615_));
  MUX2_X1    g479(.I0(new_n615_), .I1(new_n612_), .S(new_n613_), .Z(new_n616_));
  NOR2_X1    g480(.A1(\A[92] ), .A2(\A[93] ), .ZN(new_n617_));
  NOR2_X1    g481(.A1(\A[94] ), .A2(\A[95] ), .ZN(new_n618_));
  MUX2_X1    g482(.I0(new_n616_), .I1(new_n615_), .S(new_n618_), .Z(new_n619_));
  MUX2_X1    g483(.I0(new_n619_), .I1(new_n616_), .S(new_n617_), .Z(new_n620_));
  NOR2_X1    g484(.A1(\A[88] ), .A2(\A[89] ), .ZN(new_n621_));
  NOR2_X1    g485(.A1(\A[90] ), .A2(\A[91] ), .ZN(new_n622_));
  MUX2_X1    g486(.I0(new_n620_), .I1(new_n619_), .S(new_n622_), .Z(new_n623_));
  MUX2_X1    g487(.I0(new_n623_), .I1(new_n620_), .S(new_n621_), .Z(new_n624_));
  NOR2_X1    g488(.A1(\A[84] ), .A2(\A[85] ), .ZN(new_n625_));
  NOR2_X1    g489(.A1(\A[86] ), .A2(\A[87] ), .ZN(new_n626_));
  MUX2_X1    g490(.I0(new_n624_), .I1(new_n623_), .S(new_n626_), .Z(new_n627_));
  MUX2_X1    g491(.I0(new_n627_), .I1(new_n624_), .S(new_n625_), .Z(new_n628_));
  INV_X1     g492(.I(new_n628_), .ZN(new_n629_));
  NOR2_X1    g493(.A1(\A[80] ), .A2(\A[81] ), .ZN(new_n630_));
  NAND2_X1   g494(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1    g495(.A1(\A[82] ), .A2(\A[83] ), .ZN(new_n632_));
  MUX2_X1    g496(.I0(new_n628_), .I1(new_n627_), .S(new_n632_), .Z(new_n633_));
  NOR2_X1    g497(.A1(new_n633_), .A2(new_n630_), .ZN(new_n634_));
  XOR2_X1    g498(.A1(new_n634_), .A2(new_n631_), .Z(new_n635_));
  NAND2_X1   g499(.A1(new_n635_), .A2(new_n573_), .ZN(new_n636_));
  NOR2_X1    g500(.A1(\A[78] ), .A2(\A[79] ), .ZN(new_n637_));
  INV_X1     g501(.I(new_n637_), .ZN(new_n638_));
  NOR2_X1    g502(.A1(new_n633_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1     g503(.I(new_n639_), .ZN(new_n640_));
  OAI21_X1   g504(.A1(new_n635_), .A2(new_n637_), .B(new_n640_), .ZN(new_n641_));
  OAI21_X1   g505(.A1(new_n641_), .A2(new_n573_), .B(new_n636_), .ZN(new_n642_));
  NOR2_X1    g506(.A1(\A[72] ), .A2(\A[73] ), .ZN(new_n643_));
  INV_X1     g507(.I(new_n641_), .ZN(new_n644_));
  NOR2_X1    g508(.A1(\A[74] ), .A2(\A[75] ), .ZN(new_n645_));
  MUX2_X1    g509(.I0(new_n642_), .I1(new_n644_), .S(new_n645_), .Z(new_n646_));
  MUX2_X1    g510(.I0(new_n646_), .I1(new_n642_), .S(new_n643_), .Z(new_n647_));
  NOR2_X1    g511(.A1(\A[68] ), .A2(\A[69] ), .ZN(new_n648_));
  NOR2_X1    g512(.A1(\A[70] ), .A2(\A[71] ), .ZN(new_n649_));
  MUX2_X1    g513(.I0(new_n647_), .I1(new_n646_), .S(new_n649_), .Z(new_n650_));
  MUX2_X1    g514(.I0(new_n650_), .I1(new_n647_), .S(new_n648_), .Z(new_n651_));
  NOR2_X1    g515(.A1(\A[64] ), .A2(\A[65] ), .ZN(new_n652_));
  NOR2_X1    g516(.A1(\A[66] ), .A2(\A[67] ), .ZN(new_n653_));
  MUX2_X1    g517(.I0(new_n651_), .I1(new_n650_), .S(new_n653_), .Z(new_n654_));
  MUX2_X1    g518(.I0(new_n654_), .I1(new_n651_), .S(new_n652_), .Z(new_n655_));
  NOR2_X1    g519(.A1(\A[60] ), .A2(\A[61] ), .ZN(new_n656_));
  NOR2_X1    g520(.A1(\A[62] ), .A2(\A[63] ), .ZN(new_n657_));
  MUX2_X1    g521(.I0(new_n655_), .I1(new_n654_), .S(new_n657_), .Z(new_n658_));
  MUX2_X1    g522(.I0(new_n658_), .I1(new_n655_), .S(new_n656_), .Z(new_n659_));
  NOR2_X1    g523(.A1(\A[56] ), .A2(\A[57] ), .ZN(new_n660_));
  NOR2_X1    g524(.A1(\A[58] ), .A2(\A[59] ), .ZN(new_n661_));
  MUX2_X1    g525(.I0(new_n659_), .I1(new_n658_), .S(new_n661_), .Z(new_n662_));
  MUX2_X1    g526(.I0(new_n662_), .I1(new_n659_), .S(new_n660_), .Z(new_n663_));
  NOR2_X1    g527(.A1(\A[52] ), .A2(\A[53] ), .ZN(new_n664_));
  NOR2_X1    g528(.A1(\A[54] ), .A2(\A[55] ), .ZN(new_n665_));
  MUX2_X1    g529(.I0(new_n663_), .I1(new_n662_), .S(new_n665_), .Z(new_n666_));
  MUX2_X1    g530(.I0(new_n666_), .I1(new_n663_), .S(new_n664_), .Z(new_n667_));
  NOR2_X1    g531(.A1(\A[48] ), .A2(\A[49] ), .ZN(new_n668_));
  NOR2_X1    g532(.A1(\A[50] ), .A2(\A[51] ), .ZN(new_n669_));
  MUX2_X1    g533(.I0(new_n667_), .I1(new_n666_), .S(new_n669_), .Z(new_n670_));
  MUX2_X1    g534(.I0(new_n670_), .I1(new_n667_), .S(new_n668_), .Z(new_n671_));
  NOR2_X1    g535(.A1(\A[44] ), .A2(\A[45] ), .ZN(new_n672_));
  NOR2_X1    g536(.A1(\A[46] ), .A2(\A[47] ), .ZN(new_n673_));
  MUX2_X1    g537(.I0(new_n671_), .I1(new_n670_), .S(new_n673_), .Z(new_n674_));
  MUX2_X1    g538(.I0(new_n674_), .I1(new_n671_), .S(new_n672_), .Z(new_n675_));
  NOR2_X1    g539(.A1(\A[40] ), .A2(\A[41] ), .ZN(new_n676_));
  NOR2_X1    g540(.A1(\A[42] ), .A2(\A[43] ), .ZN(new_n677_));
  MUX2_X1    g541(.I0(new_n675_), .I1(new_n674_), .S(new_n677_), .Z(new_n678_));
  MUX2_X1    g542(.I0(new_n678_), .I1(new_n675_), .S(new_n676_), .Z(new_n679_));
  NOR2_X1    g543(.A1(\A[36] ), .A2(\A[37] ), .ZN(new_n680_));
  NOR2_X1    g544(.A1(\A[38] ), .A2(\A[39] ), .ZN(new_n681_));
  MUX2_X1    g545(.I0(new_n679_), .I1(new_n678_), .S(new_n681_), .Z(new_n682_));
  MUX2_X1    g546(.I0(new_n682_), .I1(new_n679_), .S(new_n680_), .Z(new_n683_));
  NOR2_X1    g547(.A1(\A[32] ), .A2(\A[33] ), .ZN(new_n684_));
  NOR2_X1    g548(.A1(\A[34] ), .A2(\A[35] ), .ZN(new_n685_));
  MUX2_X1    g549(.I0(new_n683_), .I1(new_n682_), .S(new_n685_), .Z(new_n686_));
  MUX2_X1    g550(.I0(new_n686_), .I1(new_n683_), .S(new_n684_), .Z(new_n687_));
  NOR2_X1    g551(.A1(\A[28] ), .A2(\A[29] ), .ZN(new_n688_));
  NOR2_X1    g552(.A1(\A[30] ), .A2(\A[31] ), .ZN(new_n689_));
  MUX2_X1    g553(.I0(new_n687_), .I1(new_n686_), .S(new_n689_), .Z(new_n690_));
  MUX2_X1    g554(.I0(new_n690_), .I1(new_n687_), .S(new_n688_), .Z(new_n691_));
  NOR2_X1    g555(.A1(\A[24] ), .A2(\A[25] ), .ZN(new_n692_));
  NOR2_X1    g556(.A1(\A[26] ), .A2(\A[27] ), .ZN(new_n693_));
  MUX2_X1    g557(.I0(new_n691_), .I1(new_n690_), .S(new_n693_), .Z(new_n694_));
  MUX2_X1    g558(.I0(new_n694_), .I1(new_n691_), .S(new_n692_), .Z(new_n695_));
  NOR2_X1    g559(.A1(\A[20] ), .A2(\A[21] ), .ZN(new_n696_));
  NOR2_X1    g560(.A1(\A[22] ), .A2(\A[23] ), .ZN(new_n697_));
  MUX2_X1    g561(.I0(new_n695_), .I1(new_n694_), .S(new_n697_), .Z(new_n698_));
  MUX2_X1    g562(.I0(new_n698_), .I1(new_n695_), .S(new_n696_), .Z(new_n699_));
  NOR2_X1    g563(.A1(\A[16] ), .A2(\A[17] ), .ZN(new_n700_));
  NOR2_X1    g564(.A1(\A[18] ), .A2(\A[19] ), .ZN(new_n701_));
  MUX2_X1    g565(.I0(new_n699_), .I1(new_n698_), .S(new_n701_), .Z(new_n702_));
  MUX2_X1    g566(.I0(new_n702_), .I1(new_n699_), .S(new_n700_), .Z(new_n703_));
  NOR2_X1    g567(.A1(\A[12] ), .A2(\A[13] ), .ZN(new_n704_));
  NOR2_X1    g568(.A1(\A[14] ), .A2(\A[15] ), .ZN(new_n705_));
  MUX2_X1    g569(.I0(new_n703_), .I1(new_n702_), .S(new_n705_), .Z(new_n706_));
  MUX2_X1    g570(.I0(new_n706_), .I1(new_n703_), .S(new_n704_), .Z(new_n707_));
  INV_X1     g571(.I(new_n707_), .ZN(new_n708_));
  NOR2_X1    g572(.A1(\A[8] ), .A2(\A[9] ), .ZN(new_n709_));
  NOR2_X1    g573(.A1(\A[10] ), .A2(\A[11] ), .ZN(new_n710_));
  INV_X1     g574(.I(new_n710_), .ZN(new_n711_));
  OR2_X2     g575(.A1(new_n706_), .A2(new_n711_), .Z(new_n712_));
  OAI21_X1   g576(.A1(new_n707_), .A2(new_n710_), .B(new_n712_), .ZN(new_n713_));
  MUX2_X1    g577(.I0(new_n713_), .I1(new_n708_), .S(new_n709_), .Z(new_n714_));
  NOR2_X1    g578(.A1(\A[6] ), .A2(\A[7] ), .ZN(new_n715_));
  MUX2_X1    g579(.I0(new_n714_), .I1(new_n713_), .S(new_n715_), .Z(new_n716_));
  NOR2_X1    g580(.A1(\A[2] ), .A2(\A[3] ), .ZN(new_n717_));
  NOR3_X1    g581(.A1(new_n717_), .A2(\A[4] ), .A3(\A[5] ), .ZN(new_n718_));
  MUX2_X1    g582(.I0(new_n716_), .I1(new_n714_), .S(new_n718_), .Z(\P[1] ));
  NAND2_X1   g583(.A1(new_n700_), .A2(new_n701_), .ZN(new_n720_));
  INV_X1     g584(.I(new_n720_), .ZN(new_n721_));
  NAND2_X1   g585(.A1(new_n692_), .A2(new_n693_), .ZN(new_n722_));
  INV_X1     g586(.I(new_n722_), .ZN(new_n723_));
  NAND2_X1   g587(.A1(new_n684_), .A2(new_n685_), .ZN(new_n724_));
  INV_X1     g588(.I(new_n724_), .ZN(new_n725_));
  NAND2_X1   g589(.A1(new_n676_), .A2(new_n677_), .ZN(new_n726_));
  INV_X1     g590(.I(new_n726_), .ZN(new_n727_));
  NAND2_X1   g591(.A1(new_n668_), .A2(new_n669_), .ZN(new_n728_));
  INV_X1     g592(.I(new_n728_), .ZN(new_n729_));
  NAND2_X1   g593(.A1(new_n660_), .A2(new_n661_), .ZN(new_n730_));
  INV_X1     g594(.I(new_n730_), .ZN(new_n731_));
  NAND2_X1   g595(.A1(new_n652_), .A2(new_n653_), .ZN(new_n732_));
  INV_X1     g596(.I(new_n732_), .ZN(new_n733_));
  NAND2_X1   g597(.A1(new_n643_), .A2(new_n645_), .ZN(new_n734_));
  INV_X1     g598(.I(new_n734_), .ZN(new_n735_));
  NAND2_X1   g599(.A1(new_n630_), .A2(new_n632_), .ZN(new_n736_));
  INV_X1     g600(.I(new_n736_), .ZN(new_n737_));
  NAND2_X1   g601(.A1(new_n621_), .A2(new_n622_), .ZN(new_n738_));
  INV_X1     g602(.I(new_n738_), .ZN(new_n739_));
  NAND2_X1   g603(.A1(new_n613_), .A2(new_n614_), .ZN(new_n740_));
  INV_X1     g604(.I(new_n740_), .ZN(new_n741_));
  NAND2_X1   g605(.A1(new_n601_), .A2(new_n602_), .ZN(new_n742_));
  INV_X1     g606(.I(new_n742_), .ZN(new_n743_));
  NAND3_X1   g607(.A1(new_n574_), .A2(new_n575_), .A3(new_n185_), .ZN(new_n744_));
  NAND2_X1   g608(.A1(new_n584_), .A2(new_n585_), .ZN(new_n745_));
  INV_X1     g609(.I(new_n745_), .ZN(new_n746_));
  NOR2_X1    g610(.A1(new_n746_), .A2(new_n216_), .ZN(new_n747_));
  NOR3_X1    g611(.A1(new_n579_), .A2(\A[126] ), .A3(\A[127] ), .ZN(new_n748_));
  OAI21_X1   g612(.A1(new_n747_), .A2(new_n744_), .B(new_n748_), .ZN(new_n749_));
  NOR3_X1    g613(.A1(\A[112] ), .A2(\A[113] ), .A3(\A[114] ), .ZN(new_n750_));
  OAI21_X1   g614(.A1(new_n744_), .A2(new_n745_), .B(new_n748_), .ZN(new_n751_));
  MUX2_X1    g615(.I0(new_n751_), .I1(new_n749_), .S(new_n750_), .Z(new_n752_));
  NOR2_X1    g616(.A1(new_n752_), .A2(new_n743_), .ZN(new_n753_));
  NAND2_X1   g617(.A1(new_n596_), .A2(new_n598_), .ZN(new_n754_));
  INV_X1     g618(.I(new_n754_), .ZN(new_n755_));
  NOR2_X1    g619(.A1(new_n751_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1   g620(.A1(new_n752_), .A2(new_n755_), .B(new_n756_), .ZN(new_n757_));
  AOI21_X1   g621(.A1(new_n757_), .A2(new_n743_), .B(new_n753_), .ZN(new_n758_));
  NOR2_X1    g622(.A1(new_n758_), .A2(new_n741_), .ZN(new_n759_));
  NAND2_X1   g623(.A1(new_n606_), .A2(new_n607_), .ZN(new_n760_));
  NOR2_X1    g624(.A1(new_n757_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1   g625(.A1(new_n758_), .A2(new_n760_), .B(new_n761_), .ZN(new_n762_));
  AOI21_X1   g626(.A1(new_n762_), .A2(new_n741_), .B(new_n759_), .ZN(new_n763_));
  NOR2_X1    g627(.A1(new_n763_), .A2(new_n739_), .ZN(new_n764_));
  NAND2_X1   g628(.A1(new_n617_), .A2(new_n618_), .ZN(new_n765_));
  INV_X1     g629(.I(new_n765_), .ZN(new_n766_));
  NOR2_X1    g630(.A1(new_n762_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1   g631(.A1(new_n763_), .A2(new_n766_), .B(new_n767_), .ZN(new_n768_));
  AOI21_X1   g632(.A1(new_n768_), .A2(new_n739_), .B(new_n764_), .ZN(new_n769_));
  NOR2_X1    g633(.A1(new_n769_), .A2(new_n737_), .ZN(new_n770_));
  NAND2_X1   g634(.A1(new_n625_), .A2(new_n626_), .ZN(new_n771_));
  INV_X1     g635(.I(new_n771_), .ZN(new_n772_));
  NOR2_X1    g636(.A1(new_n768_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1   g637(.A1(new_n769_), .A2(new_n772_), .B(new_n773_), .ZN(new_n774_));
  AOI21_X1   g638(.A1(new_n774_), .A2(new_n737_), .B(new_n770_), .ZN(new_n775_));
  NOR2_X1    g639(.A1(new_n775_), .A2(new_n735_), .ZN(new_n776_));
  INV_X1     g640(.I(new_n573_), .ZN(new_n777_));
  NOR2_X1    g641(.A1(new_n777_), .A2(new_n638_), .ZN(new_n778_));
  INV_X1     g642(.I(new_n778_), .ZN(new_n779_));
  NOR2_X1    g643(.A1(new_n774_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1   g644(.A1(new_n775_), .A2(new_n779_), .B(new_n780_), .ZN(new_n781_));
  AOI21_X1   g645(.A1(new_n781_), .A2(new_n735_), .B(new_n776_), .ZN(new_n782_));
  NOR2_X1    g646(.A1(new_n782_), .A2(new_n733_), .ZN(new_n783_));
  NAND2_X1   g647(.A1(new_n648_), .A2(new_n649_), .ZN(new_n784_));
  INV_X1     g648(.I(new_n784_), .ZN(new_n785_));
  NOR2_X1    g649(.A1(new_n781_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1   g650(.A1(new_n782_), .A2(new_n785_), .B(new_n786_), .ZN(new_n787_));
  AOI21_X1   g651(.A1(new_n787_), .A2(new_n733_), .B(new_n783_), .ZN(new_n788_));
  NOR2_X1    g652(.A1(new_n788_), .A2(new_n731_), .ZN(new_n789_));
  NAND2_X1   g653(.A1(new_n656_), .A2(new_n657_), .ZN(new_n790_));
  INV_X1     g654(.I(new_n790_), .ZN(new_n791_));
  NOR2_X1    g655(.A1(new_n787_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1   g656(.A1(new_n788_), .A2(new_n791_), .B(new_n792_), .ZN(new_n793_));
  AOI21_X1   g657(.A1(new_n793_), .A2(new_n731_), .B(new_n789_), .ZN(new_n794_));
  NOR2_X1    g658(.A1(new_n794_), .A2(new_n729_), .ZN(new_n795_));
  NAND2_X1   g659(.A1(new_n664_), .A2(new_n665_), .ZN(new_n796_));
  INV_X1     g660(.I(new_n796_), .ZN(new_n797_));
  NOR2_X1    g661(.A1(new_n793_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1   g662(.A1(new_n794_), .A2(new_n797_), .B(new_n798_), .ZN(new_n799_));
  AOI21_X1   g663(.A1(new_n799_), .A2(new_n729_), .B(new_n795_), .ZN(new_n800_));
  NOR2_X1    g664(.A1(new_n800_), .A2(new_n727_), .ZN(new_n801_));
  NAND2_X1   g665(.A1(new_n672_), .A2(new_n673_), .ZN(new_n802_));
  INV_X1     g666(.I(new_n802_), .ZN(new_n803_));
  NOR2_X1    g667(.A1(new_n799_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1   g668(.A1(new_n800_), .A2(new_n803_), .B(new_n804_), .ZN(new_n805_));
  AOI21_X1   g669(.A1(new_n805_), .A2(new_n727_), .B(new_n801_), .ZN(new_n806_));
  NOR2_X1    g670(.A1(new_n806_), .A2(new_n725_), .ZN(new_n807_));
  NAND2_X1   g671(.A1(new_n680_), .A2(new_n681_), .ZN(new_n808_));
  INV_X1     g672(.I(new_n808_), .ZN(new_n809_));
  NOR2_X1    g673(.A1(new_n805_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1   g674(.A1(new_n806_), .A2(new_n809_), .B(new_n810_), .ZN(new_n811_));
  AOI21_X1   g675(.A1(new_n811_), .A2(new_n725_), .B(new_n807_), .ZN(new_n812_));
  NOR2_X1    g676(.A1(new_n812_), .A2(new_n723_), .ZN(new_n813_));
  NAND2_X1   g677(.A1(new_n688_), .A2(new_n689_), .ZN(new_n814_));
  INV_X1     g678(.I(new_n814_), .ZN(new_n815_));
  NOR2_X1    g679(.A1(new_n811_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1   g680(.A1(new_n812_), .A2(new_n815_), .B(new_n816_), .ZN(new_n817_));
  AOI21_X1   g681(.A1(new_n817_), .A2(new_n723_), .B(new_n813_), .ZN(new_n818_));
  NOR2_X1    g682(.A1(new_n818_), .A2(new_n721_), .ZN(new_n819_));
  NAND2_X1   g683(.A1(new_n696_), .A2(new_n697_), .ZN(new_n820_));
  INV_X1     g684(.I(new_n820_), .ZN(new_n821_));
  NOR2_X1    g685(.A1(new_n817_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1   g686(.A1(new_n818_), .A2(new_n821_), .B(new_n822_), .ZN(new_n823_));
  AOI21_X1   g687(.A1(new_n823_), .A2(new_n721_), .B(new_n819_), .ZN(new_n824_));
  NAND2_X1   g688(.A1(new_n704_), .A2(new_n705_), .ZN(new_n825_));
  INV_X1     g689(.I(new_n825_), .ZN(new_n826_));
  NAND2_X1   g690(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1   g691(.A1(new_n823_), .A2(new_n826_), .B(new_n827_), .ZN(new_n828_));
  NOR4_X1    g692(.A1(\A[4] ), .A2(\A[5] ), .A3(\A[6] ), .A4(\A[7] ), .ZN(new_n829_));
  INV_X1     g693(.I(new_n829_), .ZN(new_n830_));
  NOR3_X1    g694(.A1(new_n711_), .A2(\A[8] ), .A3(\A[9] ), .ZN(new_n831_));
  NAND2_X1   g695(.A1(new_n831_), .A2(new_n830_), .ZN(new_n832_));
  MUX2_X1    g696(.I0(new_n824_), .I1(new_n828_), .S(new_n832_), .Z(\P[2] ));
  NOR2_X1    g697(.A1(new_n725_), .A2(new_n809_), .ZN(new_n834_));
  INV_X1     g698(.I(new_n834_), .ZN(new_n835_));
  AOI21_X1   g699(.A1(new_n588_), .A2(new_n591_), .B(new_n746_), .ZN(new_n836_));
  NOR2_X1    g700(.A1(new_n743_), .A2(new_n755_), .ZN(new_n837_));
  INV_X1     g701(.I(new_n837_), .ZN(new_n838_));
  OAI21_X1   g702(.A1(new_n838_), .A2(new_n259_), .B(new_n836_), .ZN(new_n839_));
  NOR4_X1    g703(.A1(new_n744_), .A2(\A[126] ), .A3(new_n579_), .A4(\A[127] ), .ZN(new_n840_));
  NAND2_X1   g704(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NOR4_X1    g705(.A1(new_n741_), .A2(\A[100] ), .A3(\A[101] ), .A4(\A[102] ), .ZN(new_n842_));
  INV_X1     g706(.I(new_n840_), .ZN(new_n843_));
  AOI21_X1   g707(.A1(new_n838_), .A2(new_n836_), .B(new_n843_), .ZN(new_n844_));
  INV_X1     g708(.I(new_n844_), .ZN(new_n845_));
  MUX2_X1    g709(.I0(new_n845_), .I1(new_n841_), .S(new_n842_), .Z(new_n846_));
  NOR2_X1    g710(.A1(new_n737_), .A2(new_n772_), .ZN(new_n847_));
  INV_X1     g711(.I(new_n847_), .ZN(new_n848_));
  NOR2_X1    g712(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1    g713(.A1(new_n739_), .A2(new_n766_), .ZN(new_n850_));
  INV_X1     g714(.I(new_n850_), .ZN(new_n851_));
  NAND2_X1   g715(.A1(new_n846_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1   g716(.A1(new_n845_), .A2(new_n851_), .B(new_n852_), .ZN(new_n853_));
  NOR2_X1    g717(.A1(new_n853_), .A2(new_n847_), .ZN(new_n854_));
  NOR2_X1    g718(.A1(new_n854_), .A2(new_n849_), .ZN(new_n855_));
  NOR2_X1    g719(.A1(new_n733_), .A2(new_n785_), .ZN(new_n856_));
  INV_X1     g720(.I(new_n856_), .ZN(new_n857_));
  NOR2_X1    g721(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1    g722(.A1(new_n779_), .A2(new_n735_), .ZN(new_n859_));
  NAND2_X1   g723(.A1(new_n853_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1     g724(.I(new_n859_), .ZN(new_n861_));
  NAND2_X1   g725(.A1(new_n855_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1   g726(.A1(new_n862_), .A2(new_n860_), .ZN(new_n863_));
  NOR2_X1    g727(.A1(new_n863_), .A2(new_n856_), .ZN(new_n864_));
  NOR2_X1    g728(.A1(new_n864_), .A2(new_n858_), .ZN(new_n865_));
  NOR2_X1    g729(.A1(new_n729_), .A2(new_n797_), .ZN(new_n866_));
  INV_X1     g730(.I(new_n866_), .ZN(new_n867_));
  NOR2_X1    g731(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1    g732(.A1(new_n731_), .A2(new_n791_), .ZN(new_n869_));
  NAND2_X1   g733(.A1(new_n863_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1     g734(.I(new_n869_), .ZN(new_n871_));
  NAND2_X1   g735(.A1(new_n865_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1   g736(.A1(new_n872_), .A2(new_n870_), .ZN(new_n873_));
  NOR2_X1    g737(.A1(new_n873_), .A2(new_n866_), .ZN(new_n874_));
  NOR2_X1    g738(.A1(new_n874_), .A2(new_n868_), .ZN(new_n875_));
  NOR2_X1    g739(.A1(new_n875_), .A2(new_n835_), .ZN(new_n876_));
  NOR2_X1    g740(.A1(new_n727_), .A2(new_n803_), .ZN(new_n877_));
  NOR3_X1    g741(.A1(new_n874_), .A2(new_n868_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1   g742(.A1(new_n873_), .A2(new_n877_), .B(new_n878_), .ZN(new_n879_));
  AOI21_X1   g743(.A1(new_n879_), .A2(new_n835_), .B(new_n876_), .ZN(new_n880_));
  NOR2_X1    g744(.A1(new_n723_), .A2(new_n815_), .ZN(new_n881_));
  INV_X1     g745(.I(new_n881_), .ZN(new_n882_));
  NAND2_X1   g746(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1   g747(.A1(new_n879_), .A2(new_n882_), .B(new_n883_), .ZN(new_n884_));
  NAND2_X1   g748(.A1(new_n831_), .A2(new_n825_), .ZN(new_n885_));
  NOR2_X1    g749(.A1(new_n721_), .A2(new_n821_), .ZN(new_n886_));
  NAND2_X1   g750(.A1(new_n886_), .A2(new_n885_), .ZN(new_n887_));
  MUX2_X1    g751(.I0(new_n880_), .I1(new_n884_), .S(new_n887_), .Z(\P[3] ));
  NOR3_X1    g752(.A1(new_n838_), .A2(new_n741_), .A3(new_n760_), .ZN(new_n889_));
  NOR2_X1    g753(.A1(new_n848_), .A2(new_n851_), .ZN(new_n890_));
  INV_X1     g754(.I(new_n890_), .ZN(new_n891_));
  OAI21_X1   g755(.A1(new_n891_), .A2(new_n170_), .B(new_n889_), .ZN(new_n892_));
  INV_X1     g756(.I(new_n836_), .ZN(new_n893_));
  NOR2_X1    g757(.A1(new_n893_), .A2(new_n843_), .ZN(new_n894_));
  NAND2_X1   g758(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NOR4_X1    g759(.A1(new_n857_), .A2(\A[78] ), .A3(new_n735_), .A4(new_n777_), .ZN(new_n896_));
  INV_X1     g760(.I(new_n894_), .ZN(new_n897_));
  AOI21_X1   g761(.A1(new_n891_), .A2(new_n889_), .B(new_n897_), .ZN(new_n898_));
  INV_X1     g762(.I(new_n898_), .ZN(new_n899_));
  MUX2_X1    g763(.I0(new_n899_), .I1(new_n895_), .S(new_n896_), .Z(new_n900_));
  NOR2_X1    g764(.A1(new_n867_), .A2(new_n871_), .ZN(new_n901_));
  INV_X1     g765(.I(new_n901_), .ZN(new_n902_));
  NAND2_X1   g766(.A1(new_n900_), .A2(new_n902_), .ZN(new_n903_));
  OAI21_X1   g767(.A1(new_n899_), .A2(new_n902_), .B(new_n903_), .ZN(new_n904_));
  NAND2_X1   g768(.A1(new_n834_), .A2(new_n877_), .ZN(new_n905_));
  AOI21_X1   g769(.A1(new_n881_), .A2(new_n886_), .B(new_n905_), .ZN(new_n906_));
  MUX2_X1    g770(.I0(new_n904_), .I1(new_n900_), .S(new_n906_), .Z(\P[4] ));
  AND2_X2    g771(.A1(new_n894_), .A2(new_n889_), .Z(new_n908_));
  NOR2_X1    g772(.A1(new_n902_), .A2(new_n905_), .ZN(new_n909_));
  NOR3_X1    g773(.A1(new_n891_), .A2(new_n857_), .A3(new_n861_), .ZN(new_n910_));
  INV_X1     g774(.I(new_n910_), .ZN(new_n911_));
  OAI21_X1   g775(.A1(new_n911_), .A2(new_n909_), .B(new_n908_), .ZN(\P[5] ));
  NAND2_X1   g776(.A1(new_n910_), .A2(new_n908_), .ZN(\P[6] ));
  NAND2_X1   g777(.A1(new_n881_), .A2(new_n886_), .ZN(new_n914_));
  NOR2_X1    g778(.A1(\A[0] ), .A2(\A[1] ), .ZN(new_n915_));
  NAND2_X1   g779(.A1(new_n717_), .A2(new_n915_), .ZN(new_n916_));
  NOR4_X1    g780(.A1(new_n914_), .A2(new_n830_), .A3(new_n885_), .A4(new_n916_), .ZN(new_n917_));
  NAND4_X1   g781(.A1(new_n910_), .A2(new_n908_), .A3(new_n909_), .A4(new_n917_), .ZN(F));
endmodule


