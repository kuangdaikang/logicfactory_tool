// Benchmark "testing" written by ABC on Fri Feb 25 15:12:33 2022

module 25_4 ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A139  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A139;
  wire new_n27_, new_n28_, new_n29_, new_n30_, new_n31_, new_n32_, new_n33_,
    new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_,
    new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_,
    new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_,
    new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_,
    new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_,
    new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_,
    new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_,
    new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_,
    new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_,
    new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_,
    new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_,
    new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_,
    new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_,
    new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_,
    new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_,
    new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_,
    new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_,
    new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_,
    new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_,
    new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_,
    new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_,
    new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_,
    new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_,
    new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_,
    new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_,
    new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_,
    new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_,
    new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_,
    new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_,
    new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_,
    new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_,
    new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_,
    new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_,
    new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_,
    new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_,
    new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_,
    new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_,
    new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_,
    new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_,
    new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_,
    new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_,
    new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_,
    new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_,
    new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_,
    new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_,
    new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_,
    new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_,
    new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_,
    new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_,
    new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_,
    new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_,
    new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_,
    new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_,
    new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_,
    new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_,
    new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_,
    new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_,
    new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_,
    new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_,
    new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_,
    new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_,
    new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_,
    new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_,
    new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_,
    new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_,
    new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_,
    new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_,
    new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_,
    new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_,
    new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_,
    new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_,
    new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_,
    new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_,
    new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_,
    new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_,
    new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_,
    new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_,
    new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_,
    new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_,
    new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_,
    new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_,
    new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_,
    new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_,
    new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_,
    new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_,
    new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_,
    new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_,
    new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_,
    new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_,
    new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_,
    new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_,
    new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_,
    new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_,
    new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_,
    new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_,
    new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_,
    new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_,
    new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_,
    new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_,
    new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_,
    new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_,
    new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_,
    new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_,
    new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_,
    new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_,
    new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_,
    new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_,
    new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_,
    new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_,
    new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_,
    new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_,
    new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_,
    new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_,
    new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_,
    new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_,
    new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_,
    new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_,
    new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_,
    new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_,
    new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_,
    new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_,
    new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_,
    new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_,
    new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_,
    new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_,
    new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_,
    new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_,
    new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_,
    new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_,
    new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_,
    new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_,
    new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_,
    new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_,
    new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_,
    new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_,
    new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_,
    new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_,
    new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_,
    new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_,
    new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_,
    new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_,
    new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_,
    new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_,
    new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_,
    new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_,
    new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_,
    new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_,
    new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_,
    new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_,
    new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_,
    new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_,
    new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_,
    new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_,
    new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_,
    new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_,
    new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_,
    new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_,
    new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_,
    new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_,
    new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_,
    new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_,
    new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_,
    new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_,
    new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_,
    new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_,
    new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_,
    new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_,
    new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_,
    new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_,
    new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_,
    new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_,
    new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_,
    new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_,
    new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_,
    new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_,
    new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_,
    new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_,
    new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_,
    new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_,
    new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_,
    new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_,
    new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_,
    new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_,
    new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_,
    new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_,
    new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_,
    new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_,
    new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_,
    new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_,
    new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_,
    new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_,
    new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_,
    new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_,
    new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_,
    new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_,
    new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_,
    new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_,
    new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_,
    new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_,
    new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_,
    new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_,
    new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_,
    new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_,
    new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_,
    new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_,
    new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_,
    new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_,
    new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_,
    new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_,
    new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_,
    new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_,
    new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_,
    new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_,
    new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_,
    new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_,
    new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_,
    new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_,
    new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_,
    new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_,
    new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_,
    new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_,
    new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_,
    new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_,
    new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_,
    new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_,
    new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_,
    new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_,
    new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_,
    new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_,
    new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_,
    new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_,
    new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_,
    new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_,
    new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_,
    new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_,
    new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_,
    new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_,
    new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_,
    new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_,
    new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_,
    new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_,
    new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_,
    new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_,
    new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_,
    new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_,
    new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_,
    new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_,
    new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_,
    new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_,
    new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_,
    new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_,
    new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_,
    new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_,
    new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_,
    new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_,
    new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_,
    new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_,
    new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_,
    new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_,
    new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_,
    new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_,
    new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_,
    new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_,
    new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_,
    new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_,
    new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_,
    new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_,
    new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_,
    new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_,
    new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_,
    new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_,
    new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_,
    new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_,
    new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_,
    new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_,
    new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_,
    new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_,
    new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_,
    new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_,
    new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_,
    new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_,
    new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_,
    new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_,
    new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_,
    new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_,
    new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_,
    new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_,
    new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_,
    new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_,
    new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_,
    new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_,
    new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_,
    new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_,
    new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_,
    new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_,
    new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_,
    new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_,
    new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_,
    new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_,
    new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_,
    new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_,
    new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_,
    new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_,
    new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_,
    new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_,
    new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_,
    new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_,
    new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_,
    new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_,
    new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_,
    new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_,
    new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_,
    new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_,
    new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_,
    new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_,
    new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_,
    new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_,
    new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_,
    new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_,
    new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_,
    new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_,
    new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_,
    new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_,
    new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_,
    new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_,
    new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_,
    new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_,
    new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_,
    new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_,
    new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_,
    new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_,
    new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_,
    new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_,
    new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_,
    new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_,
    new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_,
    new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_,
    new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_,
    new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_,
    new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_,
    new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_,
    new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_,
    new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_,
    new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_,
    new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_,
    new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_,
    new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_,
    new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_,
    new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_,
    new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_,
    new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_,
    new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_,
    new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_,
    new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_,
    new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_,
    new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_,
    new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_,
    new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_,
    new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_,
    new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_,
    new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_,
    new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_,
    new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_,
    new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_,
    new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_,
    new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_,
    new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_,
    new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_,
    new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_,
    new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_,
    new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_,
    new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_,
    new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_,
    new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_,
    new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_,
    new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_,
    new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_,
    new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_,
    new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_,
    new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_,
    new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_,
    new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_,
    new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_,
    new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_,
    new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_,
    new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_,
    new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_,
    new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_,
    new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_,
    new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_,
    new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_,
    new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_,
    new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_,
    new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_,
    new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_,
    new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_,
    new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_,
    new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_,
    new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_,
    new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_,
    new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_,
    new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_,
    new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_,
    new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_,
    new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_,
    new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_,
    new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_,
    new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_,
    new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_,
    new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_,
    new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_,
    new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_,
    new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_,
    new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_,
    new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_,
    new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_,
    new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_,
    new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_,
    new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_,
    new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_,
    new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_,
    new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_,
    new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_,
    new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_,
    new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_,
    new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_,
    new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_,
    new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_,
    new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_,
    new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_,
    new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_,
    new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_,
    new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_,
    new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_,
    new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_,
    new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_,
    new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_,
    new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_,
    new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_,
    new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_,
    new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_,
    new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_,
    new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_,
    new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_,
    new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_,
    new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_,
    new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_,
    new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_,
    new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_,
    new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_,
    new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_,
    new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_,
    new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_,
    new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_,
    new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_,
    new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_,
    new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_,
    new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_,
    new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_,
    new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_,
    new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_,
    new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_,
    new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_,
    new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_,
    new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_,
    new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_,
    new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_,
    new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_,
    new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_,
    new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_,
    new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_,
    new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_,
    new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_,
    new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_,
    new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_,
    new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_,
    new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_,
    new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_,
    new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_,
    new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_,
    new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_,
    new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_,
    new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_,
    new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_,
    new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_,
    new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_,
    new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_,
    new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_,
    new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_,
    new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_,
    new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_,
    new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_,
    new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_,
    new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_,
    new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_,
    new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_,
    new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_,
    new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_,
    new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_,
    new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_,
    new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_,
    new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_,
    new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_,
    new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_,
    new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_,
    new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_,
    new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_,
    new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_,
    new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_,
    new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_,
    new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_,
    new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_,
    new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_,
    new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_,
    new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_,
    new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_,
    new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_,
    new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_,
    new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_,
    new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_,
    new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_,
    new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_,
    new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_,
    new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_,
    new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_,
    new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_,
    new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_,
    new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_,
    new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_,
    new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_,
    new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_,
    new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_,
    new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_,
    new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_,
    new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_,
    new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_,
    new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_,
    new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_,
    new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_,
    new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_,
    new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_,
    new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_,
    new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_,
    new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_,
    new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_,
    new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_,
    new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_,
    new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_,
    new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_,
    new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_,
    new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_,
    new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_,
    new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_,
    new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_,
    new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_,
    new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_,
    new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_,
    new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_,
    new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_,
    new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_,
    new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_,
    new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_,
    new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_,
    new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_,
    new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_,
    new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_,
    new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_,
    new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_,
    new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_,
    new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_,
    new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_,
    new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_,
    new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_,
    new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_,
    new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_,
    new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_,
    new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_,
    new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_,
    new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_,
    new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_,
    new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_,
    new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_,
    new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_,
    new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_,
    new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_,
    new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_,
    new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_,
    new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_,
    new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_,
    new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_,
    new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_,
    new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_,
    new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_,
    new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_,
    new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_,
    new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_,
    new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_,
    new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_,
    new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_,
    new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_,
    new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_,
    new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_,
    new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_,
    new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_,
    new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_,
    new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_,
    new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_,
    new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_,
    new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_,
    new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_,
    new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_,
    new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_,
    new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_,
    new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_,
    new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_,
    new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_,
    new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_,
    new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_,
    new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_,
    new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_,
    new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_,
    new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_,
    new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_,
    new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_,
    new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_,
    new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_,
    new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_,
    new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_,
    new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_,
    new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_,
    new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_,
    new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_,
    new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_,
    new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_,
    new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_,
    new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_,
    new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_,
    new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_,
    new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_,
    new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_,
    new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_,
    new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_,
    new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_,
    new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_,
    new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_,
    new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_,
    new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_,
    new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_,
    new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_,
    new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_,
    new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_,
    new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_,
    new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_,
    new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_,
    new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_,
    new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_,
    new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_,
    new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_,
    new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_,
    new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_,
    new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_,
    new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_,
    new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_,
    new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_,
    new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_,
    new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_,
    new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_,
    new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_,
    new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_,
    new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_,
    new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_,
    new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_,
    new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_,
    new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_,
    new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_,
    new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_,
    new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_,
    new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_,
    new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_,
    new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_,
    new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_,
    new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_,
    new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_,
    new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_,
    new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_,
    new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_,
    new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_,
    new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_,
    new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_,
    new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_,
    new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_,
    new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_,
    new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_,
    new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_,
    new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_,
    new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_,
    new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_,
    new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_,
    new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_,
    new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_,
    new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_,
    new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_,
    new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_,
    new_n7531_, new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_,
    new_n7537_, new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_,
    new_n7543_, new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_,
    new_n7549_, new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_,
    new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_,
    new_n7561_, new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_,
    new_n7567_, new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_,
    new_n7573_, new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_,
    new_n7579_, new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_,
    new_n7585_, new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_,
    new_n7591_, new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_,
    new_n7597_, new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_,
    new_n7603_, new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_,
    new_n7609_, new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_,
    new_n7615_, new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_,
    new_n7621_, new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_,
    new_n7627_, new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_,
    new_n7633_, new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_,
    new_n7639_, new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_,
    new_n7645_, new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_,
    new_n7651_, new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_,
    new_n7657_, new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_,
    new_n7663_, new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_,
    new_n7669_, new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_,
    new_n7675_, new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_,
    new_n7681_, new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_,
    new_n7687_, new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_,
    new_n7693_, new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_,
    new_n7699_, new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_,
    new_n7705_, new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_,
    new_n7711_, new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_,
    new_n7717_, new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_,
    new_n7723_, new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_,
    new_n7729_, new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_,
    new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_,
    new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_,
    new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_,
    new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7758_,
    new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_,
    new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7770_,
    new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_,
    new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_,
    new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_,
    new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_, new_n7794_,
    new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_, new_n7800_,
    new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_, new_n7806_,
    new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_, new_n7812_,
    new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_, new_n7818_,
    new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_,
    new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_,
    new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_,
    new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_,
    new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_, new_n7848_,
    new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_,
    new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_,
    new_n7861_, new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_,
    new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_,
    new_n7873_, new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_,
    new_n7879_, new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_,
    new_n7885_, new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_,
    new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_,
    new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_,
    new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_,
    new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_,
    new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_, new_n7920_,
    new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_,
    new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_,
    new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_,
    new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_,
    new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_, new_n7950_,
    new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_,
    new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_,
    new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_,
    new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_,
    new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_,
    new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_,
    new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_,
    new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_,
    new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_,
    new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_,
    new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_,
    new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_,
    new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_,
    new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_,
    new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_,
    new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_,
    new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_, new_n8052_,
    new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_,
    new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_,
    new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_, new_n8070_,
    new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_, new_n8076_,
    new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_,
    new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_,
    new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_,
    new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_,
    new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_,
    new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_,
    new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_,
    new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_,
    new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_,
    new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_,
    new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_,
    new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_,
    new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_,
    new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_,
    new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_,
    new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_,
    new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_,
    new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_,
    new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_,
    new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_,
    new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_,
    new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_,
    new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_,
    new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_,
    new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_,
    new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_,
    new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_,
    new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_,
    new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_,
    new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_,
    new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_,
    new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_,
    new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_,
    new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_,
    new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_,
    new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_,
    new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_,
    new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_,
    new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_,
    new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_,
    new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_,
    new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_,
    new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_,
    new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_,
    new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_,
    new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_,
    new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_,
    new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_,
    new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_,
    new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_,
    new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_,
    new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_,
    new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_,
    new_n8395_;
  assign new_n27_ = ~A302 & ~A301;
  assign new_n28_ = A300 & new_n27_;
  assign new_n29_ = ~A269 & ~A268;
  assign new_n30_ = new_n28_ & new_n29_;
  assign new_n31_ = ~A267 & ~A266;
  assign new_n32_ = A265 & ~A203;
  assign new_n33_ = new_n31_ & new_n32_;
  assign new_n34_ = new_n30_ & new_n33_;
  assign new_n35_ = ~A202 & ~A201;
  assign new_n36_ = ~A200 & new_n35_;
  assign new_n37_ = A199 & A166;
  assign new_n38_ = new_n36_ & new_n37_;
  assign new_n39_ = ~A167 & ~A168;
  assign new_n40_ = ~A169 & A170;
  assign new_n41_ = new_n39_ & new_n40_;
  assign new_n42_ = new_n38_ & new_n41_;
  assign new_n43_ = new_n34_ & new_n42_;
  assign new_n44_ = ~A267 & A266;
  assign new_n45_ = ~A265 & ~A203;
  assign new_n46_ = new_n44_ & new_n45_;
  assign new_n47_ = new_n30_ & new_n46_;
  assign new_n48_ = new_n42_ & new_n47_;
  assign new_n49_ = ~new_n43_ & ~new_n48_;
  assign new_n50_ = A200 & new_n35_;
  assign new_n51_ = ~A199 & A166;
  assign new_n52_ = new_n50_ & new_n51_;
  assign new_n53_ = new_n41_ & new_n52_;
  assign new_n54_ = new_n34_ & new_n53_;
  assign new_n55_ = new_n47_ & new_n53_;
  assign new_n56_ = ~new_n54_ & ~new_n55_;
  assign new_n57_ = new_n49_ & new_n56_;
  assign new_n58_ = A199 & ~A166;
  assign new_n59_ = new_n36_ & new_n58_;
  assign new_n60_ = A167 & ~A168;
  assign new_n61_ = new_n40_ & new_n60_;
  assign new_n62_ = new_n59_ & new_n61_;
  assign new_n63_ = new_n34_ & new_n62_;
  assign new_n64_ = new_n47_ & new_n62_;
  assign new_n65_ = ~new_n63_ & ~new_n64_;
  assign new_n66_ = ~A199 & ~A166;
  assign new_n67_ = new_n50_ & new_n66_;
  assign new_n68_ = new_n61_ & new_n67_;
  assign new_n69_ = new_n34_ & new_n68_;
  assign new_n70_ = new_n47_ & new_n68_;
  assign new_n71_ = ~new_n69_ & ~new_n70_;
  assign new_n72_ = new_n65_ & new_n71_;
  assign new_n73_ = new_n57_ & new_n72_;
  assign new_n74_ = ~A299 & ~A298;
  assign new_n75_ = ~A269 & new_n74_;
  assign new_n76_ = ~A268 & ~A267;
  assign new_n77_ = new_n75_ & new_n76_;
  assign new_n78_ = ~A266 & A265;
  assign new_n79_ = ~A203 & ~A202;
  assign new_n80_ = new_n78_ & new_n79_;
  assign new_n81_ = new_n77_ & new_n80_;
  assign new_n82_ = ~A201 & ~A200;
  assign new_n83_ = new_n37_ & new_n82_;
  assign new_n84_ = new_n41_ & new_n83_;
  assign new_n85_ = new_n81_ & new_n84_;
  assign new_n86_ = A299 & A298;
  assign new_n87_ = ~A269 & new_n86_;
  assign new_n88_ = new_n76_ & new_n87_;
  assign new_n89_ = new_n80_ & new_n88_;
  assign new_n90_ = new_n84_ & new_n89_;
  assign new_n91_ = ~new_n85_ & ~new_n90_;
  assign new_n92_ = A302 & ~A300;
  assign new_n93_ = ~A269 & new_n92_;
  assign new_n94_ = new_n76_ & new_n93_;
  assign new_n95_ = new_n80_ & new_n94_;
  assign new_n96_ = new_n84_ & new_n95_;
  assign new_n97_ = A301 & ~A300;
  assign new_n98_ = ~A269 & new_n97_;
  assign new_n99_ = new_n76_ & new_n98_;
  assign new_n100_ = new_n80_ & new_n99_;
  assign new_n101_ = new_n84_ & new_n100_;
  assign new_n102_ = ~new_n96_ & ~new_n101_;
  assign new_n103_ = new_n91_ & new_n102_;
  assign new_n104_ = A266 & ~A265;
  assign new_n105_ = new_n79_ & new_n104_;
  assign new_n106_ = new_n77_ & new_n105_;
  assign new_n107_ = new_n84_ & new_n106_;
  assign new_n108_ = A269 & A267;
  assign new_n109_ = new_n28_ & new_n108_;
  assign new_n110_ = new_n80_ & new_n109_;
  assign new_n111_ = new_n84_ & new_n110_;
  assign new_n112_ = A268 & A267;
  assign new_n113_ = new_n28_ & new_n112_;
  assign new_n114_ = new_n80_ & new_n113_;
  assign new_n115_ = new_n84_ & new_n114_;
  assign new_n116_ = ~new_n111_ & ~new_n115_;
  assign new_n117_ = ~new_n107_ & new_n116_;
  assign new_n118_ = new_n103_ & new_n117_;
  assign new_n119_ = new_n73_ & new_n118_;
  assign new_n120_ = new_n88_ & new_n105_;
  assign new_n121_ = new_n84_ & new_n120_;
  assign new_n122_ = new_n94_ & new_n105_;
  assign new_n123_ = new_n84_ & new_n122_;
  assign new_n124_ = ~new_n121_ & ~new_n123_;
  assign new_n125_ = new_n99_ & new_n105_;
  assign new_n126_ = new_n84_ & new_n125_;
  assign new_n127_ = new_n105_ & new_n109_;
  assign new_n128_ = new_n84_ & new_n127_;
  assign new_n129_ = ~new_n126_ & ~new_n128_;
  assign new_n130_ = new_n124_ & new_n129_;
  assign new_n131_ = ~A265 & A203;
  assign new_n132_ = new_n44_ & new_n131_;
  assign new_n133_ = new_n30_ & new_n132_;
  assign new_n134_ = A201 & ~A200;
  assign new_n135_ = new_n37_ & new_n134_;
  assign new_n136_ = new_n41_ & new_n135_;
  assign new_n137_ = new_n133_ & new_n136_;
  assign new_n138_ = new_n105_ & new_n113_;
  assign new_n139_ = new_n84_ & new_n138_;
  assign new_n140_ = A265 & A203;
  assign new_n141_ = new_n31_ & new_n140_;
  assign new_n142_ = new_n30_ & new_n141_;
  assign new_n143_ = new_n136_ & new_n142_;
  assign new_n144_ = ~new_n139_ & ~new_n143_;
  assign new_n145_ = ~new_n137_ & new_n144_;
  assign new_n146_ = new_n130_ & new_n145_;
  assign new_n147_ = A265 & A202;
  assign new_n148_ = new_n31_ & new_n147_;
  assign new_n149_ = new_n30_ & new_n148_;
  assign new_n150_ = new_n136_ & new_n149_;
  assign new_n151_ = ~A265 & A202;
  assign new_n152_ = new_n44_ & new_n151_;
  assign new_n153_ = new_n30_ & new_n152_;
  assign new_n154_ = new_n136_ & new_n153_;
  assign new_n155_ = ~new_n150_ & ~new_n154_;
  assign new_n156_ = ~A201 & A200;
  assign new_n157_ = new_n51_ & new_n156_;
  assign new_n158_ = new_n41_ & new_n157_;
  assign new_n159_ = new_n81_ & new_n158_;
  assign new_n160_ = new_n89_ & new_n158_;
  assign new_n161_ = ~new_n159_ & ~new_n160_;
  assign new_n162_ = new_n155_ & new_n161_;
  assign new_n163_ = new_n110_ & new_n158_;
  assign new_n164_ = new_n95_ & new_n158_;
  assign new_n165_ = new_n100_ & new_n158_;
  assign new_n166_ = ~new_n164_ & ~new_n165_;
  assign new_n167_ = ~new_n163_ & new_n166_;
  assign new_n168_ = new_n162_ & new_n167_;
  assign new_n169_ = new_n146_ & new_n168_;
  assign new_n170_ = new_n119_ & new_n169_;
  assign new_n171_ = new_n114_ & new_n158_;
  assign new_n172_ = new_n106_ & new_n158_;
  assign new_n173_ = ~new_n171_ & ~new_n172_;
  assign new_n174_ = new_n120_ & new_n158_;
  assign new_n175_ = new_n122_ & new_n158_;
  assign new_n176_ = ~new_n174_ & ~new_n175_;
  assign new_n177_ = new_n173_ & new_n176_;
  assign new_n178_ = new_n125_ & new_n158_;
  assign new_n179_ = new_n127_ & new_n158_;
  assign new_n180_ = ~new_n178_ & ~new_n179_;
  assign new_n181_ = new_n138_ & new_n158_;
  assign new_n182_ = A201 & A200;
  assign new_n183_ = new_n51_ & new_n182_;
  assign new_n184_ = new_n41_ & new_n183_;
  assign new_n185_ = new_n142_ & new_n184_;
  assign new_n186_ = ~new_n181_ & ~new_n185_;
  assign new_n187_ = new_n180_ & new_n186_;
  assign new_n188_ = new_n177_ & new_n187_;
  assign new_n189_ = new_n133_ & new_n184_;
  assign new_n190_ = new_n149_ & new_n184_;
  assign new_n191_ = ~new_n189_ & ~new_n190_;
  assign new_n192_ = new_n153_ & new_n184_;
  assign new_n193_ = new_n58_ & new_n82_;
  assign new_n194_ = new_n61_ & new_n193_;
  assign new_n195_ = new_n81_ & new_n194_;
  assign new_n196_ = ~new_n192_ & ~new_n195_;
  assign new_n197_ = new_n191_ & new_n196_;
  assign new_n198_ = new_n100_ & new_n194_;
  assign new_n199_ = new_n89_ & new_n194_;
  assign new_n200_ = new_n95_ & new_n194_;
  assign new_n201_ = ~new_n199_ & ~new_n200_;
  assign new_n202_ = ~new_n198_ & new_n201_;
  assign new_n203_ = new_n197_ & new_n202_;
  assign new_n204_ = new_n188_ & new_n203_;
  assign new_n205_ = new_n110_ & new_n194_;
  assign new_n206_ = new_n114_ & new_n194_;
  assign new_n207_ = ~new_n205_ & ~new_n206_;
  assign new_n208_ = new_n106_ & new_n194_;
  assign new_n209_ = new_n120_ & new_n194_;
  assign new_n210_ = ~new_n208_ & ~new_n209_;
  assign new_n211_ = new_n207_ & new_n210_;
  assign new_n212_ = new_n127_ & new_n194_;
  assign new_n213_ = new_n122_ & new_n194_;
  assign new_n214_ = new_n125_ & new_n194_;
  assign new_n215_ = ~new_n213_ & ~new_n214_;
  assign new_n216_ = ~new_n212_ & new_n215_;
  assign new_n217_ = new_n211_ & new_n216_;
  assign new_n218_ = new_n138_ & new_n194_;
  assign new_n219_ = new_n58_ & new_n134_;
  assign new_n220_ = new_n61_ & new_n219_;
  assign new_n221_ = new_n142_ & new_n220_;
  assign new_n222_ = ~new_n218_ & ~new_n221_;
  assign new_n223_ = new_n133_ & new_n220_;
  assign new_n224_ = new_n149_ & new_n220_;
  assign new_n225_ = ~new_n223_ & ~new_n224_;
  assign new_n226_ = new_n222_ & new_n225_;
  assign new_n227_ = new_n66_ & new_n156_;
  assign new_n228_ = new_n61_ & new_n227_;
  assign new_n229_ = new_n89_ & new_n228_;
  assign new_n230_ = new_n153_ & new_n220_;
  assign new_n231_ = new_n81_ & new_n228_;
  assign new_n232_ = ~new_n230_ & ~new_n231_;
  assign new_n233_ = ~new_n229_ & new_n232_;
  assign new_n234_ = new_n226_ & new_n233_;
  assign new_n235_ = new_n217_ & new_n234_;
  assign new_n236_ = new_n204_ & new_n235_;
  assign new_n237_ = new_n170_ & new_n236_;
  assign new_n238_ = new_n95_ & new_n228_;
  assign new_n239_ = new_n100_ & new_n228_;
  assign new_n240_ = ~new_n238_ & ~new_n239_;
  assign new_n241_ = new_n110_ & new_n228_;
  assign new_n242_ = new_n114_ & new_n228_;
  assign new_n243_ = ~new_n241_ & ~new_n242_;
  assign new_n244_ = new_n240_ & new_n243_;
  assign new_n245_ = new_n106_ & new_n228_;
  assign new_n246_ = new_n120_ & new_n228_;
  assign new_n247_ = ~new_n245_ & ~new_n246_;
  assign new_n248_ = new_n122_ & new_n228_;
  assign new_n249_ = new_n125_ & new_n228_;
  assign new_n250_ = ~new_n248_ & ~new_n249_;
  assign new_n251_ = new_n247_ & new_n250_;
  assign new_n252_ = new_n244_ & new_n251_;
  assign new_n253_ = new_n127_ & new_n228_;
  assign new_n254_ = new_n138_ & new_n228_;
  assign new_n255_ = ~new_n253_ & ~new_n254_;
  assign new_n256_ = new_n66_ & new_n182_;
  assign new_n257_ = new_n61_ & new_n256_;
  assign new_n258_ = new_n142_ & new_n257_;
  assign new_n259_ = new_n133_ & new_n257_;
  assign new_n260_ = ~new_n258_ & ~new_n259_;
  assign new_n261_ = new_n255_ & new_n260_;
  assign new_n262_ = ~A200 & A199;
  assign new_n263_ = new_n35_ & new_n262_;
  assign new_n264_ = A166 & ~A167;
  assign new_n265_ = A168 & A169;
  assign new_n266_ = new_n264_ & new_n265_;
  assign new_n267_ = new_n263_ & new_n266_;
  assign new_n268_ = new_n34_ & new_n267_;
  assign new_n269_ = new_n149_ & new_n257_;
  assign new_n270_ = new_n153_ & new_n257_;
  assign new_n271_ = ~new_n269_ & ~new_n270_;
  assign new_n272_ = ~new_n268_ & new_n271_;
  assign new_n273_ = new_n261_ & new_n272_;
  assign new_n274_ = new_n252_ & new_n273_;
  assign new_n275_ = new_n47_ & new_n267_;
  assign new_n276_ = A200 & ~A199;
  assign new_n277_ = new_n35_ & new_n276_;
  assign new_n278_ = new_n266_ & new_n277_;
  assign new_n279_ = new_n34_ & new_n278_;
  assign new_n280_ = ~new_n275_ & ~new_n279_;
  assign new_n281_ = new_n47_ & new_n278_;
  assign new_n282_ = ~A166 & A167;
  assign new_n283_ = new_n265_ & new_n282_;
  assign new_n284_ = new_n263_ & new_n283_;
  assign new_n285_ = new_n34_ & new_n284_;
  assign new_n286_ = ~new_n281_ & ~new_n285_;
  assign new_n287_ = new_n280_ & new_n286_;
  assign new_n288_ = new_n277_ & new_n283_;
  assign new_n289_ = new_n47_ & new_n288_;
  assign new_n290_ = new_n47_ & new_n284_;
  assign new_n291_ = new_n34_ & new_n288_;
  assign new_n292_ = ~new_n290_ & ~new_n291_;
  assign new_n293_ = ~new_n289_ & new_n292_;
  assign new_n294_ = new_n287_ & new_n293_;
  assign new_n295_ = A168 & ~A170;
  assign new_n296_ = new_n264_ & new_n295_;
  assign new_n297_ = new_n263_ & new_n296_;
  assign new_n298_ = new_n34_ & new_n297_;
  assign new_n299_ = new_n47_ & new_n297_;
  assign new_n300_ = ~new_n298_ & ~new_n299_;
  assign new_n301_ = new_n277_ & new_n296_;
  assign new_n302_ = new_n34_ & new_n301_;
  assign new_n303_ = new_n47_ & new_n301_;
  assign new_n304_ = ~new_n302_ & ~new_n303_;
  assign new_n305_ = new_n300_ & new_n304_;
  assign new_n306_ = new_n282_ & new_n295_;
  assign new_n307_ = new_n277_ & new_n306_;
  assign new_n308_ = new_n34_ & new_n307_;
  assign new_n309_ = new_n263_ & new_n306_;
  assign new_n310_ = new_n34_ & new_n309_;
  assign new_n311_ = new_n47_ & new_n309_;
  assign new_n312_ = ~new_n310_ & ~new_n311_;
  assign new_n313_ = ~new_n308_ & new_n312_;
  assign new_n314_ = new_n305_ & new_n313_;
  assign new_n315_ = new_n294_ & new_n314_;
  assign new_n316_ = new_n274_ & new_n315_;
  assign new_n317_ = new_n47_ & new_n307_;
  assign new_n318_ = new_n74_ & new_n108_;
  assign new_n319_ = new_n80_ & new_n318_;
  assign new_n320_ = new_n84_ & new_n319_;
  assign new_n321_ = ~new_n317_ & ~new_n320_;
  assign new_n322_ = new_n86_ & new_n108_;
  assign new_n323_ = new_n80_ & new_n322_;
  assign new_n324_ = new_n84_ & new_n323_;
  assign new_n325_ = new_n92_ & new_n108_;
  assign new_n326_ = new_n80_ & new_n325_;
  assign new_n327_ = new_n84_ & new_n326_;
  assign new_n328_ = ~new_n324_ & ~new_n327_;
  assign new_n329_ = new_n321_ & new_n328_;
  assign new_n330_ = new_n97_ & new_n108_;
  assign new_n331_ = new_n80_ & new_n330_;
  assign new_n332_ = new_n84_ & new_n331_;
  assign new_n333_ = new_n74_ & new_n112_;
  assign new_n334_ = new_n80_ & new_n333_;
  assign new_n335_ = new_n84_ & new_n334_;
  assign new_n336_ = ~new_n332_ & ~new_n335_;
  assign new_n337_ = new_n86_ & new_n112_;
  assign new_n338_ = new_n80_ & new_n337_;
  assign new_n339_ = new_n84_ & new_n338_;
  assign new_n340_ = new_n92_ & new_n112_;
  assign new_n341_ = new_n80_ & new_n340_;
  assign new_n342_ = new_n84_ & new_n341_;
  assign new_n343_ = ~new_n339_ & ~new_n342_;
  assign new_n344_ = new_n336_ & new_n343_;
  assign new_n345_ = new_n329_ & new_n344_;
  assign new_n346_ = new_n97_ & new_n112_;
  assign new_n347_ = new_n80_ & new_n346_;
  assign new_n348_ = new_n84_ & new_n347_;
  assign new_n349_ = new_n105_ & new_n318_;
  assign new_n350_ = new_n84_ & new_n349_;
  assign new_n351_ = ~new_n348_ & ~new_n350_;
  assign new_n352_ = new_n105_ & new_n322_;
  assign new_n353_ = new_n84_ & new_n352_;
  assign new_n354_ = new_n105_ & new_n325_;
  assign new_n355_ = new_n84_ & new_n354_;
  assign new_n356_ = ~new_n353_ & ~new_n355_;
  assign new_n357_ = new_n351_ & new_n356_;
  assign new_n358_ = new_n105_ & new_n337_;
  assign new_n359_ = new_n84_ & new_n358_;
  assign new_n360_ = new_n105_ & new_n330_;
  assign new_n361_ = new_n84_ & new_n360_;
  assign new_n362_ = new_n105_ & new_n333_;
  assign new_n363_ = new_n84_ & new_n362_;
  assign new_n364_ = ~new_n361_ & ~new_n363_;
  assign new_n365_ = ~new_n359_ & new_n364_;
  assign new_n366_ = new_n357_ & new_n365_;
  assign new_n367_ = new_n345_ & new_n366_;
  assign new_n368_ = new_n105_ & new_n340_;
  assign new_n369_ = new_n84_ & new_n368_;
  assign new_n370_ = new_n105_ & new_n346_;
  assign new_n371_ = new_n84_ & new_n370_;
  assign new_n372_ = ~new_n369_ & ~new_n371_;
  assign new_n373_ = new_n29_ & new_n74_;
  assign new_n374_ = new_n141_ & new_n373_;
  assign new_n375_ = new_n136_ & new_n374_;
  assign new_n376_ = new_n29_ & new_n86_;
  assign new_n377_ = new_n141_ & new_n376_;
  assign new_n378_ = new_n136_ & new_n377_;
  assign new_n379_ = ~new_n375_ & ~new_n378_;
  assign new_n380_ = new_n372_ & new_n379_;
  assign new_n381_ = A300 & A269;
  assign new_n382_ = new_n27_ & new_n381_;
  assign new_n383_ = A267 & ~A266;
  assign new_n384_ = new_n140_ & new_n383_;
  assign new_n385_ = new_n382_ & new_n384_;
  assign new_n386_ = new_n136_ & new_n385_;
  assign new_n387_ = new_n29_ & new_n92_;
  assign new_n388_ = new_n141_ & new_n387_;
  assign new_n389_ = new_n136_ & new_n388_;
  assign new_n390_ = new_n29_ & new_n97_;
  assign new_n391_ = new_n141_ & new_n390_;
  assign new_n392_ = new_n136_ & new_n391_;
  assign new_n393_ = ~new_n389_ & ~new_n392_;
  assign new_n394_ = ~new_n386_ & new_n393_;
  assign new_n395_ = new_n380_ & new_n394_;
  assign new_n396_ = A300 & A268;
  assign new_n397_ = new_n27_ & new_n396_;
  assign new_n398_ = new_n384_ & new_n397_;
  assign new_n399_ = new_n136_ & new_n398_;
  assign new_n400_ = new_n132_ & new_n373_;
  assign new_n401_ = new_n136_ & new_n400_;
  assign new_n402_ = ~new_n399_ & ~new_n401_;
  assign new_n403_ = new_n132_ & new_n376_;
  assign new_n404_ = new_n136_ & new_n403_;
  assign new_n405_ = new_n132_ & new_n387_;
  assign new_n406_ = new_n136_ & new_n405_;
  assign new_n407_ = ~new_n404_ & ~new_n406_;
  assign new_n408_ = new_n402_ & new_n407_;
  assign new_n409_ = A267 & A266;
  assign new_n410_ = new_n131_ & new_n409_;
  assign new_n411_ = new_n397_ & new_n410_;
  assign new_n412_ = new_n136_ & new_n411_;
  assign new_n413_ = new_n132_ & new_n390_;
  assign new_n414_ = new_n136_ & new_n413_;
  assign new_n415_ = new_n382_ & new_n410_;
  assign new_n416_ = new_n136_ & new_n415_;
  assign new_n417_ = ~new_n414_ & ~new_n416_;
  assign new_n418_ = ~new_n412_ & new_n417_;
  assign new_n419_ = new_n408_ & new_n418_;
  assign new_n420_ = new_n395_ & new_n419_;
  assign new_n421_ = new_n367_ & new_n420_;
  assign new_n422_ = new_n316_ & new_n421_;
  assign new_n423_ = new_n237_ & new_n422_;
  assign new_n424_ = new_n148_ & new_n373_;
  assign new_n425_ = new_n136_ & new_n424_;
  assign new_n426_ = new_n148_ & new_n376_;
  assign new_n427_ = new_n136_ & new_n426_;
  assign new_n428_ = ~new_n425_ & ~new_n427_;
  assign new_n429_ = new_n148_ & new_n387_;
  assign new_n430_ = new_n136_ & new_n429_;
  assign new_n431_ = new_n148_ & new_n390_;
  assign new_n432_ = new_n136_ & new_n431_;
  assign new_n433_ = ~new_n430_ & ~new_n432_;
  assign new_n434_ = new_n428_ & new_n433_;
  assign new_n435_ = new_n147_ & new_n383_;
  assign new_n436_ = new_n382_ & new_n435_;
  assign new_n437_ = new_n136_ & new_n436_;
  assign new_n438_ = new_n397_ & new_n435_;
  assign new_n439_ = new_n136_ & new_n438_;
  assign new_n440_ = ~new_n437_ & ~new_n439_;
  assign new_n441_ = new_n152_ & new_n373_;
  assign new_n442_ = new_n136_ & new_n441_;
  assign new_n443_ = new_n152_ & new_n376_;
  assign new_n444_ = new_n136_ & new_n443_;
  assign new_n445_ = ~new_n442_ & ~new_n444_;
  assign new_n446_ = new_n440_ & new_n445_;
  assign new_n447_ = new_n434_ & new_n446_;
  assign new_n448_ = new_n152_ & new_n387_;
  assign new_n449_ = new_n136_ & new_n448_;
  assign new_n450_ = new_n152_ & new_n390_;
  assign new_n451_ = new_n136_ & new_n450_;
  assign new_n452_ = ~new_n449_ & ~new_n451_;
  assign new_n453_ = new_n151_ & new_n409_;
  assign new_n454_ = new_n382_ & new_n453_;
  assign new_n455_ = new_n136_ & new_n454_;
  assign new_n456_ = new_n397_ & new_n453_;
  assign new_n457_ = new_n136_ & new_n456_;
  assign new_n458_ = ~new_n455_ & ~new_n457_;
  assign new_n459_ = new_n452_ & new_n458_;
  assign new_n460_ = new_n158_ & new_n326_;
  assign new_n461_ = new_n158_ & new_n319_;
  assign new_n462_ = new_n158_ & new_n323_;
  assign new_n463_ = ~new_n461_ & ~new_n462_;
  assign new_n464_ = ~new_n460_ & new_n463_;
  assign new_n465_ = new_n459_ & new_n464_;
  assign new_n466_ = new_n447_ & new_n465_;
  assign new_n467_ = new_n158_ & new_n331_;
  assign new_n468_ = new_n158_ & new_n334_;
  assign new_n469_ = ~new_n467_ & ~new_n468_;
  assign new_n470_ = new_n158_ & new_n338_;
  assign new_n471_ = new_n158_ & new_n341_;
  assign new_n472_ = ~new_n470_ & ~new_n471_;
  assign new_n473_ = new_n469_ & new_n472_;
  assign new_n474_ = new_n158_ & new_n352_;
  assign new_n475_ = new_n158_ & new_n347_;
  assign new_n476_ = new_n158_ & new_n349_;
  assign new_n477_ = ~new_n475_ & ~new_n476_;
  assign new_n478_ = ~new_n474_ & new_n477_;
  assign new_n479_ = new_n473_ & new_n478_;
  assign new_n480_ = new_n158_ & new_n354_;
  assign new_n481_ = new_n158_ & new_n360_;
  assign new_n482_ = ~new_n480_ & ~new_n481_;
  assign new_n483_ = new_n158_ & new_n362_;
  assign new_n484_ = new_n158_ & new_n358_;
  assign new_n485_ = ~new_n483_ & ~new_n484_;
  assign new_n486_ = new_n482_ & new_n485_;
  assign new_n487_ = new_n184_ & new_n374_;
  assign new_n488_ = new_n158_ & new_n368_;
  assign new_n489_ = new_n158_ & new_n370_;
  assign new_n490_ = ~new_n488_ & ~new_n489_;
  assign new_n491_ = ~new_n487_ & new_n490_;
  assign new_n492_ = new_n486_ & new_n491_;
  assign new_n493_ = new_n479_ & new_n492_;
  assign new_n494_ = new_n466_ & new_n493_;
  assign new_n495_ = new_n184_ & new_n377_;
  assign new_n496_ = new_n184_ & new_n388_;
  assign new_n497_ = ~new_n495_ & ~new_n496_;
  assign new_n498_ = new_n184_ & new_n391_;
  assign new_n499_ = new_n184_ & new_n385_;
  assign new_n500_ = ~new_n498_ & ~new_n499_;
  assign new_n501_ = new_n497_ & new_n500_;
  assign new_n502_ = new_n184_ & new_n398_;
  assign new_n503_ = new_n184_ & new_n400_;
  assign new_n504_ = ~new_n502_ & ~new_n503_;
  assign new_n505_ = new_n184_ & new_n403_;
  assign new_n506_ = new_n184_ & new_n405_;
  assign new_n507_ = ~new_n505_ & ~new_n506_;
  assign new_n508_ = new_n504_ & new_n507_;
  assign new_n509_ = new_n501_ & new_n508_;
  assign new_n510_ = new_n184_ & new_n413_;
  assign new_n511_ = new_n184_ & new_n415_;
  assign new_n512_ = ~new_n510_ & ~new_n511_;
  assign new_n513_ = new_n184_ & new_n411_;
  assign new_n514_ = new_n184_ & new_n424_;
  assign new_n515_ = ~new_n513_ & ~new_n514_;
  assign new_n516_ = new_n512_ & new_n515_;
  assign new_n517_ = new_n184_ & new_n431_;
  assign new_n518_ = new_n184_ & new_n426_;
  assign new_n519_ = new_n184_ & new_n429_;
  assign new_n520_ = ~new_n518_ & ~new_n519_;
  assign new_n521_ = ~new_n517_ & new_n520_;
  assign new_n522_ = new_n516_ & new_n521_;
  assign new_n523_ = new_n509_ & new_n522_;
  assign new_n524_ = new_n184_ & new_n436_;
  assign new_n525_ = new_n184_ & new_n438_;
  assign new_n526_ = ~new_n524_ & ~new_n525_;
  assign new_n527_ = new_n184_ & new_n441_;
  assign new_n528_ = new_n184_ & new_n443_;
  assign new_n529_ = ~new_n527_ & ~new_n528_;
  assign new_n530_ = new_n526_ & new_n529_;
  assign new_n531_ = new_n184_ & new_n454_;
  assign new_n532_ = new_n184_ & new_n448_;
  assign new_n533_ = new_n184_ & new_n450_;
  assign new_n534_ = ~new_n532_ & ~new_n533_;
  assign new_n535_ = ~new_n531_ & new_n534_;
  assign new_n536_ = new_n530_ & new_n535_;
  assign new_n537_ = new_n184_ & new_n456_;
  assign new_n538_ = ~A300 & A299;
  assign new_n539_ = new_n27_ & new_n538_;
  assign new_n540_ = ~A298 & ~A269;
  assign new_n541_ = ~A268 & A267;
  assign new_n542_ = new_n540_ & new_n541_;
  assign new_n543_ = new_n539_ & new_n542_;
  assign new_n544_ = A201 & A166;
  assign new_n545_ = new_n79_ & new_n544_;
  assign new_n546_ = new_n41_ & new_n545_;
  assign new_n547_ = new_n543_ & new_n546_;
  assign new_n548_ = ~new_n537_ & ~new_n547_;
  assign new_n549_ = ~A300 & ~A299;
  assign new_n550_ = new_n27_ & new_n549_;
  assign new_n551_ = A298 & ~A269;
  assign new_n552_ = new_n541_ & new_n551_;
  assign new_n553_ = new_n550_ & new_n552_;
  assign new_n554_ = new_n546_ & new_n553_;
  assign new_n555_ = new_n194_ & new_n319_;
  assign new_n556_ = ~new_n554_ & ~new_n555_;
  assign new_n557_ = new_n548_ & new_n556_;
  assign new_n558_ = new_n194_ & new_n331_;
  assign new_n559_ = new_n194_ & new_n323_;
  assign new_n560_ = new_n194_ & new_n326_;
  assign new_n561_ = ~new_n559_ & ~new_n560_;
  assign new_n562_ = ~new_n558_ & new_n561_;
  assign new_n563_ = new_n557_ & new_n562_;
  assign new_n564_ = new_n536_ & new_n563_;
  assign new_n565_ = new_n523_ & new_n564_;
  assign new_n566_ = new_n494_ & new_n565_;
  assign new_n567_ = new_n194_ & new_n334_;
  assign new_n568_ = new_n194_ & new_n338_;
  assign new_n569_ = ~new_n567_ & ~new_n568_;
  assign new_n570_ = new_n194_ & new_n341_;
  assign new_n571_ = new_n194_ & new_n347_;
  assign new_n572_ = ~new_n570_ & ~new_n571_;
  assign new_n573_ = new_n569_ & new_n572_;
  assign new_n574_ = new_n194_ & new_n349_;
  assign new_n575_ = new_n194_ & new_n352_;
  assign new_n576_ = ~new_n574_ & ~new_n575_;
  assign new_n577_ = new_n194_ & new_n354_;
  assign new_n578_ = new_n194_ & new_n360_;
  assign new_n579_ = ~new_n577_ & ~new_n578_;
  assign new_n580_ = new_n576_ & new_n579_;
  assign new_n581_ = new_n573_ & new_n580_;
  assign new_n582_ = new_n194_ & new_n362_;
  assign new_n583_ = new_n194_ & new_n358_;
  assign new_n584_ = ~new_n582_ & ~new_n583_;
  assign new_n585_ = new_n194_ & new_n368_;
  assign new_n586_ = new_n194_ & new_n370_;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = new_n584_ & new_n587_;
  assign new_n589_ = new_n220_ & new_n388_;
  assign new_n590_ = new_n220_ & new_n374_;
  assign new_n591_ = new_n220_ & new_n377_;
  assign new_n592_ = ~new_n590_ & ~new_n591_;
  assign new_n593_ = ~new_n589_ & new_n592_;
  assign new_n594_ = new_n588_ & new_n593_;
  assign new_n595_ = new_n581_ & new_n594_;
  assign new_n596_ = new_n220_ & new_n391_;
  assign new_n597_ = new_n220_ & new_n385_;
  assign new_n598_ = ~new_n596_ & ~new_n597_;
  assign new_n599_ = new_n220_ & new_n398_;
  assign new_n600_ = new_n220_ & new_n400_;
  assign new_n601_ = ~new_n599_ & ~new_n600_;
  assign new_n602_ = new_n598_ & new_n601_;
  assign new_n603_ = new_n220_ & new_n413_;
  assign new_n604_ = new_n220_ & new_n403_;
  assign new_n605_ = new_n220_ & new_n405_;
  assign new_n606_ = ~new_n604_ & ~new_n605_;
  assign new_n607_ = ~new_n603_ & new_n606_;
  assign new_n608_ = new_n602_ & new_n607_;
  assign new_n609_ = new_n220_ & new_n415_;
  assign new_n610_ = new_n220_ & new_n411_;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign new_n612_ = new_n220_ & new_n424_;
  assign new_n613_ = new_n220_ & new_n426_;
  assign new_n614_ = ~new_n612_ & ~new_n613_;
  assign new_n615_ = new_n611_ & new_n614_;
  assign new_n616_ = new_n220_ & new_n436_;
  assign new_n617_ = new_n220_ & new_n429_;
  assign new_n618_ = new_n220_ & new_n431_;
  assign new_n619_ = ~new_n617_ & ~new_n618_;
  assign new_n620_ = ~new_n616_ & new_n619_;
  assign new_n621_ = new_n615_ & new_n620_;
  assign new_n622_ = new_n608_ & new_n621_;
  assign new_n623_ = new_n595_ & new_n622_;
  assign new_n624_ = new_n220_ & new_n438_;
  assign new_n625_ = new_n220_ & new_n441_;
  assign new_n626_ = ~new_n624_ & ~new_n625_;
  assign new_n627_ = new_n220_ & new_n443_;
  assign new_n628_ = new_n220_ & new_n448_;
  assign new_n629_ = ~new_n627_ & ~new_n628_;
  assign new_n630_ = new_n626_ & new_n629_;
  assign new_n631_ = new_n220_ & new_n450_;
  assign new_n632_ = new_n220_ & new_n454_;
  assign new_n633_ = ~new_n631_ & ~new_n632_;
  assign new_n634_ = new_n220_ & new_n456_;
  assign new_n635_ = new_n228_ & new_n319_;
  assign new_n636_ = ~new_n634_ & ~new_n635_;
  assign new_n637_ = new_n633_ & new_n636_;
  assign new_n638_ = new_n630_ & new_n637_;
  assign new_n639_ = new_n228_ & new_n323_;
  assign new_n640_ = new_n228_ & new_n326_;
  assign new_n641_ = ~new_n639_ & ~new_n640_;
  assign new_n642_ = new_n228_ & new_n331_;
  assign new_n643_ = new_n228_ & new_n334_;
  assign new_n644_ = ~new_n642_ & ~new_n643_;
  assign new_n645_ = new_n641_ & new_n644_;
  assign new_n646_ = new_n228_ & new_n347_;
  assign new_n647_ = new_n228_ & new_n338_;
  assign new_n648_ = new_n228_ & new_n341_;
  assign new_n649_ = ~new_n647_ & ~new_n648_;
  assign new_n650_ = ~new_n646_ & new_n649_;
  assign new_n651_ = new_n645_ & new_n650_;
  assign new_n652_ = new_n638_ & new_n651_;
  assign new_n653_ = new_n228_ & new_n349_;
  assign new_n654_ = new_n228_ & new_n352_;
  assign new_n655_ = ~new_n653_ & ~new_n654_;
  assign new_n656_ = new_n228_ & new_n354_;
  assign new_n657_ = new_n228_ & new_n360_;
  assign new_n658_ = ~new_n656_ & ~new_n657_;
  assign new_n659_ = new_n655_ & new_n658_;
  assign new_n660_ = new_n228_ & new_n368_;
  assign new_n661_ = new_n228_ & new_n362_;
  assign new_n662_ = new_n228_ & new_n358_;
  assign new_n663_ = ~new_n661_ & ~new_n662_;
  assign new_n664_ = ~new_n660_ & new_n663_;
  assign new_n665_ = new_n659_ & new_n664_;
  assign new_n666_ = new_n228_ & new_n370_;
  assign new_n667_ = new_n257_ & new_n374_;
  assign new_n668_ = ~new_n666_ & ~new_n667_;
  assign new_n669_ = new_n257_ & new_n377_;
  assign new_n670_ = new_n257_ & new_n388_;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign new_n672_ = new_n668_ & new_n671_;
  assign new_n673_ = new_n257_ & new_n398_;
  assign new_n674_ = new_n257_ & new_n391_;
  assign new_n675_ = new_n257_ & new_n385_;
  assign new_n676_ = ~new_n674_ & ~new_n675_;
  assign new_n677_ = ~new_n673_ & new_n676_;
  assign new_n678_ = new_n672_ & new_n677_;
  assign new_n679_ = new_n665_ & new_n678_;
  assign new_n680_ = new_n652_ & new_n679_;
  assign new_n681_ = new_n623_ & new_n680_;
  assign new_n682_ = new_n566_ & new_n681_;
  assign new_n683_ = new_n423_ & new_n682_;
  assign new_n684_ = new_n257_ & new_n400_;
  assign new_n685_ = new_n257_ & new_n403_;
  assign new_n686_ = ~new_n684_ & ~new_n685_;
  assign new_n687_ = new_n257_ & new_n405_;
  assign new_n688_ = new_n257_ & new_n413_;
  assign new_n689_ = ~new_n687_ & ~new_n688_;
  assign new_n690_ = new_n686_ & new_n689_;
  assign new_n691_ = new_n257_ & new_n415_;
  assign new_n692_ = new_n257_ & new_n411_;
  assign new_n693_ = ~new_n691_ & ~new_n692_;
  assign new_n694_ = new_n257_ & new_n424_;
  assign new_n695_ = new_n257_ & new_n426_;
  assign new_n696_ = ~new_n694_ & ~new_n695_;
  assign new_n697_ = new_n693_ & new_n696_;
  assign new_n698_ = new_n690_ & new_n697_;
  assign new_n699_ = new_n257_ & new_n429_;
  assign new_n700_ = new_n257_ & new_n431_;
  assign new_n701_ = ~new_n699_ & ~new_n700_;
  assign new_n702_ = new_n257_ & new_n436_;
  assign new_n703_ = new_n257_ & new_n438_;
  assign new_n704_ = ~new_n702_ & ~new_n703_;
  assign new_n705_ = new_n701_ & new_n704_;
  assign new_n706_ = new_n257_ & new_n448_;
  assign new_n707_ = new_n257_ & new_n441_;
  assign new_n708_ = new_n257_ & new_n443_;
  assign new_n709_ = ~new_n707_ & ~new_n708_;
  assign new_n710_ = ~new_n706_ & new_n709_;
  assign new_n711_ = new_n705_ & new_n710_;
  assign new_n712_ = new_n698_ & new_n711_;
  assign new_n713_ = new_n257_ & new_n450_;
  assign new_n714_ = new_n257_ & new_n454_;
  assign new_n715_ = ~new_n713_ & ~new_n714_;
  assign new_n716_ = new_n257_ & new_n456_;
  assign new_n717_ = A201 & ~A166;
  assign new_n718_ = new_n79_ & new_n717_;
  assign new_n719_ = new_n61_ & new_n718_;
  assign new_n720_ = new_n543_ & new_n719_;
  assign new_n721_ = ~new_n716_ & ~new_n720_;
  assign new_n722_ = new_n715_ & new_n721_;
  assign new_n723_ = new_n79_ & new_n82_;
  assign new_n724_ = A199 & A168;
  assign new_n725_ = new_n40_ & new_n724_;
  assign new_n726_ = new_n723_ & new_n725_;
  assign new_n727_ = new_n553_ & new_n726_;
  assign new_n728_ = new_n553_ & new_n719_;
  assign new_n729_ = new_n543_ & new_n726_;
  assign new_n730_ = ~new_n728_ & ~new_n729_;
  assign new_n731_ = ~new_n727_ & new_n730_;
  assign new_n732_ = new_n722_ & new_n731_;
  assign new_n733_ = new_n79_ & new_n156_;
  assign new_n734_ = ~A199 & A168;
  assign new_n735_ = new_n40_ & new_n734_;
  assign new_n736_ = new_n733_ & new_n735_;
  assign new_n737_ = new_n543_ & new_n736_;
  assign new_n738_ = new_n553_ & new_n736_;
  assign new_n739_ = ~new_n737_ & ~new_n738_;
  assign new_n740_ = new_n33_ & new_n373_;
  assign new_n741_ = new_n267_ & new_n740_;
  assign new_n742_ = new_n33_ & new_n376_;
  assign new_n743_ = new_n267_ & new_n742_;
  assign new_n744_ = ~new_n741_ & ~new_n743_;
  assign new_n745_ = new_n739_ & new_n744_;
  assign new_n746_ = new_n32_ & new_n383_;
  assign new_n747_ = new_n382_ & new_n746_;
  assign new_n748_ = new_n267_ & new_n747_;
  assign new_n749_ = new_n33_ & new_n387_;
  assign new_n750_ = new_n267_ & new_n749_;
  assign new_n751_ = new_n33_ & new_n390_;
  assign new_n752_ = new_n267_ & new_n751_;
  assign new_n753_ = ~new_n750_ & ~new_n752_;
  assign new_n754_ = ~new_n748_ & new_n753_;
  assign new_n755_ = new_n745_ & new_n754_;
  assign new_n756_ = new_n732_ & new_n755_;
  assign new_n757_ = new_n712_ & new_n756_;
  assign new_n758_ = new_n397_ & new_n746_;
  assign new_n759_ = new_n267_ & new_n758_;
  assign new_n760_ = new_n46_ & new_n373_;
  assign new_n761_ = new_n267_ & new_n760_;
  assign new_n762_ = ~new_n759_ & ~new_n761_;
  assign new_n763_ = new_n46_ & new_n376_;
  assign new_n764_ = new_n267_ & new_n763_;
  assign new_n765_ = new_n46_ & new_n387_;
  assign new_n766_ = new_n267_ & new_n765_;
  assign new_n767_ = ~new_n764_ & ~new_n766_;
  assign new_n768_ = new_n762_ & new_n767_;
  assign new_n769_ = new_n46_ & new_n390_;
  assign new_n770_ = new_n267_ & new_n769_;
  assign new_n771_ = new_n45_ & new_n409_;
  assign new_n772_ = new_n382_ & new_n771_;
  assign new_n773_ = new_n267_ & new_n772_;
  assign new_n774_ = ~new_n770_ & ~new_n773_;
  assign new_n775_ = new_n397_ & new_n771_;
  assign new_n776_ = new_n267_ & new_n775_;
  assign new_n777_ = A300 & ~A269;
  assign new_n778_ = new_n27_ & new_n777_;
  assign new_n779_ = new_n76_ & new_n78_;
  assign new_n780_ = new_n778_ & new_n779_;
  assign new_n781_ = A203 & A201;
  assign new_n782_ = new_n262_ & new_n781_;
  assign new_n783_ = new_n266_ & new_n782_;
  assign new_n784_ = new_n780_ & new_n783_;
  assign new_n785_ = ~new_n776_ & ~new_n784_;
  assign new_n786_ = new_n774_ & new_n785_;
  assign new_n787_ = new_n768_ & new_n786_;
  assign new_n788_ = new_n76_ & new_n104_;
  assign new_n789_ = new_n778_ & new_n788_;
  assign new_n790_ = new_n783_ & new_n789_;
  assign new_n791_ = A202 & A201;
  assign new_n792_ = new_n262_ & new_n791_;
  assign new_n793_ = new_n266_ & new_n792_;
  assign new_n794_ = new_n780_ & new_n793_;
  assign new_n795_ = ~new_n790_ & ~new_n794_;
  assign new_n796_ = new_n789_ & new_n793_;
  assign new_n797_ = new_n278_ & new_n740_;
  assign new_n798_ = ~new_n796_ & ~new_n797_;
  assign new_n799_ = new_n795_ & new_n798_;
  assign new_n800_ = new_n278_ & new_n751_;
  assign new_n801_ = new_n278_ & new_n742_;
  assign new_n802_ = new_n278_ & new_n749_;
  assign new_n803_ = ~new_n801_ & ~new_n802_;
  assign new_n804_ = ~new_n800_ & new_n803_;
  assign new_n805_ = new_n799_ & new_n804_;
  assign new_n806_ = new_n787_ & new_n805_;
  assign new_n807_ = new_n278_ & new_n747_;
  assign new_n808_ = new_n278_ & new_n758_;
  assign new_n809_ = ~new_n807_ & ~new_n808_;
  assign new_n810_ = new_n278_ & new_n760_;
  assign new_n811_ = new_n278_ & new_n763_;
  assign new_n812_ = ~new_n810_ & ~new_n811_;
  assign new_n813_ = new_n809_ & new_n812_;
  assign new_n814_ = new_n278_ & new_n772_;
  assign new_n815_ = new_n278_ & new_n765_;
  assign new_n816_ = new_n278_ & new_n769_;
  assign new_n817_ = ~new_n815_ & ~new_n816_;
  assign new_n818_ = ~new_n814_ & new_n817_;
  assign new_n819_ = new_n813_ & new_n818_;
  assign new_n820_ = new_n278_ & new_n775_;
  assign new_n821_ = new_n276_ & new_n781_;
  assign new_n822_ = new_n266_ & new_n821_;
  assign new_n823_ = new_n780_ & new_n822_;
  assign new_n824_ = ~new_n820_ & ~new_n823_;
  assign new_n825_ = new_n789_ & new_n822_;
  assign new_n826_ = new_n276_ & new_n791_;
  assign new_n827_ = new_n266_ & new_n826_;
  assign new_n828_ = new_n780_ & new_n827_;
  assign new_n829_ = ~new_n825_ & ~new_n828_;
  assign new_n830_ = new_n824_ & new_n829_;
  assign new_n831_ = new_n284_ & new_n742_;
  assign new_n832_ = new_n789_ & new_n827_;
  assign new_n833_ = new_n284_ & new_n740_;
  assign new_n834_ = ~new_n832_ & ~new_n833_;
  assign new_n835_ = ~new_n831_ & new_n834_;
  assign new_n836_ = new_n830_ & new_n835_;
  assign new_n837_ = new_n819_ & new_n836_;
  assign new_n838_ = new_n806_ & new_n837_;
  assign new_n839_ = new_n757_ & new_n838_;
  assign new_n840_ = new_n284_ & new_n749_;
  assign new_n841_ = new_n284_ & new_n751_;
  assign new_n842_ = ~new_n840_ & ~new_n841_;
  assign new_n843_ = new_n284_ & new_n747_;
  assign new_n844_ = new_n284_ & new_n758_;
  assign new_n845_ = ~new_n843_ & ~new_n844_;
  assign new_n846_ = new_n842_ & new_n845_;
  assign new_n847_ = new_n284_ & new_n760_;
  assign new_n848_ = new_n284_ & new_n763_;
  assign new_n849_ = ~new_n847_ & ~new_n848_;
  assign new_n850_ = new_n284_ & new_n765_;
  assign new_n851_ = new_n284_ & new_n769_;
  assign new_n852_ = ~new_n850_ & ~new_n851_;
  assign new_n853_ = new_n849_ & new_n852_;
  assign new_n854_ = new_n846_ & new_n853_;
  assign new_n855_ = new_n284_ & new_n772_;
  assign new_n856_ = new_n284_ & new_n775_;
  assign new_n857_ = ~new_n855_ & ~new_n856_;
  assign new_n858_ = new_n283_ & new_n782_;
  assign new_n859_ = new_n780_ & new_n858_;
  assign new_n860_ = new_n789_ & new_n858_;
  assign new_n861_ = ~new_n859_ & ~new_n860_;
  assign new_n862_ = new_n857_ & new_n861_;
  assign new_n863_ = new_n288_ & new_n740_;
  assign new_n864_ = new_n283_ & new_n792_;
  assign new_n865_ = new_n780_ & new_n864_;
  assign new_n866_ = new_n789_ & new_n864_;
  assign new_n867_ = ~new_n865_ & ~new_n866_;
  assign new_n868_ = ~new_n863_ & new_n867_;
  assign new_n869_ = new_n862_ & new_n868_;
  assign new_n870_ = new_n854_ & new_n869_;
  assign new_n871_ = new_n288_ & new_n742_;
  assign new_n872_ = new_n288_ & new_n749_;
  assign new_n873_ = ~new_n871_ & ~new_n872_;
  assign new_n874_ = new_n288_ & new_n751_;
  assign new_n875_ = new_n288_ & new_n747_;
  assign new_n876_ = ~new_n874_ & ~new_n875_;
  assign new_n877_ = new_n873_ & new_n876_;
  assign new_n878_ = new_n288_ & new_n763_;
  assign new_n879_ = new_n288_ & new_n758_;
  assign new_n880_ = new_n288_ & new_n760_;
  assign new_n881_ = ~new_n879_ & ~new_n880_;
  assign new_n882_ = ~new_n878_ & new_n881_;
  assign new_n883_ = new_n877_ & new_n882_;
  assign new_n884_ = new_n288_ & new_n765_;
  assign new_n885_ = new_n288_ & new_n769_;
  assign new_n886_ = ~new_n884_ & ~new_n885_;
  assign new_n887_ = new_n288_ & new_n772_;
  assign new_n888_ = new_n288_ & new_n775_;
  assign new_n889_ = ~new_n887_ & ~new_n888_;
  assign new_n890_ = new_n886_ & new_n889_;
  assign new_n891_ = new_n283_ & new_n826_;
  assign new_n892_ = new_n780_ & new_n891_;
  assign new_n893_ = new_n283_ & new_n821_;
  assign new_n894_ = new_n780_ & new_n893_;
  assign new_n895_ = new_n789_ & new_n893_;
  assign new_n896_ = ~new_n894_ & ~new_n895_;
  assign new_n897_ = ~new_n892_ & new_n896_;
  assign new_n898_ = new_n890_ & new_n897_;
  assign new_n899_ = new_n883_ & new_n898_;
  assign new_n900_ = new_n870_ & new_n899_;
  assign new_n901_ = new_n789_ & new_n891_;
  assign new_n902_ = new_n297_ & new_n740_;
  assign new_n903_ = ~new_n901_ & ~new_n902_;
  assign new_n904_ = new_n297_ & new_n742_;
  assign new_n905_ = new_n297_ & new_n749_;
  assign new_n906_ = ~new_n904_ & ~new_n905_;
  assign new_n907_ = new_n903_ & new_n906_;
  assign new_n908_ = new_n297_ & new_n751_;
  assign new_n909_ = new_n297_ & new_n747_;
  assign new_n910_ = ~new_n908_ & ~new_n909_;
  assign new_n911_ = new_n297_ & new_n758_;
  assign new_n912_ = new_n297_ & new_n760_;
  assign new_n913_ = ~new_n911_ & ~new_n912_;
  assign new_n914_ = new_n910_ & new_n913_;
  assign new_n915_ = new_n907_ & new_n914_;
  assign new_n916_ = new_n297_ & new_n763_;
  assign new_n917_ = new_n297_ & new_n765_;
  assign new_n918_ = ~new_n916_ & ~new_n917_;
  assign new_n919_ = new_n297_ & new_n769_;
  assign new_n920_ = new_n297_ & new_n772_;
  assign new_n921_ = ~new_n919_ & ~new_n920_;
  assign new_n922_ = new_n918_ & new_n921_;
  assign new_n923_ = new_n296_ & new_n782_;
  assign new_n924_ = new_n789_ & new_n923_;
  assign new_n925_ = new_n297_ & new_n775_;
  assign new_n926_ = new_n780_ & new_n923_;
  assign new_n927_ = ~new_n925_ & ~new_n926_;
  assign new_n928_ = ~new_n924_ & new_n927_;
  assign new_n929_ = new_n922_ & new_n928_;
  assign new_n930_ = new_n915_ & new_n929_;
  assign new_n931_ = new_n296_ & new_n792_;
  assign new_n932_ = new_n780_ & new_n931_;
  assign new_n933_ = new_n789_ & new_n931_;
  assign new_n934_ = ~new_n932_ & ~new_n933_;
  assign new_n935_ = new_n301_ & new_n740_;
  assign new_n936_ = new_n301_ & new_n742_;
  assign new_n937_ = ~new_n935_ & ~new_n936_;
  assign new_n938_ = new_n934_ & new_n937_;
  assign new_n939_ = new_n301_ & new_n747_;
  assign new_n940_ = new_n301_ & new_n749_;
  assign new_n941_ = new_n301_ & new_n751_;
  assign new_n942_ = ~new_n940_ & ~new_n941_;
  assign new_n943_ = ~new_n939_ & new_n942_;
  assign new_n944_ = new_n938_ & new_n943_;
  assign new_n945_ = new_n301_ & new_n758_;
  assign new_n946_ = new_n301_ & new_n760_;
  assign new_n947_ = ~new_n945_ & ~new_n946_;
  assign new_n948_ = new_n301_ & new_n763_;
  assign new_n949_ = new_n301_ & new_n765_;
  assign new_n950_ = ~new_n948_ & ~new_n949_;
  assign new_n951_ = new_n947_ & new_n950_;
  assign new_n952_ = new_n301_ & new_n775_;
  assign new_n953_ = new_n301_ & new_n769_;
  assign new_n954_ = new_n301_ & new_n772_;
  assign new_n955_ = ~new_n953_ & ~new_n954_;
  assign new_n956_ = ~new_n952_ & new_n955_;
  assign new_n957_ = new_n951_ & new_n956_;
  assign new_n958_ = new_n944_ & new_n957_;
  assign new_n959_ = new_n930_ & new_n958_;
  assign new_n960_ = new_n900_ & new_n959_;
  assign new_n961_ = new_n839_ & new_n960_;
  assign new_n962_ = new_n296_ & new_n821_;
  assign new_n963_ = new_n780_ & new_n962_;
  assign new_n964_ = new_n789_ & new_n962_;
  assign new_n965_ = ~new_n963_ & ~new_n964_;
  assign new_n966_ = new_n296_ & new_n826_;
  assign new_n967_ = new_n780_ & new_n966_;
  assign new_n968_ = new_n789_ & new_n966_;
  assign new_n969_ = ~new_n967_ & ~new_n968_;
  assign new_n970_ = new_n965_ & new_n969_;
  assign new_n971_ = new_n309_ & new_n740_;
  assign new_n972_ = new_n309_ & new_n742_;
  assign new_n973_ = ~new_n971_ & ~new_n972_;
  assign new_n974_ = new_n309_ & new_n749_;
  assign new_n975_ = new_n309_ & new_n751_;
  assign new_n976_ = ~new_n974_ & ~new_n975_;
  assign new_n977_ = new_n973_ & new_n976_;
  assign new_n978_ = new_n970_ & new_n977_;
  assign new_n979_ = new_n309_ & new_n747_;
  assign new_n980_ = new_n309_ & new_n758_;
  assign new_n981_ = ~new_n979_ & ~new_n980_;
  assign new_n982_ = new_n309_ & new_n760_;
  assign new_n983_ = new_n309_ & new_n763_;
  assign new_n984_ = ~new_n982_ & ~new_n983_;
  assign new_n985_ = new_n981_ & new_n984_;
  assign new_n986_ = new_n309_ & new_n772_;
  assign new_n987_ = new_n309_ & new_n765_;
  assign new_n988_ = new_n309_ & new_n769_;
  assign new_n989_ = ~new_n987_ & ~new_n988_;
  assign new_n990_ = ~new_n986_ & new_n989_;
  assign new_n991_ = new_n985_ & new_n990_;
  assign new_n992_ = new_n978_ & new_n991_;
  assign new_n993_ = new_n309_ & new_n775_;
  assign new_n994_ = new_n306_ & new_n782_;
  assign new_n995_ = new_n780_ & new_n994_;
  assign new_n996_ = ~new_n993_ & ~new_n995_;
  assign new_n997_ = new_n789_ & new_n994_;
  assign new_n998_ = new_n306_ & new_n792_;
  assign new_n999_ = new_n780_ & new_n998_;
  assign new_n1000_ = ~new_n997_ & ~new_n999_;
  assign new_n1001_ = new_n996_ & new_n1000_;
  assign new_n1002_ = new_n307_ & new_n742_;
  assign new_n1003_ = new_n789_ & new_n998_;
  assign new_n1004_ = new_n307_ & new_n740_;
  assign new_n1005_ = ~new_n1003_ & ~new_n1004_;
  assign new_n1006_ = ~new_n1002_ & new_n1005_;
  assign new_n1007_ = new_n1001_ & new_n1006_;
  assign new_n1008_ = new_n307_ & new_n749_;
  assign new_n1009_ = new_n307_ & new_n751_;
  assign new_n1010_ = ~new_n1008_ & ~new_n1009_;
  assign new_n1011_ = new_n307_ & new_n747_;
  assign new_n1012_ = new_n307_ & new_n758_;
  assign new_n1013_ = ~new_n1011_ & ~new_n1012_;
  assign new_n1014_ = new_n1010_ & new_n1013_;
  assign new_n1015_ = new_n307_ & new_n765_;
  assign new_n1016_ = new_n307_ & new_n760_;
  assign new_n1017_ = new_n307_ & new_n763_;
  assign new_n1018_ = ~new_n1016_ & ~new_n1017_;
  assign new_n1019_ = ~new_n1015_ & new_n1018_;
  assign new_n1020_ = new_n1014_ & new_n1019_;
  assign new_n1021_ = new_n1007_ & new_n1020_;
  assign new_n1022_ = new_n992_ & new_n1021_;
  assign new_n1023_ = new_n307_ & new_n769_;
  assign new_n1024_ = new_n307_ & new_n772_;
  assign new_n1025_ = ~new_n1023_ & ~new_n1024_;
  assign new_n1026_ = new_n307_ & new_n775_;
  assign new_n1027_ = new_n306_ & new_n821_;
  assign new_n1028_ = new_n780_ & new_n1027_;
  assign new_n1029_ = ~new_n1026_ & ~new_n1028_;
  assign new_n1030_ = new_n1025_ & new_n1029_;
  assign new_n1031_ = new_n789_ & new_n1027_;
  assign new_n1032_ = new_n306_ & new_n826_;
  assign new_n1033_ = new_n780_ & new_n1032_;
  assign new_n1034_ = ~new_n1031_ & ~new_n1033_;
  assign new_n1035_ = new_n789_ & new_n1032_;
  assign new_n1036_ = ~A200 & ~A199;
  assign new_n1037_ = new_n264_ & new_n1036_;
  assign new_n1038_ = ~A168 & ~A169;
  assign new_n1039_ = A170 & new_n1038_;
  assign new_n1040_ = new_n1037_ & new_n1039_;
  assign new_n1041_ = new_n543_ & new_n1040_;
  assign new_n1042_ = ~new_n1035_ & ~new_n1041_;
  assign new_n1043_ = new_n1034_ & new_n1042_;
  assign new_n1044_ = new_n1030_ & new_n1043_;
  assign new_n1045_ = new_n553_ & new_n1040_;
  assign new_n1046_ = new_n78_ & new_n781_;
  assign new_n1047_ = new_n318_ & new_n1046_;
  assign new_n1048_ = new_n262_ & new_n264_;
  assign new_n1049_ = new_n1039_ & new_n1048_;
  assign new_n1050_ = new_n1047_ & new_n1049_;
  assign new_n1051_ = ~new_n1045_ & ~new_n1050_;
  assign new_n1052_ = new_n322_ & new_n1046_;
  assign new_n1053_ = new_n1049_ & new_n1052_;
  assign new_n1054_ = new_n325_ & new_n1046_;
  assign new_n1055_ = new_n1049_ & new_n1054_;
  assign new_n1056_ = ~new_n1053_ & ~new_n1055_;
  assign new_n1057_ = new_n1051_ & new_n1056_;
  assign new_n1058_ = new_n337_ & new_n1046_;
  assign new_n1059_ = new_n1049_ & new_n1058_;
  assign new_n1060_ = new_n330_ & new_n1046_;
  assign new_n1061_ = new_n1049_ & new_n1060_;
  assign new_n1062_ = new_n333_ & new_n1046_;
  assign new_n1063_ = new_n1049_ & new_n1062_;
  assign new_n1064_ = ~new_n1061_ & ~new_n1063_;
  assign new_n1065_ = ~new_n1059_ & new_n1064_;
  assign new_n1066_ = new_n1057_ & new_n1065_;
  assign new_n1067_ = new_n1044_ & new_n1066_;
  assign new_n1068_ = new_n340_ & new_n1046_;
  assign new_n1069_ = new_n1049_ & new_n1068_;
  assign new_n1070_ = new_n346_ & new_n1046_;
  assign new_n1071_ = new_n1049_ & new_n1070_;
  assign new_n1072_ = ~new_n1069_ & ~new_n1071_;
  assign new_n1073_ = new_n104_ & new_n781_;
  assign new_n1074_ = new_n318_ & new_n1073_;
  assign new_n1075_ = new_n1049_ & new_n1074_;
  assign new_n1076_ = new_n322_ & new_n1073_;
  assign new_n1077_ = new_n1049_ & new_n1076_;
  assign new_n1078_ = ~new_n1075_ & ~new_n1077_;
  assign new_n1079_ = new_n1072_ & new_n1078_;
  assign new_n1080_ = new_n333_ & new_n1073_;
  assign new_n1081_ = new_n1049_ & new_n1080_;
  assign new_n1082_ = new_n325_ & new_n1073_;
  assign new_n1083_ = new_n1049_ & new_n1082_;
  assign new_n1084_ = new_n330_ & new_n1073_;
  assign new_n1085_ = new_n1049_ & new_n1084_;
  assign new_n1086_ = ~new_n1083_ & ~new_n1085_;
  assign new_n1087_ = ~new_n1081_ & new_n1086_;
  assign new_n1088_ = new_n1079_ & new_n1087_;
  assign new_n1089_ = new_n337_ & new_n1073_;
  assign new_n1090_ = new_n1049_ & new_n1089_;
  assign new_n1091_ = new_n340_ & new_n1073_;
  assign new_n1092_ = new_n1049_ & new_n1091_;
  assign new_n1093_ = ~new_n1090_ & ~new_n1092_;
  assign new_n1094_ = new_n346_ & new_n1073_;
  assign new_n1095_ = new_n1049_ & new_n1094_;
  assign new_n1096_ = new_n78_ & new_n791_;
  assign new_n1097_ = new_n318_ & new_n1096_;
  assign new_n1098_ = new_n1049_ & new_n1097_;
  assign new_n1099_ = ~new_n1095_ & ~new_n1098_;
  assign new_n1100_ = new_n1093_ & new_n1099_;
  assign new_n1101_ = new_n330_ & new_n1096_;
  assign new_n1102_ = new_n1049_ & new_n1101_;
  assign new_n1103_ = new_n322_ & new_n1096_;
  assign new_n1104_ = new_n1049_ & new_n1103_;
  assign new_n1105_ = new_n325_ & new_n1096_;
  assign new_n1106_ = new_n1049_ & new_n1105_;
  assign new_n1107_ = ~new_n1104_ & ~new_n1106_;
  assign new_n1108_ = ~new_n1102_ & new_n1107_;
  assign new_n1109_ = new_n1100_ & new_n1108_;
  assign new_n1110_ = new_n1088_ & new_n1109_;
  assign new_n1111_ = new_n1067_ & new_n1110_;
  assign new_n1112_ = new_n1022_ & new_n1111_;
  assign new_n1113_ = new_n333_ & new_n1096_;
  assign new_n1114_ = new_n1049_ & new_n1113_;
  assign new_n1115_ = new_n337_ & new_n1096_;
  assign new_n1116_ = new_n1049_ & new_n1115_;
  assign new_n1117_ = ~new_n1114_ & ~new_n1116_;
  assign new_n1118_ = new_n340_ & new_n1096_;
  assign new_n1119_ = new_n1049_ & new_n1118_;
  assign new_n1120_ = new_n346_ & new_n1096_;
  assign new_n1121_ = new_n1049_ & new_n1120_;
  assign new_n1122_ = ~new_n1119_ & ~new_n1121_;
  assign new_n1123_ = new_n1117_ & new_n1122_;
  assign new_n1124_ = new_n104_ & new_n791_;
  assign new_n1125_ = new_n318_ & new_n1124_;
  assign new_n1126_ = new_n1049_ & new_n1125_;
  assign new_n1127_ = new_n322_ & new_n1124_;
  assign new_n1128_ = new_n1049_ & new_n1127_;
  assign new_n1129_ = ~new_n1126_ & ~new_n1128_;
  assign new_n1130_ = new_n325_ & new_n1124_;
  assign new_n1131_ = new_n1049_ & new_n1130_;
  assign new_n1132_ = new_n330_ & new_n1124_;
  assign new_n1133_ = new_n1049_ & new_n1132_;
  assign new_n1134_ = ~new_n1131_ & ~new_n1133_;
  assign new_n1135_ = new_n1129_ & new_n1134_;
  assign new_n1136_ = new_n1123_ & new_n1135_;
  assign new_n1137_ = new_n333_ & new_n1124_;
  assign new_n1138_ = new_n1049_ & new_n1137_;
  assign new_n1139_ = new_n337_ & new_n1124_;
  assign new_n1140_ = new_n1049_ & new_n1139_;
  assign new_n1141_ = ~new_n1138_ & ~new_n1140_;
  assign new_n1142_ = new_n340_ & new_n1124_;
  assign new_n1143_ = new_n1049_ & new_n1142_;
  assign new_n1144_ = new_n346_ & new_n1124_;
  assign new_n1145_ = new_n1049_ & new_n1144_;
  assign new_n1146_ = ~new_n1143_ & ~new_n1145_;
  assign new_n1147_ = new_n1141_ & new_n1146_;
  assign new_n1148_ = new_n264_ & new_n276_;
  assign new_n1149_ = new_n1039_ & new_n1148_;
  assign new_n1150_ = new_n1054_ & new_n1149_;
  assign new_n1151_ = new_n1047_ & new_n1149_;
  assign new_n1152_ = new_n1052_ & new_n1149_;
  assign new_n1153_ = ~new_n1151_ & ~new_n1152_;
  assign new_n1154_ = ~new_n1150_ & new_n1153_;
  assign new_n1155_ = new_n1147_ & new_n1154_;
  assign new_n1156_ = new_n1136_ & new_n1155_;
  assign new_n1157_ = new_n1060_ & new_n1149_;
  assign new_n1158_ = new_n1062_ & new_n1149_;
  assign new_n1159_ = ~new_n1157_ & ~new_n1158_;
  assign new_n1160_ = new_n1058_ & new_n1149_;
  assign new_n1161_ = new_n1068_ & new_n1149_;
  assign new_n1162_ = ~new_n1160_ & ~new_n1161_;
  assign new_n1163_ = new_n1159_ & new_n1162_;
  assign new_n1164_ = new_n1076_ & new_n1149_;
  assign new_n1165_ = new_n1070_ & new_n1149_;
  assign new_n1166_ = new_n1074_ & new_n1149_;
  assign new_n1167_ = ~new_n1165_ & ~new_n1166_;
  assign new_n1168_ = ~new_n1164_ & new_n1167_;
  assign new_n1169_ = new_n1163_ & new_n1168_;
  assign new_n1170_ = new_n1082_ & new_n1149_;
  assign new_n1171_ = new_n1084_ & new_n1149_;
  assign new_n1172_ = ~new_n1170_ & ~new_n1171_;
  assign new_n1173_ = new_n1080_ & new_n1149_;
  assign new_n1174_ = new_n1089_ & new_n1149_;
  assign new_n1175_ = ~new_n1173_ & ~new_n1174_;
  assign new_n1176_ = new_n1172_ & new_n1175_;
  assign new_n1177_ = new_n1097_ & new_n1149_;
  assign new_n1178_ = new_n1091_ & new_n1149_;
  assign new_n1179_ = new_n1094_ & new_n1149_;
  assign new_n1180_ = ~new_n1178_ & ~new_n1179_;
  assign new_n1181_ = ~new_n1177_ & new_n1180_;
  assign new_n1182_ = new_n1176_ & new_n1181_;
  assign new_n1183_ = new_n1169_ & new_n1182_;
  assign new_n1184_ = new_n1156_ & new_n1183_;
  assign new_n1185_ = new_n1103_ & new_n1149_;
  assign new_n1186_ = new_n1105_ & new_n1149_;
  assign new_n1187_ = ~new_n1185_ & ~new_n1186_;
  assign new_n1188_ = new_n1101_ & new_n1149_;
  assign new_n1189_ = new_n1113_ & new_n1149_;
  assign new_n1190_ = ~new_n1188_ & ~new_n1189_;
  assign new_n1191_ = new_n1187_ & new_n1190_;
  assign new_n1192_ = new_n1120_ & new_n1149_;
  assign new_n1193_ = new_n1115_ & new_n1149_;
  assign new_n1194_ = new_n1118_ & new_n1149_;
  assign new_n1195_ = ~new_n1193_ & ~new_n1194_;
  assign new_n1196_ = ~new_n1192_ & new_n1195_;
  assign new_n1197_ = new_n1191_ & new_n1196_;
  assign new_n1198_ = new_n1125_ & new_n1149_;
  assign new_n1199_ = new_n1127_ & new_n1149_;
  assign new_n1200_ = ~new_n1198_ & ~new_n1199_;
  assign new_n1201_ = new_n1130_ & new_n1149_;
  assign new_n1202_ = new_n1132_ & new_n1149_;
  assign new_n1203_ = ~new_n1201_ & ~new_n1202_;
  assign new_n1204_ = new_n1200_ & new_n1203_;
  assign new_n1205_ = new_n1142_ & new_n1149_;
  assign new_n1206_ = new_n1137_ & new_n1149_;
  assign new_n1207_ = new_n1139_ & new_n1149_;
  assign new_n1208_ = ~new_n1206_ & ~new_n1207_;
  assign new_n1209_ = ~new_n1205_ & new_n1208_;
  assign new_n1210_ = new_n1204_ & new_n1209_;
  assign new_n1211_ = new_n1197_ & new_n1210_;
  assign new_n1212_ = new_n1144_ & new_n1149_;
  assign new_n1213_ = A200 & A199;
  assign new_n1214_ = new_n264_ & new_n1213_;
  assign new_n1215_ = new_n1039_ & new_n1214_;
  assign new_n1216_ = new_n543_ & new_n1215_;
  assign new_n1217_ = ~new_n1212_ & ~new_n1216_;
  assign new_n1218_ = new_n553_ & new_n1215_;
  assign new_n1219_ = A203 & ~A201;
  assign new_n1220_ = new_n264_ & new_n1219_;
  assign new_n1221_ = new_n1039_ & new_n1220_;
  assign new_n1222_ = new_n543_ & new_n1221_;
  assign new_n1223_ = ~new_n1218_ & ~new_n1222_;
  assign new_n1224_ = new_n1217_ & new_n1223_;
  assign new_n1225_ = A202 & ~A201;
  assign new_n1226_ = new_n264_ & new_n1225_;
  assign new_n1227_ = new_n1039_ & new_n1226_;
  assign new_n1228_ = new_n553_ & new_n1227_;
  assign new_n1229_ = new_n553_ & new_n1221_;
  assign new_n1230_ = new_n543_ & new_n1227_;
  assign new_n1231_ = ~new_n1229_ & ~new_n1230_;
  assign new_n1232_ = ~new_n1228_ & new_n1231_;
  assign new_n1233_ = new_n1224_ & new_n1232_;
  assign new_n1234_ = ~A298 & ~A266;
  assign new_n1235_ = new_n45_ & new_n1234_;
  assign new_n1236_ = new_n539_ & new_n1235_;
  assign new_n1237_ = ~A202 & A201;
  assign new_n1238_ = new_n264_ & new_n1237_;
  assign new_n1239_ = new_n1039_ & new_n1238_;
  assign new_n1240_ = new_n1236_ & new_n1239_;
  assign new_n1241_ = A298 & ~A266;
  assign new_n1242_ = new_n45_ & new_n1241_;
  assign new_n1243_ = new_n550_ & new_n1242_;
  assign new_n1244_ = new_n1239_ & new_n1243_;
  assign new_n1245_ = ~new_n1240_ & ~new_n1244_;
  assign new_n1246_ = ~A298 & A266;
  assign new_n1247_ = new_n32_ & new_n1246_;
  assign new_n1248_ = new_n539_ & new_n1247_;
  assign new_n1249_ = new_n1239_ & new_n1248_;
  assign new_n1250_ = A298 & A266;
  assign new_n1251_ = new_n32_ & new_n1250_;
  assign new_n1252_ = new_n550_ & new_n1251_;
  assign new_n1253_ = new_n1239_ & new_n1252_;
  assign new_n1254_ = ~new_n1249_ & ~new_n1253_;
  assign new_n1255_ = new_n1245_ & new_n1254_;
  assign new_n1256_ = ~A298 & A268;
  assign new_n1257_ = ~A267 & ~A203;
  assign new_n1258_ = new_n1256_ & new_n1257_;
  assign new_n1259_ = new_n539_ & new_n1258_;
  assign new_n1260_ = new_n1239_ & new_n1259_;
  assign new_n1261_ = ~A298 & A269;
  assign new_n1262_ = new_n1257_ & new_n1261_;
  assign new_n1263_ = new_n539_ & new_n1262_;
  assign new_n1264_ = new_n1239_ & new_n1263_;
  assign new_n1265_ = A298 & A269;
  assign new_n1266_ = new_n1257_ & new_n1265_;
  assign new_n1267_ = new_n550_ & new_n1266_;
  assign new_n1268_ = new_n1239_ & new_n1267_;
  assign new_n1269_ = ~new_n1264_ & ~new_n1268_;
  assign new_n1270_ = ~new_n1260_ & new_n1269_;
  assign new_n1271_ = new_n1255_ & new_n1270_;
  assign new_n1272_ = new_n1233_ & new_n1271_;
  assign new_n1273_ = new_n1211_ & new_n1272_;
  assign new_n1274_ = new_n1184_ & new_n1273_;
  assign new_n1275_ = new_n1112_ & new_n1274_;
  assign new_n1276_ = new_n961_ & new_n1275_;
  assign new_n1277_ = new_n683_ & new_n1276_;
  assign new_n1278_ = A298 & A268;
  assign new_n1279_ = new_n1257_ & new_n1278_;
  assign new_n1280_ = new_n550_ & new_n1279_;
  assign new_n1281_ = new_n1239_ & new_n1280_;
  assign new_n1282_ = A302 & A300;
  assign new_n1283_ = A299 & ~A298;
  assign new_n1284_ = new_n1282_ & new_n1283_;
  assign new_n1285_ = A267 & ~A203;
  assign new_n1286_ = new_n29_ & new_n1285_;
  assign new_n1287_ = new_n1284_ & new_n1286_;
  assign new_n1288_ = new_n1239_ & new_n1287_;
  assign new_n1289_ = ~new_n1281_ & ~new_n1288_;
  assign new_n1290_ = A301 & A300;
  assign new_n1291_ = new_n1283_ & new_n1290_;
  assign new_n1292_ = new_n1286_ & new_n1291_;
  assign new_n1293_ = new_n1239_ & new_n1292_;
  assign new_n1294_ = ~A299 & A298;
  assign new_n1295_ = new_n1282_ & new_n1294_;
  assign new_n1296_ = new_n1286_ & new_n1295_;
  assign new_n1297_ = new_n1239_ & new_n1296_;
  assign new_n1298_ = ~new_n1293_ & ~new_n1297_;
  assign new_n1299_ = new_n1289_ & new_n1298_;
  assign new_n1300_ = new_n1290_ & new_n1294_;
  assign new_n1301_ = new_n1286_ & new_n1300_;
  assign new_n1302_ = new_n1239_ & new_n1301_;
  assign new_n1303_ = new_n282_ & new_n1036_;
  assign new_n1304_ = new_n1039_ & new_n1303_;
  assign new_n1305_ = new_n543_ & new_n1304_;
  assign new_n1306_ = ~new_n1302_ & ~new_n1305_;
  assign new_n1307_ = new_n553_ & new_n1304_;
  assign new_n1308_ = new_n262_ & new_n282_;
  assign new_n1309_ = new_n1039_ & new_n1308_;
  assign new_n1310_ = new_n1047_ & new_n1309_;
  assign new_n1311_ = ~new_n1307_ & ~new_n1310_;
  assign new_n1312_ = new_n1306_ & new_n1311_;
  assign new_n1313_ = new_n1299_ & new_n1312_;
  assign new_n1314_ = new_n1052_ & new_n1309_;
  assign new_n1315_ = new_n1054_ & new_n1309_;
  assign new_n1316_ = ~new_n1314_ & ~new_n1315_;
  assign new_n1317_ = new_n1060_ & new_n1309_;
  assign new_n1318_ = new_n1062_ & new_n1309_;
  assign new_n1319_ = ~new_n1317_ & ~new_n1318_;
  assign new_n1320_ = new_n1316_ & new_n1319_;
  assign new_n1321_ = new_n1070_ & new_n1309_;
  assign new_n1322_ = new_n1058_ & new_n1309_;
  assign new_n1323_ = new_n1068_ & new_n1309_;
  assign new_n1324_ = ~new_n1322_ & ~new_n1323_;
  assign new_n1325_ = ~new_n1321_ & new_n1324_;
  assign new_n1326_ = new_n1320_ & new_n1325_;
  assign new_n1327_ = new_n1313_ & new_n1326_;
  assign new_n1328_ = new_n1074_ & new_n1309_;
  assign new_n1329_ = new_n1076_ & new_n1309_;
  assign new_n1330_ = ~new_n1328_ & ~new_n1329_;
  assign new_n1331_ = new_n1082_ & new_n1309_;
  assign new_n1332_ = new_n1084_ & new_n1309_;
  assign new_n1333_ = ~new_n1331_ & ~new_n1332_;
  assign new_n1334_ = new_n1330_ & new_n1333_;
  assign new_n1335_ = new_n1091_ & new_n1309_;
  assign new_n1336_ = new_n1080_ & new_n1309_;
  assign new_n1337_ = new_n1089_ & new_n1309_;
  assign new_n1338_ = ~new_n1336_ & ~new_n1337_;
  assign new_n1339_ = ~new_n1335_ & new_n1338_;
  assign new_n1340_ = new_n1334_ & new_n1339_;
  assign new_n1341_ = new_n1094_ & new_n1309_;
  assign new_n1342_ = new_n1097_ & new_n1309_;
  assign new_n1343_ = ~new_n1341_ & ~new_n1342_;
  assign new_n1344_ = new_n1103_ & new_n1309_;
  assign new_n1345_ = new_n1105_ & new_n1309_;
  assign new_n1346_ = ~new_n1344_ & ~new_n1345_;
  assign new_n1347_ = new_n1343_ & new_n1346_;
  assign new_n1348_ = new_n1115_ & new_n1309_;
  assign new_n1349_ = new_n1101_ & new_n1309_;
  assign new_n1350_ = new_n1113_ & new_n1309_;
  assign new_n1351_ = ~new_n1349_ & ~new_n1350_;
  assign new_n1352_ = ~new_n1348_ & new_n1351_;
  assign new_n1353_ = new_n1347_ & new_n1352_;
  assign new_n1354_ = new_n1340_ & new_n1353_;
  assign new_n1355_ = new_n1327_ & new_n1354_;
  assign new_n1356_ = new_n1118_ & new_n1309_;
  assign new_n1357_ = new_n1120_ & new_n1309_;
  assign new_n1358_ = ~new_n1356_ & ~new_n1357_;
  assign new_n1359_ = new_n1125_ & new_n1309_;
  assign new_n1360_ = new_n1127_ & new_n1309_;
  assign new_n1361_ = ~new_n1359_ & ~new_n1360_;
  assign new_n1362_ = new_n1358_ & new_n1361_;
  assign new_n1363_ = new_n1130_ & new_n1309_;
  assign new_n1364_ = new_n1132_ & new_n1309_;
  assign new_n1365_ = ~new_n1363_ & ~new_n1364_;
  assign new_n1366_ = new_n1137_ & new_n1309_;
  assign new_n1367_ = new_n1139_ & new_n1309_;
  assign new_n1368_ = ~new_n1366_ & ~new_n1367_;
  assign new_n1369_ = new_n1365_ & new_n1368_;
  assign new_n1370_ = new_n1362_ & new_n1369_;
  assign new_n1371_ = new_n1142_ & new_n1309_;
  assign new_n1372_ = new_n1144_ & new_n1309_;
  assign new_n1373_ = ~new_n1371_ & ~new_n1372_;
  assign new_n1374_ = new_n276_ & new_n282_;
  assign new_n1375_ = new_n1039_ & new_n1374_;
  assign new_n1376_ = new_n1047_ & new_n1375_;
  assign new_n1377_ = new_n1052_ & new_n1375_;
  assign new_n1378_ = ~new_n1376_ & ~new_n1377_;
  assign new_n1379_ = new_n1373_ & new_n1378_;
  assign new_n1380_ = new_n1062_ & new_n1375_;
  assign new_n1381_ = new_n1054_ & new_n1375_;
  assign new_n1382_ = new_n1060_ & new_n1375_;
  assign new_n1383_ = ~new_n1381_ & ~new_n1382_;
  assign new_n1384_ = ~new_n1380_ & new_n1383_;
  assign new_n1385_ = new_n1379_ & new_n1384_;
  assign new_n1386_ = new_n1370_ & new_n1385_;
  assign new_n1387_ = new_n1058_ & new_n1375_;
  assign new_n1388_ = new_n1068_ & new_n1375_;
  assign new_n1389_ = ~new_n1387_ & ~new_n1388_;
  assign new_n1390_ = new_n1070_ & new_n1375_;
  assign new_n1391_ = new_n1074_ & new_n1375_;
  assign new_n1392_ = ~new_n1390_ & ~new_n1391_;
  assign new_n1393_ = new_n1389_ & new_n1392_;
  assign new_n1394_ = new_n1084_ & new_n1375_;
  assign new_n1395_ = new_n1076_ & new_n1375_;
  assign new_n1396_ = new_n1082_ & new_n1375_;
  assign new_n1397_ = ~new_n1395_ & ~new_n1396_;
  assign new_n1398_ = ~new_n1394_ & new_n1397_;
  assign new_n1399_ = new_n1393_ & new_n1398_;
  assign new_n1400_ = new_n1080_ & new_n1375_;
  assign new_n1401_ = new_n1089_ & new_n1375_;
  assign new_n1402_ = ~new_n1400_ & ~new_n1401_;
  assign new_n1403_ = new_n1091_ & new_n1375_;
  assign new_n1404_ = new_n1094_ & new_n1375_;
  assign new_n1405_ = ~new_n1403_ & ~new_n1404_;
  assign new_n1406_ = new_n1402_ & new_n1405_;
  assign new_n1407_ = new_n1105_ & new_n1375_;
  assign new_n1408_ = new_n1097_ & new_n1375_;
  assign new_n1409_ = new_n1103_ & new_n1375_;
  assign new_n1410_ = ~new_n1408_ & ~new_n1409_;
  assign new_n1411_ = ~new_n1407_ & new_n1410_;
  assign new_n1412_ = new_n1406_ & new_n1411_;
  assign new_n1413_ = new_n1399_ & new_n1412_;
  assign new_n1414_ = new_n1386_ & new_n1413_;
  assign new_n1415_ = new_n1355_ & new_n1414_;
  assign new_n1416_ = new_n1101_ & new_n1375_;
  assign new_n1417_ = new_n1113_ & new_n1375_;
  assign new_n1418_ = ~new_n1416_ & ~new_n1417_;
  assign new_n1419_ = new_n1115_ & new_n1375_;
  assign new_n1420_ = new_n1118_ & new_n1375_;
  assign new_n1421_ = ~new_n1419_ & ~new_n1420_;
  assign new_n1422_ = new_n1418_ & new_n1421_;
  assign new_n1423_ = new_n1120_ & new_n1375_;
  assign new_n1424_ = new_n1125_ & new_n1375_;
  assign new_n1425_ = ~new_n1423_ & ~new_n1424_;
  assign new_n1426_ = new_n1127_ & new_n1375_;
  assign new_n1427_ = new_n1130_ & new_n1375_;
  assign new_n1428_ = ~new_n1426_ & ~new_n1427_;
  assign new_n1429_ = new_n1425_ & new_n1428_;
  assign new_n1430_ = new_n1422_ & new_n1429_;
  assign new_n1431_ = new_n1132_ & new_n1375_;
  assign new_n1432_ = new_n1137_ & new_n1375_;
  assign new_n1433_ = ~new_n1431_ & ~new_n1432_;
  assign new_n1434_ = new_n1139_ & new_n1375_;
  assign new_n1435_ = new_n1142_ & new_n1375_;
  assign new_n1436_ = ~new_n1434_ & ~new_n1435_;
  assign new_n1437_ = new_n1433_ & new_n1436_;
  assign new_n1438_ = new_n282_ & new_n1213_;
  assign new_n1439_ = new_n1039_ & new_n1438_;
  assign new_n1440_ = new_n553_ & new_n1439_;
  assign new_n1441_ = new_n1144_ & new_n1375_;
  assign new_n1442_ = new_n543_ & new_n1439_;
  assign new_n1443_ = ~new_n1441_ & ~new_n1442_;
  assign new_n1444_ = ~new_n1440_ & new_n1443_;
  assign new_n1445_ = new_n1437_ & new_n1444_;
  assign new_n1446_ = new_n1430_ & new_n1445_;
  assign new_n1447_ = new_n282_ & new_n1219_;
  assign new_n1448_ = new_n1039_ & new_n1447_;
  assign new_n1449_ = new_n543_ & new_n1448_;
  assign new_n1450_ = new_n553_ & new_n1448_;
  assign new_n1451_ = ~new_n1449_ & ~new_n1450_;
  assign new_n1452_ = new_n282_ & new_n1225_;
  assign new_n1453_ = new_n1039_ & new_n1452_;
  assign new_n1454_ = new_n543_ & new_n1453_;
  assign new_n1455_ = new_n553_ & new_n1453_;
  assign new_n1456_ = ~new_n1454_ & ~new_n1455_;
  assign new_n1457_ = new_n1451_ & new_n1456_;
  assign new_n1458_ = new_n282_ & new_n1237_;
  assign new_n1459_ = new_n1039_ & new_n1458_;
  assign new_n1460_ = new_n1248_ & new_n1459_;
  assign new_n1461_ = new_n1236_ & new_n1459_;
  assign new_n1462_ = new_n1243_ & new_n1459_;
  assign new_n1463_ = ~new_n1461_ & ~new_n1462_;
  assign new_n1464_ = ~new_n1460_ & new_n1463_;
  assign new_n1465_ = new_n1457_ & new_n1464_;
  assign new_n1466_ = new_n1252_ & new_n1459_;
  assign new_n1467_ = new_n1263_ & new_n1459_;
  assign new_n1468_ = ~new_n1466_ & ~new_n1467_;
  assign new_n1469_ = new_n1267_ & new_n1459_;
  assign new_n1470_ = new_n1259_ & new_n1459_;
  assign new_n1471_ = ~new_n1469_ & ~new_n1470_;
  assign new_n1472_ = new_n1468_ & new_n1471_;
  assign new_n1473_ = new_n1292_ & new_n1459_;
  assign new_n1474_ = new_n1280_ & new_n1459_;
  assign new_n1475_ = new_n1287_ & new_n1459_;
  assign new_n1476_ = ~new_n1474_ & ~new_n1475_;
  assign new_n1477_ = ~new_n1473_ & new_n1476_;
  assign new_n1478_ = new_n1472_ & new_n1477_;
  assign new_n1479_ = new_n1465_ & new_n1478_;
  assign new_n1480_ = new_n1446_ & new_n1479_;
  assign new_n1481_ = new_n1296_ & new_n1459_;
  assign new_n1482_ = new_n1301_ & new_n1459_;
  assign new_n1483_ = ~new_n1481_ & ~new_n1482_;
  assign new_n1484_ = A168 & ~A169;
  assign new_n1485_ = A170 & new_n1484_;
  assign new_n1486_ = new_n263_ & new_n1485_;
  assign new_n1487_ = new_n1236_ & new_n1486_;
  assign new_n1488_ = new_n1243_ & new_n1486_;
  assign new_n1489_ = ~new_n1487_ & ~new_n1488_;
  assign new_n1490_ = new_n1483_ & new_n1489_;
  assign new_n1491_ = new_n1248_ & new_n1486_;
  assign new_n1492_ = new_n1252_ & new_n1486_;
  assign new_n1493_ = ~new_n1491_ & ~new_n1492_;
  assign new_n1494_ = new_n1263_ & new_n1486_;
  assign new_n1495_ = new_n1267_ & new_n1486_;
  assign new_n1496_ = ~new_n1494_ & ~new_n1495_;
  assign new_n1497_ = new_n1493_ & new_n1496_;
  assign new_n1498_ = new_n1490_ & new_n1497_;
  assign new_n1499_ = new_n1259_ & new_n1486_;
  assign new_n1500_ = new_n1280_ & new_n1486_;
  assign new_n1501_ = ~new_n1499_ & ~new_n1500_;
  assign new_n1502_ = new_n1287_ & new_n1486_;
  assign new_n1503_ = new_n1292_ & new_n1486_;
  assign new_n1504_ = ~new_n1502_ & ~new_n1503_;
  assign new_n1505_ = new_n1501_ & new_n1504_;
  assign new_n1506_ = new_n782_ & new_n1485_;
  assign new_n1507_ = new_n543_ & new_n1506_;
  assign new_n1508_ = new_n1296_ & new_n1486_;
  assign new_n1509_ = new_n1301_ & new_n1486_;
  assign new_n1510_ = ~new_n1508_ & ~new_n1509_;
  assign new_n1511_ = ~new_n1507_ & new_n1510_;
  assign new_n1512_ = new_n1505_ & new_n1511_;
  assign new_n1513_ = new_n1498_ & new_n1512_;
  assign new_n1514_ = new_n553_ & new_n1506_;
  assign new_n1515_ = new_n792_ & new_n1485_;
  assign new_n1516_ = new_n543_ & new_n1515_;
  assign new_n1517_ = ~new_n1514_ & ~new_n1516_;
  assign new_n1518_ = new_n553_ & new_n1515_;
  assign new_n1519_ = new_n277_ & new_n1485_;
  assign new_n1520_ = new_n1236_ & new_n1519_;
  assign new_n1521_ = ~new_n1518_ & ~new_n1520_;
  assign new_n1522_ = new_n1517_ & new_n1521_;
  assign new_n1523_ = new_n1252_ & new_n1519_;
  assign new_n1524_ = new_n1243_ & new_n1519_;
  assign new_n1525_ = new_n1248_ & new_n1519_;
  assign new_n1526_ = ~new_n1524_ & ~new_n1525_;
  assign new_n1527_ = ~new_n1523_ & new_n1526_;
  assign new_n1528_ = new_n1522_ & new_n1527_;
  assign new_n1529_ = new_n1263_ & new_n1519_;
  assign new_n1530_ = new_n1267_ & new_n1519_;
  assign new_n1531_ = ~new_n1529_ & ~new_n1530_;
  assign new_n1532_ = new_n1259_ & new_n1519_;
  assign new_n1533_ = new_n1280_ & new_n1519_;
  assign new_n1534_ = ~new_n1532_ & ~new_n1533_;
  assign new_n1535_ = new_n1531_ & new_n1534_;
  assign new_n1536_ = new_n1296_ & new_n1519_;
  assign new_n1537_ = new_n1287_ & new_n1519_;
  assign new_n1538_ = new_n1292_ & new_n1519_;
  assign new_n1539_ = ~new_n1537_ & ~new_n1538_;
  assign new_n1540_ = ~new_n1536_ & new_n1539_;
  assign new_n1541_ = new_n1535_ & new_n1540_;
  assign new_n1542_ = new_n1528_ & new_n1541_;
  assign new_n1543_ = new_n1513_ & new_n1542_;
  assign new_n1544_ = new_n1480_ & new_n1543_;
  assign new_n1545_ = new_n1415_ & new_n1544_;
  assign new_n1546_ = new_n1301_ & new_n1519_;
  assign new_n1547_ = new_n821_ & new_n1485_;
  assign new_n1548_ = new_n543_ & new_n1547_;
  assign new_n1549_ = ~new_n1546_ & ~new_n1548_;
  assign new_n1550_ = new_n553_ & new_n1547_;
  assign new_n1551_ = new_n826_ & new_n1485_;
  assign new_n1552_ = new_n543_ & new_n1551_;
  assign new_n1553_ = ~new_n1550_ & ~new_n1552_;
  assign new_n1554_ = new_n1549_ & new_n1553_;
  assign new_n1555_ = new_n553_ & new_n1551_;
  assign new_n1556_ = A199 & ~A168;
  assign new_n1557_ = A169 & new_n1556_;
  assign new_n1558_ = new_n723_ & new_n1557_;
  assign new_n1559_ = new_n543_ & new_n1558_;
  assign new_n1560_ = ~new_n1555_ & ~new_n1559_;
  assign new_n1561_ = new_n553_ & new_n1558_;
  assign new_n1562_ = ~A199 & ~A168;
  assign new_n1563_ = A169 & new_n1562_;
  assign new_n1564_ = new_n733_ & new_n1563_;
  assign new_n1565_ = new_n543_ & new_n1564_;
  assign new_n1566_ = ~new_n1561_ & ~new_n1565_;
  assign new_n1567_ = new_n1560_ & new_n1566_;
  assign new_n1568_ = new_n1554_ & new_n1567_;
  assign new_n1569_ = new_n553_ & new_n1564_;
  assign new_n1570_ = ~A167 & A168;
  assign new_n1571_ = A169 & new_n1570_;
  assign new_n1572_ = new_n83_ & new_n1571_;
  assign new_n1573_ = new_n319_ & new_n1572_;
  assign new_n1574_ = ~new_n1569_ & ~new_n1573_;
  assign new_n1575_ = new_n323_ & new_n1572_;
  assign new_n1576_ = new_n326_ & new_n1572_;
  assign new_n1577_ = ~new_n1575_ & ~new_n1576_;
  assign new_n1578_ = new_n1574_ & new_n1577_;
  assign new_n1579_ = new_n338_ & new_n1572_;
  assign new_n1580_ = new_n331_ & new_n1572_;
  assign new_n1581_ = new_n334_ & new_n1572_;
  assign new_n1582_ = ~new_n1580_ & ~new_n1581_;
  assign new_n1583_ = ~new_n1579_ & new_n1582_;
  assign new_n1584_ = new_n1578_ & new_n1583_;
  assign new_n1585_ = new_n1568_ & new_n1584_;
  assign new_n1586_ = new_n341_ & new_n1572_;
  assign new_n1587_ = new_n347_ & new_n1572_;
  assign new_n1588_ = ~new_n1586_ & ~new_n1587_;
  assign new_n1589_ = new_n349_ & new_n1572_;
  assign new_n1590_ = new_n352_ & new_n1572_;
  assign new_n1591_ = ~new_n1589_ & ~new_n1590_;
  assign new_n1592_ = new_n1588_ & new_n1591_;
  assign new_n1593_ = new_n362_ & new_n1572_;
  assign new_n1594_ = new_n354_ & new_n1572_;
  assign new_n1595_ = new_n360_ & new_n1572_;
  assign new_n1596_ = ~new_n1594_ & ~new_n1595_;
  assign new_n1597_ = ~new_n1593_ & new_n1596_;
  assign new_n1598_ = new_n1592_ & new_n1597_;
  assign new_n1599_ = new_n358_ & new_n1572_;
  assign new_n1600_ = new_n368_ & new_n1572_;
  assign new_n1601_ = ~new_n1599_ & ~new_n1600_;
  assign new_n1602_ = new_n370_ & new_n1572_;
  assign new_n1603_ = new_n135_ & new_n1571_;
  assign new_n1604_ = new_n374_ & new_n1603_;
  assign new_n1605_ = ~new_n1602_ & ~new_n1604_;
  assign new_n1606_ = new_n1601_ & new_n1605_;
  assign new_n1607_ = new_n391_ & new_n1603_;
  assign new_n1608_ = new_n377_ & new_n1603_;
  assign new_n1609_ = new_n388_ & new_n1603_;
  assign new_n1610_ = ~new_n1608_ & ~new_n1609_;
  assign new_n1611_ = ~new_n1607_ & new_n1610_;
  assign new_n1612_ = new_n1606_ & new_n1611_;
  assign new_n1613_ = new_n1598_ & new_n1612_;
  assign new_n1614_ = new_n1585_ & new_n1613_;
  assign new_n1615_ = new_n385_ & new_n1603_;
  assign new_n1616_ = new_n398_ & new_n1603_;
  assign new_n1617_ = ~new_n1615_ & ~new_n1616_;
  assign new_n1618_ = new_n400_ & new_n1603_;
  assign new_n1619_ = new_n403_ & new_n1603_;
  assign new_n1620_ = ~new_n1618_ & ~new_n1619_;
  assign new_n1621_ = new_n1617_ & new_n1620_;
  assign new_n1622_ = new_n405_ & new_n1603_;
  assign new_n1623_ = new_n413_ & new_n1603_;
  assign new_n1624_ = ~new_n1622_ & ~new_n1623_;
  assign new_n1625_ = new_n415_ & new_n1603_;
  assign new_n1626_ = new_n411_ & new_n1603_;
  assign new_n1627_ = ~new_n1625_ & ~new_n1626_;
  assign new_n1628_ = new_n1624_ & new_n1627_;
  assign new_n1629_ = new_n1621_ & new_n1628_;
  assign new_n1630_ = new_n424_ & new_n1603_;
  assign new_n1631_ = new_n426_ & new_n1603_;
  assign new_n1632_ = ~new_n1630_ & ~new_n1631_;
  assign new_n1633_ = new_n429_ & new_n1603_;
  assign new_n1634_ = new_n431_ & new_n1603_;
  assign new_n1635_ = ~new_n1633_ & ~new_n1634_;
  assign new_n1636_ = new_n1632_ & new_n1635_;
  assign new_n1637_ = new_n441_ & new_n1603_;
  assign new_n1638_ = new_n436_ & new_n1603_;
  assign new_n1639_ = new_n438_ & new_n1603_;
  assign new_n1640_ = ~new_n1638_ & ~new_n1639_;
  assign new_n1641_ = ~new_n1637_ & new_n1640_;
  assign new_n1642_ = new_n1636_ & new_n1641_;
  assign new_n1643_ = new_n1629_ & new_n1642_;
  assign new_n1644_ = new_n443_ & new_n1603_;
  assign new_n1645_ = new_n448_ & new_n1603_;
  assign new_n1646_ = ~new_n1644_ & ~new_n1645_;
  assign new_n1647_ = new_n450_ & new_n1603_;
  assign new_n1648_ = new_n454_ & new_n1603_;
  assign new_n1649_ = ~new_n1647_ & ~new_n1648_;
  assign new_n1650_ = new_n1646_ & new_n1649_;
  assign new_n1651_ = new_n157_ & new_n1571_;
  assign new_n1652_ = new_n323_ & new_n1651_;
  assign new_n1653_ = new_n456_ & new_n1603_;
  assign new_n1654_ = new_n319_ & new_n1651_;
  assign new_n1655_ = ~new_n1653_ & ~new_n1654_;
  assign new_n1656_ = ~new_n1652_ & new_n1655_;
  assign new_n1657_ = new_n1650_ & new_n1656_;
  assign new_n1658_ = new_n326_ & new_n1651_;
  assign new_n1659_ = new_n331_ & new_n1651_;
  assign new_n1660_ = ~new_n1658_ & ~new_n1659_;
  assign new_n1661_ = new_n334_ & new_n1651_;
  assign new_n1662_ = new_n338_ & new_n1651_;
  assign new_n1663_ = ~new_n1661_ & ~new_n1662_;
  assign new_n1664_ = new_n1660_ & new_n1663_;
  assign new_n1665_ = new_n349_ & new_n1651_;
  assign new_n1666_ = new_n341_ & new_n1651_;
  assign new_n1667_ = new_n347_ & new_n1651_;
  assign new_n1668_ = ~new_n1666_ & ~new_n1667_;
  assign new_n1669_ = ~new_n1665_ & new_n1668_;
  assign new_n1670_ = new_n1664_ & new_n1669_;
  assign new_n1671_ = new_n1657_ & new_n1670_;
  assign new_n1672_ = new_n1643_ & new_n1671_;
  assign new_n1673_ = new_n1614_ & new_n1672_;
  assign new_n1674_ = new_n352_ & new_n1651_;
  assign new_n1675_ = new_n354_ & new_n1651_;
  assign new_n1676_ = ~new_n1674_ & ~new_n1675_;
  assign new_n1677_ = new_n360_ & new_n1651_;
  assign new_n1678_ = new_n362_ & new_n1651_;
  assign new_n1679_ = ~new_n1677_ & ~new_n1678_;
  assign new_n1680_ = new_n1676_ & new_n1679_;
  assign new_n1681_ = new_n358_ & new_n1651_;
  assign new_n1682_ = new_n368_ & new_n1651_;
  assign new_n1683_ = ~new_n1681_ & ~new_n1682_;
  assign new_n1684_ = new_n370_ & new_n1651_;
  assign new_n1685_ = new_n183_ & new_n1571_;
  assign new_n1686_ = new_n374_ & new_n1685_;
  assign new_n1687_ = ~new_n1684_ & ~new_n1686_;
  assign new_n1688_ = new_n1683_ & new_n1687_;
  assign new_n1689_ = new_n1680_ & new_n1688_;
  assign new_n1690_ = new_n377_ & new_n1685_;
  assign new_n1691_ = new_n388_ & new_n1685_;
  assign new_n1692_ = ~new_n1690_ & ~new_n1691_;
  assign new_n1693_ = new_n391_ & new_n1685_;
  assign new_n1694_ = new_n385_ & new_n1685_;
  assign new_n1695_ = ~new_n1693_ & ~new_n1694_;
  assign new_n1696_ = new_n1692_ & new_n1695_;
  assign new_n1697_ = new_n403_ & new_n1685_;
  assign new_n1698_ = new_n398_ & new_n1685_;
  assign new_n1699_ = new_n400_ & new_n1685_;
  assign new_n1700_ = ~new_n1698_ & ~new_n1699_;
  assign new_n1701_ = ~new_n1697_ & new_n1700_;
  assign new_n1702_ = new_n1696_ & new_n1701_;
  assign new_n1703_ = new_n1689_ & new_n1702_;
  assign new_n1704_ = new_n405_ & new_n1685_;
  assign new_n1705_ = new_n413_ & new_n1685_;
  assign new_n1706_ = ~new_n1704_ & ~new_n1705_;
  assign new_n1707_ = new_n415_ & new_n1685_;
  assign new_n1708_ = new_n411_ & new_n1685_;
  assign new_n1709_ = ~new_n1707_ & ~new_n1708_;
  assign new_n1710_ = new_n1706_ & new_n1709_;
  assign new_n1711_ = new_n429_ & new_n1685_;
  assign new_n1712_ = new_n424_ & new_n1685_;
  assign new_n1713_ = new_n426_ & new_n1685_;
  assign new_n1714_ = ~new_n1712_ & ~new_n1713_;
  assign new_n1715_ = ~new_n1711_ & new_n1714_;
  assign new_n1716_ = new_n1710_ & new_n1715_;
  assign new_n1717_ = new_n431_ & new_n1685_;
  assign new_n1718_ = new_n436_ & new_n1685_;
  assign new_n1719_ = ~new_n1717_ & ~new_n1718_;
  assign new_n1720_ = new_n438_ & new_n1685_;
  assign new_n1721_ = new_n441_ & new_n1685_;
  assign new_n1722_ = ~new_n1720_ & ~new_n1721_;
  assign new_n1723_ = new_n1719_ & new_n1722_;
  assign new_n1724_ = new_n450_ & new_n1685_;
  assign new_n1725_ = new_n443_ & new_n1685_;
  assign new_n1726_ = new_n448_ & new_n1685_;
  assign new_n1727_ = ~new_n1725_ & ~new_n1726_;
  assign new_n1728_ = ~new_n1724_ & new_n1727_;
  assign new_n1729_ = new_n1723_ & new_n1728_;
  assign new_n1730_ = new_n1716_ & new_n1729_;
  assign new_n1731_ = new_n1703_ & new_n1730_;
  assign new_n1732_ = new_n454_ & new_n1685_;
  assign new_n1733_ = new_n456_ & new_n1685_;
  assign new_n1734_ = ~new_n1732_ & ~new_n1733_;
  assign new_n1735_ = new_n545_ & new_n1571_;
  assign new_n1736_ = new_n543_ & new_n1735_;
  assign new_n1737_ = new_n553_ & new_n1735_;
  assign new_n1738_ = ~new_n1736_ & ~new_n1737_;
  assign new_n1739_ = new_n1734_ & new_n1738_;
  assign new_n1740_ = A167 & A168;
  assign new_n1741_ = A169 & new_n1740_;
  assign new_n1742_ = new_n193_ & new_n1741_;
  assign new_n1743_ = new_n319_ & new_n1742_;
  assign new_n1744_ = new_n323_ & new_n1742_;
  assign new_n1745_ = ~new_n1743_ & ~new_n1744_;
  assign new_n1746_ = new_n326_ & new_n1742_;
  assign new_n1747_ = new_n331_ & new_n1742_;
  assign new_n1748_ = ~new_n1746_ & ~new_n1747_;
  assign new_n1749_ = new_n1745_ & new_n1748_;
  assign new_n1750_ = new_n1739_ & new_n1749_;
  assign new_n1751_ = new_n334_ & new_n1742_;
  assign new_n1752_ = new_n338_ & new_n1742_;
  assign new_n1753_ = ~new_n1751_ & ~new_n1752_;
  assign new_n1754_ = new_n341_ & new_n1742_;
  assign new_n1755_ = new_n347_ & new_n1742_;
  assign new_n1756_ = ~new_n1754_ & ~new_n1755_;
  assign new_n1757_ = new_n1753_ & new_n1756_;
  assign new_n1758_ = new_n354_ & new_n1742_;
  assign new_n1759_ = new_n349_ & new_n1742_;
  assign new_n1760_ = new_n352_ & new_n1742_;
  assign new_n1761_ = ~new_n1759_ & ~new_n1760_;
  assign new_n1762_ = ~new_n1758_ & new_n1761_;
  assign new_n1763_ = new_n1757_ & new_n1762_;
  assign new_n1764_ = new_n1750_ & new_n1763_;
  assign new_n1765_ = new_n360_ & new_n1742_;
  assign new_n1766_ = new_n362_ & new_n1742_;
  assign new_n1767_ = ~new_n1765_ & ~new_n1766_;
  assign new_n1768_ = new_n358_ & new_n1742_;
  assign new_n1769_ = new_n368_ & new_n1742_;
  assign new_n1770_ = ~new_n1768_ & ~new_n1769_;
  assign new_n1771_ = new_n1767_ & new_n1770_;
  assign new_n1772_ = new_n219_ & new_n1741_;
  assign new_n1773_ = new_n377_ & new_n1772_;
  assign new_n1774_ = new_n370_ & new_n1742_;
  assign new_n1775_ = new_n374_ & new_n1772_;
  assign new_n1776_ = ~new_n1774_ & ~new_n1775_;
  assign new_n1777_ = ~new_n1773_ & new_n1776_;
  assign new_n1778_ = new_n1771_ & new_n1777_;
  assign new_n1779_ = new_n388_ & new_n1772_;
  assign new_n1780_ = new_n391_ & new_n1772_;
  assign new_n1781_ = ~new_n1779_ & ~new_n1780_;
  assign new_n1782_ = new_n385_ & new_n1772_;
  assign new_n1783_ = new_n398_ & new_n1772_;
  assign new_n1784_ = ~new_n1782_ & ~new_n1783_;
  assign new_n1785_ = new_n1781_ & new_n1784_;
  assign new_n1786_ = new_n405_ & new_n1772_;
  assign new_n1787_ = new_n400_ & new_n1772_;
  assign new_n1788_ = new_n403_ & new_n1772_;
  assign new_n1789_ = ~new_n1787_ & ~new_n1788_;
  assign new_n1790_ = ~new_n1786_ & new_n1789_;
  assign new_n1791_ = new_n1785_ & new_n1790_;
  assign new_n1792_ = new_n1778_ & new_n1791_;
  assign new_n1793_ = new_n1764_ & new_n1792_;
  assign new_n1794_ = new_n1731_ & new_n1793_;
  assign new_n1795_ = new_n1673_ & new_n1794_;
  assign new_n1796_ = new_n1545_ & new_n1795_;
  assign new_n1797_ = new_n413_ & new_n1772_;
  assign new_n1798_ = new_n415_ & new_n1772_;
  assign new_n1799_ = ~new_n1797_ & ~new_n1798_;
  assign new_n1800_ = new_n411_ & new_n1772_;
  assign new_n1801_ = new_n424_ & new_n1772_;
  assign new_n1802_ = ~new_n1800_ & ~new_n1801_;
  assign new_n1803_ = new_n1799_ & new_n1802_;
  assign new_n1804_ = new_n426_ & new_n1772_;
  assign new_n1805_ = new_n429_ & new_n1772_;
  assign new_n1806_ = ~new_n1804_ & ~new_n1805_;
  assign new_n1807_ = new_n431_ & new_n1772_;
  assign new_n1808_ = new_n436_ & new_n1772_;
  assign new_n1809_ = ~new_n1807_ & ~new_n1808_;
  assign new_n1810_ = new_n1806_ & new_n1809_;
  assign new_n1811_ = new_n1803_ & new_n1810_;
  assign new_n1812_ = new_n438_ & new_n1772_;
  assign new_n1813_ = new_n441_ & new_n1772_;
  assign new_n1814_ = ~new_n1812_ & ~new_n1813_;
  assign new_n1815_ = new_n443_ & new_n1772_;
  assign new_n1816_ = new_n448_ & new_n1772_;
  assign new_n1817_ = ~new_n1815_ & ~new_n1816_;
  assign new_n1818_ = new_n1814_ & new_n1817_;
  assign new_n1819_ = new_n456_ & new_n1772_;
  assign new_n1820_ = new_n450_ & new_n1772_;
  assign new_n1821_ = new_n454_ & new_n1772_;
  assign new_n1822_ = ~new_n1820_ & ~new_n1821_;
  assign new_n1823_ = ~new_n1819_ & new_n1822_;
  assign new_n1824_ = new_n1818_ & new_n1823_;
  assign new_n1825_ = new_n1811_ & new_n1824_;
  assign new_n1826_ = new_n227_ & new_n1741_;
  assign new_n1827_ = new_n319_ & new_n1826_;
  assign new_n1828_ = new_n323_ & new_n1826_;
  assign new_n1829_ = ~new_n1827_ & ~new_n1828_;
  assign new_n1830_ = new_n326_ & new_n1826_;
  assign new_n1831_ = new_n331_ & new_n1826_;
  assign new_n1832_ = ~new_n1830_ & ~new_n1831_;
  assign new_n1833_ = new_n1829_ & new_n1832_;
  assign new_n1834_ = new_n341_ & new_n1826_;
  assign new_n1835_ = new_n334_ & new_n1826_;
  assign new_n1836_ = new_n338_ & new_n1826_;
  assign new_n1837_ = ~new_n1835_ & ~new_n1836_;
  assign new_n1838_ = ~new_n1834_ & new_n1837_;
  assign new_n1839_ = new_n1833_ & new_n1838_;
  assign new_n1840_ = new_n347_ & new_n1826_;
  assign new_n1841_ = new_n349_ & new_n1826_;
  assign new_n1842_ = ~new_n1840_ & ~new_n1841_;
  assign new_n1843_ = new_n352_ & new_n1826_;
  assign new_n1844_ = new_n354_ & new_n1826_;
  assign new_n1845_ = ~new_n1843_ & ~new_n1844_;
  assign new_n1846_ = new_n1842_ & new_n1845_;
  assign new_n1847_ = new_n358_ & new_n1826_;
  assign new_n1848_ = new_n360_ & new_n1826_;
  assign new_n1849_ = new_n362_ & new_n1826_;
  assign new_n1850_ = ~new_n1848_ & ~new_n1849_;
  assign new_n1851_ = ~new_n1847_ & new_n1850_;
  assign new_n1852_ = new_n1846_ & new_n1851_;
  assign new_n1853_ = new_n1839_ & new_n1852_;
  assign new_n1854_ = new_n1825_ & new_n1853_;
  assign new_n1855_ = new_n368_ & new_n1826_;
  assign new_n1856_ = new_n370_ & new_n1826_;
  assign new_n1857_ = ~new_n1855_ & ~new_n1856_;
  assign new_n1858_ = new_n256_ & new_n1741_;
  assign new_n1859_ = new_n374_ & new_n1858_;
  assign new_n1860_ = new_n377_ & new_n1858_;
  assign new_n1861_ = ~new_n1859_ & ~new_n1860_;
  assign new_n1862_ = new_n1857_ & new_n1861_;
  assign new_n1863_ = new_n388_ & new_n1858_;
  assign new_n1864_ = new_n391_ & new_n1858_;
  assign new_n1865_ = ~new_n1863_ & ~new_n1864_;
  assign new_n1866_ = new_n385_ & new_n1858_;
  assign new_n1867_ = new_n398_ & new_n1858_;
  assign new_n1868_ = ~new_n1866_ & ~new_n1867_;
  assign new_n1869_ = new_n1865_ & new_n1868_;
  assign new_n1870_ = new_n1862_ & new_n1869_;
  assign new_n1871_ = new_n400_ & new_n1858_;
  assign new_n1872_ = new_n403_ & new_n1858_;
  assign new_n1873_ = ~new_n1871_ & ~new_n1872_;
  assign new_n1874_ = new_n405_ & new_n1858_;
  assign new_n1875_ = new_n413_ & new_n1858_;
  assign new_n1876_ = ~new_n1874_ & ~new_n1875_;
  assign new_n1877_ = new_n1873_ & new_n1876_;
  assign new_n1878_ = new_n424_ & new_n1858_;
  assign new_n1879_ = new_n415_ & new_n1858_;
  assign new_n1880_ = new_n411_ & new_n1858_;
  assign new_n1881_ = ~new_n1879_ & ~new_n1880_;
  assign new_n1882_ = ~new_n1878_ & new_n1881_;
  assign new_n1883_ = new_n1877_ & new_n1882_;
  assign new_n1884_ = new_n1870_ & new_n1883_;
  assign new_n1885_ = new_n426_ & new_n1858_;
  assign new_n1886_ = new_n429_ & new_n1858_;
  assign new_n1887_ = ~new_n1885_ & ~new_n1886_;
  assign new_n1888_ = new_n431_ & new_n1858_;
  assign new_n1889_ = new_n436_ & new_n1858_;
  assign new_n1890_ = ~new_n1888_ & ~new_n1889_;
  assign new_n1891_ = new_n1887_ & new_n1890_;
  assign new_n1892_ = new_n443_ & new_n1858_;
  assign new_n1893_ = new_n438_ & new_n1858_;
  assign new_n1894_ = new_n441_ & new_n1858_;
  assign new_n1895_ = ~new_n1893_ & ~new_n1894_;
  assign new_n1896_ = ~new_n1892_ & new_n1895_;
  assign new_n1897_ = new_n1891_ & new_n1896_;
  assign new_n1898_ = new_n448_ & new_n1858_;
  assign new_n1899_ = new_n450_ & new_n1858_;
  assign new_n1900_ = ~new_n1898_ & ~new_n1899_;
  assign new_n1901_ = new_n454_ & new_n1858_;
  assign new_n1902_ = new_n456_ & new_n1858_;
  assign new_n1903_ = ~new_n1901_ & ~new_n1902_;
  assign new_n1904_ = new_n1900_ & new_n1903_;
  assign new_n1905_ = ~A170 & new_n1556_;
  assign new_n1906_ = new_n723_ & new_n1905_;
  assign new_n1907_ = new_n543_ & new_n1906_;
  assign new_n1908_ = new_n718_ & new_n1741_;
  assign new_n1909_ = new_n543_ & new_n1908_;
  assign new_n1910_ = new_n553_ & new_n1908_;
  assign new_n1911_ = ~new_n1909_ & ~new_n1910_;
  assign new_n1912_ = ~new_n1907_ & new_n1911_;
  assign new_n1913_ = new_n1904_ & new_n1912_;
  assign new_n1914_ = new_n1897_ & new_n1913_;
  assign new_n1915_ = new_n1884_ & new_n1914_;
  assign new_n1916_ = new_n1854_ & new_n1915_;
  assign new_n1917_ = new_n553_ & new_n1906_;
  assign new_n1918_ = ~A170 & new_n1562_;
  assign new_n1919_ = new_n733_ & new_n1918_;
  assign new_n1920_ = new_n543_ & new_n1919_;
  assign new_n1921_ = ~new_n1917_ & ~new_n1920_;
  assign new_n1922_ = new_n553_ & new_n1919_;
  assign new_n1923_ = ~A170 & new_n1570_;
  assign new_n1924_ = new_n83_ & new_n1923_;
  assign new_n1925_ = new_n319_ & new_n1924_;
  assign new_n1926_ = ~new_n1922_ & ~new_n1925_;
  assign new_n1927_ = new_n1921_ & new_n1926_;
  assign new_n1928_ = new_n323_ & new_n1924_;
  assign new_n1929_ = new_n326_ & new_n1924_;
  assign new_n1930_ = ~new_n1928_ & ~new_n1929_;
  assign new_n1931_ = new_n331_ & new_n1924_;
  assign new_n1932_ = new_n334_ & new_n1924_;
  assign new_n1933_ = ~new_n1931_ & ~new_n1932_;
  assign new_n1934_ = new_n1930_ & new_n1933_;
  assign new_n1935_ = new_n1927_ & new_n1934_;
  assign new_n1936_ = new_n338_ & new_n1924_;
  assign new_n1937_ = new_n341_ & new_n1924_;
  assign new_n1938_ = ~new_n1936_ & ~new_n1937_;
  assign new_n1939_ = new_n347_ & new_n1924_;
  assign new_n1940_ = new_n349_ & new_n1924_;
  assign new_n1941_ = ~new_n1939_ & ~new_n1940_;
  assign new_n1942_ = new_n1938_ & new_n1941_;
  assign new_n1943_ = new_n360_ & new_n1924_;
  assign new_n1944_ = new_n352_ & new_n1924_;
  assign new_n1945_ = new_n354_ & new_n1924_;
  assign new_n1946_ = ~new_n1944_ & ~new_n1945_;
  assign new_n1947_ = ~new_n1943_ & new_n1946_;
  assign new_n1948_ = new_n1942_ & new_n1947_;
  assign new_n1949_ = new_n1935_ & new_n1948_;
  assign new_n1950_ = new_n362_ & new_n1924_;
  assign new_n1951_ = new_n358_ & new_n1924_;
  assign new_n1952_ = ~new_n1950_ & ~new_n1951_;
  assign new_n1953_ = new_n368_ & new_n1924_;
  assign new_n1954_ = new_n370_ & new_n1924_;
  assign new_n1955_ = ~new_n1953_ & ~new_n1954_;
  assign new_n1956_ = new_n1952_ & new_n1955_;
  assign new_n1957_ = new_n135_ & new_n1923_;
  assign new_n1958_ = new_n388_ & new_n1957_;
  assign new_n1959_ = new_n374_ & new_n1957_;
  assign new_n1960_ = new_n377_ & new_n1957_;
  assign new_n1961_ = ~new_n1959_ & ~new_n1960_;
  assign new_n1962_ = ~new_n1958_ & new_n1961_;
  assign new_n1963_ = new_n1956_ & new_n1962_;
  assign new_n1964_ = new_n391_ & new_n1957_;
  assign new_n1965_ = new_n385_ & new_n1957_;
  assign new_n1966_ = ~new_n1964_ & ~new_n1965_;
  assign new_n1967_ = new_n398_ & new_n1957_;
  assign new_n1968_ = new_n400_ & new_n1957_;
  assign new_n1969_ = ~new_n1967_ & ~new_n1968_;
  assign new_n1970_ = new_n1966_ & new_n1969_;
  assign new_n1971_ = new_n413_ & new_n1957_;
  assign new_n1972_ = new_n403_ & new_n1957_;
  assign new_n1973_ = new_n405_ & new_n1957_;
  assign new_n1974_ = ~new_n1972_ & ~new_n1973_;
  assign new_n1975_ = ~new_n1971_ & new_n1974_;
  assign new_n1976_ = new_n1970_ & new_n1975_;
  assign new_n1977_ = new_n1963_ & new_n1976_;
  assign new_n1978_ = new_n1949_ & new_n1977_;
  assign new_n1979_ = new_n415_ & new_n1957_;
  assign new_n1980_ = new_n411_ & new_n1957_;
  assign new_n1981_ = ~new_n1979_ & ~new_n1980_;
  assign new_n1982_ = new_n424_ & new_n1957_;
  assign new_n1983_ = new_n426_ & new_n1957_;
  assign new_n1984_ = ~new_n1982_ & ~new_n1983_;
  assign new_n1985_ = new_n1981_ & new_n1984_;
  assign new_n1986_ = new_n429_ & new_n1957_;
  assign new_n1987_ = new_n431_ & new_n1957_;
  assign new_n1988_ = ~new_n1986_ & ~new_n1987_;
  assign new_n1989_ = new_n436_ & new_n1957_;
  assign new_n1990_ = new_n438_ & new_n1957_;
  assign new_n1991_ = ~new_n1989_ & ~new_n1990_;
  assign new_n1992_ = new_n1988_ & new_n1991_;
  assign new_n1993_ = new_n1985_ & new_n1992_;
  assign new_n1994_ = new_n441_ & new_n1957_;
  assign new_n1995_ = new_n443_ & new_n1957_;
  assign new_n1996_ = ~new_n1994_ & ~new_n1995_;
  assign new_n1997_ = new_n448_ & new_n1957_;
  assign new_n1998_ = new_n450_ & new_n1957_;
  assign new_n1999_ = ~new_n1997_ & ~new_n1998_;
  assign new_n2000_ = new_n1996_ & new_n1999_;
  assign new_n2001_ = new_n157_ & new_n1923_;
  assign new_n2002_ = new_n319_ & new_n2001_;
  assign new_n2003_ = new_n454_ & new_n1957_;
  assign new_n2004_ = new_n456_ & new_n1957_;
  assign new_n2005_ = ~new_n2003_ & ~new_n2004_;
  assign new_n2006_ = ~new_n2002_ & new_n2005_;
  assign new_n2007_ = new_n2000_ & new_n2006_;
  assign new_n2008_ = new_n1993_ & new_n2007_;
  assign new_n2009_ = new_n323_ & new_n2001_;
  assign new_n2010_ = new_n326_ & new_n2001_;
  assign new_n2011_ = ~new_n2009_ & ~new_n2010_;
  assign new_n2012_ = new_n331_ & new_n2001_;
  assign new_n2013_ = new_n334_ & new_n2001_;
  assign new_n2014_ = ~new_n2012_ & ~new_n2013_;
  assign new_n2015_ = new_n2011_ & new_n2014_;
  assign new_n2016_ = new_n347_ & new_n2001_;
  assign new_n2017_ = new_n338_ & new_n2001_;
  assign new_n2018_ = new_n341_ & new_n2001_;
  assign new_n2019_ = ~new_n2017_ & ~new_n2018_;
  assign new_n2020_ = ~new_n2016_ & new_n2019_;
  assign new_n2021_ = new_n2015_ & new_n2020_;
  assign new_n2022_ = new_n349_ & new_n2001_;
  assign new_n2023_ = new_n352_ & new_n2001_;
  assign new_n2024_ = ~new_n2022_ & ~new_n2023_;
  assign new_n2025_ = new_n354_ & new_n2001_;
  assign new_n2026_ = new_n360_ & new_n2001_;
  assign new_n2027_ = ~new_n2025_ & ~new_n2026_;
  assign new_n2028_ = new_n2024_ & new_n2027_;
  assign new_n2029_ = new_n368_ & new_n2001_;
  assign new_n2030_ = new_n362_ & new_n2001_;
  assign new_n2031_ = new_n358_ & new_n2001_;
  assign new_n2032_ = ~new_n2030_ & ~new_n2031_;
  assign new_n2033_ = ~new_n2029_ & new_n2032_;
  assign new_n2034_ = new_n2028_ & new_n2033_;
  assign new_n2035_ = new_n2021_ & new_n2034_;
  assign new_n2036_ = new_n2008_ & new_n2035_;
  assign new_n2037_ = new_n1978_ & new_n2036_;
  assign new_n2038_ = new_n1916_ & new_n2037_;
  assign new_n2039_ = new_n370_ & new_n2001_;
  assign new_n2040_ = new_n183_ & new_n1923_;
  assign new_n2041_ = new_n374_ & new_n2040_;
  assign new_n2042_ = ~new_n2039_ & ~new_n2041_;
  assign new_n2043_ = new_n377_ & new_n2040_;
  assign new_n2044_ = new_n388_ & new_n2040_;
  assign new_n2045_ = ~new_n2043_ & ~new_n2044_;
  assign new_n2046_ = new_n2042_ & new_n2045_;
  assign new_n2047_ = new_n391_ & new_n2040_;
  assign new_n2048_ = new_n385_ & new_n2040_;
  assign new_n2049_ = ~new_n2047_ & ~new_n2048_;
  assign new_n2050_ = new_n398_ & new_n2040_;
  assign new_n2051_ = new_n400_ & new_n2040_;
  assign new_n2052_ = ~new_n2050_ & ~new_n2051_;
  assign new_n2053_ = new_n2049_ & new_n2052_;
  assign new_n2054_ = new_n2046_ & new_n2053_;
  assign new_n2055_ = new_n403_ & new_n2040_;
  assign new_n2056_ = new_n405_ & new_n2040_;
  assign new_n2057_ = ~new_n2055_ & ~new_n2056_;
  assign new_n2058_ = new_n413_ & new_n2040_;
  assign new_n2059_ = new_n415_ & new_n2040_;
  assign new_n2060_ = ~new_n2058_ & ~new_n2059_;
  assign new_n2061_ = new_n2057_ & new_n2060_;
  assign new_n2062_ = new_n426_ & new_n2040_;
  assign new_n2063_ = new_n411_ & new_n2040_;
  assign new_n2064_ = new_n424_ & new_n2040_;
  assign new_n2065_ = ~new_n2063_ & ~new_n2064_;
  assign new_n2066_ = ~new_n2062_ & new_n2065_;
  assign new_n2067_ = new_n2061_ & new_n2066_;
  assign new_n2068_ = new_n2054_ & new_n2067_;
  assign new_n2069_ = new_n429_ & new_n2040_;
  assign new_n2070_ = new_n431_ & new_n2040_;
  assign new_n2071_ = ~new_n2069_ & ~new_n2070_;
  assign new_n2072_ = new_n436_ & new_n2040_;
  assign new_n2073_ = new_n438_ & new_n2040_;
  assign new_n2074_ = ~new_n2072_ & ~new_n2073_;
  assign new_n2075_ = new_n2071_ & new_n2074_;
  assign new_n2076_ = new_n448_ & new_n2040_;
  assign new_n2077_ = new_n441_ & new_n2040_;
  assign new_n2078_ = new_n443_ & new_n2040_;
  assign new_n2079_ = ~new_n2077_ & ~new_n2078_;
  assign new_n2080_ = ~new_n2076_ & new_n2079_;
  assign new_n2081_ = new_n2075_ & new_n2080_;
  assign new_n2082_ = new_n450_ & new_n2040_;
  assign new_n2083_ = new_n454_ & new_n2040_;
  assign new_n2084_ = ~new_n2082_ & ~new_n2083_;
  assign new_n2085_ = new_n456_ & new_n2040_;
  assign new_n2086_ = new_n545_ & new_n1923_;
  assign new_n2087_ = new_n543_ & new_n2086_;
  assign new_n2088_ = ~new_n2085_ & ~new_n2087_;
  assign new_n2089_ = new_n2084_ & new_n2088_;
  assign new_n2090_ = ~A170 & new_n1740_;
  assign new_n2091_ = new_n193_ & new_n2090_;
  assign new_n2092_ = new_n323_ & new_n2091_;
  assign new_n2093_ = new_n553_ & new_n2086_;
  assign new_n2094_ = new_n319_ & new_n2091_;
  assign new_n2095_ = ~new_n2093_ & ~new_n2094_;
  assign new_n2096_ = ~new_n2092_ & new_n2095_;
  assign new_n2097_ = new_n2089_ & new_n2096_;
  assign new_n2098_ = new_n2081_ & new_n2097_;
  assign new_n2099_ = new_n2068_ & new_n2098_;
  assign new_n2100_ = new_n326_ & new_n2091_;
  assign new_n2101_ = new_n331_ & new_n2091_;
  assign new_n2102_ = ~new_n2100_ & ~new_n2101_;
  assign new_n2103_ = new_n334_ & new_n2091_;
  assign new_n2104_ = new_n338_ & new_n2091_;
  assign new_n2105_ = ~new_n2103_ & ~new_n2104_;
  assign new_n2106_ = new_n2102_ & new_n2105_;
  assign new_n2107_ = new_n341_ & new_n2091_;
  assign new_n2108_ = new_n347_ & new_n2091_;
  assign new_n2109_ = ~new_n2107_ & ~new_n2108_;
  assign new_n2110_ = new_n349_ & new_n2091_;
  assign new_n2111_ = new_n352_ & new_n2091_;
  assign new_n2112_ = ~new_n2110_ & ~new_n2111_;
  assign new_n2113_ = new_n2109_ & new_n2112_;
  assign new_n2114_ = new_n2106_ & new_n2113_;
  assign new_n2115_ = new_n354_ & new_n2091_;
  assign new_n2116_ = new_n360_ & new_n2091_;
  assign new_n2117_ = ~new_n2115_ & ~new_n2116_;
  assign new_n2118_ = new_n362_ & new_n2091_;
  assign new_n2119_ = new_n358_ & new_n2091_;
  assign new_n2120_ = ~new_n2118_ & ~new_n2119_;
  assign new_n2121_ = new_n2117_ & new_n2120_;
  assign new_n2122_ = new_n219_ & new_n2090_;
  assign new_n2123_ = new_n374_ & new_n2122_;
  assign new_n2124_ = new_n368_ & new_n2091_;
  assign new_n2125_ = new_n370_ & new_n2091_;
  assign new_n2126_ = ~new_n2124_ & ~new_n2125_;
  assign new_n2127_ = ~new_n2123_ & new_n2126_;
  assign new_n2128_ = new_n2121_ & new_n2127_;
  assign new_n2129_ = new_n2114_ & new_n2128_;
  assign new_n2130_ = new_n377_ & new_n2122_;
  assign new_n2131_ = new_n388_ & new_n2122_;
  assign new_n2132_ = ~new_n2130_ & ~new_n2131_;
  assign new_n2133_ = new_n391_ & new_n2122_;
  assign new_n2134_ = new_n385_ & new_n2122_;
  assign new_n2135_ = ~new_n2133_ & ~new_n2134_;
  assign new_n2136_ = new_n2132_ & new_n2135_;
  assign new_n2137_ = new_n403_ & new_n2122_;
  assign new_n2138_ = new_n398_ & new_n2122_;
  assign new_n2139_ = new_n400_ & new_n2122_;
  assign new_n2140_ = ~new_n2138_ & ~new_n2139_;
  assign new_n2141_ = ~new_n2137_ & new_n2140_;
  assign new_n2142_ = new_n2136_ & new_n2141_;
  assign new_n2143_ = new_n405_ & new_n2122_;
  assign new_n2144_ = new_n413_ & new_n2122_;
  assign new_n2145_ = ~new_n2143_ & ~new_n2144_;
  assign new_n2146_ = new_n415_ & new_n2122_;
  assign new_n2147_ = new_n411_ & new_n2122_;
  assign new_n2148_ = ~new_n2146_ & ~new_n2147_;
  assign new_n2149_ = new_n2145_ & new_n2148_;
  assign new_n2150_ = new_n429_ & new_n2122_;
  assign new_n2151_ = new_n424_ & new_n2122_;
  assign new_n2152_ = new_n426_ & new_n2122_;
  assign new_n2153_ = ~new_n2151_ & ~new_n2152_;
  assign new_n2154_ = ~new_n2150_ & new_n2153_;
  assign new_n2155_ = new_n2149_ & new_n2154_;
  assign new_n2156_ = new_n2142_ & new_n2155_;
  assign new_n2157_ = new_n2129_ & new_n2156_;
  assign new_n2158_ = new_n2099_ & new_n2157_;
  assign new_n2159_ = new_n431_ & new_n2122_;
  assign new_n2160_ = new_n436_ & new_n2122_;
  assign new_n2161_ = ~new_n2159_ & ~new_n2160_;
  assign new_n2162_ = new_n438_ & new_n2122_;
  assign new_n2163_ = new_n441_ & new_n2122_;
  assign new_n2164_ = ~new_n2162_ & ~new_n2163_;
  assign new_n2165_ = new_n2161_ & new_n2164_;
  assign new_n2166_ = new_n443_ & new_n2122_;
  assign new_n2167_ = new_n448_ & new_n2122_;
  assign new_n2168_ = ~new_n2166_ & ~new_n2167_;
  assign new_n2169_ = new_n450_ & new_n2122_;
  assign new_n2170_ = new_n454_ & new_n2122_;
  assign new_n2171_ = ~new_n2169_ & ~new_n2170_;
  assign new_n2172_ = new_n2168_ & new_n2171_;
  assign new_n2173_ = new_n2165_ & new_n2172_;
  assign new_n2174_ = new_n456_ & new_n2122_;
  assign new_n2175_ = new_n227_ & new_n2090_;
  assign new_n2176_ = new_n319_ & new_n2175_;
  assign new_n2177_ = ~new_n2174_ & ~new_n2176_;
  assign new_n2178_ = new_n323_ & new_n2175_;
  assign new_n2179_ = new_n326_ & new_n2175_;
  assign new_n2180_ = ~new_n2178_ & ~new_n2179_;
  assign new_n2181_ = new_n2177_ & new_n2180_;
  assign new_n2182_ = new_n338_ & new_n2175_;
  assign new_n2183_ = new_n331_ & new_n2175_;
  assign new_n2184_ = new_n334_ & new_n2175_;
  assign new_n2185_ = ~new_n2183_ & ~new_n2184_;
  assign new_n2186_ = ~new_n2182_ & new_n2185_;
  assign new_n2187_ = new_n2181_ & new_n2186_;
  assign new_n2188_ = new_n2173_ & new_n2187_;
  assign new_n2189_ = new_n341_ & new_n2175_;
  assign new_n2190_ = new_n347_ & new_n2175_;
  assign new_n2191_ = ~new_n2189_ & ~new_n2190_;
  assign new_n2192_ = new_n349_ & new_n2175_;
  assign new_n2193_ = new_n352_ & new_n2175_;
  assign new_n2194_ = ~new_n2192_ & ~new_n2193_;
  assign new_n2195_ = new_n2191_ & new_n2194_;
  assign new_n2196_ = new_n362_ & new_n2175_;
  assign new_n2197_ = new_n354_ & new_n2175_;
  assign new_n2198_ = new_n360_ & new_n2175_;
  assign new_n2199_ = ~new_n2197_ & ~new_n2198_;
  assign new_n2200_ = ~new_n2196_ & new_n2199_;
  assign new_n2201_ = new_n2195_ & new_n2200_;
  assign new_n2202_ = new_n358_ & new_n2175_;
  assign new_n2203_ = new_n368_ & new_n2175_;
  assign new_n2204_ = ~new_n2202_ & ~new_n2203_;
  assign new_n2205_ = new_n370_ & new_n2175_;
  assign new_n2206_ = new_n256_ & new_n2090_;
  assign new_n2207_ = new_n374_ & new_n2206_;
  assign new_n2208_ = ~new_n2205_ & ~new_n2207_;
  assign new_n2209_ = new_n2204_ & new_n2208_;
  assign new_n2210_ = new_n391_ & new_n2206_;
  assign new_n2211_ = new_n377_ & new_n2206_;
  assign new_n2212_ = new_n388_ & new_n2206_;
  assign new_n2213_ = ~new_n2211_ & ~new_n2212_;
  assign new_n2214_ = ~new_n2210_ & new_n2213_;
  assign new_n2215_ = new_n2209_ & new_n2214_;
  assign new_n2216_ = new_n2201_ & new_n2215_;
  assign new_n2217_ = new_n2188_ & new_n2216_;
  assign new_n2218_ = new_n385_ & new_n2206_;
  assign new_n2219_ = new_n398_ & new_n2206_;
  assign new_n2220_ = ~new_n2218_ & ~new_n2219_;
  assign new_n2221_ = new_n400_ & new_n2206_;
  assign new_n2222_ = new_n403_ & new_n2206_;
  assign new_n2223_ = ~new_n2221_ & ~new_n2222_;
  assign new_n2224_ = new_n2220_ & new_n2223_;
  assign new_n2225_ = new_n415_ & new_n2206_;
  assign new_n2226_ = new_n405_ & new_n2206_;
  assign new_n2227_ = new_n413_ & new_n2206_;
  assign new_n2228_ = ~new_n2226_ & ~new_n2227_;
  assign new_n2229_ = ~new_n2225_ & new_n2228_;
  assign new_n2230_ = new_n2224_ & new_n2229_;
  assign new_n2231_ = new_n411_ & new_n2206_;
  assign new_n2232_ = new_n424_ & new_n2206_;
  assign new_n2233_ = ~new_n2231_ & ~new_n2232_;
  assign new_n2234_ = new_n426_ & new_n2206_;
  assign new_n2235_ = new_n429_ & new_n2206_;
  assign new_n2236_ = ~new_n2234_ & ~new_n2235_;
  assign new_n2237_ = new_n2233_ & new_n2236_;
  assign new_n2238_ = new_n438_ & new_n2206_;
  assign new_n2239_ = new_n431_ & new_n2206_;
  assign new_n2240_ = new_n436_ & new_n2206_;
  assign new_n2241_ = ~new_n2239_ & ~new_n2240_;
  assign new_n2242_ = ~new_n2238_ & new_n2241_;
  assign new_n2243_ = new_n2237_ & new_n2242_;
  assign new_n2244_ = new_n2230_ & new_n2243_;
  assign new_n2245_ = new_n441_ & new_n2206_;
  assign new_n2246_ = new_n443_ & new_n2206_;
  assign new_n2247_ = ~new_n2245_ & ~new_n2246_;
  assign new_n2248_ = new_n448_ & new_n2206_;
  assign new_n2249_ = new_n450_ & new_n2206_;
  assign new_n2250_ = ~new_n2248_ & ~new_n2249_;
  assign new_n2251_ = new_n2247_ & new_n2250_;
  assign new_n2252_ = new_n718_ & new_n2090_;
  assign new_n2253_ = new_n543_ & new_n2252_;
  assign new_n2254_ = new_n454_ & new_n2206_;
  assign new_n2255_ = new_n456_ & new_n2206_;
  assign new_n2256_ = ~new_n2254_ & ~new_n2255_;
  assign new_n2257_ = ~new_n2253_ & new_n2256_;
  assign new_n2258_ = new_n2251_ & new_n2257_;
  assign new_n2259_ = new_n553_ & new_n2252_;
  assign new_n2260_ = ~A167 & new_n58_;
  assign new_n2261_ = new_n723_ & new_n2260_;
  assign new_n2262_ = new_n543_ & new_n2261_;
  assign new_n2263_ = ~new_n2259_ & ~new_n2262_;
  assign new_n2264_ = new_n553_ & new_n2261_;
  assign new_n2265_ = ~A167 & new_n66_;
  assign new_n2266_ = new_n733_ & new_n2265_;
  assign new_n2267_ = new_n543_ & new_n2266_;
  assign new_n2268_ = ~new_n2264_ & ~new_n2267_;
  assign new_n2269_ = new_n2263_ & new_n2268_;
  assign new_n2270_ = A167 & new_n37_;
  assign new_n2271_ = new_n723_ & new_n2270_;
  assign new_n2272_ = new_n553_ & new_n2271_;
  assign new_n2273_ = new_n553_ & new_n2266_;
  assign new_n2274_ = new_n543_ & new_n2271_;
  assign new_n2275_ = ~new_n2273_ & ~new_n2274_;
  assign new_n2276_ = ~new_n2272_ & new_n2275_;
  assign new_n2277_ = new_n2269_ & new_n2276_;
  assign new_n2278_ = new_n2258_ & new_n2277_;
  assign new_n2279_ = new_n2244_ & new_n2278_;
  assign new_n2280_ = new_n2217_ & new_n2279_;
  assign new_n2281_ = new_n2158_ & new_n2280_;
  assign new_n2282_ = new_n2038_ & new_n2281_;
  assign new_n2283_ = new_n1796_ & new_n2282_;
  assign new_n2284_ = new_n1277_ & new_n2283_;
  assign new_n2285_ = A167 & new_n51_;
  assign new_n2286_ = new_n733_ & new_n2285_;
  assign new_n2287_ = new_n543_ & new_n2286_;
  assign new_n2288_ = new_n553_ & new_n2286_;
  assign new_n2289_ = ~new_n2287_ & ~new_n2288_;
  assign new_n2290_ = ~A265 & new_n1234_;
  assign new_n2291_ = new_n539_ & new_n2290_;
  assign new_n2292_ = new_n1040_ & new_n2291_;
  assign new_n2293_ = ~A265 & new_n1241_;
  assign new_n2294_ = new_n550_ & new_n2293_;
  assign new_n2295_ = new_n1040_ & new_n2294_;
  assign new_n2296_ = ~new_n2292_ & ~new_n2295_;
  assign new_n2297_ = new_n2289_ & new_n2296_;
  assign new_n2298_ = A265 & new_n1246_;
  assign new_n2299_ = new_n539_ & new_n2298_;
  assign new_n2300_ = new_n1040_ & new_n2299_;
  assign new_n2301_ = A265 & new_n1250_;
  assign new_n2302_ = new_n550_ & new_n2301_;
  assign new_n2303_ = new_n1040_ & new_n2302_;
  assign new_n2304_ = ~new_n2300_ & ~new_n2303_;
  assign new_n2305_ = ~A267 & new_n1261_;
  assign new_n2306_ = new_n539_ & new_n2305_;
  assign new_n2307_ = new_n1040_ & new_n2306_;
  assign new_n2308_ = ~A267 & new_n1265_;
  assign new_n2309_ = new_n550_ & new_n2308_;
  assign new_n2310_ = new_n1040_ & new_n2309_;
  assign new_n2311_ = ~new_n2307_ & ~new_n2310_;
  assign new_n2312_ = new_n2304_ & new_n2311_;
  assign new_n2313_ = new_n2297_ & new_n2312_;
  assign new_n2314_ = ~A267 & new_n1256_;
  assign new_n2315_ = new_n539_ & new_n2314_;
  assign new_n2316_ = new_n1040_ & new_n2315_;
  assign new_n2317_ = ~A267 & new_n1278_;
  assign new_n2318_ = new_n550_ & new_n2317_;
  assign new_n2319_ = new_n1040_ & new_n2318_;
  assign new_n2320_ = ~new_n2316_ & ~new_n2319_;
  assign new_n2321_ = A267 & new_n29_;
  assign new_n2322_ = new_n1284_ & new_n2321_;
  assign new_n2323_ = new_n1040_ & new_n2322_;
  assign new_n2324_ = new_n1291_ & new_n2321_;
  assign new_n2325_ = new_n1040_ & new_n2324_;
  assign new_n2326_ = ~new_n2323_ & ~new_n2325_;
  assign new_n2327_ = new_n2320_ & new_n2326_;
  assign new_n2328_ = new_n1215_ & new_n2291_;
  assign new_n2329_ = new_n1295_ & new_n2321_;
  assign new_n2330_ = new_n1040_ & new_n2329_;
  assign new_n2331_ = new_n1300_ & new_n2321_;
  assign new_n2332_ = new_n1040_ & new_n2331_;
  assign new_n2333_ = ~new_n2330_ & ~new_n2332_;
  assign new_n2334_ = ~new_n2328_ & new_n2333_;
  assign new_n2335_ = new_n2327_ & new_n2334_;
  assign new_n2336_ = new_n2313_ & new_n2335_;
  assign new_n2337_ = new_n1215_ & new_n2294_;
  assign new_n2338_ = new_n1215_ & new_n2299_;
  assign new_n2339_ = ~new_n2337_ & ~new_n2338_;
  assign new_n2340_ = new_n1215_ & new_n2302_;
  assign new_n2341_ = new_n1215_ & new_n2306_;
  assign new_n2342_ = ~new_n2340_ & ~new_n2341_;
  assign new_n2343_ = new_n2339_ & new_n2342_;
  assign new_n2344_ = new_n1215_ & new_n2318_;
  assign new_n2345_ = new_n1215_ & new_n2309_;
  assign new_n2346_ = new_n1215_ & new_n2315_;
  assign new_n2347_ = ~new_n2345_ & ~new_n2346_;
  assign new_n2348_ = ~new_n2344_ & new_n2347_;
  assign new_n2349_ = new_n2343_ & new_n2348_;
  assign new_n2350_ = new_n1215_ & new_n2322_;
  assign new_n2351_ = new_n1215_ & new_n2324_;
  assign new_n2352_ = ~new_n2350_ & ~new_n2351_;
  assign new_n2353_ = new_n1215_ & new_n2329_;
  assign new_n2354_ = new_n1215_ & new_n2331_;
  assign new_n2355_ = ~new_n2353_ & ~new_n2354_;
  assign new_n2356_ = new_n2352_ & new_n2355_;
  assign new_n2357_ = new_n1221_ & new_n2299_;
  assign new_n2358_ = new_n1221_ & new_n2291_;
  assign new_n2359_ = new_n1221_ & new_n2294_;
  assign new_n2360_ = ~new_n2358_ & ~new_n2359_;
  assign new_n2361_ = ~new_n2357_ & new_n2360_;
  assign new_n2362_ = new_n2356_ & new_n2361_;
  assign new_n2363_ = new_n2349_ & new_n2362_;
  assign new_n2364_ = new_n2336_ & new_n2363_;
  assign new_n2365_ = new_n1221_ & new_n2302_;
  assign new_n2366_ = new_n1221_ & new_n2306_;
  assign new_n2367_ = ~new_n2365_ & ~new_n2366_;
  assign new_n2368_ = new_n1221_ & new_n2309_;
  assign new_n2369_ = new_n1221_ & new_n2315_;
  assign new_n2370_ = ~new_n2368_ & ~new_n2369_;
  assign new_n2371_ = new_n2367_ & new_n2370_;
  assign new_n2372_ = new_n1221_ & new_n2318_;
  assign new_n2373_ = new_n1221_ & new_n2322_;
  assign new_n2374_ = ~new_n2372_ & ~new_n2373_;
  assign new_n2375_ = new_n1221_ & new_n2324_;
  assign new_n2376_ = new_n1221_ & new_n2329_;
  assign new_n2377_ = ~new_n2375_ & ~new_n2376_;
  assign new_n2378_ = new_n2374_ & new_n2377_;
  assign new_n2379_ = new_n2371_ & new_n2378_;
  assign new_n2380_ = new_n1221_ & new_n2331_;
  assign new_n2381_ = new_n1227_ & new_n2291_;
  assign new_n2382_ = ~new_n2380_ & ~new_n2381_;
  assign new_n2383_ = new_n1227_ & new_n2294_;
  assign new_n2384_ = new_n1227_ & new_n2299_;
  assign new_n2385_ = ~new_n2383_ & ~new_n2384_;
  assign new_n2386_ = new_n2382_ & new_n2385_;
  assign new_n2387_ = new_n1227_ & new_n2309_;
  assign new_n2388_ = new_n1227_ & new_n2302_;
  assign new_n2389_ = new_n1227_ & new_n2306_;
  assign new_n2390_ = ~new_n2388_ & ~new_n2389_;
  assign new_n2391_ = ~new_n2387_ & new_n2390_;
  assign new_n2392_ = new_n2386_ & new_n2391_;
  assign new_n2393_ = new_n2379_ & new_n2392_;
  assign new_n2394_ = new_n1227_ & new_n2315_;
  assign new_n2395_ = new_n1227_ & new_n2318_;
  assign new_n2396_ = ~new_n2394_ & ~new_n2395_;
  assign new_n2397_ = new_n1227_ & new_n2322_;
  assign new_n2398_ = new_n1227_ & new_n2324_;
  assign new_n2399_ = ~new_n2397_ & ~new_n2398_;
  assign new_n2400_ = new_n2396_ & new_n2399_;
  assign new_n2401_ = ~A266 & ~A265;
  assign new_n2402_ = ~A203 & new_n2401_;
  assign new_n2403_ = new_n1284_ & new_n2402_;
  assign new_n2404_ = new_n1239_ & new_n2403_;
  assign new_n2405_ = new_n1227_ & new_n2329_;
  assign new_n2406_ = new_n1227_ & new_n2331_;
  assign new_n2407_ = ~new_n2405_ & ~new_n2406_;
  assign new_n2408_ = ~new_n2404_ & new_n2407_;
  assign new_n2409_ = new_n2400_ & new_n2408_;
  assign new_n2410_ = new_n1291_ & new_n2402_;
  assign new_n2411_ = new_n1239_ & new_n2410_;
  assign new_n2412_ = new_n1295_ & new_n2402_;
  assign new_n2413_ = new_n1239_ & new_n2412_;
  assign new_n2414_ = ~new_n2411_ & ~new_n2413_;
  assign new_n2415_ = new_n1300_ & new_n2402_;
  assign new_n2416_ = new_n1239_ & new_n2415_;
  assign new_n2417_ = A266 & A265;
  assign new_n2418_ = ~A203 & new_n2417_;
  assign new_n2419_ = new_n1284_ & new_n2418_;
  assign new_n2420_ = new_n1239_ & new_n2419_;
  assign new_n2421_ = ~new_n2416_ & ~new_n2420_;
  assign new_n2422_ = new_n2414_ & new_n2421_;
  assign new_n2423_ = new_n1300_ & new_n2418_;
  assign new_n2424_ = new_n1239_ & new_n2423_;
  assign new_n2425_ = new_n1291_ & new_n2418_;
  assign new_n2426_ = new_n1239_ & new_n2425_;
  assign new_n2427_ = new_n1295_ & new_n2418_;
  assign new_n2428_ = new_n1239_ & new_n2427_;
  assign new_n2429_ = ~new_n2426_ & ~new_n2428_;
  assign new_n2430_ = ~new_n2424_ & new_n2429_;
  assign new_n2431_ = new_n2422_ & new_n2430_;
  assign new_n2432_ = new_n2409_ & new_n2431_;
  assign new_n2433_ = new_n2393_ & new_n2432_;
  assign new_n2434_ = new_n2364_ & new_n2433_;
  assign new_n2435_ = A269 & ~A267;
  assign new_n2436_ = ~A203 & new_n2435_;
  assign new_n2437_ = new_n1284_ & new_n2436_;
  assign new_n2438_ = new_n1239_ & new_n2437_;
  assign new_n2439_ = new_n1291_ & new_n2436_;
  assign new_n2440_ = new_n1239_ & new_n2439_;
  assign new_n2441_ = ~new_n2438_ & ~new_n2440_;
  assign new_n2442_ = new_n1295_ & new_n2436_;
  assign new_n2443_ = new_n1239_ & new_n2442_;
  assign new_n2444_ = new_n1300_ & new_n2436_;
  assign new_n2445_ = new_n1239_ & new_n2444_;
  assign new_n2446_ = ~new_n2443_ & ~new_n2445_;
  assign new_n2447_ = new_n2441_ & new_n2446_;
  assign new_n2448_ = A268 & ~A267;
  assign new_n2449_ = ~A203 & new_n2448_;
  assign new_n2450_ = new_n1284_ & new_n2449_;
  assign new_n2451_ = new_n1239_ & new_n2450_;
  assign new_n2452_ = new_n1291_ & new_n2449_;
  assign new_n2453_ = new_n1239_ & new_n2452_;
  assign new_n2454_ = ~new_n2451_ & ~new_n2453_;
  assign new_n2455_ = new_n1295_ & new_n2449_;
  assign new_n2456_ = new_n1239_ & new_n2455_;
  assign new_n2457_ = new_n1300_ & new_n2449_;
  assign new_n2458_ = new_n1239_ & new_n2457_;
  assign new_n2459_ = ~new_n2456_ & ~new_n2458_;
  assign new_n2460_ = new_n2454_ & new_n2459_;
  assign new_n2461_ = new_n2447_ & new_n2460_;
  assign new_n2462_ = new_n1304_ & new_n2291_;
  assign new_n2463_ = new_n1304_ & new_n2294_;
  assign new_n2464_ = ~new_n2462_ & ~new_n2463_;
  assign new_n2465_ = new_n1304_ & new_n2299_;
  assign new_n2466_ = new_n1304_ & new_n2302_;
  assign new_n2467_ = ~new_n2465_ & ~new_n2466_;
  assign new_n2468_ = new_n2464_ & new_n2467_;
  assign new_n2469_ = new_n1304_ & new_n2315_;
  assign new_n2470_ = new_n1304_ & new_n2306_;
  assign new_n2471_ = new_n1304_ & new_n2309_;
  assign new_n2472_ = ~new_n2470_ & ~new_n2471_;
  assign new_n2473_ = ~new_n2469_ & new_n2472_;
  assign new_n2474_ = new_n2468_ & new_n2473_;
  assign new_n2475_ = new_n2461_ & new_n2474_;
  assign new_n2476_ = new_n1304_ & new_n2318_;
  assign new_n2477_ = new_n1304_ & new_n2322_;
  assign new_n2478_ = ~new_n2476_ & ~new_n2477_;
  assign new_n2479_ = new_n1304_ & new_n2324_;
  assign new_n2480_ = new_n1304_ & new_n2329_;
  assign new_n2481_ = ~new_n2479_ & ~new_n2480_;
  assign new_n2482_ = new_n2478_ & new_n2481_;
  assign new_n2483_ = new_n1439_ & new_n2294_;
  assign new_n2484_ = new_n1304_ & new_n2331_;
  assign new_n2485_ = new_n1439_ & new_n2291_;
  assign new_n2486_ = ~new_n2484_ & ~new_n2485_;
  assign new_n2487_ = ~new_n2483_ & new_n2486_;
  assign new_n2488_ = new_n2482_ & new_n2487_;
  assign new_n2489_ = new_n1439_ & new_n2299_;
  assign new_n2490_ = new_n1439_ & new_n2302_;
  assign new_n2491_ = ~new_n2489_ & ~new_n2490_;
  assign new_n2492_ = new_n1439_ & new_n2306_;
  assign new_n2493_ = new_n1439_ & new_n2309_;
  assign new_n2494_ = ~new_n2492_ & ~new_n2493_;
  assign new_n2495_ = new_n2491_ & new_n2494_;
  assign new_n2496_ = new_n1439_ & new_n2322_;
  assign new_n2497_ = new_n1439_ & new_n2315_;
  assign new_n2498_ = new_n1439_ & new_n2318_;
  assign new_n2499_ = ~new_n2497_ & ~new_n2498_;
  assign new_n2500_ = ~new_n2496_ & new_n2499_;
  assign new_n2501_ = new_n2495_ & new_n2500_;
  assign new_n2502_ = new_n2488_ & new_n2501_;
  assign new_n2503_ = new_n2475_ & new_n2502_;
  assign new_n2504_ = new_n1439_ & new_n2324_;
  assign new_n2505_ = new_n1439_ & new_n2329_;
  assign new_n2506_ = ~new_n2504_ & ~new_n2505_;
  assign new_n2507_ = new_n1439_ & new_n2331_;
  assign new_n2508_ = new_n1448_ & new_n2291_;
  assign new_n2509_ = ~new_n2507_ & ~new_n2508_;
  assign new_n2510_ = new_n2506_ & new_n2509_;
  assign new_n2511_ = new_n1448_ & new_n2294_;
  assign new_n2512_ = new_n1448_ & new_n2299_;
  assign new_n2513_ = ~new_n2511_ & ~new_n2512_;
  assign new_n2514_ = new_n1448_ & new_n2302_;
  assign new_n2515_ = new_n1448_ & new_n2306_;
  assign new_n2516_ = ~new_n2514_ & ~new_n2515_;
  assign new_n2517_ = new_n2513_ & new_n2516_;
  assign new_n2518_ = new_n2510_ & new_n2517_;
  assign new_n2519_ = new_n1448_ & new_n2309_;
  assign new_n2520_ = new_n1448_ & new_n2315_;
  assign new_n2521_ = ~new_n2519_ & ~new_n2520_;
  assign new_n2522_ = new_n1448_ & new_n2318_;
  assign new_n2523_ = new_n1448_ & new_n2322_;
  assign new_n2524_ = ~new_n2522_ & ~new_n2523_;
  assign new_n2525_ = new_n2521_ & new_n2524_;
  assign new_n2526_ = new_n1448_ & new_n2331_;
  assign new_n2527_ = new_n1448_ & new_n2324_;
  assign new_n2528_ = new_n1448_ & new_n2329_;
  assign new_n2529_ = ~new_n2527_ & ~new_n2528_;
  assign new_n2530_ = ~new_n2526_ & new_n2529_;
  assign new_n2531_ = new_n2525_ & new_n2530_;
  assign new_n2532_ = new_n2518_ & new_n2531_;
  assign new_n2533_ = new_n1453_ & new_n2291_;
  assign new_n2534_ = new_n1453_ & new_n2294_;
  assign new_n2535_ = ~new_n2533_ & ~new_n2534_;
  assign new_n2536_ = new_n1453_ & new_n2299_;
  assign new_n2537_ = new_n1453_ & new_n2302_;
  assign new_n2538_ = ~new_n2536_ & ~new_n2537_;
  assign new_n2539_ = new_n2535_ & new_n2538_;
  assign new_n2540_ = new_n1453_ & new_n2315_;
  assign new_n2541_ = new_n1453_ & new_n2306_;
  assign new_n2542_ = new_n1453_ & new_n2309_;
  assign new_n2543_ = ~new_n2541_ & ~new_n2542_;
  assign new_n2544_ = ~new_n2540_ & new_n2543_;
  assign new_n2545_ = new_n2539_ & new_n2544_;
  assign new_n2546_ = new_n1453_ & new_n2318_;
  assign new_n2547_ = new_n1453_ & new_n2322_;
  assign new_n2548_ = ~new_n2546_ & ~new_n2547_;
  assign new_n2549_ = new_n1453_ & new_n2324_;
  assign new_n2550_ = new_n1453_ & new_n2329_;
  assign new_n2551_ = ~new_n2549_ & ~new_n2550_;
  assign new_n2552_ = new_n2548_ & new_n2551_;
  assign new_n2553_ = new_n1459_ & new_n2410_;
  assign new_n2554_ = new_n1453_ & new_n2331_;
  assign new_n2555_ = new_n1459_ & new_n2403_;
  assign new_n2556_ = ~new_n2554_ & ~new_n2555_;
  assign new_n2557_ = ~new_n2553_ & new_n2556_;
  assign new_n2558_ = new_n2552_ & new_n2557_;
  assign new_n2559_ = new_n2545_ & new_n2558_;
  assign new_n2560_ = new_n2532_ & new_n2559_;
  assign new_n2561_ = new_n2503_ & new_n2560_;
  assign new_n2562_ = new_n2434_ & new_n2561_;
  assign new_n2563_ = new_n1459_ & new_n2412_;
  assign new_n2564_ = new_n1459_ & new_n2415_;
  assign new_n2565_ = ~new_n2563_ & ~new_n2564_;
  assign new_n2566_ = new_n1459_ & new_n2419_;
  assign new_n2567_ = new_n1459_ & new_n2425_;
  assign new_n2568_ = ~new_n2566_ & ~new_n2567_;
  assign new_n2569_ = new_n2565_ & new_n2568_;
  assign new_n2570_ = new_n1459_ & new_n2427_;
  assign new_n2571_ = new_n1459_ & new_n2423_;
  assign new_n2572_ = ~new_n2570_ & ~new_n2571_;
  assign new_n2573_ = new_n1459_ & new_n2437_;
  assign new_n2574_ = new_n1459_ & new_n2439_;
  assign new_n2575_ = ~new_n2573_ & ~new_n2574_;
  assign new_n2576_ = new_n2572_ & new_n2575_;
  assign new_n2577_ = new_n2569_ & new_n2576_;
  assign new_n2578_ = new_n1459_ & new_n2442_;
  assign new_n2579_ = new_n1459_ & new_n2444_;
  assign new_n2580_ = ~new_n2578_ & ~new_n2579_;
  assign new_n2581_ = new_n1459_ & new_n2450_;
  assign new_n2582_ = new_n1459_ & new_n2452_;
  assign new_n2583_ = ~new_n2581_ & ~new_n2582_;
  assign new_n2584_ = new_n2580_ & new_n2583_;
  assign new_n2585_ = new_n1486_ & new_n2403_;
  assign new_n2586_ = new_n1459_ & new_n2455_;
  assign new_n2587_ = new_n1459_ & new_n2457_;
  assign new_n2588_ = ~new_n2586_ & ~new_n2587_;
  assign new_n2589_ = ~new_n2585_ & new_n2588_;
  assign new_n2590_ = new_n2584_ & new_n2589_;
  assign new_n2591_ = new_n2577_ & new_n2590_;
  assign new_n2592_ = new_n1486_ & new_n2410_;
  assign new_n2593_ = new_n1486_ & new_n2412_;
  assign new_n2594_ = ~new_n2592_ & ~new_n2593_;
  assign new_n2595_ = new_n1486_ & new_n2415_;
  assign new_n2596_ = new_n1486_ & new_n2419_;
  assign new_n2597_ = ~new_n2595_ & ~new_n2596_;
  assign new_n2598_ = new_n2594_ & new_n2597_;
  assign new_n2599_ = new_n1486_ & new_n2423_;
  assign new_n2600_ = new_n1486_ & new_n2425_;
  assign new_n2601_ = new_n1486_ & new_n2427_;
  assign new_n2602_ = ~new_n2600_ & ~new_n2601_;
  assign new_n2603_ = ~new_n2599_ & new_n2602_;
  assign new_n2604_ = new_n2598_ & new_n2603_;
  assign new_n2605_ = new_n1486_ & new_n2437_;
  assign new_n2606_ = new_n1486_ & new_n2439_;
  assign new_n2607_ = ~new_n2605_ & ~new_n2606_;
  assign new_n2608_ = new_n1486_ & new_n2442_;
  assign new_n2609_ = new_n1486_ & new_n2444_;
  assign new_n2610_ = ~new_n2608_ & ~new_n2609_;
  assign new_n2611_ = new_n2607_ & new_n2610_;
  assign new_n2612_ = new_n1486_ & new_n2455_;
  assign new_n2613_ = new_n1486_ & new_n2450_;
  assign new_n2614_ = new_n1486_ & new_n2452_;
  assign new_n2615_ = ~new_n2613_ & ~new_n2614_;
  assign new_n2616_ = ~new_n2612_ & new_n2615_;
  assign new_n2617_ = new_n2611_ & new_n2616_;
  assign new_n2618_ = new_n2604_ & new_n2617_;
  assign new_n2619_ = new_n2591_ & new_n2618_;
  assign new_n2620_ = new_n1486_ & new_n2457_;
  assign new_n2621_ = new_n1506_ & new_n2291_;
  assign new_n2622_ = ~new_n2620_ & ~new_n2621_;
  assign new_n2623_ = new_n1506_ & new_n2294_;
  assign new_n2624_ = new_n1506_ & new_n2299_;
  assign new_n2625_ = ~new_n2623_ & ~new_n2624_;
  assign new_n2626_ = new_n2622_ & new_n2625_;
  assign new_n2627_ = new_n1506_ & new_n2302_;
  assign new_n2628_ = new_n1506_ & new_n2306_;
  assign new_n2629_ = ~new_n2627_ & ~new_n2628_;
  assign new_n2630_ = new_n1506_ & new_n2309_;
  assign new_n2631_ = new_n1506_ & new_n2315_;
  assign new_n2632_ = ~new_n2630_ & ~new_n2631_;
  assign new_n2633_ = new_n2629_ & new_n2632_;
  assign new_n2634_ = new_n2626_ & new_n2633_;
  assign new_n2635_ = new_n1506_ & new_n2318_;
  assign new_n2636_ = new_n1506_ & new_n2322_;
  assign new_n2637_ = ~new_n2635_ & ~new_n2636_;
  assign new_n2638_ = new_n1506_ & new_n2324_;
  assign new_n2639_ = new_n1506_ & new_n2329_;
  assign new_n2640_ = ~new_n2638_ & ~new_n2639_;
  assign new_n2641_ = new_n2637_ & new_n2640_;
  assign new_n2642_ = new_n1515_ & new_n2294_;
  assign new_n2643_ = new_n1506_ & new_n2331_;
  assign new_n2644_ = new_n1515_ & new_n2291_;
  assign new_n2645_ = ~new_n2643_ & ~new_n2644_;
  assign new_n2646_ = ~new_n2642_ & new_n2645_;
  assign new_n2647_ = new_n2641_ & new_n2646_;
  assign new_n2648_ = new_n2634_ & new_n2647_;
  assign new_n2649_ = new_n1515_ & new_n2299_;
  assign new_n2650_ = new_n1515_ & new_n2302_;
  assign new_n2651_ = ~new_n2649_ & ~new_n2650_;
  assign new_n2652_ = new_n1515_ & new_n2306_;
  assign new_n2653_ = new_n1515_ & new_n2309_;
  assign new_n2654_ = ~new_n2652_ & ~new_n2653_;
  assign new_n2655_ = new_n2651_ & new_n2654_;
  assign new_n2656_ = new_n1515_ & new_n2322_;
  assign new_n2657_ = new_n1515_ & new_n2315_;
  assign new_n2658_ = new_n1515_ & new_n2318_;
  assign new_n2659_ = ~new_n2657_ & ~new_n2658_;
  assign new_n2660_ = ~new_n2656_ & new_n2659_;
  assign new_n2661_ = new_n2655_ & new_n2660_;
  assign new_n2662_ = new_n1515_ & new_n2324_;
  assign new_n2663_ = new_n1515_ & new_n2329_;
  assign new_n2664_ = ~new_n2662_ & ~new_n2663_;
  assign new_n2665_ = new_n1515_ & new_n2331_;
  assign new_n2666_ = new_n1519_ & new_n2403_;
  assign new_n2667_ = ~new_n2665_ & ~new_n2666_;
  assign new_n2668_ = new_n2664_ & new_n2667_;
  assign new_n2669_ = new_n1519_ & new_n2415_;
  assign new_n2670_ = new_n1519_ & new_n2410_;
  assign new_n2671_ = new_n1519_ & new_n2412_;
  assign new_n2672_ = ~new_n2670_ & ~new_n2671_;
  assign new_n2673_ = ~new_n2669_ & new_n2672_;
  assign new_n2674_ = new_n2668_ & new_n2673_;
  assign new_n2675_ = new_n2661_ & new_n2674_;
  assign new_n2676_ = new_n2648_ & new_n2675_;
  assign new_n2677_ = new_n2619_ & new_n2676_;
  assign new_n2678_ = new_n1519_ & new_n2419_;
  assign new_n2679_ = new_n1519_ & new_n2425_;
  assign new_n2680_ = ~new_n2678_ & ~new_n2679_;
  assign new_n2681_ = new_n1519_ & new_n2427_;
  assign new_n2682_ = new_n1519_ & new_n2423_;
  assign new_n2683_ = ~new_n2681_ & ~new_n2682_;
  assign new_n2684_ = new_n2680_ & new_n2683_;
  assign new_n2685_ = new_n1519_ & new_n2437_;
  assign new_n2686_ = new_n1519_ & new_n2439_;
  assign new_n2687_ = ~new_n2685_ & ~new_n2686_;
  assign new_n2688_ = new_n1519_ & new_n2442_;
  assign new_n2689_ = new_n1519_ & new_n2444_;
  assign new_n2690_ = ~new_n2688_ & ~new_n2689_;
  assign new_n2691_ = new_n2687_ & new_n2690_;
  assign new_n2692_ = new_n2684_ & new_n2691_;
  assign new_n2693_ = new_n1519_ & new_n2450_;
  assign new_n2694_ = new_n1519_ & new_n2452_;
  assign new_n2695_ = ~new_n2693_ & ~new_n2694_;
  assign new_n2696_ = new_n1519_ & new_n2455_;
  assign new_n2697_ = new_n1519_ & new_n2457_;
  assign new_n2698_ = ~new_n2696_ & ~new_n2697_;
  assign new_n2699_ = new_n2695_ & new_n2698_;
  assign new_n2700_ = new_n1547_ & new_n2299_;
  assign new_n2701_ = new_n1547_ & new_n2291_;
  assign new_n2702_ = new_n1547_ & new_n2294_;
  assign new_n2703_ = ~new_n2701_ & ~new_n2702_;
  assign new_n2704_ = ~new_n2700_ & new_n2703_;
  assign new_n2705_ = new_n2699_ & new_n2704_;
  assign new_n2706_ = new_n2692_ & new_n2705_;
  assign new_n2707_ = new_n1547_ & new_n2302_;
  assign new_n2708_ = new_n1547_ & new_n2306_;
  assign new_n2709_ = ~new_n2707_ & ~new_n2708_;
  assign new_n2710_ = new_n1547_ & new_n2309_;
  assign new_n2711_ = new_n1547_ & new_n2315_;
  assign new_n2712_ = ~new_n2710_ & ~new_n2711_;
  assign new_n2713_ = new_n2709_ & new_n2712_;
  assign new_n2714_ = new_n1547_ & new_n2324_;
  assign new_n2715_ = new_n1547_ & new_n2318_;
  assign new_n2716_ = new_n1547_ & new_n2322_;
  assign new_n2717_ = ~new_n2715_ & ~new_n2716_;
  assign new_n2718_ = ~new_n2714_ & new_n2717_;
  assign new_n2719_ = new_n2713_ & new_n2718_;
  assign new_n2720_ = new_n1547_ & new_n2329_;
  assign new_n2721_ = new_n1547_ & new_n2331_;
  assign new_n2722_ = ~new_n2720_ & ~new_n2721_;
  assign new_n2723_ = new_n1551_ & new_n2291_;
  assign new_n2724_ = new_n1551_ & new_n2294_;
  assign new_n2725_ = ~new_n2723_ & ~new_n2724_;
  assign new_n2726_ = new_n2722_ & new_n2725_;
  assign new_n2727_ = new_n1551_ & new_n2306_;
  assign new_n2728_ = new_n1551_ & new_n2299_;
  assign new_n2729_ = new_n1551_ & new_n2302_;
  assign new_n2730_ = ~new_n2728_ & ~new_n2729_;
  assign new_n2731_ = ~new_n2727_ & new_n2730_;
  assign new_n2732_ = new_n2726_ & new_n2731_;
  assign new_n2733_ = new_n2719_ & new_n2732_;
  assign new_n2734_ = new_n2706_ & new_n2733_;
  assign new_n2735_ = new_n1551_ & new_n2309_;
  assign new_n2736_ = new_n1551_ & new_n2315_;
  assign new_n2737_ = ~new_n2735_ & ~new_n2736_;
  assign new_n2738_ = new_n1551_ & new_n2318_;
  assign new_n2739_ = new_n1551_ & new_n2322_;
  assign new_n2740_ = ~new_n2738_ & ~new_n2739_;
  assign new_n2741_ = new_n2737_ & new_n2740_;
  assign new_n2742_ = new_n1551_ & new_n2324_;
  assign new_n2743_ = new_n1551_ & new_n2329_;
  assign new_n2744_ = ~new_n2742_ & ~new_n2743_;
  assign new_n2745_ = new_n1551_ & new_n2331_;
  assign new_n2746_ = ~A266 & new_n76_;
  assign new_n2747_ = new_n778_ & new_n2746_;
  assign new_n2748_ = new_n32_ & new_n1237_;
  assign new_n2749_ = new_n1485_ & new_n2748_;
  assign new_n2750_ = new_n2747_ & new_n2749_;
  assign new_n2751_ = ~new_n2745_ & ~new_n2750_;
  assign new_n2752_ = new_n2744_ & new_n2751_;
  assign new_n2753_ = new_n2741_ & new_n2752_;
  assign new_n2754_ = A266 & new_n76_;
  assign new_n2755_ = new_n778_ & new_n2754_;
  assign new_n2756_ = new_n45_ & new_n1237_;
  assign new_n2757_ = new_n1485_ & new_n2756_;
  assign new_n2758_ = new_n2755_ & new_n2757_;
  assign new_n2759_ = new_n1558_ & new_n2291_;
  assign new_n2760_ = ~new_n2758_ & ~new_n2759_;
  assign new_n2761_ = new_n1558_ & new_n2294_;
  assign new_n2762_ = new_n1558_ & new_n2299_;
  assign new_n2763_ = ~new_n2761_ & ~new_n2762_;
  assign new_n2764_ = new_n2760_ & new_n2763_;
  assign new_n2765_ = new_n1558_ & new_n2309_;
  assign new_n2766_ = new_n1558_ & new_n2302_;
  assign new_n2767_ = new_n1558_ & new_n2306_;
  assign new_n2768_ = ~new_n2766_ & ~new_n2767_;
  assign new_n2769_ = ~new_n2765_ & new_n2768_;
  assign new_n2770_ = new_n2764_ & new_n2769_;
  assign new_n2771_ = new_n2753_ & new_n2770_;
  assign new_n2772_ = new_n1558_ & new_n2315_;
  assign new_n2773_ = new_n1558_ & new_n2318_;
  assign new_n2774_ = ~new_n2772_ & ~new_n2773_;
  assign new_n2775_ = new_n1558_ & new_n2322_;
  assign new_n2776_ = new_n1558_ & new_n2324_;
  assign new_n2777_ = ~new_n2775_ & ~new_n2776_;
  assign new_n2778_ = new_n2774_ & new_n2777_;
  assign new_n2779_ = ~A268 & new_n540_;
  assign new_n2780_ = new_n539_ & new_n2779_;
  assign new_n2781_ = A267 & A203;
  assign new_n2782_ = new_n134_ & new_n2781_;
  assign new_n2783_ = new_n1557_ & new_n2782_;
  assign new_n2784_ = new_n2780_ & new_n2783_;
  assign new_n2785_ = new_n1558_ & new_n2329_;
  assign new_n2786_ = new_n1558_ & new_n2331_;
  assign new_n2787_ = ~new_n2785_ & ~new_n2786_;
  assign new_n2788_ = ~new_n2784_ & new_n2787_;
  assign new_n2789_ = new_n2778_ & new_n2788_;
  assign new_n2790_ = ~A268 & new_n551_;
  assign new_n2791_ = new_n550_ & new_n2790_;
  assign new_n2792_ = new_n2783_ & new_n2791_;
  assign new_n2793_ = A267 & A202;
  assign new_n2794_ = new_n134_ & new_n2793_;
  assign new_n2795_ = new_n1557_ & new_n2794_;
  assign new_n2796_ = new_n2780_ & new_n2795_;
  assign new_n2797_ = ~new_n2792_ & ~new_n2796_;
  assign new_n2798_ = new_n2791_ & new_n2795_;
  assign new_n2799_ = new_n1564_ & new_n2291_;
  assign new_n2800_ = ~new_n2798_ & ~new_n2799_;
  assign new_n2801_ = new_n2797_ & new_n2800_;
  assign new_n2802_ = new_n1564_ & new_n2302_;
  assign new_n2803_ = new_n1564_ & new_n2294_;
  assign new_n2804_ = new_n1564_ & new_n2299_;
  assign new_n2805_ = ~new_n2803_ & ~new_n2804_;
  assign new_n2806_ = ~new_n2802_ & new_n2805_;
  assign new_n2807_ = new_n2801_ & new_n2806_;
  assign new_n2808_ = new_n2789_ & new_n2807_;
  assign new_n2809_ = new_n2771_ & new_n2808_;
  assign new_n2810_ = new_n2734_ & new_n2809_;
  assign new_n2811_ = new_n2677_ & new_n2810_;
  assign new_n2812_ = new_n2562_ & new_n2811_;
  assign new_n2813_ = new_n1564_ & new_n2306_;
  assign new_n2814_ = new_n1564_ & new_n2309_;
  assign new_n2815_ = ~new_n2813_ & ~new_n2814_;
  assign new_n2816_ = new_n1564_ & new_n2315_;
  assign new_n2817_ = new_n1564_ & new_n2318_;
  assign new_n2818_ = ~new_n2816_ & ~new_n2817_;
  assign new_n2819_ = new_n2815_ & new_n2818_;
  assign new_n2820_ = new_n1564_ & new_n2322_;
  assign new_n2821_ = new_n1564_ & new_n2324_;
  assign new_n2822_ = ~new_n2820_ & ~new_n2821_;
  assign new_n2823_ = new_n1564_ & new_n2329_;
  assign new_n2824_ = new_n1564_ & new_n2331_;
  assign new_n2825_ = ~new_n2823_ & ~new_n2824_;
  assign new_n2826_ = new_n2822_ & new_n2825_;
  assign new_n2827_ = new_n2819_ & new_n2826_;
  assign new_n2828_ = new_n182_ & new_n2781_;
  assign new_n2829_ = new_n1563_ & new_n2828_;
  assign new_n2830_ = new_n2780_ & new_n2829_;
  assign new_n2831_ = new_n2791_ & new_n2829_;
  assign new_n2832_ = ~new_n2830_ & ~new_n2831_;
  assign new_n2833_ = new_n182_ & new_n2793_;
  assign new_n2834_ = new_n1563_ & new_n2833_;
  assign new_n2835_ = new_n2780_ & new_n2834_;
  assign new_n2836_ = new_n2791_ & new_n2834_;
  assign new_n2837_ = ~new_n2835_ & ~new_n2836_;
  assign new_n2838_ = new_n2832_ & new_n2837_;
  assign new_n2839_ = A203 & new_n78_;
  assign new_n2840_ = new_n318_ & new_n2839_;
  assign new_n2841_ = new_n1603_ & new_n2840_;
  assign new_n2842_ = A267 & ~A200;
  assign new_n2843_ = new_n51_ & new_n2842_;
  assign new_n2844_ = new_n1571_ & new_n2843_;
  assign new_n2845_ = new_n2780_ & new_n2844_;
  assign new_n2846_ = new_n2791_ & new_n2844_;
  assign new_n2847_ = ~new_n2845_ & ~new_n2846_;
  assign new_n2848_ = ~new_n2841_ & new_n2847_;
  assign new_n2849_ = new_n2838_ & new_n2848_;
  assign new_n2850_ = new_n2827_ & new_n2849_;
  assign new_n2851_ = new_n322_ & new_n2839_;
  assign new_n2852_ = new_n1603_ & new_n2851_;
  assign new_n2853_ = new_n325_ & new_n2839_;
  assign new_n2854_ = new_n1603_ & new_n2853_;
  assign new_n2855_ = ~new_n2852_ & ~new_n2854_;
  assign new_n2856_ = new_n330_ & new_n2839_;
  assign new_n2857_ = new_n1603_ & new_n2856_;
  assign new_n2858_ = new_n333_ & new_n2839_;
  assign new_n2859_ = new_n1603_ & new_n2858_;
  assign new_n2860_ = ~new_n2857_ & ~new_n2859_;
  assign new_n2861_ = new_n2855_ & new_n2860_;
  assign new_n2862_ = new_n346_ & new_n2839_;
  assign new_n2863_ = new_n1603_ & new_n2862_;
  assign new_n2864_ = new_n337_ & new_n2839_;
  assign new_n2865_ = new_n1603_ & new_n2864_;
  assign new_n2866_ = new_n340_ & new_n2839_;
  assign new_n2867_ = new_n1603_ & new_n2866_;
  assign new_n2868_ = ~new_n2865_ & ~new_n2867_;
  assign new_n2869_ = ~new_n2863_ & new_n2868_;
  assign new_n2870_ = new_n2861_ & new_n2869_;
  assign new_n2871_ = A203 & new_n104_;
  assign new_n2872_ = new_n318_ & new_n2871_;
  assign new_n2873_ = new_n1603_ & new_n2872_;
  assign new_n2874_ = new_n322_ & new_n2871_;
  assign new_n2875_ = new_n1603_ & new_n2874_;
  assign new_n2876_ = ~new_n2873_ & ~new_n2875_;
  assign new_n2877_ = new_n325_ & new_n2871_;
  assign new_n2878_ = new_n1603_ & new_n2877_;
  assign new_n2879_ = new_n330_ & new_n2871_;
  assign new_n2880_ = new_n1603_ & new_n2879_;
  assign new_n2881_ = ~new_n2878_ & ~new_n2880_;
  assign new_n2882_ = new_n2876_ & new_n2881_;
  assign new_n2883_ = new_n340_ & new_n2871_;
  assign new_n2884_ = new_n1603_ & new_n2883_;
  assign new_n2885_ = new_n333_ & new_n2871_;
  assign new_n2886_ = new_n1603_ & new_n2885_;
  assign new_n2887_ = new_n337_ & new_n2871_;
  assign new_n2888_ = new_n1603_ & new_n2887_;
  assign new_n2889_ = ~new_n2886_ & ~new_n2888_;
  assign new_n2890_ = ~new_n2884_ & new_n2889_;
  assign new_n2891_ = new_n2882_ & new_n2890_;
  assign new_n2892_ = new_n2870_ & new_n2891_;
  assign new_n2893_ = new_n2850_ & new_n2892_;
  assign new_n2894_ = new_n346_ & new_n2871_;
  assign new_n2895_ = new_n1603_ & new_n2894_;
  assign new_n2896_ = A202 & new_n78_;
  assign new_n2897_ = new_n318_ & new_n2896_;
  assign new_n2898_ = new_n1603_ & new_n2897_;
  assign new_n2899_ = ~new_n2895_ & ~new_n2898_;
  assign new_n2900_ = new_n322_ & new_n2896_;
  assign new_n2901_ = new_n1603_ & new_n2900_;
  assign new_n2902_ = new_n325_ & new_n2896_;
  assign new_n2903_ = new_n1603_ & new_n2902_;
  assign new_n2904_ = ~new_n2901_ & ~new_n2903_;
  assign new_n2905_ = new_n2899_ & new_n2904_;
  assign new_n2906_ = new_n330_ & new_n2896_;
  assign new_n2907_ = new_n1603_ & new_n2906_;
  assign new_n2908_ = new_n333_ & new_n2896_;
  assign new_n2909_ = new_n1603_ & new_n2908_;
  assign new_n2910_ = ~new_n2907_ & ~new_n2909_;
  assign new_n2911_ = new_n337_ & new_n2896_;
  assign new_n2912_ = new_n1603_ & new_n2911_;
  assign new_n2913_ = new_n340_ & new_n2896_;
  assign new_n2914_ = new_n1603_ & new_n2913_;
  assign new_n2915_ = ~new_n2912_ & ~new_n2914_;
  assign new_n2916_ = new_n2910_ & new_n2915_;
  assign new_n2917_ = new_n2905_ & new_n2916_;
  assign new_n2918_ = new_n346_ & new_n2896_;
  assign new_n2919_ = new_n1603_ & new_n2918_;
  assign new_n2920_ = A202 & new_n104_;
  assign new_n2921_ = new_n318_ & new_n2920_;
  assign new_n2922_ = new_n1603_ & new_n2921_;
  assign new_n2923_ = ~new_n2919_ & ~new_n2922_;
  assign new_n2924_ = new_n322_ & new_n2920_;
  assign new_n2925_ = new_n1603_ & new_n2924_;
  assign new_n2926_ = new_n325_ & new_n2920_;
  assign new_n2927_ = new_n1603_ & new_n2926_;
  assign new_n2928_ = ~new_n2925_ & ~new_n2927_;
  assign new_n2929_ = new_n2923_ & new_n2928_;
  assign new_n2930_ = new_n337_ & new_n2920_;
  assign new_n2931_ = new_n1603_ & new_n2930_;
  assign new_n2932_ = new_n330_ & new_n2920_;
  assign new_n2933_ = new_n1603_ & new_n2932_;
  assign new_n2934_ = new_n333_ & new_n2920_;
  assign new_n2935_ = new_n1603_ & new_n2934_;
  assign new_n2936_ = ~new_n2933_ & ~new_n2935_;
  assign new_n2937_ = ~new_n2931_ & new_n2936_;
  assign new_n2938_ = new_n2929_ & new_n2937_;
  assign new_n2939_ = new_n2917_ & new_n2938_;
  assign new_n2940_ = new_n340_ & new_n2920_;
  assign new_n2941_ = new_n1603_ & new_n2940_;
  assign new_n2942_ = new_n346_ & new_n2920_;
  assign new_n2943_ = new_n1603_ & new_n2942_;
  assign new_n2944_ = ~new_n2941_ & ~new_n2943_;
  assign new_n2945_ = new_n1685_ & new_n2840_;
  assign new_n2946_ = new_n1685_ & new_n2851_;
  assign new_n2947_ = ~new_n2945_ & ~new_n2946_;
  assign new_n2948_ = new_n2944_ & new_n2947_;
  assign new_n2949_ = new_n1685_ & new_n2858_;
  assign new_n2950_ = new_n1685_ & new_n2853_;
  assign new_n2951_ = new_n1685_ & new_n2856_;
  assign new_n2952_ = ~new_n2950_ & ~new_n2951_;
  assign new_n2953_ = ~new_n2949_ & new_n2952_;
  assign new_n2954_ = new_n2948_ & new_n2953_;
  assign new_n2955_ = new_n1685_ & new_n2864_;
  assign new_n2956_ = new_n1685_ & new_n2866_;
  assign new_n2957_ = ~new_n2955_ & ~new_n2956_;
  assign new_n2958_ = new_n1685_ & new_n2862_;
  assign new_n2959_ = new_n1685_ & new_n2872_;
  assign new_n2960_ = ~new_n2958_ & ~new_n2959_;
  assign new_n2961_ = new_n2957_ & new_n2960_;
  assign new_n2962_ = new_n1685_ & new_n2879_;
  assign new_n2963_ = new_n1685_ & new_n2874_;
  assign new_n2964_ = new_n1685_ & new_n2877_;
  assign new_n2965_ = ~new_n2963_ & ~new_n2964_;
  assign new_n2966_ = ~new_n2962_ & new_n2965_;
  assign new_n2967_ = new_n2961_ & new_n2966_;
  assign new_n2968_ = new_n2954_ & new_n2967_;
  assign new_n2969_ = new_n2939_ & new_n2968_;
  assign new_n2970_ = new_n2893_ & new_n2969_;
  assign new_n2971_ = new_n1685_ & new_n2885_;
  assign new_n2972_ = new_n1685_ & new_n2887_;
  assign new_n2973_ = ~new_n2971_ & ~new_n2972_;
  assign new_n2974_ = new_n1685_ & new_n2883_;
  assign new_n2975_ = new_n1685_ & new_n2894_;
  assign new_n2976_ = ~new_n2974_ & ~new_n2975_;
  assign new_n2977_ = new_n2973_ & new_n2976_;
  assign new_n2978_ = new_n1685_ & new_n2897_;
  assign new_n2979_ = new_n1685_ & new_n2900_;
  assign new_n2980_ = ~new_n2978_ & ~new_n2979_;
  assign new_n2981_ = new_n1685_ & new_n2902_;
  assign new_n2982_ = new_n1685_ & new_n2906_;
  assign new_n2983_ = ~new_n2981_ & ~new_n2982_;
  assign new_n2984_ = new_n2980_ & new_n2983_;
  assign new_n2985_ = new_n2977_ & new_n2984_;
  assign new_n2986_ = new_n1685_ & new_n2908_;
  assign new_n2987_ = new_n1685_ & new_n2911_;
  assign new_n2988_ = ~new_n2986_ & ~new_n2987_;
  assign new_n2989_ = new_n1685_ & new_n2913_;
  assign new_n2990_ = new_n1685_ & new_n2918_;
  assign new_n2991_ = ~new_n2989_ & ~new_n2990_;
  assign new_n2992_ = new_n2988_ & new_n2991_;
  assign new_n2993_ = new_n1685_ & new_n2926_;
  assign new_n2994_ = new_n1685_ & new_n2921_;
  assign new_n2995_ = new_n1685_ & new_n2924_;
  assign new_n2996_ = ~new_n2994_ & ~new_n2995_;
  assign new_n2997_ = ~new_n2993_ & new_n2996_;
  assign new_n2998_ = new_n2992_ & new_n2997_;
  assign new_n2999_ = new_n2985_ & new_n2998_;
  assign new_n3000_ = new_n1685_ & new_n2932_;
  assign new_n3001_ = new_n1685_ & new_n2934_;
  assign new_n3002_ = ~new_n3000_ & ~new_n3001_;
  assign new_n3003_ = new_n1685_ & new_n2930_;
  assign new_n3004_ = new_n1685_ & new_n2940_;
  assign new_n3005_ = ~new_n3003_ & ~new_n3004_;
  assign new_n3006_ = new_n3002_ & new_n3005_;
  assign new_n3007_ = A267 & A200;
  assign new_n3008_ = new_n37_ & new_n3007_;
  assign new_n3009_ = new_n1571_ & new_n3008_;
  assign new_n3010_ = new_n2791_ & new_n3009_;
  assign new_n3011_ = new_n1685_ & new_n2942_;
  assign new_n3012_ = new_n2780_ & new_n3009_;
  assign new_n3013_ = ~new_n3011_ & ~new_n3012_;
  assign new_n3014_ = ~new_n3010_ & new_n3013_;
  assign new_n3015_ = new_n3006_ & new_n3014_;
  assign new_n3016_ = ~A201 & A166;
  assign new_n3017_ = new_n2781_ & new_n3016_;
  assign new_n3018_ = new_n1571_ & new_n3017_;
  assign new_n3019_ = new_n2780_ & new_n3018_;
  assign new_n3020_ = new_n2791_ & new_n3018_;
  assign new_n3021_ = ~new_n3019_ & ~new_n3020_;
  assign new_n3022_ = new_n2793_ & new_n3016_;
  assign new_n3023_ = new_n1571_ & new_n3022_;
  assign new_n3024_ = new_n2780_ & new_n3023_;
  assign new_n3025_ = new_n2791_ & new_n3023_;
  assign new_n3026_ = ~new_n3024_ & ~new_n3025_;
  assign new_n3027_ = new_n3021_ & new_n3026_;
  assign new_n3028_ = new_n1735_ & new_n2299_;
  assign new_n3029_ = new_n1735_ & new_n2291_;
  assign new_n3030_ = new_n1735_ & new_n2294_;
  assign new_n3031_ = ~new_n3029_ & ~new_n3030_;
  assign new_n3032_ = ~new_n3028_ & new_n3031_;
  assign new_n3033_ = new_n3027_ & new_n3032_;
  assign new_n3034_ = new_n3015_ & new_n3033_;
  assign new_n3035_ = new_n2999_ & new_n3034_;
  assign new_n3036_ = new_n1735_ & new_n2302_;
  assign new_n3037_ = new_n1735_ & new_n2306_;
  assign new_n3038_ = ~new_n3036_ & ~new_n3037_;
  assign new_n3039_ = new_n1735_ & new_n2309_;
  assign new_n3040_ = new_n1735_ & new_n2315_;
  assign new_n3041_ = ~new_n3039_ & ~new_n3040_;
  assign new_n3042_ = new_n3038_ & new_n3041_;
  assign new_n3043_ = new_n1735_ & new_n2318_;
  assign new_n3044_ = new_n1735_ & new_n2322_;
  assign new_n3045_ = ~new_n3043_ & ~new_n3044_;
  assign new_n3046_ = new_n1735_ & new_n2324_;
  assign new_n3047_ = new_n1735_ & new_n2329_;
  assign new_n3048_ = ~new_n3046_ & ~new_n3047_;
  assign new_n3049_ = new_n3045_ & new_n3048_;
  assign new_n3050_ = new_n3042_ & new_n3049_;
  assign new_n3051_ = new_n1735_ & new_n2331_;
  assign new_n3052_ = new_n66_ & new_n2842_;
  assign new_n3053_ = new_n1741_ & new_n3052_;
  assign new_n3054_ = new_n2780_ & new_n3053_;
  assign new_n3055_ = ~new_n3051_ & ~new_n3054_;
  assign new_n3056_ = new_n2791_ & new_n3053_;
  assign new_n3057_ = new_n1772_ & new_n2840_;
  assign new_n3058_ = ~new_n3056_ & ~new_n3057_;
  assign new_n3059_ = new_n3055_ & new_n3058_;
  assign new_n3060_ = new_n1772_ & new_n2856_;
  assign new_n3061_ = new_n1772_ & new_n2851_;
  assign new_n3062_ = new_n1772_ & new_n2853_;
  assign new_n3063_ = ~new_n3061_ & ~new_n3062_;
  assign new_n3064_ = ~new_n3060_ & new_n3063_;
  assign new_n3065_ = new_n3059_ & new_n3064_;
  assign new_n3066_ = new_n3050_ & new_n3065_;
  assign new_n3067_ = new_n1772_ & new_n2858_;
  assign new_n3068_ = new_n1772_ & new_n2864_;
  assign new_n3069_ = ~new_n3067_ & ~new_n3068_;
  assign new_n3070_ = new_n1772_ & new_n2866_;
  assign new_n3071_ = new_n1772_ & new_n2862_;
  assign new_n3072_ = ~new_n3070_ & ~new_n3071_;
  assign new_n3073_ = new_n3069_ & new_n3072_;
  assign new_n3074_ = new_n1772_ & new_n2877_;
  assign new_n3075_ = new_n1772_ & new_n2872_;
  assign new_n3076_ = new_n1772_ & new_n2874_;
  assign new_n3077_ = ~new_n3075_ & ~new_n3076_;
  assign new_n3078_ = ~new_n3074_ & new_n3077_;
  assign new_n3079_ = new_n3073_ & new_n3078_;
  assign new_n3080_ = new_n1772_ & new_n2879_;
  assign new_n3081_ = new_n1772_ & new_n2885_;
  assign new_n3082_ = ~new_n3080_ & ~new_n3081_;
  assign new_n3083_ = new_n1772_ & new_n2887_;
  assign new_n3084_ = new_n1772_ & new_n2883_;
  assign new_n3085_ = ~new_n3083_ & ~new_n3084_;
  assign new_n3086_ = new_n3082_ & new_n3085_;
  assign new_n3087_ = new_n1772_ & new_n2900_;
  assign new_n3088_ = new_n1772_ & new_n2894_;
  assign new_n3089_ = new_n1772_ & new_n2897_;
  assign new_n3090_ = ~new_n3088_ & ~new_n3089_;
  assign new_n3091_ = ~new_n3087_ & new_n3090_;
  assign new_n3092_ = new_n3086_ & new_n3091_;
  assign new_n3093_ = new_n3079_ & new_n3092_;
  assign new_n3094_ = new_n3066_ & new_n3093_;
  assign new_n3095_ = new_n3035_ & new_n3094_;
  assign new_n3096_ = new_n2970_ & new_n3095_;
  assign new_n3097_ = new_n1772_ & new_n2902_;
  assign new_n3098_ = new_n1772_ & new_n2906_;
  assign new_n3099_ = ~new_n3097_ & ~new_n3098_;
  assign new_n3100_ = new_n1772_ & new_n2908_;
  assign new_n3101_ = new_n1772_ & new_n2911_;
  assign new_n3102_ = ~new_n3100_ & ~new_n3101_;
  assign new_n3103_ = new_n3099_ & new_n3102_;
  assign new_n3104_ = new_n1772_ & new_n2913_;
  assign new_n3105_ = new_n1772_ & new_n2918_;
  assign new_n3106_ = ~new_n3104_ & ~new_n3105_;
  assign new_n3107_ = new_n1772_ & new_n2921_;
  assign new_n3108_ = new_n1772_ & new_n2924_;
  assign new_n3109_ = ~new_n3107_ & ~new_n3108_;
  assign new_n3110_ = new_n3106_ & new_n3109_;
  assign new_n3111_ = new_n3103_ & new_n3110_;
  assign new_n3112_ = new_n1772_ & new_n2926_;
  assign new_n3113_ = new_n1772_ & new_n2932_;
  assign new_n3114_ = ~new_n3112_ & ~new_n3113_;
  assign new_n3115_ = new_n1772_ & new_n2934_;
  assign new_n3116_ = new_n1772_ & new_n2930_;
  assign new_n3117_ = ~new_n3115_ & ~new_n3116_;
  assign new_n3118_ = new_n3114_ & new_n3117_;
  assign new_n3119_ = new_n1858_ & new_n2840_;
  assign new_n3120_ = new_n1772_ & new_n2940_;
  assign new_n3121_ = new_n1772_ & new_n2942_;
  assign new_n3122_ = ~new_n3120_ & ~new_n3121_;
  assign new_n3123_ = ~new_n3119_ & new_n3122_;
  assign new_n3124_ = new_n3118_ & new_n3123_;
  assign new_n3125_ = new_n3111_ & new_n3124_;
  assign new_n3126_ = new_n1858_ & new_n2851_;
  assign new_n3127_ = new_n1858_ & new_n2853_;
  assign new_n3128_ = ~new_n3126_ & ~new_n3127_;
  assign new_n3129_ = new_n1858_ & new_n2856_;
  assign new_n3130_ = new_n1858_ & new_n2858_;
  assign new_n3131_ = ~new_n3129_ & ~new_n3130_;
  assign new_n3132_ = new_n3128_ & new_n3131_;
  assign new_n3133_ = new_n1858_ & new_n2862_;
  assign new_n3134_ = new_n1858_ & new_n2864_;
  assign new_n3135_ = new_n1858_ & new_n2866_;
  assign new_n3136_ = ~new_n3134_ & ~new_n3135_;
  assign new_n3137_ = ~new_n3133_ & new_n3136_;
  assign new_n3138_ = new_n3132_ & new_n3137_;
  assign new_n3139_ = new_n1858_ & new_n2872_;
  assign new_n3140_ = new_n1858_ & new_n2874_;
  assign new_n3141_ = ~new_n3139_ & ~new_n3140_;
  assign new_n3142_ = new_n1858_ & new_n2877_;
  assign new_n3143_ = new_n1858_ & new_n2879_;
  assign new_n3144_ = ~new_n3142_ & ~new_n3143_;
  assign new_n3145_ = new_n3141_ & new_n3144_;
  assign new_n3146_ = new_n1858_ & new_n2883_;
  assign new_n3147_ = new_n1858_ & new_n2885_;
  assign new_n3148_ = new_n1858_ & new_n2887_;
  assign new_n3149_ = ~new_n3147_ & ~new_n3148_;
  assign new_n3150_ = ~new_n3146_ & new_n3149_;
  assign new_n3151_ = new_n3145_ & new_n3150_;
  assign new_n3152_ = new_n3138_ & new_n3151_;
  assign new_n3153_ = new_n3125_ & new_n3152_;
  assign new_n3154_ = new_n1858_ & new_n2894_;
  assign new_n3155_ = new_n1858_ & new_n2897_;
  assign new_n3156_ = ~new_n3154_ & ~new_n3155_;
  assign new_n3157_ = new_n1858_ & new_n2900_;
  assign new_n3158_ = new_n1858_ & new_n2902_;
  assign new_n3159_ = ~new_n3157_ & ~new_n3158_;
  assign new_n3160_ = new_n3156_ & new_n3159_;
  assign new_n3161_ = new_n1858_ & new_n2906_;
  assign new_n3162_ = new_n1858_ & new_n2908_;
  assign new_n3163_ = ~new_n3161_ & ~new_n3162_;
  assign new_n3164_ = new_n1858_ & new_n2911_;
  assign new_n3165_ = new_n1858_ & new_n2913_;
  assign new_n3166_ = ~new_n3164_ & ~new_n3165_;
  assign new_n3167_ = new_n3163_ & new_n3166_;
  assign new_n3168_ = new_n3160_ & new_n3167_;
  assign new_n3169_ = new_n1858_ & new_n2918_;
  assign new_n3170_ = new_n1858_ & new_n2921_;
  assign new_n3171_ = ~new_n3169_ & ~new_n3170_;
  assign new_n3172_ = new_n1858_ & new_n2924_;
  assign new_n3173_ = new_n1858_ & new_n2926_;
  assign new_n3174_ = ~new_n3172_ & ~new_n3173_;
  assign new_n3175_ = new_n3171_ & new_n3174_;
  assign new_n3176_ = new_n1858_ & new_n2930_;
  assign new_n3177_ = new_n1858_ & new_n2932_;
  assign new_n3178_ = new_n1858_ & new_n2934_;
  assign new_n3179_ = ~new_n3177_ & ~new_n3178_;
  assign new_n3180_ = ~new_n3176_ & new_n3179_;
  assign new_n3181_ = new_n3175_ & new_n3180_;
  assign new_n3182_ = new_n3168_ & new_n3181_;
  assign new_n3183_ = new_n1858_ & new_n2940_;
  assign new_n3184_ = new_n1858_ & new_n2942_;
  assign new_n3185_ = ~new_n3183_ & ~new_n3184_;
  assign new_n3186_ = new_n58_ & new_n3007_;
  assign new_n3187_ = new_n1741_ & new_n3186_;
  assign new_n3188_ = new_n2780_ & new_n3187_;
  assign new_n3189_ = new_n2791_ & new_n3187_;
  assign new_n3190_ = ~new_n3188_ & ~new_n3189_;
  assign new_n3191_ = new_n3185_ & new_n3190_;
  assign new_n3192_ = ~A201 & ~A166;
  assign new_n3193_ = new_n2793_ & new_n3192_;
  assign new_n3194_ = new_n1741_ & new_n3193_;
  assign new_n3195_ = new_n2780_ & new_n3194_;
  assign new_n3196_ = new_n2781_ & new_n3192_;
  assign new_n3197_ = new_n1741_ & new_n3196_;
  assign new_n3198_ = new_n2780_ & new_n3197_;
  assign new_n3199_ = new_n2791_ & new_n3197_;
  assign new_n3200_ = ~new_n3198_ & ~new_n3199_;
  assign new_n3201_ = ~new_n3195_ & new_n3200_;
  assign new_n3202_ = new_n3191_ & new_n3201_;
  assign new_n3203_ = new_n2791_ & new_n3194_;
  assign new_n3204_ = new_n1908_ & new_n2291_;
  assign new_n3205_ = ~new_n3203_ & ~new_n3204_;
  assign new_n3206_ = new_n1908_ & new_n2294_;
  assign new_n3207_ = new_n1908_ & new_n2299_;
  assign new_n3208_ = ~new_n3206_ & ~new_n3207_;
  assign new_n3209_ = new_n3205_ & new_n3208_;
  assign new_n3210_ = new_n1908_ & new_n2309_;
  assign new_n3211_ = new_n1908_ & new_n2302_;
  assign new_n3212_ = new_n1908_ & new_n2306_;
  assign new_n3213_ = ~new_n3211_ & ~new_n3212_;
  assign new_n3214_ = ~new_n3210_ & new_n3213_;
  assign new_n3215_ = new_n3209_ & new_n3214_;
  assign new_n3216_ = new_n3202_ & new_n3215_;
  assign new_n3217_ = new_n3182_ & new_n3216_;
  assign new_n3218_ = new_n3153_ & new_n3217_;
  assign new_n3219_ = new_n1908_ & new_n2315_;
  assign new_n3220_ = new_n1908_ & new_n2318_;
  assign new_n3221_ = ~new_n3219_ & ~new_n3220_;
  assign new_n3222_ = new_n1908_ & new_n2322_;
  assign new_n3223_ = new_n1908_ & new_n2324_;
  assign new_n3224_ = ~new_n3222_ & ~new_n3223_;
  assign new_n3225_ = new_n3221_ & new_n3224_;
  assign new_n3226_ = new_n1908_ & new_n2329_;
  assign new_n3227_ = new_n1908_ & new_n2331_;
  assign new_n3228_ = ~new_n3226_ & ~new_n3227_;
  assign new_n3229_ = new_n1906_ & new_n2291_;
  assign new_n3230_ = new_n1906_ & new_n2294_;
  assign new_n3231_ = ~new_n3229_ & ~new_n3230_;
  assign new_n3232_ = new_n3228_ & new_n3231_;
  assign new_n3233_ = new_n3225_ & new_n3232_;
  assign new_n3234_ = new_n1906_ & new_n2299_;
  assign new_n3235_ = new_n1906_ & new_n2302_;
  assign new_n3236_ = ~new_n3234_ & ~new_n3235_;
  assign new_n3237_ = new_n1906_ & new_n2306_;
  assign new_n3238_ = new_n1906_ & new_n2309_;
  assign new_n3239_ = ~new_n3237_ & ~new_n3238_;
  assign new_n3240_ = new_n3236_ & new_n3239_;
  assign new_n3241_ = new_n1906_ & new_n2322_;
  assign new_n3242_ = new_n1906_ & new_n2315_;
  assign new_n3243_ = new_n1906_ & new_n2318_;
  assign new_n3244_ = ~new_n3242_ & ~new_n3243_;
  assign new_n3245_ = ~new_n3241_ & new_n3244_;
  assign new_n3246_ = new_n3240_ & new_n3245_;
  assign new_n3247_ = new_n3233_ & new_n3246_;
  assign new_n3248_ = new_n1906_ & new_n2324_;
  assign new_n3249_ = new_n1906_ & new_n2329_;
  assign new_n3250_ = ~new_n3248_ & ~new_n3249_;
  assign new_n3251_ = new_n1906_ & new_n2331_;
  assign new_n3252_ = new_n1905_ & new_n2782_;
  assign new_n3253_ = new_n2780_ & new_n3252_;
  assign new_n3254_ = ~new_n3251_ & ~new_n3253_;
  assign new_n3255_ = new_n3250_ & new_n3254_;
  assign new_n3256_ = new_n1905_ & new_n2794_;
  assign new_n3257_ = new_n2791_ & new_n3256_;
  assign new_n3258_ = new_n2791_ & new_n3252_;
  assign new_n3259_ = new_n2780_ & new_n3256_;
  assign new_n3260_ = ~new_n3258_ & ~new_n3259_;
  assign new_n3261_ = ~new_n3257_ & new_n3260_;
  assign new_n3262_ = new_n3255_ & new_n3261_;
  assign new_n3263_ = new_n1919_ & new_n2291_;
  assign new_n3264_ = new_n1919_ & new_n2294_;
  assign new_n3265_ = ~new_n3263_ & ~new_n3264_;
  assign new_n3266_ = new_n1919_ & new_n2299_;
  assign new_n3267_ = new_n1919_ & new_n2302_;
  assign new_n3268_ = ~new_n3266_ & ~new_n3267_;
  assign new_n3269_ = new_n3265_ & new_n3268_;
  assign new_n3270_ = new_n1919_ & new_n2315_;
  assign new_n3271_ = new_n1919_ & new_n2306_;
  assign new_n3272_ = new_n1919_ & new_n2309_;
  assign new_n3273_ = ~new_n3271_ & ~new_n3272_;
  assign new_n3274_ = ~new_n3270_ & new_n3273_;
  assign new_n3275_ = new_n3269_ & new_n3274_;
  assign new_n3276_ = new_n3262_ & new_n3275_;
  assign new_n3277_ = new_n3247_ & new_n3276_;
  assign new_n3278_ = new_n1919_ & new_n2318_;
  assign new_n3279_ = new_n1919_ & new_n2322_;
  assign new_n3280_ = ~new_n3278_ & ~new_n3279_;
  assign new_n3281_ = new_n1919_ & new_n2324_;
  assign new_n3282_ = new_n1919_ & new_n2329_;
  assign new_n3283_ = ~new_n3281_ & ~new_n3282_;
  assign new_n3284_ = new_n3280_ & new_n3283_;
  assign new_n3285_ = new_n1918_ & new_n2828_;
  assign new_n3286_ = new_n2791_ & new_n3285_;
  assign new_n3287_ = new_n1919_ & new_n2331_;
  assign new_n3288_ = new_n2780_ & new_n3285_;
  assign new_n3289_ = ~new_n3287_ & ~new_n3288_;
  assign new_n3290_ = ~new_n3286_ & new_n3289_;
  assign new_n3291_ = new_n3284_ & new_n3290_;
  assign new_n3292_ = new_n1918_ & new_n2833_;
  assign new_n3293_ = new_n2780_ & new_n3292_;
  assign new_n3294_ = new_n2791_ & new_n3292_;
  assign new_n3295_ = ~new_n3293_ & ~new_n3294_;
  assign new_n3296_ = new_n1923_ & new_n2843_;
  assign new_n3297_ = new_n2780_ & new_n3296_;
  assign new_n3298_ = new_n2791_ & new_n3296_;
  assign new_n3299_ = ~new_n3297_ & ~new_n3298_;
  assign new_n3300_ = new_n3295_ & new_n3299_;
  assign new_n3301_ = new_n1957_ & new_n2853_;
  assign new_n3302_ = new_n1957_ & new_n2840_;
  assign new_n3303_ = new_n1957_ & new_n2851_;
  assign new_n3304_ = ~new_n3302_ & ~new_n3303_;
  assign new_n3305_ = ~new_n3301_ & new_n3304_;
  assign new_n3306_ = new_n3300_ & new_n3305_;
  assign new_n3307_ = new_n3291_ & new_n3306_;
  assign new_n3308_ = new_n1957_ & new_n2856_;
  assign new_n3309_ = new_n1957_ & new_n2858_;
  assign new_n3310_ = ~new_n3308_ & ~new_n3309_;
  assign new_n3311_ = new_n1957_ & new_n2864_;
  assign new_n3312_ = new_n1957_ & new_n2866_;
  assign new_n3313_ = ~new_n3311_ & ~new_n3312_;
  assign new_n3314_ = new_n3310_ & new_n3313_;
  assign new_n3315_ = new_n1957_ & new_n2874_;
  assign new_n3316_ = new_n1957_ & new_n2862_;
  assign new_n3317_ = new_n1957_ & new_n2872_;
  assign new_n3318_ = ~new_n3316_ & ~new_n3317_;
  assign new_n3319_ = ~new_n3315_ & new_n3318_;
  assign new_n3320_ = new_n3314_ & new_n3319_;
  assign new_n3321_ = new_n1957_ & new_n2877_;
  assign new_n3322_ = new_n1957_ & new_n2879_;
  assign new_n3323_ = ~new_n3321_ & ~new_n3322_;
  assign new_n3324_ = new_n1957_ & new_n2885_;
  assign new_n3325_ = new_n1957_ & new_n2887_;
  assign new_n3326_ = ~new_n3324_ & ~new_n3325_;
  assign new_n3327_ = new_n3323_ & new_n3326_;
  assign new_n3328_ = new_n1957_ & new_n2897_;
  assign new_n3329_ = new_n1957_ & new_n2883_;
  assign new_n3330_ = new_n1957_ & new_n2894_;
  assign new_n3331_ = ~new_n3329_ & ~new_n3330_;
  assign new_n3332_ = ~new_n3328_ & new_n3331_;
  assign new_n3333_ = new_n3327_ & new_n3332_;
  assign new_n3334_ = new_n3320_ & new_n3333_;
  assign new_n3335_ = new_n3307_ & new_n3334_;
  assign new_n3336_ = new_n3277_ & new_n3335_;
  assign new_n3337_ = new_n3218_ & new_n3336_;
  assign new_n3338_ = new_n3096_ & new_n3337_;
  assign new_n3339_ = new_n2812_ & new_n3338_;
  assign new_n3340_ = new_n1957_ & new_n2900_;
  assign new_n3341_ = new_n1957_ & new_n2902_;
  assign new_n3342_ = ~new_n3340_ & ~new_n3341_;
  assign new_n3343_ = new_n1957_ & new_n2906_;
  assign new_n3344_ = new_n1957_ & new_n2908_;
  assign new_n3345_ = ~new_n3343_ & ~new_n3344_;
  assign new_n3346_ = new_n3342_ & new_n3345_;
  assign new_n3347_ = new_n1957_ & new_n2911_;
  assign new_n3348_ = new_n1957_ & new_n2913_;
  assign new_n3349_ = ~new_n3347_ & ~new_n3348_;
  assign new_n3350_ = new_n1957_ & new_n2918_;
  assign new_n3351_ = new_n1957_ & new_n2921_;
  assign new_n3352_ = ~new_n3350_ & ~new_n3351_;
  assign new_n3353_ = new_n3349_ & new_n3352_;
  assign new_n3354_ = new_n3346_ & new_n3353_;
  assign new_n3355_ = new_n1957_ & new_n2924_;
  assign new_n3356_ = new_n1957_ & new_n2926_;
  assign new_n3357_ = ~new_n3355_ & ~new_n3356_;
  assign new_n3358_ = new_n1957_ & new_n2932_;
  assign new_n3359_ = new_n1957_ & new_n2934_;
  assign new_n3360_ = ~new_n3358_ & ~new_n3359_;
  assign new_n3361_ = new_n3357_ & new_n3360_;
  assign new_n3362_ = new_n1957_ & new_n2942_;
  assign new_n3363_ = new_n1957_ & new_n2930_;
  assign new_n3364_ = new_n1957_ & new_n2940_;
  assign new_n3365_ = ~new_n3363_ & ~new_n3364_;
  assign new_n3366_ = ~new_n3362_ & new_n3365_;
  assign new_n3367_ = new_n3361_ & new_n3366_;
  assign new_n3368_ = new_n3354_ & new_n3367_;
  assign new_n3369_ = new_n2040_ & new_n2840_;
  assign new_n3370_ = new_n2040_ & new_n2851_;
  assign new_n3371_ = ~new_n3369_ & ~new_n3370_;
  assign new_n3372_ = new_n2040_ & new_n2853_;
  assign new_n3373_ = new_n2040_ & new_n2856_;
  assign new_n3374_ = ~new_n3372_ & ~new_n3373_;
  assign new_n3375_ = new_n3371_ & new_n3374_;
  assign new_n3376_ = new_n2040_ & new_n2866_;
  assign new_n3377_ = new_n2040_ & new_n2858_;
  assign new_n3378_ = new_n2040_ & new_n2864_;
  assign new_n3379_ = ~new_n3377_ & ~new_n3378_;
  assign new_n3380_ = ~new_n3376_ & new_n3379_;
  assign new_n3381_ = new_n3375_ & new_n3380_;
  assign new_n3382_ = new_n2040_ & new_n2862_;
  assign new_n3383_ = new_n2040_ & new_n2872_;
  assign new_n3384_ = ~new_n3382_ & ~new_n3383_;
  assign new_n3385_ = new_n2040_ & new_n2874_;
  assign new_n3386_ = new_n2040_ & new_n2877_;
  assign new_n3387_ = ~new_n3385_ & ~new_n3386_;
  assign new_n3388_ = new_n3384_ & new_n3387_;
  assign new_n3389_ = new_n2040_ & new_n2887_;
  assign new_n3390_ = new_n2040_ & new_n2879_;
  assign new_n3391_ = new_n2040_ & new_n2885_;
  assign new_n3392_ = ~new_n3390_ & ~new_n3391_;
  assign new_n3393_ = ~new_n3389_ & new_n3392_;
  assign new_n3394_ = new_n3388_ & new_n3393_;
  assign new_n3395_ = new_n3381_ & new_n3394_;
  assign new_n3396_ = new_n3368_ & new_n3395_;
  assign new_n3397_ = new_n2040_ & new_n2883_;
  assign new_n3398_ = new_n2040_ & new_n2894_;
  assign new_n3399_ = ~new_n3397_ & ~new_n3398_;
  assign new_n3400_ = new_n2040_ & new_n2897_;
  assign new_n3401_ = new_n2040_ & new_n2900_;
  assign new_n3402_ = ~new_n3400_ & ~new_n3401_;
  assign new_n3403_ = new_n3399_ & new_n3402_;
  assign new_n3404_ = new_n2040_ & new_n2902_;
  assign new_n3405_ = new_n2040_ & new_n2906_;
  assign new_n3406_ = ~new_n3404_ & ~new_n3405_;
  assign new_n3407_ = new_n2040_ & new_n2908_;
  assign new_n3408_ = new_n2040_ & new_n2911_;
  assign new_n3409_ = ~new_n3407_ & ~new_n3408_;
  assign new_n3410_ = new_n3406_ & new_n3409_;
  assign new_n3411_ = new_n3403_ & new_n3410_;
  assign new_n3412_ = new_n2040_ & new_n2913_;
  assign new_n3413_ = new_n2040_ & new_n2918_;
  assign new_n3414_ = ~new_n3412_ & ~new_n3413_;
  assign new_n3415_ = new_n2040_ & new_n2921_;
  assign new_n3416_ = new_n2040_ & new_n2924_;
  assign new_n3417_ = ~new_n3415_ & ~new_n3416_;
  assign new_n3418_ = new_n3414_ & new_n3417_;
  assign new_n3419_ = new_n2040_ & new_n2934_;
  assign new_n3420_ = new_n2040_ & new_n2926_;
  assign new_n3421_ = new_n2040_ & new_n2932_;
  assign new_n3422_ = ~new_n3420_ & ~new_n3421_;
  assign new_n3423_ = ~new_n3419_ & new_n3422_;
  assign new_n3424_ = new_n3418_ & new_n3423_;
  assign new_n3425_ = new_n3411_ & new_n3424_;
  assign new_n3426_ = new_n2040_ & new_n2930_;
  assign new_n3427_ = new_n2040_ & new_n2940_;
  assign new_n3428_ = ~new_n3426_ & ~new_n3427_;
  assign new_n3429_ = new_n2040_ & new_n2942_;
  assign new_n3430_ = new_n1923_ & new_n3008_;
  assign new_n3431_ = new_n2780_ & new_n3430_;
  assign new_n3432_ = ~new_n3429_ & ~new_n3431_;
  assign new_n3433_ = new_n3428_ & new_n3432_;
  assign new_n3434_ = new_n1923_ & new_n3017_;
  assign new_n3435_ = new_n2791_ & new_n3434_;
  assign new_n3436_ = new_n2791_ & new_n3430_;
  assign new_n3437_ = new_n2780_ & new_n3434_;
  assign new_n3438_ = ~new_n3436_ & ~new_n3437_;
  assign new_n3439_ = ~new_n3435_ & new_n3438_;
  assign new_n3440_ = new_n3433_ & new_n3439_;
  assign new_n3441_ = new_n1923_ & new_n3022_;
  assign new_n3442_ = new_n2780_ & new_n3441_;
  assign new_n3443_ = new_n2791_ & new_n3441_;
  assign new_n3444_ = ~new_n3442_ & ~new_n3443_;
  assign new_n3445_ = new_n2086_ & new_n2291_;
  assign new_n3446_ = new_n2086_ & new_n2294_;
  assign new_n3447_ = ~new_n3445_ & ~new_n3446_;
  assign new_n3448_ = new_n3444_ & new_n3447_;
  assign new_n3449_ = new_n2086_ & new_n2306_;
  assign new_n3450_ = new_n2086_ & new_n2299_;
  assign new_n3451_ = new_n2086_ & new_n2302_;
  assign new_n3452_ = ~new_n3450_ & ~new_n3451_;
  assign new_n3453_ = ~new_n3449_ & new_n3452_;
  assign new_n3454_ = new_n3448_ & new_n3453_;
  assign new_n3455_ = new_n3440_ & new_n3454_;
  assign new_n3456_ = new_n3425_ & new_n3455_;
  assign new_n3457_ = new_n3396_ & new_n3456_;
  assign new_n3458_ = new_n2086_ & new_n2309_;
  assign new_n3459_ = new_n2086_ & new_n2315_;
  assign new_n3460_ = ~new_n3458_ & ~new_n3459_;
  assign new_n3461_ = new_n2086_ & new_n2318_;
  assign new_n3462_ = new_n2086_ & new_n2322_;
  assign new_n3463_ = ~new_n3461_ & ~new_n3462_;
  assign new_n3464_ = new_n3460_ & new_n3463_;
  assign new_n3465_ = new_n2086_ & new_n2324_;
  assign new_n3466_ = new_n2086_ & new_n2329_;
  assign new_n3467_ = ~new_n3465_ & ~new_n3466_;
  assign new_n3468_ = new_n2086_ & new_n2331_;
  assign new_n3469_ = new_n2090_ & new_n3052_;
  assign new_n3470_ = new_n2780_ & new_n3469_;
  assign new_n3471_ = ~new_n3468_ & ~new_n3470_;
  assign new_n3472_ = new_n3467_ & new_n3471_;
  assign new_n3473_ = new_n3464_ & new_n3472_;
  assign new_n3474_ = new_n2791_ & new_n3469_;
  assign new_n3475_ = new_n2122_ & new_n2840_;
  assign new_n3476_ = ~new_n3474_ & ~new_n3475_;
  assign new_n3477_ = new_n2122_ & new_n2851_;
  assign new_n3478_ = new_n2122_ & new_n2853_;
  assign new_n3479_ = ~new_n3477_ & ~new_n3478_;
  assign new_n3480_ = new_n3476_ & new_n3479_;
  assign new_n3481_ = new_n2122_ & new_n2864_;
  assign new_n3482_ = new_n2122_ & new_n2856_;
  assign new_n3483_ = new_n2122_ & new_n2858_;
  assign new_n3484_ = ~new_n3482_ & ~new_n3483_;
  assign new_n3485_ = ~new_n3481_ & new_n3484_;
  assign new_n3486_ = new_n3480_ & new_n3485_;
  assign new_n3487_ = new_n3473_ & new_n3486_;
  assign new_n3488_ = new_n2122_ & new_n2866_;
  assign new_n3489_ = new_n2122_ & new_n2862_;
  assign new_n3490_ = ~new_n3488_ & ~new_n3489_;
  assign new_n3491_ = new_n2122_ & new_n2872_;
  assign new_n3492_ = new_n2122_ & new_n2874_;
  assign new_n3493_ = ~new_n3491_ & ~new_n3492_;
  assign new_n3494_ = new_n3490_ & new_n3493_;
  assign new_n3495_ = new_n2122_ & new_n2885_;
  assign new_n3496_ = new_n2122_ & new_n2877_;
  assign new_n3497_ = new_n2122_ & new_n2879_;
  assign new_n3498_ = ~new_n3496_ & ~new_n3497_;
  assign new_n3499_ = ~new_n3495_ & new_n3498_;
  assign new_n3500_ = new_n3494_ & new_n3499_;
  assign new_n3501_ = new_n2122_ & new_n2887_;
  assign new_n3502_ = new_n2122_ & new_n2883_;
  assign new_n3503_ = ~new_n3501_ & ~new_n3502_;
  assign new_n3504_ = new_n2122_ & new_n2894_;
  assign new_n3505_ = new_n2122_ & new_n2897_;
  assign new_n3506_ = ~new_n3504_ & ~new_n3505_;
  assign new_n3507_ = new_n3503_ & new_n3506_;
  assign new_n3508_ = new_n2122_ & new_n2906_;
  assign new_n3509_ = new_n2122_ & new_n2900_;
  assign new_n3510_ = new_n2122_ & new_n2902_;
  assign new_n3511_ = ~new_n3509_ & ~new_n3510_;
  assign new_n3512_ = ~new_n3508_ & new_n3511_;
  assign new_n3513_ = new_n3507_ & new_n3512_;
  assign new_n3514_ = new_n3500_ & new_n3513_;
  assign new_n3515_ = new_n3487_ & new_n3514_;
  assign new_n3516_ = new_n2122_ & new_n2908_;
  assign new_n3517_ = new_n2122_ & new_n2911_;
  assign new_n3518_ = ~new_n3516_ & ~new_n3517_;
  assign new_n3519_ = new_n2122_ & new_n2913_;
  assign new_n3520_ = new_n2122_ & new_n2918_;
  assign new_n3521_ = ~new_n3519_ & ~new_n3520_;
  assign new_n3522_ = new_n3518_ & new_n3521_;
  assign new_n3523_ = new_n2122_ & new_n2921_;
  assign new_n3524_ = new_n2122_ & new_n2924_;
  assign new_n3525_ = ~new_n3523_ & ~new_n3524_;
  assign new_n3526_ = new_n2122_ & new_n2926_;
  assign new_n3527_ = new_n2122_ & new_n2932_;
  assign new_n3528_ = ~new_n3526_ & ~new_n3527_;
  assign new_n3529_ = new_n3525_ & new_n3528_;
  assign new_n3530_ = new_n3522_ & new_n3529_;
  assign new_n3531_ = new_n2122_ & new_n2934_;
  assign new_n3532_ = new_n2122_ & new_n2930_;
  assign new_n3533_ = ~new_n3531_ & ~new_n3532_;
  assign new_n3534_ = new_n2122_ & new_n2940_;
  assign new_n3535_ = new_n2122_ & new_n2942_;
  assign new_n3536_ = ~new_n3534_ & ~new_n3535_;
  assign new_n3537_ = new_n3533_ & new_n3536_;
  assign new_n3538_ = new_n2206_ & new_n2853_;
  assign new_n3539_ = new_n2206_ & new_n2840_;
  assign new_n3540_ = new_n2206_ & new_n2851_;
  assign new_n3541_ = ~new_n3539_ & ~new_n3540_;
  assign new_n3542_ = ~new_n3538_ & new_n3541_;
  assign new_n3543_ = new_n3537_ & new_n3542_;
  assign new_n3544_ = new_n3530_ & new_n3543_;
  assign new_n3545_ = new_n2206_ & new_n2856_;
  assign new_n3546_ = new_n2206_ & new_n2858_;
  assign new_n3547_ = ~new_n3545_ & ~new_n3546_;
  assign new_n3548_ = new_n2206_ & new_n2864_;
  assign new_n3549_ = new_n2206_ & new_n2866_;
  assign new_n3550_ = ~new_n3548_ & ~new_n3549_;
  assign new_n3551_ = new_n3547_ & new_n3550_;
  assign new_n3552_ = new_n2206_ & new_n2874_;
  assign new_n3553_ = new_n2206_ & new_n2862_;
  assign new_n3554_ = new_n2206_ & new_n2872_;
  assign new_n3555_ = ~new_n3553_ & ~new_n3554_;
  assign new_n3556_ = ~new_n3552_ & new_n3555_;
  assign new_n3557_ = new_n3551_ & new_n3556_;
  assign new_n3558_ = new_n2206_ & new_n2877_;
  assign new_n3559_ = new_n2206_ & new_n2879_;
  assign new_n3560_ = ~new_n3558_ & ~new_n3559_;
  assign new_n3561_ = new_n2206_ & new_n2885_;
  assign new_n3562_ = new_n2206_ & new_n2887_;
  assign new_n3563_ = ~new_n3561_ & ~new_n3562_;
  assign new_n3564_ = new_n3560_ & new_n3563_;
  assign new_n3565_ = new_n2206_ & new_n2897_;
  assign new_n3566_ = new_n2206_ & new_n2883_;
  assign new_n3567_ = new_n2206_ & new_n2894_;
  assign new_n3568_ = ~new_n3566_ & ~new_n3567_;
  assign new_n3569_ = ~new_n3565_ & new_n3568_;
  assign new_n3570_ = new_n3564_ & new_n3569_;
  assign new_n3571_ = new_n3557_ & new_n3570_;
  assign new_n3572_ = new_n3544_ & new_n3571_;
  assign new_n3573_ = new_n3515_ & new_n3572_;
  assign new_n3574_ = new_n3457_ & new_n3573_;
  assign new_n3575_ = new_n2206_ & new_n2900_;
  assign new_n3576_ = new_n2206_ & new_n2902_;
  assign new_n3577_ = ~new_n3575_ & ~new_n3576_;
  assign new_n3578_ = new_n2206_ & new_n2906_;
  assign new_n3579_ = new_n2206_ & new_n2908_;
  assign new_n3580_ = ~new_n3578_ & ~new_n3579_;
  assign new_n3581_ = new_n3577_ & new_n3580_;
  assign new_n3582_ = new_n2206_ & new_n2911_;
  assign new_n3583_ = new_n2206_ & new_n2913_;
  assign new_n3584_ = ~new_n3582_ & ~new_n3583_;
  assign new_n3585_ = new_n2206_ & new_n2918_;
  assign new_n3586_ = new_n2206_ & new_n2921_;
  assign new_n3587_ = ~new_n3585_ & ~new_n3586_;
  assign new_n3588_ = new_n3584_ & new_n3587_;
  assign new_n3589_ = new_n3581_ & new_n3588_;
  assign new_n3590_ = new_n2206_ & new_n2924_;
  assign new_n3591_ = new_n2206_ & new_n2926_;
  assign new_n3592_ = ~new_n3590_ & ~new_n3591_;
  assign new_n3593_ = new_n2206_ & new_n2932_;
  assign new_n3594_ = new_n2206_ & new_n2934_;
  assign new_n3595_ = ~new_n3593_ & ~new_n3594_;
  assign new_n3596_ = new_n3592_ & new_n3595_;
  assign new_n3597_ = new_n2206_ & new_n2942_;
  assign new_n3598_ = new_n2206_ & new_n2930_;
  assign new_n3599_ = new_n2206_ & new_n2940_;
  assign new_n3600_ = ~new_n3598_ & ~new_n3599_;
  assign new_n3601_ = ~new_n3597_ & new_n3600_;
  assign new_n3602_ = new_n3596_ & new_n3601_;
  assign new_n3603_ = new_n3589_ & new_n3602_;
  assign new_n3604_ = new_n2090_ & new_n3186_;
  assign new_n3605_ = new_n2780_ & new_n3604_;
  assign new_n3606_ = new_n2791_ & new_n3604_;
  assign new_n3607_ = ~new_n3605_ & ~new_n3606_;
  assign new_n3608_ = new_n2090_ & new_n3196_;
  assign new_n3609_ = new_n2780_ & new_n3608_;
  assign new_n3610_ = new_n2791_ & new_n3608_;
  assign new_n3611_ = ~new_n3609_ & ~new_n3610_;
  assign new_n3612_ = new_n3607_ & new_n3611_;
  assign new_n3613_ = new_n2252_ & new_n2291_;
  assign new_n3614_ = new_n2090_ & new_n3193_;
  assign new_n3615_ = new_n2780_ & new_n3614_;
  assign new_n3616_ = new_n2791_ & new_n3614_;
  assign new_n3617_ = ~new_n3615_ & ~new_n3616_;
  assign new_n3618_ = ~new_n3613_ & new_n3617_;
  assign new_n3619_ = new_n3612_ & new_n3618_;
  assign new_n3620_ = new_n2252_ & new_n2294_;
  assign new_n3621_ = new_n2252_ & new_n2299_;
  assign new_n3622_ = ~new_n3620_ & ~new_n3621_;
  assign new_n3623_ = new_n2252_ & new_n2302_;
  assign new_n3624_ = new_n2252_ & new_n2306_;
  assign new_n3625_ = ~new_n3623_ & ~new_n3624_;
  assign new_n3626_ = new_n3622_ & new_n3625_;
  assign new_n3627_ = new_n2252_ & new_n2318_;
  assign new_n3628_ = new_n2252_ & new_n2309_;
  assign new_n3629_ = new_n2252_ & new_n2315_;
  assign new_n3630_ = ~new_n3628_ & ~new_n3629_;
  assign new_n3631_ = ~new_n3627_ & new_n3630_;
  assign new_n3632_ = new_n3626_ & new_n3631_;
  assign new_n3633_ = new_n3619_ & new_n3632_;
  assign new_n3634_ = new_n3603_ & new_n3633_;
  assign new_n3635_ = new_n2252_ & new_n2322_;
  assign new_n3636_ = new_n2252_ & new_n2324_;
  assign new_n3637_ = ~new_n3635_ & ~new_n3636_;
  assign new_n3638_ = new_n2252_ & new_n2329_;
  assign new_n3639_ = new_n2252_ & new_n2331_;
  assign new_n3640_ = ~new_n3638_ & ~new_n3639_;
  assign new_n3641_ = new_n3637_ & new_n3640_;
  assign new_n3642_ = new_n2261_ & new_n2291_;
  assign new_n3643_ = new_n2261_ & new_n2294_;
  assign new_n3644_ = ~new_n3642_ & ~new_n3643_;
  assign new_n3645_ = new_n2261_ & new_n2299_;
  assign new_n3646_ = new_n2261_ & new_n2302_;
  assign new_n3647_ = ~new_n3645_ & ~new_n3646_;
  assign new_n3648_ = new_n3644_ & new_n3647_;
  assign new_n3649_ = new_n3641_ & new_n3648_;
  assign new_n3650_ = new_n2261_ & new_n2306_;
  assign new_n3651_ = new_n2261_ & new_n2309_;
  assign new_n3652_ = ~new_n3650_ & ~new_n3651_;
  assign new_n3653_ = new_n2261_ & new_n2315_;
  assign new_n3654_ = new_n2261_ & new_n2318_;
  assign new_n3655_ = ~new_n3653_ & ~new_n3654_;
  assign new_n3656_ = new_n3652_ & new_n3655_;
  assign new_n3657_ = new_n2261_ & new_n2329_;
  assign new_n3658_ = new_n2261_ & new_n2322_;
  assign new_n3659_ = new_n2261_ & new_n2324_;
  assign new_n3660_ = ~new_n3658_ & ~new_n3659_;
  assign new_n3661_ = ~new_n3657_ & new_n3660_;
  assign new_n3662_ = new_n3656_ & new_n3661_;
  assign new_n3663_ = new_n3649_ & new_n3662_;
  assign new_n3664_ = new_n2261_ & new_n2331_;
  assign new_n3665_ = new_n2260_ & new_n2782_;
  assign new_n3666_ = new_n2780_ & new_n3665_;
  assign new_n3667_ = ~new_n3664_ & ~new_n3666_;
  assign new_n3668_ = new_n2791_ & new_n3665_;
  assign new_n3669_ = new_n2260_ & new_n2794_;
  assign new_n3670_ = new_n2780_ & new_n3669_;
  assign new_n3671_ = ~new_n3668_ & ~new_n3670_;
  assign new_n3672_ = new_n3667_ & new_n3671_;
  assign new_n3673_ = new_n2266_ & new_n2294_;
  assign new_n3674_ = new_n2791_ & new_n3669_;
  assign new_n3675_ = new_n2266_ & new_n2291_;
  assign new_n3676_ = ~new_n3674_ & ~new_n3675_;
  assign new_n3677_ = ~new_n3673_ & new_n3676_;
  assign new_n3678_ = new_n3672_ & new_n3677_;
  assign new_n3679_ = new_n2266_ & new_n2299_;
  assign new_n3680_ = new_n2266_ & new_n2302_;
  assign new_n3681_ = ~new_n3679_ & ~new_n3680_;
  assign new_n3682_ = new_n2266_ & new_n2306_;
  assign new_n3683_ = new_n2266_ & new_n2309_;
  assign new_n3684_ = ~new_n3682_ & ~new_n3683_;
  assign new_n3685_ = new_n3681_ & new_n3684_;
  assign new_n3686_ = new_n2266_ & new_n2322_;
  assign new_n3687_ = new_n2266_ & new_n2315_;
  assign new_n3688_ = new_n2266_ & new_n2318_;
  assign new_n3689_ = ~new_n3687_ & ~new_n3688_;
  assign new_n3690_ = ~new_n3686_ & new_n3689_;
  assign new_n3691_ = new_n3685_ & new_n3690_;
  assign new_n3692_ = new_n3678_ & new_n3691_;
  assign new_n3693_ = new_n3663_ & new_n3692_;
  assign new_n3694_ = new_n3634_ & new_n3693_;
  assign new_n3695_ = new_n2266_ & new_n2324_;
  assign new_n3696_ = new_n2266_ & new_n2329_;
  assign new_n3697_ = ~new_n3695_ & ~new_n3696_;
  assign new_n3698_ = new_n2266_ & new_n2331_;
  assign new_n3699_ = new_n2265_ & new_n2828_;
  assign new_n3700_ = new_n2780_ & new_n3699_;
  assign new_n3701_ = ~new_n3698_ & ~new_n3700_;
  assign new_n3702_ = new_n3697_ & new_n3701_;
  assign new_n3703_ = new_n2791_ & new_n3699_;
  assign new_n3704_ = new_n2265_ & new_n2833_;
  assign new_n3705_ = new_n2780_ & new_n3704_;
  assign new_n3706_ = ~new_n3703_ & ~new_n3705_;
  assign new_n3707_ = new_n2791_ & new_n3704_;
  assign new_n3708_ = new_n2271_ & new_n2291_;
  assign new_n3709_ = ~new_n3707_ & ~new_n3708_;
  assign new_n3710_ = new_n3706_ & new_n3709_;
  assign new_n3711_ = new_n3702_ & new_n3710_;
  assign new_n3712_ = new_n2271_ & new_n2294_;
  assign new_n3713_ = new_n2271_ & new_n2299_;
  assign new_n3714_ = ~new_n3712_ & ~new_n3713_;
  assign new_n3715_ = new_n2271_ & new_n2302_;
  assign new_n3716_ = new_n2271_ & new_n2306_;
  assign new_n3717_ = ~new_n3715_ & ~new_n3716_;
  assign new_n3718_ = new_n3714_ & new_n3717_;
  assign new_n3719_ = new_n2271_ & new_n2318_;
  assign new_n3720_ = new_n2271_ & new_n2309_;
  assign new_n3721_ = new_n2271_ & new_n2315_;
  assign new_n3722_ = ~new_n3720_ & ~new_n3721_;
  assign new_n3723_ = ~new_n3719_ & new_n3722_;
  assign new_n3724_ = new_n3718_ & new_n3723_;
  assign new_n3725_ = new_n3711_ & new_n3724_;
  assign new_n3726_ = new_n2271_ & new_n2322_;
  assign new_n3727_ = new_n2271_ & new_n2324_;
  assign new_n3728_ = ~new_n3726_ & ~new_n3727_;
  assign new_n3729_ = new_n2271_ & new_n2329_;
  assign new_n3730_ = new_n2271_ & new_n2331_;
  assign new_n3731_ = ~new_n3729_ & ~new_n3730_;
  assign new_n3732_ = new_n3728_ & new_n3731_;
  assign new_n3733_ = new_n2270_ & new_n2794_;
  assign new_n3734_ = new_n2780_ & new_n3733_;
  assign new_n3735_ = new_n2270_ & new_n2782_;
  assign new_n3736_ = new_n2780_ & new_n3735_;
  assign new_n3737_ = new_n2791_ & new_n3735_;
  assign new_n3738_ = ~new_n3736_ & ~new_n3737_;
  assign new_n3739_ = ~new_n3734_ & new_n3738_;
  assign new_n3740_ = new_n3732_ & new_n3739_;
  assign new_n3741_ = new_n2791_ & new_n3733_;
  assign new_n3742_ = new_n2286_ & new_n2291_;
  assign new_n3743_ = ~new_n3741_ & ~new_n3742_;
  assign new_n3744_ = new_n2286_ & new_n2294_;
  assign new_n3745_ = new_n2286_ & new_n2299_;
  assign new_n3746_ = ~new_n3744_ & ~new_n3745_;
  assign new_n3747_ = new_n3743_ & new_n3746_;
  assign new_n3748_ = new_n2286_ & new_n2309_;
  assign new_n3749_ = new_n2286_ & new_n2302_;
  assign new_n3750_ = new_n2286_ & new_n2306_;
  assign new_n3751_ = ~new_n3749_ & ~new_n3750_;
  assign new_n3752_ = ~new_n3748_ & new_n3751_;
  assign new_n3753_ = new_n3747_ & new_n3752_;
  assign new_n3754_ = new_n3740_ & new_n3753_;
  assign new_n3755_ = new_n3725_ & new_n3754_;
  assign new_n3756_ = new_n2286_ & new_n2315_;
  assign new_n3757_ = new_n2286_ & new_n2318_;
  assign new_n3758_ = ~new_n3756_ & ~new_n3757_;
  assign new_n3759_ = new_n2286_ & new_n2322_;
  assign new_n3760_ = new_n2286_ & new_n2324_;
  assign new_n3761_ = ~new_n3759_ & ~new_n3760_;
  assign new_n3762_ = new_n3758_ & new_n3761_;
  assign new_n3763_ = new_n2285_ & new_n2828_;
  assign new_n3764_ = new_n2780_ & new_n3763_;
  assign new_n3765_ = new_n2286_ & new_n2329_;
  assign new_n3766_ = new_n2286_ & new_n2331_;
  assign new_n3767_ = ~new_n3765_ & ~new_n3766_;
  assign new_n3768_ = ~new_n3764_ & new_n3767_;
  assign new_n3769_ = new_n3762_ & new_n3768_;
  assign new_n3770_ = new_n2791_ & new_n3763_;
  assign new_n3771_ = new_n2285_ & new_n2833_;
  assign new_n3772_ = new_n2780_ & new_n3771_;
  assign new_n3773_ = ~new_n3770_ & ~new_n3772_;
  assign new_n3774_ = new_n2791_ & new_n3771_;
  assign new_n3775_ = ~A200 & new_n2401_;
  assign new_n3776_ = new_n1284_ & new_n3775_;
  assign new_n3777_ = ~A167 & new_n51_;
  assign new_n3778_ = new_n1039_ & new_n3777_;
  assign new_n3779_ = new_n3776_ & new_n3778_;
  assign new_n3780_ = ~new_n3774_ & ~new_n3779_;
  assign new_n3781_ = new_n3773_ & new_n3780_;
  assign new_n3782_ = new_n1300_ & new_n3775_;
  assign new_n3783_ = new_n3778_ & new_n3782_;
  assign new_n3784_ = new_n1291_ & new_n3775_;
  assign new_n3785_ = new_n3778_ & new_n3784_;
  assign new_n3786_ = new_n1295_ & new_n3775_;
  assign new_n3787_ = new_n3778_ & new_n3786_;
  assign new_n3788_ = ~new_n3785_ & ~new_n3787_;
  assign new_n3789_ = ~new_n3783_ & new_n3788_;
  assign new_n3790_ = new_n3781_ & new_n3789_;
  assign new_n3791_ = new_n3769_ & new_n3790_;
  assign new_n3792_ = ~A200 & new_n2417_;
  assign new_n3793_ = new_n1284_ & new_n3792_;
  assign new_n3794_ = new_n3778_ & new_n3793_;
  assign new_n3795_ = new_n1291_ & new_n3792_;
  assign new_n3796_ = new_n3778_ & new_n3795_;
  assign new_n3797_ = ~new_n3794_ & ~new_n3796_;
  assign new_n3798_ = new_n1295_ & new_n3792_;
  assign new_n3799_ = new_n3778_ & new_n3798_;
  assign new_n3800_ = new_n1300_ & new_n3792_;
  assign new_n3801_ = new_n3778_ & new_n3800_;
  assign new_n3802_ = ~new_n3799_ & ~new_n3801_;
  assign new_n3803_ = new_n3797_ & new_n3802_;
  assign new_n3804_ = ~A200 & new_n2435_;
  assign new_n3805_ = new_n1295_ & new_n3804_;
  assign new_n3806_ = new_n3778_ & new_n3805_;
  assign new_n3807_ = new_n1284_ & new_n3804_;
  assign new_n3808_ = new_n3778_ & new_n3807_;
  assign new_n3809_ = new_n1291_ & new_n3804_;
  assign new_n3810_ = new_n3778_ & new_n3809_;
  assign new_n3811_ = ~new_n3808_ & ~new_n3810_;
  assign new_n3812_ = ~new_n3806_ & new_n3811_;
  assign new_n3813_ = new_n3803_ & new_n3812_;
  assign new_n3814_ = new_n1300_ & new_n3804_;
  assign new_n3815_ = new_n3778_ & new_n3814_;
  assign new_n3816_ = ~A200 & new_n2448_;
  assign new_n3817_ = new_n1284_ & new_n3816_;
  assign new_n3818_ = new_n3778_ & new_n3817_;
  assign new_n3819_ = ~new_n3815_ & ~new_n3818_;
  assign new_n3820_ = new_n1291_ & new_n3816_;
  assign new_n3821_ = new_n3778_ & new_n3820_;
  assign new_n3822_ = new_n1295_ & new_n3816_;
  assign new_n3823_ = new_n3778_ & new_n3822_;
  assign new_n3824_ = ~new_n3821_ & ~new_n3823_;
  assign new_n3825_ = new_n3819_ & new_n3824_;
  assign new_n3826_ = A200 & new_n2401_;
  assign new_n3827_ = new_n1291_ & new_n3826_;
  assign new_n3828_ = ~A167 & new_n37_;
  assign new_n3829_ = new_n1039_ & new_n3828_;
  assign new_n3830_ = new_n3827_ & new_n3829_;
  assign new_n3831_ = new_n1300_ & new_n3816_;
  assign new_n3832_ = new_n3778_ & new_n3831_;
  assign new_n3833_ = new_n1284_ & new_n3826_;
  assign new_n3834_ = new_n3829_ & new_n3833_;
  assign new_n3835_ = ~new_n3832_ & ~new_n3834_;
  assign new_n3836_ = ~new_n3830_ & new_n3835_;
  assign new_n3837_ = new_n3825_ & new_n3836_;
  assign new_n3838_ = new_n3813_ & new_n3837_;
  assign new_n3839_ = new_n3791_ & new_n3838_;
  assign new_n3840_ = new_n3755_ & new_n3839_;
  assign new_n3841_ = new_n3694_ & new_n3840_;
  assign new_n3842_ = new_n3574_ & new_n3841_;
  assign new_n3843_ = new_n1295_ & new_n3826_;
  assign new_n3844_ = new_n3829_ & new_n3843_;
  assign new_n3845_ = new_n1300_ & new_n3826_;
  assign new_n3846_ = new_n3829_ & new_n3845_;
  assign new_n3847_ = ~new_n3844_ & ~new_n3846_;
  assign new_n3848_ = A200 & new_n2417_;
  assign new_n3849_ = new_n1284_ & new_n3848_;
  assign new_n3850_ = new_n3829_ & new_n3849_;
  assign new_n3851_ = new_n1291_ & new_n3848_;
  assign new_n3852_ = new_n3829_ & new_n3851_;
  assign new_n3853_ = ~new_n3850_ & ~new_n3852_;
  assign new_n3854_ = new_n3847_ & new_n3853_;
  assign new_n3855_ = new_n1295_ & new_n3848_;
  assign new_n3856_ = new_n3829_ & new_n3855_;
  assign new_n3857_ = new_n1300_ & new_n3848_;
  assign new_n3858_ = new_n3829_ & new_n3857_;
  assign new_n3859_ = ~new_n3856_ & ~new_n3858_;
  assign new_n3860_ = A200 & new_n2435_;
  assign new_n3861_ = new_n1284_ & new_n3860_;
  assign new_n3862_ = new_n3829_ & new_n3861_;
  assign new_n3863_ = new_n1291_ & new_n3860_;
  assign new_n3864_ = new_n3829_ & new_n3863_;
  assign new_n3865_ = ~new_n3862_ & ~new_n3864_;
  assign new_n3866_ = new_n3859_ & new_n3865_;
  assign new_n3867_ = new_n3854_ & new_n3866_;
  assign new_n3868_ = new_n1295_ & new_n3860_;
  assign new_n3869_ = new_n3829_ & new_n3868_;
  assign new_n3870_ = new_n1300_ & new_n3860_;
  assign new_n3871_ = new_n3829_ & new_n3870_;
  assign new_n3872_ = ~new_n3869_ & ~new_n3871_;
  assign new_n3873_ = A200 & new_n2448_;
  assign new_n3874_ = new_n1284_ & new_n3873_;
  assign new_n3875_ = new_n3829_ & new_n3874_;
  assign new_n3876_ = new_n1291_ & new_n3873_;
  assign new_n3877_ = new_n3829_ & new_n3876_;
  assign new_n3878_ = ~new_n3875_ & ~new_n3877_;
  assign new_n3879_ = new_n3872_ & new_n3878_;
  assign new_n3880_ = A203 & new_n2401_;
  assign new_n3881_ = new_n1284_ & new_n3880_;
  assign new_n3882_ = ~A167 & new_n3016_;
  assign new_n3883_ = new_n1039_ & new_n3882_;
  assign new_n3884_ = new_n3881_ & new_n3883_;
  assign new_n3885_ = new_n1295_ & new_n3873_;
  assign new_n3886_ = new_n3829_ & new_n3885_;
  assign new_n3887_ = new_n1300_ & new_n3873_;
  assign new_n3888_ = new_n3829_ & new_n3887_;
  assign new_n3889_ = ~new_n3886_ & ~new_n3888_;
  assign new_n3890_ = ~new_n3884_ & new_n3889_;
  assign new_n3891_ = new_n3879_ & new_n3890_;
  assign new_n3892_ = new_n3867_ & new_n3891_;
  assign new_n3893_ = new_n1291_ & new_n3880_;
  assign new_n3894_ = new_n3883_ & new_n3893_;
  assign new_n3895_ = new_n1295_ & new_n3880_;
  assign new_n3896_ = new_n3883_ & new_n3895_;
  assign new_n3897_ = ~new_n3894_ & ~new_n3896_;
  assign new_n3898_ = new_n1300_ & new_n3880_;
  assign new_n3899_ = new_n3883_ & new_n3898_;
  assign new_n3900_ = A203 & new_n2417_;
  assign new_n3901_ = new_n1284_ & new_n3900_;
  assign new_n3902_ = new_n3883_ & new_n3901_;
  assign new_n3903_ = ~new_n3899_ & ~new_n3902_;
  assign new_n3904_ = new_n3897_ & new_n3903_;
  assign new_n3905_ = new_n1300_ & new_n3900_;
  assign new_n3906_ = new_n3883_ & new_n3905_;
  assign new_n3907_ = new_n1291_ & new_n3900_;
  assign new_n3908_ = new_n3883_ & new_n3907_;
  assign new_n3909_ = new_n1295_ & new_n3900_;
  assign new_n3910_ = new_n3883_ & new_n3909_;
  assign new_n3911_ = ~new_n3908_ & ~new_n3910_;
  assign new_n3912_ = ~new_n3906_ & new_n3911_;
  assign new_n3913_ = new_n3904_ & new_n3912_;
  assign new_n3914_ = A203 & new_n2435_;
  assign new_n3915_ = new_n1284_ & new_n3914_;
  assign new_n3916_ = new_n3883_ & new_n3915_;
  assign new_n3917_ = new_n1291_ & new_n3914_;
  assign new_n3918_ = new_n3883_ & new_n3917_;
  assign new_n3919_ = ~new_n3916_ & ~new_n3918_;
  assign new_n3920_ = new_n1295_ & new_n3914_;
  assign new_n3921_ = new_n3883_ & new_n3920_;
  assign new_n3922_ = new_n1300_ & new_n3914_;
  assign new_n3923_ = new_n3883_ & new_n3922_;
  assign new_n3924_ = ~new_n3921_ & ~new_n3923_;
  assign new_n3925_ = new_n3919_ & new_n3924_;
  assign new_n3926_ = A203 & new_n2448_;
  assign new_n3927_ = new_n1295_ & new_n3926_;
  assign new_n3928_ = new_n3883_ & new_n3927_;
  assign new_n3929_ = new_n1284_ & new_n3926_;
  assign new_n3930_ = new_n3883_ & new_n3929_;
  assign new_n3931_ = new_n1291_ & new_n3926_;
  assign new_n3932_ = new_n3883_ & new_n3931_;
  assign new_n3933_ = ~new_n3930_ & ~new_n3932_;
  assign new_n3934_ = ~new_n3928_ & new_n3933_;
  assign new_n3935_ = new_n3925_ & new_n3934_;
  assign new_n3936_ = new_n3913_ & new_n3935_;
  assign new_n3937_ = new_n3892_ & new_n3936_;
  assign new_n3938_ = new_n1300_ & new_n3926_;
  assign new_n3939_ = new_n3883_ & new_n3938_;
  assign new_n3940_ = A202 & new_n2401_;
  assign new_n3941_ = new_n1284_ & new_n3940_;
  assign new_n3942_ = new_n3883_ & new_n3941_;
  assign new_n3943_ = ~new_n3939_ & ~new_n3942_;
  assign new_n3944_ = new_n1291_ & new_n3940_;
  assign new_n3945_ = new_n3883_ & new_n3944_;
  assign new_n3946_ = new_n1295_ & new_n3940_;
  assign new_n3947_ = new_n3883_ & new_n3946_;
  assign new_n3948_ = ~new_n3945_ & ~new_n3947_;
  assign new_n3949_ = new_n3943_ & new_n3948_;
  assign new_n3950_ = new_n1300_ & new_n3940_;
  assign new_n3951_ = new_n3883_ & new_n3950_;
  assign new_n3952_ = A202 & new_n2417_;
  assign new_n3953_ = new_n1284_ & new_n3952_;
  assign new_n3954_ = new_n3883_ & new_n3953_;
  assign new_n3955_ = ~new_n3951_ & ~new_n3954_;
  assign new_n3956_ = new_n1291_ & new_n3952_;
  assign new_n3957_ = new_n3883_ & new_n3956_;
  assign new_n3958_ = new_n1295_ & new_n3952_;
  assign new_n3959_ = new_n3883_ & new_n3958_;
  assign new_n3960_ = ~new_n3957_ & ~new_n3959_;
  assign new_n3961_ = new_n3955_ & new_n3960_;
  assign new_n3962_ = new_n3949_ & new_n3961_;
  assign new_n3963_ = new_n1300_ & new_n3952_;
  assign new_n3964_ = new_n3883_ & new_n3963_;
  assign new_n3965_ = A202 & new_n2435_;
  assign new_n3966_ = new_n1284_ & new_n3965_;
  assign new_n3967_ = new_n3883_ & new_n3966_;
  assign new_n3968_ = ~new_n3964_ & ~new_n3967_;
  assign new_n3969_ = new_n1291_ & new_n3965_;
  assign new_n3970_ = new_n3883_ & new_n3969_;
  assign new_n3971_ = new_n1295_ & new_n3965_;
  assign new_n3972_ = new_n3883_ & new_n3971_;
  assign new_n3973_ = ~new_n3970_ & ~new_n3972_;
  assign new_n3974_ = new_n3968_ & new_n3973_;
  assign new_n3975_ = A202 & new_n2448_;
  assign new_n3976_ = new_n1291_ & new_n3975_;
  assign new_n3977_ = new_n3883_ & new_n3976_;
  assign new_n3978_ = new_n1300_ & new_n3965_;
  assign new_n3979_ = new_n3883_ & new_n3978_;
  assign new_n3980_ = new_n1284_ & new_n3975_;
  assign new_n3981_ = new_n3883_ & new_n3980_;
  assign new_n3982_ = ~new_n3979_ & ~new_n3981_;
  assign new_n3983_ = ~new_n3977_ & new_n3982_;
  assign new_n3984_ = new_n3974_ & new_n3983_;
  assign new_n3985_ = new_n3962_ & new_n3984_;
  assign new_n3986_ = new_n1295_ & new_n3975_;
  assign new_n3987_ = new_n3883_ & new_n3986_;
  assign new_n3988_ = new_n1300_ & new_n3975_;
  assign new_n3989_ = new_n3883_ & new_n3988_;
  assign new_n3990_ = ~new_n3987_ & ~new_n3989_;
  assign new_n3991_ = A167 & new_n66_;
  assign new_n3992_ = new_n1039_ & new_n3991_;
  assign new_n3993_ = new_n3776_ & new_n3992_;
  assign new_n3994_ = new_n3784_ & new_n3992_;
  assign new_n3995_ = ~new_n3993_ & ~new_n3994_;
  assign new_n3996_ = new_n3990_ & new_n3995_;
  assign new_n3997_ = new_n3793_ & new_n3992_;
  assign new_n3998_ = new_n3786_ & new_n3992_;
  assign new_n3999_ = new_n3782_ & new_n3992_;
  assign new_n4000_ = ~new_n3998_ & ~new_n3999_;
  assign new_n4001_ = ~new_n3997_ & new_n4000_;
  assign new_n4002_ = new_n3996_ & new_n4001_;
  assign new_n4003_ = new_n3795_ & new_n3992_;
  assign new_n4004_ = new_n3798_ & new_n3992_;
  assign new_n4005_ = ~new_n4003_ & ~new_n4004_;
  assign new_n4006_ = new_n3800_ & new_n3992_;
  assign new_n4007_ = new_n3807_ & new_n3992_;
  assign new_n4008_ = ~new_n4006_ & ~new_n4007_;
  assign new_n4009_ = new_n4005_ & new_n4008_;
  assign new_n4010_ = new_n3814_ & new_n3992_;
  assign new_n4011_ = new_n3809_ & new_n3992_;
  assign new_n4012_ = new_n3805_ & new_n3992_;
  assign new_n4013_ = ~new_n4011_ & ~new_n4012_;
  assign new_n4014_ = ~new_n4010_ & new_n4013_;
  assign new_n4015_ = new_n4009_ & new_n4014_;
  assign new_n4016_ = new_n4002_ & new_n4015_;
  assign new_n4017_ = new_n3985_ & new_n4016_;
  assign new_n4018_ = new_n3937_ & new_n4017_;
  assign new_n4019_ = new_n3817_ & new_n3992_;
  assign new_n4020_ = new_n3820_ & new_n3992_;
  assign new_n4021_ = ~new_n4019_ & ~new_n4020_;
  assign new_n4022_ = new_n3822_ & new_n3992_;
  assign new_n4023_ = new_n3831_ & new_n3992_;
  assign new_n4024_ = ~new_n4022_ & ~new_n4023_;
  assign new_n4025_ = new_n4021_ & new_n4024_;
  assign new_n4026_ = A167 & new_n58_;
  assign new_n4027_ = new_n1039_ & new_n4026_;
  assign new_n4028_ = new_n3833_ & new_n4027_;
  assign new_n4029_ = new_n3827_ & new_n4027_;
  assign new_n4030_ = ~new_n4028_ & ~new_n4029_;
  assign new_n4031_ = new_n3843_ & new_n4027_;
  assign new_n4032_ = new_n3845_ & new_n4027_;
  assign new_n4033_ = ~new_n4031_ & ~new_n4032_;
  assign new_n4034_ = new_n4030_ & new_n4033_;
  assign new_n4035_ = new_n4025_ & new_n4034_;
  assign new_n4036_ = new_n3849_ & new_n4027_;
  assign new_n4037_ = new_n3851_ & new_n4027_;
  assign new_n4038_ = ~new_n4036_ & ~new_n4037_;
  assign new_n4039_ = new_n3855_ & new_n4027_;
  assign new_n4040_ = new_n3857_ & new_n4027_;
  assign new_n4041_ = ~new_n4039_ & ~new_n4040_;
  assign new_n4042_ = new_n4038_ & new_n4041_;
  assign new_n4043_ = new_n3868_ & new_n4027_;
  assign new_n4044_ = new_n3861_ & new_n4027_;
  assign new_n4045_ = new_n3863_ & new_n4027_;
  assign new_n4046_ = ~new_n4044_ & ~new_n4045_;
  assign new_n4047_ = ~new_n4043_ & new_n4046_;
  assign new_n4048_ = new_n4042_ & new_n4047_;
  assign new_n4049_ = new_n4035_ & new_n4048_;
  assign new_n4050_ = new_n3870_ & new_n4027_;
  assign new_n4051_ = new_n3874_ & new_n4027_;
  assign new_n4052_ = ~new_n4050_ & ~new_n4051_;
  assign new_n4053_ = new_n3876_ & new_n4027_;
  assign new_n4054_ = new_n3885_ & new_n4027_;
  assign new_n4055_ = ~new_n4053_ & ~new_n4054_;
  assign new_n4056_ = new_n4052_ & new_n4055_;
  assign new_n4057_ = A167 & new_n3192_;
  assign new_n4058_ = new_n1039_ & new_n4057_;
  assign new_n4059_ = new_n3893_ & new_n4058_;
  assign new_n4060_ = new_n3887_ & new_n4027_;
  assign new_n4061_ = new_n3881_ & new_n4058_;
  assign new_n4062_ = ~new_n4060_ & ~new_n4061_;
  assign new_n4063_ = ~new_n4059_ & new_n4062_;
  assign new_n4064_ = new_n4056_ & new_n4063_;
  assign new_n4065_ = new_n3895_ & new_n4058_;
  assign new_n4066_ = new_n3898_ & new_n4058_;
  assign new_n4067_ = ~new_n4065_ & ~new_n4066_;
  assign new_n4068_ = new_n3901_ & new_n4058_;
  assign new_n4069_ = new_n3907_ & new_n4058_;
  assign new_n4070_ = ~new_n4068_ & ~new_n4069_;
  assign new_n4071_ = new_n4067_ & new_n4070_;
  assign new_n4072_ = new_n3915_ & new_n4058_;
  assign new_n4073_ = new_n3909_ & new_n4058_;
  assign new_n4074_ = new_n3905_ & new_n4058_;
  assign new_n4075_ = ~new_n4073_ & ~new_n4074_;
  assign new_n4076_ = ~new_n4072_ & new_n4075_;
  assign new_n4077_ = new_n4071_ & new_n4076_;
  assign new_n4078_ = new_n4064_ & new_n4077_;
  assign new_n4079_ = new_n4049_ & new_n4078_;
  assign new_n4080_ = new_n3917_ & new_n4058_;
  assign new_n4081_ = new_n3920_ & new_n4058_;
  assign new_n4082_ = ~new_n4080_ & ~new_n4081_;
  assign new_n4083_ = new_n3922_ & new_n4058_;
  assign new_n4084_ = new_n3929_ & new_n4058_;
  assign new_n4085_ = ~new_n4083_ & ~new_n4084_;
  assign new_n4086_ = new_n4082_ & new_n4085_;
  assign new_n4087_ = new_n3931_ & new_n4058_;
  assign new_n4088_ = new_n3927_ & new_n4058_;
  assign new_n4089_ = ~new_n4087_ & ~new_n4088_;
  assign new_n4090_ = new_n3938_ & new_n4058_;
  assign new_n4091_ = new_n3941_ & new_n4058_;
  assign new_n4092_ = ~new_n4090_ & ~new_n4091_;
  assign new_n4093_ = new_n4089_ & new_n4092_;
  assign new_n4094_ = new_n4086_ & new_n4093_;
  assign new_n4095_ = new_n3944_ & new_n4058_;
  assign new_n4096_ = new_n3946_ & new_n4058_;
  assign new_n4097_ = ~new_n4095_ & ~new_n4096_;
  assign new_n4098_ = new_n3950_ & new_n4058_;
  assign new_n4099_ = new_n3953_ & new_n4058_;
  assign new_n4100_ = ~new_n4098_ & ~new_n4099_;
  assign new_n4101_ = new_n4097_ & new_n4100_;
  assign new_n4102_ = new_n3963_ & new_n4058_;
  assign new_n4103_ = new_n3956_ & new_n4058_;
  assign new_n4104_ = new_n3958_ & new_n4058_;
  assign new_n4105_ = ~new_n4103_ & ~new_n4104_;
  assign new_n4106_ = ~new_n4102_ & new_n4105_;
  assign new_n4107_ = new_n4101_ & new_n4106_;
  assign new_n4108_ = new_n4094_ & new_n4107_;
  assign new_n4109_ = new_n3966_ & new_n4058_;
  assign new_n4110_ = new_n3969_ & new_n4058_;
  assign new_n4111_ = ~new_n4109_ & ~new_n4110_;
  assign new_n4112_ = new_n3971_ & new_n4058_;
  assign new_n4113_ = new_n3978_ & new_n4058_;
  assign new_n4114_ = ~new_n4112_ & ~new_n4113_;
  assign new_n4115_ = new_n4111_ & new_n4114_;
  assign new_n4116_ = new_n3986_ & new_n4058_;
  assign new_n4117_ = new_n3980_ & new_n4058_;
  assign new_n4118_ = new_n3976_ & new_n4058_;
  assign new_n4119_ = ~new_n4117_ & ~new_n4118_;
  assign new_n4120_ = ~new_n4116_ & new_n4119_;
  assign new_n4121_ = new_n4115_ & new_n4120_;
  assign new_n4122_ = new_n3988_ & new_n4058_;
  assign new_n4123_ = A265 & ~A200;
  assign new_n4124_ = ~A199 & new_n4123_;
  assign new_n4125_ = new_n1485_ & new_n4124_;
  assign new_n4126_ = new_n2747_ & new_n4125_;
  assign new_n4127_ = ~new_n4122_ & ~new_n4126_;
  assign new_n4128_ = ~A265 & ~A200;
  assign new_n4129_ = ~A199 & new_n4128_;
  assign new_n4130_ = new_n1485_ & new_n4129_;
  assign new_n4131_ = new_n2755_ & new_n4130_;
  assign new_n4132_ = A199 & new_n134_;
  assign new_n4133_ = new_n1485_ & new_n4132_;
  assign new_n4134_ = new_n3881_ & new_n4133_;
  assign new_n4135_ = ~new_n4131_ & ~new_n4134_;
  assign new_n4136_ = new_n4127_ & new_n4135_;
  assign new_n4137_ = new_n3898_ & new_n4133_;
  assign new_n4138_ = new_n3893_ & new_n4133_;
  assign new_n4139_ = new_n3895_ & new_n4133_;
  assign new_n4140_ = ~new_n4138_ & ~new_n4139_;
  assign new_n4141_ = ~new_n4137_ & new_n4140_;
  assign new_n4142_ = new_n4136_ & new_n4141_;
  assign new_n4143_ = new_n4121_ & new_n4142_;
  assign new_n4144_ = new_n4108_ & new_n4143_;
  assign new_n4145_ = new_n4079_ & new_n4144_;
  assign new_n4146_ = new_n4018_ & new_n4145_;
  assign new_n4147_ = new_n3901_ & new_n4133_;
  assign new_n4148_ = new_n3907_ & new_n4133_;
  assign new_n4149_ = ~new_n4147_ & ~new_n4148_;
  assign new_n4150_ = new_n3909_ & new_n4133_;
  assign new_n4151_ = new_n3905_ & new_n4133_;
  assign new_n4152_ = ~new_n4150_ & ~new_n4151_;
  assign new_n4153_ = new_n4149_ & new_n4152_;
  assign new_n4154_ = new_n3915_ & new_n4133_;
  assign new_n4155_ = new_n3917_ & new_n4133_;
  assign new_n4156_ = ~new_n4154_ & ~new_n4155_;
  assign new_n4157_ = new_n3920_ & new_n4133_;
  assign new_n4158_ = new_n3922_ & new_n4133_;
  assign new_n4159_ = ~new_n4157_ & ~new_n4158_;
  assign new_n4160_ = new_n4156_ & new_n4159_;
  assign new_n4161_ = new_n4153_ & new_n4160_;
  assign new_n4162_ = new_n3929_ & new_n4133_;
  assign new_n4163_ = new_n3931_ & new_n4133_;
  assign new_n4164_ = ~new_n4162_ & ~new_n4163_;
  assign new_n4165_ = new_n3927_ & new_n4133_;
  assign new_n4166_ = new_n3938_ & new_n4133_;
  assign new_n4167_ = ~new_n4165_ & ~new_n4166_;
  assign new_n4168_ = new_n4164_ & new_n4167_;
  assign new_n4169_ = new_n3946_ & new_n4133_;
  assign new_n4170_ = new_n3941_ & new_n4133_;
  assign new_n4171_ = new_n3944_ & new_n4133_;
  assign new_n4172_ = ~new_n4170_ & ~new_n4171_;
  assign new_n4173_ = ~new_n4169_ & new_n4172_;
  assign new_n4174_ = new_n4168_ & new_n4173_;
  assign new_n4175_ = new_n4161_ & new_n4174_;
  assign new_n4176_ = new_n3950_ & new_n4133_;
  assign new_n4177_ = new_n3953_ & new_n4133_;
  assign new_n4178_ = ~new_n4176_ & ~new_n4177_;
  assign new_n4179_ = new_n3956_ & new_n4133_;
  assign new_n4180_ = new_n3958_ & new_n4133_;
  assign new_n4181_ = ~new_n4179_ & ~new_n4180_;
  assign new_n4182_ = new_n4178_ & new_n4181_;
  assign new_n4183_ = new_n3969_ & new_n4133_;
  assign new_n4184_ = new_n3963_ & new_n4133_;
  assign new_n4185_ = new_n3966_ & new_n4133_;
  assign new_n4186_ = ~new_n4184_ & ~new_n4185_;
  assign new_n4187_ = ~new_n4183_ & new_n4186_;
  assign new_n4188_ = new_n4182_ & new_n4187_;
  assign new_n4189_ = new_n3971_ & new_n4133_;
  assign new_n4190_ = new_n3978_ & new_n4133_;
  assign new_n4191_ = ~new_n4189_ & ~new_n4190_;
  assign new_n4192_ = new_n3980_ & new_n4133_;
  assign new_n4193_ = new_n3976_ & new_n4133_;
  assign new_n4194_ = ~new_n4192_ & ~new_n4193_;
  assign new_n4195_ = new_n4191_ & new_n4194_;
  assign new_n4196_ = ~A199 & new_n182_;
  assign new_n4197_ = new_n1485_ & new_n4196_;
  assign new_n4198_ = new_n3881_ & new_n4197_;
  assign new_n4199_ = new_n3986_ & new_n4133_;
  assign new_n4200_ = new_n3988_ & new_n4133_;
  assign new_n4201_ = ~new_n4199_ & ~new_n4200_;
  assign new_n4202_ = ~new_n4198_ & new_n4201_;
  assign new_n4203_ = new_n4195_ & new_n4202_;
  assign new_n4204_ = new_n4188_ & new_n4203_;
  assign new_n4205_ = new_n4175_ & new_n4204_;
  assign new_n4206_ = new_n3893_ & new_n4197_;
  assign new_n4207_ = new_n3895_ & new_n4197_;
  assign new_n4208_ = ~new_n4206_ & ~new_n4207_;
  assign new_n4209_ = new_n3898_ & new_n4197_;
  assign new_n4210_ = new_n3901_ & new_n4197_;
  assign new_n4211_ = ~new_n4209_ & ~new_n4210_;
  assign new_n4212_ = new_n4208_ & new_n4211_;
  assign new_n4213_ = new_n3907_ & new_n4197_;
  assign new_n4214_ = new_n3909_ & new_n4197_;
  assign new_n4215_ = ~new_n4213_ & ~new_n4214_;
  assign new_n4216_ = new_n3905_ & new_n4197_;
  assign new_n4217_ = new_n3915_ & new_n4197_;
  assign new_n4218_ = ~new_n4216_ & ~new_n4217_;
  assign new_n4219_ = new_n4215_ & new_n4218_;
  assign new_n4220_ = new_n4212_ & new_n4219_;
  assign new_n4221_ = new_n3917_ & new_n4197_;
  assign new_n4222_ = new_n3920_ & new_n4197_;
  assign new_n4223_ = ~new_n4221_ & ~new_n4222_;
  assign new_n4224_ = new_n3922_ & new_n4197_;
  assign new_n4225_ = new_n3929_ & new_n4197_;
  assign new_n4226_ = ~new_n4224_ & ~new_n4225_;
  assign new_n4227_ = new_n4223_ & new_n4226_;
  assign new_n4228_ = new_n3938_ & new_n4197_;
  assign new_n4229_ = new_n3931_ & new_n4197_;
  assign new_n4230_ = new_n3927_ & new_n4197_;
  assign new_n4231_ = ~new_n4229_ & ~new_n4230_;
  assign new_n4232_ = ~new_n4228_ & new_n4231_;
  assign new_n4233_ = new_n4227_ & new_n4232_;
  assign new_n4234_ = new_n4220_ & new_n4233_;
  assign new_n4235_ = new_n3941_ & new_n4197_;
  assign new_n4236_ = new_n3944_ & new_n4197_;
  assign new_n4237_ = ~new_n4235_ & ~new_n4236_;
  assign new_n4238_ = new_n3946_ & new_n4197_;
  assign new_n4239_ = new_n3950_ & new_n4197_;
  assign new_n4240_ = ~new_n4238_ & ~new_n4239_;
  assign new_n4241_ = new_n4237_ & new_n4240_;
  assign new_n4242_ = new_n3958_ & new_n4197_;
  assign new_n4243_ = new_n3953_ & new_n4197_;
  assign new_n4244_ = new_n3956_ & new_n4197_;
  assign new_n4245_ = ~new_n4243_ & ~new_n4244_;
  assign new_n4246_ = ~new_n4242_ & new_n4245_;
  assign new_n4247_ = new_n4241_ & new_n4246_;
  assign new_n4248_ = new_n3963_ & new_n4197_;
  assign new_n4249_ = new_n3966_ & new_n4197_;
  assign new_n4250_ = ~new_n4248_ & ~new_n4249_;
  assign new_n4251_ = new_n3969_ & new_n4197_;
  assign new_n4252_ = new_n3971_ & new_n4197_;
  assign new_n4253_ = ~new_n4251_ & ~new_n4252_;
  assign new_n4254_ = new_n4250_ & new_n4253_;
  assign new_n4255_ = new_n3976_ & new_n4197_;
  assign new_n4256_ = new_n3978_ & new_n4197_;
  assign new_n4257_ = new_n3980_ & new_n4197_;
  assign new_n4258_ = ~new_n4256_ & ~new_n4257_;
  assign new_n4259_ = ~new_n4255_ & new_n4258_;
  assign new_n4260_ = new_n4254_ & new_n4259_;
  assign new_n4261_ = new_n4247_ & new_n4260_;
  assign new_n4262_ = new_n4234_ & new_n4261_;
  assign new_n4263_ = new_n4205_ & new_n4262_;
  assign new_n4264_ = new_n3986_ & new_n4197_;
  assign new_n4265_ = new_n3988_ & new_n4197_;
  assign new_n4266_ = ~new_n4264_ & ~new_n4265_;
  assign new_n4267_ = A265 & A200;
  assign new_n4268_ = A199 & new_n4267_;
  assign new_n4269_ = new_n1485_ & new_n4268_;
  assign new_n4270_ = new_n2747_ & new_n4269_;
  assign new_n4271_ = ~A265 & A200;
  assign new_n4272_ = A199 & new_n4271_;
  assign new_n4273_ = new_n1485_ & new_n4272_;
  assign new_n4274_ = new_n2755_ & new_n4273_;
  assign new_n4275_ = ~new_n4270_ & ~new_n4274_;
  assign new_n4276_ = new_n4266_ & new_n4275_;
  assign new_n4277_ = ~A201 & new_n140_;
  assign new_n4278_ = new_n1485_ & new_n4277_;
  assign new_n4279_ = new_n2747_ & new_n4278_;
  assign new_n4280_ = ~A201 & new_n131_;
  assign new_n4281_ = new_n1485_ & new_n4280_;
  assign new_n4282_ = new_n2755_ & new_n4281_;
  assign new_n4283_ = ~new_n4279_ & ~new_n4282_;
  assign new_n4284_ = ~A201 & new_n147_;
  assign new_n4285_ = new_n1485_ & new_n4284_;
  assign new_n4286_ = new_n2747_ & new_n4285_;
  assign new_n4287_ = ~A201 & new_n151_;
  assign new_n4288_ = new_n1485_ & new_n4287_;
  assign new_n4289_ = new_n2755_ & new_n4288_;
  assign new_n4290_ = ~new_n4286_ & ~new_n4289_;
  assign new_n4291_ = new_n4283_ & new_n4290_;
  assign new_n4292_ = new_n4276_ & new_n4291_;
  assign new_n4293_ = A265 & new_n31_;
  assign new_n4294_ = new_n373_ & new_n4293_;
  assign new_n4295_ = A201 & new_n79_;
  assign new_n4296_ = new_n1485_ & new_n4295_;
  assign new_n4297_ = new_n4294_ & new_n4296_;
  assign new_n4298_ = new_n376_ & new_n4293_;
  assign new_n4299_ = new_n4296_ & new_n4298_;
  assign new_n4300_ = ~new_n4297_ & ~new_n4299_;
  assign new_n4301_ = new_n387_ & new_n4293_;
  assign new_n4302_ = new_n4296_ & new_n4301_;
  assign new_n4303_ = new_n390_ & new_n4293_;
  assign new_n4304_ = new_n4296_ & new_n4303_;
  assign new_n4305_ = ~new_n4302_ & ~new_n4304_;
  assign new_n4306_ = new_n4300_ & new_n4305_;
  assign new_n4307_ = ~A265 & new_n44_;
  assign new_n4308_ = new_n373_ & new_n4307_;
  assign new_n4309_ = new_n4296_ & new_n4308_;
  assign new_n4310_ = A265 & new_n383_;
  assign new_n4311_ = new_n382_ & new_n4310_;
  assign new_n4312_ = new_n4296_ & new_n4311_;
  assign new_n4313_ = new_n397_ & new_n4310_;
  assign new_n4314_ = new_n4296_ & new_n4313_;
  assign new_n4315_ = ~new_n4312_ & ~new_n4314_;
  assign new_n4316_ = ~new_n4309_ & new_n4315_;
  assign new_n4317_ = new_n4306_ & new_n4316_;
  assign new_n4318_ = new_n4292_ & new_n4317_;
  assign new_n4319_ = new_n376_ & new_n4307_;
  assign new_n4320_ = new_n4296_ & new_n4319_;
  assign new_n4321_ = new_n387_ & new_n4307_;
  assign new_n4322_ = new_n4296_ & new_n4321_;
  assign new_n4323_ = ~new_n4320_ & ~new_n4322_;
  assign new_n4324_ = new_n390_ & new_n4307_;
  assign new_n4325_ = new_n4296_ & new_n4324_;
  assign new_n4326_ = ~A265 & new_n409_;
  assign new_n4327_ = new_n382_ & new_n4326_;
  assign new_n4328_ = new_n4296_ & new_n4327_;
  assign new_n4329_ = ~new_n4325_ & ~new_n4328_;
  assign new_n4330_ = new_n4323_ & new_n4329_;
  assign new_n4331_ = new_n36_ & new_n1557_;
  assign new_n4332_ = new_n2410_ & new_n4331_;
  assign new_n4333_ = new_n397_ & new_n4326_;
  assign new_n4334_ = new_n4296_ & new_n4333_;
  assign new_n4335_ = new_n2403_ & new_n4331_;
  assign new_n4336_ = ~new_n4334_ & ~new_n4335_;
  assign new_n4337_ = ~new_n4332_ & new_n4336_;
  assign new_n4338_ = new_n4330_ & new_n4337_;
  assign new_n4339_ = new_n2412_ & new_n4331_;
  assign new_n4340_ = new_n2415_ & new_n4331_;
  assign new_n4341_ = ~new_n4339_ & ~new_n4340_;
  assign new_n4342_ = new_n2419_ & new_n4331_;
  assign new_n4343_ = new_n2425_ & new_n4331_;
  assign new_n4344_ = ~new_n4342_ & ~new_n4343_;
  assign new_n4345_ = new_n4341_ & new_n4344_;
  assign new_n4346_ = new_n2437_ & new_n4331_;
  assign new_n4347_ = new_n2427_ & new_n4331_;
  assign new_n4348_ = new_n2423_ & new_n4331_;
  assign new_n4349_ = ~new_n4347_ & ~new_n4348_;
  assign new_n4350_ = ~new_n4346_ & new_n4349_;
  assign new_n4351_ = new_n4345_ & new_n4350_;
  assign new_n4352_ = new_n4338_ & new_n4351_;
  assign new_n4353_ = new_n4318_ & new_n4352_;
  assign new_n4354_ = new_n2439_ & new_n4331_;
  assign new_n4355_ = new_n2442_ & new_n4331_;
  assign new_n4356_ = ~new_n4354_ & ~new_n4355_;
  assign new_n4357_ = new_n2444_ & new_n4331_;
  assign new_n4358_ = new_n2450_ & new_n4331_;
  assign new_n4359_ = ~new_n4357_ & ~new_n4358_;
  assign new_n4360_ = new_n4356_ & new_n4359_;
  assign new_n4361_ = new_n2457_ & new_n4331_;
  assign new_n4362_ = new_n2452_ & new_n4331_;
  assign new_n4363_ = new_n2455_ & new_n4331_;
  assign new_n4364_ = ~new_n4362_ & ~new_n4363_;
  assign new_n4365_ = ~new_n4361_ & new_n4364_;
  assign new_n4366_ = new_n4360_ & new_n4365_;
  assign new_n4367_ = ~A200 & new_n781_;
  assign new_n4368_ = new_n1557_ & new_n4367_;
  assign new_n4369_ = new_n2291_ & new_n4368_;
  assign new_n4370_ = new_n2294_ & new_n4368_;
  assign new_n4371_ = ~new_n4369_ & ~new_n4370_;
  assign new_n4372_ = new_n2299_ & new_n4368_;
  assign new_n4373_ = new_n2302_ & new_n4368_;
  assign new_n4374_ = ~new_n4372_ & ~new_n4373_;
  assign new_n4375_ = new_n4371_ & new_n4374_;
  assign new_n4376_ = new_n2315_ & new_n4368_;
  assign new_n4377_ = new_n2306_ & new_n4368_;
  assign new_n4378_ = new_n2309_ & new_n4368_;
  assign new_n4379_ = ~new_n4377_ & ~new_n4378_;
  assign new_n4380_ = ~new_n4376_ & new_n4379_;
  assign new_n4381_ = new_n4375_ & new_n4380_;
  assign new_n4382_ = new_n4366_ & new_n4381_;
  assign new_n4383_ = new_n2318_ & new_n4368_;
  assign new_n4384_ = new_n2322_ & new_n4368_;
  assign new_n4385_ = ~new_n4383_ & ~new_n4384_;
  assign new_n4386_ = new_n2324_ & new_n4368_;
  assign new_n4387_ = new_n2329_ & new_n4368_;
  assign new_n4388_ = ~new_n4386_ & ~new_n4387_;
  assign new_n4389_ = new_n4385_ & new_n4388_;
  assign new_n4390_ = ~A200 & new_n791_;
  assign new_n4391_ = new_n1557_ & new_n4390_;
  assign new_n4392_ = new_n2294_ & new_n4391_;
  assign new_n4393_ = new_n2331_ & new_n4368_;
  assign new_n4394_ = new_n2291_ & new_n4391_;
  assign new_n4395_ = ~new_n4393_ & ~new_n4394_;
  assign new_n4396_ = ~new_n4392_ & new_n4395_;
  assign new_n4397_ = new_n4389_ & new_n4396_;
  assign new_n4398_ = new_n2299_ & new_n4391_;
  assign new_n4399_ = new_n2302_ & new_n4391_;
  assign new_n4400_ = ~new_n4398_ & ~new_n4399_;
  assign new_n4401_ = new_n2306_ & new_n4391_;
  assign new_n4402_ = new_n2309_ & new_n4391_;
  assign new_n4403_ = ~new_n4401_ & ~new_n4402_;
  assign new_n4404_ = new_n4400_ & new_n4403_;
  assign new_n4405_ = new_n2322_ & new_n4391_;
  assign new_n4406_ = new_n2315_ & new_n4391_;
  assign new_n4407_ = new_n2318_ & new_n4391_;
  assign new_n4408_ = ~new_n4406_ & ~new_n4407_;
  assign new_n4409_ = ~new_n4405_ & new_n4408_;
  assign new_n4410_ = new_n4404_ & new_n4409_;
  assign new_n4411_ = new_n4397_ & new_n4410_;
  assign new_n4412_ = new_n4382_ & new_n4411_;
  assign new_n4413_ = new_n4353_ & new_n4412_;
  assign new_n4414_ = new_n4263_ & new_n4413_;
  assign new_n4415_ = new_n4146_ & new_n4414_;
  assign new_n4416_ = new_n3842_ & new_n4415_;
  assign new_n4417_ = new_n3339_ & new_n4416_;
  assign new_n4418_ = new_n2284_ & new_n4417_;
  assign new_n4419_ = new_n2324_ & new_n4391_;
  assign new_n4420_ = new_n2329_ & new_n4391_;
  assign new_n4421_ = ~new_n4419_ & ~new_n4420_;
  assign new_n4422_ = new_n2331_ & new_n4391_;
  assign new_n4423_ = new_n50_ & new_n1563_;
  assign new_n4424_ = new_n2403_ & new_n4423_;
  assign new_n4425_ = ~new_n4422_ & ~new_n4424_;
  assign new_n4426_ = new_n4421_ & new_n4425_;
  assign new_n4427_ = new_n2410_ & new_n4423_;
  assign new_n4428_ = new_n2412_ & new_n4423_;
  assign new_n4429_ = ~new_n4427_ & ~new_n4428_;
  assign new_n4430_ = new_n2415_ & new_n4423_;
  assign new_n4431_ = new_n2419_ & new_n4423_;
  assign new_n4432_ = ~new_n4430_ & ~new_n4431_;
  assign new_n4433_ = new_n4429_ & new_n4432_;
  assign new_n4434_ = new_n4426_ & new_n4433_;
  assign new_n4435_ = new_n2425_ & new_n4423_;
  assign new_n4436_ = new_n2427_ & new_n4423_;
  assign new_n4437_ = ~new_n4435_ & ~new_n4436_;
  assign new_n4438_ = new_n2423_ & new_n4423_;
  assign new_n4439_ = new_n2437_ & new_n4423_;
  assign new_n4440_ = ~new_n4438_ & ~new_n4439_;
  assign new_n4441_ = new_n4437_ & new_n4440_;
  assign new_n4442_ = new_n2444_ & new_n4423_;
  assign new_n4443_ = new_n2439_ & new_n4423_;
  assign new_n4444_ = new_n2442_ & new_n4423_;
  assign new_n4445_ = ~new_n4443_ & ~new_n4444_;
  assign new_n4446_ = ~new_n4442_ & new_n4445_;
  assign new_n4447_ = new_n4441_ & new_n4446_;
  assign new_n4448_ = new_n4434_ & new_n4447_;
  assign new_n4449_ = new_n2450_ & new_n4423_;
  assign new_n4450_ = new_n2452_ & new_n4423_;
  assign new_n4451_ = ~new_n4449_ & ~new_n4450_;
  assign new_n4452_ = new_n2455_ & new_n4423_;
  assign new_n4453_ = new_n2457_ & new_n4423_;
  assign new_n4454_ = ~new_n4452_ & ~new_n4453_;
  assign new_n4455_ = new_n4451_ & new_n4454_;
  assign new_n4456_ = A200 & new_n781_;
  assign new_n4457_ = new_n1563_ & new_n4456_;
  assign new_n4458_ = new_n2299_ & new_n4457_;
  assign new_n4459_ = new_n2291_ & new_n4457_;
  assign new_n4460_ = new_n2294_ & new_n4457_;
  assign new_n4461_ = ~new_n4459_ & ~new_n4460_;
  assign new_n4462_ = ~new_n4458_ & new_n4461_;
  assign new_n4463_ = new_n4455_ & new_n4462_;
  assign new_n4464_ = new_n2302_ & new_n4457_;
  assign new_n4465_ = new_n2306_ & new_n4457_;
  assign new_n4466_ = ~new_n4464_ & ~new_n4465_;
  assign new_n4467_ = new_n2309_ & new_n4457_;
  assign new_n4468_ = new_n2315_ & new_n4457_;
  assign new_n4469_ = ~new_n4467_ & ~new_n4468_;
  assign new_n4470_ = new_n4466_ & new_n4469_;
  assign new_n4471_ = new_n2324_ & new_n4457_;
  assign new_n4472_ = new_n2318_ & new_n4457_;
  assign new_n4473_ = new_n2322_ & new_n4457_;
  assign new_n4474_ = ~new_n4472_ & ~new_n4473_;
  assign new_n4475_ = ~new_n4471_ & new_n4474_;
  assign new_n4476_ = new_n4470_ & new_n4475_;
  assign new_n4477_ = new_n4463_ & new_n4476_;
  assign new_n4478_ = new_n4448_ & new_n4477_;
  assign new_n4479_ = new_n2329_ & new_n4457_;
  assign new_n4480_ = new_n2331_ & new_n4457_;
  assign new_n4481_ = ~new_n4479_ & ~new_n4480_;
  assign new_n4482_ = A200 & new_n791_;
  assign new_n4483_ = new_n1563_ & new_n4482_;
  assign new_n4484_ = new_n2291_ & new_n4483_;
  assign new_n4485_ = new_n2294_ & new_n4483_;
  assign new_n4486_ = ~new_n4484_ & ~new_n4485_;
  assign new_n4487_ = new_n4481_ & new_n4486_;
  assign new_n4488_ = new_n2299_ & new_n4483_;
  assign new_n4489_ = new_n2302_ & new_n4483_;
  assign new_n4490_ = ~new_n4488_ & ~new_n4489_;
  assign new_n4491_ = new_n2306_ & new_n4483_;
  assign new_n4492_ = new_n2309_ & new_n4483_;
  assign new_n4493_ = ~new_n4491_ & ~new_n4492_;
  assign new_n4494_ = new_n4490_ & new_n4493_;
  assign new_n4495_ = new_n4487_ & new_n4494_;
  assign new_n4496_ = new_n2315_ & new_n4483_;
  assign new_n4497_ = new_n2318_ & new_n4483_;
  assign new_n4498_ = ~new_n4496_ & ~new_n4497_;
  assign new_n4499_ = new_n2322_ & new_n4483_;
  assign new_n4500_ = new_n2324_ & new_n4483_;
  assign new_n4501_ = ~new_n4499_ & ~new_n4500_;
  assign new_n4502_ = new_n4498_ & new_n4501_;
  assign new_n4503_ = ~A202 & new_n32_;
  assign new_n4504_ = A201 & ~A168;
  assign new_n4505_ = A169 & new_n4504_;
  assign new_n4506_ = new_n4503_ & new_n4505_;
  assign new_n4507_ = new_n2747_ & new_n4506_;
  assign new_n4508_ = new_n2329_ & new_n4483_;
  assign new_n4509_ = new_n2331_ & new_n4483_;
  assign new_n4510_ = ~new_n4508_ & ~new_n4509_;
  assign new_n4511_ = ~new_n4507_ & new_n4510_;
  assign new_n4512_ = new_n4502_ & new_n4511_;
  assign new_n4513_ = new_n4495_ & new_n4512_;
  assign new_n4514_ = ~A202 & new_n45_;
  assign new_n4515_ = new_n4505_ & new_n4514_;
  assign new_n4516_ = new_n2755_ & new_n4515_;
  assign new_n4517_ = A166 & new_n1036_;
  assign new_n4518_ = new_n1571_ & new_n4517_;
  assign new_n4519_ = new_n2291_ & new_n4518_;
  assign new_n4520_ = ~new_n4516_ & ~new_n4519_;
  assign new_n4521_ = new_n2294_ & new_n4518_;
  assign new_n4522_ = new_n2299_ & new_n4518_;
  assign new_n4523_ = ~new_n4521_ & ~new_n4522_;
  assign new_n4524_ = new_n4520_ & new_n4523_;
  assign new_n4525_ = new_n2309_ & new_n4518_;
  assign new_n4526_ = new_n2302_ & new_n4518_;
  assign new_n4527_ = new_n2306_ & new_n4518_;
  assign new_n4528_ = ~new_n4526_ & ~new_n4527_;
  assign new_n4529_ = ~new_n4525_ & new_n4528_;
  assign new_n4530_ = new_n4524_ & new_n4529_;
  assign new_n4531_ = new_n2315_ & new_n4518_;
  assign new_n4532_ = new_n2318_ & new_n4518_;
  assign new_n4533_ = ~new_n4531_ & ~new_n4532_;
  assign new_n4534_ = new_n2322_ & new_n4518_;
  assign new_n4535_ = new_n2324_ & new_n4518_;
  assign new_n4536_ = ~new_n4534_ & ~new_n4535_;
  assign new_n4537_ = new_n4533_ & new_n4536_;
  assign new_n4538_ = A166 & new_n1213_;
  assign new_n4539_ = new_n1571_ & new_n4538_;
  assign new_n4540_ = new_n2291_ & new_n4539_;
  assign new_n4541_ = new_n2329_ & new_n4518_;
  assign new_n4542_ = new_n2331_ & new_n4518_;
  assign new_n4543_ = ~new_n4541_ & ~new_n4542_;
  assign new_n4544_ = ~new_n4540_ & new_n4543_;
  assign new_n4545_ = new_n4537_ & new_n4544_;
  assign new_n4546_ = new_n4530_ & new_n4545_;
  assign new_n4547_ = new_n4513_ & new_n4546_;
  assign new_n4548_ = new_n4478_ & new_n4547_;
  assign new_n4549_ = new_n2294_ & new_n4539_;
  assign new_n4550_ = new_n2299_ & new_n4539_;
  assign new_n4551_ = ~new_n4549_ & ~new_n4550_;
  assign new_n4552_ = new_n2302_ & new_n4539_;
  assign new_n4553_ = new_n2306_ & new_n4539_;
  assign new_n4554_ = ~new_n4552_ & ~new_n4553_;
  assign new_n4555_ = new_n4551_ & new_n4554_;
  assign new_n4556_ = new_n2309_ & new_n4539_;
  assign new_n4557_ = new_n2315_ & new_n4539_;
  assign new_n4558_ = ~new_n4556_ & ~new_n4557_;
  assign new_n4559_ = new_n2318_ & new_n4539_;
  assign new_n4560_ = new_n2322_ & new_n4539_;
  assign new_n4561_ = ~new_n4559_ & ~new_n4560_;
  assign new_n4562_ = new_n4558_ & new_n4561_;
  assign new_n4563_ = new_n4555_ & new_n4562_;
  assign new_n4564_ = new_n2324_ & new_n4539_;
  assign new_n4565_ = new_n2329_ & new_n4539_;
  assign new_n4566_ = ~new_n4564_ & ~new_n4565_;
  assign new_n4567_ = new_n2331_ & new_n4539_;
  assign new_n4568_ = A166 & new_n1219_;
  assign new_n4569_ = new_n1571_ & new_n4568_;
  assign new_n4570_ = new_n2291_ & new_n4569_;
  assign new_n4571_ = ~new_n4567_ & ~new_n4570_;
  assign new_n4572_ = new_n4566_ & new_n4571_;
  assign new_n4573_ = new_n2302_ & new_n4569_;
  assign new_n4574_ = new_n2294_ & new_n4569_;
  assign new_n4575_ = new_n2299_ & new_n4569_;
  assign new_n4576_ = ~new_n4574_ & ~new_n4575_;
  assign new_n4577_ = ~new_n4573_ & new_n4576_;
  assign new_n4578_ = new_n4572_ & new_n4577_;
  assign new_n4579_ = new_n4563_ & new_n4578_;
  assign new_n4580_ = new_n2306_ & new_n4569_;
  assign new_n4581_ = new_n2309_ & new_n4569_;
  assign new_n4582_ = ~new_n4580_ & ~new_n4581_;
  assign new_n4583_ = new_n2315_ & new_n4569_;
  assign new_n4584_ = new_n2318_ & new_n4569_;
  assign new_n4585_ = ~new_n4583_ & ~new_n4584_;
  assign new_n4586_ = new_n4582_ & new_n4585_;
  assign new_n4587_ = new_n2329_ & new_n4569_;
  assign new_n4588_ = new_n2322_ & new_n4569_;
  assign new_n4589_ = new_n2324_ & new_n4569_;
  assign new_n4590_ = ~new_n4588_ & ~new_n4589_;
  assign new_n4591_ = ~new_n4587_ & new_n4590_;
  assign new_n4592_ = new_n4586_ & new_n4591_;
  assign new_n4593_ = new_n2331_ & new_n4569_;
  assign new_n4594_ = A166 & new_n1225_;
  assign new_n4595_ = new_n1571_ & new_n4594_;
  assign new_n4596_ = new_n2291_ & new_n4595_;
  assign new_n4597_ = ~new_n4593_ & ~new_n4596_;
  assign new_n4598_ = new_n2294_ & new_n4595_;
  assign new_n4599_ = new_n2299_ & new_n4595_;
  assign new_n4600_ = ~new_n4598_ & ~new_n4599_;
  assign new_n4601_ = new_n4597_ & new_n4600_;
  assign new_n4602_ = new_n2309_ & new_n4595_;
  assign new_n4603_ = new_n2302_ & new_n4595_;
  assign new_n4604_ = new_n2306_ & new_n4595_;
  assign new_n4605_ = ~new_n4603_ & ~new_n4604_;
  assign new_n4606_ = ~new_n4602_ & new_n4605_;
  assign new_n4607_ = new_n4601_ & new_n4606_;
  assign new_n4608_ = new_n4592_ & new_n4607_;
  assign new_n4609_ = new_n4579_ & new_n4608_;
  assign new_n4610_ = new_n2315_ & new_n4595_;
  assign new_n4611_ = new_n2318_ & new_n4595_;
  assign new_n4612_ = ~new_n4610_ & ~new_n4611_;
  assign new_n4613_ = new_n2322_ & new_n4595_;
  assign new_n4614_ = new_n2324_ & new_n4595_;
  assign new_n4615_ = ~new_n4613_ & ~new_n4614_;
  assign new_n4616_ = new_n4612_ & new_n4615_;
  assign new_n4617_ = new_n2329_ & new_n4595_;
  assign new_n4618_ = new_n2331_ & new_n4595_;
  assign new_n4619_ = ~new_n4617_ & ~new_n4618_;
  assign new_n4620_ = A166 & new_n1237_;
  assign new_n4621_ = new_n1571_ & new_n4620_;
  assign new_n4622_ = new_n2403_ & new_n4621_;
  assign new_n4623_ = new_n2410_ & new_n4621_;
  assign new_n4624_ = ~new_n4622_ & ~new_n4623_;
  assign new_n4625_ = new_n4619_ & new_n4624_;
  assign new_n4626_ = new_n4616_ & new_n4625_;
  assign new_n4627_ = new_n2412_ & new_n4621_;
  assign new_n4628_ = new_n2415_ & new_n4621_;
  assign new_n4629_ = ~new_n4627_ & ~new_n4628_;
  assign new_n4630_ = new_n2419_ & new_n4621_;
  assign new_n4631_ = new_n2425_ & new_n4621_;
  assign new_n4632_ = ~new_n4630_ & ~new_n4631_;
  assign new_n4633_ = new_n4629_ & new_n4632_;
  assign new_n4634_ = new_n2437_ & new_n4621_;
  assign new_n4635_ = new_n2427_ & new_n4621_;
  assign new_n4636_ = new_n2423_ & new_n4621_;
  assign new_n4637_ = ~new_n4635_ & ~new_n4636_;
  assign new_n4638_ = ~new_n4634_ & new_n4637_;
  assign new_n4639_ = new_n4633_ & new_n4638_;
  assign new_n4640_ = new_n4626_ & new_n4639_;
  assign new_n4641_ = new_n2439_ & new_n4621_;
  assign new_n4642_ = new_n2442_ & new_n4621_;
  assign new_n4643_ = ~new_n4641_ & ~new_n4642_;
  assign new_n4644_ = new_n2444_ & new_n4621_;
  assign new_n4645_ = new_n2450_ & new_n4621_;
  assign new_n4646_ = ~new_n4644_ & ~new_n4645_;
  assign new_n4647_ = new_n4643_ & new_n4646_;
  assign new_n4648_ = new_n2457_ & new_n4621_;
  assign new_n4649_ = new_n2452_ & new_n4621_;
  assign new_n4650_ = new_n2455_ & new_n4621_;
  assign new_n4651_ = ~new_n4649_ & ~new_n4650_;
  assign new_n4652_ = ~new_n4648_ & new_n4651_;
  assign new_n4653_ = new_n4647_ & new_n4652_;
  assign new_n4654_ = ~A166 & new_n1036_;
  assign new_n4655_ = new_n1741_ & new_n4654_;
  assign new_n4656_ = new_n2291_ & new_n4655_;
  assign new_n4657_ = new_n2294_ & new_n4655_;
  assign new_n4658_ = ~new_n4656_ & ~new_n4657_;
  assign new_n4659_ = new_n2299_ & new_n4655_;
  assign new_n4660_ = new_n2302_ & new_n4655_;
  assign new_n4661_ = ~new_n4659_ & ~new_n4660_;
  assign new_n4662_ = new_n4658_ & new_n4661_;
  assign new_n4663_ = new_n2315_ & new_n4655_;
  assign new_n4664_ = new_n2306_ & new_n4655_;
  assign new_n4665_ = new_n2309_ & new_n4655_;
  assign new_n4666_ = ~new_n4664_ & ~new_n4665_;
  assign new_n4667_ = ~new_n4663_ & new_n4666_;
  assign new_n4668_ = new_n4662_ & new_n4667_;
  assign new_n4669_ = new_n4653_ & new_n4668_;
  assign new_n4670_ = new_n4640_ & new_n4669_;
  assign new_n4671_ = new_n4609_ & new_n4670_;
  assign new_n4672_ = new_n4548_ & new_n4671_;
  assign new_n4673_ = new_n2318_ & new_n4655_;
  assign new_n4674_ = new_n2322_ & new_n4655_;
  assign new_n4675_ = ~new_n4673_ & ~new_n4674_;
  assign new_n4676_ = new_n2324_ & new_n4655_;
  assign new_n4677_ = new_n2329_ & new_n4655_;
  assign new_n4678_ = ~new_n4676_ & ~new_n4677_;
  assign new_n4679_ = new_n4675_ & new_n4678_;
  assign new_n4680_ = new_n2331_ & new_n4655_;
  assign new_n4681_ = ~A166 & new_n1213_;
  assign new_n4682_ = new_n1741_ & new_n4681_;
  assign new_n4683_ = new_n2291_ & new_n4682_;
  assign new_n4684_ = ~new_n4680_ & ~new_n4683_;
  assign new_n4685_ = new_n2294_ & new_n4682_;
  assign new_n4686_ = new_n2299_ & new_n4682_;
  assign new_n4687_ = ~new_n4685_ & ~new_n4686_;
  assign new_n4688_ = new_n4684_ & new_n4687_;
  assign new_n4689_ = new_n4679_ & new_n4688_;
  assign new_n4690_ = new_n2302_ & new_n4682_;
  assign new_n4691_ = new_n2306_ & new_n4682_;
  assign new_n4692_ = ~new_n4690_ & ~new_n4691_;
  assign new_n4693_ = new_n2309_ & new_n4682_;
  assign new_n4694_ = new_n2315_ & new_n4682_;
  assign new_n4695_ = ~new_n4693_ & ~new_n4694_;
  assign new_n4696_ = new_n4692_ & new_n4695_;
  assign new_n4697_ = new_n2324_ & new_n4682_;
  assign new_n4698_ = new_n2318_ & new_n4682_;
  assign new_n4699_ = new_n2322_ & new_n4682_;
  assign new_n4700_ = ~new_n4698_ & ~new_n4699_;
  assign new_n4701_ = ~new_n4697_ & new_n4700_;
  assign new_n4702_ = new_n4696_ & new_n4701_;
  assign new_n4703_ = new_n4689_ & new_n4702_;
  assign new_n4704_ = new_n2329_ & new_n4682_;
  assign new_n4705_ = new_n2331_ & new_n4682_;
  assign new_n4706_ = ~new_n4704_ & ~new_n4705_;
  assign new_n4707_ = ~A166 & new_n1219_;
  assign new_n4708_ = new_n1741_ & new_n4707_;
  assign new_n4709_ = new_n2291_ & new_n4708_;
  assign new_n4710_ = new_n2294_ & new_n4708_;
  assign new_n4711_ = ~new_n4709_ & ~new_n4710_;
  assign new_n4712_ = new_n4706_ & new_n4711_;
  assign new_n4713_ = new_n2306_ & new_n4708_;
  assign new_n4714_ = new_n2299_ & new_n4708_;
  assign new_n4715_ = new_n2302_ & new_n4708_;
  assign new_n4716_ = ~new_n4714_ & ~new_n4715_;
  assign new_n4717_ = ~new_n4713_ & new_n4716_;
  assign new_n4718_ = new_n4712_ & new_n4717_;
  assign new_n4719_ = new_n2309_ & new_n4708_;
  assign new_n4720_ = new_n2315_ & new_n4708_;
  assign new_n4721_ = ~new_n4719_ & ~new_n4720_;
  assign new_n4722_ = new_n2318_ & new_n4708_;
  assign new_n4723_ = new_n2322_ & new_n4708_;
  assign new_n4724_ = ~new_n4722_ & ~new_n4723_;
  assign new_n4725_ = new_n4721_ & new_n4724_;
  assign new_n4726_ = new_n2331_ & new_n4708_;
  assign new_n4727_ = new_n2324_ & new_n4708_;
  assign new_n4728_ = new_n2329_ & new_n4708_;
  assign new_n4729_ = ~new_n4727_ & ~new_n4728_;
  assign new_n4730_ = ~new_n4726_ & new_n4729_;
  assign new_n4731_ = new_n4725_ & new_n4730_;
  assign new_n4732_ = new_n4718_ & new_n4731_;
  assign new_n4733_ = new_n4703_ & new_n4732_;
  assign new_n4734_ = ~A166 & new_n1225_;
  assign new_n4735_ = new_n1741_ & new_n4734_;
  assign new_n4736_ = new_n2291_ & new_n4735_;
  assign new_n4737_ = new_n2294_ & new_n4735_;
  assign new_n4738_ = ~new_n4736_ & ~new_n4737_;
  assign new_n4739_ = new_n2299_ & new_n4735_;
  assign new_n4740_ = new_n2302_ & new_n4735_;
  assign new_n4741_ = ~new_n4739_ & ~new_n4740_;
  assign new_n4742_ = new_n4738_ & new_n4741_;
  assign new_n4743_ = new_n2306_ & new_n4735_;
  assign new_n4744_ = new_n2309_ & new_n4735_;
  assign new_n4745_ = ~new_n4743_ & ~new_n4744_;
  assign new_n4746_ = new_n2315_ & new_n4735_;
  assign new_n4747_ = new_n2318_ & new_n4735_;
  assign new_n4748_ = ~new_n4746_ & ~new_n4747_;
  assign new_n4749_ = new_n4745_ & new_n4748_;
  assign new_n4750_ = new_n4742_ & new_n4749_;
  assign new_n4751_ = new_n2322_ & new_n4735_;
  assign new_n4752_ = new_n2324_ & new_n4735_;
  assign new_n4753_ = ~new_n4751_ & ~new_n4752_;
  assign new_n4754_ = new_n2329_ & new_n4735_;
  assign new_n4755_ = new_n2331_ & new_n4735_;
  assign new_n4756_ = ~new_n4754_ & ~new_n4755_;
  assign new_n4757_ = new_n4753_ & new_n4756_;
  assign new_n4758_ = ~A166 & new_n1237_;
  assign new_n4759_ = new_n1741_ & new_n4758_;
  assign new_n4760_ = new_n2412_ & new_n4759_;
  assign new_n4761_ = new_n2403_ & new_n4759_;
  assign new_n4762_ = new_n2410_ & new_n4759_;
  assign new_n4763_ = ~new_n4761_ & ~new_n4762_;
  assign new_n4764_ = ~new_n4760_ & new_n4763_;
  assign new_n4765_ = new_n4757_ & new_n4764_;
  assign new_n4766_ = new_n4750_ & new_n4765_;
  assign new_n4767_ = new_n2415_ & new_n4759_;
  assign new_n4768_ = new_n2419_ & new_n4759_;
  assign new_n4769_ = ~new_n4767_ & ~new_n4768_;
  assign new_n4770_ = new_n2425_ & new_n4759_;
  assign new_n4771_ = new_n2427_ & new_n4759_;
  assign new_n4772_ = ~new_n4770_ & ~new_n4771_;
  assign new_n4773_ = new_n4769_ & new_n4772_;
  assign new_n4774_ = new_n2439_ & new_n4759_;
  assign new_n4775_ = new_n2423_ & new_n4759_;
  assign new_n4776_ = new_n2437_ & new_n4759_;
  assign new_n4777_ = ~new_n4775_ & ~new_n4776_;
  assign new_n4778_ = ~new_n4774_ & new_n4777_;
  assign new_n4779_ = new_n4773_ & new_n4778_;
  assign new_n4780_ = new_n2442_ & new_n4759_;
  assign new_n4781_ = new_n2444_ & new_n4759_;
  assign new_n4782_ = ~new_n4780_ & ~new_n4781_;
  assign new_n4783_ = new_n2450_ & new_n4759_;
  assign new_n4784_ = new_n2452_ & new_n4759_;
  assign new_n4785_ = ~new_n4783_ & ~new_n4784_;
  assign new_n4786_ = new_n4782_ & new_n4785_;
  assign new_n4787_ = new_n36_ & new_n1905_;
  assign new_n4788_ = new_n2403_ & new_n4787_;
  assign new_n4789_ = new_n2455_ & new_n4759_;
  assign new_n4790_ = new_n2457_ & new_n4759_;
  assign new_n4791_ = ~new_n4789_ & ~new_n4790_;
  assign new_n4792_ = ~new_n4788_ & new_n4791_;
  assign new_n4793_ = new_n4786_ & new_n4792_;
  assign new_n4794_ = new_n4779_ & new_n4793_;
  assign new_n4795_ = new_n4766_ & new_n4794_;
  assign new_n4796_ = new_n4733_ & new_n4795_;
  assign new_n4797_ = new_n2410_ & new_n4787_;
  assign new_n4798_ = new_n2412_ & new_n4787_;
  assign new_n4799_ = ~new_n4797_ & ~new_n4798_;
  assign new_n4800_ = new_n2415_ & new_n4787_;
  assign new_n4801_ = new_n2419_ & new_n4787_;
  assign new_n4802_ = ~new_n4800_ & ~new_n4801_;
  assign new_n4803_ = new_n4799_ & new_n4802_;
  assign new_n4804_ = new_n2425_ & new_n4787_;
  assign new_n4805_ = new_n2427_ & new_n4787_;
  assign new_n4806_ = ~new_n4804_ & ~new_n4805_;
  assign new_n4807_ = new_n2423_ & new_n4787_;
  assign new_n4808_ = new_n2437_ & new_n4787_;
  assign new_n4809_ = ~new_n4807_ & ~new_n4808_;
  assign new_n4810_ = new_n4806_ & new_n4809_;
  assign new_n4811_ = new_n4803_ & new_n4810_;
  assign new_n4812_ = new_n2439_ & new_n4787_;
  assign new_n4813_ = new_n2442_ & new_n4787_;
  assign new_n4814_ = ~new_n4812_ & ~new_n4813_;
  assign new_n4815_ = new_n2444_ & new_n4787_;
  assign new_n4816_ = new_n2450_ & new_n4787_;
  assign new_n4817_ = ~new_n4815_ & ~new_n4816_;
  assign new_n4818_ = new_n4814_ & new_n4817_;
  assign new_n4819_ = new_n2457_ & new_n4787_;
  assign new_n4820_ = new_n2452_ & new_n4787_;
  assign new_n4821_ = new_n2455_ & new_n4787_;
  assign new_n4822_ = ~new_n4820_ & ~new_n4821_;
  assign new_n4823_ = ~new_n4819_ & new_n4822_;
  assign new_n4824_ = new_n4818_ & new_n4823_;
  assign new_n4825_ = new_n4811_ & new_n4824_;
  assign new_n4826_ = new_n1905_ & new_n4367_;
  assign new_n4827_ = new_n2291_ & new_n4826_;
  assign new_n4828_ = new_n2294_ & new_n4826_;
  assign new_n4829_ = ~new_n4827_ & ~new_n4828_;
  assign new_n4830_ = new_n2299_ & new_n4826_;
  assign new_n4831_ = new_n2302_ & new_n4826_;
  assign new_n4832_ = ~new_n4830_ & ~new_n4831_;
  assign new_n4833_ = new_n4829_ & new_n4832_;
  assign new_n4834_ = new_n2315_ & new_n4826_;
  assign new_n4835_ = new_n2306_ & new_n4826_;
  assign new_n4836_ = new_n2309_ & new_n4826_;
  assign new_n4837_ = ~new_n4835_ & ~new_n4836_;
  assign new_n4838_ = ~new_n4834_ & new_n4837_;
  assign new_n4839_ = new_n4833_ & new_n4838_;
  assign new_n4840_ = new_n2318_ & new_n4826_;
  assign new_n4841_ = new_n2322_ & new_n4826_;
  assign new_n4842_ = ~new_n4840_ & ~new_n4841_;
  assign new_n4843_ = new_n2324_ & new_n4826_;
  assign new_n4844_ = new_n2329_ & new_n4826_;
  assign new_n4845_ = ~new_n4843_ & ~new_n4844_;
  assign new_n4846_ = new_n4842_ & new_n4845_;
  assign new_n4847_ = new_n1905_ & new_n4390_;
  assign new_n4848_ = new_n2294_ & new_n4847_;
  assign new_n4849_ = new_n2331_ & new_n4826_;
  assign new_n4850_ = new_n2291_ & new_n4847_;
  assign new_n4851_ = ~new_n4849_ & ~new_n4850_;
  assign new_n4852_ = ~new_n4848_ & new_n4851_;
  assign new_n4853_ = new_n4846_ & new_n4852_;
  assign new_n4854_ = new_n4839_ & new_n4853_;
  assign new_n4855_ = new_n4825_ & new_n4854_;
  assign new_n4856_ = new_n2299_ & new_n4847_;
  assign new_n4857_ = new_n2302_ & new_n4847_;
  assign new_n4858_ = ~new_n4856_ & ~new_n4857_;
  assign new_n4859_ = new_n2306_ & new_n4847_;
  assign new_n4860_ = new_n2309_ & new_n4847_;
  assign new_n4861_ = ~new_n4859_ & ~new_n4860_;
  assign new_n4862_ = new_n4858_ & new_n4861_;
  assign new_n4863_ = new_n2315_ & new_n4847_;
  assign new_n4864_ = new_n2318_ & new_n4847_;
  assign new_n4865_ = ~new_n4863_ & ~new_n4864_;
  assign new_n4866_ = new_n2322_ & new_n4847_;
  assign new_n4867_ = new_n2324_ & new_n4847_;
  assign new_n4868_ = ~new_n4866_ & ~new_n4867_;
  assign new_n4869_ = new_n4865_ & new_n4868_;
  assign new_n4870_ = new_n4862_ & new_n4869_;
  assign new_n4871_ = new_n2329_ & new_n4847_;
  assign new_n4872_ = new_n2331_ & new_n4847_;
  assign new_n4873_ = ~new_n4871_ & ~new_n4872_;
  assign new_n4874_ = new_n50_ & new_n1918_;
  assign new_n4875_ = new_n2403_ & new_n4874_;
  assign new_n4876_ = new_n2410_ & new_n4874_;
  assign new_n4877_ = ~new_n4875_ & ~new_n4876_;
  assign new_n4878_ = new_n4873_ & new_n4877_;
  assign new_n4879_ = new_n2419_ & new_n4874_;
  assign new_n4880_ = new_n2412_ & new_n4874_;
  assign new_n4881_ = new_n2415_ & new_n4874_;
  assign new_n4882_ = ~new_n4880_ & ~new_n4881_;
  assign new_n4883_ = ~new_n4879_ & new_n4882_;
  assign new_n4884_ = new_n4878_ & new_n4883_;
  assign new_n4885_ = new_n4870_ & new_n4884_;
  assign new_n4886_ = new_n2425_ & new_n4874_;
  assign new_n4887_ = new_n2427_ & new_n4874_;
  assign new_n4888_ = ~new_n4886_ & ~new_n4887_;
  assign new_n4889_ = new_n2423_ & new_n4874_;
  assign new_n4890_ = new_n2437_ & new_n4874_;
  assign new_n4891_ = ~new_n4889_ & ~new_n4890_;
  assign new_n4892_ = new_n4888_ & new_n4891_;
  assign new_n4893_ = new_n2444_ & new_n4874_;
  assign new_n4894_ = new_n2439_ & new_n4874_;
  assign new_n4895_ = new_n2442_ & new_n4874_;
  assign new_n4896_ = ~new_n4894_ & ~new_n4895_;
  assign new_n4897_ = ~new_n4893_ & new_n4896_;
  assign new_n4898_ = new_n4892_ & new_n4897_;
  assign new_n4899_ = new_n2450_ & new_n4874_;
  assign new_n4900_ = new_n2452_ & new_n4874_;
  assign new_n4901_ = ~new_n4899_ & ~new_n4900_;
  assign new_n4902_ = new_n2455_ & new_n4874_;
  assign new_n4903_ = new_n2457_ & new_n4874_;
  assign new_n4904_ = ~new_n4902_ & ~new_n4903_;
  assign new_n4905_ = new_n4901_ & new_n4904_;
  assign new_n4906_ = new_n1918_ & new_n4456_;
  assign new_n4907_ = new_n2299_ & new_n4906_;
  assign new_n4908_ = new_n2291_ & new_n4906_;
  assign new_n4909_ = new_n2294_ & new_n4906_;
  assign new_n4910_ = ~new_n4908_ & ~new_n4909_;
  assign new_n4911_ = ~new_n4907_ & new_n4910_;
  assign new_n4912_ = new_n4905_ & new_n4911_;
  assign new_n4913_ = new_n4898_ & new_n4912_;
  assign new_n4914_ = new_n4885_ & new_n4913_;
  assign new_n4915_ = new_n4855_ & new_n4914_;
  assign new_n4916_ = new_n4796_ & new_n4915_;
  assign new_n4917_ = new_n4672_ & new_n4916_;
  assign new_n4918_ = new_n2302_ & new_n4906_;
  assign new_n4919_ = new_n2306_ & new_n4906_;
  assign new_n4920_ = ~new_n4918_ & ~new_n4919_;
  assign new_n4921_ = new_n2309_ & new_n4906_;
  assign new_n4922_ = new_n2315_ & new_n4906_;
  assign new_n4923_ = ~new_n4921_ & ~new_n4922_;
  assign new_n4924_ = new_n4920_ & new_n4923_;
  assign new_n4925_ = new_n2318_ & new_n4906_;
  assign new_n4926_ = new_n2322_ & new_n4906_;
  assign new_n4927_ = ~new_n4925_ & ~new_n4926_;
  assign new_n4928_ = new_n2324_ & new_n4906_;
  assign new_n4929_ = new_n2329_ & new_n4906_;
  assign new_n4930_ = ~new_n4928_ & ~new_n4929_;
  assign new_n4931_ = new_n4927_ & new_n4930_;
  assign new_n4932_ = new_n4924_ & new_n4931_;
  assign new_n4933_ = new_n2331_ & new_n4906_;
  assign new_n4934_ = new_n1918_ & new_n4482_;
  assign new_n4935_ = new_n2291_ & new_n4934_;
  assign new_n4936_ = ~new_n4933_ & ~new_n4935_;
  assign new_n4937_ = new_n2294_ & new_n4934_;
  assign new_n4938_ = new_n2299_ & new_n4934_;
  assign new_n4939_ = ~new_n4937_ & ~new_n4938_;
  assign new_n4940_ = new_n4936_ & new_n4939_;
  assign new_n4941_ = new_n2309_ & new_n4934_;
  assign new_n4942_ = new_n2302_ & new_n4934_;
  assign new_n4943_ = new_n2306_ & new_n4934_;
  assign new_n4944_ = ~new_n4942_ & ~new_n4943_;
  assign new_n4945_ = ~new_n4941_ & new_n4944_;
  assign new_n4946_ = new_n4940_ & new_n4945_;
  assign new_n4947_ = new_n4932_ & new_n4946_;
  assign new_n4948_ = new_n2315_ & new_n4934_;
  assign new_n4949_ = new_n2318_ & new_n4934_;
  assign new_n4950_ = ~new_n4948_ & ~new_n4949_;
  assign new_n4951_ = new_n2322_ & new_n4934_;
  assign new_n4952_ = new_n2324_ & new_n4934_;
  assign new_n4953_ = ~new_n4951_ & ~new_n4952_;
  assign new_n4954_ = new_n4950_ & new_n4953_;
  assign new_n4955_ = ~A170 & new_n4504_;
  assign new_n4956_ = new_n4503_ & new_n4955_;
  assign new_n4957_ = new_n2747_ & new_n4956_;
  assign new_n4958_ = new_n2329_ & new_n4934_;
  assign new_n4959_ = new_n2331_ & new_n4934_;
  assign new_n4960_ = ~new_n4958_ & ~new_n4959_;
  assign new_n4961_ = ~new_n4957_ & new_n4960_;
  assign new_n4962_ = new_n4954_ & new_n4961_;
  assign new_n4963_ = new_n4514_ & new_n4955_;
  assign new_n4964_ = new_n2755_ & new_n4963_;
  assign new_n4965_ = new_n1923_ & new_n4517_;
  assign new_n4966_ = new_n2291_ & new_n4965_;
  assign new_n4967_ = ~new_n4964_ & ~new_n4966_;
  assign new_n4968_ = new_n2294_ & new_n4965_;
  assign new_n4969_ = new_n2299_ & new_n4965_;
  assign new_n4970_ = ~new_n4968_ & ~new_n4969_;
  assign new_n4971_ = new_n4967_ & new_n4970_;
  assign new_n4972_ = new_n2309_ & new_n4965_;
  assign new_n4973_ = new_n2302_ & new_n4965_;
  assign new_n4974_ = new_n2306_ & new_n4965_;
  assign new_n4975_ = ~new_n4973_ & ~new_n4974_;
  assign new_n4976_ = ~new_n4972_ & new_n4975_;
  assign new_n4977_ = new_n4971_ & new_n4976_;
  assign new_n4978_ = new_n4962_ & new_n4977_;
  assign new_n4979_ = new_n4947_ & new_n4978_;
  assign new_n4980_ = new_n2315_ & new_n4965_;
  assign new_n4981_ = new_n2318_ & new_n4965_;
  assign new_n4982_ = ~new_n4980_ & ~new_n4981_;
  assign new_n4983_ = new_n2322_ & new_n4965_;
  assign new_n4984_ = new_n2324_ & new_n4965_;
  assign new_n4985_ = ~new_n4983_ & ~new_n4984_;
  assign new_n4986_ = new_n4982_ & new_n4985_;
  assign new_n4987_ = new_n2329_ & new_n4965_;
  assign new_n4988_ = new_n2331_ & new_n4965_;
  assign new_n4989_ = ~new_n4987_ & ~new_n4988_;
  assign new_n4990_ = new_n1923_ & new_n4538_;
  assign new_n4991_ = new_n2291_ & new_n4990_;
  assign new_n4992_ = new_n2294_ & new_n4990_;
  assign new_n4993_ = ~new_n4991_ & ~new_n4992_;
  assign new_n4994_ = new_n4989_ & new_n4993_;
  assign new_n4995_ = new_n4986_ & new_n4994_;
  assign new_n4996_ = new_n2299_ & new_n4990_;
  assign new_n4997_ = new_n2302_ & new_n4990_;
  assign new_n4998_ = ~new_n4996_ & ~new_n4997_;
  assign new_n4999_ = new_n2306_ & new_n4990_;
  assign new_n5000_ = new_n2309_ & new_n4990_;
  assign new_n5001_ = ~new_n4999_ & ~new_n5000_;
  assign new_n5002_ = new_n4998_ & new_n5001_;
  assign new_n5003_ = new_n2322_ & new_n4990_;
  assign new_n5004_ = new_n2315_ & new_n4990_;
  assign new_n5005_ = new_n2318_ & new_n4990_;
  assign new_n5006_ = ~new_n5004_ & ~new_n5005_;
  assign new_n5007_ = ~new_n5003_ & new_n5006_;
  assign new_n5008_ = new_n5002_ & new_n5007_;
  assign new_n5009_ = new_n4995_ & new_n5008_;
  assign new_n5010_ = new_n2324_ & new_n4990_;
  assign new_n5011_ = new_n2329_ & new_n4990_;
  assign new_n5012_ = ~new_n5010_ & ~new_n5011_;
  assign new_n5013_ = new_n2331_ & new_n4990_;
  assign new_n5014_ = new_n1923_ & new_n4568_;
  assign new_n5015_ = new_n2291_ & new_n5014_;
  assign new_n5016_ = ~new_n5013_ & ~new_n5015_;
  assign new_n5017_ = new_n5012_ & new_n5016_;
  assign new_n5018_ = new_n2302_ & new_n5014_;
  assign new_n5019_ = new_n2294_ & new_n5014_;
  assign new_n5020_ = new_n2299_ & new_n5014_;
  assign new_n5021_ = ~new_n5019_ & ~new_n5020_;
  assign new_n5022_ = ~new_n5018_ & new_n5021_;
  assign new_n5023_ = new_n5017_ & new_n5022_;
  assign new_n5024_ = new_n2306_ & new_n5014_;
  assign new_n5025_ = new_n2309_ & new_n5014_;
  assign new_n5026_ = ~new_n5024_ & ~new_n5025_;
  assign new_n5027_ = new_n2315_ & new_n5014_;
  assign new_n5028_ = new_n2318_ & new_n5014_;
  assign new_n5029_ = ~new_n5027_ & ~new_n5028_;
  assign new_n5030_ = new_n5026_ & new_n5029_;
  assign new_n5031_ = new_n2329_ & new_n5014_;
  assign new_n5032_ = new_n2322_ & new_n5014_;
  assign new_n5033_ = new_n2324_ & new_n5014_;
  assign new_n5034_ = ~new_n5032_ & ~new_n5033_;
  assign new_n5035_ = ~new_n5031_ & new_n5034_;
  assign new_n5036_ = new_n5030_ & new_n5035_;
  assign new_n5037_ = new_n5023_ & new_n5036_;
  assign new_n5038_ = new_n5009_ & new_n5037_;
  assign new_n5039_ = new_n4979_ & new_n5038_;
  assign new_n5040_ = new_n2331_ & new_n5014_;
  assign new_n5041_ = new_n1923_ & new_n4594_;
  assign new_n5042_ = new_n2291_ & new_n5041_;
  assign new_n5043_ = ~new_n5040_ & ~new_n5042_;
  assign new_n5044_ = new_n2294_ & new_n5041_;
  assign new_n5045_ = new_n2299_ & new_n5041_;
  assign new_n5046_ = ~new_n5044_ & ~new_n5045_;
  assign new_n5047_ = new_n5043_ & new_n5046_;
  assign new_n5048_ = new_n2302_ & new_n5041_;
  assign new_n5049_ = new_n2306_ & new_n5041_;
  assign new_n5050_ = ~new_n5048_ & ~new_n5049_;
  assign new_n5051_ = new_n2309_ & new_n5041_;
  assign new_n5052_ = new_n2315_ & new_n5041_;
  assign new_n5053_ = ~new_n5051_ & ~new_n5052_;
  assign new_n5054_ = new_n5050_ & new_n5053_;
  assign new_n5055_ = new_n5047_ & new_n5054_;
  assign new_n5056_ = new_n2318_ & new_n5041_;
  assign new_n5057_ = new_n2322_ & new_n5041_;
  assign new_n5058_ = ~new_n5056_ & ~new_n5057_;
  assign new_n5059_ = new_n2324_ & new_n5041_;
  assign new_n5060_ = new_n2329_ & new_n5041_;
  assign new_n5061_ = ~new_n5059_ & ~new_n5060_;
  assign new_n5062_ = new_n5058_ & new_n5061_;
  assign new_n5063_ = new_n1923_ & new_n4620_;
  assign new_n5064_ = new_n2410_ & new_n5063_;
  assign new_n5065_ = new_n2331_ & new_n5041_;
  assign new_n5066_ = new_n2403_ & new_n5063_;
  assign new_n5067_ = ~new_n5065_ & ~new_n5066_;
  assign new_n5068_ = ~new_n5064_ & new_n5067_;
  assign new_n5069_ = new_n5062_ & new_n5068_;
  assign new_n5070_ = new_n5055_ & new_n5069_;
  assign new_n5071_ = new_n2412_ & new_n5063_;
  assign new_n5072_ = new_n2415_ & new_n5063_;
  assign new_n5073_ = ~new_n5071_ & ~new_n5072_;
  assign new_n5074_ = new_n2419_ & new_n5063_;
  assign new_n5075_ = new_n2425_ & new_n5063_;
  assign new_n5076_ = ~new_n5074_ & ~new_n5075_;
  assign new_n5077_ = new_n5073_ & new_n5076_;
  assign new_n5078_ = new_n2437_ & new_n5063_;
  assign new_n5079_ = new_n2427_ & new_n5063_;
  assign new_n5080_ = new_n2423_ & new_n5063_;
  assign new_n5081_ = ~new_n5079_ & ~new_n5080_;
  assign new_n5082_ = ~new_n5078_ & new_n5081_;
  assign new_n5083_ = new_n5077_ & new_n5082_;
  assign new_n5084_ = new_n2439_ & new_n5063_;
  assign new_n5085_ = new_n2442_ & new_n5063_;
  assign new_n5086_ = ~new_n5084_ & ~new_n5085_;
  assign new_n5087_ = new_n2444_ & new_n5063_;
  assign new_n5088_ = new_n2450_ & new_n5063_;
  assign new_n5089_ = ~new_n5087_ & ~new_n5088_;
  assign new_n5090_ = new_n5086_ & new_n5089_;
  assign new_n5091_ = new_n2457_ & new_n5063_;
  assign new_n5092_ = new_n2452_ & new_n5063_;
  assign new_n5093_ = new_n2455_ & new_n5063_;
  assign new_n5094_ = ~new_n5092_ & ~new_n5093_;
  assign new_n5095_ = ~new_n5091_ & new_n5094_;
  assign new_n5096_ = new_n5090_ & new_n5095_;
  assign new_n5097_ = new_n5083_ & new_n5096_;
  assign new_n5098_ = new_n5070_ & new_n5097_;
  assign new_n5099_ = new_n2090_ & new_n4654_;
  assign new_n5100_ = new_n2291_ & new_n5099_;
  assign new_n5101_ = new_n2294_ & new_n5099_;
  assign new_n5102_ = ~new_n5100_ & ~new_n5101_;
  assign new_n5103_ = new_n2299_ & new_n5099_;
  assign new_n5104_ = new_n2302_ & new_n5099_;
  assign new_n5105_ = ~new_n5103_ & ~new_n5104_;
  assign new_n5106_ = new_n5102_ & new_n5105_;
  assign new_n5107_ = new_n2306_ & new_n5099_;
  assign new_n5108_ = new_n2309_ & new_n5099_;
  assign new_n5109_ = ~new_n5107_ & ~new_n5108_;
  assign new_n5110_ = new_n2315_ & new_n5099_;
  assign new_n5111_ = new_n2318_ & new_n5099_;
  assign new_n5112_ = ~new_n5110_ & ~new_n5111_;
  assign new_n5113_ = new_n5109_ & new_n5112_;
  assign new_n5114_ = new_n5106_ & new_n5113_;
  assign new_n5115_ = new_n2322_ & new_n5099_;
  assign new_n5116_ = new_n2324_ & new_n5099_;
  assign new_n5117_ = ~new_n5115_ & ~new_n5116_;
  assign new_n5118_ = new_n2329_ & new_n5099_;
  assign new_n5119_ = new_n2331_ & new_n5099_;
  assign new_n5120_ = ~new_n5118_ & ~new_n5119_;
  assign new_n5121_ = new_n5117_ & new_n5120_;
  assign new_n5122_ = new_n2090_ & new_n4681_;
  assign new_n5123_ = new_n2299_ & new_n5122_;
  assign new_n5124_ = new_n2291_ & new_n5122_;
  assign new_n5125_ = new_n2294_ & new_n5122_;
  assign new_n5126_ = ~new_n5124_ & ~new_n5125_;
  assign new_n5127_ = ~new_n5123_ & new_n5126_;
  assign new_n5128_ = new_n5121_ & new_n5127_;
  assign new_n5129_ = new_n5114_ & new_n5128_;
  assign new_n5130_ = new_n2302_ & new_n5122_;
  assign new_n5131_ = new_n2306_ & new_n5122_;
  assign new_n5132_ = ~new_n5130_ & ~new_n5131_;
  assign new_n5133_ = new_n2309_ & new_n5122_;
  assign new_n5134_ = new_n2315_ & new_n5122_;
  assign new_n5135_ = ~new_n5133_ & ~new_n5134_;
  assign new_n5136_ = new_n5132_ & new_n5135_;
  assign new_n5137_ = new_n2324_ & new_n5122_;
  assign new_n5138_ = new_n2318_ & new_n5122_;
  assign new_n5139_ = new_n2322_ & new_n5122_;
  assign new_n5140_ = ~new_n5138_ & ~new_n5139_;
  assign new_n5141_ = ~new_n5137_ & new_n5140_;
  assign new_n5142_ = new_n5136_ & new_n5141_;
  assign new_n5143_ = new_n2329_ & new_n5122_;
  assign new_n5144_ = new_n2331_ & new_n5122_;
  assign new_n5145_ = ~new_n5143_ & ~new_n5144_;
  assign new_n5146_ = new_n2090_ & new_n4707_;
  assign new_n5147_ = new_n2291_ & new_n5146_;
  assign new_n5148_ = new_n2294_ & new_n5146_;
  assign new_n5149_ = ~new_n5147_ & ~new_n5148_;
  assign new_n5150_ = new_n5145_ & new_n5149_;
  assign new_n5151_ = new_n2306_ & new_n5146_;
  assign new_n5152_ = new_n2299_ & new_n5146_;
  assign new_n5153_ = new_n2302_ & new_n5146_;
  assign new_n5154_ = ~new_n5152_ & ~new_n5153_;
  assign new_n5155_ = ~new_n5151_ & new_n5154_;
  assign new_n5156_ = new_n5150_ & new_n5155_;
  assign new_n5157_ = new_n5142_ & new_n5156_;
  assign new_n5158_ = new_n5129_ & new_n5157_;
  assign new_n5159_ = new_n5098_ & new_n5158_;
  assign new_n5160_ = new_n5039_ & new_n5159_;
  assign new_n5161_ = new_n2309_ & new_n5146_;
  assign new_n5162_ = new_n2315_ & new_n5146_;
  assign new_n5163_ = ~new_n5161_ & ~new_n5162_;
  assign new_n5164_ = new_n2318_ & new_n5146_;
  assign new_n5165_ = new_n2322_ & new_n5146_;
  assign new_n5166_ = ~new_n5164_ & ~new_n5165_;
  assign new_n5167_ = new_n5163_ & new_n5166_;
  assign new_n5168_ = new_n2324_ & new_n5146_;
  assign new_n5169_ = new_n2329_ & new_n5146_;
  assign new_n5170_ = ~new_n5168_ & ~new_n5169_;
  assign new_n5171_ = new_n2331_ & new_n5146_;
  assign new_n5172_ = new_n2090_ & new_n4734_;
  assign new_n5173_ = new_n2291_ & new_n5172_;
  assign new_n5174_ = ~new_n5171_ & ~new_n5173_;
  assign new_n5175_ = new_n5170_ & new_n5174_;
  assign new_n5176_ = new_n5167_ & new_n5175_;
  assign new_n5177_ = new_n2294_ & new_n5172_;
  assign new_n5178_ = new_n2299_ & new_n5172_;
  assign new_n5179_ = ~new_n5177_ & ~new_n5178_;
  assign new_n5180_ = new_n2302_ & new_n5172_;
  assign new_n5181_ = new_n2306_ & new_n5172_;
  assign new_n5182_ = ~new_n5180_ & ~new_n5181_;
  assign new_n5183_ = new_n5179_ & new_n5182_;
  assign new_n5184_ = new_n2318_ & new_n5172_;
  assign new_n5185_ = new_n2309_ & new_n5172_;
  assign new_n5186_ = new_n2315_ & new_n5172_;
  assign new_n5187_ = ~new_n5185_ & ~new_n5186_;
  assign new_n5188_ = ~new_n5184_ & new_n5187_;
  assign new_n5189_ = new_n5183_ & new_n5188_;
  assign new_n5190_ = new_n5176_ & new_n5189_;
  assign new_n5191_ = new_n2322_ & new_n5172_;
  assign new_n5192_ = new_n2324_ & new_n5172_;
  assign new_n5193_ = ~new_n5191_ & ~new_n5192_;
  assign new_n5194_ = new_n2329_ & new_n5172_;
  assign new_n5195_ = new_n2331_ & new_n5172_;
  assign new_n5196_ = ~new_n5194_ & ~new_n5195_;
  assign new_n5197_ = new_n5193_ & new_n5196_;
  assign new_n5198_ = new_n2090_ & new_n4758_;
  assign new_n5199_ = new_n2412_ & new_n5198_;
  assign new_n5200_ = new_n2403_ & new_n5198_;
  assign new_n5201_ = new_n2410_ & new_n5198_;
  assign new_n5202_ = ~new_n5200_ & ~new_n5201_;
  assign new_n5203_ = ~new_n5199_ & new_n5202_;
  assign new_n5204_ = new_n5197_ & new_n5203_;
  assign new_n5205_ = new_n2415_ & new_n5198_;
  assign new_n5206_ = new_n2419_ & new_n5198_;
  assign new_n5207_ = ~new_n5205_ & ~new_n5206_;
  assign new_n5208_ = new_n2425_ & new_n5198_;
  assign new_n5209_ = new_n2427_ & new_n5198_;
  assign new_n5210_ = ~new_n5208_ & ~new_n5209_;
  assign new_n5211_ = new_n5207_ & new_n5210_;
  assign new_n5212_ = new_n2439_ & new_n5198_;
  assign new_n5213_ = new_n2423_ & new_n5198_;
  assign new_n5214_ = new_n2437_ & new_n5198_;
  assign new_n5215_ = ~new_n5213_ & ~new_n5214_;
  assign new_n5216_ = ~new_n5212_ & new_n5215_;
  assign new_n5217_ = new_n5211_ & new_n5216_;
  assign new_n5218_ = new_n5204_ & new_n5217_;
  assign new_n5219_ = new_n5190_ & new_n5218_;
  assign new_n5220_ = new_n2442_ & new_n5198_;
  assign new_n5221_ = new_n2444_ & new_n5198_;
  assign new_n5222_ = ~new_n5220_ & ~new_n5221_;
  assign new_n5223_ = new_n2450_ & new_n5198_;
  assign new_n5224_ = new_n2452_ & new_n5198_;
  assign new_n5225_ = ~new_n5223_ & ~new_n5224_;
  assign new_n5226_ = new_n5222_ & new_n5225_;
  assign new_n5227_ = new_n2455_ & new_n5198_;
  assign new_n5228_ = new_n2457_ & new_n5198_;
  assign new_n5229_ = ~new_n5227_ & ~new_n5228_;
  assign new_n5230_ = new_n36_ & new_n2260_;
  assign new_n5231_ = new_n2403_ & new_n5230_;
  assign new_n5232_ = new_n2410_ & new_n5230_;
  assign new_n5233_ = ~new_n5231_ & ~new_n5232_;
  assign new_n5234_ = new_n5229_ & new_n5233_;
  assign new_n5235_ = new_n5226_ & new_n5234_;
  assign new_n5236_ = new_n2412_ & new_n5230_;
  assign new_n5237_ = new_n2415_ & new_n5230_;
  assign new_n5238_ = ~new_n5236_ & ~new_n5237_;
  assign new_n5239_ = new_n2419_ & new_n5230_;
  assign new_n5240_ = new_n2425_ & new_n5230_;
  assign new_n5241_ = ~new_n5239_ & ~new_n5240_;
  assign new_n5242_ = new_n5238_ & new_n5241_;
  assign new_n5243_ = new_n2437_ & new_n5230_;
  assign new_n5244_ = new_n2427_ & new_n5230_;
  assign new_n5245_ = new_n2423_ & new_n5230_;
  assign new_n5246_ = ~new_n5244_ & ~new_n5245_;
  assign new_n5247_ = ~new_n5243_ & new_n5246_;
  assign new_n5248_ = new_n5242_ & new_n5247_;
  assign new_n5249_ = new_n5235_ & new_n5248_;
  assign new_n5250_ = new_n2439_ & new_n5230_;
  assign new_n5251_ = new_n2442_ & new_n5230_;
  assign new_n5252_ = ~new_n5250_ & ~new_n5251_;
  assign new_n5253_ = new_n2444_ & new_n5230_;
  assign new_n5254_ = new_n2450_ & new_n5230_;
  assign new_n5255_ = ~new_n5253_ & ~new_n5254_;
  assign new_n5256_ = new_n5252_ & new_n5255_;
  assign new_n5257_ = new_n2457_ & new_n5230_;
  assign new_n5258_ = new_n2452_ & new_n5230_;
  assign new_n5259_ = new_n2455_ & new_n5230_;
  assign new_n5260_ = ~new_n5258_ & ~new_n5259_;
  assign new_n5261_ = ~new_n5257_ & new_n5260_;
  assign new_n5262_ = new_n5256_ & new_n5261_;
  assign new_n5263_ = new_n2260_ & new_n4367_;
  assign new_n5264_ = new_n2291_ & new_n5263_;
  assign new_n5265_ = new_n2294_ & new_n5263_;
  assign new_n5266_ = ~new_n5264_ & ~new_n5265_;
  assign new_n5267_ = new_n2299_ & new_n5263_;
  assign new_n5268_ = new_n2302_ & new_n5263_;
  assign new_n5269_ = ~new_n5267_ & ~new_n5268_;
  assign new_n5270_ = new_n5266_ & new_n5269_;
  assign new_n5271_ = new_n2315_ & new_n5263_;
  assign new_n5272_ = new_n2306_ & new_n5263_;
  assign new_n5273_ = new_n2309_ & new_n5263_;
  assign new_n5274_ = ~new_n5272_ & ~new_n5273_;
  assign new_n5275_ = ~new_n5271_ & new_n5274_;
  assign new_n5276_ = new_n5270_ & new_n5275_;
  assign new_n5277_ = new_n5262_ & new_n5276_;
  assign new_n5278_ = new_n5249_ & new_n5277_;
  assign new_n5279_ = new_n5219_ & new_n5278_;
  assign new_n5280_ = new_n2318_ & new_n5263_;
  assign new_n5281_ = new_n2322_ & new_n5263_;
  assign new_n5282_ = ~new_n5280_ & ~new_n5281_;
  assign new_n5283_ = new_n2324_ & new_n5263_;
  assign new_n5284_ = new_n2329_ & new_n5263_;
  assign new_n5285_ = ~new_n5283_ & ~new_n5284_;
  assign new_n5286_ = new_n5282_ & new_n5285_;
  assign new_n5287_ = new_n2331_ & new_n5263_;
  assign new_n5288_ = new_n2260_ & new_n4390_;
  assign new_n5289_ = new_n2291_ & new_n5288_;
  assign new_n5290_ = ~new_n5287_ & ~new_n5289_;
  assign new_n5291_ = new_n2294_ & new_n5288_;
  assign new_n5292_ = new_n2299_ & new_n5288_;
  assign new_n5293_ = ~new_n5291_ & ~new_n5292_;
  assign new_n5294_ = new_n5290_ & new_n5293_;
  assign new_n5295_ = new_n5286_ & new_n5294_;
  assign new_n5296_ = new_n2302_ & new_n5288_;
  assign new_n5297_ = new_n2306_ & new_n5288_;
  assign new_n5298_ = ~new_n5296_ & ~new_n5297_;
  assign new_n5299_ = new_n2309_ & new_n5288_;
  assign new_n5300_ = new_n2315_ & new_n5288_;
  assign new_n5301_ = ~new_n5299_ & ~new_n5300_;
  assign new_n5302_ = new_n5298_ & new_n5301_;
  assign new_n5303_ = new_n2324_ & new_n5288_;
  assign new_n5304_ = new_n2318_ & new_n5288_;
  assign new_n5305_ = new_n2322_ & new_n5288_;
  assign new_n5306_ = ~new_n5304_ & ~new_n5305_;
  assign new_n5307_ = ~new_n5303_ & new_n5306_;
  assign new_n5308_ = new_n5302_ & new_n5307_;
  assign new_n5309_ = new_n5295_ & new_n5308_;
  assign new_n5310_ = new_n2329_ & new_n5288_;
  assign new_n5311_ = new_n2331_ & new_n5288_;
  assign new_n5312_ = ~new_n5310_ & ~new_n5311_;
  assign new_n5313_ = new_n50_ & new_n2265_;
  assign new_n5314_ = new_n2403_ & new_n5313_;
  assign new_n5315_ = new_n2410_ & new_n5313_;
  assign new_n5316_ = ~new_n5314_ & ~new_n5315_;
  assign new_n5317_ = new_n5312_ & new_n5316_;
  assign new_n5318_ = new_n2419_ & new_n5313_;
  assign new_n5319_ = new_n2412_ & new_n5313_;
  assign new_n5320_ = new_n2415_ & new_n5313_;
  assign new_n5321_ = ~new_n5319_ & ~new_n5320_;
  assign new_n5322_ = ~new_n5318_ & new_n5321_;
  assign new_n5323_ = new_n5317_ & new_n5322_;
  assign new_n5324_ = new_n2425_ & new_n5313_;
  assign new_n5325_ = new_n2427_ & new_n5313_;
  assign new_n5326_ = ~new_n5324_ & ~new_n5325_;
  assign new_n5327_ = new_n2423_ & new_n5313_;
  assign new_n5328_ = new_n2437_ & new_n5313_;
  assign new_n5329_ = ~new_n5327_ & ~new_n5328_;
  assign new_n5330_ = new_n5326_ & new_n5329_;
  assign new_n5331_ = new_n2444_ & new_n5313_;
  assign new_n5332_ = new_n2439_ & new_n5313_;
  assign new_n5333_ = new_n2442_ & new_n5313_;
  assign new_n5334_ = ~new_n5332_ & ~new_n5333_;
  assign new_n5335_ = ~new_n5331_ & new_n5334_;
  assign new_n5336_ = new_n5330_ & new_n5335_;
  assign new_n5337_ = new_n5323_ & new_n5336_;
  assign new_n5338_ = new_n5309_ & new_n5337_;
  assign new_n5339_ = new_n2450_ & new_n5313_;
  assign new_n5340_ = new_n2452_ & new_n5313_;
  assign new_n5341_ = ~new_n5339_ & ~new_n5340_;
  assign new_n5342_ = new_n2455_ & new_n5313_;
  assign new_n5343_ = new_n2457_ & new_n5313_;
  assign new_n5344_ = ~new_n5342_ & ~new_n5343_;
  assign new_n5345_ = new_n5341_ & new_n5344_;
  assign new_n5346_ = new_n2265_ & new_n4456_;
  assign new_n5347_ = new_n2299_ & new_n5346_;
  assign new_n5348_ = new_n2291_ & new_n5346_;
  assign new_n5349_ = new_n2294_ & new_n5346_;
  assign new_n5350_ = ~new_n5348_ & ~new_n5349_;
  assign new_n5351_ = ~new_n5347_ & new_n5350_;
  assign new_n5352_ = new_n5345_ & new_n5351_;
  assign new_n5353_ = new_n2302_ & new_n5346_;
  assign new_n5354_ = new_n2306_ & new_n5346_;
  assign new_n5355_ = ~new_n5353_ & ~new_n5354_;
  assign new_n5356_ = new_n2309_ & new_n5346_;
  assign new_n5357_ = new_n2315_ & new_n5346_;
  assign new_n5358_ = ~new_n5356_ & ~new_n5357_;
  assign new_n5359_ = new_n5355_ & new_n5358_;
  assign new_n5360_ = new_n2324_ & new_n5346_;
  assign new_n5361_ = new_n2318_ & new_n5346_;
  assign new_n5362_ = new_n2322_ & new_n5346_;
  assign new_n5363_ = ~new_n5361_ & ~new_n5362_;
  assign new_n5364_ = ~new_n5360_ & new_n5363_;
  assign new_n5365_ = new_n5359_ & new_n5364_;
  assign new_n5366_ = new_n5352_ & new_n5365_;
  assign new_n5367_ = new_n2329_ & new_n5346_;
  assign new_n5368_ = new_n2331_ & new_n5346_;
  assign new_n5369_ = ~new_n5367_ & ~new_n5368_;
  assign new_n5370_ = new_n2265_ & new_n4482_;
  assign new_n5371_ = new_n2291_ & new_n5370_;
  assign new_n5372_ = new_n2294_ & new_n5370_;
  assign new_n5373_ = ~new_n5371_ & ~new_n5372_;
  assign new_n5374_ = new_n5369_ & new_n5373_;
  assign new_n5375_ = new_n2306_ & new_n5370_;
  assign new_n5376_ = new_n2299_ & new_n5370_;
  assign new_n5377_ = new_n2302_ & new_n5370_;
  assign new_n5378_ = ~new_n5376_ & ~new_n5377_;
  assign new_n5379_ = ~new_n5375_ & new_n5378_;
  assign new_n5380_ = new_n5374_ & new_n5379_;
  assign new_n5381_ = new_n2309_ & new_n5370_;
  assign new_n5382_ = new_n2315_ & new_n5370_;
  assign new_n5383_ = ~new_n5381_ & ~new_n5382_;
  assign new_n5384_ = new_n2318_ & new_n5370_;
  assign new_n5385_ = new_n2322_ & new_n5370_;
  assign new_n5386_ = ~new_n5384_ & ~new_n5385_;
  assign new_n5387_ = new_n5383_ & new_n5386_;
  assign new_n5388_ = new_n2331_ & new_n5370_;
  assign new_n5389_ = new_n2324_ & new_n5370_;
  assign new_n5390_ = new_n2329_ & new_n5370_;
  assign new_n5391_ = ~new_n5389_ & ~new_n5390_;
  assign new_n5392_ = ~new_n5388_ & new_n5391_;
  assign new_n5393_ = new_n5387_ & new_n5392_;
  assign new_n5394_ = new_n5380_ & new_n5393_;
  assign new_n5395_ = new_n5366_ & new_n5394_;
  assign new_n5396_ = new_n5338_ & new_n5395_;
  assign new_n5397_ = new_n5279_ & new_n5396_;
  assign new_n5398_ = new_n5160_ & new_n5397_;
  assign new_n5399_ = new_n4917_ & new_n5398_;
  assign new_n5400_ = ~A167 & new_n717_;
  assign new_n5401_ = new_n4503_ & new_n5400_;
  assign new_n5402_ = new_n2747_ & new_n5401_;
  assign new_n5403_ = new_n4514_ & new_n5400_;
  assign new_n5404_ = new_n2755_ & new_n5403_;
  assign new_n5405_ = ~new_n5402_ & ~new_n5404_;
  assign new_n5406_ = new_n36_ & new_n2270_;
  assign new_n5407_ = new_n2403_ & new_n5406_;
  assign new_n5408_ = new_n2410_ & new_n5406_;
  assign new_n5409_ = ~new_n5407_ & ~new_n5408_;
  assign new_n5410_ = new_n5405_ & new_n5409_;
  assign new_n5411_ = new_n2412_ & new_n5406_;
  assign new_n5412_ = new_n2415_ & new_n5406_;
  assign new_n5413_ = ~new_n5411_ & ~new_n5412_;
  assign new_n5414_ = new_n2419_ & new_n5406_;
  assign new_n5415_ = new_n2425_ & new_n5406_;
  assign new_n5416_ = ~new_n5414_ & ~new_n5415_;
  assign new_n5417_ = new_n5413_ & new_n5416_;
  assign new_n5418_ = new_n5410_ & new_n5417_;
  assign new_n5419_ = new_n2427_ & new_n5406_;
  assign new_n5420_ = new_n2423_ & new_n5406_;
  assign new_n5421_ = ~new_n5419_ & ~new_n5420_;
  assign new_n5422_ = new_n2437_ & new_n5406_;
  assign new_n5423_ = new_n2439_ & new_n5406_;
  assign new_n5424_ = ~new_n5422_ & ~new_n5423_;
  assign new_n5425_ = new_n5421_ & new_n5424_;
  assign new_n5426_ = new_n2450_ & new_n5406_;
  assign new_n5427_ = new_n2442_ & new_n5406_;
  assign new_n5428_ = new_n2444_ & new_n5406_;
  assign new_n5429_ = ~new_n5427_ & ~new_n5428_;
  assign new_n5430_ = ~new_n5426_ & new_n5429_;
  assign new_n5431_ = new_n5425_ & new_n5430_;
  assign new_n5432_ = new_n5418_ & new_n5431_;
  assign new_n5433_ = new_n2452_ & new_n5406_;
  assign new_n5434_ = new_n2455_ & new_n5406_;
  assign new_n5435_ = ~new_n5433_ & ~new_n5434_;
  assign new_n5436_ = new_n2457_ & new_n5406_;
  assign new_n5437_ = new_n2270_ & new_n4367_;
  assign new_n5438_ = new_n2291_ & new_n5437_;
  assign new_n5439_ = ~new_n5436_ & ~new_n5438_;
  assign new_n5440_ = new_n5435_ & new_n5439_;
  assign new_n5441_ = new_n2302_ & new_n5437_;
  assign new_n5442_ = new_n2294_ & new_n5437_;
  assign new_n5443_ = new_n2299_ & new_n5437_;
  assign new_n5444_ = ~new_n5442_ & ~new_n5443_;
  assign new_n5445_ = ~new_n5441_ & new_n5444_;
  assign new_n5446_ = new_n5440_ & new_n5445_;
  assign new_n5447_ = new_n2306_ & new_n5437_;
  assign new_n5448_ = new_n2309_ & new_n5437_;
  assign new_n5449_ = ~new_n5447_ & ~new_n5448_;
  assign new_n5450_ = new_n2315_ & new_n5437_;
  assign new_n5451_ = new_n2318_ & new_n5437_;
  assign new_n5452_ = ~new_n5450_ & ~new_n5451_;
  assign new_n5453_ = new_n5449_ & new_n5452_;
  assign new_n5454_ = new_n2329_ & new_n5437_;
  assign new_n5455_ = new_n2322_ & new_n5437_;
  assign new_n5456_ = new_n2324_ & new_n5437_;
  assign new_n5457_ = ~new_n5455_ & ~new_n5456_;
  assign new_n5458_ = ~new_n5454_ & new_n5457_;
  assign new_n5459_ = new_n5453_ & new_n5458_;
  assign new_n5460_ = new_n5446_ & new_n5459_;
  assign new_n5461_ = new_n5432_ & new_n5460_;
  assign new_n5462_ = new_n2331_ & new_n5437_;
  assign new_n5463_ = new_n2270_ & new_n4390_;
  assign new_n5464_ = new_n2291_ & new_n5463_;
  assign new_n5465_ = ~new_n5462_ & ~new_n5464_;
  assign new_n5466_ = new_n2294_ & new_n5463_;
  assign new_n5467_ = new_n2299_ & new_n5463_;
  assign new_n5468_ = ~new_n5466_ & ~new_n5467_;
  assign new_n5469_ = new_n5465_ & new_n5468_;
  assign new_n5470_ = new_n2302_ & new_n5463_;
  assign new_n5471_ = new_n2306_ & new_n5463_;
  assign new_n5472_ = ~new_n5470_ & ~new_n5471_;
  assign new_n5473_ = new_n2309_ & new_n5463_;
  assign new_n5474_ = new_n2315_ & new_n5463_;
  assign new_n5475_ = ~new_n5473_ & ~new_n5474_;
  assign new_n5476_ = new_n5472_ & new_n5475_;
  assign new_n5477_ = new_n5469_ & new_n5476_;
  assign new_n5478_ = new_n2318_ & new_n5463_;
  assign new_n5479_ = new_n2322_ & new_n5463_;
  assign new_n5480_ = ~new_n5478_ & ~new_n5479_;
  assign new_n5481_ = new_n2324_ & new_n5463_;
  assign new_n5482_ = new_n2329_ & new_n5463_;
  assign new_n5483_ = ~new_n5481_ & ~new_n5482_;
  assign new_n5484_ = new_n5480_ & new_n5483_;
  assign new_n5485_ = new_n50_ & new_n2285_;
  assign new_n5486_ = new_n2410_ & new_n5485_;
  assign new_n5487_ = new_n2331_ & new_n5463_;
  assign new_n5488_ = new_n2403_ & new_n5485_;
  assign new_n5489_ = ~new_n5487_ & ~new_n5488_;
  assign new_n5490_ = ~new_n5486_ & new_n5489_;
  assign new_n5491_ = new_n5484_ & new_n5490_;
  assign new_n5492_ = new_n5477_ & new_n5491_;
  assign new_n5493_ = new_n2412_ & new_n5485_;
  assign new_n5494_ = new_n2415_ & new_n5485_;
  assign new_n5495_ = ~new_n5493_ & ~new_n5494_;
  assign new_n5496_ = new_n2419_ & new_n5485_;
  assign new_n5497_ = new_n2425_ & new_n5485_;
  assign new_n5498_ = ~new_n5496_ & ~new_n5497_;
  assign new_n5499_ = new_n5495_ & new_n5498_;
  assign new_n5500_ = new_n2437_ & new_n5485_;
  assign new_n5501_ = new_n2427_ & new_n5485_;
  assign new_n5502_ = new_n2423_ & new_n5485_;
  assign new_n5503_ = ~new_n5501_ & ~new_n5502_;
  assign new_n5504_ = ~new_n5500_ & new_n5503_;
  assign new_n5505_ = new_n5499_ & new_n5504_;
  assign new_n5506_ = new_n2439_ & new_n5485_;
  assign new_n5507_ = new_n2442_ & new_n5485_;
  assign new_n5508_ = ~new_n5506_ & ~new_n5507_;
  assign new_n5509_ = new_n2444_ & new_n5485_;
  assign new_n5510_ = new_n2450_ & new_n5485_;
  assign new_n5511_ = ~new_n5509_ & ~new_n5510_;
  assign new_n5512_ = new_n5508_ & new_n5511_;
  assign new_n5513_ = new_n2457_ & new_n5485_;
  assign new_n5514_ = new_n2452_ & new_n5485_;
  assign new_n5515_ = new_n2455_ & new_n5485_;
  assign new_n5516_ = ~new_n5514_ & ~new_n5515_;
  assign new_n5517_ = ~new_n5513_ & new_n5516_;
  assign new_n5518_ = new_n5512_ & new_n5517_;
  assign new_n5519_ = new_n5505_ & new_n5518_;
  assign new_n5520_ = new_n5492_ & new_n5519_;
  assign new_n5521_ = new_n5461_ & new_n5520_;
  assign new_n5522_ = new_n2285_ & new_n4456_;
  assign new_n5523_ = new_n2291_ & new_n5522_;
  assign new_n5524_ = new_n2294_ & new_n5522_;
  assign new_n5525_ = ~new_n5523_ & ~new_n5524_;
  assign new_n5526_ = new_n2299_ & new_n5522_;
  assign new_n5527_ = new_n2302_ & new_n5522_;
  assign new_n5528_ = ~new_n5526_ & ~new_n5527_;
  assign new_n5529_ = new_n5525_ & new_n5528_;
  assign new_n5530_ = new_n2306_ & new_n5522_;
  assign new_n5531_ = new_n2309_ & new_n5522_;
  assign new_n5532_ = ~new_n5530_ & ~new_n5531_;
  assign new_n5533_ = new_n2315_ & new_n5522_;
  assign new_n5534_ = new_n2318_ & new_n5522_;
  assign new_n5535_ = ~new_n5533_ & ~new_n5534_;
  assign new_n5536_ = new_n5532_ & new_n5535_;
  assign new_n5537_ = new_n5529_ & new_n5536_;
  assign new_n5538_ = new_n2322_ & new_n5522_;
  assign new_n5539_ = new_n2324_ & new_n5522_;
  assign new_n5540_ = ~new_n5538_ & ~new_n5539_;
  assign new_n5541_ = new_n2329_ & new_n5522_;
  assign new_n5542_ = new_n2331_ & new_n5522_;
  assign new_n5543_ = ~new_n5541_ & ~new_n5542_;
  assign new_n5544_ = new_n5540_ & new_n5543_;
  assign new_n5545_ = new_n2285_ & new_n4482_;
  assign new_n5546_ = new_n2299_ & new_n5545_;
  assign new_n5547_ = new_n2291_ & new_n5545_;
  assign new_n5548_ = new_n2294_ & new_n5545_;
  assign new_n5549_ = ~new_n5547_ & ~new_n5548_;
  assign new_n5550_ = ~new_n5546_ & new_n5549_;
  assign new_n5551_ = new_n5544_ & new_n5550_;
  assign new_n5552_ = new_n5537_ & new_n5551_;
  assign new_n5553_ = new_n2302_ & new_n5545_;
  assign new_n5554_ = new_n2306_ & new_n5545_;
  assign new_n5555_ = ~new_n5553_ & ~new_n5554_;
  assign new_n5556_ = new_n2309_ & new_n5545_;
  assign new_n5557_ = new_n2315_ & new_n5545_;
  assign new_n5558_ = ~new_n5556_ & ~new_n5557_;
  assign new_n5559_ = new_n5555_ & new_n5558_;
  assign new_n5560_ = new_n2324_ & new_n5545_;
  assign new_n5561_ = new_n2318_ & new_n5545_;
  assign new_n5562_ = new_n2322_ & new_n5545_;
  assign new_n5563_ = ~new_n5561_ & ~new_n5562_;
  assign new_n5564_ = ~new_n5560_ & new_n5563_;
  assign new_n5565_ = new_n5559_ & new_n5564_;
  assign new_n5566_ = new_n2329_ & new_n5545_;
  assign new_n5567_ = new_n2331_ & new_n5545_;
  assign new_n5568_ = ~new_n5566_ & ~new_n5567_;
  assign new_n5569_ = A167 & new_n544_;
  assign new_n5570_ = new_n4503_ & new_n5569_;
  assign new_n5571_ = new_n2747_ & new_n5570_;
  assign new_n5572_ = new_n4514_ & new_n5569_;
  assign new_n5573_ = new_n2755_ & new_n5572_;
  assign new_n5574_ = ~new_n5571_ & ~new_n5573_;
  assign new_n5575_ = new_n5568_ & new_n5574_;
  assign new_n5576_ = new_n93_ & new_n2746_;
  assign new_n5577_ = new_n4125_ & new_n5576_;
  assign new_n5578_ = new_n75_ & new_n2746_;
  assign new_n5579_ = new_n4125_ & new_n5578_;
  assign new_n5580_ = new_n87_ & new_n2746_;
  assign new_n5581_ = new_n4125_ & new_n5580_;
  assign new_n5582_ = ~new_n5579_ & ~new_n5581_;
  assign new_n5583_ = ~new_n5577_ & new_n5582_;
  assign new_n5584_ = new_n5575_ & new_n5583_;
  assign new_n5585_ = new_n5565_ & new_n5584_;
  assign new_n5586_ = new_n5552_ & new_n5585_;
  assign new_n5587_ = new_n98_ & new_n2746_;
  assign new_n5588_ = new_n4125_ & new_n5587_;
  assign new_n5589_ = ~A266 & new_n108_;
  assign new_n5590_ = new_n28_ & new_n5589_;
  assign new_n5591_ = new_n4125_ & new_n5590_;
  assign new_n5592_ = ~new_n5588_ & ~new_n5591_;
  assign new_n5593_ = ~A266 & new_n112_;
  assign new_n5594_ = new_n28_ & new_n5593_;
  assign new_n5595_ = new_n4125_ & new_n5594_;
  assign new_n5596_ = new_n75_ & new_n2754_;
  assign new_n5597_ = new_n4130_ & new_n5596_;
  assign new_n5598_ = ~new_n5595_ & ~new_n5597_;
  assign new_n5599_ = new_n5592_ & new_n5598_;
  assign new_n5600_ = new_n87_ & new_n2754_;
  assign new_n5601_ = new_n4130_ & new_n5600_;
  assign new_n5602_ = new_n93_ & new_n2754_;
  assign new_n5603_ = new_n4130_ & new_n5602_;
  assign new_n5604_ = ~new_n5601_ & ~new_n5603_;
  assign new_n5605_ = new_n98_ & new_n2754_;
  assign new_n5606_ = new_n4130_ & new_n5605_;
  assign new_n5607_ = A266 & new_n108_;
  assign new_n5608_ = new_n28_ & new_n5607_;
  assign new_n5609_ = new_n4130_ & new_n5608_;
  assign new_n5610_ = ~new_n5606_ & ~new_n5609_;
  assign new_n5611_ = new_n5604_ & new_n5610_;
  assign new_n5612_ = new_n5599_ & new_n5611_;
  assign new_n5613_ = A266 & new_n112_;
  assign new_n5614_ = new_n28_ & new_n5613_;
  assign new_n5615_ = new_n4130_ & new_n5614_;
  assign new_n5616_ = new_n4269_ & new_n5578_;
  assign new_n5617_ = ~new_n5615_ & ~new_n5616_;
  assign new_n5618_ = new_n4269_ & new_n5580_;
  assign new_n5619_ = new_n4269_ & new_n5576_;
  assign new_n5620_ = ~new_n5618_ & ~new_n5619_;
  assign new_n5621_ = new_n5617_ & new_n5620_;
  assign new_n5622_ = new_n4269_ & new_n5594_;
  assign new_n5623_ = new_n4269_ & new_n5587_;
  assign new_n5624_ = new_n4269_ & new_n5590_;
  assign new_n5625_ = ~new_n5623_ & ~new_n5624_;
  assign new_n5626_ = ~new_n5622_ & new_n5625_;
  assign new_n5627_ = new_n5621_ & new_n5626_;
  assign new_n5628_ = new_n5612_ & new_n5627_;
  assign new_n5629_ = new_n4273_ & new_n5596_;
  assign new_n5630_ = new_n4273_ & new_n5600_;
  assign new_n5631_ = ~new_n5629_ & ~new_n5630_;
  assign new_n5632_ = new_n4273_ & new_n5602_;
  assign new_n5633_ = new_n4273_ & new_n5605_;
  assign new_n5634_ = ~new_n5632_ & ~new_n5633_;
  assign new_n5635_ = new_n5631_ & new_n5634_;
  assign new_n5636_ = new_n4278_ & new_n5578_;
  assign new_n5637_ = new_n4273_ & new_n5608_;
  assign new_n5638_ = new_n4273_ & new_n5614_;
  assign new_n5639_ = ~new_n5637_ & ~new_n5638_;
  assign new_n5640_ = ~new_n5636_ & new_n5639_;
  assign new_n5641_ = new_n5635_ & new_n5640_;
  assign new_n5642_ = new_n4278_ & new_n5580_;
  assign new_n5643_ = new_n4278_ & new_n5576_;
  assign new_n5644_ = ~new_n5642_ & ~new_n5643_;
  assign new_n5645_ = new_n4278_ & new_n5587_;
  assign new_n5646_ = new_n4278_ & new_n5590_;
  assign new_n5647_ = ~new_n5645_ & ~new_n5646_;
  assign new_n5648_ = new_n5644_ & new_n5647_;
  assign new_n5649_ = new_n4281_ & new_n5600_;
  assign new_n5650_ = new_n4278_ & new_n5594_;
  assign new_n5651_ = new_n4281_ & new_n5596_;
  assign new_n5652_ = ~new_n5650_ & ~new_n5651_;
  assign new_n5653_ = ~new_n5649_ & new_n5652_;
  assign new_n5654_ = new_n5648_ & new_n5653_;
  assign new_n5655_ = new_n5641_ & new_n5654_;
  assign new_n5656_ = new_n5628_ & new_n5655_;
  assign new_n5657_ = new_n5586_ & new_n5656_;
  assign new_n5658_ = new_n5521_ & new_n5657_;
  assign new_n5659_ = new_n4281_ & new_n5602_;
  assign new_n5660_ = new_n4281_ & new_n5605_;
  assign new_n5661_ = ~new_n5659_ & ~new_n5660_;
  assign new_n5662_ = new_n4281_ & new_n5608_;
  assign new_n5663_ = new_n4281_ & new_n5614_;
  assign new_n5664_ = ~new_n5662_ & ~new_n5663_;
  assign new_n5665_ = new_n5661_ & new_n5664_;
  assign new_n5666_ = new_n4285_ & new_n5578_;
  assign new_n5667_ = new_n4285_ & new_n5580_;
  assign new_n5668_ = ~new_n5666_ & ~new_n5667_;
  assign new_n5669_ = new_n4285_ & new_n5576_;
  assign new_n5670_ = new_n4285_ & new_n5587_;
  assign new_n5671_ = ~new_n5669_ & ~new_n5670_;
  assign new_n5672_ = new_n5668_ & new_n5671_;
  assign new_n5673_ = new_n5665_ & new_n5672_;
  assign new_n5674_ = new_n4285_ & new_n5590_;
  assign new_n5675_ = new_n4285_ & new_n5594_;
  assign new_n5676_ = ~new_n5674_ & ~new_n5675_;
  assign new_n5677_ = new_n4288_ & new_n5596_;
  assign new_n5678_ = new_n4288_ & new_n5600_;
  assign new_n5679_ = ~new_n5677_ & ~new_n5678_;
  assign new_n5680_ = new_n5676_ & new_n5679_;
  assign new_n5681_ = new_n4288_ & new_n5608_;
  assign new_n5682_ = new_n4288_ & new_n5602_;
  assign new_n5683_ = new_n4288_ & new_n5605_;
  assign new_n5684_ = ~new_n5682_ & ~new_n5683_;
  assign new_n5685_ = ~new_n5681_ & new_n5684_;
  assign new_n5686_ = new_n5680_ & new_n5685_;
  assign new_n5687_ = new_n5673_ & new_n5686_;
  assign new_n5688_ = new_n4288_ & new_n5614_;
  assign new_n5689_ = A269 & new_n74_;
  assign new_n5690_ = new_n4310_ & new_n5689_;
  assign new_n5691_ = new_n4296_ & new_n5690_;
  assign new_n5692_ = ~new_n5688_ & ~new_n5691_;
  assign new_n5693_ = A269 & new_n86_;
  assign new_n5694_ = new_n4310_ & new_n5693_;
  assign new_n5695_ = new_n4296_ & new_n5694_;
  assign new_n5696_ = A269 & new_n92_;
  assign new_n5697_ = new_n4310_ & new_n5696_;
  assign new_n5698_ = new_n4296_ & new_n5697_;
  assign new_n5699_ = ~new_n5695_ & ~new_n5698_;
  assign new_n5700_ = new_n5692_ & new_n5699_;
  assign new_n5701_ = A268 & new_n86_;
  assign new_n5702_ = new_n4310_ & new_n5701_;
  assign new_n5703_ = new_n4296_ & new_n5702_;
  assign new_n5704_ = A269 & new_n97_;
  assign new_n5705_ = new_n4310_ & new_n5704_;
  assign new_n5706_ = new_n4296_ & new_n5705_;
  assign new_n5707_ = A268 & new_n74_;
  assign new_n5708_ = new_n4310_ & new_n5707_;
  assign new_n5709_ = new_n4296_ & new_n5708_;
  assign new_n5710_ = ~new_n5706_ & ~new_n5709_;
  assign new_n5711_ = ~new_n5703_ & new_n5710_;
  assign new_n5712_ = new_n5700_ & new_n5711_;
  assign new_n5713_ = A268 & new_n92_;
  assign new_n5714_ = new_n4310_ & new_n5713_;
  assign new_n5715_ = new_n4296_ & new_n5714_;
  assign new_n5716_ = A268 & new_n97_;
  assign new_n5717_ = new_n4310_ & new_n5716_;
  assign new_n5718_ = new_n4296_ & new_n5717_;
  assign new_n5719_ = ~new_n5715_ & ~new_n5718_;
  assign new_n5720_ = new_n4326_ & new_n5689_;
  assign new_n5721_ = new_n4296_ & new_n5720_;
  assign new_n5722_ = new_n4326_ & new_n5693_;
  assign new_n5723_ = new_n4296_ & new_n5722_;
  assign new_n5724_ = ~new_n5721_ & ~new_n5723_;
  assign new_n5725_ = new_n5719_ & new_n5724_;
  assign new_n5726_ = new_n4326_ & new_n5707_;
  assign new_n5727_ = new_n4296_ & new_n5726_;
  assign new_n5728_ = new_n4326_ & new_n5696_;
  assign new_n5729_ = new_n4296_ & new_n5728_;
  assign new_n5730_ = new_n4326_ & new_n5704_;
  assign new_n5731_ = new_n4296_ & new_n5730_;
  assign new_n5732_ = ~new_n5729_ & ~new_n5731_;
  assign new_n5733_ = ~new_n5727_ & new_n5732_;
  assign new_n5734_ = new_n5725_ & new_n5733_;
  assign new_n5735_ = new_n5712_ & new_n5734_;
  assign new_n5736_ = new_n5687_ & new_n5735_;
  assign new_n5737_ = new_n4326_ & new_n5701_;
  assign new_n5738_ = new_n4296_ & new_n5737_;
  assign new_n5739_ = new_n4326_ & new_n5713_;
  assign new_n5740_ = new_n4296_ & new_n5739_;
  assign new_n5741_ = ~new_n5738_ & ~new_n5740_;
  assign new_n5742_ = new_n4326_ & new_n5716_;
  assign new_n5743_ = new_n4296_ & new_n5742_;
  assign new_n5744_ = ~A267 & new_n29_;
  assign new_n5745_ = new_n28_ & new_n5744_;
  assign new_n5746_ = ~A200 & new_n78_;
  assign new_n5747_ = new_n1563_ & new_n5746_;
  assign new_n5748_ = new_n5745_ & new_n5747_;
  assign new_n5749_ = ~new_n5743_ & ~new_n5748_;
  assign new_n5750_ = new_n5741_ & new_n5749_;
  assign new_n5751_ = ~A200 & new_n104_;
  assign new_n5752_ = new_n1563_ & new_n5751_;
  assign new_n5753_ = new_n5745_ & new_n5752_;
  assign new_n5754_ = A299 & new_n1282_;
  assign new_n5755_ = new_n2290_ & new_n5754_;
  assign new_n5756_ = new_n4368_ & new_n5755_;
  assign new_n5757_ = ~new_n5753_ & ~new_n5756_;
  assign new_n5758_ = A299 & new_n1290_;
  assign new_n5759_ = new_n2290_ & new_n5758_;
  assign new_n5760_ = new_n4368_ & new_n5759_;
  assign new_n5761_ = ~A299 & new_n1282_;
  assign new_n5762_ = new_n2293_ & new_n5761_;
  assign new_n5763_ = new_n4368_ & new_n5762_;
  assign new_n5764_ = ~new_n5760_ & ~new_n5763_;
  assign new_n5765_ = new_n5757_ & new_n5764_;
  assign new_n5766_ = new_n5750_ & new_n5765_;
  assign new_n5767_ = ~A299 & new_n1290_;
  assign new_n5768_ = new_n2293_ & new_n5767_;
  assign new_n5769_ = new_n4368_ & new_n5768_;
  assign new_n5770_ = new_n2298_ & new_n5754_;
  assign new_n5771_ = new_n4368_ & new_n5770_;
  assign new_n5772_ = ~new_n5769_ & ~new_n5771_;
  assign new_n5773_ = new_n2298_ & new_n5758_;
  assign new_n5774_ = new_n4368_ & new_n5773_;
  assign new_n5775_ = new_n2301_ & new_n5761_;
  assign new_n5776_ = new_n4368_ & new_n5775_;
  assign new_n5777_ = ~new_n5774_ & ~new_n5776_;
  assign new_n5778_ = new_n5772_ & new_n5777_;
  assign new_n5779_ = new_n2305_ & new_n5758_;
  assign new_n5780_ = new_n4368_ & new_n5779_;
  assign new_n5781_ = new_n2301_ & new_n5767_;
  assign new_n5782_ = new_n4368_ & new_n5781_;
  assign new_n5783_ = new_n2305_ & new_n5754_;
  assign new_n5784_ = new_n4368_ & new_n5783_;
  assign new_n5785_ = ~new_n5782_ & ~new_n5784_;
  assign new_n5786_ = ~new_n5780_ & new_n5785_;
  assign new_n5787_ = new_n5778_ & new_n5786_;
  assign new_n5788_ = new_n5766_ & new_n5787_;
  assign new_n5789_ = new_n2308_ & new_n5761_;
  assign new_n5790_ = new_n4368_ & new_n5789_;
  assign new_n5791_ = new_n2308_ & new_n5767_;
  assign new_n5792_ = new_n4368_ & new_n5791_;
  assign new_n5793_ = ~new_n5790_ & ~new_n5792_;
  assign new_n5794_ = new_n2314_ & new_n5754_;
  assign new_n5795_ = new_n4368_ & new_n5794_;
  assign new_n5796_ = new_n2314_ & new_n5758_;
  assign new_n5797_ = new_n4368_ & new_n5796_;
  assign new_n5798_ = ~new_n5795_ & ~new_n5797_;
  assign new_n5799_ = new_n5793_ & new_n5798_;
  assign new_n5800_ = new_n4391_ & new_n5755_;
  assign new_n5801_ = new_n2317_ & new_n5761_;
  assign new_n5802_ = new_n4368_ & new_n5801_;
  assign new_n5803_ = new_n2317_ & new_n5767_;
  assign new_n5804_ = new_n4368_ & new_n5803_;
  assign new_n5805_ = ~new_n5802_ & ~new_n5804_;
  assign new_n5806_ = ~new_n5800_ & new_n5805_;
  assign new_n5807_ = new_n5799_ & new_n5806_;
  assign new_n5808_ = new_n4391_ & new_n5759_;
  assign new_n5809_ = new_n4391_ & new_n5762_;
  assign new_n5810_ = ~new_n5808_ & ~new_n5809_;
  assign new_n5811_ = new_n4391_ & new_n5768_;
  assign new_n5812_ = new_n4391_ & new_n5770_;
  assign new_n5813_ = ~new_n5811_ & ~new_n5812_;
  assign new_n5814_ = new_n5810_ & new_n5813_;
  assign new_n5815_ = new_n4391_ & new_n5781_;
  assign new_n5816_ = new_n4391_ & new_n5773_;
  assign new_n5817_ = new_n4391_ & new_n5775_;
  assign new_n5818_ = ~new_n5816_ & ~new_n5817_;
  assign new_n5819_ = ~new_n5815_ & new_n5818_;
  assign new_n5820_ = new_n5814_ & new_n5819_;
  assign new_n5821_ = new_n5807_ & new_n5820_;
  assign new_n5822_ = new_n5788_ & new_n5821_;
  assign new_n5823_ = new_n5736_ & new_n5822_;
  assign new_n5824_ = new_n4391_ & new_n5783_;
  assign new_n5825_ = new_n4391_ & new_n5779_;
  assign new_n5826_ = ~new_n5824_ & ~new_n5825_;
  assign new_n5827_ = new_n4391_ & new_n5789_;
  assign new_n5828_ = new_n4391_ & new_n5791_;
  assign new_n5829_ = ~new_n5827_ & ~new_n5828_;
  assign new_n5830_ = new_n5826_ & new_n5829_;
  assign new_n5831_ = new_n4391_ & new_n5794_;
  assign new_n5832_ = new_n4391_ & new_n5796_;
  assign new_n5833_ = ~new_n5831_ & ~new_n5832_;
  assign new_n5834_ = new_n4391_ & new_n5801_;
  assign new_n5835_ = new_n4391_ & new_n5803_;
  assign new_n5836_ = ~new_n5834_ & ~new_n5835_;
  assign new_n5837_ = new_n5833_ & new_n5836_;
  assign new_n5838_ = new_n5830_ & new_n5837_;
  assign new_n5839_ = new_n4457_ & new_n5755_;
  assign new_n5840_ = new_n4457_ & new_n5759_;
  assign new_n5841_ = ~new_n5839_ & ~new_n5840_;
  assign new_n5842_ = new_n4457_ & new_n5762_;
  assign new_n5843_ = new_n4457_ & new_n5768_;
  assign new_n5844_ = ~new_n5842_ & ~new_n5843_;
  assign new_n5845_ = new_n5841_ & new_n5844_;
  assign new_n5846_ = new_n4457_ & new_n5775_;
  assign new_n5847_ = new_n4457_ & new_n5770_;
  assign new_n5848_ = new_n4457_ & new_n5773_;
  assign new_n5849_ = ~new_n5847_ & ~new_n5848_;
  assign new_n5850_ = ~new_n5846_ & new_n5849_;
  assign new_n5851_ = new_n5845_ & new_n5850_;
  assign new_n5852_ = new_n5838_ & new_n5851_;
  assign new_n5853_ = new_n4457_ & new_n5781_;
  assign new_n5854_ = new_n4457_ & new_n5783_;
  assign new_n5855_ = ~new_n5853_ & ~new_n5854_;
  assign new_n5856_ = new_n4457_ & new_n5779_;
  assign new_n5857_ = new_n4457_ & new_n5789_;
  assign new_n5858_ = ~new_n5856_ & ~new_n5857_;
  assign new_n5859_ = new_n5855_ & new_n5858_;
  assign new_n5860_ = new_n4457_ & new_n5796_;
  assign new_n5861_ = new_n4457_ & new_n5791_;
  assign new_n5862_ = new_n4457_ & new_n5794_;
  assign new_n5863_ = ~new_n5861_ & ~new_n5862_;
  assign new_n5864_ = ~new_n5860_ & new_n5863_;
  assign new_n5865_ = new_n5859_ & new_n5864_;
  assign new_n5866_ = new_n4457_ & new_n5801_;
  assign new_n5867_ = new_n4457_ & new_n5803_;
  assign new_n5868_ = ~new_n5866_ & ~new_n5867_;
  assign new_n5869_ = new_n4483_ & new_n5755_;
  assign new_n5870_ = new_n4483_ & new_n5759_;
  assign new_n5871_ = ~new_n5869_ & ~new_n5870_;
  assign new_n5872_ = new_n5868_ & new_n5871_;
  assign new_n5873_ = new_n4483_ & new_n5770_;
  assign new_n5874_ = new_n4483_ & new_n5762_;
  assign new_n5875_ = new_n4483_ & new_n5768_;
  assign new_n5876_ = ~new_n5874_ & ~new_n5875_;
  assign new_n5877_ = ~new_n5873_ & new_n5876_;
  assign new_n5878_ = new_n5872_ & new_n5877_;
  assign new_n5879_ = new_n5865_ & new_n5878_;
  assign new_n5880_ = new_n5852_ & new_n5879_;
  assign new_n5881_ = new_n4483_ & new_n5773_;
  assign new_n5882_ = new_n4483_ & new_n5775_;
  assign new_n5883_ = ~new_n5881_ & ~new_n5882_;
  assign new_n5884_ = new_n4483_ & new_n5781_;
  assign new_n5885_ = new_n4483_ & new_n5783_;
  assign new_n5886_ = ~new_n5884_ & ~new_n5885_;
  assign new_n5887_ = new_n5883_ & new_n5886_;
  assign new_n5888_ = new_n4483_ & new_n5779_;
  assign new_n5889_ = new_n4483_ & new_n5789_;
  assign new_n5890_ = ~new_n5888_ & ~new_n5889_;
  assign new_n5891_ = new_n4483_ & new_n5791_;
  assign new_n5892_ = new_n4483_ & new_n5794_;
  assign new_n5893_ = ~new_n5891_ & ~new_n5892_;
  assign new_n5894_ = new_n5890_ & new_n5893_;
  assign new_n5895_ = new_n5887_ & new_n5894_;
  assign new_n5896_ = new_n4483_ & new_n5796_;
  assign new_n5897_ = new_n4483_ & new_n5801_;
  assign new_n5898_ = ~new_n5896_ & ~new_n5897_;
  assign new_n5899_ = new_n4483_ & new_n5803_;
  assign new_n5900_ = A200 & new_n78_;
  assign new_n5901_ = new_n1557_ & new_n5900_;
  assign new_n5902_ = new_n5745_ & new_n5901_;
  assign new_n5903_ = ~new_n5899_ & ~new_n5902_;
  assign new_n5904_ = new_n5898_ & new_n5903_;
  assign new_n5905_ = ~A201 & ~A168;
  assign new_n5906_ = A169 & new_n5905_;
  assign new_n5907_ = new_n2871_ & new_n5906_;
  assign new_n5908_ = new_n5745_ & new_n5907_;
  assign new_n5909_ = A200 & new_n104_;
  assign new_n5910_ = new_n1557_ & new_n5909_;
  assign new_n5911_ = new_n5745_ & new_n5910_;
  assign new_n5912_ = new_n2839_ & new_n5906_;
  assign new_n5913_ = new_n5745_ & new_n5912_;
  assign new_n5914_ = ~new_n5911_ & ~new_n5913_;
  assign new_n5915_ = ~new_n5908_ & new_n5914_;
  assign new_n5916_ = new_n5904_ & new_n5915_;
  assign new_n5917_ = new_n5895_ & new_n5916_;
  assign new_n5918_ = new_n2896_ & new_n5906_;
  assign new_n5919_ = new_n5745_ & new_n5918_;
  assign new_n5920_ = new_n2920_ & new_n5906_;
  assign new_n5921_ = new_n5745_ & new_n5920_;
  assign new_n5922_ = ~new_n5919_ & ~new_n5921_;
  assign new_n5923_ = new_n4506_ & new_n5578_;
  assign new_n5924_ = new_n4506_ & new_n5580_;
  assign new_n5925_ = ~new_n5923_ & ~new_n5924_;
  assign new_n5926_ = new_n5922_ & new_n5925_;
  assign new_n5927_ = new_n4506_ & new_n5590_;
  assign new_n5928_ = new_n4506_ & new_n5576_;
  assign new_n5929_ = new_n4506_ & new_n5587_;
  assign new_n5930_ = ~new_n5928_ & ~new_n5929_;
  assign new_n5931_ = ~new_n5927_ & new_n5930_;
  assign new_n5932_ = new_n5926_ & new_n5931_;
  assign new_n5933_ = new_n4506_ & new_n5594_;
  assign new_n5934_ = new_n4515_ & new_n5596_;
  assign new_n5935_ = ~new_n5933_ & ~new_n5934_;
  assign new_n5936_ = new_n4515_ & new_n5600_;
  assign new_n5937_ = new_n4515_ & new_n5602_;
  assign new_n5938_ = ~new_n5936_ & ~new_n5937_;
  assign new_n5939_ = new_n5935_ & new_n5938_;
  assign new_n5940_ = new_n4515_ & new_n5614_;
  assign new_n5941_ = new_n4515_ & new_n5605_;
  assign new_n5942_ = new_n4515_ & new_n5608_;
  assign new_n5943_ = ~new_n5941_ & ~new_n5942_;
  assign new_n5944_ = ~new_n5940_ & new_n5943_;
  assign new_n5945_ = new_n5939_ & new_n5944_;
  assign new_n5946_ = new_n5932_ & new_n5945_;
  assign new_n5947_ = new_n5917_ & new_n5946_;
  assign new_n5948_ = new_n5880_ & new_n5947_;
  assign new_n5949_ = new_n5823_ & new_n5948_;
  assign new_n5950_ = new_n5658_ & new_n5949_;
  assign new_n5951_ = new_n4518_ & new_n5755_;
  assign new_n5952_ = new_n4518_ & new_n5759_;
  assign new_n5953_ = ~new_n5951_ & ~new_n5952_;
  assign new_n5954_ = new_n4518_ & new_n5762_;
  assign new_n5955_ = new_n4518_ & new_n5768_;
  assign new_n5956_ = ~new_n5954_ & ~new_n5955_;
  assign new_n5957_ = new_n5953_ & new_n5956_;
  assign new_n5958_ = new_n4518_ & new_n5770_;
  assign new_n5959_ = new_n4518_ & new_n5773_;
  assign new_n5960_ = ~new_n5958_ & ~new_n5959_;
  assign new_n5961_ = new_n4518_ & new_n5775_;
  assign new_n5962_ = new_n4518_ & new_n5781_;
  assign new_n5963_ = ~new_n5961_ & ~new_n5962_;
  assign new_n5964_ = new_n5960_ & new_n5963_;
  assign new_n5965_ = new_n5957_ & new_n5964_;
  assign new_n5966_ = new_n4518_ & new_n5783_;
  assign new_n5967_ = new_n4518_ & new_n5779_;
  assign new_n5968_ = ~new_n5966_ & ~new_n5967_;
  assign new_n5969_ = new_n4518_ & new_n5789_;
  assign new_n5970_ = new_n4518_ & new_n5791_;
  assign new_n5971_ = ~new_n5969_ & ~new_n5970_;
  assign new_n5972_ = new_n5968_ & new_n5971_;
  assign new_n5973_ = new_n4518_ & new_n5801_;
  assign new_n5974_ = new_n4518_ & new_n5794_;
  assign new_n5975_ = new_n4518_ & new_n5796_;
  assign new_n5976_ = ~new_n5974_ & ~new_n5975_;
  assign new_n5977_ = ~new_n5973_ & new_n5976_;
  assign new_n5978_ = new_n5972_ & new_n5977_;
  assign new_n5979_ = new_n5965_ & new_n5978_;
  assign new_n5980_ = new_n4518_ & new_n5803_;
  assign new_n5981_ = new_n4539_ & new_n5755_;
  assign new_n5982_ = ~new_n5980_ & ~new_n5981_;
  assign new_n5983_ = new_n4539_ & new_n5759_;
  assign new_n5984_ = new_n4539_ & new_n5762_;
  assign new_n5985_ = ~new_n5983_ & ~new_n5984_;
  assign new_n5986_ = new_n5982_ & new_n5985_;
  assign new_n5987_ = new_n4539_ & new_n5773_;
  assign new_n5988_ = new_n4539_ & new_n5768_;
  assign new_n5989_ = new_n4539_ & new_n5770_;
  assign new_n5990_ = ~new_n5988_ & ~new_n5989_;
  assign new_n5991_ = ~new_n5987_ & new_n5990_;
  assign new_n5992_ = new_n5986_ & new_n5991_;
  assign new_n5993_ = new_n4539_ & new_n5775_;
  assign new_n5994_ = new_n4539_ & new_n5781_;
  assign new_n5995_ = ~new_n5993_ & ~new_n5994_;
  assign new_n5996_ = new_n4539_ & new_n5783_;
  assign new_n5997_ = new_n4539_ & new_n5779_;
  assign new_n5998_ = ~new_n5996_ & ~new_n5997_;
  assign new_n5999_ = new_n5995_ & new_n5998_;
  assign new_n6000_ = new_n4539_ & new_n5794_;
  assign new_n6001_ = new_n4539_ & new_n5789_;
  assign new_n6002_ = new_n4539_ & new_n5791_;
  assign new_n6003_ = ~new_n6001_ & ~new_n6002_;
  assign new_n6004_ = ~new_n6000_ & new_n6003_;
  assign new_n6005_ = new_n5999_ & new_n6004_;
  assign new_n6006_ = new_n5992_ & new_n6005_;
  assign new_n6007_ = new_n5979_ & new_n6006_;
  assign new_n6008_ = new_n4539_ & new_n5796_;
  assign new_n6009_ = new_n4539_ & new_n5801_;
  assign new_n6010_ = ~new_n6008_ & ~new_n6009_;
  assign new_n6011_ = new_n4539_ & new_n5803_;
  assign new_n6012_ = new_n4569_ & new_n5755_;
  assign new_n6013_ = ~new_n6011_ & ~new_n6012_;
  assign new_n6014_ = new_n6010_ & new_n6013_;
  assign new_n6015_ = new_n4569_ & new_n5759_;
  assign new_n6016_ = new_n4569_ & new_n5762_;
  assign new_n6017_ = ~new_n6015_ & ~new_n6016_;
  assign new_n6018_ = new_n4569_ & new_n5768_;
  assign new_n6019_ = new_n4569_ & new_n5770_;
  assign new_n6020_ = ~new_n6018_ & ~new_n6019_;
  assign new_n6021_ = new_n6017_ & new_n6020_;
  assign new_n6022_ = new_n6014_ & new_n6021_;
  assign new_n6023_ = new_n4569_ & new_n5773_;
  assign new_n6024_ = new_n4569_ & new_n5775_;
  assign new_n6025_ = ~new_n6023_ & ~new_n6024_;
  assign new_n6026_ = new_n4569_ & new_n5781_;
  assign new_n6027_ = new_n4569_ & new_n5783_;
  assign new_n6028_ = ~new_n6026_ & ~new_n6027_;
  assign new_n6029_ = new_n6025_ & new_n6028_;
  assign new_n6030_ = new_n4569_ & new_n5791_;
  assign new_n6031_ = new_n4569_ & new_n5779_;
  assign new_n6032_ = new_n4569_ & new_n5789_;
  assign new_n6033_ = ~new_n6031_ & ~new_n6032_;
  assign new_n6034_ = ~new_n6030_ & new_n6033_;
  assign new_n6035_ = new_n6029_ & new_n6034_;
  assign new_n6036_ = new_n6022_ & new_n6035_;
  assign new_n6037_ = new_n4569_ & new_n5794_;
  assign new_n6038_ = new_n4569_ & new_n5796_;
  assign new_n6039_ = ~new_n6037_ & ~new_n6038_;
  assign new_n6040_ = new_n4569_ & new_n5801_;
  assign new_n6041_ = new_n4569_ & new_n5803_;
  assign new_n6042_ = ~new_n6040_ & ~new_n6041_;
  assign new_n6043_ = new_n6039_ & new_n6042_;
  assign new_n6044_ = new_n4595_ & new_n5762_;
  assign new_n6045_ = new_n4595_ & new_n5755_;
  assign new_n6046_ = new_n4595_ & new_n5759_;
  assign new_n6047_ = ~new_n6045_ & ~new_n6046_;
  assign new_n6048_ = ~new_n6044_ & new_n6047_;
  assign new_n6049_ = new_n6043_ & new_n6048_;
  assign new_n6050_ = new_n4595_ & new_n5768_;
  assign new_n6051_ = new_n4595_ & new_n5770_;
  assign new_n6052_ = ~new_n6050_ & ~new_n6051_;
  assign new_n6053_ = new_n4595_ & new_n5773_;
  assign new_n6054_ = new_n4595_ & new_n5775_;
  assign new_n6055_ = ~new_n6053_ & ~new_n6054_;
  assign new_n6056_ = new_n6052_ & new_n6055_;
  assign new_n6057_ = new_n4595_ & new_n5779_;
  assign new_n6058_ = new_n4595_ & new_n5781_;
  assign new_n6059_ = new_n4595_ & new_n5783_;
  assign new_n6060_ = ~new_n6058_ & ~new_n6059_;
  assign new_n6061_ = ~new_n6057_ & new_n6060_;
  assign new_n6062_ = new_n6056_ & new_n6061_;
  assign new_n6063_ = new_n6049_ & new_n6062_;
  assign new_n6064_ = new_n6036_ & new_n6063_;
  assign new_n6065_ = new_n6007_ & new_n6064_;
  assign new_n6066_ = new_n4595_ & new_n5789_;
  assign new_n6067_ = new_n4595_ & new_n5791_;
  assign new_n6068_ = ~new_n6066_ & ~new_n6067_;
  assign new_n6069_ = new_n4595_ & new_n5794_;
  assign new_n6070_ = new_n4595_ & new_n5796_;
  assign new_n6071_ = ~new_n6069_ & ~new_n6070_;
  assign new_n6072_ = new_n6068_ & new_n6071_;
  assign new_n6073_ = new_n4595_ & new_n5801_;
  assign new_n6074_ = new_n4595_ & new_n5803_;
  assign new_n6075_ = ~new_n6073_ & ~new_n6074_;
  assign new_n6076_ = new_n4655_ & new_n5755_;
  assign new_n6077_ = new_n4655_ & new_n5759_;
  assign new_n6078_ = ~new_n6076_ & ~new_n6077_;
  assign new_n6079_ = new_n6075_ & new_n6078_;
  assign new_n6080_ = new_n6072_ & new_n6079_;
  assign new_n6081_ = new_n4655_ & new_n5762_;
  assign new_n6082_ = new_n4655_ & new_n5768_;
  assign new_n6083_ = ~new_n6081_ & ~new_n6082_;
  assign new_n6084_ = new_n4655_ & new_n5770_;
  assign new_n6085_ = new_n4655_ & new_n5773_;
  assign new_n6086_ = ~new_n6084_ & ~new_n6085_;
  assign new_n6087_ = new_n6083_ & new_n6086_;
  assign new_n6088_ = new_n4655_ & new_n5783_;
  assign new_n6089_ = new_n4655_ & new_n5775_;
  assign new_n6090_ = new_n4655_ & new_n5781_;
  assign new_n6091_ = ~new_n6089_ & ~new_n6090_;
  assign new_n6092_ = ~new_n6088_ & new_n6091_;
  assign new_n6093_ = new_n6087_ & new_n6092_;
  assign new_n6094_ = new_n6080_ & new_n6093_;
  assign new_n6095_ = new_n4655_ & new_n5779_;
  assign new_n6096_ = new_n4655_ & new_n5789_;
  assign new_n6097_ = ~new_n6095_ & ~new_n6096_;
  assign new_n6098_ = new_n4655_ & new_n5791_;
  assign new_n6099_ = new_n4655_ & new_n5794_;
  assign new_n6100_ = ~new_n6098_ & ~new_n6099_;
  assign new_n6101_ = new_n6097_ & new_n6100_;
  assign new_n6102_ = new_n4655_ & new_n5803_;
  assign new_n6103_ = new_n4655_ & new_n5796_;
  assign new_n6104_ = new_n4655_ & new_n5801_;
  assign new_n6105_ = ~new_n6103_ & ~new_n6104_;
  assign new_n6106_ = ~new_n6102_ & new_n6105_;
  assign new_n6107_ = new_n6101_ & new_n6106_;
  assign new_n6108_ = new_n4682_ & new_n5755_;
  assign new_n6109_ = new_n4682_ & new_n5759_;
  assign new_n6110_ = ~new_n6108_ & ~new_n6109_;
  assign new_n6111_ = new_n4682_ & new_n5762_;
  assign new_n6112_ = new_n4682_ & new_n5768_;
  assign new_n6113_ = ~new_n6111_ & ~new_n6112_;
  assign new_n6114_ = new_n6110_ & new_n6113_;
  assign new_n6115_ = new_n4682_ & new_n5775_;
  assign new_n6116_ = new_n4682_ & new_n5770_;
  assign new_n6117_ = new_n4682_ & new_n5773_;
  assign new_n6118_ = ~new_n6116_ & ~new_n6117_;
  assign new_n6119_ = ~new_n6115_ & new_n6118_;
  assign new_n6120_ = new_n6114_ & new_n6119_;
  assign new_n6121_ = new_n6107_ & new_n6120_;
  assign new_n6122_ = new_n6094_ & new_n6121_;
  assign new_n6123_ = new_n4682_ & new_n5781_;
  assign new_n6124_ = new_n4682_ & new_n5783_;
  assign new_n6125_ = ~new_n6123_ & ~new_n6124_;
  assign new_n6126_ = new_n4682_ & new_n5779_;
  assign new_n6127_ = new_n4682_ & new_n5789_;
  assign new_n6128_ = ~new_n6126_ & ~new_n6127_;
  assign new_n6129_ = new_n6125_ & new_n6128_;
  assign new_n6130_ = new_n4682_ & new_n5791_;
  assign new_n6131_ = new_n4682_ & new_n5794_;
  assign new_n6132_ = ~new_n6130_ & ~new_n6131_;
  assign new_n6133_ = new_n4682_ & new_n5796_;
  assign new_n6134_ = new_n4682_ & new_n5801_;
  assign new_n6135_ = ~new_n6133_ & ~new_n6134_;
  assign new_n6136_ = new_n6132_ & new_n6135_;
  assign new_n6137_ = new_n6129_ & new_n6136_;
  assign new_n6138_ = new_n4682_ & new_n5803_;
  assign new_n6139_ = new_n4708_ & new_n5755_;
  assign new_n6140_ = ~new_n6138_ & ~new_n6139_;
  assign new_n6141_ = new_n4708_ & new_n5759_;
  assign new_n6142_ = new_n4708_ & new_n5762_;
  assign new_n6143_ = ~new_n6141_ & ~new_n6142_;
  assign new_n6144_ = new_n6140_ & new_n6143_;
  assign new_n6145_ = new_n4708_ & new_n5773_;
  assign new_n6146_ = new_n4708_ & new_n5768_;
  assign new_n6147_ = new_n4708_ & new_n5770_;
  assign new_n6148_ = ~new_n6146_ & ~new_n6147_;
  assign new_n6149_ = ~new_n6145_ & new_n6148_;
  assign new_n6150_ = new_n6144_ & new_n6149_;
  assign new_n6151_ = new_n6137_ & new_n6150_;
  assign new_n6152_ = new_n4708_ & new_n5775_;
  assign new_n6153_ = new_n4708_ & new_n5781_;
  assign new_n6154_ = ~new_n6152_ & ~new_n6153_;
  assign new_n6155_ = new_n4708_ & new_n5783_;
  assign new_n6156_ = new_n4708_ & new_n5779_;
  assign new_n6157_ = ~new_n6155_ & ~new_n6156_;
  assign new_n6158_ = new_n6154_ & new_n6157_;
  assign new_n6159_ = new_n4708_ & new_n5794_;
  assign new_n6160_ = new_n4708_ & new_n5789_;
  assign new_n6161_ = new_n4708_ & new_n5791_;
  assign new_n6162_ = ~new_n6160_ & ~new_n6161_;
  assign new_n6163_ = ~new_n6159_ & new_n6162_;
  assign new_n6164_ = new_n6158_ & new_n6163_;
  assign new_n6165_ = new_n4708_ & new_n5796_;
  assign new_n6166_ = new_n4708_ & new_n5801_;
  assign new_n6167_ = ~new_n6165_ & ~new_n6166_;
  assign new_n6168_ = new_n4708_ & new_n5803_;
  assign new_n6169_ = new_n4735_ & new_n5755_;
  assign new_n6170_ = ~new_n6168_ & ~new_n6169_;
  assign new_n6171_ = new_n6167_ & new_n6170_;
  assign new_n6172_ = new_n4735_ & new_n5768_;
  assign new_n6173_ = new_n4735_ & new_n5759_;
  assign new_n6174_ = new_n4735_ & new_n5762_;
  assign new_n6175_ = ~new_n6173_ & ~new_n6174_;
  assign new_n6176_ = ~new_n6172_ & new_n6175_;
  assign new_n6177_ = new_n6171_ & new_n6176_;
  assign new_n6178_ = new_n6164_ & new_n6177_;
  assign new_n6179_ = new_n6151_ & new_n6178_;
  assign new_n6180_ = new_n6122_ & new_n6179_;
  assign new_n6181_ = new_n6065_ & new_n6180_;
  assign new_n6182_ = new_n4735_ & new_n5770_;
  assign new_n6183_ = new_n4735_ & new_n5773_;
  assign new_n6184_ = ~new_n6182_ & ~new_n6183_;
  assign new_n6185_ = new_n4735_ & new_n5775_;
  assign new_n6186_ = new_n4735_ & new_n5781_;
  assign new_n6187_ = ~new_n6185_ & ~new_n6186_;
  assign new_n6188_ = new_n6184_ & new_n6187_;
  assign new_n6189_ = new_n4735_ & new_n5783_;
  assign new_n6190_ = new_n4735_ & new_n5779_;
  assign new_n6191_ = ~new_n6189_ & ~new_n6190_;
  assign new_n6192_ = new_n4735_ & new_n5789_;
  assign new_n6193_ = new_n4735_ & new_n5791_;
  assign new_n6194_ = ~new_n6192_ & ~new_n6193_;
  assign new_n6195_ = new_n6191_ & new_n6194_;
  assign new_n6196_ = new_n6188_ & new_n6195_;
  assign new_n6197_ = new_n4735_ & new_n5794_;
  assign new_n6198_ = new_n4735_ & new_n5796_;
  assign new_n6199_ = ~new_n6197_ & ~new_n6198_;
  assign new_n6200_ = new_n4735_ & new_n5801_;
  assign new_n6201_ = new_n4735_ & new_n5803_;
  assign new_n6202_ = ~new_n6200_ & ~new_n6201_;
  assign new_n6203_ = new_n6199_ & new_n6202_;
  assign new_n6204_ = new_n4826_ & new_n5755_;
  assign new_n6205_ = new_n1918_ & new_n5746_;
  assign new_n6206_ = new_n5745_ & new_n6205_;
  assign new_n6207_ = new_n1918_ & new_n5751_;
  assign new_n6208_ = new_n5745_ & new_n6207_;
  assign new_n6209_ = ~new_n6206_ & ~new_n6208_;
  assign new_n6210_ = ~new_n6204_ & new_n6209_;
  assign new_n6211_ = new_n6203_ & new_n6210_;
  assign new_n6212_ = new_n6196_ & new_n6211_;
  assign new_n6213_ = new_n4826_ & new_n5759_;
  assign new_n6214_ = new_n4826_ & new_n5762_;
  assign new_n6215_ = ~new_n6213_ & ~new_n6214_;
  assign new_n6216_ = new_n4826_ & new_n5768_;
  assign new_n6217_ = new_n4826_ & new_n5770_;
  assign new_n6218_ = ~new_n6216_ & ~new_n6217_;
  assign new_n6219_ = new_n6215_ & new_n6218_;
  assign new_n6220_ = new_n4826_ & new_n5781_;
  assign new_n6221_ = new_n4826_ & new_n5773_;
  assign new_n6222_ = new_n4826_ & new_n5775_;
  assign new_n6223_ = ~new_n6221_ & ~new_n6222_;
  assign new_n6224_ = ~new_n6220_ & new_n6223_;
  assign new_n6225_ = new_n6219_ & new_n6224_;
  assign new_n6226_ = new_n4826_ & new_n5783_;
  assign new_n6227_ = new_n4826_ & new_n5779_;
  assign new_n6228_ = ~new_n6226_ & ~new_n6227_;
  assign new_n6229_ = new_n4826_ & new_n5789_;
  assign new_n6230_ = new_n4826_ & new_n5791_;
  assign new_n6231_ = ~new_n6229_ & ~new_n6230_;
  assign new_n6232_ = new_n6228_ & new_n6231_;
  assign new_n6233_ = new_n4826_ & new_n5801_;
  assign new_n6234_ = new_n4826_ & new_n5794_;
  assign new_n6235_ = new_n4826_ & new_n5796_;
  assign new_n6236_ = ~new_n6234_ & ~new_n6235_;
  assign new_n6237_ = ~new_n6233_ & new_n6236_;
  assign new_n6238_ = new_n6232_ & new_n6237_;
  assign new_n6239_ = new_n6225_ & new_n6238_;
  assign new_n6240_ = new_n6212_ & new_n6239_;
  assign new_n6241_ = new_n4826_ & new_n5803_;
  assign new_n6242_ = new_n4847_ & new_n5755_;
  assign new_n6243_ = ~new_n6241_ & ~new_n6242_;
  assign new_n6244_ = new_n4847_ & new_n5759_;
  assign new_n6245_ = new_n4847_ & new_n5762_;
  assign new_n6246_ = ~new_n6244_ & ~new_n6245_;
  assign new_n6247_ = new_n6243_ & new_n6246_;
  assign new_n6248_ = new_n4847_ & new_n5768_;
  assign new_n6249_ = new_n4847_ & new_n5770_;
  assign new_n6250_ = ~new_n6248_ & ~new_n6249_;
  assign new_n6251_ = new_n4847_ & new_n5773_;
  assign new_n6252_ = new_n4847_ & new_n5775_;
  assign new_n6253_ = ~new_n6251_ & ~new_n6252_;
  assign new_n6254_ = new_n6250_ & new_n6253_;
  assign new_n6255_ = new_n6247_ & new_n6254_;
  assign new_n6256_ = new_n4847_ & new_n5781_;
  assign new_n6257_ = new_n4847_ & new_n5783_;
  assign new_n6258_ = ~new_n6256_ & ~new_n6257_;
  assign new_n6259_ = new_n4847_ & new_n5779_;
  assign new_n6260_ = new_n4847_ & new_n5789_;
  assign new_n6261_ = ~new_n6259_ & ~new_n6260_;
  assign new_n6262_ = new_n6258_ & new_n6261_;
  assign new_n6263_ = new_n4847_ & new_n5796_;
  assign new_n6264_ = new_n4847_ & new_n5791_;
  assign new_n6265_ = new_n4847_ & new_n5794_;
  assign new_n6266_ = ~new_n6264_ & ~new_n6265_;
  assign new_n6267_ = ~new_n6263_ & new_n6266_;
  assign new_n6268_ = new_n6262_ & new_n6267_;
  assign new_n6269_ = new_n6255_ & new_n6268_;
  assign new_n6270_ = new_n4847_ & new_n5801_;
  assign new_n6271_ = new_n4847_ & new_n5803_;
  assign new_n6272_ = ~new_n6270_ & ~new_n6271_;
  assign new_n6273_ = new_n4906_ & new_n5755_;
  assign new_n6274_ = new_n4906_ & new_n5759_;
  assign new_n6275_ = ~new_n6273_ & ~new_n6274_;
  assign new_n6276_ = new_n6272_ & new_n6275_;
  assign new_n6277_ = new_n4906_ & new_n5770_;
  assign new_n6278_ = new_n4906_ & new_n5762_;
  assign new_n6279_ = new_n4906_ & new_n5768_;
  assign new_n6280_ = ~new_n6278_ & ~new_n6279_;
  assign new_n6281_ = ~new_n6277_ & new_n6280_;
  assign new_n6282_ = new_n6276_ & new_n6281_;
  assign new_n6283_ = new_n4906_ & new_n5773_;
  assign new_n6284_ = new_n4906_ & new_n5775_;
  assign new_n6285_ = ~new_n6283_ & ~new_n6284_;
  assign new_n6286_ = new_n4906_ & new_n5781_;
  assign new_n6287_ = new_n4906_ & new_n5783_;
  assign new_n6288_ = ~new_n6286_ & ~new_n6287_;
  assign new_n6289_ = new_n6285_ & new_n6288_;
  assign new_n6290_ = new_n4906_ & new_n5791_;
  assign new_n6291_ = new_n4906_ & new_n5779_;
  assign new_n6292_ = new_n4906_ & new_n5789_;
  assign new_n6293_ = ~new_n6291_ & ~new_n6292_;
  assign new_n6294_ = ~new_n6290_ & new_n6293_;
  assign new_n6295_ = new_n6289_ & new_n6294_;
  assign new_n6296_ = new_n6282_ & new_n6295_;
  assign new_n6297_ = new_n6269_ & new_n6296_;
  assign new_n6298_ = new_n6240_ & new_n6297_;
  assign new_n6299_ = new_n4906_ & new_n5794_;
  assign new_n6300_ = new_n4906_ & new_n5796_;
  assign new_n6301_ = ~new_n6299_ & ~new_n6300_;
  assign new_n6302_ = new_n4906_ & new_n5801_;
  assign new_n6303_ = new_n4906_ & new_n5803_;
  assign new_n6304_ = ~new_n6302_ & ~new_n6303_;
  assign new_n6305_ = new_n6301_ & new_n6304_;
  assign new_n6306_ = new_n4934_ & new_n5755_;
  assign new_n6307_ = new_n4934_ & new_n5759_;
  assign new_n6308_ = ~new_n6306_ & ~new_n6307_;
  assign new_n6309_ = new_n4934_ & new_n5762_;
  assign new_n6310_ = new_n4934_ & new_n5768_;
  assign new_n6311_ = ~new_n6309_ & ~new_n6310_;
  assign new_n6312_ = new_n6308_ & new_n6311_;
  assign new_n6313_ = new_n6305_ & new_n6312_;
  assign new_n6314_ = new_n4934_ & new_n5770_;
  assign new_n6315_ = new_n4934_ & new_n5773_;
  assign new_n6316_ = ~new_n6314_ & ~new_n6315_;
  assign new_n6317_ = new_n4934_ & new_n5775_;
  assign new_n6318_ = new_n4934_ & new_n5781_;
  assign new_n6319_ = ~new_n6317_ & ~new_n6318_;
  assign new_n6320_ = new_n6316_ & new_n6319_;
  assign new_n6321_ = new_n4934_ & new_n5789_;
  assign new_n6322_ = new_n4934_ & new_n5783_;
  assign new_n6323_ = new_n4934_ & new_n5779_;
  assign new_n6324_ = ~new_n6322_ & ~new_n6323_;
  assign new_n6325_ = ~new_n6321_ & new_n6324_;
  assign new_n6326_ = new_n6320_ & new_n6325_;
  assign new_n6327_ = new_n6313_ & new_n6326_;
  assign new_n6328_ = new_n4934_ & new_n5791_;
  assign new_n6329_ = new_n4934_ & new_n5794_;
  assign new_n6330_ = ~new_n6328_ & ~new_n6329_;
  assign new_n6331_ = new_n4934_ & new_n5796_;
  assign new_n6332_ = new_n4934_ & new_n5801_;
  assign new_n6333_ = ~new_n6331_ & ~new_n6332_;
  assign new_n6334_ = new_n6330_ & new_n6333_;
  assign new_n6335_ = new_n1905_ & new_n5909_;
  assign new_n6336_ = new_n5745_ & new_n6335_;
  assign new_n6337_ = new_n4934_ & new_n5803_;
  assign new_n6338_ = new_n1905_ & new_n5900_;
  assign new_n6339_ = new_n5745_ & new_n6338_;
  assign new_n6340_ = ~new_n6337_ & ~new_n6339_;
  assign new_n6341_ = ~new_n6336_ & new_n6340_;
  assign new_n6342_ = new_n6334_ & new_n6341_;
  assign new_n6343_ = ~A170 & new_n5905_;
  assign new_n6344_ = new_n2839_ & new_n6343_;
  assign new_n6345_ = new_n5745_ & new_n6344_;
  assign new_n6346_ = new_n2871_ & new_n6343_;
  assign new_n6347_ = new_n5745_ & new_n6346_;
  assign new_n6348_ = ~new_n6345_ & ~new_n6347_;
  assign new_n6349_ = new_n2896_ & new_n6343_;
  assign new_n6350_ = new_n5745_ & new_n6349_;
  assign new_n6351_ = new_n2920_ & new_n6343_;
  assign new_n6352_ = new_n5745_ & new_n6351_;
  assign new_n6353_ = ~new_n6350_ & ~new_n6352_;
  assign new_n6354_ = new_n6348_ & new_n6353_;
  assign new_n6355_ = new_n4956_ & new_n5576_;
  assign new_n6356_ = new_n4956_ & new_n5578_;
  assign new_n6357_ = new_n4956_ & new_n5580_;
  assign new_n6358_ = ~new_n6356_ & ~new_n6357_;
  assign new_n6359_ = ~new_n6355_ & new_n6358_;
  assign new_n6360_ = new_n6354_ & new_n6359_;
  assign new_n6361_ = new_n6342_ & new_n6360_;
  assign new_n6362_ = new_n6327_ & new_n6361_;
  assign new_n6363_ = new_n4956_ & new_n5587_;
  assign new_n6364_ = new_n4956_ & new_n5590_;
  assign new_n6365_ = ~new_n6363_ & ~new_n6364_;
  assign new_n6366_ = new_n4956_ & new_n5594_;
  assign new_n6367_ = new_n4963_ & new_n5596_;
  assign new_n6368_ = ~new_n6366_ & ~new_n6367_;
  assign new_n6369_ = new_n6365_ & new_n6368_;
  assign new_n6370_ = new_n4963_ & new_n5605_;
  assign new_n6371_ = new_n4963_ & new_n5600_;
  assign new_n6372_ = new_n4963_ & new_n5602_;
  assign new_n6373_ = ~new_n6371_ & ~new_n6372_;
  assign new_n6374_ = ~new_n6370_ & new_n6373_;
  assign new_n6375_ = new_n6369_ & new_n6374_;
  assign new_n6376_ = new_n4963_ & new_n5608_;
  assign new_n6377_ = new_n4963_ & new_n5614_;
  assign new_n6378_ = ~new_n6376_ & ~new_n6377_;
  assign new_n6379_ = new_n4965_ & new_n5755_;
  assign new_n6380_ = new_n4965_ & new_n5759_;
  assign new_n6381_ = ~new_n6379_ & ~new_n6380_;
  assign new_n6382_ = new_n6378_ & new_n6381_;
  assign new_n6383_ = new_n4965_ & new_n5770_;
  assign new_n6384_ = new_n4965_ & new_n5762_;
  assign new_n6385_ = new_n4965_ & new_n5768_;
  assign new_n6386_ = ~new_n6384_ & ~new_n6385_;
  assign new_n6387_ = ~new_n6383_ & new_n6386_;
  assign new_n6388_ = new_n6382_ & new_n6387_;
  assign new_n6389_ = new_n6375_ & new_n6388_;
  assign new_n6390_ = new_n4965_ & new_n5773_;
  assign new_n6391_ = new_n4965_ & new_n5775_;
  assign new_n6392_ = ~new_n6390_ & ~new_n6391_;
  assign new_n6393_ = new_n4965_ & new_n5781_;
  assign new_n6394_ = new_n4965_ & new_n5783_;
  assign new_n6395_ = ~new_n6393_ & ~new_n6394_;
  assign new_n6396_ = new_n6392_ & new_n6395_;
  assign new_n6397_ = new_n4965_ & new_n5791_;
  assign new_n6398_ = new_n4965_ & new_n5779_;
  assign new_n6399_ = new_n4965_ & new_n5789_;
  assign new_n6400_ = ~new_n6398_ & ~new_n6399_;
  assign new_n6401_ = ~new_n6397_ & new_n6400_;
  assign new_n6402_ = new_n6396_ & new_n6401_;
  assign new_n6403_ = new_n4965_ & new_n5794_;
  assign new_n6404_ = new_n4965_ & new_n5796_;
  assign new_n6405_ = ~new_n6403_ & ~new_n6404_;
  assign new_n6406_ = new_n4965_ & new_n5801_;
  assign new_n6407_ = new_n4965_ & new_n5803_;
  assign new_n6408_ = ~new_n6406_ & ~new_n6407_;
  assign new_n6409_ = new_n6405_ & new_n6408_;
  assign new_n6410_ = new_n4990_ & new_n5762_;
  assign new_n6411_ = new_n4990_ & new_n5755_;
  assign new_n6412_ = new_n4990_ & new_n5759_;
  assign new_n6413_ = ~new_n6411_ & ~new_n6412_;
  assign new_n6414_ = ~new_n6410_ & new_n6413_;
  assign new_n6415_ = new_n6409_ & new_n6414_;
  assign new_n6416_ = new_n6402_ & new_n6415_;
  assign new_n6417_ = new_n6389_ & new_n6416_;
  assign new_n6418_ = new_n6362_ & new_n6417_;
  assign new_n6419_ = new_n6298_ & new_n6418_;
  assign new_n6420_ = new_n6181_ & new_n6419_;
  assign new_n6421_ = new_n5950_ & new_n6420_;
  assign new_n6422_ = new_n5399_ & new_n6421_;
  assign new_n6423_ = new_n4990_ & new_n5768_;
  assign new_n6424_ = new_n4990_ & new_n5770_;
  assign new_n6425_ = ~new_n6423_ & ~new_n6424_;
  assign new_n6426_ = new_n4990_ & new_n5773_;
  assign new_n6427_ = new_n4990_ & new_n5775_;
  assign new_n6428_ = ~new_n6426_ & ~new_n6427_;
  assign new_n6429_ = new_n6425_ & new_n6428_;
  assign new_n6430_ = new_n4990_ & new_n5781_;
  assign new_n6431_ = new_n4990_ & new_n5783_;
  assign new_n6432_ = ~new_n6430_ & ~new_n6431_;
  assign new_n6433_ = new_n4990_ & new_n5779_;
  assign new_n6434_ = new_n4990_ & new_n5789_;
  assign new_n6435_ = ~new_n6433_ & ~new_n6434_;
  assign new_n6436_ = new_n6432_ & new_n6435_;
  assign new_n6437_ = new_n6429_ & new_n6436_;
  assign new_n6438_ = new_n4990_ & new_n5791_;
  assign new_n6439_ = new_n4990_ & new_n5794_;
  assign new_n6440_ = ~new_n6438_ & ~new_n6439_;
  assign new_n6441_ = new_n4990_ & new_n5796_;
  assign new_n6442_ = new_n4990_ & new_n5801_;
  assign new_n6443_ = ~new_n6441_ & ~new_n6442_;
  assign new_n6444_ = new_n6440_ & new_n6443_;
  assign new_n6445_ = new_n5014_ & new_n5759_;
  assign new_n6446_ = new_n4990_ & new_n5803_;
  assign new_n6447_ = new_n5014_ & new_n5755_;
  assign new_n6448_ = ~new_n6446_ & ~new_n6447_;
  assign new_n6449_ = ~new_n6445_ & new_n6448_;
  assign new_n6450_ = new_n6444_ & new_n6449_;
  assign new_n6451_ = new_n6437_ & new_n6450_;
  assign new_n6452_ = new_n5014_ & new_n5762_;
  assign new_n6453_ = new_n5014_ & new_n5768_;
  assign new_n6454_ = ~new_n6452_ & ~new_n6453_;
  assign new_n6455_ = new_n5014_ & new_n5770_;
  assign new_n6456_ = new_n5014_ & new_n5773_;
  assign new_n6457_ = ~new_n6455_ & ~new_n6456_;
  assign new_n6458_ = new_n6454_ & new_n6457_;
  assign new_n6459_ = new_n5014_ & new_n5783_;
  assign new_n6460_ = new_n5014_ & new_n5775_;
  assign new_n6461_ = new_n5014_ & new_n5781_;
  assign new_n6462_ = ~new_n6460_ & ~new_n6461_;
  assign new_n6463_ = ~new_n6459_ & new_n6462_;
  assign new_n6464_ = new_n6458_ & new_n6463_;
  assign new_n6465_ = new_n5014_ & new_n5779_;
  assign new_n6466_ = new_n5014_ & new_n5789_;
  assign new_n6467_ = ~new_n6465_ & ~new_n6466_;
  assign new_n6468_ = new_n5014_ & new_n5791_;
  assign new_n6469_ = new_n5014_ & new_n5794_;
  assign new_n6470_ = ~new_n6468_ & ~new_n6469_;
  assign new_n6471_ = new_n6467_ & new_n6470_;
  assign new_n6472_ = new_n5014_ & new_n5803_;
  assign new_n6473_ = new_n5014_ & new_n5796_;
  assign new_n6474_ = new_n5014_ & new_n5801_;
  assign new_n6475_ = ~new_n6473_ & ~new_n6474_;
  assign new_n6476_ = ~new_n6472_ & new_n6475_;
  assign new_n6477_ = new_n6471_ & new_n6476_;
  assign new_n6478_ = new_n6464_ & new_n6477_;
  assign new_n6479_ = new_n6451_ & new_n6478_;
  assign new_n6480_ = new_n5041_ & new_n5755_;
  assign new_n6481_ = new_n5041_ & new_n5759_;
  assign new_n6482_ = ~new_n6480_ & ~new_n6481_;
  assign new_n6483_ = new_n5041_ & new_n5762_;
  assign new_n6484_ = new_n5041_ & new_n5768_;
  assign new_n6485_ = ~new_n6483_ & ~new_n6484_;
  assign new_n6486_ = new_n6482_ & new_n6485_;
  assign new_n6487_ = new_n5041_ & new_n5770_;
  assign new_n6488_ = new_n5041_ & new_n5773_;
  assign new_n6489_ = ~new_n6487_ & ~new_n6488_;
  assign new_n6490_ = new_n5041_ & new_n5775_;
  assign new_n6491_ = new_n5041_ & new_n5781_;
  assign new_n6492_ = ~new_n6490_ & ~new_n6491_;
  assign new_n6493_ = new_n6489_ & new_n6492_;
  assign new_n6494_ = new_n6486_ & new_n6493_;
  assign new_n6495_ = new_n5041_ & new_n5783_;
  assign new_n6496_ = new_n5041_ & new_n5779_;
  assign new_n6497_ = ~new_n6495_ & ~new_n6496_;
  assign new_n6498_ = new_n5041_ & new_n5789_;
  assign new_n6499_ = new_n5041_ & new_n5791_;
  assign new_n6500_ = ~new_n6498_ & ~new_n6499_;
  assign new_n6501_ = new_n6497_ & new_n6500_;
  assign new_n6502_ = new_n5041_ & new_n5801_;
  assign new_n6503_ = new_n5041_ & new_n5794_;
  assign new_n6504_ = new_n5041_ & new_n5796_;
  assign new_n6505_ = ~new_n6503_ & ~new_n6504_;
  assign new_n6506_ = ~new_n6502_ & new_n6505_;
  assign new_n6507_ = new_n6501_ & new_n6506_;
  assign new_n6508_ = new_n6494_ & new_n6507_;
  assign new_n6509_ = new_n5041_ & new_n5803_;
  assign new_n6510_ = new_n5099_ & new_n5755_;
  assign new_n6511_ = ~new_n6509_ & ~new_n6510_;
  assign new_n6512_ = new_n5099_ & new_n5759_;
  assign new_n6513_ = new_n5099_ & new_n5762_;
  assign new_n6514_ = ~new_n6512_ & ~new_n6513_;
  assign new_n6515_ = new_n6511_ & new_n6514_;
  assign new_n6516_ = new_n5099_ & new_n5773_;
  assign new_n6517_ = new_n5099_ & new_n5768_;
  assign new_n6518_ = new_n5099_ & new_n5770_;
  assign new_n6519_ = ~new_n6517_ & ~new_n6518_;
  assign new_n6520_ = ~new_n6516_ & new_n6519_;
  assign new_n6521_ = new_n6515_ & new_n6520_;
  assign new_n6522_ = new_n5099_ & new_n5775_;
  assign new_n6523_ = new_n5099_ & new_n5781_;
  assign new_n6524_ = ~new_n6522_ & ~new_n6523_;
  assign new_n6525_ = new_n5099_ & new_n5783_;
  assign new_n6526_ = new_n5099_ & new_n5779_;
  assign new_n6527_ = ~new_n6525_ & ~new_n6526_;
  assign new_n6528_ = new_n6524_ & new_n6527_;
  assign new_n6529_ = new_n5099_ & new_n5794_;
  assign new_n6530_ = new_n5099_ & new_n5789_;
  assign new_n6531_ = new_n5099_ & new_n5791_;
  assign new_n6532_ = ~new_n6530_ & ~new_n6531_;
  assign new_n6533_ = ~new_n6529_ & new_n6532_;
  assign new_n6534_ = new_n6528_ & new_n6533_;
  assign new_n6535_ = new_n6521_ & new_n6534_;
  assign new_n6536_ = new_n6508_ & new_n6535_;
  assign new_n6537_ = new_n6479_ & new_n6536_;
  assign new_n6538_ = new_n5099_ & new_n5796_;
  assign new_n6539_ = new_n5099_ & new_n5801_;
  assign new_n6540_ = ~new_n6538_ & ~new_n6539_;
  assign new_n6541_ = new_n5099_ & new_n5803_;
  assign new_n6542_ = new_n5122_ & new_n5755_;
  assign new_n6543_ = ~new_n6541_ & ~new_n6542_;
  assign new_n6544_ = new_n6540_ & new_n6543_;
  assign new_n6545_ = new_n5122_ & new_n5759_;
  assign new_n6546_ = new_n5122_ & new_n5762_;
  assign new_n6547_ = ~new_n6545_ & ~new_n6546_;
  assign new_n6548_ = new_n5122_ & new_n5768_;
  assign new_n6549_ = new_n5122_ & new_n5770_;
  assign new_n6550_ = ~new_n6548_ & ~new_n6549_;
  assign new_n6551_ = new_n6547_ & new_n6550_;
  assign new_n6552_ = new_n6544_ & new_n6551_;
  assign new_n6553_ = new_n5122_ & new_n5773_;
  assign new_n6554_ = new_n5122_ & new_n5775_;
  assign new_n6555_ = ~new_n6553_ & ~new_n6554_;
  assign new_n6556_ = new_n5122_ & new_n5781_;
  assign new_n6557_ = new_n5122_ & new_n5783_;
  assign new_n6558_ = ~new_n6556_ & ~new_n6557_;
  assign new_n6559_ = new_n6555_ & new_n6558_;
  assign new_n6560_ = new_n5122_ & new_n5791_;
  assign new_n6561_ = new_n5122_ & new_n5779_;
  assign new_n6562_ = new_n5122_ & new_n5789_;
  assign new_n6563_ = ~new_n6561_ & ~new_n6562_;
  assign new_n6564_ = ~new_n6560_ & new_n6563_;
  assign new_n6565_ = new_n6559_ & new_n6564_;
  assign new_n6566_ = new_n6552_ & new_n6565_;
  assign new_n6567_ = new_n5122_ & new_n5794_;
  assign new_n6568_ = new_n5122_ & new_n5796_;
  assign new_n6569_ = ~new_n6567_ & ~new_n6568_;
  assign new_n6570_ = new_n5122_ & new_n5801_;
  assign new_n6571_ = new_n5122_ & new_n5803_;
  assign new_n6572_ = ~new_n6570_ & ~new_n6571_;
  assign new_n6573_ = new_n6569_ & new_n6572_;
  assign new_n6574_ = new_n5146_ & new_n5762_;
  assign new_n6575_ = new_n5146_ & new_n5755_;
  assign new_n6576_ = new_n5146_ & new_n5759_;
  assign new_n6577_ = ~new_n6575_ & ~new_n6576_;
  assign new_n6578_ = ~new_n6574_ & new_n6577_;
  assign new_n6579_ = new_n6573_ & new_n6578_;
  assign new_n6580_ = new_n5146_ & new_n5768_;
  assign new_n6581_ = new_n5146_ & new_n5770_;
  assign new_n6582_ = ~new_n6580_ & ~new_n6581_;
  assign new_n6583_ = new_n5146_ & new_n5773_;
  assign new_n6584_ = new_n5146_ & new_n5775_;
  assign new_n6585_ = ~new_n6583_ & ~new_n6584_;
  assign new_n6586_ = new_n6582_ & new_n6585_;
  assign new_n6587_ = new_n5146_ & new_n5779_;
  assign new_n6588_ = new_n5146_ & new_n5781_;
  assign new_n6589_ = new_n5146_ & new_n5783_;
  assign new_n6590_ = ~new_n6588_ & ~new_n6589_;
  assign new_n6591_ = ~new_n6587_ & new_n6590_;
  assign new_n6592_ = new_n6586_ & new_n6591_;
  assign new_n6593_ = new_n6579_ & new_n6592_;
  assign new_n6594_ = new_n6566_ & new_n6593_;
  assign new_n6595_ = new_n5146_ & new_n5789_;
  assign new_n6596_ = new_n5146_ & new_n5791_;
  assign new_n6597_ = ~new_n6595_ & ~new_n6596_;
  assign new_n6598_ = new_n5146_ & new_n5794_;
  assign new_n6599_ = new_n5146_ & new_n5796_;
  assign new_n6600_ = ~new_n6598_ & ~new_n6599_;
  assign new_n6601_ = new_n6597_ & new_n6600_;
  assign new_n6602_ = new_n5146_ & new_n5801_;
  assign new_n6603_ = new_n5146_ & new_n5803_;
  assign new_n6604_ = ~new_n6602_ & ~new_n6603_;
  assign new_n6605_ = new_n5172_ & new_n5755_;
  assign new_n6606_ = new_n5172_ & new_n5759_;
  assign new_n6607_ = ~new_n6605_ & ~new_n6606_;
  assign new_n6608_ = new_n6604_ & new_n6607_;
  assign new_n6609_ = new_n6601_ & new_n6608_;
  assign new_n6610_ = new_n5172_ & new_n5762_;
  assign new_n6611_ = new_n5172_ & new_n5768_;
  assign new_n6612_ = ~new_n6610_ & ~new_n6611_;
  assign new_n6613_ = new_n5172_ & new_n5770_;
  assign new_n6614_ = new_n5172_ & new_n5773_;
  assign new_n6615_ = ~new_n6613_ & ~new_n6614_;
  assign new_n6616_ = new_n6612_ & new_n6615_;
  assign new_n6617_ = new_n5172_ & new_n5783_;
  assign new_n6618_ = new_n5172_ & new_n5775_;
  assign new_n6619_ = new_n5172_ & new_n5781_;
  assign new_n6620_ = ~new_n6618_ & ~new_n6619_;
  assign new_n6621_ = ~new_n6617_ & new_n6620_;
  assign new_n6622_ = new_n6616_ & new_n6621_;
  assign new_n6623_ = new_n6609_ & new_n6622_;
  assign new_n6624_ = new_n5172_ & new_n5779_;
  assign new_n6625_ = new_n5172_ & new_n5789_;
  assign new_n6626_ = ~new_n6624_ & ~new_n6625_;
  assign new_n6627_ = new_n5172_ & new_n5791_;
  assign new_n6628_ = new_n5172_ & new_n5794_;
  assign new_n6629_ = ~new_n6627_ & ~new_n6628_;
  assign new_n6630_ = new_n6626_ & new_n6629_;
  assign new_n6631_ = new_n5172_ & new_n5803_;
  assign new_n6632_ = new_n5172_ & new_n5796_;
  assign new_n6633_ = new_n5172_ & new_n5801_;
  assign new_n6634_ = ~new_n6632_ & ~new_n6633_;
  assign new_n6635_ = ~new_n6631_ & new_n6634_;
  assign new_n6636_ = new_n6630_ & new_n6635_;
  assign new_n6637_ = new_n2265_ & new_n5746_;
  assign new_n6638_ = new_n5745_ & new_n6637_;
  assign new_n6639_ = new_n2265_ & new_n5751_;
  assign new_n6640_ = new_n5745_ & new_n6639_;
  assign new_n6641_ = ~new_n6638_ & ~new_n6640_;
  assign new_n6642_ = new_n5263_ & new_n5755_;
  assign new_n6643_ = new_n5263_ & new_n5759_;
  assign new_n6644_ = ~new_n6642_ & ~new_n6643_;
  assign new_n6645_ = new_n6641_ & new_n6644_;
  assign new_n6646_ = new_n5263_ & new_n5770_;
  assign new_n6647_ = new_n5263_ & new_n5762_;
  assign new_n6648_ = new_n5263_ & new_n5768_;
  assign new_n6649_ = ~new_n6647_ & ~new_n6648_;
  assign new_n6650_ = ~new_n6646_ & new_n6649_;
  assign new_n6651_ = new_n6645_ & new_n6650_;
  assign new_n6652_ = new_n6636_ & new_n6651_;
  assign new_n6653_ = new_n6623_ & new_n6652_;
  assign new_n6654_ = new_n6594_ & new_n6653_;
  assign new_n6655_ = new_n6537_ & new_n6654_;
  assign new_n6656_ = new_n5263_ & new_n5773_;
  assign new_n6657_ = new_n5263_ & new_n5775_;
  assign new_n6658_ = ~new_n6656_ & ~new_n6657_;
  assign new_n6659_ = new_n5263_ & new_n5781_;
  assign new_n6660_ = new_n5263_ & new_n5783_;
  assign new_n6661_ = ~new_n6659_ & ~new_n6660_;
  assign new_n6662_ = new_n6658_ & new_n6661_;
  assign new_n6663_ = new_n5263_ & new_n5779_;
  assign new_n6664_ = new_n5263_ & new_n5789_;
  assign new_n6665_ = ~new_n6663_ & ~new_n6664_;
  assign new_n6666_ = new_n5263_ & new_n5791_;
  assign new_n6667_ = new_n5263_ & new_n5794_;
  assign new_n6668_ = ~new_n6666_ & ~new_n6667_;
  assign new_n6669_ = new_n6665_ & new_n6668_;
  assign new_n6670_ = new_n6662_ & new_n6669_;
  assign new_n6671_ = new_n5263_ & new_n5796_;
  assign new_n6672_ = new_n5263_ & new_n5801_;
  assign new_n6673_ = ~new_n6671_ & ~new_n6672_;
  assign new_n6674_ = new_n5263_ & new_n5803_;
  assign new_n6675_ = new_n5288_ & new_n5755_;
  assign new_n6676_ = ~new_n6674_ & ~new_n6675_;
  assign new_n6677_ = new_n6673_ & new_n6676_;
  assign new_n6678_ = new_n5288_ & new_n5768_;
  assign new_n6679_ = new_n5288_ & new_n5759_;
  assign new_n6680_ = new_n5288_ & new_n5762_;
  assign new_n6681_ = ~new_n6679_ & ~new_n6680_;
  assign new_n6682_ = ~new_n6678_ & new_n6681_;
  assign new_n6683_ = new_n6677_ & new_n6682_;
  assign new_n6684_ = new_n6670_ & new_n6683_;
  assign new_n6685_ = new_n5288_ & new_n5770_;
  assign new_n6686_ = new_n5288_ & new_n5773_;
  assign new_n6687_ = ~new_n6685_ & ~new_n6686_;
  assign new_n6688_ = new_n5288_ & new_n5775_;
  assign new_n6689_ = new_n5288_ & new_n5781_;
  assign new_n6690_ = ~new_n6688_ & ~new_n6689_;
  assign new_n6691_ = new_n6687_ & new_n6690_;
  assign new_n6692_ = new_n5288_ & new_n5789_;
  assign new_n6693_ = new_n5288_ & new_n5783_;
  assign new_n6694_ = new_n5288_ & new_n5779_;
  assign new_n6695_ = ~new_n6693_ & ~new_n6694_;
  assign new_n6696_ = ~new_n6692_ & new_n6695_;
  assign new_n6697_ = new_n6691_ & new_n6696_;
  assign new_n6698_ = new_n5288_ & new_n5791_;
  assign new_n6699_ = new_n5288_ & new_n5794_;
  assign new_n6700_ = ~new_n6698_ & ~new_n6699_;
  assign new_n6701_ = new_n5288_ & new_n5796_;
  assign new_n6702_ = new_n5288_ & new_n5801_;
  assign new_n6703_ = ~new_n6701_ & ~new_n6702_;
  assign new_n6704_ = new_n6700_ & new_n6703_;
  assign new_n6705_ = new_n5346_ & new_n5759_;
  assign new_n6706_ = new_n5288_ & new_n5803_;
  assign new_n6707_ = new_n5346_ & new_n5755_;
  assign new_n6708_ = ~new_n6706_ & ~new_n6707_;
  assign new_n6709_ = ~new_n6705_ & new_n6708_;
  assign new_n6710_ = new_n6704_ & new_n6709_;
  assign new_n6711_ = new_n6697_ & new_n6710_;
  assign new_n6712_ = new_n6684_ & new_n6711_;
  assign new_n6713_ = new_n5346_ & new_n5762_;
  assign new_n6714_ = new_n5346_ & new_n5768_;
  assign new_n6715_ = ~new_n6713_ & ~new_n6714_;
  assign new_n6716_ = new_n5346_ & new_n5770_;
  assign new_n6717_ = new_n5346_ & new_n5773_;
  assign new_n6718_ = ~new_n6716_ & ~new_n6717_;
  assign new_n6719_ = new_n6715_ & new_n6718_;
  assign new_n6720_ = new_n5346_ & new_n5775_;
  assign new_n6721_ = new_n5346_ & new_n5781_;
  assign new_n6722_ = ~new_n6720_ & ~new_n6721_;
  assign new_n6723_ = new_n5346_ & new_n5783_;
  assign new_n6724_ = new_n5346_ & new_n5779_;
  assign new_n6725_ = ~new_n6723_ & ~new_n6724_;
  assign new_n6726_ = new_n6722_ & new_n6725_;
  assign new_n6727_ = new_n6719_ & new_n6726_;
  assign new_n6728_ = new_n5346_ & new_n5789_;
  assign new_n6729_ = new_n5346_ & new_n5791_;
  assign new_n6730_ = ~new_n6728_ & ~new_n6729_;
  assign new_n6731_ = new_n5346_ & new_n5794_;
  assign new_n6732_ = new_n5346_ & new_n5796_;
  assign new_n6733_ = ~new_n6731_ & ~new_n6732_;
  assign new_n6734_ = new_n6730_ & new_n6733_;
  assign new_n6735_ = new_n5370_ & new_n5755_;
  assign new_n6736_ = new_n5346_ & new_n5801_;
  assign new_n6737_ = new_n5346_ & new_n5803_;
  assign new_n6738_ = ~new_n6736_ & ~new_n6737_;
  assign new_n6739_ = ~new_n6735_ & new_n6738_;
  assign new_n6740_ = new_n6734_ & new_n6739_;
  assign new_n6741_ = new_n6727_ & new_n6740_;
  assign new_n6742_ = new_n5370_ & new_n5759_;
  assign new_n6743_ = new_n5370_ & new_n5762_;
  assign new_n6744_ = ~new_n6742_ & ~new_n6743_;
  assign new_n6745_ = new_n5370_ & new_n5768_;
  assign new_n6746_ = new_n5370_ & new_n5770_;
  assign new_n6747_ = ~new_n6745_ & ~new_n6746_;
  assign new_n6748_ = new_n6744_ & new_n6747_;
  assign new_n6749_ = new_n5370_ & new_n5781_;
  assign new_n6750_ = new_n5370_ & new_n5773_;
  assign new_n6751_ = new_n5370_ & new_n5775_;
  assign new_n6752_ = ~new_n6750_ & ~new_n6751_;
  assign new_n6753_ = ~new_n6749_ & new_n6752_;
  assign new_n6754_ = new_n6748_ & new_n6753_;
  assign new_n6755_ = new_n5370_ & new_n5783_;
  assign new_n6756_ = new_n5370_ & new_n5779_;
  assign new_n6757_ = ~new_n6755_ & ~new_n6756_;
  assign new_n6758_ = new_n5370_ & new_n5789_;
  assign new_n6759_ = new_n5370_ & new_n5791_;
  assign new_n6760_ = ~new_n6758_ & ~new_n6759_;
  assign new_n6761_ = new_n6757_ & new_n6760_;
  assign new_n6762_ = new_n5370_ & new_n5801_;
  assign new_n6763_ = new_n5370_ & new_n5794_;
  assign new_n6764_ = new_n5370_ & new_n5796_;
  assign new_n6765_ = ~new_n6763_ & ~new_n6764_;
  assign new_n6766_ = ~new_n6762_ & new_n6765_;
  assign new_n6767_ = new_n6761_ & new_n6766_;
  assign new_n6768_ = new_n6754_ & new_n6767_;
  assign new_n6769_ = new_n6741_ & new_n6768_;
  assign new_n6770_ = new_n6712_ & new_n6769_;
  assign new_n6771_ = new_n5370_ & new_n5803_;
  assign new_n6772_ = new_n2260_ & new_n5900_;
  assign new_n6773_ = new_n5745_ & new_n6772_;
  assign new_n6774_ = ~new_n6771_ & ~new_n6773_;
  assign new_n6775_ = new_n2260_ & new_n5909_;
  assign new_n6776_ = new_n5745_ & new_n6775_;
  assign new_n6777_ = ~A167 & new_n3192_;
  assign new_n6778_ = new_n2839_ & new_n6777_;
  assign new_n6779_ = new_n5745_ & new_n6778_;
  assign new_n6780_ = ~new_n6776_ & ~new_n6779_;
  assign new_n6781_ = new_n6774_ & new_n6780_;
  assign new_n6782_ = new_n2871_ & new_n6777_;
  assign new_n6783_ = new_n5745_ & new_n6782_;
  assign new_n6784_ = new_n2896_ & new_n6777_;
  assign new_n6785_ = new_n5745_ & new_n6784_;
  assign new_n6786_ = ~new_n6783_ & ~new_n6785_;
  assign new_n6787_ = new_n2920_ & new_n6777_;
  assign new_n6788_ = new_n5745_ & new_n6787_;
  assign new_n6789_ = new_n5401_ & new_n5578_;
  assign new_n6790_ = ~new_n6788_ & ~new_n6789_;
  assign new_n6791_ = new_n6786_ & new_n6790_;
  assign new_n6792_ = new_n6781_ & new_n6791_;
  assign new_n6793_ = new_n5401_ & new_n5580_;
  assign new_n6794_ = new_n5401_ & new_n5576_;
  assign new_n6795_ = ~new_n6793_ & ~new_n6794_;
  assign new_n6796_ = new_n5401_ & new_n5587_;
  assign new_n6797_ = new_n5401_ & new_n5590_;
  assign new_n6798_ = ~new_n6796_ & ~new_n6797_;
  assign new_n6799_ = new_n6795_ & new_n6798_;
  assign new_n6800_ = new_n5403_ & new_n5600_;
  assign new_n6801_ = new_n5401_ & new_n5594_;
  assign new_n6802_ = new_n5403_ & new_n5596_;
  assign new_n6803_ = ~new_n6801_ & ~new_n6802_;
  assign new_n6804_ = ~new_n6800_ & new_n6803_;
  assign new_n6805_ = new_n6799_ & new_n6804_;
  assign new_n6806_ = new_n6792_ & new_n6805_;
  assign new_n6807_ = new_n5403_ & new_n5602_;
  assign new_n6808_ = new_n5403_ & new_n5605_;
  assign new_n6809_ = ~new_n6807_ & ~new_n6808_;
  assign new_n6810_ = new_n5403_ & new_n5608_;
  assign new_n6811_ = new_n5403_ & new_n5614_;
  assign new_n6812_ = ~new_n6810_ & ~new_n6811_;
  assign new_n6813_ = new_n6809_ & new_n6812_;
  assign new_n6814_ = new_n5437_ & new_n5755_;
  assign new_n6815_ = new_n2285_ & new_n5746_;
  assign new_n6816_ = new_n5745_ & new_n6815_;
  assign new_n6817_ = new_n2285_ & new_n5751_;
  assign new_n6818_ = new_n5745_ & new_n6817_;
  assign new_n6819_ = ~new_n6816_ & ~new_n6818_;
  assign new_n6820_ = ~new_n6814_ & new_n6819_;
  assign new_n6821_ = new_n6813_ & new_n6820_;
  assign new_n6822_ = new_n5437_ & new_n5759_;
  assign new_n6823_ = new_n5437_ & new_n5762_;
  assign new_n6824_ = ~new_n6822_ & ~new_n6823_;
  assign new_n6825_ = new_n5437_ & new_n5768_;
  assign new_n6826_ = new_n5437_ & new_n5770_;
  assign new_n6827_ = ~new_n6825_ & ~new_n6826_;
  assign new_n6828_ = new_n6824_ & new_n6827_;
  assign new_n6829_ = new_n5437_ & new_n5781_;
  assign new_n6830_ = new_n5437_ & new_n5773_;
  assign new_n6831_ = new_n5437_ & new_n5775_;
  assign new_n6832_ = ~new_n6830_ & ~new_n6831_;
  assign new_n6833_ = ~new_n6829_ & new_n6832_;
  assign new_n6834_ = new_n6828_ & new_n6833_;
  assign new_n6835_ = new_n6821_ & new_n6834_;
  assign new_n6836_ = new_n6806_ & new_n6835_;
  assign new_n6837_ = new_n5437_ & new_n5783_;
  assign new_n6838_ = new_n5437_ & new_n5779_;
  assign new_n6839_ = ~new_n6837_ & ~new_n6838_;
  assign new_n6840_ = new_n5437_ & new_n5789_;
  assign new_n6841_ = new_n5437_ & new_n5791_;
  assign new_n6842_ = ~new_n6840_ & ~new_n6841_;
  assign new_n6843_ = new_n6839_ & new_n6842_;
  assign new_n6844_ = new_n5437_ & new_n5794_;
  assign new_n6845_ = new_n5437_ & new_n5796_;
  assign new_n6846_ = ~new_n6844_ & ~new_n6845_;
  assign new_n6847_ = new_n5437_ & new_n5801_;
  assign new_n6848_ = new_n5437_ & new_n5803_;
  assign new_n6849_ = ~new_n6847_ & ~new_n6848_;
  assign new_n6850_ = new_n6846_ & new_n6849_;
  assign new_n6851_ = new_n6843_ & new_n6850_;
  assign new_n6852_ = new_n5463_ & new_n5755_;
  assign new_n6853_ = new_n5463_ & new_n5759_;
  assign new_n6854_ = ~new_n6852_ & ~new_n6853_;
  assign new_n6855_ = new_n5463_ & new_n5762_;
  assign new_n6856_ = new_n5463_ & new_n5768_;
  assign new_n6857_ = ~new_n6855_ & ~new_n6856_;
  assign new_n6858_ = new_n6854_ & new_n6857_;
  assign new_n6859_ = new_n5463_ & new_n5775_;
  assign new_n6860_ = new_n5463_ & new_n5770_;
  assign new_n6861_ = new_n5463_ & new_n5773_;
  assign new_n6862_ = ~new_n6860_ & ~new_n6861_;
  assign new_n6863_ = ~new_n6859_ & new_n6862_;
  assign new_n6864_ = new_n6858_ & new_n6863_;
  assign new_n6865_ = new_n6851_ & new_n6864_;
  assign new_n6866_ = new_n5463_ & new_n5781_;
  assign new_n6867_ = new_n5463_ & new_n5783_;
  assign new_n6868_ = ~new_n6866_ & ~new_n6867_;
  assign new_n6869_ = new_n5463_ & new_n5779_;
  assign new_n6870_ = new_n5463_ & new_n5789_;
  assign new_n6871_ = ~new_n6869_ & ~new_n6870_;
  assign new_n6872_ = new_n6868_ & new_n6871_;
  assign new_n6873_ = new_n5463_ & new_n5796_;
  assign new_n6874_ = new_n5463_ & new_n5791_;
  assign new_n6875_ = new_n5463_ & new_n5794_;
  assign new_n6876_ = ~new_n6874_ & ~new_n6875_;
  assign new_n6877_ = ~new_n6873_ & new_n6876_;
  assign new_n6878_ = new_n6872_ & new_n6877_;
  assign new_n6879_ = new_n5463_ & new_n5801_;
  assign new_n6880_ = new_n5463_ & new_n5803_;
  assign new_n6881_ = ~new_n6879_ & ~new_n6880_;
  assign new_n6882_ = new_n5522_ & new_n5755_;
  assign new_n6883_ = new_n5522_ & new_n5759_;
  assign new_n6884_ = ~new_n6882_ & ~new_n6883_;
  assign new_n6885_ = new_n6881_ & new_n6884_;
  assign new_n6886_ = new_n5522_ & new_n5770_;
  assign new_n6887_ = new_n5522_ & new_n5762_;
  assign new_n6888_ = new_n5522_ & new_n5768_;
  assign new_n6889_ = ~new_n6887_ & ~new_n6888_;
  assign new_n6890_ = ~new_n6886_ & new_n6889_;
  assign new_n6891_ = new_n6885_ & new_n6890_;
  assign new_n6892_ = new_n6878_ & new_n6891_;
  assign new_n6893_ = new_n6865_ & new_n6892_;
  assign new_n6894_ = new_n6836_ & new_n6893_;
  assign new_n6895_ = new_n6770_ & new_n6894_;
  assign new_n6896_ = new_n6655_ & new_n6895_;
  assign new_n6897_ = new_n5522_ & new_n5773_;
  assign new_n6898_ = new_n5522_ & new_n5775_;
  assign new_n6899_ = ~new_n6897_ & ~new_n6898_;
  assign new_n6900_ = new_n5522_ & new_n5781_;
  assign new_n6901_ = new_n5522_ & new_n5783_;
  assign new_n6902_ = ~new_n6900_ & ~new_n6901_;
  assign new_n6903_ = new_n6899_ & new_n6902_;
  assign new_n6904_ = new_n5522_ & new_n5779_;
  assign new_n6905_ = new_n5522_ & new_n5789_;
  assign new_n6906_ = ~new_n6904_ & ~new_n6905_;
  assign new_n6907_ = new_n5522_ & new_n5791_;
  assign new_n6908_ = new_n5522_ & new_n5794_;
  assign new_n6909_ = ~new_n6907_ & ~new_n6908_;
  assign new_n6910_ = new_n6906_ & new_n6909_;
  assign new_n6911_ = new_n6903_ & new_n6910_;
  assign new_n6912_ = new_n5522_ & new_n5796_;
  assign new_n6913_ = new_n5522_ & new_n5801_;
  assign new_n6914_ = ~new_n6912_ & ~new_n6913_;
  assign new_n6915_ = new_n5522_ & new_n5803_;
  assign new_n6916_ = new_n5545_ & new_n5755_;
  assign new_n6917_ = ~new_n6915_ & ~new_n6916_;
  assign new_n6918_ = new_n6914_ & new_n6917_;
  assign new_n6919_ = new_n5545_ & new_n5768_;
  assign new_n6920_ = new_n5545_ & new_n5759_;
  assign new_n6921_ = new_n5545_ & new_n5762_;
  assign new_n6922_ = ~new_n6920_ & ~new_n6921_;
  assign new_n6923_ = ~new_n6919_ & new_n6922_;
  assign new_n6924_ = new_n6918_ & new_n6923_;
  assign new_n6925_ = new_n6911_ & new_n6924_;
  assign new_n6926_ = new_n5545_ & new_n5770_;
  assign new_n6927_ = new_n5545_ & new_n5773_;
  assign new_n6928_ = ~new_n6926_ & ~new_n6927_;
  assign new_n6929_ = new_n5545_ & new_n5775_;
  assign new_n6930_ = new_n5545_ & new_n5781_;
  assign new_n6931_ = ~new_n6929_ & ~new_n6930_;
  assign new_n6932_ = new_n6928_ & new_n6931_;
  assign new_n6933_ = new_n5545_ & new_n5789_;
  assign new_n6934_ = new_n5545_ & new_n5783_;
  assign new_n6935_ = new_n5545_ & new_n5779_;
  assign new_n6936_ = ~new_n6934_ & ~new_n6935_;
  assign new_n6937_ = ~new_n6933_ & new_n6936_;
  assign new_n6938_ = new_n6932_ & new_n6937_;
  assign new_n6939_ = new_n5545_ & new_n5791_;
  assign new_n6940_ = new_n5545_ & new_n5794_;
  assign new_n6941_ = ~new_n6939_ & ~new_n6940_;
  assign new_n6942_ = new_n5545_ & new_n5796_;
  assign new_n6943_ = new_n5545_ & new_n5801_;
  assign new_n6944_ = ~new_n6942_ & ~new_n6943_;
  assign new_n6945_ = new_n6941_ & new_n6944_;
  assign new_n6946_ = new_n2270_ & new_n5909_;
  assign new_n6947_ = new_n5745_ & new_n6946_;
  assign new_n6948_ = new_n5545_ & new_n5803_;
  assign new_n6949_ = new_n2270_ & new_n5900_;
  assign new_n6950_ = new_n5745_ & new_n6949_;
  assign new_n6951_ = ~new_n6948_ & ~new_n6950_;
  assign new_n6952_ = ~new_n6947_ & new_n6951_;
  assign new_n6953_ = new_n6945_ & new_n6952_;
  assign new_n6954_ = new_n6938_ & new_n6953_;
  assign new_n6955_ = new_n6925_ & new_n6954_;
  assign new_n6956_ = A167 & new_n3016_;
  assign new_n6957_ = new_n2839_ & new_n6956_;
  assign new_n6958_ = new_n5745_ & new_n6957_;
  assign new_n6959_ = new_n2871_ & new_n6956_;
  assign new_n6960_ = new_n5745_ & new_n6959_;
  assign new_n6961_ = ~new_n6958_ & ~new_n6960_;
  assign new_n6962_ = new_n2896_ & new_n6956_;
  assign new_n6963_ = new_n5745_ & new_n6962_;
  assign new_n6964_ = new_n2920_ & new_n6956_;
  assign new_n6965_ = new_n5745_ & new_n6964_;
  assign new_n6966_ = ~new_n6963_ & ~new_n6965_;
  assign new_n6967_ = new_n6961_ & new_n6966_;
  assign new_n6968_ = new_n5570_ & new_n5578_;
  assign new_n6969_ = new_n5570_ & new_n5580_;
  assign new_n6970_ = ~new_n6968_ & ~new_n6969_;
  assign new_n6971_ = new_n5570_ & new_n5576_;
  assign new_n6972_ = new_n5570_ & new_n5587_;
  assign new_n6973_ = ~new_n6971_ & ~new_n6972_;
  assign new_n6974_ = new_n6970_ & new_n6973_;
  assign new_n6975_ = new_n6967_ & new_n6974_;
  assign new_n6976_ = new_n5570_ & new_n5590_;
  assign new_n6977_ = new_n5570_ & new_n5594_;
  assign new_n6978_ = ~new_n6976_ & ~new_n6977_;
  assign new_n6979_ = new_n5572_ & new_n5596_;
  assign new_n6980_ = new_n5572_ & new_n5600_;
  assign new_n6981_ = ~new_n6979_ & ~new_n6980_;
  assign new_n6982_ = new_n6978_ & new_n6981_;
  assign new_n6983_ = new_n5572_ & new_n5608_;
  assign new_n6984_ = new_n5572_ & new_n5602_;
  assign new_n6985_ = new_n5572_ & new_n5605_;
  assign new_n6986_ = ~new_n6984_ & ~new_n6985_;
  assign new_n6987_ = ~new_n6983_ & new_n6986_;
  assign new_n6988_ = new_n6982_ & new_n6987_;
  assign new_n6989_ = new_n6975_ & new_n6988_;
  assign new_n6990_ = new_n5572_ & new_n5614_;
  assign new_n6991_ = A168 & new_n1036_;
  assign new_n6992_ = new_n40_ & new_n6991_;
  assign new_n6993_ = new_n5690_ & new_n6992_;
  assign new_n6994_ = ~new_n6990_ & ~new_n6993_;
  assign new_n6995_ = new_n5694_ & new_n6992_;
  assign new_n6996_ = new_n5697_ & new_n6992_;
  assign new_n6997_ = ~new_n6995_ & ~new_n6996_;
  assign new_n6998_ = new_n6994_ & new_n6997_;
  assign new_n6999_ = new_n5702_ & new_n6992_;
  assign new_n7000_ = new_n5705_ & new_n6992_;
  assign new_n7001_ = new_n5708_ & new_n6992_;
  assign new_n7002_ = ~new_n7000_ & ~new_n7001_;
  assign new_n7003_ = ~new_n6999_ & new_n7002_;
  assign new_n7004_ = new_n6998_ & new_n7003_;
  assign new_n7005_ = new_n5714_ & new_n6992_;
  assign new_n7006_ = new_n5717_ & new_n6992_;
  assign new_n7007_ = ~new_n7005_ & ~new_n7006_;
  assign new_n7008_ = new_n5720_ & new_n6992_;
  assign new_n7009_ = new_n5722_ & new_n6992_;
  assign new_n7010_ = ~new_n7008_ & ~new_n7009_;
  assign new_n7011_ = new_n7007_ & new_n7010_;
  assign new_n7012_ = new_n5726_ & new_n6992_;
  assign new_n7013_ = new_n5728_ & new_n6992_;
  assign new_n7014_ = new_n5730_ & new_n6992_;
  assign new_n7015_ = ~new_n7013_ & ~new_n7014_;
  assign new_n7016_ = ~new_n7012_ & new_n7015_;
  assign new_n7017_ = new_n7011_ & new_n7016_;
  assign new_n7018_ = new_n7004_ & new_n7017_;
  assign new_n7019_ = new_n6989_ & new_n7018_;
  assign new_n7020_ = new_n6955_ & new_n7019_;
  assign new_n7021_ = new_n5737_ & new_n6992_;
  assign new_n7022_ = new_n5739_ & new_n6992_;
  assign new_n7023_ = ~new_n7021_ & ~new_n7022_;
  assign new_n7024_ = new_n5742_ & new_n6992_;
  assign new_n7025_ = A168 & new_n1213_;
  assign new_n7026_ = new_n40_ & new_n7025_;
  assign new_n7027_ = new_n5690_ & new_n7026_;
  assign new_n7028_ = ~new_n7024_ & ~new_n7027_;
  assign new_n7029_ = new_n7023_ & new_n7028_;
  assign new_n7030_ = new_n5694_ & new_n7026_;
  assign new_n7031_ = new_n5697_ & new_n7026_;
  assign new_n7032_ = ~new_n7030_ & ~new_n7031_;
  assign new_n7033_ = new_n5705_ & new_n7026_;
  assign new_n7034_ = new_n5708_ & new_n7026_;
  assign new_n7035_ = ~new_n7033_ & ~new_n7034_;
  assign new_n7036_ = new_n7032_ & new_n7035_;
  assign new_n7037_ = new_n7029_ & new_n7036_;
  assign new_n7038_ = new_n5702_ & new_n7026_;
  assign new_n7039_ = new_n5714_ & new_n7026_;
  assign new_n7040_ = ~new_n7038_ & ~new_n7039_;
  assign new_n7041_ = new_n5717_ & new_n7026_;
  assign new_n7042_ = new_n5720_ & new_n7026_;
  assign new_n7043_ = ~new_n7041_ & ~new_n7042_;
  assign new_n7044_ = new_n7040_ & new_n7043_;
  assign new_n7045_ = new_n5730_ & new_n7026_;
  assign new_n7046_ = new_n5722_ & new_n7026_;
  assign new_n7047_ = new_n5728_ & new_n7026_;
  assign new_n7048_ = ~new_n7046_ & ~new_n7047_;
  assign new_n7049_ = ~new_n7045_ & new_n7048_;
  assign new_n7050_ = new_n7044_ & new_n7049_;
  assign new_n7051_ = new_n7037_ & new_n7050_;
  assign new_n7052_ = new_n5726_ & new_n7026_;
  assign new_n7053_ = new_n5737_ & new_n7026_;
  assign new_n7054_ = ~new_n7052_ & ~new_n7053_;
  assign new_n7055_ = new_n5739_ & new_n7026_;
  assign new_n7056_ = new_n5742_ & new_n7026_;
  assign new_n7057_ = ~new_n7055_ & ~new_n7056_;
  assign new_n7058_ = new_n7054_ & new_n7057_;
  assign new_n7059_ = A168 & new_n1219_;
  assign new_n7060_ = new_n40_ & new_n7059_;
  assign new_n7061_ = new_n5697_ & new_n7060_;
  assign new_n7062_ = new_n5690_ & new_n7060_;
  assign new_n7063_ = new_n5694_ & new_n7060_;
  assign new_n7064_ = ~new_n7062_ & ~new_n7063_;
  assign new_n7065_ = ~new_n7061_ & new_n7064_;
  assign new_n7066_ = new_n7058_ & new_n7065_;
  assign new_n7067_ = new_n5705_ & new_n7060_;
  assign new_n7068_ = new_n5708_ & new_n7060_;
  assign new_n7069_ = ~new_n7067_ & ~new_n7068_;
  assign new_n7070_ = new_n5702_ & new_n7060_;
  assign new_n7071_ = new_n5714_ & new_n7060_;
  assign new_n7072_ = ~new_n7070_ & ~new_n7071_;
  assign new_n7073_ = new_n7069_ & new_n7072_;
  assign new_n7074_ = new_n5722_ & new_n7060_;
  assign new_n7075_ = new_n5717_ & new_n7060_;
  assign new_n7076_ = new_n5720_ & new_n7060_;
  assign new_n7077_ = ~new_n7075_ & ~new_n7076_;
  assign new_n7078_ = ~new_n7074_ & new_n7077_;
  assign new_n7079_ = new_n7073_ & new_n7078_;
  assign new_n7080_ = new_n7066_ & new_n7079_;
  assign new_n7081_ = new_n7051_ & new_n7080_;
  assign new_n7082_ = new_n5728_ & new_n7060_;
  assign new_n7083_ = new_n5730_ & new_n7060_;
  assign new_n7084_ = ~new_n7082_ & ~new_n7083_;
  assign new_n7085_ = new_n5726_ & new_n7060_;
  assign new_n7086_ = new_n5737_ & new_n7060_;
  assign new_n7087_ = ~new_n7085_ & ~new_n7086_;
  assign new_n7088_ = new_n7084_ & new_n7087_;
  assign new_n7089_ = new_n5739_ & new_n7060_;
  assign new_n7090_ = new_n5742_ & new_n7060_;
  assign new_n7091_ = ~new_n7089_ & ~new_n7090_;
  assign new_n7092_ = A168 & new_n1225_;
  assign new_n7093_ = new_n40_ & new_n7092_;
  assign new_n7094_ = new_n5690_ & new_n7093_;
  assign new_n7095_ = new_n5694_ & new_n7093_;
  assign new_n7096_ = ~new_n7094_ & ~new_n7095_;
  assign new_n7097_ = new_n7091_ & new_n7096_;
  assign new_n7098_ = new_n7088_ & new_n7097_;
  assign new_n7099_ = new_n5697_ & new_n7093_;
  assign new_n7100_ = new_n5705_ & new_n7093_;
  assign new_n7101_ = ~new_n7099_ & ~new_n7100_;
  assign new_n7102_ = new_n5708_ & new_n7093_;
  assign new_n7103_ = new_n5702_ & new_n7093_;
  assign new_n7104_ = ~new_n7102_ & ~new_n7103_;
  assign new_n7105_ = new_n7101_ & new_n7104_;
  assign new_n7106_ = new_n5720_ & new_n7093_;
  assign new_n7107_ = new_n5714_ & new_n7093_;
  assign new_n7108_ = new_n5717_ & new_n7093_;
  assign new_n7109_ = ~new_n7107_ & ~new_n7108_;
  assign new_n7110_ = ~new_n7106_ & new_n7109_;
  assign new_n7111_ = new_n7105_ & new_n7110_;
  assign new_n7112_ = new_n7098_ & new_n7111_;
  assign new_n7113_ = new_n5722_ & new_n7093_;
  assign new_n7114_ = new_n5728_ & new_n7093_;
  assign new_n7115_ = ~new_n7113_ & ~new_n7114_;
  assign new_n7116_ = new_n5730_ & new_n7093_;
  assign new_n7117_ = new_n5726_ & new_n7093_;
  assign new_n7118_ = ~new_n7116_ & ~new_n7117_;
  assign new_n7119_ = new_n7115_ & new_n7118_;
  assign new_n7120_ = new_n5742_ & new_n7093_;
  assign new_n7121_ = new_n5737_ & new_n7093_;
  assign new_n7122_ = new_n5739_ & new_n7093_;
  assign new_n7123_ = ~new_n7121_ & ~new_n7122_;
  assign new_n7124_ = ~new_n7120_ & new_n7123_;
  assign new_n7125_ = new_n7119_ & new_n7124_;
  assign new_n7126_ = ~A168 & A169;
  assign new_n7127_ = new_n4124_ & new_n7126_;
  assign new_n7128_ = new_n5578_ & new_n7127_;
  assign new_n7129_ = new_n5580_ & new_n7127_;
  assign new_n7130_ = ~new_n7128_ & ~new_n7129_;
  assign new_n7131_ = new_n5576_ & new_n7127_;
  assign new_n7132_ = new_n5587_ & new_n7127_;
  assign new_n7133_ = ~new_n7131_ & ~new_n7132_;
  assign new_n7134_ = new_n7130_ & new_n7133_;
  assign new_n7135_ = new_n4129_ & new_n7126_;
  assign new_n7136_ = new_n5596_ & new_n7135_;
  assign new_n7137_ = new_n5590_ & new_n7127_;
  assign new_n7138_ = new_n5594_ & new_n7127_;
  assign new_n7139_ = ~new_n7137_ & ~new_n7138_;
  assign new_n7140_ = ~new_n7136_ & new_n7139_;
  assign new_n7141_ = new_n7134_ & new_n7140_;
  assign new_n7142_ = new_n7125_ & new_n7141_;
  assign new_n7143_ = new_n7112_ & new_n7142_;
  assign new_n7144_ = new_n7081_ & new_n7143_;
  assign new_n7145_ = new_n7020_ & new_n7144_;
  assign new_n7146_ = new_n5600_ & new_n7135_;
  assign new_n7147_ = new_n5602_ & new_n7135_;
  assign new_n7148_ = ~new_n7146_ & ~new_n7147_;
  assign new_n7149_ = new_n5605_ & new_n7135_;
  assign new_n7150_ = new_n5608_ & new_n7135_;
  assign new_n7151_ = ~new_n7149_ & ~new_n7150_;
  assign new_n7152_ = new_n7148_ & new_n7151_;
  assign new_n7153_ = new_n5614_ & new_n7135_;
  assign new_n7154_ = new_n4268_ & new_n7126_;
  assign new_n7155_ = new_n5578_ & new_n7154_;
  assign new_n7156_ = ~new_n7153_ & ~new_n7155_;
  assign new_n7157_ = new_n5580_ & new_n7154_;
  assign new_n7158_ = new_n5576_ & new_n7154_;
  assign new_n7159_ = ~new_n7157_ & ~new_n7158_;
  assign new_n7160_ = new_n7156_ & new_n7159_;
  assign new_n7161_ = new_n7152_ & new_n7160_;
  assign new_n7162_ = new_n5587_ & new_n7154_;
  assign new_n7163_ = new_n5590_ & new_n7154_;
  assign new_n7164_ = ~new_n7162_ & ~new_n7163_;
  assign new_n7165_ = new_n5594_ & new_n7154_;
  assign new_n7166_ = new_n4272_ & new_n7126_;
  assign new_n7167_ = new_n5596_ & new_n7166_;
  assign new_n7168_ = ~new_n7165_ & ~new_n7167_;
  assign new_n7169_ = new_n7164_ & new_n7168_;
  assign new_n7170_ = new_n5605_ & new_n7166_;
  assign new_n7171_ = new_n5600_ & new_n7166_;
  assign new_n7172_ = new_n5602_ & new_n7166_;
  assign new_n7173_ = ~new_n7171_ & ~new_n7172_;
  assign new_n7174_ = ~new_n7170_ & new_n7173_;
  assign new_n7175_ = new_n7169_ & new_n7174_;
  assign new_n7176_ = new_n7161_ & new_n7175_;
  assign new_n7177_ = new_n5608_ & new_n7166_;
  assign new_n7178_ = new_n5614_ & new_n7166_;
  assign new_n7179_ = ~new_n7177_ & ~new_n7178_;
  assign new_n7180_ = new_n4277_ & new_n7126_;
  assign new_n7181_ = new_n5578_ & new_n7180_;
  assign new_n7182_ = new_n5580_ & new_n7180_;
  assign new_n7183_ = ~new_n7181_ & ~new_n7182_;
  assign new_n7184_ = new_n7179_ & new_n7183_;
  assign new_n7185_ = new_n5590_ & new_n7180_;
  assign new_n7186_ = new_n5576_ & new_n7180_;
  assign new_n7187_ = new_n5587_ & new_n7180_;
  assign new_n7188_ = ~new_n7186_ & ~new_n7187_;
  assign new_n7189_ = ~new_n7185_ & new_n7188_;
  assign new_n7190_ = new_n7184_ & new_n7189_;
  assign new_n7191_ = new_n5594_ & new_n7180_;
  assign new_n7192_ = new_n4280_ & new_n7126_;
  assign new_n7193_ = new_n5596_ & new_n7192_;
  assign new_n7194_ = ~new_n7191_ & ~new_n7193_;
  assign new_n7195_ = new_n5600_ & new_n7192_;
  assign new_n7196_ = new_n5602_ & new_n7192_;
  assign new_n7197_ = ~new_n7195_ & ~new_n7196_;
  assign new_n7198_ = new_n7194_ & new_n7197_;
  assign new_n7199_ = new_n5614_ & new_n7192_;
  assign new_n7200_ = new_n5605_ & new_n7192_;
  assign new_n7201_ = new_n5608_ & new_n7192_;
  assign new_n7202_ = ~new_n7200_ & ~new_n7201_;
  assign new_n7203_ = ~new_n7199_ & new_n7202_;
  assign new_n7204_ = new_n7198_ & new_n7203_;
  assign new_n7205_ = new_n7190_ & new_n7204_;
  assign new_n7206_ = new_n7176_ & new_n7205_;
  assign new_n7207_ = new_n4284_ & new_n7126_;
  assign new_n7208_ = new_n5578_ & new_n7207_;
  assign new_n7209_ = new_n5580_ & new_n7207_;
  assign new_n7210_ = ~new_n7208_ & ~new_n7209_;
  assign new_n7211_ = new_n5576_ & new_n7207_;
  assign new_n7212_ = new_n5587_ & new_n7207_;
  assign new_n7213_ = ~new_n7211_ & ~new_n7212_;
  assign new_n7214_ = new_n7210_ & new_n7213_;
  assign new_n7215_ = new_n5590_ & new_n7207_;
  assign new_n7216_ = new_n5594_ & new_n7207_;
  assign new_n7217_ = ~new_n7215_ & ~new_n7216_;
  assign new_n7218_ = new_n4287_ & new_n7126_;
  assign new_n7219_ = new_n5596_ & new_n7218_;
  assign new_n7220_ = new_n5600_ & new_n7218_;
  assign new_n7221_ = ~new_n7219_ & ~new_n7220_;
  assign new_n7222_ = new_n7217_ & new_n7221_;
  assign new_n7223_ = new_n7214_ & new_n7222_;
  assign new_n7224_ = new_n5602_ & new_n7218_;
  assign new_n7225_ = new_n5605_ & new_n7218_;
  assign new_n7226_ = ~new_n7224_ & ~new_n7225_;
  assign new_n7227_ = new_n5608_ & new_n7218_;
  assign new_n7228_ = new_n5614_ & new_n7218_;
  assign new_n7229_ = ~new_n7227_ & ~new_n7228_;
  assign new_n7230_ = new_n7226_ & new_n7229_;
  assign new_n7231_ = new_n4295_ & new_n7126_;
  assign new_n7232_ = new_n5697_ & new_n7231_;
  assign new_n7233_ = new_n5690_ & new_n7231_;
  assign new_n7234_ = new_n5694_ & new_n7231_;
  assign new_n7235_ = ~new_n7233_ & ~new_n7234_;
  assign new_n7236_ = ~new_n7232_ & new_n7235_;
  assign new_n7237_ = new_n7230_ & new_n7236_;
  assign new_n7238_ = new_n7223_ & new_n7237_;
  assign new_n7239_ = new_n5705_ & new_n7231_;
  assign new_n7240_ = new_n5708_ & new_n7231_;
  assign new_n7241_ = ~new_n7239_ & ~new_n7240_;
  assign new_n7242_ = new_n5702_ & new_n7231_;
  assign new_n7243_ = new_n5714_ & new_n7231_;
  assign new_n7244_ = ~new_n7242_ & ~new_n7243_;
  assign new_n7245_ = new_n7241_ & new_n7244_;
  assign new_n7246_ = new_n5722_ & new_n7231_;
  assign new_n7247_ = new_n5717_ & new_n7231_;
  assign new_n7248_ = new_n5720_ & new_n7231_;
  assign new_n7249_ = ~new_n7247_ & ~new_n7248_;
  assign new_n7250_ = ~new_n7246_ & new_n7249_;
  assign new_n7251_ = new_n7245_ & new_n7250_;
  assign new_n7252_ = new_n5728_ & new_n7231_;
  assign new_n7253_ = new_n5730_ & new_n7231_;
  assign new_n7254_ = ~new_n7252_ & ~new_n7253_;
  assign new_n7255_ = new_n5726_ & new_n7231_;
  assign new_n7256_ = new_n5737_ & new_n7231_;
  assign new_n7257_ = ~new_n7255_ & ~new_n7256_;
  assign new_n7258_ = new_n7254_ & new_n7257_;
  assign new_n7259_ = ~A168 & ~A170;
  assign new_n7260_ = new_n4124_ & new_n7259_;
  assign new_n7261_ = new_n5578_ & new_n7260_;
  assign new_n7262_ = new_n5739_ & new_n7231_;
  assign new_n7263_ = new_n5742_ & new_n7231_;
  assign new_n7264_ = ~new_n7262_ & ~new_n7263_;
  assign new_n7265_ = ~new_n7261_ & new_n7264_;
  assign new_n7266_ = new_n7258_ & new_n7265_;
  assign new_n7267_ = new_n7251_ & new_n7266_;
  assign new_n7268_ = new_n7238_ & new_n7267_;
  assign new_n7269_ = new_n7206_ & new_n7268_;
  assign new_n7270_ = new_n5580_ & new_n7260_;
  assign new_n7271_ = new_n5576_ & new_n7260_;
  assign new_n7272_ = ~new_n7270_ & ~new_n7271_;
  assign new_n7273_ = new_n5587_ & new_n7260_;
  assign new_n7274_ = new_n5590_ & new_n7260_;
  assign new_n7275_ = ~new_n7273_ & ~new_n7274_;
  assign new_n7276_ = new_n7272_ & new_n7275_;
  assign new_n7277_ = new_n5594_ & new_n7260_;
  assign new_n7278_ = new_n4129_ & new_n7259_;
  assign new_n7279_ = new_n5596_ & new_n7278_;
  assign new_n7280_ = ~new_n7277_ & ~new_n7279_;
  assign new_n7281_ = new_n5600_ & new_n7278_;
  assign new_n7282_ = new_n5602_ & new_n7278_;
  assign new_n7283_ = ~new_n7281_ & ~new_n7282_;
  assign new_n7284_ = new_n7280_ & new_n7283_;
  assign new_n7285_ = new_n7276_ & new_n7284_;
  assign new_n7286_ = new_n5605_ & new_n7278_;
  assign new_n7287_ = new_n5608_ & new_n7278_;
  assign new_n7288_ = ~new_n7286_ & ~new_n7287_;
  assign new_n7289_ = new_n5614_ & new_n7278_;
  assign new_n7290_ = new_n4268_ & new_n7259_;
  assign new_n7291_ = new_n5578_ & new_n7290_;
  assign new_n7292_ = ~new_n7289_ & ~new_n7291_;
  assign new_n7293_ = new_n7288_ & new_n7292_;
  assign new_n7294_ = new_n5587_ & new_n7290_;
  assign new_n7295_ = new_n5580_ & new_n7290_;
  assign new_n7296_ = new_n5576_ & new_n7290_;
  assign new_n7297_ = ~new_n7295_ & ~new_n7296_;
  assign new_n7298_ = ~new_n7294_ & new_n7297_;
  assign new_n7299_ = new_n7293_ & new_n7298_;
  assign new_n7300_ = new_n7285_ & new_n7299_;
  assign new_n7301_ = new_n5590_ & new_n7290_;
  assign new_n7302_ = new_n5594_ & new_n7290_;
  assign new_n7303_ = ~new_n7301_ & ~new_n7302_;
  assign new_n7304_ = new_n4272_ & new_n7259_;
  assign new_n7305_ = new_n5596_ & new_n7304_;
  assign new_n7306_ = new_n5600_ & new_n7304_;
  assign new_n7307_ = ~new_n7305_ & ~new_n7306_;
  assign new_n7308_ = new_n7303_ & new_n7307_;
  assign new_n7309_ = new_n5608_ & new_n7304_;
  assign new_n7310_ = new_n5602_ & new_n7304_;
  assign new_n7311_ = new_n5605_ & new_n7304_;
  assign new_n7312_ = ~new_n7310_ & ~new_n7311_;
  assign new_n7313_ = ~new_n7309_ & new_n7312_;
  assign new_n7314_ = new_n7308_ & new_n7313_;
  assign new_n7315_ = new_n5614_ & new_n7304_;
  assign new_n7316_ = new_n4277_ & new_n7259_;
  assign new_n7317_ = new_n5578_ & new_n7316_;
  assign new_n7318_ = ~new_n7315_ & ~new_n7317_;
  assign new_n7319_ = new_n5580_ & new_n7316_;
  assign new_n7320_ = new_n5576_ & new_n7316_;
  assign new_n7321_ = ~new_n7319_ & ~new_n7320_;
  assign new_n7322_ = new_n7318_ & new_n7321_;
  assign new_n7323_ = new_n5594_ & new_n7316_;
  assign new_n7324_ = new_n5587_ & new_n7316_;
  assign new_n7325_ = new_n5590_ & new_n7316_;
  assign new_n7326_ = ~new_n7324_ & ~new_n7325_;
  assign new_n7327_ = ~new_n7323_ & new_n7326_;
  assign new_n7328_ = new_n7322_ & new_n7327_;
  assign new_n7329_ = new_n7314_ & new_n7328_;
  assign new_n7330_ = new_n7300_ & new_n7329_;
  assign new_n7331_ = new_n4280_ & new_n7259_;
  assign new_n7332_ = new_n5596_ & new_n7331_;
  assign new_n7333_ = new_n5600_ & new_n7331_;
  assign new_n7334_ = ~new_n7332_ & ~new_n7333_;
  assign new_n7335_ = new_n5602_ & new_n7331_;
  assign new_n7336_ = new_n5605_ & new_n7331_;
  assign new_n7337_ = ~new_n7335_ & ~new_n7336_;
  assign new_n7338_ = new_n7334_ & new_n7337_;
  assign new_n7339_ = new_n4284_ & new_n7259_;
  assign new_n7340_ = new_n5578_ & new_n7339_;
  assign new_n7341_ = new_n5608_ & new_n7331_;
  assign new_n7342_ = new_n5614_ & new_n7331_;
  assign new_n7343_ = ~new_n7341_ & ~new_n7342_;
  assign new_n7344_ = ~new_n7340_ & new_n7343_;
  assign new_n7345_ = new_n7338_ & new_n7344_;
  assign new_n7346_ = new_n5580_ & new_n7339_;
  assign new_n7347_ = new_n5576_ & new_n7339_;
  assign new_n7348_ = ~new_n7346_ & ~new_n7347_;
  assign new_n7349_ = new_n5587_ & new_n7339_;
  assign new_n7350_ = new_n5590_ & new_n7339_;
  assign new_n7351_ = ~new_n7349_ & ~new_n7350_;
  assign new_n7352_ = new_n7348_ & new_n7351_;
  assign new_n7353_ = new_n4287_ & new_n7259_;
  assign new_n7354_ = new_n5600_ & new_n7353_;
  assign new_n7355_ = new_n5594_ & new_n7339_;
  assign new_n7356_ = new_n5596_ & new_n7353_;
  assign new_n7357_ = ~new_n7355_ & ~new_n7356_;
  assign new_n7358_ = ~new_n7354_ & new_n7357_;
  assign new_n7359_ = new_n7352_ & new_n7358_;
  assign new_n7360_ = new_n7345_ & new_n7359_;
  assign new_n7361_ = new_n5602_ & new_n7353_;
  assign new_n7362_ = new_n5605_ & new_n7353_;
  assign new_n7363_ = ~new_n7361_ & ~new_n7362_;
  assign new_n7364_ = new_n5608_ & new_n7353_;
  assign new_n7365_ = new_n5614_ & new_n7353_;
  assign new_n7366_ = ~new_n7364_ & ~new_n7365_;
  assign new_n7367_ = new_n7363_ & new_n7366_;
  assign new_n7368_ = new_n4295_ & new_n7259_;
  assign new_n7369_ = new_n5697_ & new_n7368_;
  assign new_n7370_ = new_n5690_ & new_n7368_;
  assign new_n7371_ = new_n5694_ & new_n7368_;
  assign new_n7372_ = ~new_n7370_ & ~new_n7371_;
  assign new_n7373_ = ~new_n7369_ & new_n7372_;
  assign new_n7374_ = new_n7367_ & new_n7373_;
  assign new_n7375_ = new_n5705_ & new_n7368_;
  assign new_n7376_ = new_n5708_ & new_n7368_;
  assign new_n7377_ = ~new_n7375_ & ~new_n7376_;
  assign new_n7378_ = new_n5702_ & new_n7368_;
  assign new_n7379_ = new_n5714_ & new_n7368_;
  assign new_n7380_ = ~new_n7378_ & ~new_n7379_;
  assign new_n7381_ = new_n7377_ & new_n7380_;
  assign new_n7382_ = new_n5722_ & new_n7368_;
  assign new_n7383_ = new_n5717_ & new_n7368_;
  assign new_n7384_ = new_n5720_ & new_n7368_;
  assign new_n7385_ = ~new_n7383_ & ~new_n7384_;
  assign new_n7386_ = ~new_n7382_ & new_n7385_;
  assign new_n7387_ = new_n7381_ & new_n7386_;
  assign new_n7388_ = new_n7374_ & new_n7387_;
  assign new_n7389_ = new_n7360_ & new_n7388_;
  assign new_n7390_ = new_n7330_ & new_n7389_;
  assign new_n7391_ = new_n7269_ & new_n7390_;
  assign new_n7392_ = new_n7145_ & new_n7391_;
  assign new_n7393_ = new_n6896_ & new_n7392_;
  assign new_n7394_ = new_n5728_ & new_n7368_;
  assign new_n7395_ = new_n5730_ & new_n7368_;
  assign new_n7396_ = ~new_n7394_ & ~new_n7395_;
  assign new_n7397_ = new_n5726_ & new_n7368_;
  assign new_n7398_ = new_n5737_ & new_n7368_;
  assign new_n7399_ = ~new_n7397_ & ~new_n7398_;
  assign new_n7400_ = new_n7396_ & new_n7399_;
  assign new_n7401_ = new_n5739_ & new_n7368_;
  assign new_n7402_ = new_n5742_ & new_n7368_;
  assign new_n7403_ = ~new_n7401_ & ~new_n7402_;
  assign new_n7404_ = ~A166 & ~A167;
  assign new_n7405_ = new_n4124_ & new_n7404_;
  assign new_n7406_ = new_n5578_ & new_n7405_;
  assign new_n7407_ = new_n5580_ & new_n7405_;
  assign new_n7408_ = ~new_n7406_ & ~new_n7407_;
  assign new_n7409_ = new_n7403_ & new_n7408_;
  assign new_n7410_ = new_n7400_ & new_n7409_;
  assign new_n7411_ = new_n5576_ & new_n7405_;
  assign new_n7412_ = new_n5587_ & new_n7405_;
  assign new_n7413_ = ~new_n7411_ & ~new_n7412_;
  assign new_n7414_ = new_n5590_ & new_n7405_;
  assign new_n7415_ = new_n5594_ & new_n7405_;
  assign new_n7416_ = ~new_n7414_ & ~new_n7415_;
  assign new_n7417_ = new_n7413_ & new_n7416_;
  assign new_n7418_ = new_n4129_ & new_n7404_;
  assign new_n7419_ = new_n5602_ & new_n7418_;
  assign new_n7420_ = new_n5596_ & new_n7418_;
  assign new_n7421_ = new_n5600_ & new_n7418_;
  assign new_n7422_ = ~new_n7420_ & ~new_n7421_;
  assign new_n7423_ = ~new_n7419_ & new_n7422_;
  assign new_n7424_ = new_n7417_ & new_n7423_;
  assign new_n7425_ = new_n7410_ & new_n7424_;
  assign new_n7426_ = new_n5605_ & new_n7418_;
  assign new_n7427_ = new_n5608_ & new_n7418_;
  assign new_n7428_ = ~new_n7426_ & ~new_n7427_;
  assign new_n7429_ = new_n5614_ & new_n7418_;
  assign new_n7430_ = new_n4268_ & new_n7404_;
  assign new_n7431_ = new_n5578_ & new_n7430_;
  assign new_n7432_ = ~new_n7429_ & ~new_n7431_;
  assign new_n7433_ = new_n7428_ & new_n7432_;
  assign new_n7434_ = new_n5587_ & new_n7430_;
  assign new_n7435_ = new_n5580_ & new_n7430_;
  assign new_n7436_ = new_n5576_ & new_n7430_;
  assign new_n7437_ = ~new_n7435_ & ~new_n7436_;
  assign new_n7438_ = ~new_n7434_ & new_n7437_;
  assign new_n7439_ = new_n7433_ & new_n7438_;
  assign new_n7440_ = new_n5590_ & new_n7430_;
  assign new_n7441_ = new_n5594_ & new_n7430_;
  assign new_n7442_ = ~new_n7440_ & ~new_n7441_;
  assign new_n7443_ = new_n4272_ & new_n7404_;
  assign new_n7444_ = new_n5596_ & new_n7443_;
  assign new_n7445_ = new_n5600_ & new_n7443_;
  assign new_n7446_ = ~new_n7444_ & ~new_n7445_;
  assign new_n7447_ = new_n7442_ & new_n7446_;
  assign new_n7448_ = new_n5608_ & new_n7443_;
  assign new_n7449_ = new_n5602_ & new_n7443_;
  assign new_n7450_ = new_n5605_ & new_n7443_;
  assign new_n7451_ = ~new_n7449_ & ~new_n7450_;
  assign new_n7452_ = ~new_n7448_ & new_n7451_;
  assign new_n7453_ = new_n7447_ & new_n7452_;
  assign new_n7454_ = new_n7439_ & new_n7453_;
  assign new_n7455_ = new_n7425_ & new_n7454_;
  assign new_n7456_ = new_n5614_ & new_n7443_;
  assign new_n7457_ = new_n4277_ & new_n7404_;
  assign new_n7458_ = new_n5578_ & new_n7457_;
  assign new_n7459_ = ~new_n7456_ & ~new_n7458_;
  assign new_n7460_ = new_n5580_ & new_n7457_;
  assign new_n7461_ = new_n5576_ & new_n7457_;
  assign new_n7462_ = ~new_n7460_ & ~new_n7461_;
  assign new_n7463_ = new_n7459_ & new_n7462_;
  assign new_n7464_ = new_n5587_ & new_n7457_;
  assign new_n7465_ = new_n5590_ & new_n7457_;
  assign new_n7466_ = ~new_n7464_ & ~new_n7465_;
  assign new_n7467_ = new_n5594_ & new_n7457_;
  assign new_n7468_ = new_n4280_ & new_n7404_;
  assign new_n7469_ = new_n5596_ & new_n7468_;
  assign new_n7470_ = ~new_n7467_ & ~new_n7469_;
  assign new_n7471_ = new_n7466_ & new_n7470_;
  assign new_n7472_ = new_n7463_ & new_n7471_;
  assign new_n7473_ = new_n5600_ & new_n7468_;
  assign new_n7474_ = new_n5602_ & new_n7468_;
  assign new_n7475_ = ~new_n7473_ & ~new_n7474_;
  assign new_n7476_ = new_n5605_ & new_n7468_;
  assign new_n7477_ = new_n5608_ & new_n7468_;
  assign new_n7478_ = ~new_n7476_ & ~new_n7477_;
  assign new_n7479_ = new_n7475_ & new_n7478_;
  assign new_n7480_ = new_n4284_ & new_n7404_;
  assign new_n7481_ = new_n5580_ & new_n7480_;
  assign new_n7482_ = new_n5614_ & new_n7468_;
  assign new_n7483_ = new_n5578_ & new_n7480_;
  assign new_n7484_ = ~new_n7482_ & ~new_n7483_;
  assign new_n7485_ = ~new_n7481_ & new_n7484_;
  assign new_n7486_ = new_n7479_ & new_n7485_;
  assign new_n7487_ = new_n7472_ & new_n7486_;
  assign new_n7488_ = new_n5576_ & new_n7480_;
  assign new_n7489_ = new_n5587_ & new_n7480_;
  assign new_n7490_ = ~new_n7488_ & ~new_n7489_;
  assign new_n7491_ = new_n5590_ & new_n7480_;
  assign new_n7492_ = new_n5594_ & new_n7480_;
  assign new_n7493_ = ~new_n7491_ & ~new_n7492_;
  assign new_n7494_ = new_n7490_ & new_n7493_;
  assign new_n7495_ = new_n4287_ & new_n7404_;
  assign new_n7496_ = new_n5602_ & new_n7495_;
  assign new_n7497_ = new_n5596_ & new_n7495_;
  assign new_n7498_ = new_n5600_ & new_n7495_;
  assign new_n7499_ = ~new_n7497_ & ~new_n7498_;
  assign new_n7500_ = ~new_n7496_ & new_n7499_;
  assign new_n7501_ = new_n7494_ & new_n7500_;
  assign new_n7502_ = new_n5605_ & new_n7495_;
  assign new_n7503_ = new_n5608_ & new_n7495_;
  assign new_n7504_ = ~new_n7502_ & ~new_n7503_;
  assign new_n7505_ = new_n5614_ & new_n7495_;
  assign new_n7506_ = new_n4295_ & new_n7404_;
  assign new_n7507_ = new_n5690_ & new_n7506_;
  assign new_n7508_ = ~new_n7505_ & ~new_n7507_;
  assign new_n7509_ = new_n7504_ & new_n7508_;
  assign new_n7510_ = new_n5705_ & new_n7506_;
  assign new_n7511_ = new_n5694_ & new_n7506_;
  assign new_n7512_ = new_n5697_ & new_n7506_;
  assign new_n7513_ = ~new_n7511_ & ~new_n7512_;
  assign new_n7514_ = ~new_n7510_ & new_n7513_;
  assign new_n7515_ = new_n7509_ & new_n7514_;
  assign new_n7516_ = new_n7501_ & new_n7515_;
  assign new_n7517_ = new_n7487_ & new_n7516_;
  assign new_n7518_ = new_n7455_ & new_n7517_;
  assign new_n7519_ = new_n5708_ & new_n7506_;
  assign new_n7520_ = new_n5702_ & new_n7506_;
  assign new_n7521_ = ~new_n7519_ & ~new_n7520_;
  assign new_n7522_ = new_n5714_ & new_n7506_;
  assign new_n7523_ = new_n5717_ & new_n7506_;
  assign new_n7524_ = ~new_n7522_ & ~new_n7523_;
  assign new_n7525_ = new_n7521_ & new_n7524_;
  assign new_n7526_ = new_n5720_ & new_n7506_;
  assign new_n7527_ = new_n5722_ & new_n7506_;
  assign new_n7528_ = ~new_n7526_ & ~new_n7527_;
  assign new_n7529_ = new_n5728_ & new_n7506_;
  assign new_n7530_ = new_n5730_ & new_n7506_;
  assign new_n7531_ = ~new_n7529_ & ~new_n7530_;
  assign new_n7532_ = new_n7528_ & new_n7531_;
  assign new_n7533_ = new_n7525_ & new_n7532_;
  assign new_n7534_ = new_n5726_ & new_n7506_;
  assign new_n7535_ = new_n5737_ & new_n7506_;
  assign new_n7536_ = ~new_n7534_ & ~new_n7535_;
  assign new_n7537_ = new_n5739_ & new_n7506_;
  assign new_n7538_ = new_n5742_ & new_n7506_;
  assign new_n7539_ = ~new_n7537_ & ~new_n7538_;
  assign new_n7540_ = new_n7536_ & new_n7539_;
  assign new_n7541_ = A166 & A167;
  assign new_n7542_ = new_n4124_ & new_n7541_;
  assign new_n7543_ = new_n5576_ & new_n7542_;
  assign new_n7544_ = new_n5578_ & new_n7542_;
  assign new_n7545_ = new_n5580_ & new_n7542_;
  assign new_n7546_ = ~new_n7544_ & ~new_n7545_;
  assign new_n7547_ = ~new_n7543_ & new_n7546_;
  assign new_n7548_ = new_n7540_ & new_n7547_;
  assign new_n7549_ = new_n7533_ & new_n7548_;
  assign new_n7550_ = new_n5587_ & new_n7542_;
  assign new_n7551_ = new_n5590_ & new_n7542_;
  assign new_n7552_ = ~new_n7550_ & ~new_n7551_;
  assign new_n7553_ = new_n5594_ & new_n7542_;
  assign new_n7554_ = new_n4129_ & new_n7541_;
  assign new_n7555_ = new_n5596_ & new_n7554_;
  assign new_n7556_ = ~new_n7553_ & ~new_n7555_;
  assign new_n7557_ = new_n7552_ & new_n7556_;
  assign new_n7558_ = new_n5605_ & new_n7554_;
  assign new_n7559_ = new_n5600_ & new_n7554_;
  assign new_n7560_ = new_n5602_ & new_n7554_;
  assign new_n7561_ = ~new_n7559_ & ~new_n7560_;
  assign new_n7562_ = ~new_n7558_ & new_n7561_;
  assign new_n7563_ = new_n7557_ & new_n7562_;
  assign new_n7564_ = new_n5608_ & new_n7554_;
  assign new_n7565_ = new_n5614_ & new_n7554_;
  assign new_n7566_ = ~new_n7564_ & ~new_n7565_;
  assign new_n7567_ = new_n4268_ & new_n7541_;
  assign new_n7568_ = new_n5578_ & new_n7567_;
  assign new_n7569_ = new_n5580_ & new_n7567_;
  assign new_n7570_ = ~new_n7568_ & ~new_n7569_;
  assign new_n7571_ = new_n7566_ & new_n7570_;
  assign new_n7572_ = new_n5590_ & new_n7567_;
  assign new_n7573_ = new_n5576_ & new_n7567_;
  assign new_n7574_ = new_n5587_ & new_n7567_;
  assign new_n7575_ = ~new_n7573_ & ~new_n7574_;
  assign new_n7576_ = ~new_n7572_ & new_n7575_;
  assign new_n7577_ = new_n7571_ & new_n7576_;
  assign new_n7578_ = new_n7563_ & new_n7577_;
  assign new_n7579_ = new_n7549_ & new_n7578_;
  assign new_n7580_ = new_n5594_ & new_n7567_;
  assign new_n7581_ = new_n4272_ & new_n7541_;
  assign new_n7582_ = new_n5596_ & new_n7581_;
  assign new_n7583_ = ~new_n7580_ & ~new_n7582_;
  assign new_n7584_ = new_n5600_ & new_n7581_;
  assign new_n7585_ = new_n5602_ & new_n7581_;
  assign new_n7586_ = ~new_n7584_ & ~new_n7585_;
  assign new_n7587_ = new_n7583_ & new_n7586_;
  assign new_n7588_ = new_n5605_ & new_n7581_;
  assign new_n7589_ = new_n5608_ & new_n7581_;
  assign new_n7590_ = ~new_n7588_ & ~new_n7589_;
  assign new_n7591_ = new_n5614_ & new_n7581_;
  assign new_n7592_ = new_n4277_ & new_n7541_;
  assign new_n7593_ = new_n5578_ & new_n7592_;
  assign new_n7594_ = ~new_n7591_ & ~new_n7593_;
  assign new_n7595_ = new_n7590_ & new_n7594_;
  assign new_n7596_ = new_n7587_ & new_n7595_;
  assign new_n7597_ = new_n5580_ & new_n7592_;
  assign new_n7598_ = new_n5576_ & new_n7592_;
  assign new_n7599_ = ~new_n7597_ & ~new_n7598_;
  assign new_n7600_ = new_n5587_ & new_n7592_;
  assign new_n7601_ = new_n5590_ & new_n7592_;
  assign new_n7602_ = ~new_n7600_ & ~new_n7601_;
  assign new_n7603_ = new_n7599_ & new_n7602_;
  assign new_n7604_ = new_n4280_ & new_n7541_;
  assign new_n7605_ = new_n5600_ & new_n7604_;
  assign new_n7606_ = new_n5594_ & new_n7592_;
  assign new_n7607_ = new_n5596_ & new_n7604_;
  assign new_n7608_ = ~new_n7606_ & ~new_n7607_;
  assign new_n7609_ = ~new_n7605_ & new_n7608_;
  assign new_n7610_ = new_n7603_ & new_n7609_;
  assign new_n7611_ = new_n7596_ & new_n7610_;
  assign new_n7612_ = new_n5602_ & new_n7604_;
  assign new_n7613_ = new_n5605_ & new_n7604_;
  assign new_n7614_ = ~new_n7612_ & ~new_n7613_;
  assign new_n7615_ = new_n5608_ & new_n7604_;
  assign new_n7616_ = new_n5614_ & new_n7604_;
  assign new_n7617_ = ~new_n7615_ & ~new_n7616_;
  assign new_n7618_ = new_n7614_ & new_n7617_;
  assign new_n7619_ = new_n4284_ & new_n7541_;
  assign new_n7620_ = new_n5576_ & new_n7619_;
  assign new_n7621_ = new_n5578_ & new_n7619_;
  assign new_n7622_ = new_n5580_ & new_n7619_;
  assign new_n7623_ = ~new_n7621_ & ~new_n7622_;
  assign new_n7624_ = ~new_n7620_ & new_n7623_;
  assign new_n7625_ = new_n7618_ & new_n7624_;
  assign new_n7626_ = new_n5587_ & new_n7619_;
  assign new_n7627_ = new_n5590_ & new_n7619_;
  assign new_n7628_ = ~new_n7626_ & ~new_n7627_;
  assign new_n7629_ = new_n5594_ & new_n7619_;
  assign new_n7630_ = new_n4287_ & new_n7541_;
  assign new_n7631_ = new_n5596_ & new_n7630_;
  assign new_n7632_ = ~new_n7629_ & ~new_n7631_;
  assign new_n7633_ = new_n7628_ & new_n7632_;
  assign new_n7634_ = new_n5605_ & new_n7630_;
  assign new_n7635_ = new_n5600_ & new_n7630_;
  assign new_n7636_ = new_n5602_ & new_n7630_;
  assign new_n7637_ = ~new_n7635_ & ~new_n7636_;
  assign new_n7638_ = ~new_n7634_ & new_n7637_;
  assign new_n7639_ = new_n7633_ & new_n7638_;
  assign new_n7640_ = new_n7625_ & new_n7639_;
  assign new_n7641_ = new_n7611_ & new_n7640_;
  assign new_n7642_ = new_n7579_ & new_n7641_;
  assign new_n7643_ = new_n7518_ & new_n7642_;
  assign new_n7644_ = new_n5608_ & new_n7630_;
  assign new_n7645_ = new_n5614_ & new_n7630_;
  assign new_n7646_ = ~new_n7644_ & ~new_n7645_;
  assign new_n7647_ = new_n4295_ & new_n7541_;
  assign new_n7648_ = new_n5690_ & new_n7647_;
  assign new_n7649_ = new_n5694_ & new_n7647_;
  assign new_n7650_ = ~new_n7648_ & ~new_n7649_;
  assign new_n7651_ = new_n7646_ & new_n7650_;
  assign new_n7652_ = new_n5697_ & new_n7647_;
  assign new_n7653_ = new_n5705_ & new_n7647_;
  assign new_n7654_ = ~new_n7652_ & ~new_n7653_;
  assign new_n7655_ = new_n5708_ & new_n7647_;
  assign new_n7656_ = new_n5702_ & new_n7647_;
  assign new_n7657_ = ~new_n7655_ & ~new_n7656_;
  assign new_n7658_ = new_n7654_ & new_n7657_;
  assign new_n7659_ = new_n7651_ & new_n7658_;
  assign new_n7660_ = new_n5714_ & new_n7647_;
  assign new_n7661_ = new_n5717_ & new_n7647_;
  assign new_n7662_ = ~new_n7660_ & ~new_n7661_;
  assign new_n7663_ = new_n5720_ & new_n7647_;
  assign new_n7664_ = new_n5722_ & new_n7647_;
  assign new_n7665_ = ~new_n7663_ & ~new_n7664_;
  assign new_n7666_ = new_n7662_ & new_n7665_;
  assign new_n7667_ = new_n5726_ & new_n7647_;
  assign new_n7668_ = new_n5728_ & new_n7647_;
  assign new_n7669_ = new_n5730_ & new_n7647_;
  assign new_n7670_ = ~new_n7668_ & ~new_n7669_;
  assign new_n7671_ = ~new_n7667_ & new_n7670_;
  assign new_n7672_ = new_n7666_ & new_n7671_;
  assign new_n7673_ = new_n7659_ & new_n7672_;
  assign new_n7674_ = new_n5737_ & new_n7647_;
  assign new_n7675_ = new_n5739_ & new_n7647_;
  assign new_n7676_ = ~new_n7674_ & ~new_n7675_;
  assign new_n7677_ = new_n5742_ & new_n7647_;
  assign new_n7678_ = ~A236 & ~A235;
  assign new_n7679_ = ~A234 & new_n7678_;
  assign new_n7680_ = ~A233 & A232;
  assign new_n7681_ = new_n7679_ & new_n7680_;
  assign new_n7682_ = ~A168 & new_n264_;
  assign new_n7683_ = new_n40_ & new_n7682_;
  assign new_n7684_ = new_n7681_ & new_n7683_;
  assign new_n7685_ = ~new_n7677_ & ~new_n7684_;
  assign new_n7686_ = new_n7676_ & new_n7685_;
  assign new_n7687_ = A233 & ~A232;
  assign new_n7688_ = new_n7679_ & new_n7687_;
  assign new_n7689_ = ~A168 & new_n282_;
  assign new_n7690_ = new_n40_ & new_n7689_;
  assign new_n7691_ = new_n7688_ & new_n7690_;
  assign new_n7692_ = new_n7683_ & new_n7688_;
  assign new_n7693_ = new_n7681_ & new_n7690_;
  assign new_n7694_ = ~new_n7692_ & ~new_n7693_;
  assign new_n7695_ = ~new_n7691_ & new_n7694_;
  assign new_n7696_ = new_n7686_ & new_n7695_;
  assign new_n7697_ = new_n383_ & new_n5689_;
  assign new_n7698_ = new_n7127_ & new_n7697_;
  assign new_n7699_ = new_n383_ & new_n5693_;
  assign new_n7700_ = new_n7127_ & new_n7699_;
  assign new_n7701_ = ~new_n7698_ & ~new_n7700_;
  assign new_n7702_ = new_n383_ & new_n5696_;
  assign new_n7703_ = new_n7127_ & new_n7702_;
  assign new_n7704_ = new_n383_ & new_n5704_;
  assign new_n7705_ = new_n7127_ & new_n7704_;
  assign new_n7706_ = ~new_n7703_ & ~new_n7705_;
  assign new_n7707_ = new_n7701_ & new_n7706_;
  assign new_n7708_ = new_n383_ & new_n5713_;
  assign new_n7709_ = new_n7127_ & new_n7708_;
  assign new_n7710_ = new_n383_ & new_n5707_;
  assign new_n7711_ = new_n7127_ & new_n7710_;
  assign new_n7712_ = new_n383_ & new_n5701_;
  assign new_n7713_ = new_n7127_ & new_n7712_;
  assign new_n7714_ = ~new_n7711_ & ~new_n7713_;
  assign new_n7715_ = ~new_n7709_ & new_n7714_;
  assign new_n7716_ = new_n7707_ & new_n7715_;
  assign new_n7717_ = new_n7696_ & new_n7716_;
  assign new_n7718_ = new_n7673_ & new_n7717_;
  assign new_n7719_ = new_n383_ & new_n5716_;
  assign new_n7720_ = new_n7127_ & new_n7719_;
  assign new_n7721_ = new_n409_ & new_n5689_;
  assign new_n7722_ = new_n7135_ & new_n7721_;
  assign new_n7723_ = ~new_n7720_ & ~new_n7722_;
  assign new_n7724_ = new_n409_ & new_n5693_;
  assign new_n7725_ = new_n7135_ & new_n7724_;
  assign new_n7726_ = new_n409_ & new_n5696_;
  assign new_n7727_ = new_n7135_ & new_n7726_;
  assign new_n7728_ = ~new_n7725_ & ~new_n7727_;
  assign new_n7729_ = new_n7723_ & new_n7728_;
  assign new_n7730_ = new_n409_ & new_n5704_;
  assign new_n7731_ = new_n7135_ & new_n7730_;
  assign new_n7732_ = new_n409_ & new_n5707_;
  assign new_n7733_ = new_n7135_ & new_n7732_;
  assign new_n7734_ = ~new_n7731_ & ~new_n7733_;
  assign new_n7735_ = new_n409_ & new_n5701_;
  assign new_n7736_ = new_n7135_ & new_n7735_;
  assign new_n7737_ = new_n409_ & new_n5713_;
  assign new_n7738_ = new_n7135_ & new_n7737_;
  assign new_n7739_ = ~new_n7736_ & ~new_n7738_;
  assign new_n7740_ = new_n7734_ & new_n7739_;
  assign new_n7741_ = new_n7729_ & new_n7740_;
  assign new_n7742_ = new_n409_ & new_n5716_;
  assign new_n7743_ = new_n7135_ & new_n7742_;
  assign new_n7744_ = new_n7154_ & new_n7697_;
  assign new_n7745_ = ~new_n7743_ & ~new_n7744_;
  assign new_n7746_ = new_n7154_ & new_n7699_;
  assign new_n7747_ = new_n7154_ & new_n7702_;
  assign new_n7748_ = ~new_n7746_ & ~new_n7747_;
  assign new_n7749_ = new_n7745_ & new_n7748_;
  assign new_n7750_ = new_n7154_ & new_n7712_;
  assign new_n7751_ = new_n7154_ & new_n7704_;
  assign new_n7752_ = new_n7154_ & new_n7710_;
  assign new_n7753_ = ~new_n7751_ & ~new_n7752_;
  assign new_n7754_ = ~new_n7750_ & new_n7753_;
  assign new_n7755_ = new_n7749_ & new_n7754_;
  assign new_n7756_ = new_n7741_ & new_n7755_;
  assign new_n7757_ = new_n7154_ & new_n7708_;
  assign new_n7758_ = new_n7154_ & new_n7719_;
  assign new_n7759_ = ~new_n7757_ & ~new_n7758_;
  assign new_n7760_ = new_n7166_ & new_n7721_;
  assign new_n7761_ = new_n7166_ & new_n7724_;
  assign new_n7762_ = ~new_n7760_ & ~new_n7761_;
  assign new_n7763_ = new_n7759_ & new_n7762_;
  assign new_n7764_ = new_n7166_ & new_n7732_;
  assign new_n7765_ = new_n7166_ & new_n7726_;
  assign new_n7766_ = new_n7166_ & new_n7730_;
  assign new_n7767_ = ~new_n7765_ & ~new_n7766_;
  assign new_n7768_ = ~new_n7764_ & new_n7767_;
  assign new_n7769_ = new_n7763_ & new_n7768_;
  assign new_n7770_ = new_n7166_ & new_n7735_;
  assign new_n7771_ = new_n7166_ & new_n7737_;
  assign new_n7772_ = ~new_n7770_ & ~new_n7771_;
  assign new_n7773_ = new_n7166_ & new_n7742_;
  assign new_n7774_ = new_n7180_ & new_n7697_;
  assign new_n7775_ = ~new_n7773_ & ~new_n7774_;
  assign new_n7776_ = new_n7772_ & new_n7775_;
  assign new_n7777_ = new_n7180_ & new_n7704_;
  assign new_n7778_ = new_n7180_ & new_n7699_;
  assign new_n7779_ = new_n7180_ & new_n7702_;
  assign new_n7780_ = ~new_n7778_ & ~new_n7779_;
  assign new_n7781_ = ~new_n7777_ & new_n7780_;
  assign new_n7782_ = new_n7776_ & new_n7781_;
  assign new_n7783_ = new_n7769_ & new_n7782_;
  assign new_n7784_ = new_n7756_ & new_n7783_;
  assign new_n7785_ = new_n7718_ & new_n7784_;
  assign new_n7786_ = new_n7180_ & new_n7710_;
  assign new_n7787_ = new_n7180_ & new_n7712_;
  assign new_n7788_ = ~new_n7786_ & ~new_n7787_;
  assign new_n7789_ = new_n7180_ & new_n7708_;
  assign new_n7790_ = new_n7180_ & new_n7719_;
  assign new_n7791_ = ~new_n7789_ & ~new_n7790_;
  assign new_n7792_ = new_n7788_ & new_n7791_;
  assign new_n7793_ = new_n7192_ & new_n7721_;
  assign new_n7794_ = new_n7192_ & new_n7724_;
  assign new_n7795_ = ~new_n7793_ & ~new_n7794_;
  assign new_n7796_ = new_n7192_ & new_n7726_;
  assign new_n7797_ = new_n7192_ & new_n7730_;
  assign new_n7798_ = ~new_n7796_ & ~new_n7797_;
  assign new_n7799_ = new_n7795_ & new_n7798_;
  assign new_n7800_ = new_n7792_ & new_n7799_;
  assign new_n7801_ = new_n7192_ & new_n7732_;
  assign new_n7802_ = new_n7192_ & new_n7735_;
  assign new_n7803_ = ~new_n7801_ & ~new_n7802_;
  assign new_n7804_ = new_n7192_ & new_n7737_;
  assign new_n7805_ = new_n7192_ & new_n7742_;
  assign new_n7806_ = ~new_n7804_ & ~new_n7805_;
  assign new_n7807_ = new_n7803_ & new_n7806_;
  assign new_n7808_ = new_n7207_ & new_n7702_;
  assign new_n7809_ = new_n7207_ & new_n7697_;
  assign new_n7810_ = new_n7207_ & new_n7699_;
  assign new_n7811_ = ~new_n7809_ & ~new_n7810_;
  assign new_n7812_ = ~new_n7808_ & new_n7811_;
  assign new_n7813_ = new_n7807_ & new_n7812_;
  assign new_n7814_ = new_n7800_ & new_n7813_;
  assign new_n7815_ = new_n7207_ & new_n7704_;
  assign new_n7816_ = new_n7207_ & new_n7710_;
  assign new_n7817_ = ~new_n7815_ & ~new_n7816_;
  assign new_n7818_ = new_n7207_ & new_n7712_;
  assign new_n7819_ = new_n7207_ & new_n7708_;
  assign new_n7820_ = ~new_n7818_ & ~new_n7819_;
  assign new_n7821_ = new_n7817_ & new_n7820_;
  assign new_n7822_ = new_n7218_ & new_n7724_;
  assign new_n7823_ = new_n7207_ & new_n7719_;
  assign new_n7824_ = new_n7218_ & new_n7721_;
  assign new_n7825_ = ~new_n7823_ & ~new_n7824_;
  assign new_n7826_ = ~new_n7822_ & new_n7825_;
  assign new_n7827_ = new_n7821_ & new_n7826_;
  assign new_n7828_ = new_n7218_ & new_n7726_;
  assign new_n7829_ = new_n7218_ & new_n7730_;
  assign new_n7830_ = ~new_n7828_ & ~new_n7829_;
  assign new_n7831_ = new_n7218_ & new_n7732_;
  assign new_n7832_ = new_n7218_ & new_n7735_;
  assign new_n7833_ = ~new_n7831_ & ~new_n7832_;
  assign new_n7834_ = new_n7830_ & new_n7833_;
  assign new_n7835_ = new_n7260_ & new_n7697_;
  assign new_n7836_ = new_n7218_ & new_n7737_;
  assign new_n7837_ = new_n7218_ & new_n7742_;
  assign new_n7838_ = ~new_n7836_ & ~new_n7837_;
  assign new_n7839_ = ~new_n7835_ & new_n7838_;
  assign new_n7840_ = new_n7834_ & new_n7839_;
  assign new_n7841_ = new_n7827_ & new_n7840_;
  assign new_n7842_ = new_n7814_ & new_n7841_;
  assign new_n7843_ = new_n7260_ & new_n7699_;
  assign new_n7844_ = new_n7260_ & new_n7702_;
  assign new_n7845_ = ~new_n7843_ & ~new_n7844_;
  assign new_n7846_ = new_n7260_ & new_n7704_;
  assign new_n7847_ = new_n7260_ & new_n7710_;
  assign new_n7848_ = ~new_n7846_ & ~new_n7847_;
  assign new_n7849_ = new_n7845_ & new_n7848_;
  assign new_n7850_ = new_n7260_ & new_n7719_;
  assign new_n7851_ = new_n7260_ & new_n7712_;
  assign new_n7852_ = new_n7260_ & new_n7708_;
  assign new_n7853_ = ~new_n7851_ & ~new_n7852_;
  assign new_n7854_ = ~new_n7850_ & new_n7853_;
  assign new_n7855_ = new_n7849_ & new_n7854_;
  assign new_n7856_ = new_n7278_ & new_n7721_;
  assign new_n7857_ = new_n7278_ & new_n7724_;
  assign new_n7858_ = ~new_n7856_ & ~new_n7857_;
  assign new_n7859_ = new_n7278_ & new_n7726_;
  assign new_n7860_ = new_n7278_ & new_n7730_;
  assign new_n7861_ = ~new_n7859_ & ~new_n7860_;
  assign new_n7862_ = new_n7858_ & new_n7861_;
  assign new_n7863_ = new_n7278_ & new_n7737_;
  assign new_n7864_ = new_n7278_ & new_n7732_;
  assign new_n7865_ = new_n7278_ & new_n7735_;
  assign new_n7866_ = ~new_n7864_ & ~new_n7865_;
  assign new_n7867_ = ~new_n7863_ & new_n7866_;
  assign new_n7868_ = new_n7862_ & new_n7867_;
  assign new_n7869_ = new_n7855_ & new_n7868_;
  assign new_n7870_ = new_n7278_ & new_n7742_;
  assign new_n7871_ = new_n7290_ & new_n7697_;
  assign new_n7872_ = ~new_n7870_ & ~new_n7871_;
  assign new_n7873_ = new_n7290_ & new_n7699_;
  assign new_n7874_ = new_n7290_ & new_n7702_;
  assign new_n7875_ = ~new_n7873_ & ~new_n7874_;
  assign new_n7876_ = new_n7872_ & new_n7875_;
  assign new_n7877_ = new_n7290_ & new_n7712_;
  assign new_n7878_ = new_n7290_ & new_n7704_;
  assign new_n7879_ = new_n7290_ & new_n7710_;
  assign new_n7880_ = ~new_n7878_ & ~new_n7879_;
  assign new_n7881_ = ~new_n7877_ & new_n7880_;
  assign new_n7882_ = new_n7876_ & new_n7881_;
  assign new_n7883_ = new_n7290_ & new_n7708_;
  assign new_n7884_ = new_n7290_ & new_n7719_;
  assign new_n7885_ = ~new_n7883_ & ~new_n7884_;
  assign new_n7886_ = new_n7304_ & new_n7721_;
  assign new_n7887_ = new_n7304_ & new_n7724_;
  assign new_n7888_ = ~new_n7886_ & ~new_n7887_;
  assign new_n7889_ = new_n7885_ & new_n7888_;
  assign new_n7890_ = new_n7304_ & new_n7732_;
  assign new_n7891_ = new_n7304_ & new_n7726_;
  assign new_n7892_ = new_n7304_ & new_n7730_;
  assign new_n7893_ = ~new_n7891_ & ~new_n7892_;
  assign new_n7894_ = ~new_n7890_ & new_n7893_;
  assign new_n7895_ = new_n7889_ & new_n7894_;
  assign new_n7896_ = new_n7882_ & new_n7895_;
  assign new_n7897_ = new_n7869_ & new_n7896_;
  assign new_n7898_ = new_n7842_ & new_n7897_;
  assign new_n7899_ = new_n7785_ & new_n7898_;
  assign new_n7900_ = new_n7643_ & new_n7899_;
  assign new_n7901_ = new_n7304_ & new_n7735_;
  assign new_n7902_ = new_n7304_ & new_n7737_;
  assign new_n7903_ = ~new_n7901_ & ~new_n7902_;
  assign new_n7904_ = new_n7304_ & new_n7742_;
  assign new_n7905_ = new_n7316_ & new_n7697_;
  assign new_n7906_ = ~new_n7904_ & ~new_n7905_;
  assign new_n7907_ = new_n7903_ & new_n7906_;
  assign new_n7908_ = new_n7316_ & new_n7699_;
  assign new_n7909_ = new_n7316_ & new_n7702_;
  assign new_n7910_ = ~new_n7908_ & ~new_n7909_;
  assign new_n7911_ = new_n7316_ & new_n7704_;
  assign new_n7912_ = new_n7316_ & new_n7710_;
  assign new_n7913_ = ~new_n7911_ & ~new_n7912_;
  assign new_n7914_ = new_n7910_ & new_n7913_;
  assign new_n7915_ = new_n7907_ & new_n7914_;
  assign new_n7916_ = new_n7316_ & new_n7712_;
  assign new_n7917_ = new_n7316_ & new_n7708_;
  assign new_n7918_ = ~new_n7916_ & ~new_n7917_;
  assign new_n7919_ = new_n7316_ & new_n7719_;
  assign new_n7920_ = new_n7331_ & new_n7721_;
  assign new_n7921_ = ~new_n7919_ & ~new_n7920_;
  assign new_n7922_ = new_n7918_ & new_n7921_;
  assign new_n7923_ = new_n7331_ & new_n7730_;
  assign new_n7924_ = new_n7331_ & new_n7724_;
  assign new_n7925_ = new_n7331_ & new_n7726_;
  assign new_n7926_ = ~new_n7924_ & ~new_n7925_;
  assign new_n7927_ = ~new_n7923_ & new_n7926_;
  assign new_n7928_ = new_n7922_ & new_n7927_;
  assign new_n7929_ = new_n7915_ & new_n7928_;
  assign new_n7930_ = new_n7331_ & new_n7732_;
  assign new_n7931_ = new_n7331_ & new_n7735_;
  assign new_n7932_ = ~new_n7930_ & ~new_n7931_;
  assign new_n7933_ = new_n7331_ & new_n7737_;
  assign new_n7934_ = new_n7331_ & new_n7742_;
  assign new_n7935_ = ~new_n7933_ & ~new_n7934_;
  assign new_n7936_ = new_n7932_ & new_n7935_;
  assign new_n7937_ = new_n7339_ & new_n7702_;
  assign new_n7938_ = new_n7339_ & new_n7697_;
  assign new_n7939_ = new_n7339_ & new_n7699_;
  assign new_n7940_ = ~new_n7938_ & ~new_n7939_;
  assign new_n7941_ = ~new_n7937_ & new_n7940_;
  assign new_n7942_ = new_n7936_ & new_n7941_;
  assign new_n7943_ = new_n7339_ & new_n7704_;
  assign new_n7944_ = new_n7339_ & new_n7710_;
  assign new_n7945_ = ~new_n7943_ & ~new_n7944_;
  assign new_n7946_ = new_n7339_ & new_n7712_;
  assign new_n7947_ = new_n7339_ & new_n7708_;
  assign new_n7948_ = ~new_n7946_ & ~new_n7947_;
  assign new_n7949_ = new_n7945_ & new_n7948_;
  assign new_n7950_ = new_n7353_ & new_n7724_;
  assign new_n7951_ = new_n7339_ & new_n7719_;
  assign new_n7952_ = new_n7353_ & new_n7721_;
  assign new_n7953_ = ~new_n7951_ & ~new_n7952_;
  assign new_n7954_ = ~new_n7950_ & new_n7953_;
  assign new_n7955_ = new_n7949_ & new_n7954_;
  assign new_n7956_ = new_n7942_ & new_n7955_;
  assign new_n7957_ = new_n7929_ & new_n7956_;
  assign new_n7958_ = new_n7353_ & new_n7726_;
  assign new_n7959_ = new_n7353_ & new_n7730_;
  assign new_n7960_ = ~new_n7958_ & ~new_n7959_;
  assign new_n7961_ = new_n7353_ & new_n7732_;
  assign new_n7962_ = new_n7353_ & new_n7735_;
  assign new_n7963_ = ~new_n7961_ & ~new_n7962_;
  assign new_n7964_ = new_n7960_ & new_n7963_;
  assign new_n7965_ = new_n7353_ & new_n7737_;
  assign new_n7966_ = new_n7353_ & new_n7742_;
  assign new_n7967_ = ~new_n7965_ & ~new_n7966_;
  assign new_n7968_ = new_n7405_ & new_n7697_;
  assign new_n7969_ = new_n7405_ & new_n7699_;
  assign new_n7970_ = ~new_n7968_ & ~new_n7969_;
  assign new_n7971_ = new_n7967_ & new_n7970_;
  assign new_n7972_ = new_n7964_ & new_n7971_;
  assign new_n7973_ = new_n7405_ & new_n7702_;
  assign new_n7974_ = new_n7405_ & new_n7704_;
  assign new_n7975_ = ~new_n7973_ & ~new_n7974_;
  assign new_n7976_ = new_n7405_ & new_n7710_;
  assign new_n7977_ = new_n7405_ & new_n7712_;
  assign new_n7978_ = ~new_n7976_ & ~new_n7977_;
  assign new_n7979_ = new_n7975_ & new_n7978_;
  assign new_n7980_ = new_n7418_ & new_n7721_;
  assign new_n7981_ = new_n7405_ & new_n7708_;
  assign new_n7982_ = new_n7405_ & new_n7719_;
  assign new_n7983_ = ~new_n7981_ & ~new_n7982_;
  assign new_n7984_ = ~new_n7980_ & new_n7983_;
  assign new_n7985_ = new_n7979_ & new_n7984_;
  assign new_n7986_ = new_n7972_ & new_n7985_;
  assign new_n7987_ = new_n7418_ & new_n7724_;
  assign new_n7988_ = new_n7418_ & new_n7726_;
  assign new_n7989_ = ~new_n7987_ & ~new_n7988_;
  assign new_n7990_ = new_n7418_ & new_n7730_;
  assign new_n7991_ = new_n7418_ & new_n7732_;
  assign new_n7992_ = ~new_n7990_ & ~new_n7991_;
  assign new_n7993_ = new_n7989_ & new_n7992_;
  assign new_n7994_ = new_n7418_ & new_n7742_;
  assign new_n7995_ = new_n7418_ & new_n7735_;
  assign new_n7996_ = new_n7418_ & new_n7737_;
  assign new_n7997_ = ~new_n7995_ & ~new_n7996_;
  assign new_n7998_ = ~new_n7994_ & new_n7997_;
  assign new_n7999_ = new_n7993_ & new_n7998_;
  assign new_n8000_ = new_n7430_ & new_n7697_;
  assign new_n8001_ = new_n7430_ & new_n7699_;
  assign new_n8002_ = ~new_n8000_ & ~new_n8001_;
  assign new_n8003_ = new_n7430_ & new_n7702_;
  assign new_n8004_ = new_n7430_ & new_n7704_;
  assign new_n8005_ = ~new_n8003_ & ~new_n8004_;
  assign new_n8006_ = new_n8002_ & new_n8005_;
  assign new_n8007_ = new_n7430_ & new_n7708_;
  assign new_n8008_ = new_n7430_ & new_n7710_;
  assign new_n8009_ = new_n7430_ & new_n7712_;
  assign new_n8010_ = ~new_n8008_ & ~new_n8009_;
  assign new_n8011_ = ~new_n8007_ & new_n8010_;
  assign new_n8012_ = new_n8006_ & new_n8011_;
  assign new_n8013_ = new_n7999_ & new_n8012_;
  assign new_n8014_ = new_n7986_ & new_n8013_;
  assign new_n8015_ = new_n7957_ & new_n8014_;
  assign new_n8016_ = new_n7430_ & new_n7719_;
  assign new_n8017_ = new_n7443_ & new_n7721_;
  assign new_n8018_ = ~new_n8016_ & ~new_n8017_;
  assign new_n8019_ = new_n7443_ & new_n7724_;
  assign new_n8020_ = new_n7443_ & new_n7726_;
  assign new_n8021_ = ~new_n8019_ & ~new_n8020_;
  assign new_n8022_ = new_n8018_ & new_n8021_;
  assign new_n8023_ = new_n7443_ & new_n7730_;
  assign new_n8024_ = new_n7443_ & new_n7732_;
  assign new_n8025_ = ~new_n8023_ & ~new_n8024_;
  assign new_n8026_ = new_n7443_ & new_n7735_;
  assign new_n8027_ = new_n7443_ & new_n7737_;
  assign new_n8028_ = ~new_n8026_ & ~new_n8027_;
  assign new_n8029_ = new_n8025_ & new_n8028_;
  assign new_n8030_ = new_n8022_ & new_n8029_;
  assign new_n8031_ = new_n7443_ & new_n7742_;
  assign new_n8032_ = new_n7457_ & new_n7697_;
  assign new_n8033_ = ~new_n8031_ & ~new_n8032_;
  assign new_n8034_ = new_n7457_ & new_n7699_;
  assign new_n8035_ = new_n7457_ & new_n7702_;
  assign new_n8036_ = ~new_n8034_ & ~new_n8035_;
  assign new_n8037_ = new_n8033_ & new_n8036_;
  assign new_n8038_ = new_n7457_ & new_n7712_;
  assign new_n8039_ = new_n7457_ & new_n7704_;
  assign new_n8040_ = new_n7457_ & new_n7710_;
  assign new_n8041_ = ~new_n8039_ & ~new_n8040_;
  assign new_n8042_ = ~new_n8038_ & new_n8041_;
  assign new_n8043_ = new_n8037_ & new_n8042_;
  assign new_n8044_ = new_n8030_ & new_n8043_;
  assign new_n8045_ = new_n7457_ & new_n7708_;
  assign new_n8046_ = new_n7457_ & new_n7719_;
  assign new_n8047_ = ~new_n8045_ & ~new_n8046_;
  assign new_n8048_ = new_n7468_ & new_n7721_;
  assign new_n8049_ = new_n7468_ & new_n7724_;
  assign new_n8050_ = ~new_n8048_ & ~new_n8049_;
  assign new_n8051_ = new_n8047_ & new_n8050_;
  assign new_n8052_ = new_n7468_ & new_n7732_;
  assign new_n8053_ = new_n7468_ & new_n7726_;
  assign new_n8054_ = new_n7468_ & new_n7730_;
  assign new_n8055_ = ~new_n8053_ & ~new_n8054_;
  assign new_n8056_ = ~new_n8052_ & new_n8055_;
  assign new_n8057_ = new_n8051_ & new_n8056_;
  assign new_n8058_ = new_n7468_ & new_n7735_;
  assign new_n8059_ = new_n7468_ & new_n7737_;
  assign new_n8060_ = ~new_n8058_ & ~new_n8059_;
  assign new_n8061_ = new_n7468_ & new_n7742_;
  assign new_n8062_ = new_n7480_ & new_n7697_;
  assign new_n8063_ = ~new_n8061_ & ~new_n8062_;
  assign new_n8064_ = new_n8060_ & new_n8063_;
  assign new_n8065_ = new_n7480_ & new_n7704_;
  assign new_n8066_ = new_n7480_ & new_n7699_;
  assign new_n8067_ = new_n7480_ & new_n7702_;
  assign new_n8068_ = ~new_n8066_ & ~new_n8067_;
  assign new_n8069_ = ~new_n8065_ & new_n8068_;
  assign new_n8070_ = new_n8064_ & new_n8069_;
  assign new_n8071_ = new_n8057_ & new_n8070_;
  assign new_n8072_ = new_n8044_ & new_n8071_;
  assign new_n8073_ = new_n7480_ & new_n7710_;
  assign new_n8074_ = new_n7480_ & new_n7712_;
  assign new_n8075_ = ~new_n8073_ & ~new_n8074_;
  assign new_n8076_ = new_n7480_ & new_n7708_;
  assign new_n8077_ = new_n7480_ & new_n7719_;
  assign new_n8078_ = ~new_n8076_ & ~new_n8077_;
  assign new_n8079_ = new_n8075_ & new_n8078_;
  assign new_n8080_ = new_n7495_ & new_n7721_;
  assign new_n8081_ = new_n7495_ & new_n7724_;
  assign new_n8082_ = ~new_n8080_ & ~new_n8081_;
  assign new_n8083_ = new_n7495_ & new_n7726_;
  assign new_n8084_ = new_n7495_ & new_n7730_;
  assign new_n8085_ = ~new_n8083_ & ~new_n8084_;
  assign new_n8086_ = new_n8082_ & new_n8085_;
  assign new_n8087_ = new_n8079_ & new_n8086_;
  assign new_n8088_ = new_n7495_ & new_n7732_;
  assign new_n8089_ = new_n7495_ & new_n7735_;
  assign new_n8090_ = ~new_n8088_ & ~new_n8089_;
  assign new_n8091_ = new_n7495_ & new_n7737_;
  assign new_n8092_ = new_n7495_ & new_n7742_;
  assign new_n8093_ = ~new_n8091_ & ~new_n8092_;
  assign new_n8094_ = new_n8090_ & new_n8093_;
  assign new_n8095_ = new_n7542_ & new_n7702_;
  assign new_n8096_ = new_n7542_ & new_n7697_;
  assign new_n8097_ = new_n7542_ & new_n7699_;
  assign new_n8098_ = ~new_n8096_ & ~new_n8097_;
  assign new_n8099_ = ~new_n8095_ & new_n8098_;
  assign new_n8100_ = new_n8094_ & new_n8099_;
  assign new_n8101_ = new_n8087_ & new_n8100_;
  assign new_n8102_ = new_n7542_ & new_n7704_;
  assign new_n8103_ = new_n7542_ & new_n7710_;
  assign new_n8104_ = ~new_n8102_ & ~new_n8103_;
  assign new_n8105_ = new_n7542_ & new_n7712_;
  assign new_n8106_ = new_n7542_ & new_n7708_;
  assign new_n8107_ = ~new_n8105_ & ~new_n8106_;
  assign new_n8108_ = new_n8104_ & new_n8107_;
  assign new_n8109_ = new_n7554_ & new_n7724_;
  assign new_n8110_ = new_n7542_ & new_n7719_;
  assign new_n8111_ = new_n7554_ & new_n7721_;
  assign new_n8112_ = ~new_n8110_ & ~new_n8111_;
  assign new_n8113_ = ~new_n8109_ & new_n8112_;
  assign new_n8114_ = new_n8108_ & new_n8113_;
  assign new_n8115_ = new_n7554_ & new_n7726_;
  assign new_n8116_ = new_n7554_ & new_n7730_;
  assign new_n8117_ = ~new_n8115_ & ~new_n8116_;
  assign new_n8118_ = new_n7554_ & new_n7732_;
  assign new_n8119_ = new_n7554_ & new_n7735_;
  assign new_n8120_ = ~new_n8118_ & ~new_n8119_;
  assign new_n8121_ = new_n8117_ & new_n8120_;
  assign new_n8122_ = new_n7567_ & new_n7697_;
  assign new_n8123_ = new_n7554_ & new_n7737_;
  assign new_n8124_ = new_n7554_ & new_n7742_;
  assign new_n8125_ = ~new_n8123_ & ~new_n8124_;
  assign new_n8126_ = ~new_n8122_ & new_n8125_;
  assign new_n8127_ = new_n8121_ & new_n8126_;
  assign new_n8128_ = new_n8114_ & new_n8127_;
  assign new_n8129_ = new_n8101_ & new_n8128_;
  assign new_n8130_ = new_n8072_ & new_n8129_;
  assign new_n8131_ = new_n8015_ & new_n8130_;
  assign new_n8132_ = new_n7567_ & new_n7699_;
  assign new_n8133_ = new_n7567_ & new_n7702_;
  assign new_n8134_ = ~new_n8132_ & ~new_n8133_;
  assign new_n8135_ = new_n7567_ & new_n7704_;
  assign new_n8136_ = new_n7567_ & new_n7710_;
  assign new_n8137_ = ~new_n8135_ & ~new_n8136_;
  assign new_n8138_ = new_n8134_ & new_n8137_;
  assign new_n8139_ = new_n7567_ & new_n7712_;
  assign new_n8140_ = new_n7567_ & new_n7708_;
  assign new_n8141_ = ~new_n8139_ & ~new_n8140_;
  assign new_n8142_ = new_n7567_ & new_n7719_;
  assign new_n8143_ = new_n7581_ & new_n7721_;
  assign new_n8144_ = ~new_n8142_ & ~new_n8143_;
  assign new_n8145_ = new_n8141_ & new_n8144_;
  assign new_n8146_ = new_n8138_ & new_n8145_;
  assign new_n8147_ = new_n7581_ & new_n7724_;
  assign new_n8148_ = new_n7581_ & new_n7726_;
  assign new_n8149_ = ~new_n8147_ & ~new_n8148_;
  assign new_n8150_ = new_n7581_ & new_n7730_;
  assign new_n8151_ = new_n7581_ & new_n7732_;
  assign new_n8152_ = ~new_n8150_ & ~new_n8151_;
  assign new_n8153_ = new_n8149_ & new_n8152_;
  assign new_n8154_ = new_n7581_ & new_n7742_;
  assign new_n8155_ = new_n7581_ & new_n7735_;
  assign new_n8156_ = new_n7581_ & new_n7737_;
  assign new_n8157_ = ~new_n8155_ & ~new_n8156_;
  assign new_n8158_ = ~new_n8154_ & new_n8157_;
  assign new_n8159_ = new_n8153_ & new_n8158_;
  assign new_n8160_ = new_n8146_ & new_n8159_;
  assign new_n8161_ = new_n7592_ & new_n7697_;
  assign new_n8162_ = new_n7592_ & new_n7699_;
  assign new_n8163_ = ~new_n8161_ & ~new_n8162_;
  assign new_n8164_ = new_n7592_ & new_n7702_;
  assign new_n8165_ = new_n7592_ & new_n7704_;
  assign new_n8166_ = ~new_n8164_ & ~new_n8165_;
  assign new_n8167_ = new_n8163_ & new_n8166_;
  assign new_n8168_ = new_n7592_ & new_n7708_;
  assign new_n8169_ = new_n7592_ & new_n7710_;
  assign new_n8170_ = new_n7592_ & new_n7712_;
  assign new_n8171_ = ~new_n8169_ & ~new_n8170_;
  assign new_n8172_ = ~new_n8168_ & new_n8171_;
  assign new_n8173_ = new_n8167_ & new_n8172_;
  assign new_n8174_ = new_n7592_ & new_n7719_;
  assign new_n8175_ = new_n7604_ & new_n7721_;
  assign new_n8176_ = ~new_n8174_ & ~new_n8175_;
  assign new_n8177_ = new_n7604_ & new_n7724_;
  assign new_n8178_ = new_n7604_ & new_n7726_;
  assign new_n8179_ = ~new_n8177_ & ~new_n8178_;
  assign new_n8180_ = new_n8176_ & new_n8179_;
  assign new_n8181_ = new_n7604_ & new_n7735_;
  assign new_n8182_ = new_n7604_ & new_n7730_;
  assign new_n8183_ = new_n7604_ & new_n7732_;
  assign new_n8184_ = ~new_n8182_ & ~new_n8183_;
  assign new_n8185_ = ~new_n8181_ & new_n8184_;
  assign new_n8186_ = new_n8180_ & new_n8185_;
  assign new_n8187_ = new_n8173_ & new_n8186_;
  assign new_n8188_ = new_n8160_ & new_n8187_;
  assign new_n8189_ = new_n7604_ & new_n7737_;
  assign new_n8190_ = new_n7604_ & new_n7742_;
  assign new_n8191_ = ~new_n8189_ & ~new_n8190_;
  assign new_n8192_ = new_n7619_ & new_n7697_;
  assign new_n8193_ = new_n7619_ & new_n7699_;
  assign new_n8194_ = ~new_n8192_ & ~new_n8193_;
  assign new_n8195_ = new_n8191_ & new_n8194_;
  assign new_n8196_ = new_n7619_ & new_n7702_;
  assign new_n8197_ = new_n7619_ & new_n7704_;
  assign new_n8198_ = ~new_n8196_ & ~new_n8197_;
  assign new_n8199_ = new_n7619_ & new_n7710_;
  assign new_n8200_ = new_n7619_ & new_n7712_;
  assign new_n8201_ = ~new_n8199_ & ~new_n8200_;
  assign new_n8202_ = new_n8198_ & new_n8201_;
  assign new_n8203_ = new_n8195_ & new_n8202_;
  assign new_n8204_ = new_n7619_ & new_n7708_;
  assign new_n8205_ = new_n7619_ & new_n7719_;
  assign new_n8206_ = ~new_n8204_ & ~new_n8205_;
  assign new_n8207_ = new_n7630_ & new_n7721_;
  assign new_n8208_ = new_n7630_ & new_n7724_;
  assign new_n8209_ = ~new_n8207_ & ~new_n8208_;
  assign new_n8210_ = new_n8206_ & new_n8209_;
  assign new_n8211_ = new_n7630_ & new_n7732_;
  assign new_n8212_ = new_n7630_ & new_n7726_;
  assign new_n8213_ = new_n7630_ & new_n7730_;
  assign new_n8214_ = ~new_n8212_ & ~new_n8213_;
  assign new_n8215_ = ~new_n8211_ & new_n8214_;
  assign new_n8216_ = new_n8210_ & new_n8215_;
  assign new_n8217_ = new_n8203_ & new_n8216_;
  assign new_n8218_ = new_n7630_ & new_n7735_;
  assign new_n8219_ = new_n7630_ & new_n7737_;
  assign new_n8220_ = ~new_n8218_ & ~new_n8219_;
  assign new_n8221_ = new_n7630_ & new_n7742_;
  assign new_n8222_ = ~A201 & new_n79_;
  assign new_n8223_ = new_n262_ & new_n8222_;
  assign new_n8224_ = new_n7681_ & new_n8223_;
  assign new_n8225_ = ~new_n8221_ & ~new_n8224_;
  assign new_n8226_ = new_n8220_ & new_n8225_;
  assign new_n8227_ = new_n276_ & new_n8222_;
  assign new_n8228_ = new_n7688_ & new_n8227_;
  assign new_n8229_ = new_n7688_ & new_n8223_;
  assign new_n8230_ = new_n7681_ & new_n8227_;
  assign new_n8231_ = ~new_n8229_ & ~new_n8230_;
  assign new_n8232_ = ~new_n8228_ & new_n8231_;
  assign new_n8233_ = new_n8226_ & new_n8232_;
  assign new_n8234_ = A236 & A234;
  assign new_n8235_ = ~A233 & new_n8234_;
  assign new_n8236_ = A232 & A166;
  assign new_n8237_ = new_n8235_ & new_n8236_;
  assign new_n8238_ = new_n41_ & new_n8237_;
  assign new_n8239_ = A235 & A234;
  assign new_n8240_ = ~A233 & new_n8239_;
  assign new_n8241_ = new_n8236_ & new_n8240_;
  assign new_n8242_ = new_n41_ & new_n8241_;
  assign new_n8243_ = ~new_n8238_ & ~new_n8242_;
  assign new_n8244_ = A233 & new_n8234_;
  assign new_n8245_ = ~A232 & A166;
  assign new_n8246_ = new_n8244_ & new_n8245_;
  assign new_n8247_ = new_n41_ & new_n8246_;
  assign new_n8248_ = A233 & new_n8239_;
  assign new_n8249_ = new_n8245_ & new_n8248_;
  assign new_n8250_ = new_n41_ & new_n8249_;
  assign new_n8251_ = ~new_n8247_ & ~new_n8250_;
  assign new_n8252_ = new_n8243_ & new_n8251_;
  assign new_n8253_ = ~A232 & ~A166;
  assign new_n8254_ = new_n8244_ & new_n8253_;
  assign new_n8255_ = new_n61_ & new_n8254_;
  assign new_n8256_ = A232 & ~A166;
  assign new_n8257_ = new_n8235_ & new_n8256_;
  assign new_n8258_ = new_n61_ & new_n8257_;
  assign new_n8259_ = new_n8240_ & new_n8256_;
  assign new_n8260_ = new_n61_ & new_n8259_;
  assign new_n8261_ = ~new_n8258_ & ~new_n8260_;
  assign new_n8262_ = ~new_n8255_ & new_n8261_;
  assign new_n8263_ = new_n8252_ & new_n8262_;
  assign new_n8264_ = new_n8233_ & new_n8263_;
  assign new_n8265_ = new_n8217_ & new_n8264_;
  assign new_n8266_ = new_n8188_ & new_n8265_;
  assign new_n8267_ = new_n8248_ & new_n8253_;
  assign new_n8268_ = new_n61_ & new_n8267_;
  assign new_n8269_ = new_n266_ & new_n7681_;
  assign new_n8270_ = ~new_n8268_ & ~new_n8269_;
  assign new_n8271_ = new_n266_ & new_n7688_;
  assign new_n8272_ = new_n283_ & new_n7681_;
  assign new_n8273_ = ~new_n8271_ & ~new_n8272_;
  assign new_n8274_ = new_n8270_ & new_n8273_;
  assign new_n8275_ = new_n283_ & new_n7688_;
  assign new_n8276_ = new_n296_ & new_n7681_;
  assign new_n8277_ = ~new_n8275_ & ~new_n8276_;
  assign new_n8278_ = new_n296_ & new_n7688_;
  assign new_n8279_ = new_n306_ & new_n7681_;
  assign new_n8280_ = ~new_n8278_ & ~new_n8279_;
  assign new_n8281_ = new_n8277_ & new_n8280_;
  assign new_n8282_ = new_n8274_ & new_n8281_;
  assign new_n8283_ = new_n306_ & new_n7688_;
  assign new_n8284_ = A232 & ~A203;
  assign new_n8285_ = new_n8235_ & new_n8284_;
  assign new_n8286_ = new_n263_ & new_n8285_;
  assign new_n8287_ = ~new_n8283_ & ~new_n8286_;
  assign new_n8288_ = new_n8240_ & new_n8284_;
  assign new_n8289_ = new_n263_ & new_n8288_;
  assign new_n8290_ = ~A232 & ~A203;
  assign new_n8291_ = new_n8244_ & new_n8290_;
  assign new_n8292_ = new_n263_ & new_n8291_;
  assign new_n8293_ = ~new_n8289_ & ~new_n8292_;
  assign new_n8294_ = new_n8287_ & new_n8293_;
  assign new_n8295_ = new_n782_ & new_n7688_;
  assign new_n8296_ = new_n8248_ & new_n8290_;
  assign new_n8297_ = new_n263_ & new_n8296_;
  assign new_n8298_ = new_n782_ & new_n7681_;
  assign new_n8299_ = ~new_n8297_ & ~new_n8298_;
  assign new_n8300_ = ~new_n8295_ & new_n8299_;
  assign new_n8301_ = new_n8294_ & new_n8300_;
  assign new_n8302_ = new_n8282_ & new_n8301_;
  assign new_n8303_ = new_n792_ & new_n7681_;
  assign new_n8304_ = new_n792_ & new_n7688_;
  assign new_n8305_ = ~new_n8303_ & ~new_n8304_;
  assign new_n8306_ = new_n277_ & new_n8285_;
  assign new_n8307_ = new_n277_ & new_n8288_;
  assign new_n8308_ = ~new_n8306_ & ~new_n8307_;
  assign new_n8309_ = new_n8305_ & new_n8308_;
  assign new_n8310_ = new_n821_ & new_n7681_;
  assign new_n8311_ = new_n277_ & new_n8291_;
  assign new_n8312_ = new_n277_ & new_n8296_;
  assign new_n8313_ = ~new_n8311_ & ~new_n8312_;
  assign new_n8314_ = ~new_n8310_ & new_n8313_;
  assign new_n8315_ = new_n8309_ & new_n8314_;
  assign new_n8316_ = new_n821_ & new_n7688_;
  assign new_n8317_ = new_n826_ & new_n7681_;
  assign new_n8318_ = ~new_n8316_ & ~new_n8317_;
  assign new_n8319_ = new_n826_ & new_n7688_;
  assign new_n8320_ = new_n7680_ & new_n8234_;
  assign new_n8321_ = new_n266_ & new_n8320_;
  assign new_n8322_ = ~new_n8319_ & ~new_n8321_;
  assign new_n8323_ = new_n8318_ & new_n8322_;
  assign new_n8324_ = new_n7687_ & new_n8239_;
  assign new_n8325_ = new_n266_ & new_n8324_;
  assign new_n8326_ = new_n7680_ & new_n8239_;
  assign new_n8327_ = new_n266_ & new_n8326_;
  assign new_n8328_ = new_n7687_ & new_n8234_;
  assign new_n8329_ = new_n266_ & new_n8328_;
  assign new_n8330_ = ~new_n8327_ & ~new_n8329_;
  assign new_n8331_ = ~new_n8325_ & new_n8330_;
  assign new_n8332_ = new_n8323_ & new_n8331_;
  assign new_n8333_ = new_n8315_ & new_n8332_;
  assign new_n8334_ = new_n8302_ & new_n8333_;
  assign new_n8335_ = new_n283_ & new_n8320_;
  assign new_n8336_ = new_n283_ & new_n8326_;
  assign new_n8337_ = ~new_n8335_ & ~new_n8336_;
  assign new_n8338_ = new_n283_ & new_n8328_;
  assign new_n8339_ = new_n283_ & new_n8324_;
  assign new_n8340_ = ~new_n8338_ & ~new_n8339_;
  assign new_n8341_ = new_n8337_ & new_n8340_;
  assign new_n8342_ = new_n296_ & new_n8328_;
  assign new_n8343_ = new_n296_ & new_n8320_;
  assign new_n8344_ = new_n296_ & new_n8326_;
  assign new_n8345_ = ~new_n8343_ & ~new_n8344_;
  assign new_n8346_ = ~new_n8342_ & new_n8345_;
  assign new_n8347_ = new_n8341_ & new_n8346_;
  assign new_n8348_ = new_n296_ & new_n8324_;
  assign new_n8349_ = new_n306_ & new_n8320_;
  assign new_n8350_ = ~new_n8348_ & ~new_n8349_;
  assign new_n8351_ = new_n306_ & new_n8326_;
  assign new_n8352_ = new_n306_ & new_n8328_;
  assign new_n8353_ = ~new_n8351_ & ~new_n8352_;
  assign new_n8354_ = new_n8350_ & new_n8353_;
  assign new_n8355_ = new_n782_ & new_n8326_;
  assign new_n8356_ = new_n306_ & new_n8324_;
  assign new_n8357_ = new_n782_ & new_n8320_;
  assign new_n8358_ = ~new_n8356_ & ~new_n8357_;
  assign new_n8359_ = ~new_n8355_ & new_n8358_;
  assign new_n8360_ = new_n8354_ & new_n8359_;
  assign new_n8361_ = new_n8347_ & new_n8360_;
  assign new_n8362_ = new_n782_ & new_n8328_;
  assign new_n8363_ = new_n782_ & new_n8324_;
  assign new_n8364_ = ~new_n8362_ & ~new_n8363_;
  assign new_n8365_ = new_n792_ & new_n8320_;
  assign new_n8366_ = new_n792_ & new_n8326_;
  assign new_n8367_ = ~new_n8365_ & ~new_n8366_;
  assign new_n8368_ = new_n8364_ & new_n8367_;
  assign new_n8369_ = new_n821_ & new_n8320_;
  assign new_n8370_ = new_n792_ & new_n8328_;
  assign new_n8371_ = new_n792_ & new_n8324_;
  assign new_n8372_ = ~new_n8370_ & ~new_n8371_;
  assign new_n8373_ = ~new_n8369_ & new_n8372_;
  assign new_n8374_ = new_n8368_ & new_n8373_;
  assign new_n8375_ = new_n821_ & new_n8326_;
  assign new_n8376_ = new_n821_ & new_n8328_;
  assign new_n8377_ = ~new_n8375_ & ~new_n8376_;
  assign new_n8378_ = new_n821_ & new_n8324_;
  assign new_n8379_ = new_n826_ & new_n8320_;
  assign new_n8380_ = ~new_n8378_ & ~new_n8379_;
  assign new_n8381_ = new_n8377_ & new_n8380_;
  assign new_n8382_ = new_n826_ & new_n8324_;
  assign new_n8383_ = new_n826_ & new_n8326_;
  assign new_n8384_ = new_n826_ & new_n8328_;
  assign new_n8385_ = ~new_n8383_ & ~new_n8384_;
  assign new_n8386_ = ~new_n8382_ & new_n8385_;
  assign new_n8387_ = new_n8381_ & new_n8386_;
  assign new_n8388_ = new_n8374_ & new_n8387_;
  assign new_n8389_ = new_n8361_ & new_n8388_;
  assign new_n8390_ = new_n8334_ & new_n8389_;
  assign new_n8391_ = new_n8266_ & new_n8390_;
  assign new_n8392_ = new_n8131_ & new_n8391_;
  assign new_n8393_ = new_n7900_ & new_n8392_;
  assign new_n8394_ = new_n7393_ & new_n8393_;
  assign new_n8395_ = new_n6422_ & new_n8394_;
  assign A139 = ~new_n4418_ | ~new_n8395_;
endmodule


