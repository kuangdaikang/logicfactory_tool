// Benchmark "c1355.blif" written by ABC on Fri Feb 25 15:12:57 2022

module c1355  ( 
    G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat,
    G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat,
    G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat,
    G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat,
    G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat,
    G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat,
    G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat,
    G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat,
    G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat,
    G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n421_, new_n422_, new_n423_, new_n424_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n450_, new_n451_, new_n452_, new_n453_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n506_, new_n507_, new_n508_, new_n509_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n528_, new_n529_, new_n530_, new_n531_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n573_, new_n574_, new_n575_, new_n576_;
  assign new_n74_ = G1gat & G29gat;
  assign new_n75_ = G1gat & ~new_n74_;
  assign new_n76_ = G29gat & ~new_n74_;
  assign new_n77_ = ~new_n75_ & ~new_n76_;
  assign new_n78_ = G57gat & G85gat;
  assign new_n79_ = G57gat & ~new_n78_;
  assign new_n80_ = G85gat & ~new_n78_;
  assign new_n81_ = ~new_n79_ & ~new_n80_;
  assign new_n82_ = ~new_n77_ & ~new_n81_;
  assign new_n83_ = ~new_n77_ & ~new_n82_;
  assign new_n84_ = ~new_n81_ & ~new_n82_;
  assign new_n85_ = ~new_n83_ & ~new_n84_;
  assign new_n86_ = G225gat & G233gat;
  assign new_n87_ = G113gat & G120gat;
  assign new_n88_ = G113gat & ~new_n87_;
  assign new_n89_ = G120gat & ~new_n87_;
  assign new_n90_ = ~new_n88_ & ~new_n89_;
  assign new_n91_ = G127gat & G134gat;
  assign new_n92_ = G127gat & ~new_n91_;
  assign new_n93_ = G134gat & ~new_n91_;
  assign new_n94_ = ~new_n92_ & ~new_n93_;
  assign new_n95_ = ~new_n90_ & ~new_n94_;
  assign new_n96_ = ~new_n90_ & ~new_n95_;
  assign new_n97_ = ~new_n94_ & ~new_n95_;
  assign new_n98_ = ~new_n96_ & ~new_n97_;
  assign new_n99_ = G141gat & G148gat;
  assign new_n100_ = G141gat & ~new_n99_;
  assign new_n101_ = G148gat & ~new_n99_;
  assign new_n102_ = ~new_n100_ & ~new_n101_;
  assign new_n103_ = G155gat & G162gat;
  assign new_n104_ = G155gat & ~new_n103_;
  assign new_n105_ = G162gat & ~new_n103_;
  assign new_n106_ = ~new_n104_ & ~new_n105_;
  assign new_n107_ = ~new_n102_ & ~new_n106_;
  assign new_n108_ = ~new_n102_ & ~new_n107_;
  assign new_n109_ = ~new_n106_ & ~new_n107_;
  assign new_n110_ = ~new_n108_ & ~new_n109_;
  assign new_n111_ = ~new_n98_ & ~new_n110_;
  assign new_n112_ = ~new_n98_ & ~new_n111_;
  assign new_n113_ = ~new_n110_ & ~new_n111_;
  assign new_n114_ = ~new_n112_ & ~new_n113_;
  assign new_n115_ = new_n86_ & ~new_n114_;
  assign new_n116_ = new_n86_ & ~new_n115_;
  assign new_n117_ = ~new_n114_ & ~new_n115_;
  assign new_n118_ = ~new_n116_ & ~new_n117_;
  assign new_n119_ = ~new_n85_ & ~new_n118_;
  assign new_n120_ = ~new_n85_ & ~new_n119_;
  assign new_n121_ = ~new_n118_ & ~new_n119_;
  assign new_n122_ = ~new_n120_ & ~new_n121_;
  assign new_n123_ = G113gat & G141gat;
  assign new_n124_ = G113gat & ~new_n123_;
  assign new_n125_ = G141gat & ~new_n123_;
  assign new_n126_ = ~new_n124_ & ~new_n125_;
  assign new_n127_ = G169gat & G197gat;
  assign new_n128_ = G169gat & ~new_n127_;
  assign new_n129_ = G197gat & ~new_n127_;
  assign new_n130_ = ~new_n128_ & ~new_n129_;
  assign new_n131_ = ~new_n126_ & ~new_n130_;
  assign new_n132_ = ~new_n126_ & ~new_n131_;
  assign new_n133_ = ~new_n130_ & ~new_n131_;
  assign new_n134_ = ~new_n132_ & ~new_n133_;
  assign new_n135_ = G229gat & G233gat;
  assign new_n136_ = G1gat & G8gat;
  assign new_n137_ = G1gat & ~new_n136_;
  assign new_n138_ = G8gat & ~new_n136_;
  assign new_n139_ = ~new_n137_ & ~new_n138_;
  assign new_n140_ = G15gat & G22gat;
  assign new_n141_ = G15gat & ~new_n140_;
  assign new_n142_ = G22gat & ~new_n140_;
  assign new_n143_ = ~new_n141_ & ~new_n142_;
  assign new_n144_ = ~new_n139_ & ~new_n143_;
  assign new_n145_ = ~new_n139_ & ~new_n144_;
  assign new_n146_ = ~new_n143_ & ~new_n144_;
  assign new_n147_ = ~new_n145_ & ~new_n146_;
  assign new_n148_ = G29gat & G36gat;
  assign new_n149_ = G29gat & ~new_n148_;
  assign new_n150_ = G36gat & ~new_n148_;
  assign new_n151_ = ~new_n149_ & ~new_n150_;
  assign new_n152_ = G43gat & G50gat;
  assign new_n153_ = G43gat & ~new_n152_;
  assign new_n154_ = G50gat & ~new_n152_;
  assign new_n155_ = ~new_n153_ & ~new_n154_;
  assign new_n156_ = ~new_n151_ & ~new_n155_;
  assign new_n157_ = ~new_n151_ & ~new_n156_;
  assign new_n158_ = ~new_n155_ & ~new_n156_;
  assign new_n159_ = ~new_n157_ & ~new_n158_;
  assign new_n160_ = ~new_n147_ & ~new_n159_;
  assign new_n161_ = ~new_n147_ & ~new_n160_;
  assign new_n162_ = ~new_n159_ & ~new_n160_;
  assign new_n163_ = ~new_n161_ & ~new_n162_;
  assign new_n164_ = new_n135_ & ~new_n163_;
  assign new_n165_ = new_n135_ & ~new_n164_;
  assign new_n166_ = ~new_n163_ & ~new_n164_;
  assign new_n167_ = ~new_n165_ & ~new_n166_;
  assign new_n168_ = ~new_n134_ & ~new_n167_;
  assign new_n169_ = ~new_n134_ & ~new_n168_;
  assign new_n170_ = ~new_n167_ & ~new_n168_;
  assign new_n171_ = ~new_n169_ & ~new_n170_;
  assign new_n172_ = G120gat & G148gat;
  assign new_n173_ = G120gat & ~new_n172_;
  assign new_n174_ = G148gat & ~new_n172_;
  assign new_n175_ = ~new_n173_ & ~new_n174_;
  assign new_n176_ = G176gat & G204gat;
  assign new_n177_ = G176gat & ~new_n176_;
  assign new_n178_ = G204gat & ~new_n176_;
  assign new_n179_ = ~new_n177_ & ~new_n178_;
  assign new_n180_ = ~new_n175_ & ~new_n179_;
  assign new_n181_ = ~new_n175_ & ~new_n180_;
  assign new_n182_ = ~new_n179_ & ~new_n180_;
  assign new_n183_ = ~new_n181_ & ~new_n182_;
  assign new_n184_ = G230gat & G233gat;
  assign new_n185_ = G57gat & G64gat;
  assign new_n186_ = G57gat & ~new_n185_;
  assign new_n187_ = G64gat & ~new_n185_;
  assign new_n188_ = ~new_n186_ & ~new_n187_;
  assign new_n189_ = G71gat & G78gat;
  assign new_n190_ = G71gat & ~new_n189_;
  assign new_n191_ = G78gat & ~new_n189_;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign new_n193_ = ~new_n188_ & ~new_n192_;
  assign new_n194_ = ~new_n188_ & ~new_n193_;
  assign new_n195_ = ~new_n192_ & ~new_n193_;
  assign new_n196_ = ~new_n194_ & ~new_n195_;
  assign new_n197_ = G85gat & G92gat;
  assign new_n198_ = G85gat & ~new_n197_;
  assign new_n199_ = G92gat & ~new_n197_;
  assign new_n200_ = ~new_n198_ & ~new_n199_;
  assign new_n201_ = G99gat & G106gat;
  assign new_n202_ = G99gat & ~new_n201_;
  assign new_n203_ = G106gat & ~new_n201_;
  assign new_n204_ = ~new_n202_ & ~new_n203_;
  assign new_n205_ = ~new_n200_ & ~new_n204_;
  assign new_n206_ = ~new_n200_ & ~new_n205_;
  assign new_n207_ = ~new_n204_ & ~new_n205_;
  assign new_n208_ = ~new_n206_ & ~new_n207_;
  assign new_n209_ = ~new_n196_ & ~new_n208_;
  assign new_n210_ = ~new_n196_ & ~new_n209_;
  assign new_n211_ = ~new_n208_ & ~new_n209_;
  assign new_n212_ = ~new_n210_ & ~new_n211_;
  assign new_n213_ = new_n184_ & ~new_n212_;
  assign new_n214_ = new_n184_ & ~new_n213_;
  assign new_n215_ = ~new_n212_ & ~new_n213_;
  assign new_n216_ = ~new_n214_ & ~new_n215_;
  assign new_n217_ = ~new_n183_ & ~new_n216_;
  assign new_n218_ = ~new_n183_ & ~new_n217_;
  assign new_n219_ = ~new_n216_ & ~new_n217_;
  assign new_n220_ = ~new_n218_ & ~new_n219_;
  assign new_n221_ = G127gat & G155gat;
  assign new_n222_ = G127gat & ~new_n221_;
  assign new_n223_ = G155gat & ~new_n221_;
  assign new_n224_ = ~new_n222_ & ~new_n223_;
  assign new_n225_ = G183gat & G211gat;
  assign new_n226_ = G183gat & ~new_n225_;
  assign new_n227_ = G211gat & ~new_n225_;
  assign new_n228_ = ~new_n226_ & ~new_n227_;
  assign new_n229_ = ~new_n224_ & ~new_n228_;
  assign new_n230_ = ~new_n224_ & ~new_n229_;
  assign new_n231_ = ~new_n228_ & ~new_n229_;
  assign new_n232_ = ~new_n230_ & ~new_n231_;
  assign new_n233_ = G231gat & G233gat;
  assign new_n234_ = ~new_n147_ & ~new_n196_;
  assign new_n235_ = ~new_n147_ & ~new_n234_;
  assign new_n236_ = ~new_n196_ & ~new_n234_;
  assign new_n237_ = ~new_n235_ & ~new_n236_;
  assign new_n238_ = new_n233_ & ~new_n237_;
  assign new_n239_ = new_n233_ & ~new_n238_;
  assign new_n240_ = ~new_n237_ & ~new_n238_;
  assign new_n241_ = ~new_n239_ & ~new_n240_;
  assign new_n242_ = ~new_n232_ & ~new_n241_;
  assign new_n243_ = ~new_n232_ & ~new_n242_;
  assign new_n244_ = ~new_n241_ & ~new_n242_;
  assign new_n245_ = ~new_n243_ & ~new_n244_;
  assign new_n246_ = G134gat & G162gat;
  assign new_n247_ = G134gat & ~new_n246_;
  assign new_n248_ = G162gat & ~new_n246_;
  assign new_n249_ = ~new_n247_ & ~new_n248_;
  assign new_n250_ = G190gat & G218gat;
  assign new_n251_ = G190gat & ~new_n250_;
  assign new_n252_ = G218gat & ~new_n250_;
  assign new_n253_ = ~new_n251_ & ~new_n252_;
  assign new_n254_ = ~new_n249_ & ~new_n253_;
  assign new_n255_ = ~new_n249_ & ~new_n254_;
  assign new_n256_ = ~new_n253_ & ~new_n254_;
  assign new_n257_ = ~new_n255_ & ~new_n256_;
  assign new_n258_ = G232gat & G233gat;
  assign new_n259_ = ~new_n159_ & ~new_n208_;
  assign new_n260_ = ~new_n159_ & ~new_n259_;
  assign new_n261_ = ~new_n208_ & ~new_n259_;
  assign new_n262_ = ~new_n260_ & ~new_n261_;
  assign new_n263_ = new_n258_ & ~new_n262_;
  assign new_n264_ = new_n258_ & ~new_n263_;
  assign new_n265_ = ~new_n262_ & ~new_n263_;
  assign new_n266_ = ~new_n264_ & ~new_n265_;
  assign new_n267_ = ~new_n257_ & ~new_n266_;
  assign new_n268_ = ~new_n257_ & ~new_n267_;
  assign new_n269_ = ~new_n266_ & ~new_n267_;
  assign new_n270_ = ~new_n268_ & ~new_n269_;
  assign new_n271_ = G8gat & G36gat;
  assign new_n272_ = G8gat & ~new_n271_;
  assign new_n273_ = G36gat & ~new_n271_;
  assign new_n274_ = ~new_n272_ & ~new_n273_;
  assign new_n275_ = G64gat & G92gat;
  assign new_n276_ = G64gat & ~new_n275_;
  assign new_n277_ = G92gat & ~new_n275_;
  assign new_n278_ = ~new_n276_ & ~new_n277_;
  assign new_n279_ = ~new_n274_ & ~new_n278_;
  assign new_n280_ = ~new_n274_ & ~new_n279_;
  assign new_n281_ = ~new_n278_ & ~new_n279_;
  assign new_n282_ = ~new_n280_ & ~new_n281_;
  assign new_n283_ = G226gat & G233gat;
  assign new_n284_ = G169gat & G176gat;
  assign new_n285_ = G169gat & ~new_n284_;
  assign new_n286_ = G176gat & ~new_n284_;
  assign new_n287_ = ~new_n285_ & ~new_n286_;
  assign new_n288_ = G183gat & G190gat;
  assign new_n289_ = G183gat & ~new_n288_;
  assign new_n290_ = G190gat & ~new_n288_;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = ~new_n287_ & ~new_n291_;
  assign new_n293_ = ~new_n287_ & ~new_n292_;
  assign new_n294_ = ~new_n291_ & ~new_n292_;
  assign new_n295_ = ~new_n293_ & ~new_n294_;
  assign new_n296_ = G197gat & G204gat;
  assign new_n297_ = G197gat & ~new_n296_;
  assign new_n298_ = G204gat & ~new_n296_;
  assign new_n299_ = ~new_n297_ & ~new_n298_;
  assign new_n300_ = G211gat & G218gat;
  assign new_n301_ = G211gat & ~new_n300_;
  assign new_n302_ = G218gat & ~new_n300_;
  assign new_n303_ = ~new_n301_ & ~new_n302_;
  assign new_n304_ = ~new_n299_ & ~new_n303_;
  assign new_n305_ = ~new_n299_ & ~new_n304_;
  assign new_n306_ = ~new_n303_ & ~new_n304_;
  assign new_n307_ = ~new_n305_ & ~new_n306_;
  assign new_n308_ = ~new_n295_ & ~new_n307_;
  assign new_n309_ = ~new_n295_ & ~new_n308_;
  assign new_n310_ = ~new_n307_ & ~new_n308_;
  assign new_n311_ = ~new_n309_ & ~new_n310_;
  assign new_n312_ = new_n283_ & ~new_n311_;
  assign new_n313_ = new_n283_ & ~new_n312_;
  assign new_n314_ = ~new_n311_ & ~new_n312_;
  assign new_n315_ = ~new_n313_ & ~new_n314_;
  assign new_n316_ = ~new_n282_ & ~new_n315_;
  assign new_n317_ = ~new_n282_ & ~new_n316_;
  assign new_n318_ = ~new_n315_ & ~new_n316_;
  assign new_n319_ = ~new_n317_ & ~new_n318_;
  assign new_n320_ = G15gat & G43gat;
  assign new_n321_ = G15gat & ~new_n320_;
  assign new_n322_ = G43gat & ~new_n320_;
  assign new_n323_ = ~new_n321_ & ~new_n322_;
  assign new_n324_ = G71gat & G99gat;
  assign new_n325_ = G71gat & ~new_n324_;
  assign new_n326_ = G99gat & ~new_n324_;
  assign new_n327_ = ~new_n325_ & ~new_n326_;
  assign new_n328_ = ~new_n323_ & ~new_n327_;
  assign new_n329_ = ~new_n323_ & ~new_n328_;
  assign new_n330_ = ~new_n327_ & ~new_n328_;
  assign new_n331_ = ~new_n329_ & ~new_n330_;
  assign new_n332_ = G227gat & G233gat;
  assign new_n333_ = ~new_n98_ & ~new_n295_;
  assign new_n334_ = ~new_n98_ & ~new_n333_;
  assign new_n335_ = ~new_n295_ & ~new_n333_;
  assign new_n336_ = ~new_n334_ & ~new_n335_;
  assign new_n337_ = new_n332_ & ~new_n336_;
  assign new_n338_ = new_n332_ & ~new_n337_;
  assign new_n339_ = ~new_n336_ & ~new_n337_;
  assign new_n340_ = ~new_n338_ & ~new_n339_;
  assign new_n341_ = ~new_n331_ & ~new_n340_;
  assign new_n342_ = ~new_n331_ & ~new_n341_;
  assign new_n343_ = ~new_n340_ & ~new_n341_;
  assign new_n344_ = ~new_n342_ & ~new_n343_;
  assign new_n345_ = G22gat & G50gat;
  assign new_n346_ = G22gat & ~new_n345_;
  assign new_n347_ = G50gat & ~new_n345_;
  assign new_n348_ = ~new_n346_ & ~new_n347_;
  assign new_n349_ = G78gat & G106gat;
  assign new_n350_ = G78gat & ~new_n349_;
  assign new_n351_ = G106gat & ~new_n349_;
  assign new_n352_ = ~new_n350_ & ~new_n351_;
  assign new_n353_ = ~new_n348_ & ~new_n352_;
  assign new_n354_ = ~new_n348_ & ~new_n353_;
  assign new_n355_ = ~new_n352_ & ~new_n353_;
  assign new_n356_ = ~new_n354_ & ~new_n355_;
  assign new_n357_ = G228gat & G233gat;
  assign new_n358_ = ~new_n110_ & ~new_n307_;
  assign new_n359_ = ~new_n110_ & ~new_n358_;
  assign new_n360_ = ~new_n307_ & ~new_n358_;
  assign new_n361_ = ~new_n359_ & ~new_n360_;
  assign new_n362_ = new_n357_ & ~new_n361_;
  assign new_n363_ = new_n357_ & ~new_n362_;
  assign new_n364_ = ~new_n361_ & ~new_n362_;
  assign new_n365_ = ~new_n363_ & ~new_n364_;
  assign new_n366_ = ~new_n356_ & ~new_n365_;
  assign new_n367_ = ~new_n356_ & ~new_n366_;
  assign new_n368_ = ~new_n365_ & ~new_n366_;
  assign new_n369_ = ~new_n367_ & ~new_n368_;
  assign new_n370_ = new_n122_ & new_n319_;
  assign new_n371_ = new_n344_ & new_n370_;
  assign new_n372_ = ~new_n369_ & new_n371_;
  assign new_n373_ = ~new_n344_ & new_n370_;
  assign new_n374_ = new_n369_ & new_n373_;
  assign new_n375_ = new_n122_ & ~new_n319_;
  assign new_n376_ = new_n344_ & new_n375_;
  assign new_n377_ = new_n369_ & new_n376_;
  assign new_n378_ = ~new_n122_ & new_n319_;
  assign new_n379_ = new_n344_ & new_n378_;
  assign new_n380_ = new_n369_ & new_n379_;
  assign new_n381_ = ~new_n377_ & ~new_n380_;
  assign new_n382_ = ~new_n372_ & ~new_n374_;
  assign new_n383_ = new_n381_ & new_n382_;
  assign new_n384_ = ~new_n171_ & new_n220_;
  assign new_n385_ = ~new_n245_ & new_n384_;
  assign new_n386_ = new_n270_ & new_n385_;
  assign new_n387_ = ~new_n383_ & new_n386_;
  assign new_n388_ = ~new_n122_ & new_n387_;
  assign new_n389_ = G1gat & new_n388_;
  assign new_n390_ = G1gat & ~new_n389_;
  assign new_n391_ = new_n388_ & ~new_n389_;
  assign G1324gat = new_n390_ | new_n391_;
  assign new_n393_ = ~new_n319_ & new_n387_;
  assign new_n394_ = G8gat & new_n393_;
  assign new_n395_ = G8gat & ~new_n394_;
  assign new_n396_ = new_n393_ & ~new_n394_;
  assign G1325gat = new_n395_ | new_n396_;
  assign new_n398_ = ~new_n344_ & new_n387_;
  assign new_n399_ = G15gat & new_n398_;
  assign new_n400_ = G15gat & ~new_n399_;
  assign new_n401_ = new_n398_ & ~new_n399_;
  assign G1326gat = new_n400_ | new_n401_;
  assign new_n403_ = ~new_n369_ & new_n387_;
  assign new_n404_ = G22gat & new_n403_;
  assign new_n405_ = G22gat & ~new_n404_;
  assign new_n406_ = new_n403_ & ~new_n404_;
  assign G1327gat = new_n405_ | new_n406_;
  assign new_n408_ = new_n245_ & new_n384_;
  assign new_n409_ = ~new_n270_ & new_n408_;
  assign new_n410_ = ~new_n383_ & new_n409_;
  assign new_n411_ = ~new_n122_ & new_n410_;
  assign new_n412_ = G29gat & new_n411_;
  assign new_n413_ = G29gat & ~new_n412_;
  assign new_n414_ = new_n411_ & ~new_n412_;
  assign G1328gat = new_n413_ | new_n414_;
  assign new_n416_ = ~new_n319_ & new_n410_;
  assign new_n417_ = G36gat & new_n416_;
  assign new_n418_ = G36gat & ~new_n417_;
  assign new_n419_ = new_n416_ & ~new_n417_;
  assign G1329gat = new_n418_ | new_n419_;
  assign new_n421_ = ~new_n344_ & new_n410_;
  assign new_n422_ = G43gat & new_n421_;
  assign new_n423_ = G43gat & ~new_n422_;
  assign new_n424_ = new_n421_ & ~new_n422_;
  assign G1330gat = new_n423_ | new_n424_;
  assign new_n426_ = ~new_n369_ & new_n410_;
  assign new_n427_ = G50gat & new_n426_;
  assign new_n428_ = G50gat & ~new_n427_;
  assign new_n429_ = new_n426_ & ~new_n427_;
  assign G1331gat = new_n428_ | new_n429_;
  assign new_n431_ = new_n171_ & ~new_n220_;
  assign new_n432_ = ~new_n245_ & new_n431_;
  assign new_n433_ = new_n270_ & new_n432_;
  assign new_n434_ = ~new_n383_ & new_n433_;
  assign new_n435_ = ~new_n122_ & new_n434_;
  assign new_n436_ = G57gat & new_n435_;
  assign new_n437_ = G57gat & ~new_n436_;
  assign new_n438_ = new_n435_ & ~new_n436_;
  assign G1332gat = new_n437_ | new_n438_;
  assign new_n440_ = ~new_n319_ & new_n434_;
  assign new_n441_ = G64gat & new_n440_;
  assign new_n442_ = G64gat & ~new_n441_;
  assign new_n443_ = new_n440_ & ~new_n441_;
  assign G1333gat = new_n442_ | new_n443_;
  assign new_n445_ = ~new_n344_ & new_n434_;
  assign new_n446_ = G71gat & new_n445_;
  assign new_n447_ = G71gat & ~new_n446_;
  assign new_n448_ = new_n445_ & ~new_n446_;
  assign G1334gat = new_n447_ | new_n448_;
  assign new_n450_ = ~new_n369_ & new_n434_;
  assign new_n451_ = G78gat & new_n450_;
  assign new_n452_ = G78gat & ~new_n451_;
  assign new_n453_ = new_n450_ & ~new_n451_;
  assign G1335gat = new_n452_ | new_n453_;
  assign new_n455_ = new_n245_ & new_n431_;
  assign new_n456_ = ~new_n270_ & new_n455_;
  assign new_n457_ = ~new_n383_ & new_n456_;
  assign new_n458_ = ~new_n122_ & new_n457_;
  assign new_n459_ = G85gat & new_n458_;
  assign new_n460_ = G85gat & ~new_n459_;
  assign new_n461_ = new_n458_ & ~new_n459_;
  assign G1336gat = new_n460_ | new_n461_;
  assign new_n463_ = ~new_n319_ & new_n457_;
  assign new_n464_ = G92gat & new_n463_;
  assign new_n465_ = G92gat & ~new_n464_;
  assign new_n466_ = new_n463_ & ~new_n464_;
  assign G1337gat = new_n465_ | new_n466_;
  assign new_n468_ = ~new_n344_ & new_n457_;
  assign new_n469_ = G99gat & new_n468_;
  assign new_n470_ = G99gat & ~new_n469_;
  assign new_n471_ = new_n468_ & ~new_n469_;
  assign G1338gat = new_n470_ | new_n471_;
  assign new_n473_ = ~new_n369_ & new_n457_;
  assign new_n474_ = G106gat & new_n473_;
  assign new_n475_ = G106gat & ~new_n474_;
  assign new_n476_ = new_n473_ & ~new_n474_;
  assign G1339gat = new_n475_ | new_n476_;
  assign new_n478_ = new_n171_ & new_n220_;
  assign new_n479_ = new_n245_ & new_n478_;
  assign new_n480_ = ~new_n270_ & new_n479_;
  assign new_n481_ = ~new_n245_ & new_n478_;
  assign new_n482_ = new_n270_ & new_n481_;
  assign new_n483_ = new_n270_ & new_n455_;
  assign new_n484_ = new_n270_ & new_n408_;
  assign new_n485_ = ~new_n483_ & ~new_n484_;
  assign new_n486_ = ~new_n480_ & ~new_n482_;
  assign new_n487_ = new_n485_ & new_n486_;
  assign new_n488_ = ~new_n344_ & new_n378_;
  assign new_n489_ = new_n369_ & new_n488_;
  assign new_n490_ = ~new_n487_ & new_n489_;
  assign new_n491_ = ~new_n171_ & new_n490_;
  assign new_n492_ = G113gat & new_n491_;
  assign new_n493_ = G113gat & ~new_n492_;
  assign new_n494_ = new_n491_ & ~new_n492_;
  assign G1340gat = new_n493_ | new_n494_;
  assign new_n496_ = ~new_n220_ & new_n490_;
  assign new_n497_ = G120gat & new_n496_;
  assign new_n498_ = G120gat & ~new_n497_;
  assign new_n499_ = new_n496_ & ~new_n497_;
  assign G1341gat = new_n498_ | new_n499_;
  assign new_n501_ = ~new_n245_ & new_n490_;
  assign new_n502_ = G127gat & new_n501_;
  assign new_n503_ = G127gat & ~new_n502_;
  assign new_n504_ = new_n501_ & ~new_n502_;
  assign G1342gat = new_n503_ | new_n504_;
  assign new_n506_ = ~new_n270_ & new_n490_;
  assign new_n507_ = G134gat & new_n506_;
  assign new_n508_ = G134gat & ~new_n507_;
  assign new_n509_ = new_n506_ & ~new_n507_;
  assign G1343gat = new_n508_ | new_n509_;
  assign new_n511_ = ~new_n369_ & new_n379_;
  assign new_n512_ = ~new_n487_ & new_n511_;
  assign new_n513_ = ~new_n171_ & new_n512_;
  assign new_n514_ = G141gat & new_n513_;
  assign new_n515_ = G141gat & ~new_n514_;
  assign new_n516_ = new_n513_ & ~new_n514_;
  assign G1344gat = new_n515_ | new_n516_;
  assign new_n518_ = ~new_n220_ & new_n512_;
  assign new_n519_ = G148gat & new_n518_;
  assign new_n520_ = G148gat & ~new_n519_;
  assign new_n521_ = new_n518_ & ~new_n519_;
  assign G1345gat = new_n520_ | new_n521_;
  assign new_n523_ = ~new_n245_ & new_n512_;
  assign new_n524_ = G155gat & new_n523_;
  assign new_n525_ = G155gat & ~new_n524_;
  assign new_n526_ = new_n523_ & ~new_n524_;
  assign G1346gat = new_n525_ | new_n526_;
  assign new_n528_ = ~new_n270_ & new_n512_;
  assign new_n529_ = G162gat & new_n528_;
  assign new_n530_ = G162gat & ~new_n529_;
  assign new_n531_ = new_n528_ & ~new_n529_;
  assign G1347gat = new_n530_ | new_n531_;
  assign new_n533_ = ~new_n344_ & new_n375_;
  assign new_n534_ = new_n369_ & new_n533_;
  assign new_n535_ = ~new_n487_ & new_n534_;
  assign new_n536_ = ~new_n171_ & new_n535_;
  assign new_n537_ = G169gat & new_n536_;
  assign new_n538_ = G169gat & ~new_n537_;
  assign new_n539_ = new_n536_ & ~new_n537_;
  assign G1348gat = new_n538_ | new_n539_;
  assign new_n541_ = ~new_n220_ & new_n535_;
  assign new_n542_ = G176gat & new_n541_;
  assign new_n543_ = G176gat & ~new_n542_;
  assign new_n544_ = new_n541_ & ~new_n542_;
  assign G1349gat = new_n543_ | new_n544_;
  assign new_n546_ = ~new_n245_ & new_n535_;
  assign new_n547_ = G183gat & new_n546_;
  assign new_n548_ = G183gat & ~new_n547_;
  assign new_n549_ = new_n546_ & ~new_n547_;
  assign G1350gat = new_n548_ | new_n549_;
  assign new_n551_ = ~new_n270_ & new_n535_;
  assign new_n552_ = G190gat & new_n551_;
  assign new_n553_ = G190gat & ~new_n552_;
  assign new_n554_ = new_n551_ & ~new_n552_;
  assign G1351gat = new_n553_ | new_n554_;
  assign new_n556_ = ~new_n369_ & new_n376_;
  assign new_n557_ = ~new_n487_ & new_n556_;
  assign new_n558_ = ~new_n171_ & new_n557_;
  assign new_n559_ = G197gat & new_n558_;
  assign new_n560_ = G197gat & ~new_n559_;
  assign new_n561_ = new_n558_ & ~new_n559_;
  assign G1352gat = new_n560_ | new_n561_;
  assign new_n563_ = ~new_n220_ & new_n557_;
  assign new_n564_ = G204gat & new_n563_;
  assign new_n565_ = G204gat & ~new_n564_;
  assign new_n566_ = new_n563_ & ~new_n564_;
  assign G1353gat = new_n565_ | new_n566_;
  assign new_n568_ = ~new_n245_ & new_n557_;
  assign new_n569_ = G211gat & new_n568_;
  assign new_n570_ = G211gat & ~new_n569_;
  assign new_n571_ = new_n568_ & ~new_n569_;
  assign G1354gat = new_n570_ | new_n571_;
  assign new_n573_ = ~new_n270_ & new_n557_;
  assign new_n574_ = G218gat & new_n573_;
  assign new_n575_ = G218gat & ~new_n574_;
  assign new_n576_ = new_n573_ & ~new_n574_;
  assign G1355gat = new_n575_ | new_n576_;
endmodule


