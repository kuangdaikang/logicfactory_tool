// Benchmark "i2c" written by ABC on Mon Sep 11 23:41:42 2023

module i2c ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n462_, new_n463_, new_n464_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n474_, new_n475_, new_n476_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n497_, new_n498_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n512_, new_n513_,
    new_n515_, new_n516_, new_n517_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n538_, new_n539_, new_n540_, new_n541_, new_n543_,
    new_n544_, new_n545_, new_n547_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n871_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n945_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n964_, new_n965_,
    new_n966_, new_n968_, new_n969_, new_n970_, new_n972_, new_n973_,
    new_n974_, new_n976_, new_n977_, new_n978_, new_n980_, new_n982_,
    new_n983_, new_n985_, new_n986_, new_n988_, new_n990_, new_n991_,
    new_n993_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1001_, new_n1002_, new_n1004_, new_n1005_, new_n1007_, new_n1008_,
    new_n1010_, new_n1013_, new_n1014_, new_n1016_, new_n1017_, new_n1018_,
    new_n1020_, new_n1021_, new_n1023_, new_n1024_, new_n1026_, new_n1027_,
    new_n1029_, new_n1031_, new_n1033_, new_n1035_, new_n1037_, new_n1039_,
    new_n1040_, new_n1041_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1050_, new_n1052_, new_n1054_, new_n1056_,
    new_n1058_, new_n1065_, new_n1069_, new_n1072_, new_n1073_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1080_, new_n1081_, new_n1082_,
    new_n1084_, new_n1085_, new_n1087_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1096_, new_n1101_, new_n1103_, new_n1105_;
  INV_X1     g000(.I(pi054), .ZN(new_n291_));
  INV_X1     g001(.I(pi010), .ZN(new_n292_));
  NOR4_X1    g002(.A1(pi004), .A2(pi016), .A3(pi018), .A4(pi019), .ZN(new_n293_));
  NOR2_X1    g003(.A1(pi005), .A2(pi022), .ZN(new_n294_));
  INV_X1     g004(.I(new_n294_), .ZN(new_n295_));
  INV_X1     g005(.I(pi012), .ZN(new_n296_));
  INV_X1     g006(.I(pi017), .ZN(new_n297_));
  NAND2_X1   g007(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NOR4_X1    g008(.A1(new_n295_), .A2(new_n298_), .A3(new_n293_), .A4(pi006), .ZN(new_n299_));
  INV_X1     g009(.I(pi007), .ZN(new_n300_));
  INV_X1     g010(.I(pi008), .ZN(new_n301_));
  INV_X1     g011(.I(pi013), .ZN(new_n302_));
  INV_X1     g012(.I(pi021), .ZN(new_n303_));
  NAND4_X1   g013(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .A4(new_n303_), .ZN(new_n304_));
  NOR3_X1    g014(.A1(new_n304_), .A2(new_n292_), .A3(pi014), .ZN(new_n305_));
  NOR2_X1    g015(.A1(pi009), .A2(pi011), .ZN(new_n306_));
  INV_X1     g016(.I(new_n306_), .ZN(new_n307_));
  NOR4_X1    g017(.A1(new_n305_), .A2(new_n299_), .A3(new_n292_), .A4(new_n307_), .ZN(new_n308_));
  NAND2_X1   g018(.A1(new_n295_), .A2(new_n306_), .ZN(new_n309_));
  NAND2_X1   g019(.A1(new_n307_), .A2(new_n294_), .ZN(new_n310_));
  AOI21_X1   g020(.A1(new_n309_), .A2(new_n310_), .B(pi056), .ZN(new_n311_));
  NOR3_X1    g021(.A1(new_n308_), .A2(new_n291_), .A3(new_n311_), .ZN(new_n312_));
  NOR3_X1    g022(.A1(new_n295_), .A2(pi006), .A3(pi007), .ZN(new_n313_));
  NOR3_X1    g023(.A1(pi008), .A2(pi017), .A3(pi021), .ZN(new_n314_));
  NOR4_X1    g024(.A1(new_n293_), .A2(pi012), .A3(pi013), .A4(pi014), .ZN(new_n315_));
  NAND4_X1   g025(.A1(new_n315_), .A2(new_n313_), .A3(new_n306_), .A4(new_n314_), .ZN(new_n316_));
  AOI21_X1   g026(.A1(new_n316_), .A2(pi054), .B(pi000), .ZN(new_n317_));
  NOR2_X1    g027(.A1(pi003), .A2(pi129), .ZN(new_n318_));
  OAI21_X1   g028(.A1(new_n312_), .A2(new_n317_), .B(new_n318_), .ZN(po015));
  NOR2_X1    g029(.A1(pi010), .A2(pi022), .ZN(new_n320_));
  INV_X1     g030(.I(new_n320_), .ZN(new_n321_));
  NOR2_X1    g031(.A1(pi011), .A2(pi012), .ZN(new_n322_));
  INV_X1     g032(.I(new_n322_), .ZN(new_n323_));
  NOR2_X1    g033(.A1(pi008), .A2(pi021), .ZN(new_n324_));
  INV_X1     g034(.I(new_n324_), .ZN(new_n325_));
  NOR4_X1    g035(.A1(new_n321_), .A2(new_n323_), .A3(new_n325_), .A4(pi014), .ZN(new_n326_));
  NOR2_X1    g036(.A1(pi005), .A2(pi006), .ZN(new_n327_));
  INV_X1     g037(.I(new_n327_), .ZN(new_n328_));
  NOR2_X1    g038(.A1(pi007), .A2(pi013), .ZN(new_n329_));
  INV_X1     g039(.I(new_n329_), .ZN(new_n330_));
  NOR2_X1    g040(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NOR2_X1    g041(.A1(new_n331_), .A2(new_n293_), .ZN(new_n332_));
  NAND2_X1   g042(.A1(new_n332_), .A2(new_n326_), .ZN(new_n333_));
  NOR2_X1    g043(.A1(new_n291_), .A2(pi017), .ZN(new_n334_));
  AOI21_X1   g044(.A1(new_n333_), .A2(new_n334_), .B(pi001), .ZN(new_n335_));
  INV_X1     g045(.I(new_n318_), .ZN(new_n336_));
  NOR3_X1    g046(.A1(new_n321_), .A2(pi014), .A3(new_n291_), .ZN(new_n337_));
  INV_X1     g047(.I(new_n337_), .ZN(new_n338_));
  INV_X1     g048(.I(pi011), .ZN(new_n339_));
  NAND2_X1   g049(.A1(new_n301_), .A2(new_n339_), .ZN(new_n340_));
  NOR3_X1    g050(.A1(new_n340_), .A2(pi017), .A3(pi021), .ZN(new_n341_));
  NOR3_X1    g051(.A1(new_n338_), .A2(new_n293_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1     g052(.I(pi009), .ZN(new_n343_));
  NAND2_X1   g053(.A1(new_n327_), .A2(new_n296_), .ZN(new_n344_));
  NOR2_X1    g054(.A1(new_n344_), .A2(new_n330_), .ZN(new_n345_));
  NAND2_X1   g055(.A1(new_n345_), .A2(new_n343_), .ZN(new_n346_));
  OAI21_X1   g056(.A1(new_n342_), .A2(new_n346_), .B(new_n336_), .ZN(new_n347_));
  NOR2_X1    g057(.A1(new_n347_), .A2(new_n335_), .ZN(po016));
  INV_X1     g058(.I(pi082), .ZN(new_n349_));
  NAND2_X1   g059(.A1(pi122), .A2(pi127), .ZN(new_n350_));
  INV_X1     g060(.I(new_n350_), .ZN(new_n351_));
  NOR2_X1    g061(.A1(new_n351_), .A2(new_n349_), .ZN(new_n352_));
  INV_X1     g062(.I(pi041), .ZN(new_n353_));
  INV_X1     g063(.I(pi046), .ZN(new_n354_));
  INV_X1     g064(.I(pi050), .ZN(new_n355_));
  INV_X1     g065(.I(pi038), .ZN(new_n356_));
  INV_X1     g066(.I(pi040), .ZN(new_n357_));
  NOR2_X1    g067(.A1(pi042), .A2(pi044), .ZN(new_n358_));
  NAND3_X1   g068(.A1(new_n358_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n359_));
  NAND4_X1   g069(.A1(new_n359_), .A2(new_n353_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n360_));
  NOR2_X1    g070(.A1(new_n360_), .A2(pi043), .ZN(new_n361_));
  INV_X1     g071(.I(pi024), .ZN(new_n362_));
  NOR3_X1    g072(.A1(pi015), .A2(pi020), .A3(pi049), .ZN(new_n363_));
  NAND2_X1   g073(.A1(new_n363_), .A2(new_n362_), .ZN(new_n364_));
  INV_X1     g074(.I(pi047), .ZN(new_n365_));
  INV_X1     g075(.I(pi048), .ZN(new_n366_));
  NAND2_X1   g076(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NOR4_X1    g077(.A1(new_n364_), .A2(pi045), .A3(pi082), .A4(new_n367_), .ZN(new_n368_));
  NAND2_X1   g078(.A1(new_n361_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1   g079(.A1(new_n369_), .A2(new_n352_), .ZN(new_n370_));
  INV_X1     g080(.I(new_n352_), .ZN(new_n371_));
  NAND3_X1   g081(.A1(new_n361_), .A2(new_n371_), .A3(new_n368_), .ZN(new_n372_));
  NAND3_X1   g082(.A1(new_n370_), .A2(new_n372_), .A3(pi002), .ZN(new_n373_));
  INV_X1     g083(.I(new_n364_), .ZN(new_n374_));
  NOR2_X1    g084(.A1(pi043), .A2(pi047), .ZN(new_n375_));
  INV_X1     g085(.I(pi002), .ZN(new_n376_));
  INV_X1     g086(.I(pi045), .ZN(new_n377_));
  NAND2_X1   g087(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1     g088(.I(new_n378_), .ZN(new_n379_));
  NAND4_X1   g089(.A1(new_n379_), .A2(new_n366_), .A3(new_n349_), .A4(new_n375_), .ZN(new_n380_));
  NOR2_X1    g090(.A1(pi046), .A2(pi050), .ZN(new_n381_));
  NAND3_X1   g091(.A1(new_n381_), .A2(new_n356_), .A3(new_n353_), .ZN(new_n382_));
  INV_X1     g092(.I(new_n382_), .ZN(new_n383_));
  NOR2_X1    g093(.A1(pi040), .A2(pi042), .ZN(new_n384_));
  INV_X1     g094(.I(new_n384_), .ZN(new_n385_));
  NOR2_X1    g095(.A1(new_n385_), .A2(pi044), .ZN(new_n386_));
  INV_X1     g096(.I(new_n386_), .ZN(new_n387_));
  NOR4_X1    g097(.A1(new_n380_), .A2(new_n374_), .A3(new_n383_), .A4(new_n387_), .ZN(new_n388_));
  NOR3_X1    g098(.A1(new_n388_), .A2(pi065), .A3(new_n351_), .ZN(new_n389_));
  AOI21_X1   g099(.A1(new_n373_), .A2(new_n389_), .B(pi129), .ZN(po017));
  INV_X1     g100(.I(pi113), .ZN(new_n391_));
  INV_X1     g101(.I(pi123), .ZN(new_n392_));
  NAND3_X1   g102(.A1(new_n391_), .A2(new_n392_), .A3(pi000), .ZN(new_n393_));
  NOR2_X1    g103(.A1(pi009), .A2(pi014), .ZN(new_n394_));
  INV_X1     g104(.I(new_n394_), .ZN(new_n395_));
  NOR2_X1    g105(.A1(new_n321_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1   g106(.A1(new_n332_), .A2(new_n314_), .A3(new_n322_), .A4(new_n396_), .ZN(new_n397_));
  NOR2_X1    g107(.A1(pi061), .A2(pi118), .ZN(new_n398_));
  NAND2_X1   g108(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  AOI21_X1   g109(.A1(new_n399_), .A2(new_n393_), .B(pi129), .ZN(po018));
  NOR3_X1    g110(.A1(new_n341_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n401_));
  NOR2_X1    g111(.A1(new_n292_), .A2(pi022), .ZN(new_n402_));
  NAND4_X1   g112(.A1(new_n401_), .A2(new_n345_), .A3(new_n394_), .A4(new_n402_), .ZN(new_n403_));
  NAND2_X1   g113(.A1(new_n291_), .A2(pi004), .ZN(new_n404_));
  AOI21_X1   g114(.A1(new_n403_), .A2(new_n404_), .B(new_n336_), .ZN(po019));
  NAND2_X1   g115(.A1(new_n396_), .A2(new_n302_), .ZN(new_n406_));
  NOR3_X1    g116(.A1(new_n406_), .A2(pi059), .A3(new_n341_), .ZN(new_n407_));
  NOR2_X1    g117(.A1(new_n344_), .A2(pi007), .ZN(new_n408_));
  INV_X1     g118(.I(new_n408_), .ZN(new_n409_));
  NOR2_X1    g119(.A1(pi004), .A2(pi019), .ZN(new_n410_));
  INV_X1     g120(.I(new_n410_), .ZN(new_n411_));
  NOR2_X1    g121(.A1(new_n411_), .A2(pi018), .ZN(new_n412_));
  INV_X1     g122(.I(pi028), .ZN(new_n413_));
  INV_X1     g123(.I(pi016), .ZN(new_n414_));
  NAND2_X1   g124(.A1(new_n414_), .A2(pi054), .ZN(new_n415_));
  NOR4_X1    g125(.A1(new_n415_), .A2(pi025), .A3(new_n413_), .A4(pi029), .ZN(new_n416_));
  NAND4_X1   g126(.A1(new_n407_), .A2(new_n409_), .A3(new_n412_), .A4(new_n416_), .ZN(new_n417_));
  NAND2_X1   g127(.A1(new_n291_), .A2(pi005), .ZN(new_n418_));
  AOI21_X1   g128(.A1(new_n417_), .A2(new_n418_), .B(new_n336_), .ZN(po020));
  INV_X1     g129(.I(new_n412_), .ZN(new_n420_));
  NOR2_X1    g130(.A1(new_n420_), .A2(pi028), .ZN(new_n421_));
  INV_X1     g131(.I(pi025), .ZN(new_n422_));
  NOR4_X1    g132(.A1(new_n408_), .A2(new_n422_), .A3(pi029), .A4(new_n415_), .ZN(new_n423_));
  NAND3_X1   g133(.A1(new_n407_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1   g134(.A1(new_n291_), .A2(pi006), .ZN(new_n425_));
  AOI21_X1   g135(.A1(new_n424_), .A2(new_n425_), .B(new_n336_), .ZN(po021));
  INV_X1     g136(.I(new_n406_), .ZN(new_n427_));
  INV_X1     g137(.I(pi005), .ZN(new_n428_));
  NAND2_X1   g138(.A1(new_n428_), .A2(new_n300_), .ZN(new_n429_));
  NAND2_X1   g139(.A1(new_n297_), .A2(pi008), .ZN(new_n430_));
  NOR4_X1    g140(.A1(new_n429_), .A2(new_n430_), .A3(pi018), .A4(pi021), .ZN(new_n431_));
  NOR2_X1    g141(.A1(new_n323_), .A2(pi006), .ZN(new_n432_));
  NOR2_X1    g142(.A1(new_n411_), .A2(new_n415_), .ZN(new_n433_));
  NAND4_X1   g143(.A1(new_n427_), .A2(new_n431_), .A3(new_n432_), .A4(new_n433_), .ZN(new_n434_));
  NAND2_X1   g144(.A1(new_n291_), .A2(pi007), .ZN(new_n435_));
  AOI21_X1   g145(.A1(new_n434_), .A2(new_n435_), .B(new_n336_), .ZN(po022));
  INV_X1     g146(.I(new_n396_), .ZN(new_n437_));
  NOR3_X1    g147(.A1(new_n437_), .A2(new_n330_), .A3(new_n344_), .ZN(new_n438_));
  NOR4_X1    g148(.A1(new_n340_), .A2(pi017), .A3(pi018), .A4(new_n303_), .ZN(new_n439_));
  NAND3_X1   g149(.A1(new_n438_), .A2(new_n433_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1   g150(.A1(new_n291_), .A2(pi008), .ZN(new_n441_));
  AOI21_X1   g151(.A1(new_n440_), .A2(new_n441_), .B(new_n336_), .ZN(po023));
  NOR4_X1    g152(.A1(new_n321_), .A2(new_n395_), .A3(new_n339_), .A4(pi013), .ZN(new_n443_));
  INV_X1     g153(.I(new_n314_), .ZN(new_n444_));
  NOR2_X1    g154(.A1(new_n444_), .A2(pi018), .ZN(new_n445_));
  INV_X1     g155(.I(new_n445_), .ZN(new_n446_));
  NAND4_X1   g156(.A1(new_n446_), .A2(new_n409_), .A3(new_n433_), .A4(new_n443_), .ZN(new_n447_));
  NAND2_X1   g157(.A1(new_n291_), .A2(pi009), .ZN(new_n448_));
  AOI21_X1   g158(.A1(new_n447_), .A2(new_n448_), .B(new_n336_), .ZN(po024));
  NOR4_X1    g159(.A1(new_n445_), .A2(pi009), .A3(pi010), .A4(pi022), .ZN(new_n450_));
  NOR3_X1    g160(.A1(new_n323_), .A2(new_n429_), .A3(pi006), .ZN(new_n451_));
  INV_X1     g161(.I(pi014), .ZN(new_n452_));
  NOR4_X1    g162(.A1(new_n411_), .A2(new_n415_), .A3(pi013), .A4(new_n452_), .ZN(new_n453_));
  NAND3_X1   g163(.A1(new_n450_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1   g164(.A1(new_n291_), .A2(pi010), .ZN(new_n455_));
  AOI21_X1   g165(.A1(new_n454_), .A2(new_n455_), .B(new_n336_), .ZN(po025));
  NAND3_X1   g166(.A1(new_n292_), .A2(new_n339_), .A3(pi022), .ZN(new_n457_));
  NOR4_X1    g167(.A1(new_n457_), .A2(new_n395_), .A3(new_n411_), .A4(new_n415_), .ZN(new_n458_));
  NAND3_X1   g168(.A1(new_n446_), .A2(new_n345_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1   g169(.A1(new_n291_), .A2(pi011), .ZN(new_n460_));
  AOI21_X1   g170(.A1(new_n459_), .A2(new_n460_), .B(new_n336_), .ZN(po026));
  NOR4_X1    g171(.A1(new_n437_), .A2(new_n331_), .A3(new_n411_), .A4(new_n415_), .ZN(new_n462_));
  NAND4_X1   g172(.A1(new_n462_), .A2(pi018), .A3(new_n314_), .A4(new_n322_), .ZN(new_n463_));
  NAND2_X1   g173(.A1(new_n291_), .A2(pi012), .ZN(new_n464_));
  AOI21_X1   g174(.A1(new_n463_), .A2(new_n464_), .B(new_n336_), .ZN(po027));
  INV_X1     g175(.I(pi029), .ZN(new_n466_));
  NOR3_X1    g176(.A1(new_n466_), .A2(pi025), .A3(pi028), .ZN(new_n467_));
  NOR2_X1    g177(.A1(new_n437_), .A2(new_n420_), .ZN(new_n468_));
  NOR3_X1    g178(.A1(new_n330_), .A2(new_n415_), .A3(pi059), .ZN(new_n469_));
  NOR2_X1    g179(.A1(new_n341_), .A2(new_n344_), .ZN(new_n470_));
  NAND4_X1   g180(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .A4(new_n467_), .ZN(new_n471_));
  NAND2_X1   g181(.A1(new_n291_), .A2(pi013), .ZN(new_n472_));
  AOI21_X1   g182(.A1(new_n471_), .A2(new_n472_), .B(new_n336_), .ZN(po028));
  NOR4_X1    g183(.A1(new_n411_), .A2(pi009), .A3(new_n302_), .A4(pi016), .ZN(new_n474_));
  NAND4_X1   g184(.A1(new_n446_), .A2(new_n337_), .A3(new_n451_), .A4(new_n474_), .ZN(new_n475_));
  NAND2_X1   g185(.A1(new_n291_), .A2(pi014), .ZN(new_n476_));
  AOI21_X1   g186(.A1(new_n475_), .A2(new_n476_), .B(new_n336_), .ZN(po029));
  INV_X1     g187(.I(pi129), .ZN(new_n478_));
  INV_X1     g188(.I(new_n361_), .ZN(new_n479_));
  NOR2_X1    g189(.A1(pi015), .A2(pi045), .ZN(new_n480_));
  INV_X1     g190(.I(new_n480_), .ZN(new_n481_));
  NOR2_X1    g191(.A1(pi024), .A2(pi049), .ZN(new_n482_));
  OAI21_X1   g192(.A1(pi002), .A2(pi020), .B(new_n482_), .ZN(new_n483_));
  NOR4_X1    g193(.A1(new_n479_), .A2(new_n367_), .A3(new_n481_), .A4(new_n483_), .ZN(new_n484_));
  INV_X1     g194(.I(new_n360_), .ZN(new_n485_));
  NAND2_X1   g195(.A1(new_n375_), .A2(new_n366_), .ZN(new_n486_));
  INV_X1     g196(.I(new_n486_), .ZN(new_n487_));
  NAND4_X1   g197(.A1(new_n485_), .A2(new_n480_), .A3(new_n482_), .A4(new_n487_), .ZN(new_n488_));
  INV_X1     g198(.I(new_n367_), .ZN(new_n489_));
  NOR3_X1    g199(.A1(pi038), .A2(pi046), .A3(pi050), .ZN(new_n490_));
  NAND2_X1   g200(.A1(new_n386_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1    g201(.A1(new_n491_), .A2(pi045), .ZN(new_n492_));
  NOR4_X1    g202(.A1(pi015), .A2(pi041), .A3(pi043), .A4(pi082), .ZN(new_n493_));
  NAND4_X1   g203(.A1(new_n492_), .A2(new_n489_), .A3(new_n482_), .A4(new_n493_), .ZN(new_n494_));
  INV_X1     g204(.I(pi015), .ZN(new_n495_));
  NOR3_X1    g205(.A1(new_n351_), .A2(pi070), .A3(new_n349_), .ZN(new_n497_));
  NAND3_X1   g206(.A1(new_n494_), .A2(new_n488_), .A3(new_n497_), .ZN(new_n498_));
  OAI21_X1   g207(.A1(new_n498_), .A2(new_n484_), .B(new_n478_), .ZN(po030));
  INV_X1     g208(.I(pi006), .ZN(new_n500_));
  NOR4_X1    g209(.A1(new_n330_), .A2(pi005), .A3(new_n500_), .A4(pi012), .ZN(new_n501_));
  NAND3_X1   g210(.A1(new_n401_), .A2(new_n396_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1   g211(.A1(new_n291_), .A2(pi016), .ZN(new_n503_));
  AOI21_X1   g212(.A1(new_n502_), .A2(new_n503_), .B(new_n336_), .ZN(po031));
  NOR4_X1    g213(.A1(new_n325_), .A2(new_n328_), .A3(pi011), .A4(pi017), .ZN(new_n505_));
  INV_X1     g214(.I(pi059), .ZN(new_n506_));
  NOR4_X1    g215(.A1(pi007), .A2(pi012), .A3(pi016), .A4(pi025), .ZN(new_n507_));
  NOR4_X1    g216(.A1(new_n507_), .A2(pi029), .A3(new_n291_), .A4(new_n506_), .ZN(new_n508_));
  NAND4_X1   g217(.A1(new_n427_), .A2(new_n421_), .A3(new_n505_), .A4(new_n508_), .ZN(new_n509_));
  NAND2_X1   g218(.A1(new_n291_), .A2(pi017), .ZN(new_n510_));
  AOI21_X1   g219(.A1(new_n509_), .A2(new_n510_), .B(new_n336_), .ZN(po032));
  NOR4_X1    g220(.A1(new_n420_), .A2(new_n414_), .A3(new_n341_), .A4(new_n291_), .ZN(new_n512_));
  AOI22_X1   g221(.A1(new_n512_), .A2(new_n438_), .B1(pi018), .B2(new_n291_), .ZN(new_n513_));
  NOR2_X1    g222(.A1(new_n513_), .A2(new_n336_), .ZN(po033));
  NOR4_X1    g223(.A1(new_n325_), .A2(new_n415_), .A3(pi011), .A4(new_n297_), .ZN(new_n515_));
  NAND3_X1   g224(.A1(new_n438_), .A2(new_n412_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1   g225(.A1(new_n291_), .A2(pi019), .ZN(new_n517_));
  AOI21_X1   g226(.A1(new_n516_), .A2(new_n517_), .B(new_n336_), .ZN(po034));
  NOR2_X1    g227(.A1(pi041), .A2(pi043), .ZN(new_n519_));
  INV_X1     g228(.I(new_n519_), .ZN(new_n520_));
  NOR2_X1    g229(.A1(new_n520_), .A2(pi047), .ZN(new_n521_));
  NAND2_X1   g230(.A1(new_n521_), .A2(new_n354_), .ZN(new_n522_));
  NAND4_X1   g231(.A1(new_n522_), .A2(new_n362_), .A3(new_n377_), .A4(new_n366_), .ZN(new_n523_));
  INV_X1     g232(.I(pi044), .ZN(new_n524_));
  NOR2_X1    g233(.A1(pi038), .A2(pi050), .ZN(new_n525_));
  NAND4_X1   g234(.A1(new_n363_), .A2(new_n384_), .A3(new_n525_), .A4(new_n524_), .ZN(new_n526_));
  NOR2_X1    g235(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  NOR3_X1    g236(.A1(new_n351_), .A2(pi071), .A3(new_n349_), .ZN(new_n530_));
  NAND2_X1   g237(.A1(new_n527_), .A2(pi002), .ZN(new_n531_));
  INV_X1     g238(.I(pi049), .ZN(new_n532_));
  NOR3_X1    g239(.A1(pi038), .A2(pi040), .A3(pi050), .ZN(new_n533_));
  NAND4_X1   g240(.A1(new_n533_), .A2(new_n495_), .A3(new_n358_), .A4(new_n532_), .ZN(new_n534_));
  OAI21_X1   g241(.A1(new_n523_), .A2(new_n534_), .B(pi020), .ZN(new_n535_));
  NAND3_X1   g242(.A1(new_n531_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1   g243(.A1(new_n536_), .A2(new_n478_), .ZN(po035));
  NOR3_X1    g244(.A1(new_n340_), .A2(pi004), .A3(pi016), .ZN(new_n538_));
  NAND3_X1   g245(.A1(new_n303_), .A2(pi019), .A3(pi054), .ZN(new_n539_));
  NOR4_X1    g246(.A1(new_n538_), .A2(pi017), .A3(pi018), .A4(new_n539_), .ZN(new_n540_));
  AOI22_X1   g247(.A1(new_n438_), .A2(new_n540_), .B1(pi021), .B2(new_n291_), .ZN(new_n541_));
  NOR2_X1    g248(.A1(new_n541_), .A2(new_n336_), .ZN(po036));
  NOR4_X1    g249(.A1(new_n428_), .A2(pi007), .A3(pi013), .A4(pi014), .ZN(new_n543_));
  NAND4_X1   g250(.A1(new_n450_), .A2(new_n432_), .A3(new_n433_), .A4(new_n543_), .ZN(new_n544_));
  NAND2_X1   g251(.A1(new_n291_), .A2(pi022), .ZN(new_n545_));
  AOI21_X1   g252(.A1(new_n544_), .A2(new_n545_), .B(new_n336_), .ZN(po037));
  INV_X1     g253(.I(pi023), .ZN(new_n547_));
  NOR4_X1    g254(.A1(new_n547_), .A2(pi055), .A3(pi061), .A4(pi129), .ZN(po038));
  NAND3_X1   g255(.A1(new_n492_), .A2(new_n366_), .A3(new_n521_), .ZN(new_n549_));
  NAND2_X1   g256(.A1(new_n376_), .A2(new_n495_), .ZN(new_n550_));
  NOR3_X1    g257(.A1(new_n550_), .A2(pi020), .A3(pi049), .ZN(new_n551_));
  NAND2_X1   g258(.A1(new_n551_), .A2(new_n352_), .ZN(new_n552_));
  NAND2_X1   g259(.A1(new_n552_), .A2(new_n362_), .ZN(new_n553_));
  AOI21_X1   g260(.A1(new_n549_), .A2(pi082), .B(new_n553_), .ZN(new_n554_));
  INV_X1     g261(.I(new_n363_), .ZN(new_n555_));
  NOR4_X1    g262(.A1(new_n555_), .A2(new_n367_), .A3(new_n378_), .A4(pi082), .ZN(new_n556_));
  NAND2_X1   g263(.A1(new_n350_), .A2(pi063), .ZN(new_n557_));
  AOI21_X1   g264(.A1(new_n361_), .A2(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NAND2_X1   g265(.A1(new_n519_), .A2(new_n354_), .ZN(new_n559_));
  NOR3_X1    g266(.A1(new_n559_), .A2(new_n367_), .A3(pi045), .ZN(new_n560_));
  INV_X1     g267(.I(new_n358_), .ZN(new_n561_));
  INV_X1     g268(.I(new_n533_), .ZN(new_n562_));
  NOR4_X1    g269(.A1(new_n562_), .A2(new_n362_), .A3(new_n561_), .A4(new_n349_), .ZN(new_n563_));
  AOI21_X1   g270(.A1(new_n563_), .A2(new_n560_), .B(pi129), .ZN(new_n564_));
  NOR3_X1    g271(.A1(new_n554_), .A2(new_n558_), .A3(new_n564_), .ZN(po039));
  INV_X1     g272(.I(pi053), .ZN(new_n566_));
  INV_X1     g273(.I(pi085), .ZN(new_n567_));
  INV_X1     g274(.I(pi026), .ZN(new_n568_));
  NOR3_X1    g275(.A1(pi039), .A2(pi051), .A3(pi052), .ZN(new_n569_));
  INV_X1     g276(.I(pi110), .ZN(new_n570_));
  OR2_X2     g277(.A1(pi095), .A2(pi097), .Z(new_n571_));
  OAI21_X1   g278(.A1(new_n571_), .A2(pi100), .B(new_n570_), .ZN(new_n572_));
  AOI22_X1   g279(.A1(new_n572_), .A2(pi025), .B1(pi026), .B2(pi116), .ZN(new_n573_));
  INV_X1     g280(.I(pi116), .ZN(new_n574_));
  NAND2_X1   g281(.A1(new_n574_), .A2(pi025), .ZN(new_n575_));
  OAI22_X1   g282(.A1(new_n573_), .A2(new_n569_), .B1(new_n568_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1     g283(.I(pi096), .ZN(new_n577_));
  NOR2_X1    g284(.A1(new_n567_), .A2(new_n574_), .ZN(new_n578_));
  NAND4_X1   g285(.A1(new_n578_), .A2(new_n567_), .A3(new_n577_), .A4(new_n570_), .ZN(new_n579_));
  NAND2_X1   g286(.A1(new_n579_), .A2(pi100), .ZN(new_n580_));
  NOR2_X1    g287(.A1(new_n575_), .A2(new_n567_), .ZN(new_n581_));
  NOR2_X1    g288(.A1(new_n581_), .A2(pi026), .ZN(new_n582_));
  AOI22_X1   g289(.A1(new_n576_), .A2(new_n567_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1     g290(.I(pi027), .ZN(new_n584_));
  NAND3_X1   g291(.A1(new_n569_), .A2(new_n422_), .A3(pi116), .ZN(new_n585_));
  OAI21_X1   g292(.A1(new_n569_), .A2(new_n574_), .B(pi025), .ZN(new_n586_));
  AOI21_X1   g293(.A1(new_n586_), .A2(new_n585_), .B(new_n584_), .ZN(new_n587_));
  INV_X1     g294(.I(pi100), .ZN(new_n588_));
  NOR2_X1    g295(.A1(pi095), .A2(pi097), .ZN(new_n589_));
  AOI21_X1   g296(.A1(new_n589_), .A2(new_n588_), .B(pi110), .ZN(new_n590_));
  NAND2_X1   g297(.A1(new_n569_), .A2(pi025), .ZN(new_n591_));
  NOR2_X1    g298(.A1(pi026), .A2(pi085), .ZN(new_n592_));
  OAI21_X1   g299(.A1(new_n591_), .A2(new_n590_), .B(new_n592_), .ZN(new_n593_));
  OAI21_X1   g300(.A1(new_n587_), .A2(new_n593_), .B(new_n584_), .ZN(new_n594_));
  OAI21_X1   g301(.A1(new_n583_), .A2(new_n594_), .B(new_n566_), .ZN(new_n595_));
  NOR2_X1    g302(.A1(new_n575_), .A2(pi026), .ZN(new_n596_));
  NOR2_X1    g303(.A1(pi027), .A2(pi085), .ZN(new_n597_));
  INV_X1     g304(.I(new_n597_), .ZN(new_n598_));
  NOR2_X1    g305(.A1(new_n598_), .A2(new_n566_), .ZN(new_n599_));
  AOI21_X1   g306(.A1(new_n599_), .A2(new_n596_), .B(pi058), .ZN(new_n600_));
  INV_X1     g307(.I(pi058), .ZN(new_n601_));
  NOR2_X1    g308(.A1(new_n601_), .A2(pi053), .ZN(new_n602_));
  NAND3_X1   g309(.A1(new_n596_), .A2(new_n602_), .A3(new_n597_), .ZN(new_n603_));
  NAND2_X1   g310(.A1(new_n603_), .A2(new_n336_), .ZN(new_n604_));
  AOI21_X1   g311(.A1(new_n595_), .A2(new_n600_), .B(new_n604_), .ZN(po040));
  NAND3_X1   g312(.A1(new_n569_), .A2(new_n592_), .A3(pi116), .ZN(new_n606_));
  INV_X1     g313(.I(new_n578_), .ZN(new_n607_));
  NAND2_X1   g314(.A1(pi026), .A2(pi116), .ZN(new_n608_));
  NAND2_X1   g315(.A1(new_n574_), .A2(pi085), .ZN(new_n609_));
  NAND4_X1   g316(.A1(new_n609_), .A2(new_n577_), .A3(new_n570_), .A4(new_n608_), .ZN(new_n610_));
  OAI21_X1   g317(.A1(pi026), .A2(new_n607_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1   g318(.A1(new_n611_), .A2(pi100), .ZN(new_n612_));
  NOR3_X1    g319(.A1(pi027), .A2(pi053), .A3(pi058), .ZN(new_n613_));
  NAND2_X1   g320(.A1(new_n613_), .A2(new_n318_), .ZN(new_n614_));
  AOI21_X1   g321(.A1(new_n612_), .A2(new_n606_), .B(new_n614_), .ZN(po041));
  NAND2_X1   g322(.A1(new_n577_), .A2(pi095), .ZN(new_n616_));
  AOI21_X1   g323(.A1(pi027), .A2(pi116), .B(new_n616_), .ZN(new_n617_));
  NAND3_X1   g324(.A1(new_n617_), .A2(new_n570_), .A3(new_n609_), .ZN(new_n618_));
  AOI21_X1   g325(.A1(new_n578_), .A2(new_n584_), .B(pi100), .ZN(new_n619_));
  NAND2_X1   g326(.A1(new_n569_), .A2(pi116), .ZN(new_n620_));
  NOR2_X1    g327(.A1(pi053), .A2(pi058), .ZN(new_n621_));
  INV_X1     g328(.I(new_n621_), .ZN(new_n622_));
  NAND2_X1   g329(.A1(new_n318_), .A2(new_n568_), .ZN(new_n623_));
  OAI22_X1   g330(.A1(new_n620_), .A2(new_n598_), .B1(new_n623_), .B2(new_n622_), .ZN(new_n624_));
  AOI21_X1   g331(.A1(new_n618_), .A2(new_n619_), .B(new_n624_), .ZN(po042));
  INV_X1     g332(.I(new_n569_), .ZN(new_n626_));
  NOR2_X1    g333(.A1(new_n626_), .A2(new_n608_), .ZN(new_n627_));
  NOR4_X1    g334(.A1(new_n616_), .A2(pi026), .A3(pi100), .A4(pi110), .ZN(new_n628_));
  NAND2_X1   g335(.A1(new_n626_), .A2(new_n568_), .ZN(new_n629_));
  NOR3_X1    g336(.A1(new_n629_), .A2(pi027), .A3(new_n574_), .ZN(new_n630_));
  NOR4_X1    g337(.A1(new_n630_), .A2(new_n584_), .A3(new_n627_), .A4(new_n628_), .ZN(new_n631_));
  NOR4_X1    g338(.A1(new_n569_), .A2(pi026), .A3(pi027), .A4(new_n574_), .ZN(new_n632_));
  NAND2_X1   g339(.A1(new_n569_), .A2(new_n584_), .ZN(new_n633_));
  AOI21_X1   g340(.A1(new_n629_), .A2(new_n633_), .B(new_n590_), .ZN(new_n634_));
  XNOR2_X1   g341(.A1(pi026), .A2(pi027), .ZN(new_n635_));
  OAI21_X1   g342(.A1(new_n635_), .A2(pi116), .B(pi028), .ZN(new_n636_));
  NOR4_X1    g343(.A1(new_n631_), .A2(new_n632_), .A3(new_n634_), .A4(new_n636_), .ZN(new_n637_));
  OAI21_X1   g344(.A1(new_n637_), .A2(pi085), .B(new_n566_), .ZN(new_n640_));
  NOR3_X1    g345(.A1(new_n598_), .A2(new_n413_), .A3(pi116), .ZN(new_n641_));
  NOR2_X1    g346(.A1(new_n566_), .A2(pi026), .ZN(new_n642_));
  AOI21_X1   g347(.A1(new_n641_), .A2(new_n642_), .B(pi058), .ZN(new_n643_));
  NAND3_X1   g348(.A1(new_n641_), .A2(new_n568_), .A3(new_n602_), .ZN(new_n644_));
  NAND2_X1   g349(.A1(new_n644_), .A2(new_n336_), .ZN(new_n645_));
  AOI21_X1   g350(.A1(new_n640_), .A2(new_n643_), .B(new_n645_), .ZN(po043));
  NAND2_X1   g351(.A1(new_n574_), .A2(pi029), .ZN(new_n647_));
  INV_X1     g352(.I(new_n647_), .ZN(new_n648_));
  NAND3_X1   g353(.A1(new_n648_), .A2(pi085), .A3(new_n613_), .ZN(new_n649_));
  INV_X1     g354(.I(pi097), .ZN(new_n650_));
  NAND2_X1   g355(.A1(new_n466_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1   g356(.A1(pi096), .A2(pi110), .B(pi097), .ZN(new_n652_));
  AND2_X2    g357(.A1(new_n651_), .A2(new_n652_), .Z(new_n653_));
  NOR2_X1    g358(.A1(pi095), .A2(pi100), .ZN(new_n654_));
  OAI21_X1   g359(.A1(new_n651_), .A2(new_n652_), .B(new_n654_), .ZN(new_n655_));
  AOI21_X1   g360(.A1(pi029), .A2(pi110), .B(new_n601_), .ZN(new_n656_));
  OAI21_X1   g361(.A1(new_n653_), .A2(new_n655_), .B(new_n656_), .ZN(new_n657_));
  NAND2_X1   g362(.A1(new_n466_), .A2(new_n574_), .ZN(new_n658_));
  NAND2_X1   g363(.A1(new_n650_), .A2(pi116), .ZN(new_n659_));
  AOI21_X1   g364(.A1(new_n658_), .A2(new_n659_), .B(new_n601_), .ZN(new_n660_));
  NAND2_X1   g365(.A1(new_n601_), .A2(pi053), .ZN(new_n661_));
  OAI21_X1   g366(.A1(new_n647_), .A2(new_n661_), .B(new_n566_), .ZN(new_n662_));
  NOR2_X1    g367(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  AOI21_X1   g368(.A1(new_n657_), .A2(new_n663_), .B(pi027), .ZN(new_n664_));
  NAND4_X1   g369(.A1(new_n621_), .A2(pi027), .A3(new_n574_), .A4(pi029), .ZN(new_n665_));
  NAND2_X1   g370(.A1(new_n665_), .A2(new_n567_), .ZN(new_n666_));
  OAI21_X1   g371(.A1(new_n664_), .A2(new_n666_), .B(new_n649_), .ZN(new_n667_));
  NOR4_X1    g372(.A1(new_n622_), .A2(new_n568_), .A3(pi027), .A4(pi085), .ZN(new_n668_));
  AOI21_X1   g373(.A1(new_n668_), .A2(new_n648_), .B(pi026), .ZN(new_n669_));
  AOI21_X1   g374(.A1(new_n667_), .A2(new_n669_), .B(new_n336_), .ZN(po044));
  INV_X1     g375(.I(pi106), .ZN(new_n671_));
  INV_X1     g376(.I(pi060), .ZN(new_n672_));
  NAND2_X1   g377(.A1(new_n672_), .A2(pi109), .ZN(new_n673_));
  OAI21_X1   g378(.A1(pi030), .A2(pi109), .B(new_n673_), .ZN(new_n674_));
  NAND3_X1   g379(.A1(new_n674_), .A2(pi088), .A3(new_n671_), .ZN(new_n675_));
  INV_X1     g380(.I(pi088), .ZN(new_n676_));
  OAI21_X1   g381(.A1(new_n674_), .A2(pi106), .B(new_n676_), .ZN(new_n677_));
  NAND3_X1   g382(.A1(new_n677_), .A2(new_n675_), .A3(new_n478_), .ZN(po045));
  INV_X1     g383(.I(pi109), .ZN(new_n679_));
  INV_X1     g384(.I(pi031), .ZN(new_n680_));
  NAND2_X1   g385(.A1(new_n680_), .A2(new_n679_), .ZN(new_n681_));
  OAI21_X1   g386(.A1(pi030), .A2(new_n679_), .B(new_n681_), .ZN(new_n682_));
  NAND3_X1   g387(.A1(new_n682_), .A2(pi089), .A3(new_n671_), .ZN(new_n683_));
  INV_X1     g388(.I(pi089), .ZN(new_n684_));
  OAI21_X1   g389(.A1(new_n682_), .A2(pi106), .B(new_n684_), .ZN(new_n685_));
  NAND3_X1   g390(.A1(new_n685_), .A2(new_n683_), .A3(new_n478_), .ZN(po046));
  NAND2_X1   g391(.A1(new_n680_), .A2(pi109), .ZN(new_n687_));
  OAI21_X1   g392(.A1(pi032), .A2(pi109), .B(new_n687_), .ZN(new_n688_));
  NAND3_X1   g393(.A1(new_n688_), .A2(pi099), .A3(new_n671_), .ZN(new_n689_));
  INV_X1     g394(.I(pi099), .ZN(new_n690_));
  OAI21_X1   g395(.A1(new_n688_), .A2(pi106), .B(new_n690_), .ZN(new_n691_));
  NAND3_X1   g396(.A1(new_n691_), .A2(new_n689_), .A3(new_n478_), .ZN(po047));
  INV_X1     g397(.I(pi033), .ZN(new_n693_));
  NAND2_X1   g398(.A1(new_n693_), .A2(new_n679_), .ZN(new_n694_));
  OAI21_X1   g399(.A1(pi032), .A2(new_n679_), .B(new_n694_), .ZN(new_n695_));
  NAND3_X1   g400(.A1(new_n695_), .A2(pi090), .A3(new_n671_), .ZN(new_n696_));
  INV_X1     g401(.I(pi090), .ZN(new_n697_));
  OAI21_X1   g402(.A1(new_n695_), .A2(pi106), .B(new_n697_), .ZN(new_n698_));
  NAND3_X1   g403(.A1(new_n698_), .A2(new_n696_), .A3(new_n478_), .ZN(po048));
  NAND2_X1   g404(.A1(new_n693_), .A2(pi109), .ZN(new_n700_));
  OAI21_X1   g405(.A1(pi034), .A2(pi109), .B(new_n700_), .ZN(new_n701_));
  NAND3_X1   g406(.A1(new_n701_), .A2(pi091), .A3(new_n671_), .ZN(new_n702_));
  INV_X1     g407(.I(pi091), .ZN(new_n703_));
  OAI21_X1   g408(.A1(new_n701_), .A2(pi106), .B(new_n703_), .ZN(new_n704_));
  NAND3_X1   g409(.A1(new_n704_), .A2(new_n702_), .A3(new_n478_), .ZN(po049));
  INV_X1     g410(.I(pi035), .ZN(new_n706_));
  NAND2_X1   g411(.A1(new_n706_), .A2(new_n679_), .ZN(new_n707_));
  OAI21_X1   g412(.A1(pi034), .A2(new_n679_), .B(new_n707_), .ZN(new_n708_));
  NAND3_X1   g413(.A1(new_n708_), .A2(pi092), .A3(new_n671_), .ZN(new_n709_));
  INV_X1     g414(.I(pi092), .ZN(new_n710_));
  OAI21_X1   g415(.A1(new_n708_), .A2(pi106), .B(new_n710_), .ZN(new_n711_));
  NAND3_X1   g416(.A1(new_n711_), .A2(new_n709_), .A3(new_n478_), .ZN(po050));
  NAND2_X1   g417(.A1(new_n706_), .A2(pi109), .ZN(new_n713_));
  OAI21_X1   g418(.A1(pi036), .A2(pi109), .B(new_n713_), .ZN(new_n714_));
  NAND3_X1   g419(.A1(new_n714_), .A2(pi098), .A3(new_n671_), .ZN(new_n715_));
  INV_X1     g420(.I(pi098), .ZN(new_n716_));
  OAI21_X1   g421(.A1(new_n714_), .A2(pi106), .B(new_n716_), .ZN(new_n717_));
  NAND3_X1   g422(.A1(new_n717_), .A2(new_n715_), .A3(new_n478_), .ZN(po051));
  INV_X1     g423(.I(pi037), .ZN(new_n719_));
  NAND2_X1   g424(.A1(new_n719_), .A2(new_n679_), .ZN(new_n720_));
  OAI21_X1   g425(.A1(pi036), .A2(new_n679_), .B(new_n720_), .ZN(new_n721_));
  NAND3_X1   g426(.A1(new_n721_), .A2(pi093), .A3(new_n671_), .ZN(new_n722_));
  INV_X1     g427(.I(pi093), .ZN(new_n723_));
  OAI21_X1   g428(.A1(new_n721_), .A2(pi106), .B(new_n723_), .ZN(new_n724_));
  NAND3_X1   g429(.A1(new_n724_), .A2(new_n722_), .A3(new_n478_), .ZN(po052));
  NOR2_X1    g430(.A1(new_n374_), .A2(new_n378_), .ZN(new_n726_));
  NOR4_X1    g431(.A1(new_n486_), .A2(pi041), .A3(pi046), .A4(pi050), .ZN(new_n727_));
  NOR2_X1    g432(.A1(new_n351_), .A2(pi082), .ZN(new_n728_));
  AND3_X2    g433(.A1(new_n726_), .A2(new_n727_), .A3(new_n728_), .Z(new_n729_));
  NOR2_X1    g434(.A1(new_n386_), .A2(new_n349_), .ZN(new_n730_));
  OAI21_X1   g435(.A1(new_n729_), .A2(new_n730_), .B(new_n356_), .ZN(new_n731_));
  NOR2_X1    g436(.A1(pi050), .A2(pi074), .ZN(new_n732_));
  INV_X1     g437(.I(new_n522_), .ZN(new_n733_));
  NOR3_X1    g438(.A1(new_n378_), .A2(pi024), .A3(pi048), .ZN(new_n734_));
  NOR2_X1    g439(.A1(new_n734_), .A2(new_n555_), .ZN(new_n735_));
  INV_X1     g440(.I(new_n735_), .ZN(new_n736_));
  NOR2_X1    g441(.A1(new_n736_), .A2(new_n733_), .ZN(new_n737_));
  NAND4_X1   g442(.A1(new_n737_), .A2(new_n386_), .A3(new_n728_), .A4(new_n732_), .ZN(new_n738_));
  NOR2_X1    g443(.A1(new_n349_), .A2(pi044), .ZN(new_n739_));
  NAND3_X1   g444(.A1(new_n739_), .A2(pi038), .A3(new_n384_), .ZN(new_n740_));
  NAND4_X1   g445(.A1(new_n731_), .A2(new_n738_), .A3(new_n478_), .A4(new_n740_), .ZN(po053));
  INV_X1     g446(.I(pi039), .ZN(new_n742_));
  INV_X1     g447(.I(pi051), .ZN(new_n743_));
  INV_X1     g448(.I(pi052), .ZN(new_n744_));
  NAND4_X1   g449(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .A4(pi109), .ZN(new_n745_));
  NAND2_X1   g450(.A1(new_n743_), .A2(new_n744_), .ZN(new_n746_));
  NOR2_X1    g451(.A1(pi039), .A2(pi109), .ZN(new_n747_));
  AOI21_X1   g452(.A1(new_n746_), .A2(new_n747_), .B(pi106), .ZN(new_n748_));
  AOI21_X1   g453(.A1(new_n748_), .A2(new_n745_), .B(pi129), .ZN(po054));
  NAND2_X1   g454(.A1(new_n726_), .A2(new_n487_), .ZN(new_n750_));
  NAND2_X1   g455(.A1(new_n728_), .A2(new_n382_), .ZN(new_n751_));
  OAI22_X1   g456(.A1(new_n750_), .A2(new_n751_), .B1(new_n349_), .B2(new_n358_), .ZN(new_n752_));
  NOR3_X1    g457(.A1(new_n351_), .A2(pi073), .A3(pi082), .ZN(new_n753_));
  NAND4_X1   g458(.A1(new_n522_), .A2(new_n358_), .A3(new_n525_), .A4(new_n753_), .ZN(new_n754_));
  NOR3_X1    g459(.A1(new_n561_), .A2(new_n357_), .A3(new_n349_), .ZN(new_n755_));
  OAI22_X1   g460(.A1(new_n754_), .A2(new_n736_), .B1(pi129), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1   g461(.A1(new_n357_), .A2(new_n752_), .B(new_n756_), .ZN(po055));
  NAND2_X1   g462(.A1(new_n375_), .A2(new_n381_), .ZN(new_n758_));
  NOR3_X1    g463(.A1(new_n351_), .A2(pi076), .A3(pi082), .ZN(new_n759_));
  NAND4_X1   g464(.A1(new_n735_), .A2(new_n359_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n760_));
  NAND2_X1   g465(.A1(new_n533_), .A2(new_n354_), .ZN(new_n761_));
  NOR3_X1    g466(.A1(new_n561_), .A2(new_n353_), .A3(new_n349_), .ZN(new_n762_));
  AOI21_X1   g467(.A1(new_n762_), .A2(new_n761_), .B(pi129), .ZN(new_n763_));
  NAND2_X1   g468(.A1(new_n750_), .A2(new_n352_), .ZN(new_n764_));
  AOI21_X1   g469(.A1(new_n491_), .A2(pi082), .B(pi041), .ZN(new_n765_));
  AOI22_X1   g470(.A1(new_n764_), .A2(new_n765_), .B1(new_n760_), .B2(new_n763_), .ZN(po056));
  NOR3_X1    g471(.A1(new_n736_), .A2(pi047), .A3(new_n520_), .ZN(new_n767_));
  NAND2_X1   g472(.A1(new_n767_), .A2(new_n761_), .ZN(new_n768_));
  INV_X1     g473(.I(pi042), .ZN(new_n769_));
  OAI21_X1   g474(.A1(new_n524_), .A2(new_n349_), .B(new_n769_), .ZN(new_n770_));
  AOI21_X1   g475(.A1(new_n768_), .A2(new_n352_), .B(new_n770_), .ZN(new_n771_));
  INV_X1     g476(.I(pi072), .ZN(new_n772_));
  NAND4_X1   g477(.A1(new_n728_), .A2(new_n524_), .A3(new_n772_), .A4(new_n533_), .ZN(new_n773_));
  NOR3_X1    g478(.A1(new_n736_), .A2(new_n733_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1     g479(.I(new_n739_), .ZN(new_n775_));
  NOR2_X1    g480(.A1(new_n775_), .A2(new_n769_), .ZN(new_n776_));
  NOR4_X1    g481(.A1(new_n771_), .A2(pi129), .A3(new_n774_), .A4(new_n776_), .ZN(po057));
  NOR3_X1    g482(.A1(new_n374_), .A2(new_n367_), .A3(new_n378_), .ZN(new_n778_));
  NOR2_X1    g483(.A1(new_n778_), .A2(new_n371_), .ZN(new_n779_));
  NOR2_X1    g484(.A1(new_n485_), .A2(new_n349_), .ZN(new_n780_));
  AND3_X2    g485(.A1(new_n739_), .A2(pi043), .A3(new_n384_), .Z(new_n781_));
  AOI21_X1   g486(.A1(new_n781_), .A2(new_n382_), .B(pi129), .ZN(new_n782_));
  NOR4_X1    g487(.A1(new_n780_), .A2(new_n779_), .A3(pi043), .A4(new_n782_), .ZN(new_n783_));
  INV_X1     g488(.I(pi077), .ZN(new_n784_));
  NOR2_X1    g489(.A1(pi047), .A2(pi082), .ZN(new_n785_));
  NAND2_X1   g490(.A1(new_n735_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1   g491(.A1(new_n786_), .A2(new_n360_), .B(new_n350_), .ZN(new_n787_));
  NAND2_X1   g492(.A1(new_n787_), .A2(new_n784_), .ZN(new_n788_));
  NOR2_X1    g493(.A1(new_n788_), .A2(new_n783_), .ZN(po058));
  INV_X1     g494(.I(pi067), .ZN(new_n790_));
  INV_X1     g495(.I(new_n525_), .ZN(new_n791_));
  NOR4_X1    g496(.A1(new_n733_), .A2(pi082), .A3(new_n385_), .A4(new_n791_), .ZN(new_n792_));
  AOI22_X1   g497(.A1(new_n792_), .A2(new_n735_), .B1(new_n790_), .B2(new_n350_), .ZN(new_n793_));
  NAND2_X1   g498(.A1(new_n351_), .A2(pi044), .ZN(new_n794_));
  AOI21_X1   g499(.A1(pi044), .A2(pi082), .B(pi129), .ZN(new_n795_));
  OAI21_X1   g500(.A1(new_n793_), .A2(new_n794_), .B(new_n795_), .ZN(po059));
  NOR4_X1    g501(.A1(new_n551_), .A2(pi024), .A3(pi082), .A4(new_n351_), .ZN(new_n797_));
  NOR2_X1    g502(.A1(new_n387_), .A2(new_n791_), .ZN(new_n798_));
  NOR2_X1    g503(.A1(new_n559_), .A2(new_n367_), .ZN(new_n799_));
  AOI21_X1   g504(.A1(new_n798_), .A2(new_n799_), .B(new_n349_), .ZN(new_n800_));
  OAI21_X1   g505(.A1(new_n800_), .A2(new_n797_), .B(new_n377_), .ZN(new_n801_));
  NOR4_X1    g506(.A1(new_n351_), .A2(new_n367_), .A3(pi068), .A4(pi082), .ZN(new_n802_));
  NAND4_X1   g507(.A1(new_n361_), .A2(new_n376_), .A3(new_n364_), .A4(new_n802_), .ZN(new_n803_));
  NOR2_X1    g508(.A1(new_n385_), .A2(pi038), .ZN(new_n804_));
  NAND4_X1   g509(.A1(new_n727_), .A2(pi045), .A3(new_n739_), .A4(new_n804_), .ZN(new_n805_));
  NAND4_X1   g510(.A1(new_n801_), .A2(new_n478_), .A3(new_n803_), .A4(new_n805_), .ZN(po060));
  INV_X1     g511(.I(pi075), .ZN(new_n807_));
  INV_X1     g512(.I(new_n359_), .ZN(new_n808_));
  NOR2_X1    g513(.A1(new_n808_), .A2(pi050), .ZN(new_n809_));
  AOI21_X1   g514(.A1(new_n767_), .A2(new_n809_), .B(new_n349_), .ZN(new_n810_));
  NOR3_X1    g515(.A1(new_n810_), .A2(new_n807_), .A3(new_n351_), .ZN(new_n811_));
  NOR2_X1    g516(.A1(new_n354_), .A2(new_n349_), .ZN(new_n812_));
  AOI21_X1   g517(.A1(new_n809_), .A2(new_n812_), .B(pi129), .ZN(new_n813_));
  NOR2_X1    g518(.A1(new_n767_), .A2(new_n371_), .ZN(new_n814_));
  OAI21_X1   g519(.A1(new_n798_), .A2(new_n349_), .B(new_n354_), .ZN(new_n815_));
  NOR2_X1    g520(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NOR3_X1    g521(.A1(new_n811_), .A2(new_n813_), .A3(new_n816_), .ZN(po061));
  NAND2_X1   g522(.A1(new_n361_), .A2(new_n735_), .ZN(new_n818_));
  AOI21_X1   g523(.A1(new_n818_), .A2(pi082), .B(new_n351_), .ZN(new_n819_));
  NOR2_X1    g524(.A1(new_n361_), .A2(new_n349_), .ZN(new_n820_));
  NOR4_X1    g525(.A1(new_n775_), .A2(new_n365_), .A3(new_n385_), .A4(new_n520_), .ZN(new_n821_));
  AOI21_X1   g526(.A1(new_n821_), .A2(new_n490_), .B(pi129), .ZN(new_n822_));
  NOR2_X1    g527(.A1(new_n735_), .A2(new_n371_), .ZN(new_n823_));
  NOR4_X1    g528(.A1(new_n820_), .A2(pi047), .A3(new_n822_), .A4(new_n823_), .ZN(new_n824_));
  NOR3_X1    g529(.A1(new_n824_), .A2(new_n819_), .A3(pi064), .ZN(po062));
  AOI21_X1   g530(.A1(new_n798_), .A2(new_n522_), .B(new_n349_), .ZN(new_n826_));
  OAI21_X1   g531(.A1(new_n726_), .A2(new_n371_), .B(new_n366_), .ZN(new_n827_));
  NOR2_X1    g532(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1     g533(.I(pi062), .ZN(new_n829_));
  NOR3_X1    g534(.A1(new_n555_), .A2(pi024), .A3(pi045), .ZN(new_n830_));
  NAND4_X1   g535(.A1(new_n830_), .A2(new_n829_), .A3(new_n350_), .A4(new_n785_), .ZN(new_n831_));
  NOR3_X1    g536(.A1(new_n479_), .A2(pi002), .A3(new_n831_), .ZN(new_n832_));
  NOR2_X1    g537(.A1(new_n366_), .A2(pi047), .ZN(new_n833_));
  NAND4_X1   g538(.A1(new_n739_), .A2(new_n833_), .A3(new_n381_), .A4(new_n519_), .ZN(new_n834_));
  NOR3_X1    g539(.A1(new_n834_), .A2(pi038), .A3(new_n385_), .ZN(new_n835_));
  NOR4_X1    g540(.A1(new_n828_), .A2(pi129), .A3(new_n832_), .A4(new_n835_), .ZN(po063));
  NAND3_X1   g541(.A1(new_n522_), .A2(new_n377_), .A3(new_n366_), .ZN(new_n837_));
  OAI21_X1   g542(.A1(new_n550_), .A2(pi020), .B(new_n482_), .ZN(new_n838_));
  NOR4_X1    g543(.A1(new_n837_), .A2(pi050), .A3(new_n808_), .A4(new_n838_), .ZN(new_n839_));
  NAND4_X1   g544(.A1(new_n809_), .A2(new_n349_), .A3(new_n482_), .A4(new_n560_), .ZN(new_n840_));
  NAND4_X1   g545(.A1(new_n560_), .A2(new_n358_), .A3(new_n482_), .A4(new_n533_), .ZN(new_n841_));
  NOR3_X1    g546(.A1(new_n351_), .A2(pi069), .A3(new_n349_), .ZN(new_n843_));
  NAND3_X1   g547(.A1(new_n840_), .A2(new_n841_), .A3(new_n843_), .ZN(new_n844_));
  OAI21_X1   g548(.A1(new_n844_), .A2(new_n839_), .B(new_n478_), .ZN(po064));
  INV_X1     g549(.I(new_n559_), .ZN(new_n846_));
  NAND4_X1   g550(.A1(new_n830_), .A2(new_n376_), .A3(new_n489_), .A4(new_n846_), .ZN(new_n847_));
  OAI21_X1   g551(.A1(new_n359_), .A2(new_n349_), .B(new_n355_), .ZN(new_n848_));
  AOI21_X1   g552(.A1(new_n847_), .A2(new_n352_), .B(new_n848_), .ZN(new_n849_));
  NOR4_X1    g553(.A1(new_n736_), .A2(new_n808_), .A3(new_n733_), .A4(pi082), .ZN(new_n850_));
  NAND2_X1   g554(.A1(new_n350_), .A2(pi066), .ZN(new_n851_));
  NOR2_X1    g555(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1    g556(.A1(new_n775_), .A2(new_n355_), .ZN(new_n853_));
  AOI21_X1   g557(.A1(new_n853_), .A2(new_n804_), .B(pi129), .ZN(new_n854_));
  NOR3_X1    g558(.A1(new_n852_), .A2(new_n849_), .A3(new_n854_), .ZN(po065));
  NAND2_X1   g559(.A1(new_n679_), .A2(pi051), .ZN(new_n856_));
  NOR2_X1    g560(.A1(new_n679_), .A2(pi051), .ZN(new_n857_));
  NOR2_X1    g561(.A1(new_n857_), .A2(pi106), .ZN(new_n858_));
  AOI21_X1   g562(.A1(new_n858_), .A2(new_n856_), .B(pi129), .ZN(po066));
  NOR2_X1    g563(.A1(new_n857_), .A2(new_n744_), .ZN(new_n860_));
  NOR3_X1    g564(.A1(new_n679_), .A2(pi051), .A3(pi052), .ZN(new_n861_));
  NOR4_X1    g565(.A1(new_n860_), .A2(new_n861_), .A3(pi106), .A4(pi129), .ZN(po067));
  NAND2_X1   g566(.A1(pi058), .A2(pi116), .ZN(new_n863_));
  NAND4_X1   g567(.A1(new_n654_), .A2(new_n601_), .A3(new_n577_), .A4(new_n570_), .ZN(new_n864_));
  NAND2_X1   g568(.A1(new_n566_), .A2(pi097), .ZN(new_n865_));
  AOI21_X1   g569(.A1(new_n864_), .A2(new_n863_), .B(new_n865_), .ZN(new_n866_));
  AOI21_X1   g570(.A1(new_n601_), .A2(new_n574_), .B(pi053), .ZN(new_n867_));
  NOR4_X1    g571(.A1(new_n866_), .A2(new_n598_), .A3(new_n623_), .A4(new_n867_), .ZN(po068));
  AOI21_X1   g572(.A1(new_n361_), .A2(new_n778_), .B(new_n349_), .ZN(new_n869_));
  OAI21_X1   g573(.A1(new_n869_), .A2(new_n351_), .B(new_n478_), .ZN(po069));
  INV_X1     g574(.I(pi114), .ZN(new_n871_));
  NAND2_X1   g575(.A1(new_n392_), .A2(new_n478_), .ZN(po129));
  NOR3_X1    g576(.A1(po129), .A2(new_n871_), .A3(pi122), .ZN(po070));
  NAND2_X1   g577(.A1(new_n568_), .A2(pi037), .ZN(new_n874_));
  NOR3_X1    g578(.A1(new_n719_), .A2(pi058), .A3(pi116), .ZN(new_n875_));
  NAND2_X1   g579(.A1(new_n719_), .A2(new_n601_), .ZN(new_n876_));
  AOI21_X1   g580(.A1(new_n876_), .A2(new_n574_), .B(new_n601_), .ZN(new_n877_));
  OAI22_X1   g581(.A1(new_n877_), .A2(new_n875_), .B1(new_n568_), .B2(new_n601_), .ZN(new_n878_));
  NOR2_X1    g582(.A1(new_n568_), .A2(pi058), .ZN(new_n879_));
  NOR2_X1    g583(.A1(new_n601_), .A2(pi026), .ZN(new_n880_));
  INV_X1     g584(.I(pi094), .ZN(new_n881_));
  AOI21_X1   g585(.A1(new_n601_), .A2(new_n574_), .B(new_n881_), .ZN(new_n882_));
  OAI21_X1   g586(.A1(new_n879_), .A2(new_n880_), .B(new_n882_), .ZN(new_n883_));
  NAND2_X1   g587(.A1(new_n878_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1    g588(.A1(new_n874_), .A2(pi058), .ZN(new_n885_));
  AOI21_X1   g589(.A1(new_n884_), .A2(new_n566_), .B(new_n885_), .ZN(new_n886_));
  OAI22_X1   g590(.A1(new_n886_), .A2(pi085), .B1(new_n622_), .B2(new_n874_), .ZN(new_n887_));
  NAND2_X1   g591(.A1(new_n621_), .A2(new_n567_), .ZN(new_n888_));
  OAI21_X1   g592(.A1(new_n888_), .A2(new_n874_), .B(new_n336_), .ZN(new_n889_));
  AOI21_X1   g593(.A1(new_n887_), .A2(new_n584_), .B(new_n889_), .ZN(po071));
  NAND2_X1   g594(.A1(new_n592_), .A2(new_n566_), .ZN(new_n891_));
  NOR2_X1    g595(.A1(new_n891_), .A2(pi116), .ZN(new_n892_));
  OAI21_X1   g596(.A1(pi053), .A2(pi085), .B(pi026), .ZN(new_n893_));
  NAND2_X1   g597(.A1(pi053), .A2(pi085), .ZN(new_n894_));
  NAND3_X1   g598(.A1(new_n893_), .A2(new_n894_), .A3(new_n601_), .ZN(new_n895_));
  OAI21_X1   g599(.A1(new_n892_), .A2(new_n895_), .B(pi057), .ZN(new_n896_));
  NOR3_X1    g600(.A1(new_n891_), .A2(new_n672_), .A3(new_n863_), .ZN(new_n897_));
  NOR2_X1    g601(.A1(new_n897_), .A2(pi027), .ZN(new_n898_));
  NAND2_X1   g602(.A1(new_n601_), .A2(pi057), .ZN(new_n899_));
  OAI21_X1   g603(.A1(new_n891_), .A2(new_n899_), .B(new_n336_), .ZN(new_n900_));
  AOI21_X1   g604(.A1(new_n898_), .A2(new_n896_), .B(new_n900_), .ZN(po072));
  NAND3_X1   g605(.A1(new_n569_), .A2(new_n601_), .A3(pi116), .ZN(new_n902_));
  AND2_X2    g606(.A1(new_n902_), .A2(pi027), .Z(new_n903_));
  OAI21_X1   g607(.A1(new_n601_), .A2(pi116), .B(pi027), .ZN(new_n904_));
  XOR2_X1    g608(.A1(new_n902_), .A2(new_n904_), .Z(new_n905_));
  NAND2_X1   g609(.A1(new_n905_), .A2(new_n568_), .ZN(new_n906_));
  NOR3_X1    g610(.A1(new_n336_), .A2(pi053), .A3(pi085), .ZN(new_n907_));
  OAI21_X1   g611(.A1(new_n906_), .A2(new_n903_), .B(new_n907_), .ZN(new_n908_));
  AOI21_X1   g612(.A1(new_n903_), .A2(new_n906_), .B(new_n908_), .ZN(po073));
  NOR2_X1    g613(.A1(new_n506_), .A2(pi116), .ZN(new_n910_));
  INV_X1     g614(.I(new_n910_), .ZN(new_n911_));
  NOR3_X1    g615(.A1(new_n911_), .A2(new_n567_), .A3(new_n622_), .ZN(new_n912_));
  NAND3_X1   g616(.A1(new_n590_), .A2(pi096), .A3(new_n621_), .ZN(new_n913_));
  NOR2_X1    g617(.A1(pi053), .A2(pi116), .ZN(new_n914_));
  OAI21_X1   g618(.A1(new_n590_), .A2(pi053), .B(new_n574_), .ZN(new_n915_));
  NAND3_X1   g619(.A1(new_n572_), .A2(new_n566_), .A3(pi116), .ZN(new_n916_));
  AOI21_X1   g620(.A1(new_n916_), .A2(new_n915_), .B(pi058), .ZN(new_n917_));
  NOR4_X1    g621(.A1(new_n572_), .A2(pi053), .A3(pi058), .A4(pi116), .ZN(new_n918_));
  NOR2_X1    g622(.A1(new_n918_), .A2(new_n506_), .ZN(new_n919_));
  OAI21_X1   g623(.A1(new_n914_), .A2(new_n917_), .B(new_n919_), .ZN(new_n920_));
  AOI21_X1   g624(.A1(new_n920_), .A2(new_n913_), .B(pi085), .ZN(new_n921_));
  OAI21_X1   g625(.A1(new_n921_), .A2(new_n912_), .B(new_n584_), .ZN(new_n922_));
  NOR4_X1    g626(.A1(new_n911_), .A2(new_n584_), .A3(pi085), .A4(new_n622_), .ZN(new_n923_));
  NOR2_X1    g627(.A1(new_n923_), .A2(pi026), .ZN(new_n924_));
  NAND2_X1   g628(.A1(new_n668_), .A2(new_n910_), .ZN(new_n925_));
  NAND2_X1   g629(.A1(new_n925_), .A2(new_n336_), .ZN(new_n926_));
  AOI21_X1   g630(.A1(new_n922_), .A2(new_n924_), .B(new_n926_), .ZN(po074));
  NOR2_X1    g631(.A1(pi117), .A2(pi122), .ZN(new_n928_));
  MUX2_X1    g632(.I0(new_n392_), .I1(pi060), .S(new_n928_), .Z(po075));
  NOR4_X1    g633(.A1(new_n392_), .A2(pi114), .A3(pi122), .A4(pi129), .ZN(po076));
  INV_X1     g634(.I(pi140), .ZN(new_n931_));
  NAND3_X1   g635(.A1(pi131), .A2(pi132), .A3(pi133), .ZN(new_n932_));
  NOR2_X1    g636(.A1(new_n932_), .A2(pi138), .ZN(new_n933_));
  INV_X1     g637(.I(new_n933_), .ZN(new_n934_));
  NOR2_X1    g638(.A1(new_n934_), .A2(pi137), .ZN(new_n935_));
  NAND3_X1   g639(.A1(new_n935_), .A2(pi136), .A3(new_n931_), .ZN(new_n936_));
  INV_X1     g640(.I(pi137), .ZN(new_n937_));
  INV_X1     g641(.I(pi138), .ZN(new_n938_));
  INV_X1     g642(.I(new_n932_), .ZN(new_n939_));
  NAND4_X1   g643(.A1(new_n939_), .A2(pi136), .A3(new_n937_), .A4(new_n938_), .ZN(new_n940_));
  NAND2_X1   g644(.A1(new_n940_), .A2(pi062), .ZN(new_n941_));
  AOI21_X1   g645(.A1(new_n936_), .A2(new_n941_), .B(pi129), .ZN(po077));
  INV_X1     g646(.I(pi136), .ZN(new_n943_));
  NOR2_X1    g647(.A1(new_n943_), .A2(pi142), .ZN(new_n944_));
  AOI22_X1   g648(.A1(new_n935_), .A2(new_n944_), .B1(pi063), .B2(new_n940_), .ZN(new_n945_));
  NOR2_X1    g649(.A1(new_n945_), .A2(pi129), .ZN(po078));
  NOR2_X1    g650(.A1(new_n943_), .A2(pi139), .ZN(new_n947_));
  AOI22_X1   g651(.A1(new_n935_), .A2(new_n947_), .B1(pi064), .B2(new_n940_), .ZN(new_n948_));
  NOR2_X1    g652(.A1(new_n948_), .A2(pi129), .ZN(po079));
  INV_X1     g653(.I(pi146), .ZN(new_n950_));
  NAND3_X1   g654(.A1(new_n935_), .A2(pi136), .A3(new_n950_), .ZN(new_n951_));
  NAND2_X1   g655(.A1(new_n940_), .A2(pi065), .ZN(new_n952_));
  AOI21_X1   g656(.A1(new_n951_), .A2(new_n952_), .B(pi129), .ZN(po080));
  NOR2_X1    g657(.A1(pi136), .A2(pi137), .ZN(new_n954_));
  INV_X1     g658(.I(new_n954_), .ZN(new_n955_));
  NOR2_X1    g659(.A1(new_n934_), .A2(new_n955_), .ZN(new_n956_));
  OR2_X2     g660(.A1(new_n956_), .A2(pi066), .Z(new_n957_));
  NAND2_X1   g661(.A1(new_n956_), .A2(pi143), .ZN(new_n958_));
  AOI21_X1   g662(.A1(new_n957_), .A2(new_n478_), .B(new_n958_), .ZN(po081));
  INV_X1     g663(.I(new_n956_), .ZN(new_n960_));
  NAND2_X1   g664(.A1(new_n960_), .A2(new_n790_), .ZN(new_n961_));
  NAND2_X1   g665(.A1(new_n956_), .A2(pi139), .ZN(new_n962_));
  AOI21_X1   g666(.A1(new_n961_), .A2(new_n478_), .B(new_n962_), .ZN(po082));
  INV_X1     g667(.I(pi141), .ZN(new_n964_));
  NAND3_X1   g668(.A1(new_n935_), .A2(pi136), .A3(new_n964_), .ZN(new_n965_));
  NAND2_X1   g669(.A1(new_n940_), .A2(pi068), .ZN(new_n966_));
  AOI21_X1   g670(.A1(new_n965_), .A2(new_n966_), .B(pi129), .ZN(po083));
  INV_X1     g671(.I(pi143), .ZN(new_n968_));
  NAND3_X1   g672(.A1(new_n935_), .A2(pi136), .A3(new_n968_), .ZN(new_n969_));
  NAND2_X1   g673(.A1(new_n940_), .A2(pi069), .ZN(new_n970_));
  AOI21_X1   g674(.A1(new_n969_), .A2(new_n970_), .B(pi129), .ZN(po084));
  INV_X1     g675(.I(pi144), .ZN(new_n972_));
  NAND3_X1   g676(.A1(new_n935_), .A2(pi136), .A3(new_n972_), .ZN(new_n973_));
  NAND2_X1   g677(.A1(new_n940_), .A2(pi070), .ZN(new_n974_));
  AOI21_X1   g678(.A1(new_n973_), .A2(new_n974_), .B(pi129), .ZN(po085));
  INV_X1     g679(.I(pi145), .ZN(new_n976_));
  NAND3_X1   g680(.A1(new_n935_), .A2(pi136), .A3(new_n976_), .ZN(new_n977_));
  NAND2_X1   g681(.A1(new_n940_), .A2(pi071), .ZN(new_n978_));
  AOI21_X1   g682(.A1(new_n977_), .A2(new_n978_), .B(pi129), .ZN(po086));
  AOI21_X1   g683(.A1(new_n960_), .A2(new_n772_), .B(pi129), .ZN(new_n980_));
  NOR3_X1    g684(.A1(new_n980_), .A2(new_n931_), .A3(new_n960_), .ZN(po087));
  OR2_X2     g685(.A1(new_n956_), .A2(pi073), .Z(new_n982_));
  NAND2_X1   g686(.A1(new_n956_), .A2(pi141), .ZN(new_n983_));
  AOI21_X1   g687(.A1(new_n982_), .A2(new_n478_), .B(new_n983_), .ZN(po088));
  OR2_X2     g688(.A1(new_n956_), .A2(pi074), .Z(new_n985_));
  NAND2_X1   g689(.A1(new_n956_), .A2(pi142), .ZN(new_n986_));
  AOI21_X1   g690(.A1(new_n985_), .A2(new_n478_), .B(new_n986_), .ZN(po089));
  AOI21_X1   g691(.A1(new_n960_), .A2(new_n807_), .B(pi129), .ZN(new_n988_));
  NOR3_X1    g692(.A1(new_n988_), .A2(new_n972_), .A3(new_n960_), .ZN(po090));
  OR2_X2     g693(.A1(new_n956_), .A2(pi076), .Z(new_n990_));
  NAND2_X1   g694(.A1(new_n956_), .A2(pi145), .ZN(new_n991_));
  AOI21_X1   g695(.A1(new_n990_), .A2(new_n478_), .B(new_n991_), .ZN(po091));
  AOI21_X1   g696(.A1(new_n960_), .A2(new_n784_), .B(pi129), .ZN(new_n993_));
  NOR3_X1    g697(.A1(new_n993_), .A2(new_n950_), .A3(new_n960_), .ZN(po092));
  NOR2_X1    g698(.A1(new_n937_), .A2(pi136), .ZN(new_n995_));
  NAND2_X1   g699(.A1(new_n933_), .A2(new_n995_), .ZN(new_n996_));
  INV_X1     g700(.I(new_n996_), .ZN(new_n997_));
  NOR2_X1    g701(.A1(new_n997_), .A2(pi078), .ZN(new_n998_));
  OAI21_X1   g702(.A1(new_n996_), .A2(pi142), .B(new_n478_), .ZN(new_n999_));
  NOR2_X1    g703(.A1(new_n998_), .A2(new_n999_), .ZN(po093));
  NOR2_X1    g704(.A1(new_n997_), .A2(pi079), .ZN(new_n1001_));
  OAI21_X1   g705(.A1(new_n996_), .A2(pi143), .B(new_n478_), .ZN(new_n1002_));
  NOR2_X1    g706(.A1(new_n1001_), .A2(new_n1002_), .ZN(po094));
  NOR2_X1    g707(.A1(new_n997_), .A2(pi080), .ZN(new_n1004_));
  OAI21_X1   g708(.A1(new_n996_), .A2(pi144), .B(new_n478_), .ZN(new_n1005_));
  NOR2_X1    g709(.A1(new_n1004_), .A2(new_n1005_), .ZN(po095));
  NOR2_X1    g710(.A1(new_n997_), .A2(pi081), .ZN(new_n1007_));
  OAI21_X1   g711(.A1(new_n996_), .A2(pi145), .B(new_n478_), .ZN(new_n1008_));
  NOR2_X1    g712(.A1(new_n1007_), .A2(new_n1008_), .ZN(po096));
  OAI21_X1   g713(.A1(new_n996_), .A2(pi146), .B(new_n478_), .ZN(new_n1010_));
  AOI21_X1   g714(.A1(new_n349_), .A2(new_n996_), .B(new_n1010_), .ZN(po097));
  NOR2_X1    g715(.A1(new_n997_), .A2(pi084), .ZN(new_n1013_));
  OAI21_X1   g716(.A1(new_n996_), .A2(pi141), .B(new_n478_), .ZN(new_n1014_));
  NOR2_X1    g717(.A1(new_n1013_), .A2(new_n1014_), .ZN(po099));
  NAND2_X1   g718(.A1(new_n654_), .A2(new_n650_), .ZN(new_n1016_));
  NAND3_X1   g719(.A1(new_n1016_), .A2(new_n567_), .A3(new_n570_), .ZN(new_n1017_));
  NAND4_X1   g720(.A1(new_n609_), .A2(new_n568_), .A3(new_n613_), .A4(new_n318_), .ZN(new_n1018_));
  AOI21_X1   g721(.A1(new_n1017_), .A2(pi096), .B(new_n1018_), .ZN(po100));
  NOR2_X1    g722(.A1(new_n997_), .A2(pi086), .ZN(new_n1020_));
  OAI21_X1   g723(.A1(new_n996_), .A2(pi139), .B(new_n478_), .ZN(new_n1021_));
  NOR2_X1    g724(.A1(new_n1020_), .A2(new_n1021_), .ZN(po101));
  NOR2_X1    g725(.A1(new_n997_), .A2(pi087), .ZN(new_n1023_));
  OAI21_X1   g726(.A1(new_n996_), .A2(pi140), .B(new_n478_), .ZN(new_n1024_));
  NOR2_X1    g727(.A1(new_n1023_), .A2(new_n1024_), .ZN(po102));
  NAND3_X1   g728(.A1(new_n933_), .A2(pi136), .A3(pi137), .ZN(new_n1026_));
  OAI21_X1   g729(.A1(new_n1026_), .A2(pi139), .B(new_n478_), .ZN(new_n1027_));
  AOI21_X1   g730(.A1(new_n676_), .A2(new_n1026_), .B(new_n1027_), .ZN(po103));
  OAI21_X1   g731(.A1(new_n1026_), .A2(pi140), .B(new_n478_), .ZN(new_n1029_));
  AOI21_X1   g732(.A1(new_n684_), .A2(new_n1026_), .B(new_n1029_), .ZN(po104));
  OAI21_X1   g733(.A1(new_n1026_), .A2(pi142), .B(new_n478_), .ZN(new_n1031_));
  AOI21_X1   g734(.A1(new_n697_), .A2(new_n1026_), .B(new_n1031_), .ZN(po105));
  OAI21_X1   g735(.A1(new_n1026_), .A2(pi143), .B(new_n478_), .ZN(new_n1033_));
  AOI21_X1   g736(.A1(new_n703_), .A2(new_n1026_), .B(new_n1033_), .ZN(po106));
  OAI21_X1   g737(.A1(new_n1026_), .A2(pi144), .B(new_n478_), .ZN(new_n1035_));
  AOI21_X1   g738(.A1(new_n710_), .A2(new_n1026_), .B(new_n1035_), .ZN(po107));
  OAI21_X1   g739(.A1(new_n1026_), .A2(pi146), .B(new_n478_), .ZN(new_n1037_));
  AOI21_X1   g740(.A1(new_n723_), .A2(new_n1026_), .B(new_n1037_), .ZN(po108));
  NOR2_X1    g741(.A1(new_n955_), .A2(new_n349_), .ZN(new_n1039_));
  NAND3_X1   g742(.A1(new_n1039_), .A2(pi138), .A3(new_n939_), .ZN(new_n1040_));
  OAI21_X1   g743(.A1(new_n1040_), .A2(pi142), .B(new_n478_), .ZN(new_n1041_));
  AOI21_X1   g744(.A1(new_n881_), .A2(new_n1040_), .B(new_n1041_), .ZN(po109));
  NAND2_X1   g745(.A1(new_n1039_), .A2(pi138), .ZN(new_n1043_));
  INV_X1     g746(.I(new_n1043_), .ZN(new_n1044_));
  INV_X1     g747(.I(pi003), .ZN(new_n1045_));
  AOI21_X1   g748(.A1(new_n1045_), .A2(new_n570_), .B(new_n939_), .ZN(new_n1046_));
  AOI21_X1   g749(.A1(new_n1044_), .A2(new_n939_), .B(new_n1046_), .ZN(new_n1047_));
  OAI21_X1   g750(.A1(new_n1040_), .A2(new_n968_), .B(new_n478_), .ZN(new_n1048_));
  AOI21_X1   g751(.A1(new_n1047_), .A2(pi095), .B(new_n1048_), .ZN(po110));
  OAI21_X1   g752(.A1(new_n1040_), .A2(new_n950_), .B(new_n478_), .ZN(new_n1050_));
  AOI21_X1   g753(.A1(new_n1047_), .A2(pi096), .B(new_n1050_), .ZN(po111));
  OAI21_X1   g754(.A1(new_n1040_), .A2(new_n976_), .B(new_n478_), .ZN(new_n1052_));
  AOI21_X1   g755(.A1(new_n1047_), .A2(pi097), .B(new_n1052_), .ZN(po112));
  OAI21_X1   g756(.A1(new_n1026_), .A2(pi145), .B(new_n478_), .ZN(new_n1054_));
  AOI21_X1   g757(.A1(new_n716_), .A2(new_n1026_), .B(new_n1054_), .ZN(po113));
  OAI21_X1   g758(.A1(new_n1026_), .A2(pi141), .B(new_n478_), .ZN(new_n1056_));
  AOI21_X1   g759(.A1(new_n690_), .A2(new_n1026_), .B(new_n1056_), .ZN(po114));
  OAI21_X1   g760(.A1(new_n1040_), .A2(new_n972_), .B(new_n478_), .ZN(new_n1058_));
  AOI21_X1   g761(.A1(new_n1047_), .A2(pi100), .B(new_n1058_), .ZN(po115));
  NAND4_X1   g762(.A1(new_n1017_), .A2(new_n568_), .A3(new_n584_), .A4(new_n621_), .ZN(new_n1065_));
  AOI21_X1   g763(.A1(new_n1065_), .A2(new_n607_), .B(new_n336_), .ZN(po121));
  NOR2_X1    g764(.A1(new_n336_), .A2(new_n574_), .ZN(new_n1069_));
  NOR4_X1    g765(.A1(new_n1069_), .A2(new_n568_), .A3(pi027), .A4(new_n569_), .ZN(po124));
  NOR4_X1    g766(.A1(new_n1069_), .A2(new_n566_), .A3(pi058), .A4(pi097), .ZN(po125));
  NOR4_X1    g767(.A1(new_n349_), .A2(new_n938_), .A3(pi136), .A4(pi137), .ZN(new_n1072_));
  AOI22_X1   g768(.A1(new_n1043_), .A2(pi111), .B1(pi139), .B2(new_n1072_), .ZN(new_n1073_));
  NOR3_X1    g769(.A1(new_n1073_), .A2(pi129), .A3(new_n932_), .ZN(po126));
  NOR2_X1    g770(.A1(new_n932_), .A2(pi129), .ZN(new_n1075_));
  NOR2_X1    g771(.A1(new_n1044_), .A2(pi112), .ZN(new_n1076_));
  INV_X1     g772(.I(new_n1072_), .ZN(new_n1077_));
  NOR2_X1    g773(.A1(new_n1077_), .A2(new_n964_), .ZN(new_n1078_));
  NOR3_X1    g774(.A1(new_n1076_), .A2(new_n1075_), .A3(new_n1078_), .ZN(po127));
  NAND2_X1   g775(.A1(new_n291_), .A2(new_n391_), .ZN(new_n1080_));
  OAI21_X1   g776(.A1(pi011), .A2(pi022), .B(pi054), .ZN(new_n1081_));
  OAI21_X1   g777(.A1(new_n1080_), .A2(new_n1081_), .B(new_n318_), .ZN(new_n1082_));
  AOI21_X1   g778(.A1(new_n1080_), .A2(new_n1081_), .B(new_n1082_), .ZN(po128));
  NOR2_X1    g779(.A1(new_n1044_), .A2(pi115), .ZN(new_n1084_));
  NOR2_X1    g780(.A1(new_n1077_), .A2(new_n931_), .ZN(new_n1085_));
  NOR3_X1    g781(.A1(new_n1084_), .A2(new_n1075_), .A3(new_n1085_), .ZN(po130));
  NAND3_X1   g782(.A1(new_n343_), .A2(new_n296_), .A3(pi054), .ZN(new_n1087_));
  NOR4_X1    g783(.A1(new_n1087_), .A2(new_n336_), .A3(pi004), .A4(pi007), .ZN(po131));
  NAND2_X1   g784(.A1(new_n478_), .A2(pi122), .ZN(po132));
  INV_X1     g785(.I(pi118), .ZN(new_n1090_));
  NAND2_X1   g786(.A1(new_n467_), .A2(new_n506_), .ZN(new_n1091_));
  AOI21_X1   g787(.A1(new_n291_), .A2(new_n1090_), .B(new_n1091_), .ZN(new_n1092_));
  AND3_X2    g788(.A1(new_n1091_), .A2(new_n291_), .A3(pi118), .Z(new_n1093_));
  NOR3_X1    g789(.A1(new_n1093_), .A2(pi129), .A3(new_n1092_), .ZN(po133));
  NOR2_X1    g790(.A1(new_n654_), .A2(pi129), .ZN(po134));
  NOR3_X1    g791(.A1(pi003), .A2(pi110), .A3(pi120), .ZN(new_n1096_));
  NOR3_X1    g792(.A1(new_n1096_), .A2(pi111), .A3(pi129), .ZN(po135));
  AND3_X2    g793(.A1(new_n478_), .A2(pi081), .A3(pi120), .Z(po136));
  OR2_X2     g794(.A1(pi129), .A2(pi134), .Z(po137));
  OR2_X2     g795(.A1(pi129), .A2(pi135), .Z(po138));
  INV_X1     g796(.I(pi057), .ZN(new_n1101_));
  NOR2_X1    g797(.A1(new_n1101_), .A2(pi129), .ZN(po139));
  NAND2_X1   g798(.A1(new_n577_), .A2(pi125), .ZN(new_n1103_));
  AOI21_X1   g799(.A1(new_n1103_), .A2(new_n1045_), .B(pi129), .ZN(po140));
  INV_X1     g800(.I(pi126), .ZN(new_n1105_));
  AND3_X2    g801(.A1(new_n1105_), .A2(pi132), .A3(pi133), .Z(po141));
  assign     po012 = 1'b1;
  assign     po098 = 1'b0;
  assign     po116 = 1'b0;
  assign     po117 = 1'b0;
  assign     po118 = 1'b0;
  assign     po119 = 1'b0;
  assign     po120 = 1'b0;
  assign     po122 = 1'b0;
  assign     po123 = 1'b0;
  BUF_X16    g802(.I(pi108), .Z(po000));
  BUF_X16    g803(.I(pi083), .Z(po001));
  BUF_X16    g804(.I(pi104), .Z(po002));
  BUF_X16    g805(.I(pi103), .Z(po003));
  BUF_X16    g806(.I(pi102), .Z(po004));
  BUF_X16    g807(.I(pi105), .Z(po005));
  BUF_X16    g808(.I(pi107), .Z(po006));
  BUF_X16    g809(.I(pi101), .Z(po007));
  BUF_X16    g810(.I(pi126), .Z(po008));
  BUF_X16    g811(.I(pi121), .Z(po009));
  BUF_X16    g812(.I(pi001), .Z(po010));
  BUF_X16    g813(.I(pi000), .Z(po011));
  BUF_X16    g814(.I(pi130), .Z(po013));
  BUF_X16    g815(.I(pi128), .Z(po014));
endmodule


