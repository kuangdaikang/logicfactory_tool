// Benchmark "testing" written by ABC on Fri Feb 25 15:12:53 2022

module 25_14 ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A73  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A73;
  wire new_n27_, new_n28_, new_n29_, new_n30_, new_n31_, new_n32_, new_n33_,
    new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_,
    new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_,
    new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_,
    new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_;
  assign new_n27_ = ~A301 & ~A300;
  assign new_n28_ = A299 & A298;
  assign new_n29_ = new_n27_ & new_n28_;
  assign new_n30_ = A269 & ~A266;
  assign new_n31_ = A265 & ~A202;
  assign new_n32_ = new_n30_ & new_n31_;
  assign new_n33_ = new_n29_ & new_n32_;
  assign new_n34_ = ~A201 & A200;
  assign new_n35_ = A199 & A166;
  assign new_n36_ = new_n34_ & new_n35_;
  assign new_n37_ = A167 & ~A168;
  assign new_n38_ = ~A169 & new_n37_;
  assign new_n39_ = new_n36_ & new_n38_;
  assign new_n40_ = new_n33_ & new_n39_;
  assign new_n41_ = A269 & A266;
  assign new_n42_ = ~A265 & ~A202;
  assign new_n43_ = new_n41_ & new_n42_;
  assign new_n44_ = new_n29_ & new_n43_;
  assign new_n45_ = new_n39_ & new_n44_;
  assign new_n46_ = ~new_n40_ & ~new_n45_;
  assign new_n47_ = A265 & new_n30_;
  assign new_n48_ = new_n29_ & new_n47_;
  assign new_n49_ = ~A202 & ~A201;
  assign new_n50_ = A200 & A199;
  assign new_n51_ = new_n49_ & new_n50_;
  assign new_n52_ = ~A168 & ~A169;
  assign new_n53_ = ~A170 & new_n52_;
  assign new_n54_ = new_n51_ & new_n53_;
  assign new_n55_ = new_n48_ & new_n54_;
  assign new_n56_ = ~A265 & new_n41_;
  assign new_n57_ = new_n29_ & new_n56_;
  assign new_n58_ = new_n54_ & new_n57_;
  assign new_n59_ = ~new_n55_ & ~new_n58_;
  assign new_n60_ = new_n46_ & new_n59_;
  assign new_n61_ = ~A202 & ~A200;
  assign new_n62_ = ~A199 & A166;
  assign new_n63_ = new_n61_ & new_n62_;
  assign new_n64_ = new_n38_ & new_n63_;
  assign new_n65_ = new_n48_ & new_n64_;
  assign new_n66_ = new_n57_ & new_n64_;
  assign new_n67_ = ~new_n65_ & ~new_n66_;
  assign new_n68_ = A302 & A299;
  assign new_n69_ = ~A298 & ~A268;
  assign new_n70_ = new_n68_ & new_n69_;
  assign new_n71_ = ~A267 & A266;
  assign new_n72_ = A265 & new_n71_;
  assign new_n73_ = new_n70_ & new_n72_;
  assign new_n74_ = A203 & ~A200;
  assign new_n75_ = new_n35_ & new_n74_;
  assign new_n76_ = new_n38_ & new_n75_;
  assign new_n77_ = new_n73_ & new_n76_;
  assign new_n78_ = A302 & ~A299;
  assign new_n79_ = A298 & ~A268;
  assign new_n80_ = new_n78_ & new_n79_;
  assign new_n81_ = new_n72_ & new_n80_;
  assign new_n82_ = new_n76_ & new_n81_;
  assign new_n83_ = ~new_n77_ & ~new_n82_;
  assign new_n84_ = new_n67_ & new_n83_;
  assign new_n85_ = new_n60_ & new_n84_;
  assign new_n86_ = A203 & A200;
  assign new_n87_ = new_n62_ & new_n86_;
  assign new_n88_ = new_n38_ & new_n87_;
  assign new_n89_ = new_n73_ & new_n88_;
  assign new_n90_ = new_n81_ & new_n88_;
  assign new_n91_ = ~new_n89_ & ~new_n90_;
  assign new_n92_ = ~A301 & ~A299;
  assign new_n93_ = ~A298 & A269;
  assign new_n94_ = new_n92_ & new_n93_;
  assign new_n95_ = ~A266 & A265;
  assign new_n96_ = ~A202 & new_n95_;
  assign new_n97_ = new_n94_ & new_n96_;
  assign new_n98_ = new_n39_ & new_n97_;
  assign new_n99_ = ~A302 & ~A301;
  assign new_n100_ = ~A300 & A269;
  assign new_n101_ = new_n99_ & new_n100_;
  assign new_n102_ = new_n96_ & new_n101_;
  assign new_n103_ = new_n39_ & new_n102_;
  assign new_n104_ = ~new_n98_ & ~new_n103_;
  assign new_n105_ = new_n91_ & new_n104_;
  assign new_n106_ = A266 & ~A265;
  assign new_n107_ = ~A202 & new_n106_;
  assign new_n108_ = new_n94_ & new_n107_;
  assign new_n109_ = new_n39_ & new_n108_;
  assign new_n110_ = new_n101_ & new_n107_;
  assign new_n111_ = new_n39_ & new_n110_;
  assign new_n112_ = ~new_n109_ & ~new_n111_;
  assign new_n113_ = A267 & A266;
  assign new_n114_ = ~A202 & new_n113_;
  assign new_n115_ = new_n29_ & new_n114_;
  assign new_n116_ = new_n39_ & new_n115_;
  assign new_n117_ = A267 & A265;
  assign new_n118_ = ~A202 & new_n117_;
  assign new_n119_ = new_n29_ & new_n118_;
  assign new_n120_ = new_n39_ & new_n119_;
  assign new_n121_ = ~new_n116_ & ~new_n120_;
  assign new_n122_ = new_n112_ & new_n121_;
  assign new_n123_ = new_n105_ & new_n122_;
  assign new_n124_ = new_n85_ & new_n123_;
  assign new_n125_ = ~A203 & ~A202;
  assign new_n126_ = ~A201 & A166;
  assign new_n127_ = new_n125_ & new_n126_;
  assign new_n128_ = new_n38_ & new_n127_;
  assign new_n129_ = new_n48_ & new_n128_;
  assign new_n130_ = new_n57_ & new_n128_;
  assign new_n131_ = ~new_n129_ & ~new_n130_;
  assign new_n132_ = ~A166 & ~A167;
  assign new_n133_ = ~A169 & new_n132_;
  assign new_n134_ = new_n51_ & new_n133_;
  assign new_n135_ = new_n48_ & new_n134_;
  assign new_n136_ = new_n57_ & new_n134_;
  assign new_n137_ = ~new_n135_ & ~new_n136_;
  assign new_n138_ = new_n131_ & new_n137_;
  assign new_n139_ = A166 & ~A167;
  assign new_n140_ = A170 & new_n139_;
  assign new_n141_ = new_n51_ & new_n140_;
  assign new_n142_ = new_n73_ & new_n141_;
  assign new_n143_ = new_n81_ & new_n141_;
  assign new_n144_ = ~new_n142_ & ~new_n143_;
  assign new_n145_ = ~A166 & A167;
  assign new_n146_ = A170 & new_n145_;
  assign new_n147_ = new_n51_ & new_n146_;
  assign new_n148_ = new_n73_ & new_n147_;
  assign new_n149_ = new_n81_ & new_n147_;
  assign new_n150_ = ~new_n148_ & ~new_n149_;
  assign new_n151_ = new_n144_ & new_n150_;
  assign new_n152_ = new_n138_ & new_n151_;
  assign new_n153_ = ~A199 & new_n61_;
  assign new_n154_ = new_n53_ & new_n153_;
  assign new_n155_ = new_n48_ & new_n154_;
  assign new_n156_ = new_n57_ & new_n154_;
  assign new_n157_ = ~new_n155_ & ~new_n156_;
  assign new_n158_ = A199 & new_n74_;
  assign new_n159_ = new_n53_ & new_n158_;
  assign new_n160_ = new_n73_ & new_n159_;
  assign new_n161_ = new_n81_ & new_n159_;
  assign new_n162_ = ~new_n160_ & ~new_n161_;
  assign new_n163_ = new_n157_ & new_n162_;
  assign new_n164_ = ~A199 & new_n86_;
  assign new_n165_ = new_n53_ & new_n164_;
  assign new_n166_ = new_n73_ & new_n165_;
  assign new_n167_ = new_n81_ & new_n165_;
  assign new_n168_ = ~new_n166_ & ~new_n167_;
  assign new_n169_ = A199 & new_n34_;
  assign new_n170_ = new_n53_ & new_n169_;
  assign new_n171_ = new_n97_ & new_n170_;
  assign new_n172_ = new_n102_ & new_n170_;
  assign new_n173_ = ~new_n171_ & ~new_n172_;
  assign new_n174_ = new_n168_ & new_n173_;
  assign new_n175_ = new_n163_ & new_n174_;
  assign new_n176_ = new_n152_ & new_n175_;
  assign new_n177_ = new_n124_ & new_n176_;
  assign new_n178_ = new_n108_ & new_n170_;
  assign new_n179_ = new_n110_ & new_n170_;
  assign new_n180_ = ~new_n178_ & ~new_n179_;
  assign new_n181_ = new_n115_ & new_n170_;
  assign new_n182_ = new_n119_ & new_n170_;
  assign new_n183_ = ~new_n181_ & ~new_n182_;
  assign new_n184_ = new_n180_ & new_n183_;
  assign new_n185_ = ~A201 & new_n125_;
  assign new_n186_ = new_n53_ & new_n185_;
  assign new_n187_ = new_n48_ & new_n186_;
  assign new_n188_ = new_n57_ & new_n186_;
  assign new_n189_ = ~new_n187_ & ~new_n188_;
  assign new_n190_ = ~A200 & ~A199;
  assign new_n191_ = A166 & new_n190_;
  assign new_n192_ = new_n38_ & new_n191_;
  assign new_n193_ = new_n97_ & new_n192_;
  assign new_n194_ = new_n102_ & new_n192_;
  assign new_n195_ = ~new_n193_ & ~new_n194_;
  assign new_n196_ = new_n189_ & new_n195_;
  assign new_n197_ = new_n184_ & new_n196_;
  assign new_n198_ = new_n108_ & new_n192_;
  assign new_n199_ = new_n110_ & new_n192_;
  assign new_n200_ = ~new_n198_ & ~new_n199_;
  assign new_n201_ = new_n115_ & new_n192_;
  assign new_n202_ = new_n119_ & new_n192_;
  assign new_n203_ = ~new_n201_ & ~new_n202_;
  assign new_n204_ = new_n200_ & new_n203_;
  assign new_n205_ = ~A266 & ~A265;
  assign new_n206_ = A203 & new_n205_;
  assign new_n207_ = new_n70_ & new_n206_;
  assign new_n208_ = ~A200 & A199;
  assign new_n209_ = A166 & new_n208_;
  assign new_n210_ = new_n38_ & new_n209_;
  assign new_n211_ = new_n207_ & new_n210_;
  assign new_n212_ = new_n80_ & new_n206_;
  assign new_n213_ = new_n210_ & new_n212_;
  assign new_n214_ = ~new_n211_ & ~new_n213_;
  assign new_n215_ = A300 & A298;
  assign new_n216_ = ~A268 & ~A267;
  assign new_n217_ = new_n215_ & new_n216_;
  assign new_n218_ = A266 & A265;
  assign new_n219_ = A203 & new_n218_;
  assign new_n220_ = new_n217_ & new_n219_;
  assign new_n221_ = new_n210_ & new_n220_;
  assign new_n222_ = A300 & A299;
  assign new_n223_ = new_n216_ & new_n222_;
  assign new_n224_ = new_n219_ & new_n223_;
  assign new_n225_ = new_n210_ & new_n224_;
  assign new_n226_ = ~new_n221_ & ~new_n225_;
  assign new_n227_ = new_n214_ & new_n226_;
  assign new_n228_ = new_n204_ & new_n227_;
  assign new_n229_ = new_n197_ & new_n228_;
  assign new_n230_ = ~A298 & ~A269;
  assign new_n231_ = new_n68_ & new_n230_;
  assign new_n232_ = A203 & new_n216_;
  assign new_n233_ = new_n231_ & new_n232_;
  assign new_n234_ = new_n210_ & new_n233_;
  assign new_n235_ = A298 & ~A269;
  assign new_n236_ = new_n78_ & new_n235_;
  assign new_n237_ = new_n232_ & new_n236_;
  assign new_n238_ = new_n210_ & new_n237_;
  assign new_n239_ = ~new_n234_ & ~new_n238_;
  assign new_n240_ = A200 & ~A199;
  assign new_n241_ = A166 & new_n240_;
  assign new_n242_ = new_n38_ & new_n241_;
  assign new_n243_ = new_n207_ & new_n242_;
  assign new_n244_ = new_n212_ & new_n242_;
  assign new_n245_ = ~new_n243_ & ~new_n244_;
  assign new_n246_ = new_n239_ & new_n245_;
  assign new_n247_ = new_n220_ & new_n242_;
  assign new_n248_ = new_n224_ & new_n242_;
  assign new_n249_ = ~new_n247_ & ~new_n248_;
  assign new_n250_ = new_n233_ & new_n242_;
  assign new_n251_ = new_n237_ & new_n242_;
  assign new_n252_ = ~new_n250_ & ~new_n251_;
  assign new_n253_ = new_n249_ & new_n252_;
  assign new_n254_ = new_n246_ & new_n253_;
  assign new_n255_ = ~A298 & A267;
  assign new_n256_ = new_n92_ & new_n255_;
  assign new_n257_ = A266 & ~A202;
  assign new_n258_ = ~A201 & new_n257_;
  assign new_n259_ = new_n256_ & new_n258_;
  assign new_n260_ = A166 & new_n50_;
  assign new_n261_ = new_n38_ & new_n260_;
  assign new_n262_ = new_n259_ & new_n261_;
  assign new_n263_ = ~A300 & A267;
  assign new_n264_ = new_n99_ & new_n263_;
  assign new_n265_ = new_n258_ & new_n264_;
  assign new_n266_ = new_n261_ & new_n265_;
  assign new_n267_ = ~new_n262_ & ~new_n266_;
  assign new_n268_ = ~A201 & new_n31_;
  assign new_n269_ = new_n256_ & new_n268_;
  assign new_n270_ = new_n261_ & new_n269_;
  assign new_n271_ = new_n264_ & new_n268_;
  assign new_n272_ = new_n261_ & new_n271_;
  assign new_n273_ = ~new_n270_ & ~new_n272_;
  assign new_n274_ = new_n267_ & new_n273_;
  assign new_n275_ = A268 & ~A202;
  assign new_n276_ = ~A201 & new_n275_;
  assign new_n277_ = new_n29_ & new_n276_;
  assign new_n278_ = new_n261_ & new_n277_;
  assign new_n279_ = A201 & A200;
  assign new_n280_ = A166 & new_n279_;
  assign new_n281_ = new_n38_ & new_n280_;
  assign new_n282_ = new_n73_ & new_n281_;
  assign new_n283_ = ~new_n278_ & ~new_n282_;
  assign new_n284_ = new_n81_ & new_n281_;
  assign new_n285_ = A201 & A199;
  assign new_n286_ = A166 & new_n285_;
  assign new_n287_ = new_n38_ & new_n286_;
  assign new_n288_ = new_n73_ & new_n287_;
  assign new_n289_ = ~new_n284_ & ~new_n288_;
  assign new_n290_ = new_n283_ & new_n289_;
  assign new_n291_ = new_n274_ & new_n290_;
  assign new_n292_ = new_n254_ & new_n291_;
  assign new_n293_ = new_n229_ & new_n292_;
  assign new_n294_ = new_n177_ & new_n293_;
  assign new_n295_ = new_n81_ & new_n287_;
  assign new_n296_ = ~A203 & new_n95_;
  assign new_n297_ = new_n94_ & new_n296_;
  assign new_n298_ = A166 & new_n49_;
  assign new_n299_ = new_n38_ & new_n298_;
  assign new_n300_ = new_n297_ & new_n299_;
  assign new_n301_ = ~new_n295_ & ~new_n300_;
  assign new_n302_ = new_n101_ & new_n296_;
  assign new_n303_ = new_n299_ & new_n302_;
  assign new_n304_ = ~A203 & new_n106_;
  assign new_n305_ = new_n94_ & new_n304_;
  assign new_n306_ = new_n299_ & new_n305_;
  assign new_n307_ = ~new_n303_ & ~new_n306_;
  assign new_n308_ = new_n301_ & new_n307_;
  assign new_n309_ = new_n101_ & new_n304_;
  assign new_n310_ = new_n299_ & new_n309_;
  assign new_n311_ = ~A203 & new_n113_;
  assign new_n312_ = new_n29_ & new_n311_;
  assign new_n313_ = new_n299_ & new_n312_;
  assign new_n314_ = ~new_n310_ & ~new_n313_;
  assign new_n315_ = ~A203 & new_n117_;
  assign new_n316_ = new_n29_ & new_n315_;
  assign new_n317_ = new_n299_ & new_n316_;
  assign new_n318_ = new_n133_ & new_n153_;
  assign new_n319_ = new_n48_ & new_n318_;
  assign new_n320_ = ~new_n317_ & ~new_n319_;
  assign new_n321_ = new_n314_ & new_n320_;
  assign new_n322_ = new_n308_ & new_n321_;
  assign new_n323_ = new_n57_ & new_n318_;
  assign new_n324_ = new_n133_ & new_n158_;
  assign new_n325_ = new_n73_ & new_n324_;
  assign new_n326_ = ~new_n323_ & ~new_n325_;
  assign new_n327_ = new_n81_ & new_n324_;
  assign new_n328_ = new_n133_ & new_n164_;
  assign new_n329_ = new_n73_ & new_n328_;
  assign new_n330_ = ~new_n327_ & ~new_n329_;
  assign new_n331_ = new_n326_ & new_n330_;
  assign new_n332_ = new_n81_ & new_n328_;
  assign new_n333_ = new_n133_ & new_n169_;
  assign new_n334_ = new_n97_ & new_n333_;
  assign new_n335_ = ~new_n332_ & ~new_n334_;
  assign new_n336_ = new_n102_ & new_n333_;
  assign new_n337_ = new_n108_ & new_n333_;
  assign new_n338_ = ~new_n336_ & ~new_n337_;
  assign new_n339_ = new_n335_ & new_n338_;
  assign new_n340_ = new_n331_ & new_n339_;
  assign new_n341_ = new_n322_ & new_n340_;
  assign new_n342_ = new_n110_ & new_n333_;
  assign new_n343_ = new_n115_ & new_n333_;
  assign new_n344_ = ~new_n342_ & ~new_n343_;
  assign new_n345_ = new_n119_ & new_n333_;
  assign new_n346_ = new_n133_ & new_n185_;
  assign new_n347_ = new_n48_ & new_n346_;
  assign new_n348_ = ~new_n345_ & ~new_n347_;
  assign new_n349_ = new_n344_ & new_n348_;
  assign new_n350_ = new_n57_ & new_n346_;
  assign new_n351_ = new_n140_ & new_n153_;
  assign new_n352_ = new_n73_ & new_n351_;
  assign new_n353_ = ~new_n350_ & ~new_n352_;
  assign new_n354_ = new_n81_ & new_n351_;
  assign new_n355_ = new_n140_ & new_n158_;
  assign new_n356_ = new_n48_ & new_n355_;
  assign new_n357_ = ~new_n354_ & ~new_n356_;
  assign new_n358_ = new_n353_ & new_n357_;
  assign new_n359_ = new_n349_ & new_n358_;
  assign new_n360_ = new_n57_ & new_n355_;
  assign new_n361_ = new_n140_ & new_n164_;
  assign new_n362_ = new_n48_ & new_n361_;
  assign new_n363_ = ~new_n360_ & ~new_n362_;
  assign new_n364_ = new_n57_ & new_n361_;
  assign new_n365_ = ~A202 & new_n205_;
  assign new_n366_ = new_n70_ & new_n365_;
  assign new_n367_ = new_n140_ & new_n169_;
  assign new_n368_ = new_n366_ & new_n367_;
  assign new_n369_ = ~new_n364_ & ~new_n368_;
  assign new_n370_ = new_n363_ & new_n369_;
  assign new_n371_ = new_n80_ & new_n365_;
  assign new_n372_ = new_n367_ & new_n371_;
  assign new_n373_ = ~A202 & new_n218_;
  assign new_n374_ = new_n217_ & new_n373_;
  assign new_n375_ = new_n367_ & new_n374_;
  assign new_n376_ = ~new_n372_ & ~new_n375_;
  assign new_n377_ = new_n223_ & new_n373_;
  assign new_n378_ = new_n367_ & new_n377_;
  assign new_n379_ = ~A202 & new_n216_;
  assign new_n380_ = new_n231_ & new_n379_;
  assign new_n381_ = new_n367_ & new_n380_;
  assign new_n382_ = ~new_n378_ & ~new_n381_;
  assign new_n383_ = new_n376_ & new_n382_;
  assign new_n384_ = new_n370_ & new_n383_;
  assign new_n385_ = new_n359_ & new_n384_;
  assign new_n386_ = new_n341_ & new_n385_;
  assign new_n387_ = new_n236_ & new_n379_;
  assign new_n388_ = new_n367_ & new_n387_;
  assign new_n389_ = new_n140_ & new_n185_;
  assign new_n390_ = new_n73_ & new_n389_;
  assign new_n391_ = ~new_n388_ & ~new_n390_;
  assign new_n392_ = new_n81_ & new_n389_;
  assign new_n393_ = new_n146_ & new_n153_;
  assign new_n394_ = new_n73_ & new_n393_;
  assign new_n395_ = ~new_n392_ & ~new_n394_;
  assign new_n396_ = new_n391_ & new_n395_;
  assign new_n397_ = new_n81_ & new_n393_;
  assign new_n398_ = new_n146_ & new_n158_;
  assign new_n399_ = new_n48_ & new_n398_;
  assign new_n400_ = ~new_n397_ & ~new_n399_;
  assign new_n401_ = new_n57_ & new_n398_;
  assign new_n402_ = new_n146_ & new_n164_;
  assign new_n403_ = new_n48_ & new_n402_;
  assign new_n404_ = ~new_n401_ & ~new_n403_;
  assign new_n405_ = new_n400_ & new_n404_;
  assign new_n406_ = new_n396_ & new_n405_;
  assign new_n407_ = new_n57_ & new_n402_;
  assign new_n408_ = new_n146_ & new_n169_;
  assign new_n409_ = new_n366_ & new_n408_;
  assign new_n410_ = ~new_n407_ & ~new_n409_;
  assign new_n411_ = new_n371_ & new_n408_;
  assign new_n412_ = new_n374_ & new_n408_;
  assign new_n413_ = ~new_n411_ & ~new_n412_;
  assign new_n414_ = new_n410_ & new_n413_;
  assign new_n415_ = new_n377_ & new_n408_;
  assign new_n416_ = new_n380_ & new_n408_;
  assign new_n417_ = ~new_n415_ & ~new_n416_;
  assign new_n418_ = new_n387_ & new_n408_;
  assign new_n419_ = new_n146_ & new_n185_;
  assign new_n420_ = new_n73_ & new_n419_;
  assign new_n421_ = ~new_n418_ & ~new_n420_;
  assign new_n422_ = new_n417_ & new_n421_;
  assign new_n423_ = new_n414_ & new_n422_;
  assign new_n424_ = new_n406_ & new_n423_;
  assign new_n425_ = new_n81_ & new_n419_;
  assign new_n426_ = A200 & new_n49_;
  assign new_n427_ = A199 & A167;
  assign new_n428_ = A168 & new_n427_;
  assign new_n429_ = new_n426_ & new_n428_;
  assign new_n430_ = new_n73_ & new_n429_;
  assign new_n431_ = ~new_n425_ & ~new_n430_;
  assign new_n432_ = new_n81_ & new_n429_;
  assign new_n433_ = A168 & new_n35_;
  assign new_n434_ = new_n426_ & new_n433_;
  assign new_n435_ = new_n73_ & new_n434_;
  assign new_n436_ = ~new_n432_ & ~new_n435_;
  assign new_n437_ = new_n431_ & new_n436_;
  assign new_n438_ = new_n81_ & new_n434_;
  assign new_n439_ = ~A298 & new_n92_;
  assign new_n440_ = new_n47_ & new_n439_;
  assign new_n441_ = new_n154_ & new_n440_;
  assign new_n442_ = ~new_n438_ & ~new_n441_;
  assign new_n443_ = ~A300 & new_n99_;
  assign new_n444_ = new_n47_ & new_n443_;
  assign new_n445_ = new_n154_ & new_n444_;
  assign new_n446_ = new_n56_ & new_n439_;
  assign new_n447_ = new_n154_ & new_n446_;
  assign new_n448_ = ~new_n445_ & ~new_n447_;
  assign new_n449_ = new_n442_ & new_n448_;
  assign new_n450_ = new_n437_ & new_n449_;
  assign new_n451_ = new_n56_ & new_n443_;
  assign new_n452_ = new_n154_ & new_n451_;
  assign new_n453_ = A299 & new_n27_;
  assign new_n454_ = A298 & A267;
  assign new_n455_ = A266 & new_n454_;
  assign new_n456_ = new_n453_ & new_n455_;
  assign new_n457_ = new_n154_ & new_n456_;
  assign new_n458_ = ~new_n452_ & ~new_n457_;
  assign new_n459_ = A265 & new_n454_;
  assign new_n460_ = new_n453_ & new_n459_;
  assign new_n461_ = new_n154_ & new_n460_;
  assign new_n462_ = ~A298 & new_n68_;
  assign new_n463_ = ~A268 & ~A266;
  assign new_n464_ = ~A265 & new_n463_;
  assign new_n465_ = new_n462_ & new_n464_;
  assign new_n466_ = new_n159_ & new_n465_;
  assign new_n467_ = ~new_n461_ & ~new_n466_;
  assign new_n468_ = new_n458_ & new_n467_;
  assign new_n469_ = ~A268 & new_n222_;
  assign new_n470_ = new_n72_ & new_n469_;
  assign new_n471_ = new_n159_ & new_n470_;
  assign new_n472_ = A298 & new_n78_;
  assign new_n473_ = new_n464_ & new_n472_;
  assign new_n474_ = new_n159_ & new_n473_;
  assign new_n475_ = ~A268 & new_n215_;
  assign new_n476_ = new_n72_ & new_n475_;
  assign new_n477_ = new_n159_ & new_n476_;
  assign new_n478_ = ~new_n474_ & ~new_n477_;
  assign new_n479_ = ~new_n471_ & new_n478_;
  assign new_n480_ = new_n468_ & new_n479_;
  assign new_n481_ = new_n450_ & new_n480_;
  assign new_n482_ = new_n424_ & new_n481_;
  assign new_n483_ = new_n386_ & new_n482_;
  assign new_n484_ = new_n294_ & new_n483_;
  assign new_n485_ = ~A269 & ~A268;
  assign new_n486_ = ~A267 & new_n485_;
  assign new_n487_ = new_n462_ & new_n486_;
  assign new_n488_ = new_n159_ & new_n487_;
  assign new_n489_ = new_n472_ & new_n486_;
  assign new_n490_ = new_n159_ & new_n489_;
  assign new_n491_ = ~new_n488_ & ~new_n490_;
  assign new_n492_ = new_n165_ & new_n465_;
  assign new_n493_ = new_n165_ & new_n473_;
  assign new_n494_ = ~new_n492_ & ~new_n493_;
  assign new_n495_ = new_n491_ & new_n494_;
  assign new_n496_ = new_n165_ & new_n476_;
  assign new_n497_ = new_n165_ & new_n470_;
  assign new_n498_ = ~new_n496_ & ~new_n497_;
  assign new_n499_ = new_n165_ & new_n487_;
  assign new_n500_ = new_n165_ & new_n489_;
  assign new_n501_ = ~new_n499_ & ~new_n500_;
  assign new_n502_ = new_n498_ & new_n501_;
  assign new_n503_ = new_n495_ & new_n502_;
  assign new_n504_ = new_n114_ & new_n439_;
  assign new_n505_ = new_n170_ & new_n504_;
  assign new_n506_ = new_n114_ & new_n443_;
  assign new_n507_ = new_n170_ & new_n506_;
  assign new_n508_ = ~new_n505_ & ~new_n507_;
  assign new_n509_ = new_n118_ & new_n439_;
  assign new_n510_ = new_n170_ & new_n509_;
  assign new_n511_ = new_n118_ & new_n443_;
  assign new_n512_ = new_n170_ & new_n511_;
  assign new_n513_ = ~new_n510_ & ~new_n512_;
  assign new_n514_ = new_n508_ & new_n513_;
  assign new_n515_ = A298 & A268;
  assign new_n516_ = ~A202 & new_n515_;
  assign new_n517_ = new_n453_ & new_n516_;
  assign new_n518_ = new_n170_ & new_n517_;
  assign new_n519_ = A266 & new_n216_;
  assign new_n520_ = new_n462_ & new_n519_;
  assign new_n521_ = A265 & A201;
  assign new_n522_ = A200 & new_n521_;
  assign new_n523_ = new_n53_ & new_n522_;
  assign new_n524_ = new_n520_ & new_n523_;
  assign new_n525_ = ~new_n518_ & ~new_n524_;
  assign new_n526_ = new_n472_ & new_n519_;
  assign new_n527_ = new_n523_ & new_n526_;
  assign new_n528_ = A199 & new_n521_;
  assign new_n529_ = new_n53_ & new_n528_;
  assign new_n530_ = new_n520_ & new_n529_;
  assign new_n531_ = ~new_n527_ & ~new_n530_;
  assign new_n532_ = new_n525_ & new_n531_;
  assign new_n533_ = new_n514_ & new_n532_;
  assign new_n534_ = new_n503_ & new_n533_;
  assign new_n535_ = new_n526_ & new_n529_;
  assign new_n536_ = new_n186_ & new_n440_;
  assign new_n537_ = ~new_n535_ & ~new_n536_;
  assign new_n538_ = new_n186_ & new_n444_;
  assign new_n539_ = new_n186_ & new_n446_;
  assign new_n540_ = ~new_n538_ & ~new_n539_;
  assign new_n541_ = new_n537_ & new_n540_;
  assign new_n542_ = new_n186_ & new_n451_;
  assign new_n543_ = new_n186_ & new_n456_;
  assign new_n544_ = ~new_n542_ & ~new_n543_;
  assign new_n545_ = new_n186_ & new_n460_;
  assign new_n546_ = new_n192_ & new_n504_;
  assign new_n547_ = ~new_n545_ & ~new_n546_;
  assign new_n548_ = new_n544_ & new_n547_;
  assign new_n549_ = new_n541_ & new_n548_;
  assign new_n550_ = new_n192_ & new_n506_;
  assign new_n551_ = new_n192_ & new_n509_;
  assign new_n552_ = ~new_n550_ & ~new_n551_;
  assign new_n553_ = new_n192_ & new_n511_;
  assign new_n554_ = new_n192_ & new_n517_;
  assign new_n555_ = ~new_n553_ & ~new_n554_;
  assign new_n556_ = new_n552_ & new_n555_;
  assign new_n557_ = new_n206_ & new_n475_;
  assign new_n558_ = new_n210_ & new_n557_;
  assign new_n559_ = new_n206_ & new_n469_;
  assign new_n560_ = new_n210_ & new_n559_;
  assign new_n561_ = ~new_n558_ & ~new_n560_;
  assign new_n562_ = A301 & ~A268;
  assign new_n563_ = ~A267 & new_n562_;
  assign new_n564_ = new_n219_ & new_n563_;
  assign new_n565_ = new_n210_ & new_n564_;
  assign new_n566_ = ~A269 & new_n215_;
  assign new_n567_ = new_n232_ & new_n566_;
  assign new_n568_ = new_n210_ & new_n567_;
  assign new_n569_ = ~new_n565_ & ~new_n568_;
  assign new_n570_ = new_n561_ & new_n569_;
  assign new_n571_ = new_n556_ & new_n570_;
  assign new_n572_ = new_n549_ & new_n571_;
  assign new_n573_ = new_n534_ & new_n572_;
  assign new_n574_ = ~A269 & new_n222_;
  assign new_n575_ = new_n232_ & new_n574_;
  assign new_n576_ = new_n210_ & new_n575_;
  assign new_n577_ = new_n242_ & new_n557_;
  assign new_n578_ = ~new_n576_ & ~new_n577_;
  assign new_n579_ = new_n242_ & new_n559_;
  assign new_n580_ = new_n242_ & new_n564_;
  assign new_n581_ = ~new_n579_ & ~new_n580_;
  assign new_n582_ = new_n578_ & new_n581_;
  assign new_n583_ = new_n242_ & new_n567_;
  assign new_n584_ = new_n242_ & new_n575_;
  assign new_n585_ = ~new_n583_ & ~new_n584_;
  assign new_n586_ = new_n276_ & new_n439_;
  assign new_n587_ = new_n261_ & new_n586_;
  assign new_n588_ = new_n276_ & new_n443_;
  assign new_n589_ = new_n261_ & new_n588_;
  assign new_n590_ = ~new_n587_ & ~new_n589_;
  assign new_n591_ = new_n585_ & new_n590_;
  assign new_n592_ = new_n582_ & new_n591_;
  assign new_n593_ = new_n281_ & new_n465_;
  assign new_n594_ = new_n281_ & new_n473_;
  assign new_n595_ = ~new_n593_ & ~new_n594_;
  assign new_n596_ = new_n281_ & new_n476_;
  assign new_n597_ = new_n281_ & new_n470_;
  assign new_n598_ = ~new_n596_ & ~new_n597_;
  assign new_n599_ = new_n595_ & new_n598_;
  assign new_n600_ = new_n281_ & new_n487_;
  assign new_n601_ = new_n281_ & new_n489_;
  assign new_n602_ = ~new_n600_ & ~new_n601_;
  assign new_n603_ = new_n287_ & new_n465_;
  assign new_n604_ = new_n287_ & new_n473_;
  assign new_n605_ = ~new_n603_ & ~new_n604_;
  assign new_n606_ = new_n602_ & new_n605_;
  assign new_n607_ = new_n599_ & new_n606_;
  assign new_n608_ = new_n592_ & new_n607_;
  assign new_n609_ = new_n287_ & new_n476_;
  assign new_n610_ = new_n287_ & new_n470_;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign new_n612_ = new_n287_ & new_n487_;
  assign new_n613_ = new_n287_ & new_n489_;
  assign new_n614_ = ~new_n612_ & ~new_n613_;
  assign new_n615_ = new_n611_ & new_n614_;
  assign new_n616_ = new_n311_ & new_n439_;
  assign new_n617_ = new_n299_ & new_n616_;
  assign new_n618_ = new_n311_ & new_n443_;
  assign new_n619_ = new_n299_ & new_n618_;
  assign new_n620_ = ~new_n617_ & ~new_n619_;
  assign new_n621_ = new_n315_ & new_n439_;
  assign new_n622_ = new_n299_ & new_n621_;
  assign new_n623_ = new_n315_ & new_n443_;
  assign new_n624_ = new_n299_ & new_n623_;
  assign new_n625_ = ~new_n622_ & ~new_n624_;
  assign new_n626_ = new_n620_ & new_n625_;
  assign new_n627_ = new_n615_ & new_n626_;
  assign new_n628_ = ~A203 & new_n515_;
  assign new_n629_ = new_n453_ & new_n628_;
  assign new_n630_ = new_n299_ & new_n629_;
  assign new_n631_ = A265 & A202;
  assign new_n632_ = A166 & new_n631_;
  assign new_n633_ = new_n38_ & new_n632_;
  assign new_n634_ = new_n520_ & new_n633_;
  assign new_n635_ = ~new_n630_ & ~new_n634_;
  assign new_n636_ = new_n526_ & new_n633_;
  assign new_n637_ = new_n318_ & new_n440_;
  assign new_n638_ = ~new_n636_ & ~new_n637_;
  assign new_n639_ = new_n635_ & new_n638_;
  assign new_n640_ = new_n318_ & new_n451_;
  assign new_n641_ = new_n318_ & new_n444_;
  assign new_n642_ = new_n318_ & new_n446_;
  assign new_n643_ = ~new_n641_ & ~new_n642_;
  assign new_n644_ = ~new_n640_ & new_n643_;
  assign new_n645_ = new_n639_ & new_n644_;
  assign new_n646_ = new_n627_ & new_n645_;
  assign new_n647_ = new_n608_ & new_n646_;
  assign new_n648_ = new_n573_ & new_n647_;
  assign new_n649_ = new_n318_ & new_n456_;
  assign new_n650_ = new_n318_ & new_n460_;
  assign new_n651_ = ~new_n649_ & ~new_n650_;
  assign new_n652_ = new_n324_ & new_n465_;
  assign new_n653_ = new_n324_ & new_n473_;
  assign new_n654_ = ~new_n652_ & ~new_n653_;
  assign new_n655_ = new_n651_ & new_n654_;
  assign new_n656_ = new_n324_ & new_n476_;
  assign new_n657_ = new_n324_ & new_n470_;
  assign new_n658_ = ~new_n656_ & ~new_n657_;
  assign new_n659_ = new_n324_ & new_n487_;
  assign new_n660_ = new_n324_ & new_n489_;
  assign new_n661_ = ~new_n659_ & ~new_n660_;
  assign new_n662_ = new_n658_ & new_n661_;
  assign new_n663_ = new_n655_ & new_n662_;
  assign new_n664_ = new_n328_ & new_n465_;
  assign new_n665_ = new_n328_ & new_n473_;
  assign new_n666_ = ~new_n664_ & ~new_n665_;
  assign new_n667_ = new_n328_ & new_n476_;
  assign new_n668_ = new_n328_ & new_n470_;
  assign new_n669_ = ~new_n667_ & ~new_n668_;
  assign new_n670_ = new_n666_ & new_n669_;
  assign new_n671_ = new_n328_ & new_n487_;
  assign new_n672_ = new_n328_ & new_n489_;
  assign new_n673_ = ~new_n671_ & ~new_n672_;
  assign new_n674_ = new_n333_ & new_n504_;
  assign new_n675_ = new_n333_ & new_n506_;
  assign new_n676_ = ~new_n674_ & ~new_n675_;
  assign new_n677_ = new_n673_ & new_n676_;
  assign new_n678_ = new_n670_ & new_n677_;
  assign new_n679_ = new_n663_ & new_n678_;
  assign new_n680_ = new_n333_ & new_n509_;
  assign new_n681_ = new_n333_ & new_n511_;
  assign new_n682_ = ~new_n680_ & ~new_n681_;
  assign new_n683_ = new_n333_ & new_n517_;
  assign new_n684_ = new_n133_ & new_n522_;
  assign new_n685_ = new_n520_ & new_n684_;
  assign new_n686_ = ~new_n683_ & ~new_n685_;
  assign new_n687_ = new_n682_ & new_n686_;
  assign new_n688_ = new_n526_ & new_n684_;
  assign new_n689_ = new_n133_ & new_n528_;
  assign new_n690_ = new_n520_ & new_n689_;
  assign new_n691_ = ~new_n688_ & ~new_n690_;
  assign new_n692_ = new_n526_ & new_n689_;
  assign new_n693_ = new_n346_ & new_n440_;
  assign new_n694_ = ~new_n692_ & ~new_n693_;
  assign new_n695_ = new_n691_ & new_n694_;
  assign new_n696_ = new_n687_ & new_n695_;
  assign new_n697_ = new_n346_ & new_n444_;
  assign new_n698_ = new_n346_ & new_n446_;
  assign new_n699_ = ~new_n697_ & ~new_n698_;
  assign new_n700_ = new_n346_ & new_n451_;
  assign new_n701_ = new_n346_ & new_n456_;
  assign new_n702_ = ~new_n700_ & ~new_n701_;
  assign new_n703_ = new_n699_ & new_n702_;
  assign new_n704_ = new_n346_ & new_n460_;
  assign new_n705_ = A169 & new_n50_;
  assign new_n706_ = new_n268_ & new_n705_;
  assign new_n707_ = new_n520_ & new_n706_;
  assign new_n708_ = ~new_n704_ & ~new_n707_;
  assign new_n709_ = new_n526_ & new_n706_;
  assign new_n710_ = new_n351_ & new_n465_;
  assign new_n711_ = ~new_n709_ & ~new_n710_;
  assign new_n712_ = new_n708_ & new_n711_;
  assign new_n713_ = new_n703_ & new_n712_;
  assign new_n714_ = new_n696_ & new_n713_;
  assign new_n715_ = new_n679_ & new_n714_;
  assign new_n716_ = new_n351_ & new_n473_;
  assign new_n717_ = new_n351_ & new_n476_;
  assign new_n718_ = ~new_n716_ & ~new_n717_;
  assign new_n719_ = new_n351_ & new_n470_;
  assign new_n720_ = new_n351_ & new_n487_;
  assign new_n721_ = ~new_n719_ & ~new_n720_;
  assign new_n722_ = new_n718_ & new_n721_;
  assign new_n723_ = new_n351_ & new_n489_;
  assign new_n724_ = new_n355_ & new_n440_;
  assign new_n725_ = ~new_n723_ & ~new_n724_;
  assign new_n726_ = new_n355_ & new_n444_;
  assign new_n727_ = new_n355_ & new_n446_;
  assign new_n728_ = ~new_n726_ & ~new_n727_;
  assign new_n729_ = new_n725_ & new_n728_;
  assign new_n730_ = new_n722_ & new_n729_;
  assign new_n731_ = new_n355_ & new_n451_;
  assign new_n732_ = new_n355_ & new_n456_;
  assign new_n733_ = ~new_n731_ & ~new_n732_;
  assign new_n734_ = new_n355_ & new_n460_;
  assign new_n735_ = new_n361_ & new_n440_;
  assign new_n736_ = ~new_n734_ & ~new_n735_;
  assign new_n737_ = new_n733_ & new_n736_;
  assign new_n738_ = new_n361_ & new_n444_;
  assign new_n739_ = new_n361_ & new_n446_;
  assign new_n740_ = ~new_n738_ & ~new_n739_;
  assign new_n741_ = new_n361_ & new_n451_;
  assign new_n742_ = new_n361_ & new_n456_;
  assign new_n743_ = ~new_n741_ & ~new_n742_;
  assign new_n744_ = new_n740_ & new_n743_;
  assign new_n745_ = new_n737_ & new_n744_;
  assign new_n746_ = new_n730_ & new_n745_;
  assign new_n747_ = new_n361_ & new_n460_;
  assign new_n748_ = new_n365_ & new_n475_;
  assign new_n749_ = new_n367_ & new_n748_;
  assign new_n750_ = ~new_n747_ & ~new_n749_;
  assign new_n751_ = new_n365_ & new_n469_;
  assign new_n752_ = new_n367_ & new_n751_;
  assign new_n753_ = new_n373_ & new_n563_;
  assign new_n754_ = new_n367_ & new_n753_;
  assign new_n755_ = ~new_n752_ & ~new_n754_;
  assign new_n756_ = new_n750_ & new_n755_;
  assign new_n757_ = new_n379_ & new_n566_;
  assign new_n758_ = new_n367_ & new_n757_;
  assign new_n759_ = new_n379_ & new_n574_;
  assign new_n760_ = new_n367_ & new_n759_;
  assign new_n761_ = ~new_n758_ & ~new_n760_;
  assign new_n762_ = A298 & A269;
  assign new_n763_ = ~A266 & new_n762_;
  assign new_n764_ = new_n453_ & new_n763_;
  assign new_n765_ = new_n140_ & new_n522_;
  assign new_n766_ = new_n764_ & new_n765_;
  assign new_n767_ = A266 & new_n762_;
  assign new_n768_ = new_n453_ & new_n767_;
  assign new_n769_ = ~A265 & A201;
  assign new_n770_ = A200 & new_n769_;
  assign new_n771_ = new_n140_ & new_n770_;
  assign new_n772_ = new_n768_ & new_n771_;
  assign new_n773_ = ~new_n766_ & ~new_n772_;
  assign new_n774_ = new_n761_ & new_n773_;
  assign new_n775_ = new_n756_ & new_n774_;
  assign new_n776_ = new_n140_ & new_n528_;
  assign new_n777_ = new_n764_ & new_n776_;
  assign new_n778_ = A199 & new_n769_;
  assign new_n779_ = new_n140_ & new_n778_;
  assign new_n780_ = new_n768_ & new_n779_;
  assign new_n781_ = ~new_n777_ & ~new_n780_;
  assign new_n782_ = new_n389_ & new_n465_;
  assign new_n783_ = new_n389_ & new_n473_;
  assign new_n784_ = ~new_n782_ & ~new_n783_;
  assign new_n785_ = new_n781_ & new_n784_;
  assign new_n786_ = new_n389_ & new_n487_;
  assign new_n787_ = new_n389_ & new_n476_;
  assign new_n788_ = new_n389_ & new_n470_;
  assign new_n789_ = ~new_n787_ & ~new_n788_;
  assign new_n790_ = ~new_n786_ & new_n789_;
  assign new_n791_ = new_n785_ & new_n790_;
  assign new_n792_ = new_n775_ & new_n791_;
  assign new_n793_ = new_n746_ & new_n792_;
  assign new_n794_ = new_n715_ & new_n793_;
  assign new_n795_ = new_n648_ & new_n794_;
  assign new_n796_ = new_n484_ & new_n795_;
  assign new_n797_ = new_n389_ & new_n489_;
  assign new_n798_ = new_n393_ & new_n465_;
  assign new_n799_ = ~new_n797_ & ~new_n798_;
  assign new_n800_ = new_n393_ & new_n473_;
  assign new_n801_ = new_n393_ & new_n476_;
  assign new_n802_ = ~new_n800_ & ~new_n801_;
  assign new_n803_ = new_n799_ & new_n802_;
  assign new_n804_ = new_n393_ & new_n470_;
  assign new_n805_ = new_n393_ & new_n487_;
  assign new_n806_ = ~new_n804_ & ~new_n805_;
  assign new_n807_ = new_n393_ & new_n489_;
  assign new_n808_ = new_n398_ & new_n440_;
  assign new_n809_ = ~new_n807_ & ~new_n808_;
  assign new_n810_ = new_n806_ & new_n809_;
  assign new_n811_ = new_n803_ & new_n810_;
  assign new_n812_ = new_n398_ & new_n444_;
  assign new_n813_ = new_n398_ & new_n446_;
  assign new_n814_ = ~new_n812_ & ~new_n813_;
  assign new_n815_ = new_n398_ & new_n451_;
  assign new_n816_ = new_n398_ & new_n456_;
  assign new_n817_ = ~new_n815_ & ~new_n816_;
  assign new_n818_ = new_n814_ & new_n817_;
  assign new_n819_ = new_n398_ & new_n460_;
  assign new_n820_ = new_n402_ & new_n440_;
  assign new_n821_ = ~new_n819_ & ~new_n820_;
  assign new_n822_ = new_n402_ & new_n444_;
  assign new_n823_ = new_n402_ & new_n446_;
  assign new_n824_ = ~new_n822_ & ~new_n823_;
  assign new_n825_ = new_n821_ & new_n824_;
  assign new_n826_ = new_n818_ & new_n825_;
  assign new_n827_ = new_n811_ & new_n826_;
  assign new_n828_ = new_n402_ & new_n451_;
  assign new_n829_ = new_n402_ & new_n456_;
  assign new_n830_ = ~new_n828_ & ~new_n829_;
  assign new_n831_ = new_n402_ & new_n460_;
  assign new_n832_ = new_n408_ & new_n748_;
  assign new_n833_ = ~new_n831_ & ~new_n832_;
  assign new_n834_ = new_n830_ & new_n833_;
  assign new_n835_ = new_n408_ & new_n751_;
  assign new_n836_ = new_n408_ & new_n753_;
  assign new_n837_ = ~new_n835_ & ~new_n836_;
  assign new_n838_ = new_n408_ & new_n757_;
  assign new_n839_ = new_n408_ & new_n759_;
  assign new_n840_ = ~new_n838_ & ~new_n839_;
  assign new_n841_ = new_n837_ & new_n840_;
  assign new_n842_ = new_n834_ & new_n841_;
  assign new_n843_ = new_n146_ & new_n522_;
  assign new_n844_ = new_n764_ & new_n843_;
  assign new_n845_ = new_n146_ & new_n770_;
  assign new_n846_ = new_n768_ & new_n845_;
  assign new_n847_ = ~new_n844_ & ~new_n846_;
  assign new_n848_ = new_n146_ & new_n528_;
  assign new_n849_ = new_n764_ & new_n848_;
  assign new_n850_ = new_n146_ & new_n778_;
  assign new_n851_ = new_n768_ & new_n850_;
  assign new_n852_ = ~new_n849_ & ~new_n851_;
  assign new_n853_ = new_n847_ & new_n852_;
  assign new_n854_ = new_n419_ & new_n465_;
  assign new_n855_ = new_n419_ & new_n473_;
  assign new_n856_ = ~new_n854_ & ~new_n855_;
  assign new_n857_ = new_n419_ & new_n476_;
  assign new_n858_ = new_n419_ & new_n470_;
  assign new_n859_ = ~new_n857_ & ~new_n858_;
  assign new_n860_ = new_n856_ & new_n859_;
  assign new_n861_ = new_n853_ & new_n860_;
  assign new_n862_ = new_n842_ & new_n861_;
  assign new_n863_ = new_n827_ & new_n862_;
  assign new_n864_ = new_n419_ & new_n487_;
  assign new_n865_ = new_n419_ & new_n489_;
  assign new_n866_ = ~new_n864_ & ~new_n865_;
  assign new_n867_ = ~A200 & new_n31_;
  assign new_n868_ = ~A199 & A167;
  assign new_n869_ = A168 & new_n868_;
  assign new_n870_ = new_n867_ & new_n869_;
  assign new_n871_ = new_n520_ & new_n870_;
  assign new_n872_ = new_n526_ & new_n870_;
  assign new_n873_ = ~new_n871_ & ~new_n872_;
  assign new_n874_ = new_n866_ & new_n873_;
  assign new_n875_ = A265 & A203;
  assign new_n876_ = ~A200 & new_n875_;
  assign new_n877_ = new_n428_ & new_n876_;
  assign new_n878_ = new_n764_ & new_n877_;
  assign new_n879_ = ~A265 & A203;
  assign new_n880_ = ~A200 & new_n879_;
  assign new_n881_ = new_n428_ & new_n880_;
  assign new_n882_ = new_n768_ & new_n881_;
  assign new_n883_ = ~new_n878_ & ~new_n882_;
  assign new_n884_ = A200 & new_n875_;
  assign new_n885_ = new_n869_ & new_n884_;
  assign new_n886_ = new_n764_ & new_n885_;
  assign new_n887_ = A200 & new_n879_;
  assign new_n888_ = new_n869_ & new_n887_;
  assign new_n889_ = new_n768_ & new_n888_;
  assign new_n890_ = ~new_n886_ & ~new_n889_;
  assign new_n891_ = new_n883_ & new_n890_;
  assign new_n892_ = new_n874_ & new_n891_;
  assign new_n893_ = new_n429_ & new_n465_;
  assign new_n894_ = new_n429_ & new_n473_;
  assign new_n895_ = ~new_n893_ & ~new_n894_;
  assign new_n896_ = new_n429_ & new_n476_;
  assign new_n897_ = new_n429_ & new_n470_;
  assign new_n898_ = ~new_n896_ & ~new_n897_;
  assign new_n899_ = new_n895_ & new_n898_;
  assign new_n900_ = new_n429_ & new_n487_;
  assign new_n901_ = new_n429_ & new_n489_;
  assign new_n902_ = ~new_n900_ & ~new_n901_;
  assign new_n903_ = A265 & ~A203;
  assign new_n904_ = ~A202 & new_n903_;
  assign new_n905_ = ~A201 & A167;
  assign new_n906_ = A168 & new_n905_;
  assign new_n907_ = new_n904_ & new_n906_;
  assign new_n908_ = new_n520_ & new_n907_;
  assign new_n909_ = new_n526_ & new_n907_;
  assign new_n910_ = ~new_n908_ & ~new_n909_;
  assign new_n911_ = new_n902_ & new_n910_;
  assign new_n912_ = new_n899_ & new_n911_;
  assign new_n913_ = new_n892_ & new_n912_;
  assign new_n914_ = A168 & new_n62_;
  assign new_n915_ = new_n867_ & new_n914_;
  assign new_n916_ = new_n520_ & new_n915_;
  assign new_n917_ = new_n526_ & new_n915_;
  assign new_n918_ = ~new_n916_ & ~new_n917_;
  assign new_n919_ = new_n433_ & new_n876_;
  assign new_n920_ = new_n764_ & new_n919_;
  assign new_n921_ = new_n433_ & new_n880_;
  assign new_n922_ = new_n768_ & new_n921_;
  assign new_n923_ = ~new_n920_ & ~new_n922_;
  assign new_n924_ = new_n918_ & new_n923_;
  assign new_n925_ = new_n884_ & new_n914_;
  assign new_n926_ = new_n764_ & new_n925_;
  assign new_n927_ = new_n887_ & new_n914_;
  assign new_n928_ = new_n768_ & new_n927_;
  assign new_n929_ = ~new_n926_ & ~new_n928_;
  assign new_n930_ = new_n434_ & new_n465_;
  assign new_n931_ = new_n434_ & new_n473_;
  assign new_n932_ = ~new_n930_ & ~new_n931_;
  assign new_n933_ = new_n929_ & new_n932_;
  assign new_n934_ = new_n924_ & new_n933_;
  assign new_n935_ = new_n434_ & new_n476_;
  assign new_n936_ = new_n434_ & new_n470_;
  assign new_n937_ = ~new_n935_ & ~new_n936_;
  assign new_n938_ = new_n434_ & new_n487_;
  assign new_n939_ = new_n434_ & new_n489_;
  assign new_n940_ = ~new_n938_ & ~new_n939_;
  assign new_n941_ = new_n937_ & new_n940_;
  assign new_n942_ = ~A168 & new_n190_;
  assign new_n943_ = ~A169 & ~A170;
  assign new_n944_ = new_n942_ & new_n943_;
  assign new_n945_ = new_n504_ & new_n944_;
  assign new_n946_ = A168 & new_n126_;
  assign new_n947_ = new_n904_ & new_n946_;
  assign new_n948_ = new_n520_ & new_n947_;
  assign new_n949_ = new_n526_ & new_n947_;
  assign new_n950_ = ~new_n948_ & ~new_n949_;
  assign new_n951_ = ~new_n945_ & new_n950_;
  assign new_n952_ = new_n941_ & new_n951_;
  assign new_n953_ = new_n934_ & new_n952_;
  assign new_n954_ = new_n913_ & new_n953_;
  assign new_n955_ = new_n863_ & new_n954_;
  assign new_n956_ = new_n506_ & new_n944_;
  assign new_n957_ = new_n509_ & new_n944_;
  assign new_n958_ = ~new_n956_ & ~new_n957_;
  assign new_n959_ = new_n511_ & new_n944_;
  assign new_n960_ = new_n517_ & new_n944_;
  assign new_n961_ = ~new_n959_ & ~new_n960_;
  assign new_n962_ = new_n958_ & new_n961_;
  assign new_n963_ = ~A168 & new_n208_;
  assign new_n964_ = new_n943_ & new_n963_;
  assign new_n965_ = new_n557_ & new_n964_;
  assign new_n966_ = new_n559_ & new_n964_;
  assign new_n967_ = ~new_n965_ & ~new_n966_;
  assign new_n968_ = new_n564_ & new_n964_;
  assign new_n969_ = new_n567_ & new_n964_;
  assign new_n970_ = ~new_n968_ & ~new_n969_;
  assign new_n971_ = new_n967_ & new_n970_;
  assign new_n972_ = new_n962_ & new_n971_;
  assign new_n973_ = new_n575_ & new_n964_;
  assign new_n974_ = ~A168 & new_n240_;
  assign new_n975_ = new_n943_ & new_n974_;
  assign new_n976_ = new_n557_ & new_n975_;
  assign new_n977_ = ~new_n973_ & ~new_n976_;
  assign new_n978_ = new_n559_ & new_n975_;
  assign new_n979_ = new_n564_ & new_n975_;
  assign new_n980_ = ~new_n978_ & ~new_n979_;
  assign new_n981_ = new_n977_ & new_n980_;
  assign new_n982_ = new_n567_ & new_n975_;
  assign new_n983_ = new_n575_ & new_n975_;
  assign new_n984_ = ~new_n982_ & ~new_n983_;
  assign new_n985_ = ~A168 & new_n50_;
  assign new_n986_ = new_n943_ & new_n985_;
  assign new_n987_ = new_n586_ & new_n986_;
  assign new_n988_ = new_n588_ & new_n986_;
  assign new_n989_ = ~new_n987_ & ~new_n988_;
  assign new_n990_ = new_n984_ & new_n989_;
  assign new_n991_ = new_n981_ & new_n990_;
  assign new_n992_ = new_n972_ & new_n991_;
  assign new_n993_ = ~A168 & new_n279_;
  assign new_n994_ = new_n943_ & new_n993_;
  assign new_n995_ = new_n465_ & new_n994_;
  assign new_n996_ = new_n473_ & new_n994_;
  assign new_n997_ = ~new_n995_ & ~new_n996_;
  assign new_n998_ = new_n476_ & new_n994_;
  assign new_n999_ = new_n470_ & new_n994_;
  assign new_n1000_ = ~new_n998_ & ~new_n999_;
  assign new_n1001_ = new_n997_ & new_n1000_;
  assign new_n1002_ = new_n487_ & new_n994_;
  assign new_n1003_ = new_n489_ & new_n994_;
  assign new_n1004_ = ~new_n1002_ & ~new_n1003_;
  assign new_n1005_ = ~A168 & new_n285_;
  assign new_n1006_ = new_n943_ & new_n1005_;
  assign new_n1007_ = new_n465_ & new_n1006_;
  assign new_n1008_ = new_n473_ & new_n1006_;
  assign new_n1009_ = ~new_n1007_ & ~new_n1008_;
  assign new_n1010_ = new_n1004_ & new_n1009_;
  assign new_n1011_ = new_n1001_ & new_n1010_;
  assign new_n1012_ = new_n476_ & new_n1006_;
  assign new_n1013_ = new_n470_ & new_n1006_;
  assign new_n1014_ = ~new_n1012_ & ~new_n1013_;
  assign new_n1015_ = new_n487_ & new_n1006_;
  assign new_n1016_ = new_n489_ & new_n1006_;
  assign new_n1017_ = ~new_n1015_ & ~new_n1016_;
  assign new_n1018_ = new_n1014_ & new_n1017_;
  assign new_n1019_ = ~A168 & new_n49_;
  assign new_n1020_ = new_n943_ & new_n1019_;
  assign new_n1021_ = new_n616_ & new_n1020_;
  assign new_n1022_ = new_n618_ & new_n1020_;
  assign new_n1023_ = ~new_n1021_ & ~new_n1022_;
  assign new_n1024_ = new_n621_ & new_n1020_;
  assign new_n1025_ = new_n623_ & new_n1020_;
  assign new_n1026_ = ~new_n1024_ & ~new_n1025_;
  assign new_n1027_ = new_n1023_ & new_n1026_;
  assign new_n1028_ = new_n1018_ & new_n1027_;
  assign new_n1029_ = new_n1011_ & new_n1028_;
  assign new_n1030_ = new_n992_ & new_n1029_;
  assign new_n1031_ = new_n629_ & new_n1020_;
  assign new_n1032_ = ~A168 & new_n631_;
  assign new_n1033_ = new_n943_ & new_n1032_;
  assign new_n1034_ = new_n520_ & new_n1033_;
  assign new_n1035_ = ~new_n1031_ & ~new_n1034_;
  assign new_n1036_ = new_n526_ & new_n1033_;
  assign new_n1037_ = ~A200 & new_n275_;
  assign new_n1038_ = new_n439_ & new_n1037_;
  assign new_n1039_ = A167 & new_n62_;
  assign new_n1040_ = new_n52_ & new_n1039_;
  assign new_n1041_ = new_n1038_ & new_n1040_;
  assign new_n1042_ = ~new_n1036_ & ~new_n1041_;
  assign new_n1043_ = new_n1035_ & new_n1042_;
  assign new_n1044_ = new_n443_ & new_n1037_;
  assign new_n1045_ = new_n1040_ & new_n1044_;
  assign new_n1046_ = ~A266 & new_n562_;
  assign new_n1047_ = new_n880_ & new_n1046_;
  assign new_n1048_ = A167 & new_n35_;
  assign new_n1049_ = new_n52_ & new_n1048_;
  assign new_n1050_ = new_n1047_ & new_n1049_;
  assign new_n1051_ = ~new_n1045_ & ~new_n1050_;
  assign new_n1052_ = A301 & ~A269;
  assign new_n1053_ = ~A268 & new_n1052_;
  assign new_n1054_ = ~A267 & A203;
  assign new_n1055_ = ~A200 & new_n1054_;
  assign new_n1056_ = new_n1053_ & new_n1055_;
  assign new_n1057_ = new_n1049_ & new_n1056_;
  assign new_n1058_ = new_n887_ & new_n1046_;
  assign new_n1059_ = new_n1040_ & new_n1058_;
  assign new_n1060_ = ~new_n1057_ & ~new_n1059_;
  assign new_n1061_ = new_n1051_ & new_n1060_;
  assign new_n1062_ = new_n1043_ & new_n1061_;
  assign new_n1063_ = A200 & new_n1054_;
  assign new_n1064_ = new_n1053_ & new_n1063_;
  assign new_n1065_ = new_n1040_ & new_n1064_;
  assign new_n1066_ = A201 & new_n205_;
  assign new_n1067_ = new_n475_ & new_n1066_;
  assign new_n1068_ = A200 & A166;
  assign new_n1069_ = A167 & new_n1068_;
  assign new_n1070_ = new_n52_ & new_n1069_;
  assign new_n1071_ = new_n1067_ & new_n1070_;
  assign new_n1072_ = ~new_n1065_ & ~new_n1071_;
  assign new_n1073_ = new_n469_ & new_n1066_;
  assign new_n1074_ = new_n1070_ & new_n1073_;
  assign new_n1075_ = A201 & new_n218_;
  assign new_n1076_ = new_n563_ & new_n1075_;
  assign new_n1077_ = new_n1070_ & new_n1076_;
  assign new_n1078_ = ~new_n1074_ & ~new_n1077_;
  assign new_n1079_ = new_n1072_ & new_n1078_;
  assign new_n1080_ = A201 & new_n216_;
  assign new_n1081_ = new_n566_ & new_n1080_;
  assign new_n1082_ = new_n1070_ & new_n1081_;
  assign new_n1083_ = new_n574_ & new_n1080_;
  assign new_n1084_ = new_n1070_ & new_n1083_;
  assign new_n1085_ = ~new_n1082_ & ~new_n1084_;
  assign new_n1086_ = new_n1049_ & new_n1067_;
  assign new_n1087_ = new_n1049_ & new_n1073_;
  assign new_n1088_ = ~new_n1086_ & ~new_n1087_;
  assign new_n1089_ = new_n1085_ & new_n1088_;
  assign new_n1090_ = new_n1079_ & new_n1089_;
  assign new_n1091_ = new_n1062_ & new_n1090_;
  assign new_n1092_ = new_n1049_ & new_n1076_;
  assign new_n1093_ = new_n1049_ & new_n1081_;
  assign new_n1094_ = ~new_n1092_ & ~new_n1093_;
  assign new_n1095_ = new_n1049_ & new_n1083_;
  assign new_n1096_ = A268 & ~A203;
  assign new_n1097_ = ~A202 & new_n1096_;
  assign new_n1098_ = new_n439_ & new_n1097_;
  assign new_n1099_ = A167 & new_n126_;
  assign new_n1100_ = new_n52_ & new_n1099_;
  assign new_n1101_ = new_n1098_ & new_n1100_;
  assign new_n1102_ = ~new_n1095_ & ~new_n1101_;
  assign new_n1103_ = new_n1094_ & new_n1102_;
  assign new_n1104_ = new_n443_ & new_n1097_;
  assign new_n1105_ = new_n1100_ & new_n1104_;
  assign new_n1106_ = A202 & A166;
  assign new_n1107_ = A167 & new_n1106_;
  assign new_n1108_ = new_n52_ & new_n1107_;
  assign new_n1109_ = new_n465_ & new_n1108_;
  assign new_n1110_ = ~new_n1105_ & ~new_n1109_;
  assign new_n1111_ = new_n473_ & new_n1108_;
  assign new_n1112_ = new_n476_ & new_n1108_;
  assign new_n1113_ = ~new_n1111_ & ~new_n1112_;
  assign new_n1114_ = new_n1110_ & new_n1113_;
  assign new_n1115_ = new_n1103_ & new_n1114_;
  assign new_n1116_ = new_n470_ & new_n1108_;
  assign new_n1117_ = new_n487_ & new_n1108_;
  assign new_n1118_ = ~new_n1116_ & ~new_n1117_;
  assign new_n1119_ = new_n489_ & new_n1108_;
  assign new_n1120_ = ~A166 & new_n190_;
  assign new_n1121_ = ~A167 & ~A169;
  assign new_n1122_ = new_n1120_ & new_n1121_;
  assign new_n1123_ = new_n504_ & new_n1122_;
  assign new_n1124_ = ~new_n1119_ & ~new_n1123_;
  assign new_n1125_ = new_n1118_ & new_n1124_;
  assign new_n1126_ = new_n511_ & new_n1122_;
  assign new_n1127_ = new_n506_ & new_n1122_;
  assign new_n1128_ = new_n509_ & new_n1122_;
  assign new_n1129_ = ~new_n1127_ & ~new_n1128_;
  assign new_n1130_ = ~new_n1126_ & new_n1129_;
  assign new_n1131_ = new_n1125_ & new_n1130_;
  assign new_n1132_ = new_n1115_ & new_n1131_;
  assign new_n1133_ = new_n1091_ & new_n1132_;
  assign new_n1134_ = new_n1030_ & new_n1133_;
  assign new_n1135_ = new_n955_ & new_n1134_;
  assign new_n1136_ = new_n517_ & new_n1122_;
  assign new_n1137_ = ~A166 & new_n208_;
  assign new_n1138_ = new_n1121_ & new_n1137_;
  assign new_n1139_ = new_n557_ & new_n1138_;
  assign new_n1140_ = ~new_n1136_ & ~new_n1139_;
  assign new_n1141_ = new_n559_ & new_n1138_;
  assign new_n1142_ = new_n564_ & new_n1138_;
  assign new_n1143_ = ~new_n1141_ & ~new_n1142_;
  assign new_n1144_ = new_n1140_ & new_n1143_;
  assign new_n1145_ = new_n567_ & new_n1138_;
  assign new_n1146_ = new_n575_ & new_n1138_;
  assign new_n1147_ = ~new_n1145_ & ~new_n1146_;
  assign new_n1148_ = ~A166 & new_n240_;
  assign new_n1149_ = new_n1121_ & new_n1148_;
  assign new_n1150_ = new_n557_ & new_n1149_;
  assign new_n1151_ = new_n559_ & new_n1149_;
  assign new_n1152_ = ~new_n1150_ & ~new_n1151_;
  assign new_n1153_ = new_n1147_ & new_n1152_;
  assign new_n1154_ = new_n1144_ & new_n1153_;
  assign new_n1155_ = new_n564_ & new_n1149_;
  assign new_n1156_ = new_n567_ & new_n1149_;
  assign new_n1157_ = ~new_n1155_ & ~new_n1156_;
  assign new_n1158_ = new_n575_ & new_n1149_;
  assign new_n1159_ = ~A166 & new_n50_;
  assign new_n1160_ = new_n1121_ & new_n1159_;
  assign new_n1161_ = new_n586_ & new_n1160_;
  assign new_n1162_ = ~new_n1158_ & ~new_n1161_;
  assign new_n1163_ = new_n1157_ & new_n1162_;
  assign new_n1164_ = new_n588_ & new_n1160_;
  assign new_n1165_ = ~A166 & new_n279_;
  assign new_n1166_ = new_n1121_ & new_n1165_;
  assign new_n1167_ = new_n465_ & new_n1166_;
  assign new_n1168_ = ~new_n1164_ & ~new_n1167_;
  assign new_n1169_ = new_n473_ & new_n1166_;
  assign new_n1170_ = new_n476_ & new_n1166_;
  assign new_n1171_ = ~new_n1169_ & ~new_n1170_;
  assign new_n1172_ = new_n1168_ & new_n1171_;
  assign new_n1173_ = new_n1163_ & new_n1172_;
  assign new_n1174_ = new_n1154_ & new_n1173_;
  assign new_n1175_ = new_n470_ & new_n1166_;
  assign new_n1176_ = new_n487_ & new_n1166_;
  assign new_n1177_ = ~new_n1175_ & ~new_n1176_;
  assign new_n1178_ = new_n489_ & new_n1166_;
  assign new_n1179_ = ~A166 & new_n285_;
  assign new_n1180_ = new_n1121_ & new_n1179_;
  assign new_n1181_ = new_n465_ & new_n1180_;
  assign new_n1182_ = ~new_n1178_ & ~new_n1181_;
  assign new_n1183_ = new_n1177_ & new_n1182_;
  assign new_n1184_ = new_n473_ & new_n1180_;
  assign new_n1185_ = new_n476_ & new_n1180_;
  assign new_n1186_ = ~new_n1184_ & ~new_n1185_;
  assign new_n1187_ = new_n470_ & new_n1180_;
  assign new_n1188_ = new_n487_ & new_n1180_;
  assign new_n1189_ = ~new_n1187_ & ~new_n1188_;
  assign new_n1190_ = new_n1186_ & new_n1189_;
  assign new_n1191_ = new_n1183_ & new_n1190_;
  assign new_n1192_ = new_n489_ & new_n1180_;
  assign new_n1193_ = ~A166 & new_n49_;
  assign new_n1194_ = new_n1121_ & new_n1193_;
  assign new_n1195_ = new_n616_ & new_n1194_;
  assign new_n1196_ = ~new_n1192_ & ~new_n1195_;
  assign new_n1197_ = new_n618_ & new_n1194_;
  assign new_n1198_ = new_n621_ & new_n1194_;
  assign new_n1199_ = ~new_n1197_ & ~new_n1198_;
  assign new_n1200_ = new_n1196_ & new_n1199_;
  assign new_n1201_ = new_n623_ & new_n1194_;
  assign new_n1202_ = new_n629_ & new_n1194_;
  assign new_n1203_ = ~new_n1201_ & ~new_n1202_;
  assign new_n1204_ = ~A166 & new_n631_;
  assign new_n1205_ = new_n1121_ & new_n1204_;
  assign new_n1206_ = new_n520_ & new_n1205_;
  assign new_n1207_ = new_n526_ & new_n1205_;
  assign new_n1208_ = ~new_n1206_ & ~new_n1207_;
  assign new_n1209_ = new_n1203_ & new_n1208_;
  assign new_n1210_ = new_n1200_ & new_n1209_;
  assign new_n1211_ = new_n1191_ & new_n1210_;
  assign new_n1212_ = new_n1174_ & new_n1211_;
  assign new_n1213_ = ~A199 & A169;
  assign new_n1214_ = new_n867_ & new_n1213_;
  assign new_n1215_ = new_n520_ & new_n1214_;
  assign new_n1216_ = new_n526_ & new_n1214_;
  assign new_n1217_ = ~new_n1215_ & ~new_n1216_;
  assign new_n1218_ = A199 & A169;
  assign new_n1219_ = new_n876_ & new_n1218_;
  assign new_n1220_ = new_n764_ & new_n1219_;
  assign new_n1221_ = new_n880_ & new_n1218_;
  assign new_n1222_ = new_n768_ & new_n1221_;
  assign new_n1223_ = ~new_n1220_ & ~new_n1222_;
  assign new_n1224_ = new_n1217_ & new_n1223_;
  assign new_n1225_ = new_n884_ & new_n1213_;
  assign new_n1226_ = new_n764_ & new_n1225_;
  assign new_n1227_ = new_n887_ & new_n1213_;
  assign new_n1228_ = new_n768_ & new_n1227_;
  assign new_n1229_ = ~new_n1226_ & ~new_n1228_;
  assign new_n1230_ = new_n426_ & new_n1218_;
  assign new_n1231_ = new_n465_ & new_n1230_;
  assign new_n1232_ = new_n473_ & new_n1230_;
  assign new_n1233_ = ~new_n1231_ & ~new_n1232_;
  assign new_n1234_ = new_n1229_ & new_n1233_;
  assign new_n1235_ = new_n1224_ & new_n1234_;
  assign new_n1236_ = new_n476_ & new_n1230_;
  assign new_n1237_ = new_n470_ & new_n1230_;
  assign new_n1238_ = ~new_n1236_ & ~new_n1237_;
  assign new_n1239_ = new_n487_ & new_n1230_;
  assign new_n1240_ = new_n489_ & new_n1230_;
  assign new_n1241_ = ~new_n1239_ & ~new_n1240_;
  assign new_n1242_ = new_n1238_ & new_n1241_;
  assign new_n1243_ = ~A201 & A169;
  assign new_n1244_ = new_n904_ & new_n1243_;
  assign new_n1245_ = new_n520_ & new_n1244_;
  assign new_n1246_ = new_n526_ & new_n1244_;
  assign new_n1247_ = ~new_n1245_ & ~new_n1246_;
  assign new_n1248_ = ~A167 & A170;
  assign new_n1249_ = new_n191_ & new_n1248_;
  assign new_n1250_ = new_n748_ & new_n1249_;
  assign new_n1251_ = new_n751_ & new_n1249_;
  assign new_n1252_ = ~new_n1250_ & ~new_n1251_;
  assign new_n1253_ = new_n1247_ & new_n1252_;
  assign new_n1254_ = new_n1242_ & new_n1253_;
  assign new_n1255_ = new_n1235_ & new_n1254_;
  assign new_n1256_ = new_n753_ & new_n1249_;
  assign new_n1257_ = new_n757_ & new_n1249_;
  assign new_n1258_ = ~new_n1256_ & ~new_n1257_;
  assign new_n1259_ = new_n759_ & new_n1249_;
  assign new_n1260_ = A203 & new_n113_;
  assign new_n1261_ = new_n439_ & new_n1260_;
  assign new_n1262_ = new_n209_ & new_n1248_;
  assign new_n1263_ = new_n1261_ & new_n1262_;
  assign new_n1264_ = ~new_n1259_ & ~new_n1263_;
  assign new_n1265_ = new_n1258_ & new_n1264_;
  assign new_n1266_ = new_n443_ & new_n1260_;
  assign new_n1267_ = new_n1262_ & new_n1266_;
  assign new_n1268_ = A203 & new_n117_;
  assign new_n1269_ = new_n439_ & new_n1268_;
  assign new_n1270_ = new_n1262_ & new_n1269_;
  assign new_n1271_ = ~new_n1267_ & ~new_n1270_;
  assign new_n1272_ = new_n443_ & new_n1268_;
  assign new_n1273_ = new_n1262_ & new_n1272_;
  assign new_n1274_ = A203 & new_n515_;
  assign new_n1275_ = new_n453_ & new_n1274_;
  assign new_n1276_ = new_n1262_ & new_n1275_;
  assign new_n1277_ = ~new_n1273_ & ~new_n1276_;
  assign new_n1278_ = new_n1271_ & new_n1277_;
  assign new_n1279_ = new_n1265_ & new_n1278_;
  assign new_n1280_ = new_n241_ & new_n1248_;
  assign new_n1281_ = new_n1261_ & new_n1280_;
  assign new_n1282_ = new_n1266_ & new_n1280_;
  assign new_n1283_ = ~new_n1281_ & ~new_n1282_;
  assign new_n1284_ = new_n1269_ & new_n1280_;
  assign new_n1285_ = new_n1272_ & new_n1280_;
  assign new_n1286_ = ~new_n1284_ & ~new_n1285_;
  assign new_n1287_ = new_n1283_ & new_n1286_;
  assign new_n1288_ = ~A267 & ~A202;
  assign new_n1289_ = ~A201 & new_n1288_;
  assign new_n1290_ = new_n1053_ & new_n1289_;
  assign new_n1291_ = new_n260_ & new_n1248_;
  assign new_n1292_ = new_n1290_ & new_n1291_;
  assign new_n1293_ = new_n1275_ & new_n1280_;
  assign new_n1294_ = ~A201 & new_n42_;
  assign new_n1295_ = new_n1046_ & new_n1294_;
  assign new_n1296_ = new_n1291_ & new_n1295_;
  assign new_n1297_ = ~new_n1293_ & ~new_n1296_;
  assign new_n1298_ = ~new_n1292_ & new_n1297_;
  assign new_n1299_ = new_n1287_ & new_n1298_;
  assign new_n1300_ = new_n1279_ & new_n1299_;
  assign new_n1301_ = new_n1255_ & new_n1300_;
  assign new_n1302_ = new_n1212_ & new_n1301_;
  assign new_n1303_ = new_n280_ & new_n1248_;
  assign new_n1304_ = new_n440_ & new_n1303_;
  assign new_n1305_ = new_n444_ & new_n1303_;
  assign new_n1306_ = ~new_n1304_ & ~new_n1305_;
  assign new_n1307_ = new_n446_ & new_n1303_;
  assign new_n1308_ = new_n451_ & new_n1303_;
  assign new_n1309_ = ~new_n1307_ & ~new_n1308_;
  assign new_n1310_ = new_n1306_ & new_n1309_;
  assign new_n1311_ = new_n456_ & new_n1303_;
  assign new_n1312_ = new_n460_ & new_n1303_;
  assign new_n1313_ = ~new_n1311_ & ~new_n1312_;
  assign new_n1314_ = new_n286_ & new_n1248_;
  assign new_n1315_ = new_n440_ & new_n1314_;
  assign new_n1316_ = new_n444_ & new_n1314_;
  assign new_n1317_ = ~new_n1315_ & ~new_n1316_;
  assign new_n1318_ = new_n1313_ & new_n1317_;
  assign new_n1319_ = new_n1310_ & new_n1318_;
  assign new_n1320_ = new_n446_ & new_n1314_;
  assign new_n1321_ = new_n451_ & new_n1314_;
  assign new_n1322_ = ~new_n1320_ & ~new_n1321_;
  assign new_n1323_ = new_n456_ & new_n1314_;
  assign new_n1324_ = new_n460_ & new_n1314_;
  assign new_n1325_ = ~new_n1323_ & ~new_n1324_;
  assign new_n1326_ = new_n1322_ & new_n1325_;
  assign new_n1327_ = ~A203 & new_n205_;
  assign new_n1328_ = new_n475_ & new_n1327_;
  assign new_n1329_ = new_n298_ & new_n1248_;
  assign new_n1330_ = new_n1328_ & new_n1329_;
  assign new_n1331_ = new_n469_ & new_n1327_;
  assign new_n1332_ = new_n1329_ & new_n1331_;
  assign new_n1333_ = ~new_n1330_ & ~new_n1332_;
  assign new_n1334_ = ~A203 & new_n218_;
  assign new_n1335_ = new_n563_ & new_n1334_;
  assign new_n1336_ = new_n1329_ & new_n1335_;
  assign new_n1337_ = ~A203 & new_n216_;
  assign new_n1338_ = new_n566_ & new_n1337_;
  assign new_n1339_ = new_n1329_ & new_n1338_;
  assign new_n1340_ = ~new_n1336_ & ~new_n1339_;
  assign new_n1341_ = new_n1333_ & new_n1340_;
  assign new_n1342_ = new_n1326_ & new_n1341_;
  assign new_n1343_ = new_n1319_ & new_n1342_;
  assign new_n1344_ = new_n574_ & new_n1337_;
  assign new_n1345_ = new_n1329_ & new_n1344_;
  assign new_n1346_ = new_n632_ & new_n1248_;
  assign new_n1347_ = new_n764_ & new_n1346_;
  assign new_n1348_ = ~new_n1345_ & ~new_n1347_;
  assign new_n1349_ = ~A265 & A202;
  assign new_n1350_ = A166 & new_n1349_;
  assign new_n1351_ = new_n1248_ & new_n1350_;
  assign new_n1352_ = new_n768_ & new_n1351_;
  assign new_n1353_ = A167 & A170;
  assign new_n1354_ = new_n1120_ & new_n1353_;
  assign new_n1355_ = new_n748_ & new_n1354_;
  assign new_n1356_ = ~new_n1352_ & ~new_n1355_;
  assign new_n1357_ = new_n1348_ & new_n1356_;
  assign new_n1358_ = new_n751_ & new_n1354_;
  assign new_n1359_ = new_n753_ & new_n1354_;
  assign new_n1360_ = ~new_n1358_ & ~new_n1359_;
  assign new_n1361_ = new_n757_ & new_n1354_;
  assign new_n1362_ = new_n759_ & new_n1354_;
  assign new_n1363_ = ~new_n1361_ & ~new_n1362_;
  assign new_n1364_ = new_n1360_ & new_n1363_;
  assign new_n1365_ = new_n1357_ & new_n1364_;
  assign new_n1366_ = new_n1137_ & new_n1353_;
  assign new_n1367_ = new_n1261_ & new_n1366_;
  assign new_n1368_ = new_n1266_ & new_n1366_;
  assign new_n1369_ = ~new_n1367_ & ~new_n1368_;
  assign new_n1370_ = new_n1269_ & new_n1366_;
  assign new_n1371_ = new_n1272_ & new_n1366_;
  assign new_n1372_ = ~new_n1370_ & ~new_n1371_;
  assign new_n1373_ = new_n1369_ & new_n1372_;
  assign new_n1374_ = new_n1275_ & new_n1366_;
  assign new_n1375_ = new_n1148_ & new_n1353_;
  assign new_n1376_ = new_n1261_ & new_n1375_;
  assign new_n1377_ = ~new_n1374_ & ~new_n1376_;
  assign new_n1378_ = new_n1266_ & new_n1375_;
  assign new_n1379_ = new_n1269_ & new_n1375_;
  assign new_n1380_ = ~new_n1378_ & ~new_n1379_;
  assign new_n1381_ = new_n1377_ & new_n1380_;
  assign new_n1382_ = new_n1373_ & new_n1381_;
  assign new_n1383_ = new_n1365_ & new_n1382_;
  assign new_n1384_ = new_n1343_ & new_n1383_;
  assign new_n1385_ = new_n1272_ & new_n1375_;
  assign new_n1386_ = new_n1275_ & new_n1375_;
  assign new_n1387_ = ~new_n1385_ & ~new_n1386_;
  assign new_n1388_ = new_n1159_ & new_n1353_;
  assign new_n1389_ = new_n1295_ & new_n1388_;
  assign new_n1390_ = new_n1290_ & new_n1388_;
  assign new_n1391_ = ~new_n1389_ & ~new_n1390_;
  assign new_n1392_ = new_n1387_ & new_n1391_;
  assign new_n1393_ = new_n1165_ & new_n1353_;
  assign new_n1394_ = new_n440_ & new_n1393_;
  assign new_n1395_ = new_n444_ & new_n1393_;
  assign new_n1396_ = ~new_n1394_ & ~new_n1395_;
  assign new_n1397_ = new_n446_ & new_n1393_;
  assign new_n1398_ = new_n451_ & new_n1393_;
  assign new_n1399_ = ~new_n1397_ & ~new_n1398_;
  assign new_n1400_ = new_n1396_ & new_n1399_;
  assign new_n1401_ = new_n1392_ & new_n1400_;
  assign new_n1402_ = new_n456_ & new_n1393_;
  assign new_n1403_ = new_n460_ & new_n1393_;
  assign new_n1404_ = ~new_n1402_ & ~new_n1403_;
  assign new_n1405_ = new_n1179_ & new_n1353_;
  assign new_n1406_ = new_n440_ & new_n1405_;
  assign new_n1407_ = new_n444_ & new_n1405_;
  assign new_n1408_ = ~new_n1406_ & ~new_n1407_;
  assign new_n1409_ = new_n1404_ & new_n1408_;
  assign new_n1410_ = new_n446_ & new_n1405_;
  assign new_n1411_ = new_n451_ & new_n1405_;
  assign new_n1412_ = ~new_n1410_ & ~new_n1411_;
  assign new_n1413_ = new_n456_ & new_n1405_;
  assign new_n1414_ = new_n460_ & new_n1405_;
  assign new_n1415_ = ~new_n1413_ & ~new_n1414_;
  assign new_n1416_ = new_n1412_ & new_n1415_;
  assign new_n1417_ = new_n1409_ & new_n1416_;
  assign new_n1418_ = new_n1401_ & new_n1417_;
  assign new_n1419_ = new_n1193_ & new_n1353_;
  assign new_n1420_ = new_n1328_ & new_n1419_;
  assign new_n1421_ = new_n1331_ & new_n1419_;
  assign new_n1422_ = ~new_n1420_ & ~new_n1421_;
  assign new_n1423_ = new_n1335_ & new_n1419_;
  assign new_n1424_ = new_n1338_ & new_n1419_;
  assign new_n1425_ = ~new_n1423_ & ~new_n1424_;
  assign new_n1426_ = new_n1422_ & new_n1425_;
  assign new_n1427_ = new_n1344_ & new_n1419_;
  assign new_n1428_ = new_n1204_ & new_n1353_;
  assign new_n1429_ = new_n764_ & new_n1428_;
  assign new_n1430_ = ~new_n1427_ & ~new_n1429_;
  assign new_n1431_ = ~A166 & new_n1349_;
  assign new_n1432_ = new_n1353_ & new_n1431_;
  assign new_n1433_ = new_n768_ & new_n1432_;
  assign new_n1434_ = A167 & A168;
  assign new_n1435_ = new_n153_ & new_n1434_;
  assign new_n1436_ = new_n465_ & new_n1435_;
  assign new_n1437_ = ~new_n1433_ & ~new_n1436_;
  assign new_n1438_ = new_n1430_ & new_n1437_;
  assign new_n1439_ = new_n1426_ & new_n1438_;
  assign new_n1440_ = new_n473_ & new_n1435_;
  assign new_n1441_ = new_n476_ & new_n1435_;
  assign new_n1442_ = ~new_n1440_ & ~new_n1441_;
  assign new_n1443_ = new_n470_ & new_n1435_;
  assign new_n1444_ = new_n487_ & new_n1435_;
  assign new_n1445_ = ~new_n1443_ & ~new_n1444_;
  assign new_n1446_ = new_n1442_ & new_n1445_;
  assign new_n1447_ = new_n158_ & new_n1434_;
  assign new_n1448_ = new_n444_ & new_n1447_;
  assign new_n1449_ = new_n489_ & new_n1435_;
  assign new_n1450_ = new_n440_ & new_n1447_;
  assign new_n1451_ = ~new_n1449_ & ~new_n1450_;
  assign new_n1452_ = ~new_n1448_ & new_n1451_;
  assign new_n1453_ = new_n1446_ & new_n1452_;
  assign new_n1454_ = new_n1439_ & new_n1453_;
  assign new_n1455_ = new_n1418_ & new_n1454_;
  assign new_n1456_ = new_n1384_ & new_n1455_;
  assign new_n1457_ = new_n1302_ & new_n1456_;
  assign new_n1458_ = new_n1135_ & new_n1457_;
  assign new_n1459_ = new_n796_ & new_n1458_;
  assign new_n1460_ = new_n446_ & new_n1447_;
  assign new_n1461_ = new_n451_ & new_n1447_;
  assign new_n1462_ = ~new_n1460_ & ~new_n1461_;
  assign new_n1463_ = new_n456_ & new_n1447_;
  assign new_n1464_ = new_n460_ & new_n1447_;
  assign new_n1465_ = ~new_n1463_ & ~new_n1464_;
  assign new_n1466_ = new_n1462_ & new_n1465_;
  assign new_n1467_ = new_n164_ & new_n1434_;
  assign new_n1468_ = new_n440_ & new_n1467_;
  assign new_n1469_ = new_n444_ & new_n1467_;
  assign new_n1470_ = ~new_n1468_ & ~new_n1469_;
  assign new_n1471_ = new_n446_ & new_n1467_;
  assign new_n1472_ = new_n451_ & new_n1467_;
  assign new_n1473_ = ~new_n1471_ & ~new_n1472_;
  assign new_n1474_ = new_n1470_ & new_n1473_;
  assign new_n1475_ = new_n1466_ & new_n1474_;
  assign new_n1476_ = new_n456_ & new_n1467_;
  assign new_n1477_ = new_n460_ & new_n1467_;
  assign new_n1478_ = ~new_n1476_ & ~new_n1477_;
  assign new_n1479_ = new_n169_ & new_n1434_;
  assign new_n1480_ = new_n748_ & new_n1479_;
  assign new_n1481_ = new_n751_ & new_n1479_;
  assign new_n1482_ = ~new_n1480_ & ~new_n1481_;
  assign new_n1483_ = new_n1478_ & new_n1482_;
  assign new_n1484_ = new_n753_ & new_n1479_;
  assign new_n1485_ = new_n757_ & new_n1479_;
  assign new_n1486_ = ~new_n1484_ & ~new_n1485_;
  assign new_n1487_ = new_n759_ & new_n1479_;
  assign new_n1488_ = new_n522_ & new_n1434_;
  assign new_n1489_ = new_n764_ & new_n1488_;
  assign new_n1490_ = ~new_n1487_ & ~new_n1489_;
  assign new_n1491_ = new_n1486_ & new_n1490_;
  assign new_n1492_ = new_n1483_ & new_n1491_;
  assign new_n1493_ = new_n1475_ & new_n1492_;
  assign new_n1494_ = new_n770_ & new_n1434_;
  assign new_n1495_ = new_n768_ & new_n1494_;
  assign new_n1496_ = new_n528_ & new_n1434_;
  assign new_n1497_ = new_n764_ & new_n1496_;
  assign new_n1498_ = ~new_n1495_ & ~new_n1497_;
  assign new_n1499_ = new_n778_ & new_n1434_;
  assign new_n1500_ = new_n768_ & new_n1499_;
  assign new_n1501_ = new_n185_ & new_n1434_;
  assign new_n1502_ = new_n465_ & new_n1501_;
  assign new_n1503_ = ~new_n1500_ & ~new_n1502_;
  assign new_n1504_ = new_n1498_ & new_n1503_;
  assign new_n1505_ = new_n473_ & new_n1501_;
  assign new_n1506_ = new_n476_ & new_n1501_;
  assign new_n1507_ = ~new_n1505_ & ~new_n1506_;
  assign new_n1508_ = new_n470_ & new_n1501_;
  assign new_n1509_ = new_n487_ & new_n1501_;
  assign new_n1510_ = ~new_n1508_ & ~new_n1509_;
  assign new_n1511_ = new_n1507_ & new_n1510_;
  assign new_n1512_ = new_n1504_ & new_n1511_;
  assign new_n1513_ = new_n489_ & new_n1501_;
  assign new_n1514_ = A166 & A168;
  assign new_n1515_ = new_n153_ & new_n1514_;
  assign new_n1516_ = new_n465_ & new_n1515_;
  assign new_n1517_ = ~new_n1513_ & ~new_n1516_;
  assign new_n1518_ = new_n473_ & new_n1515_;
  assign new_n1519_ = new_n476_ & new_n1515_;
  assign new_n1520_ = ~new_n1518_ & ~new_n1519_;
  assign new_n1521_ = new_n1517_ & new_n1520_;
  assign new_n1522_ = new_n470_ & new_n1515_;
  assign new_n1523_ = new_n487_ & new_n1515_;
  assign new_n1524_ = ~new_n1522_ & ~new_n1523_;
  assign new_n1525_ = new_n489_ & new_n1515_;
  assign new_n1526_ = new_n158_ & new_n1514_;
  assign new_n1527_ = new_n440_ & new_n1526_;
  assign new_n1528_ = ~new_n1525_ & ~new_n1527_;
  assign new_n1529_ = new_n1524_ & new_n1528_;
  assign new_n1530_ = new_n1521_ & new_n1529_;
  assign new_n1531_ = new_n1512_ & new_n1530_;
  assign new_n1532_ = new_n1493_ & new_n1531_;
  assign new_n1533_ = new_n444_ & new_n1526_;
  assign new_n1534_ = new_n446_ & new_n1526_;
  assign new_n1535_ = ~new_n1533_ & ~new_n1534_;
  assign new_n1536_ = new_n451_ & new_n1526_;
  assign new_n1537_ = new_n456_ & new_n1526_;
  assign new_n1538_ = ~new_n1536_ & ~new_n1537_;
  assign new_n1539_ = new_n1535_ & new_n1538_;
  assign new_n1540_ = new_n460_ & new_n1526_;
  assign new_n1541_ = new_n164_ & new_n1514_;
  assign new_n1542_ = new_n440_ & new_n1541_;
  assign new_n1543_ = ~new_n1540_ & ~new_n1542_;
  assign new_n1544_ = new_n444_ & new_n1541_;
  assign new_n1545_ = new_n446_ & new_n1541_;
  assign new_n1546_ = ~new_n1544_ & ~new_n1545_;
  assign new_n1547_ = new_n1543_ & new_n1546_;
  assign new_n1548_ = new_n1539_ & new_n1547_;
  assign new_n1549_ = new_n451_ & new_n1541_;
  assign new_n1550_ = new_n456_ & new_n1541_;
  assign new_n1551_ = ~new_n1549_ & ~new_n1550_;
  assign new_n1552_ = new_n460_ & new_n1541_;
  assign new_n1553_ = new_n169_ & new_n1514_;
  assign new_n1554_ = new_n748_ & new_n1553_;
  assign new_n1555_ = ~new_n1552_ & ~new_n1554_;
  assign new_n1556_ = new_n1551_ & new_n1555_;
  assign new_n1557_ = new_n751_ & new_n1553_;
  assign new_n1558_ = new_n753_ & new_n1553_;
  assign new_n1559_ = ~new_n1557_ & ~new_n1558_;
  assign new_n1560_ = new_n757_ & new_n1553_;
  assign new_n1561_ = new_n759_ & new_n1553_;
  assign new_n1562_ = ~new_n1560_ & ~new_n1561_;
  assign new_n1563_ = new_n1559_ & new_n1562_;
  assign new_n1564_ = new_n1556_ & new_n1563_;
  assign new_n1565_ = new_n1548_ & new_n1564_;
  assign new_n1566_ = new_n522_ & new_n1514_;
  assign new_n1567_ = new_n764_ & new_n1566_;
  assign new_n1568_ = new_n770_ & new_n1514_;
  assign new_n1569_ = new_n768_ & new_n1568_;
  assign new_n1570_ = ~new_n1567_ & ~new_n1569_;
  assign new_n1571_ = new_n528_ & new_n1514_;
  assign new_n1572_ = new_n764_ & new_n1571_;
  assign new_n1573_ = new_n778_ & new_n1514_;
  assign new_n1574_ = new_n768_ & new_n1573_;
  assign new_n1575_ = ~new_n1572_ & ~new_n1574_;
  assign new_n1576_ = new_n1570_ & new_n1575_;
  assign new_n1577_ = new_n185_ & new_n1514_;
  assign new_n1578_ = new_n465_ & new_n1577_;
  assign new_n1579_ = new_n473_ & new_n1577_;
  assign new_n1580_ = ~new_n1578_ & ~new_n1579_;
  assign new_n1581_ = new_n476_ & new_n1577_;
  assign new_n1582_ = new_n470_ & new_n1577_;
  assign new_n1583_ = ~new_n1581_ & ~new_n1582_;
  assign new_n1584_ = new_n1580_ & new_n1583_;
  assign new_n1585_ = new_n1576_ & new_n1584_;
  assign new_n1586_ = new_n487_ & new_n1577_;
  assign new_n1587_ = new_n489_ & new_n1577_;
  assign new_n1588_ = ~new_n1586_ & ~new_n1587_;
  assign new_n1589_ = new_n275_ & new_n439_;
  assign new_n1590_ = new_n944_ & new_n1589_;
  assign new_n1591_ = new_n275_ & new_n443_;
  assign new_n1592_ = new_n944_ & new_n1591_;
  assign new_n1593_ = ~new_n1590_ & ~new_n1592_;
  assign new_n1594_ = new_n1588_ & new_n1593_;
  assign new_n1595_ = new_n879_ & new_n1046_;
  assign new_n1596_ = new_n964_ & new_n1595_;
  assign new_n1597_ = new_n1053_ & new_n1054_;
  assign new_n1598_ = new_n964_ & new_n1597_;
  assign new_n1599_ = ~new_n1596_ & ~new_n1598_;
  assign new_n1600_ = new_n975_ & new_n1595_;
  assign new_n1601_ = new_n975_ & new_n1597_;
  assign new_n1602_ = ~new_n1600_ & ~new_n1601_;
  assign new_n1603_ = new_n1599_ & new_n1602_;
  assign new_n1604_ = new_n1594_ & new_n1603_;
  assign new_n1605_ = new_n1585_ & new_n1604_;
  assign new_n1606_ = new_n1565_ & new_n1605_;
  assign new_n1607_ = new_n1532_ & new_n1606_;
  assign new_n1608_ = new_n205_ & new_n475_;
  assign new_n1609_ = new_n994_ & new_n1608_;
  assign new_n1610_ = new_n205_ & new_n469_;
  assign new_n1611_ = new_n994_ & new_n1610_;
  assign new_n1612_ = ~new_n1609_ & ~new_n1611_;
  assign new_n1613_ = new_n218_ & new_n563_;
  assign new_n1614_ = new_n994_ & new_n1613_;
  assign new_n1615_ = new_n216_ & new_n566_;
  assign new_n1616_ = new_n994_ & new_n1615_;
  assign new_n1617_ = ~new_n1614_ & ~new_n1616_;
  assign new_n1618_ = new_n1612_ & new_n1617_;
  assign new_n1619_ = new_n216_ & new_n574_;
  assign new_n1620_ = new_n994_ & new_n1619_;
  assign new_n1621_ = new_n1006_ & new_n1608_;
  assign new_n1622_ = ~new_n1620_ & ~new_n1621_;
  assign new_n1623_ = new_n1006_ & new_n1610_;
  assign new_n1624_ = new_n1006_ & new_n1613_;
  assign new_n1625_ = ~new_n1623_ & ~new_n1624_;
  assign new_n1626_ = new_n1622_ & new_n1625_;
  assign new_n1627_ = new_n1618_ & new_n1626_;
  assign new_n1628_ = new_n1006_ & new_n1615_;
  assign new_n1629_ = new_n1006_ & new_n1619_;
  assign new_n1630_ = ~new_n1628_ & ~new_n1629_;
  assign new_n1631_ = new_n439_ & new_n1096_;
  assign new_n1632_ = new_n1020_ & new_n1631_;
  assign new_n1633_ = new_n443_ & new_n1096_;
  assign new_n1634_ = new_n1020_ & new_n1633_;
  assign new_n1635_ = ~new_n1632_ & ~new_n1634_;
  assign new_n1636_ = new_n1630_ & new_n1635_;
  assign new_n1637_ = new_n462_ & new_n463_;
  assign new_n1638_ = ~A168 & new_n1349_;
  assign new_n1639_ = new_n943_ & new_n1638_;
  assign new_n1640_ = new_n1637_ & new_n1639_;
  assign new_n1641_ = new_n463_ & new_n472_;
  assign new_n1642_ = new_n1639_ & new_n1641_;
  assign new_n1643_ = ~new_n1640_ & ~new_n1642_;
  assign new_n1644_ = new_n71_ & new_n475_;
  assign new_n1645_ = new_n1033_ & new_n1644_;
  assign new_n1646_ = new_n71_ & new_n469_;
  assign new_n1647_ = new_n1033_ & new_n1646_;
  assign new_n1648_ = ~new_n1645_ & ~new_n1647_;
  assign new_n1649_ = new_n1643_ & new_n1648_;
  assign new_n1650_ = new_n1636_ & new_n1649_;
  assign new_n1651_ = new_n1627_ & new_n1650_;
  assign new_n1652_ = new_n462_ & new_n485_;
  assign new_n1653_ = ~A267 & A202;
  assign new_n1654_ = ~A168 & new_n1653_;
  assign new_n1655_ = new_n943_ & new_n1654_;
  assign new_n1656_ = new_n1652_ & new_n1655_;
  assign new_n1657_ = new_n472_ & new_n485_;
  assign new_n1658_ = new_n1655_ & new_n1657_;
  assign new_n1659_ = ~new_n1656_ & ~new_n1658_;
  assign new_n1660_ = new_n769_ & new_n1046_;
  assign new_n1661_ = new_n1070_ & new_n1660_;
  assign new_n1662_ = ~A267 & A201;
  assign new_n1663_ = new_n1053_ & new_n1662_;
  assign new_n1664_ = new_n1070_ & new_n1663_;
  assign new_n1665_ = ~new_n1661_ & ~new_n1664_;
  assign new_n1666_ = new_n1659_ & new_n1665_;
  assign new_n1667_ = new_n1049_ & new_n1660_;
  assign new_n1668_ = new_n1049_ & new_n1663_;
  assign new_n1669_ = ~new_n1667_ & ~new_n1668_;
  assign new_n1670_ = new_n1108_ & new_n1608_;
  assign new_n1671_ = new_n1108_ & new_n1610_;
  assign new_n1672_ = ~new_n1670_ & ~new_n1671_;
  assign new_n1673_ = new_n1669_ & new_n1672_;
  assign new_n1674_ = new_n1666_ & new_n1673_;
  assign new_n1675_ = new_n1108_ & new_n1613_;
  assign new_n1676_ = new_n1108_ & new_n1615_;
  assign new_n1677_ = ~new_n1675_ & ~new_n1676_;
  assign new_n1678_ = new_n1108_ & new_n1619_;
  assign new_n1679_ = new_n1122_ & new_n1589_;
  assign new_n1680_ = ~new_n1678_ & ~new_n1679_;
  assign new_n1681_ = new_n1677_ & new_n1680_;
  assign new_n1682_ = new_n1122_ & new_n1591_;
  assign new_n1683_ = new_n1138_ & new_n1595_;
  assign new_n1684_ = ~new_n1682_ & ~new_n1683_;
  assign new_n1685_ = new_n1138_ & new_n1597_;
  assign new_n1686_ = new_n1149_ & new_n1595_;
  assign new_n1687_ = ~new_n1685_ & ~new_n1686_;
  assign new_n1688_ = new_n1684_ & new_n1687_;
  assign new_n1689_ = new_n1681_ & new_n1688_;
  assign new_n1690_ = new_n1674_ & new_n1689_;
  assign new_n1691_ = new_n1651_ & new_n1690_;
  assign new_n1692_ = new_n1149_ & new_n1597_;
  assign new_n1693_ = new_n1166_ & new_n1608_;
  assign new_n1694_ = ~new_n1692_ & ~new_n1693_;
  assign new_n1695_ = new_n1166_ & new_n1610_;
  assign new_n1696_ = new_n1166_ & new_n1613_;
  assign new_n1697_ = ~new_n1695_ & ~new_n1696_;
  assign new_n1698_ = new_n1694_ & new_n1697_;
  assign new_n1699_ = new_n1166_ & new_n1615_;
  assign new_n1700_ = new_n1166_ & new_n1619_;
  assign new_n1701_ = ~new_n1699_ & ~new_n1700_;
  assign new_n1702_ = new_n1180_ & new_n1608_;
  assign new_n1703_ = new_n1180_ & new_n1610_;
  assign new_n1704_ = ~new_n1702_ & ~new_n1703_;
  assign new_n1705_ = new_n1701_ & new_n1704_;
  assign new_n1706_ = new_n1698_ & new_n1705_;
  assign new_n1707_ = new_n1180_ & new_n1613_;
  assign new_n1708_ = new_n1180_ & new_n1615_;
  assign new_n1709_ = ~new_n1707_ & ~new_n1708_;
  assign new_n1710_ = new_n1180_ & new_n1619_;
  assign new_n1711_ = new_n1194_ & new_n1631_;
  assign new_n1712_ = ~new_n1710_ & ~new_n1711_;
  assign new_n1713_ = new_n1709_ & new_n1712_;
  assign new_n1714_ = new_n1194_ & new_n1633_;
  assign new_n1715_ = new_n1121_ & new_n1431_;
  assign new_n1716_ = new_n1637_ & new_n1715_;
  assign new_n1717_ = ~new_n1714_ & ~new_n1716_;
  assign new_n1718_ = new_n1641_ & new_n1715_;
  assign new_n1719_ = new_n1205_ & new_n1644_;
  assign new_n1720_ = ~new_n1718_ & ~new_n1719_;
  assign new_n1721_ = new_n1717_ & new_n1720_;
  assign new_n1722_ = new_n1713_ & new_n1721_;
  assign new_n1723_ = new_n1706_ & new_n1722_;
  assign new_n1724_ = new_n1205_ & new_n1646_;
  assign new_n1725_ = ~A166 & new_n1653_;
  assign new_n1726_ = new_n1121_ & new_n1725_;
  assign new_n1727_ = new_n1652_ & new_n1726_;
  assign new_n1728_ = ~new_n1724_ & ~new_n1727_;
  assign new_n1729_ = new_n1657_ & new_n1726_;
  assign new_n1730_ = ~A200 & new_n42_;
  assign new_n1731_ = new_n1213_ & new_n1730_;
  assign new_n1732_ = new_n1637_ & new_n1731_;
  assign new_n1733_ = ~new_n1729_ & ~new_n1732_;
  assign new_n1734_ = new_n1728_ & new_n1733_;
  assign new_n1735_ = new_n1641_ & new_n1731_;
  assign new_n1736_ = new_n1214_ & new_n1644_;
  assign new_n1737_ = ~new_n1735_ & ~new_n1736_;
  assign new_n1738_ = new_n1214_ & new_n1646_;
  assign new_n1739_ = ~A200 & new_n1288_;
  assign new_n1740_ = new_n1213_ & new_n1739_;
  assign new_n1741_ = new_n1652_ & new_n1740_;
  assign new_n1742_ = ~new_n1738_ & ~new_n1741_;
  assign new_n1743_ = new_n1737_ & new_n1742_;
  assign new_n1744_ = new_n1734_ & new_n1743_;
  assign new_n1745_ = new_n1657_ & new_n1740_;
  assign new_n1746_ = new_n30_ & new_n439_;
  assign new_n1747_ = new_n1219_ & new_n1746_;
  assign new_n1748_ = ~new_n1745_ & ~new_n1747_;
  assign new_n1749_ = new_n30_ & new_n443_;
  assign new_n1750_ = new_n1219_ & new_n1749_;
  assign new_n1751_ = new_n41_ & new_n439_;
  assign new_n1752_ = new_n1221_ & new_n1751_;
  assign new_n1753_ = ~new_n1750_ & ~new_n1752_;
  assign new_n1754_ = new_n1748_ & new_n1753_;
  assign new_n1755_ = new_n453_ & new_n454_;
  assign new_n1756_ = new_n1219_ & new_n1755_;
  assign new_n1757_ = new_n41_ & new_n443_;
  assign new_n1758_ = new_n1221_ & new_n1757_;
  assign new_n1759_ = A266 & A203;
  assign new_n1760_ = ~A200 & new_n1759_;
  assign new_n1761_ = new_n1218_ & new_n1760_;
  assign new_n1762_ = new_n1755_ & new_n1761_;
  assign new_n1763_ = ~new_n1758_ & ~new_n1762_;
  assign new_n1764_ = ~new_n1756_ & new_n1763_;
  assign new_n1765_ = new_n1754_ & new_n1764_;
  assign new_n1766_ = new_n1744_ & new_n1765_;
  assign new_n1767_ = new_n1723_ & new_n1766_;
  assign new_n1768_ = new_n1691_ & new_n1767_;
  assign new_n1769_ = new_n1607_ & new_n1768_;
  assign new_n1770_ = new_n1225_ & new_n1746_;
  assign new_n1771_ = new_n1225_ & new_n1749_;
  assign new_n1772_ = ~new_n1770_ & ~new_n1771_;
  assign new_n1773_ = new_n1227_ & new_n1751_;
  assign new_n1774_ = new_n1227_ & new_n1757_;
  assign new_n1775_ = ~new_n1773_ & ~new_n1774_;
  assign new_n1776_ = new_n1772_ & new_n1775_;
  assign new_n1777_ = A200 & new_n1759_;
  assign new_n1778_ = new_n1213_ & new_n1777_;
  assign new_n1779_ = new_n1755_ & new_n1778_;
  assign new_n1780_ = new_n1225_ & new_n1755_;
  assign new_n1781_ = ~new_n1779_ & ~new_n1780_;
  assign new_n1782_ = new_n1230_ & new_n1608_;
  assign new_n1783_ = new_n1230_ & new_n1610_;
  assign new_n1784_ = ~new_n1782_ & ~new_n1783_;
  assign new_n1785_ = new_n1781_ & new_n1784_;
  assign new_n1786_ = new_n1776_ & new_n1785_;
  assign new_n1787_ = new_n1230_ & new_n1613_;
  assign new_n1788_ = new_n1230_ & new_n1615_;
  assign new_n1789_ = ~new_n1787_ & ~new_n1788_;
  assign new_n1790_ = new_n1230_ & new_n1619_;
  assign new_n1791_ = new_n453_ & new_n762_;
  assign new_n1792_ = A201 & new_n95_;
  assign new_n1793_ = A200 & A169;
  assign new_n1794_ = new_n1792_ & new_n1793_;
  assign new_n1795_ = new_n1791_ & new_n1794_;
  assign new_n1796_ = ~new_n1790_ & ~new_n1795_;
  assign new_n1797_ = new_n1789_ & new_n1796_;
  assign new_n1798_ = A201 & new_n106_;
  assign new_n1799_ = new_n1793_ & new_n1798_;
  assign new_n1800_ = new_n1791_ & new_n1799_;
  assign new_n1801_ = new_n1218_ & new_n1792_;
  assign new_n1802_ = new_n1791_ & new_n1801_;
  assign new_n1803_ = ~new_n1800_ & ~new_n1802_;
  assign new_n1804_ = new_n1218_ & new_n1798_;
  assign new_n1805_ = new_n1791_ & new_n1804_;
  assign new_n1806_ = ~A265 & ~A203;
  assign new_n1807_ = ~A202 & new_n1806_;
  assign new_n1808_ = new_n1243_ & new_n1807_;
  assign new_n1809_ = new_n1637_ & new_n1808_;
  assign new_n1810_ = ~new_n1805_ & ~new_n1809_;
  assign new_n1811_ = new_n1803_ & new_n1810_;
  assign new_n1812_ = new_n1797_ & new_n1811_;
  assign new_n1813_ = new_n1786_ & new_n1812_;
  assign new_n1814_ = new_n1641_ & new_n1808_;
  assign new_n1815_ = new_n1244_ & new_n1644_;
  assign new_n1816_ = ~new_n1814_ & ~new_n1815_;
  assign new_n1817_ = new_n1244_ & new_n1646_;
  assign new_n1818_ = ~A267 & ~A203;
  assign new_n1819_ = ~A202 & new_n1818_;
  assign new_n1820_ = new_n1243_ & new_n1819_;
  assign new_n1821_ = new_n1652_ & new_n1820_;
  assign new_n1822_ = ~new_n1817_ & ~new_n1821_;
  assign new_n1823_ = new_n1816_ & new_n1822_;
  assign new_n1824_ = new_n1657_ & new_n1820_;
  assign new_n1825_ = new_n42_ & new_n1046_;
  assign new_n1826_ = new_n1249_ & new_n1825_;
  assign new_n1827_ = ~new_n1824_ & ~new_n1826_;
  assign new_n1828_ = new_n1053_ & new_n1288_;
  assign new_n1829_ = new_n1249_ & new_n1828_;
  assign new_n1830_ = A268 & A203;
  assign new_n1831_ = new_n439_ & new_n1830_;
  assign new_n1832_ = new_n1262_ & new_n1831_;
  assign new_n1833_ = ~new_n1829_ & ~new_n1832_;
  assign new_n1834_ = new_n1827_ & new_n1833_;
  assign new_n1835_ = new_n1823_ & new_n1834_;
  assign new_n1836_ = new_n443_ & new_n1830_;
  assign new_n1837_ = new_n1262_ & new_n1836_;
  assign new_n1838_ = new_n1280_ & new_n1831_;
  assign new_n1839_ = ~new_n1837_ & ~new_n1838_;
  assign new_n1840_ = new_n1280_ & new_n1836_;
  assign new_n1841_ = new_n113_ & new_n439_;
  assign new_n1842_ = new_n1303_ & new_n1841_;
  assign new_n1843_ = ~new_n1840_ & ~new_n1842_;
  assign new_n1844_ = new_n1839_ & new_n1843_;
  assign new_n1845_ = new_n113_ & new_n443_;
  assign new_n1846_ = new_n1303_ & new_n1845_;
  assign new_n1847_ = new_n117_ & new_n439_;
  assign new_n1848_ = new_n1303_ & new_n1847_;
  assign new_n1849_ = ~new_n1846_ & ~new_n1848_;
  assign new_n1850_ = new_n117_ & new_n443_;
  assign new_n1851_ = new_n1303_ & new_n1850_;
  assign new_n1852_ = new_n453_ & new_n515_;
  assign new_n1853_ = new_n1303_ & new_n1852_;
  assign new_n1854_ = ~new_n1851_ & ~new_n1853_;
  assign new_n1855_ = new_n1849_ & new_n1854_;
  assign new_n1856_ = new_n1844_ & new_n1855_;
  assign new_n1857_ = new_n1835_ & new_n1856_;
  assign new_n1858_ = new_n1813_ & new_n1857_;
  assign new_n1859_ = new_n1314_ & new_n1841_;
  assign new_n1860_ = new_n1314_ & new_n1845_;
  assign new_n1861_ = ~new_n1859_ & ~new_n1860_;
  assign new_n1862_ = new_n1314_ & new_n1847_;
  assign new_n1863_ = new_n1314_ & new_n1850_;
  assign new_n1864_ = ~new_n1862_ & ~new_n1863_;
  assign new_n1865_ = new_n1861_ & new_n1864_;
  assign new_n1866_ = new_n1314_ & new_n1852_;
  assign new_n1867_ = new_n1046_ & new_n1806_;
  assign new_n1868_ = new_n1329_ & new_n1867_;
  assign new_n1869_ = ~new_n1866_ & ~new_n1868_;
  assign new_n1870_ = new_n1053_ & new_n1818_;
  assign new_n1871_ = new_n1329_ & new_n1870_;
  assign new_n1872_ = new_n1346_ & new_n1746_;
  assign new_n1873_ = ~new_n1871_ & ~new_n1872_;
  assign new_n1874_ = new_n1869_ & new_n1873_;
  assign new_n1875_ = new_n1865_ & new_n1874_;
  assign new_n1876_ = new_n1346_ & new_n1749_;
  assign new_n1877_ = new_n1351_ & new_n1751_;
  assign new_n1878_ = ~new_n1876_ & ~new_n1877_;
  assign new_n1879_ = new_n1351_ & new_n1757_;
  assign new_n1880_ = A266 & A202;
  assign new_n1881_ = A166 & new_n1880_;
  assign new_n1882_ = new_n1248_ & new_n1881_;
  assign new_n1883_ = new_n1755_ & new_n1882_;
  assign new_n1884_ = ~new_n1879_ & ~new_n1883_;
  assign new_n1885_ = new_n1878_ & new_n1884_;
  assign new_n1886_ = new_n1346_ & new_n1755_;
  assign new_n1887_ = new_n1354_ & new_n1825_;
  assign new_n1888_ = ~new_n1886_ & ~new_n1887_;
  assign new_n1889_ = new_n1354_ & new_n1828_;
  assign new_n1890_ = new_n1366_ & new_n1831_;
  assign new_n1891_ = ~new_n1889_ & ~new_n1890_;
  assign new_n1892_ = new_n1888_ & new_n1891_;
  assign new_n1893_ = new_n1885_ & new_n1892_;
  assign new_n1894_ = new_n1875_ & new_n1893_;
  assign new_n1895_ = new_n1366_ & new_n1836_;
  assign new_n1896_ = new_n1375_ & new_n1831_;
  assign new_n1897_ = ~new_n1895_ & ~new_n1896_;
  assign new_n1898_ = new_n1375_ & new_n1836_;
  assign new_n1899_ = new_n1393_ & new_n1841_;
  assign new_n1900_ = ~new_n1898_ & ~new_n1899_;
  assign new_n1901_ = new_n1897_ & new_n1900_;
  assign new_n1902_ = new_n1393_ & new_n1845_;
  assign new_n1903_ = new_n1393_ & new_n1847_;
  assign new_n1904_ = ~new_n1902_ & ~new_n1903_;
  assign new_n1905_ = new_n1393_ & new_n1850_;
  assign new_n1906_ = new_n1393_ & new_n1852_;
  assign new_n1907_ = ~new_n1905_ & ~new_n1906_;
  assign new_n1908_ = new_n1904_ & new_n1907_;
  assign new_n1909_ = new_n1901_ & new_n1908_;
  assign new_n1910_ = new_n1405_ & new_n1841_;
  assign new_n1911_ = new_n1405_ & new_n1845_;
  assign new_n1912_ = ~new_n1910_ & ~new_n1911_;
  assign new_n1913_ = new_n1405_ & new_n1847_;
  assign new_n1914_ = new_n1405_ & new_n1850_;
  assign new_n1915_ = ~new_n1913_ & ~new_n1914_;
  assign new_n1916_ = new_n1912_ & new_n1915_;
  assign new_n1917_ = new_n1419_ & new_n1870_;
  assign new_n1918_ = new_n1405_ & new_n1852_;
  assign new_n1919_ = new_n1419_ & new_n1867_;
  assign new_n1920_ = ~new_n1918_ & ~new_n1919_;
  assign new_n1921_ = ~new_n1917_ & new_n1920_;
  assign new_n1922_ = new_n1916_ & new_n1921_;
  assign new_n1923_ = new_n1909_ & new_n1922_;
  assign new_n1924_ = new_n1894_ & new_n1923_;
  assign new_n1925_ = new_n1858_ & new_n1924_;
  assign new_n1926_ = new_n1428_ & new_n1746_;
  assign new_n1927_ = new_n1428_ & new_n1749_;
  assign new_n1928_ = ~new_n1926_ & ~new_n1927_;
  assign new_n1929_ = new_n1432_ & new_n1751_;
  assign new_n1930_ = new_n1432_ & new_n1757_;
  assign new_n1931_ = ~new_n1929_ & ~new_n1930_;
  assign new_n1932_ = new_n1928_ & new_n1931_;
  assign new_n1933_ = ~A166 & new_n1880_;
  assign new_n1934_ = new_n1353_ & new_n1933_;
  assign new_n1935_ = new_n1755_ & new_n1934_;
  assign new_n1936_ = new_n1428_ & new_n1755_;
  assign new_n1937_ = ~new_n1935_ & ~new_n1936_;
  assign new_n1938_ = new_n1435_ & new_n1608_;
  assign new_n1939_ = new_n1435_ & new_n1610_;
  assign new_n1940_ = ~new_n1938_ & ~new_n1939_;
  assign new_n1941_ = new_n1937_ & new_n1940_;
  assign new_n1942_ = new_n1932_ & new_n1941_;
  assign new_n1943_ = new_n1435_ & new_n1613_;
  assign new_n1944_ = new_n1435_ & new_n1615_;
  assign new_n1945_ = ~new_n1943_ & ~new_n1944_;
  assign new_n1946_ = new_n1435_ & new_n1619_;
  assign new_n1947_ = new_n1447_ & new_n1841_;
  assign new_n1948_ = ~new_n1946_ & ~new_n1947_;
  assign new_n1949_ = new_n1945_ & new_n1948_;
  assign new_n1950_ = new_n1447_ & new_n1845_;
  assign new_n1951_ = new_n1447_ & new_n1847_;
  assign new_n1952_ = ~new_n1950_ & ~new_n1951_;
  assign new_n1953_ = new_n1447_ & new_n1850_;
  assign new_n1954_ = new_n1447_ & new_n1852_;
  assign new_n1955_ = ~new_n1953_ & ~new_n1954_;
  assign new_n1956_ = new_n1952_ & new_n1955_;
  assign new_n1957_ = new_n1949_ & new_n1956_;
  assign new_n1958_ = new_n1942_ & new_n1957_;
  assign new_n1959_ = new_n1467_ & new_n1841_;
  assign new_n1960_ = new_n1467_ & new_n1845_;
  assign new_n1961_ = ~new_n1959_ & ~new_n1960_;
  assign new_n1962_ = new_n1467_ & new_n1847_;
  assign new_n1963_ = new_n1467_ & new_n1850_;
  assign new_n1964_ = ~new_n1962_ & ~new_n1963_;
  assign new_n1965_ = new_n1961_ & new_n1964_;
  assign new_n1966_ = new_n1467_ & new_n1852_;
  assign new_n1967_ = new_n1479_ & new_n1825_;
  assign new_n1968_ = ~new_n1966_ & ~new_n1967_;
  assign new_n1969_ = new_n1479_ & new_n1828_;
  assign new_n1970_ = new_n1488_ & new_n1746_;
  assign new_n1971_ = ~new_n1969_ & ~new_n1970_;
  assign new_n1972_ = new_n1968_ & new_n1971_;
  assign new_n1973_ = new_n1965_ & new_n1972_;
  assign new_n1974_ = new_n1488_ & new_n1749_;
  assign new_n1975_ = new_n1494_ & new_n1751_;
  assign new_n1976_ = ~new_n1974_ & ~new_n1975_;
  assign new_n1977_ = new_n1494_ & new_n1757_;
  assign new_n1978_ = A266 & A201;
  assign new_n1979_ = A200 & new_n1978_;
  assign new_n1980_ = new_n1434_ & new_n1979_;
  assign new_n1981_ = new_n1755_ & new_n1980_;
  assign new_n1982_ = ~new_n1977_ & ~new_n1981_;
  assign new_n1983_ = new_n1976_ & new_n1982_;
  assign new_n1984_ = new_n1488_ & new_n1755_;
  assign new_n1985_ = new_n1496_ & new_n1746_;
  assign new_n1986_ = ~new_n1984_ & ~new_n1985_;
  assign new_n1987_ = new_n1496_ & new_n1749_;
  assign new_n1988_ = new_n1499_ & new_n1751_;
  assign new_n1989_ = ~new_n1987_ & ~new_n1988_;
  assign new_n1990_ = new_n1986_ & new_n1989_;
  assign new_n1991_ = new_n1983_ & new_n1990_;
  assign new_n1992_ = new_n1973_ & new_n1991_;
  assign new_n1993_ = new_n1958_ & new_n1992_;
  assign new_n1994_ = new_n1499_ & new_n1757_;
  assign new_n1995_ = A199 & new_n1978_;
  assign new_n1996_ = new_n1434_ & new_n1995_;
  assign new_n1997_ = new_n1755_ & new_n1996_;
  assign new_n1998_ = ~new_n1994_ & ~new_n1997_;
  assign new_n1999_ = new_n1496_ & new_n1755_;
  assign new_n2000_ = new_n1501_ & new_n1608_;
  assign new_n2001_ = ~new_n1999_ & ~new_n2000_;
  assign new_n2002_ = new_n1998_ & new_n2001_;
  assign new_n2003_ = new_n1501_ & new_n1610_;
  assign new_n2004_ = new_n1501_ & new_n1613_;
  assign new_n2005_ = ~new_n2003_ & ~new_n2004_;
  assign new_n2006_ = new_n1501_ & new_n1615_;
  assign new_n2007_ = new_n1501_ & new_n1619_;
  assign new_n2008_ = ~new_n2006_ & ~new_n2007_;
  assign new_n2009_ = new_n2005_ & new_n2008_;
  assign new_n2010_ = new_n2002_ & new_n2009_;
  assign new_n2011_ = A202 & new_n95_;
  assign new_n2012_ = new_n1434_ & new_n2011_;
  assign new_n2013_ = new_n1791_ & new_n2012_;
  assign new_n2014_ = A202 & new_n106_;
  assign new_n2015_ = new_n1434_ & new_n2014_;
  assign new_n2016_ = new_n1791_ & new_n2015_;
  assign new_n2017_ = ~new_n2013_ & ~new_n2016_;
  assign new_n2018_ = new_n1515_ & new_n1608_;
  assign new_n2019_ = new_n1515_ & new_n1610_;
  assign new_n2020_ = ~new_n2018_ & ~new_n2019_;
  assign new_n2021_ = new_n2017_ & new_n2020_;
  assign new_n2022_ = new_n1515_ & new_n1613_;
  assign new_n2023_ = new_n1515_ & new_n1615_;
  assign new_n2024_ = ~new_n2022_ & ~new_n2023_;
  assign new_n2025_ = new_n1515_ & new_n1619_;
  assign new_n2026_ = new_n1526_ & new_n1841_;
  assign new_n2027_ = ~new_n2025_ & ~new_n2026_;
  assign new_n2028_ = new_n2024_ & new_n2027_;
  assign new_n2029_ = new_n2021_ & new_n2028_;
  assign new_n2030_ = new_n2010_ & new_n2029_;
  assign new_n2031_ = new_n1526_ & new_n1845_;
  assign new_n2032_ = new_n1526_ & new_n1847_;
  assign new_n2033_ = ~new_n2031_ & ~new_n2032_;
  assign new_n2034_ = new_n1526_ & new_n1850_;
  assign new_n2035_ = new_n1526_ & new_n1852_;
  assign new_n2036_ = ~new_n2034_ & ~new_n2035_;
  assign new_n2037_ = new_n2033_ & new_n2036_;
  assign new_n2038_ = new_n1541_ & new_n1841_;
  assign new_n2039_ = new_n1541_ & new_n1845_;
  assign new_n2040_ = ~new_n2038_ & ~new_n2039_;
  assign new_n2041_ = new_n1541_ & new_n1847_;
  assign new_n2042_ = new_n1541_ & new_n1850_;
  assign new_n2043_ = ~new_n2041_ & ~new_n2042_;
  assign new_n2044_ = new_n2040_ & new_n2043_;
  assign new_n2045_ = new_n2037_ & new_n2044_;
  assign new_n2046_ = new_n1541_ & new_n1852_;
  assign new_n2047_ = new_n1553_ & new_n1825_;
  assign new_n2048_ = ~new_n2046_ & ~new_n2047_;
  assign new_n2049_ = new_n1553_ & new_n1828_;
  assign new_n2050_ = new_n1566_ & new_n1746_;
  assign new_n2051_ = ~new_n2049_ & ~new_n2050_;
  assign new_n2052_ = new_n2048_ & new_n2051_;
  assign new_n2053_ = new_n1568_ & new_n1757_;
  assign new_n2054_ = new_n1566_ & new_n1749_;
  assign new_n2055_ = new_n1568_ & new_n1751_;
  assign new_n2056_ = ~new_n2054_ & ~new_n2055_;
  assign new_n2057_ = ~new_n2053_ & new_n2056_;
  assign new_n2058_ = new_n2052_ & new_n2057_;
  assign new_n2059_ = new_n2045_ & new_n2058_;
  assign new_n2060_ = new_n2030_ & new_n2059_;
  assign new_n2061_ = new_n1993_ & new_n2060_;
  assign new_n2062_ = new_n1925_ & new_n2061_;
  assign new_n2063_ = new_n1769_ & new_n2062_;
  assign new_n2064_ = new_n1514_ & new_n1979_;
  assign new_n2065_ = new_n1755_ & new_n2064_;
  assign new_n2066_ = new_n1566_ & new_n1755_;
  assign new_n2067_ = ~new_n2065_ & ~new_n2066_;
  assign new_n2068_ = new_n1571_ & new_n1746_;
  assign new_n2069_ = new_n1571_ & new_n1749_;
  assign new_n2070_ = ~new_n2068_ & ~new_n2069_;
  assign new_n2071_ = new_n2067_ & new_n2070_;
  assign new_n2072_ = new_n1573_ & new_n1751_;
  assign new_n2073_ = new_n1573_ & new_n1757_;
  assign new_n2074_ = ~new_n2072_ & ~new_n2073_;
  assign new_n2075_ = new_n1514_ & new_n1995_;
  assign new_n2076_ = new_n1755_ & new_n2075_;
  assign new_n2077_ = new_n1571_ & new_n1755_;
  assign new_n2078_ = ~new_n2076_ & ~new_n2077_;
  assign new_n2079_ = new_n2074_ & new_n2078_;
  assign new_n2080_ = new_n2071_ & new_n2079_;
  assign new_n2081_ = new_n1577_ & new_n1608_;
  assign new_n2082_ = new_n1577_ & new_n1610_;
  assign new_n2083_ = ~new_n2081_ & ~new_n2082_;
  assign new_n2084_ = new_n1577_ & new_n1613_;
  assign new_n2085_ = new_n1577_ & new_n1615_;
  assign new_n2086_ = ~new_n2084_ & ~new_n2085_;
  assign new_n2087_ = new_n2083_ & new_n2086_;
  assign new_n2088_ = new_n1577_ & new_n1619_;
  assign new_n2089_ = new_n1514_ & new_n2011_;
  assign new_n2090_ = new_n1791_ & new_n2089_;
  assign new_n2091_ = ~new_n2088_ & ~new_n2090_;
  assign new_n2092_ = new_n1514_ & new_n2014_;
  assign new_n2093_ = new_n1791_ & new_n2092_;
  assign new_n2094_ = A200 & ~A168;
  assign new_n2095_ = new_n943_ & new_n2094_;
  assign new_n2096_ = new_n1660_ & new_n2095_;
  assign new_n2097_ = ~new_n2093_ & ~new_n2096_;
  assign new_n2098_ = new_n2091_ & new_n2097_;
  assign new_n2099_ = new_n2087_ & new_n2098_;
  assign new_n2100_ = new_n2080_ & new_n2099_;
  assign new_n2101_ = new_n1663_ & new_n2095_;
  assign new_n2102_ = A199 & ~A168;
  assign new_n2103_ = new_n943_ & new_n2102_;
  assign new_n2104_ = new_n1660_ & new_n2103_;
  assign new_n2105_ = ~new_n2101_ & ~new_n2104_;
  assign new_n2106_ = new_n1663_ & new_n2103_;
  assign new_n2107_ = A202 & ~A168;
  assign new_n2108_ = new_n943_ & new_n2107_;
  assign new_n2109_ = new_n1608_ & new_n2108_;
  assign new_n2110_ = ~new_n2106_ & ~new_n2109_;
  assign new_n2111_ = new_n2105_ & new_n2110_;
  assign new_n2112_ = new_n1610_ & new_n2108_;
  assign new_n2113_ = new_n1613_ & new_n2108_;
  assign new_n2114_ = ~new_n2112_ & ~new_n2113_;
  assign new_n2115_ = new_n1615_ & new_n2108_;
  assign new_n2116_ = new_n1619_ & new_n2108_;
  assign new_n2117_ = ~new_n2115_ & ~new_n2116_;
  assign new_n2118_ = new_n2114_ & new_n2117_;
  assign new_n2119_ = new_n2111_ & new_n2118_;
  assign new_n2120_ = new_n1046_ & new_n1349_;
  assign new_n2121_ = A166 & A167;
  assign new_n2122_ = new_n52_ & new_n2121_;
  assign new_n2123_ = new_n2120_ & new_n2122_;
  assign new_n2124_ = new_n1053_ & new_n1653_;
  assign new_n2125_ = new_n2122_ & new_n2124_;
  assign new_n2126_ = ~new_n2123_ & ~new_n2125_;
  assign new_n2127_ = A200 & ~A166;
  assign new_n2128_ = new_n1121_ & new_n2127_;
  assign new_n2129_ = new_n1660_ & new_n2128_;
  assign new_n2130_ = new_n1663_ & new_n2128_;
  assign new_n2131_ = ~new_n2129_ & ~new_n2130_;
  assign new_n2132_ = new_n2126_ & new_n2131_;
  assign new_n2133_ = A199 & ~A166;
  assign new_n2134_ = new_n1121_ & new_n2133_;
  assign new_n2135_ = new_n1660_ & new_n2134_;
  assign new_n2136_ = new_n1663_ & new_n2134_;
  assign new_n2137_ = ~new_n2135_ & ~new_n2136_;
  assign new_n2138_ = A202 & ~A166;
  assign new_n2139_ = new_n1121_ & new_n2138_;
  assign new_n2140_ = new_n1608_ & new_n2139_;
  assign new_n2141_ = new_n1610_ & new_n2139_;
  assign new_n2142_ = ~new_n2140_ & ~new_n2141_;
  assign new_n2143_ = new_n2137_ & new_n2142_;
  assign new_n2144_ = new_n2132_ & new_n2143_;
  assign new_n2145_ = new_n2119_ & new_n2144_;
  assign new_n2146_ = new_n2100_ & new_n2145_;
  assign new_n2147_ = new_n1613_ & new_n2139_;
  assign new_n2148_ = new_n1615_ & new_n2139_;
  assign new_n2149_ = ~new_n2147_ & ~new_n2148_;
  assign new_n2150_ = new_n1619_ & new_n2139_;
  assign new_n2151_ = new_n61_ & new_n1213_;
  assign new_n2152_ = new_n1608_ & new_n2151_;
  assign new_n2153_ = ~new_n2150_ & ~new_n2152_;
  assign new_n2154_ = new_n2149_ & new_n2153_;
  assign new_n2155_ = new_n1610_ & new_n2151_;
  assign new_n2156_ = new_n1613_ & new_n2151_;
  assign new_n2157_ = ~new_n2155_ & ~new_n2156_;
  assign new_n2158_ = new_n1615_ & new_n2151_;
  assign new_n2159_ = new_n1619_ & new_n2151_;
  assign new_n2160_ = ~new_n2158_ & ~new_n2159_;
  assign new_n2161_ = new_n2157_ & new_n2160_;
  assign new_n2162_ = new_n2154_ & new_n2161_;
  assign new_n2163_ = new_n74_ & new_n1218_;
  assign new_n2164_ = new_n1841_ & new_n2163_;
  assign new_n2165_ = new_n1845_ & new_n2163_;
  assign new_n2166_ = ~new_n2164_ & ~new_n2165_;
  assign new_n2167_ = new_n1847_ & new_n2163_;
  assign new_n2168_ = new_n1850_ & new_n2163_;
  assign new_n2169_ = ~new_n2167_ & ~new_n2168_;
  assign new_n2170_ = new_n2166_ & new_n2169_;
  assign new_n2171_ = new_n1852_ & new_n2163_;
  assign new_n2172_ = new_n86_ & new_n1213_;
  assign new_n2173_ = new_n1841_ & new_n2172_;
  assign new_n2174_ = ~new_n2171_ & ~new_n2173_;
  assign new_n2175_ = new_n1845_ & new_n2172_;
  assign new_n2176_ = new_n1847_ & new_n2172_;
  assign new_n2177_ = ~new_n2175_ & ~new_n2176_;
  assign new_n2178_ = new_n2174_ & new_n2177_;
  assign new_n2179_ = new_n2170_ & new_n2178_;
  assign new_n2180_ = new_n2162_ & new_n2179_;
  assign new_n2181_ = new_n1850_ & new_n2172_;
  assign new_n2182_ = new_n1852_ & new_n2172_;
  assign new_n2183_ = ~new_n2181_ & ~new_n2182_;
  assign new_n2184_ = new_n34_ & new_n1218_;
  assign new_n2185_ = new_n1825_ & new_n2184_;
  assign new_n2186_ = new_n1828_ & new_n2184_;
  assign new_n2187_ = ~new_n2185_ & ~new_n2186_;
  assign new_n2188_ = new_n2183_ & new_n2187_;
  assign new_n2189_ = new_n521_ & new_n1793_;
  assign new_n2190_ = new_n1746_ & new_n2189_;
  assign new_n2191_ = new_n1749_ & new_n2189_;
  assign new_n2192_ = ~new_n2190_ & ~new_n2191_;
  assign new_n2193_ = new_n769_ & new_n1793_;
  assign new_n2194_ = new_n1751_ & new_n2193_;
  assign new_n2195_ = new_n1757_ & new_n2193_;
  assign new_n2196_ = ~new_n2194_ & ~new_n2195_;
  assign new_n2197_ = new_n2192_ & new_n2196_;
  assign new_n2198_ = new_n2188_ & new_n2197_;
  assign new_n2199_ = new_n1793_ & new_n1978_;
  assign new_n2200_ = new_n1755_ & new_n2199_;
  assign new_n2201_ = new_n1755_ & new_n2189_;
  assign new_n2202_ = ~new_n2200_ & ~new_n2201_;
  assign new_n2203_ = new_n521_ & new_n1218_;
  assign new_n2204_ = new_n1746_ & new_n2203_;
  assign new_n2205_ = new_n1749_ & new_n2203_;
  assign new_n2206_ = ~new_n2204_ & ~new_n2205_;
  assign new_n2207_ = new_n2202_ & new_n2206_;
  assign new_n2208_ = new_n1218_ & new_n1978_;
  assign new_n2209_ = new_n1755_ & new_n2208_;
  assign new_n2210_ = new_n769_ & new_n1218_;
  assign new_n2211_ = new_n1751_ & new_n2210_;
  assign new_n2212_ = new_n1757_ & new_n2210_;
  assign new_n2213_ = ~new_n2211_ & ~new_n2212_;
  assign new_n2214_ = ~new_n2209_ & new_n2213_;
  assign new_n2215_ = new_n2207_ & new_n2214_;
  assign new_n2216_ = new_n2198_ & new_n2215_;
  assign new_n2217_ = new_n2180_ & new_n2216_;
  assign new_n2218_ = new_n2146_ & new_n2217_;
  assign new_n2219_ = new_n1755_ & new_n2203_;
  assign new_n2220_ = new_n125_ & new_n1243_;
  assign new_n2221_ = new_n1608_ & new_n2220_;
  assign new_n2222_ = ~new_n2219_ & ~new_n2221_;
  assign new_n2223_ = new_n1610_ & new_n2220_;
  assign new_n2224_ = new_n1613_ & new_n2220_;
  assign new_n2225_ = ~new_n2223_ & ~new_n2224_;
  assign new_n2226_ = new_n2222_ & new_n2225_;
  assign new_n2227_ = new_n1615_ & new_n2220_;
  assign new_n2228_ = new_n1619_ & new_n2220_;
  assign new_n2229_ = ~new_n2227_ & ~new_n2228_;
  assign new_n2230_ = A202 & A169;
  assign new_n2231_ = new_n95_ & new_n2230_;
  assign new_n2232_ = new_n1791_ & new_n2231_;
  assign new_n2233_ = new_n106_ & new_n2230_;
  assign new_n2234_ = new_n1791_ & new_n2233_;
  assign new_n2235_ = ~new_n2232_ & ~new_n2234_;
  assign new_n2236_ = new_n2229_ & new_n2235_;
  assign new_n2237_ = new_n2226_ & new_n2236_;
  assign new_n2238_ = A268 & A201;
  assign new_n2239_ = new_n439_ & new_n2238_;
  assign new_n2240_ = new_n1068_ & new_n1248_;
  assign new_n2241_ = new_n2239_ & new_n2240_;
  assign new_n2242_ = new_n443_ & new_n2238_;
  assign new_n2243_ = new_n2240_ & new_n2242_;
  assign new_n2244_ = ~new_n2241_ & ~new_n2243_;
  assign new_n2245_ = new_n35_ & new_n1248_;
  assign new_n2246_ = new_n2239_ & new_n2245_;
  assign new_n2247_ = new_n2242_ & new_n2245_;
  assign new_n2248_ = ~new_n2246_ & ~new_n2247_;
  assign new_n2249_ = new_n2244_ & new_n2248_;
  assign new_n2250_ = new_n1106_ & new_n1248_;
  assign new_n2251_ = new_n1841_ & new_n2250_;
  assign new_n2252_ = new_n1845_ & new_n2250_;
  assign new_n2253_ = ~new_n2251_ & ~new_n2252_;
  assign new_n2254_ = new_n1847_ & new_n2250_;
  assign new_n2255_ = new_n1850_ & new_n2250_;
  assign new_n2256_ = ~new_n2254_ & ~new_n2255_;
  assign new_n2257_ = new_n2253_ & new_n2256_;
  assign new_n2258_ = new_n2249_ & new_n2257_;
  assign new_n2259_ = new_n2237_ & new_n2258_;
  assign new_n2260_ = new_n1852_ & new_n2250_;
  assign new_n2261_ = new_n1353_ & new_n2127_;
  assign new_n2262_ = new_n2239_ & new_n2261_;
  assign new_n2263_ = ~new_n2260_ & ~new_n2262_;
  assign new_n2264_ = new_n2242_ & new_n2261_;
  assign new_n2265_ = new_n1353_ & new_n2133_;
  assign new_n2266_ = new_n2239_ & new_n2265_;
  assign new_n2267_ = ~new_n2264_ & ~new_n2266_;
  assign new_n2268_ = new_n2263_ & new_n2267_;
  assign new_n2269_ = new_n2242_ & new_n2265_;
  assign new_n2270_ = new_n1353_ & new_n2138_;
  assign new_n2271_ = new_n1841_ & new_n2270_;
  assign new_n2272_ = ~new_n2269_ & ~new_n2271_;
  assign new_n2273_ = new_n1845_ & new_n2270_;
  assign new_n2274_ = new_n1847_ & new_n2270_;
  assign new_n2275_ = ~new_n2273_ & ~new_n2274_;
  assign new_n2276_ = new_n2272_ & new_n2275_;
  assign new_n2277_ = new_n2268_ & new_n2276_;
  assign new_n2278_ = new_n1850_ & new_n2270_;
  assign new_n2279_ = new_n1852_ & new_n2270_;
  assign new_n2280_ = ~new_n2278_ & ~new_n2279_;
  assign new_n2281_ = new_n190_ & new_n1434_;
  assign new_n2282_ = new_n1825_ & new_n2281_;
  assign new_n2283_ = new_n1828_ & new_n2281_;
  assign new_n2284_ = ~new_n2282_ & ~new_n2283_;
  assign new_n2285_ = new_n2280_ & new_n2284_;
  assign new_n2286_ = new_n208_ & new_n1434_;
  assign new_n2287_ = new_n1831_ & new_n2286_;
  assign new_n2288_ = new_n1836_ & new_n2286_;
  assign new_n2289_ = ~new_n2287_ & ~new_n2288_;
  assign new_n2290_ = new_n240_ & new_n1434_;
  assign new_n2291_ = new_n1831_ & new_n2290_;
  assign new_n2292_ = new_n1836_ & new_n2290_;
  assign new_n2293_ = ~new_n2291_ & ~new_n2292_;
  assign new_n2294_ = new_n2289_ & new_n2293_;
  assign new_n2295_ = new_n2285_ & new_n2294_;
  assign new_n2296_ = new_n2277_ & new_n2295_;
  assign new_n2297_ = new_n2259_ & new_n2296_;
  assign new_n2298_ = new_n279_ & new_n1434_;
  assign new_n2299_ = new_n1841_ & new_n2298_;
  assign new_n2300_ = new_n1845_ & new_n2298_;
  assign new_n2301_ = ~new_n2299_ & ~new_n2300_;
  assign new_n2302_ = new_n1847_ & new_n2298_;
  assign new_n2303_ = new_n1850_ & new_n2298_;
  assign new_n2304_ = ~new_n2302_ & ~new_n2303_;
  assign new_n2305_ = new_n2301_ & new_n2304_;
  assign new_n2306_ = new_n1852_ & new_n2298_;
  assign new_n2307_ = new_n285_ & new_n1434_;
  assign new_n2308_ = new_n1841_ & new_n2307_;
  assign new_n2309_ = ~new_n2306_ & ~new_n2308_;
  assign new_n2310_ = new_n1845_ & new_n2307_;
  assign new_n2311_ = new_n1847_ & new_n2307_;
  assign new_n2312_ = ~new_n2310_ & ~new_n2311_;
  assign new_n2313_ = new_n2309_ & new_n2312_;
  assign new_n2314_ = new_n2305_ & new_n2313_;
  assign new_n2315_ = new_n1850_ & new_n2307_;
  assign new_n2316_ = new_n1852_ & new_n2307_;
  assign new_n2317_ = ~new_n2315_ & ~new_n2316_;
  assign new_n2318_ = new_n49_ & new_n1434_;
  assign new_n2319_ = new_n1867_ & new_n2318_;
  assign new_n2320_ = new_n1870_ & new_n2318_;
  assign new_n2321_ = ~new_n2319_ & ~new_n2320_;
  assign new_n2322_ = new_n2317_ & new_n2321_;
  assign new_n2323_ = new_n631_ & new_n1434_;
  assign new_n2324_ = new_n1746_ & new_n2323_;
  assign new_n2325_ = new_n1749_ & new_n2323_;
  assign new_n2326_ = ~new_n2324_ & ~new_n2325_;
  assign new_n2327_ = new_n1349_ & new_n1434_;
  assign new_n2328_ = new_n1751_ & new_n2327_;
  assign new_n2329_ = new_n1757_ & new_n2327_;
  assign new_n2330_ = ~new_n2328_ & ~new_n2329_;
  assign new_n2331_ = new_n2326_ & new_n2330_;
  assign new_n2332_ = new_n2322_ & new_n2331_;
  assign new_n2333_ = new_n2314_ & new_n2332_;
  assign new_n2334_ = new_n1434_ & new_n1880_;
  assign new_n2335_ = new_n1755_ & new_n2334_;
  assign new_n2336_ = new_n1755_ & new_n2323_;
  assign new_n2337_ = ~new_n2335_ & ~new_n2336_;
  assign new_n2338_ = new_n190_ & new_n1514_;
  assign new_n2339_ = new_n1825_ & new_n2338_;
  assign new_n2340_ = new_n1828_ & new_n2338_;
  assign new_n2341_ = ~new_n2339_ & ~new_n2340_;
  assign new_n2342_ = new_n2337_ & new_n2341_;
  assign new_n2343_ = new_n208_ & new_n1514_;
  assign new_n2344_ = new_n1831_ & new_n2343_;
  assign new_n2345_ = new_n1836_ & new_n2343_;
  assign new_n2346_ = ~new_n2344_ & ~new_n2345_;
  assign new_n2347_ = new_n240_ & new_n1514_;
  assign new_n2348_ = new_n1831_ & new_n2347_;
  assign new_n2349_ = new_n1836_ & new_n2347_;
  assign new_n2350_ = ~new_n2348_ & ~new_n2349_;
  assign new_n2351_ = new_n2346_ & new_n2350_;
  assign new_n2352_ = new_n2342_ & new_n2351_;
  assign new_n2353_ = new_n279_ & new_n1514_;
  assign new_n2354_ = new_n1841_ & new_n2353_;
  assign new_n2355_ = new_n1845_ & new_n2353_;
  assign new_n2356_ = ~new_n2354_ & ~new_n2355_;
  assign new_n2357_ = new_n1847_ & new_n2353_;
  assign new_n2358_ = new_n1850_ & new_n2353_;
  assign new_n2359_ = ~new_n2357_ & ~new_n2358_;
  assign new_n2360_ = new_n2356_ & new_n2359_;
  assign new_n2361_ = new_n285_ & new_n1514_;
  assign new_n2362_ = new_n1845_ & new_n2361_;
  assign new_n2363_ = new_n1852_ & new_n2353_;
  assign new_n2364_ = new_n1841_ & new_n2361_;
  assign new_n2365_ = ~new_n2363_ & ~new_n2364_;
  assign new_n2366_ = ~new_n2362_ & new_n2365_;
  assign new_n2367_ = new_n2360_ & new_n2366_;
  assign new_n2368_ = new_n2352_ & new_n2367_;
  assign new_n2369_ = new_n2333_ & new_n2368_;
  assign new_n2370_ = new_n2297_ & new_n2369_;
  assign new_n2371_ = new_n2218_ & new_n2370_;
  assign new_n2372_ = new_n1847_ & new_n2361_;
  assign new_n2373_ = new_n1850_ & new_n2361_;
  assign new_n2374_ = ~new_n2372_ & ~new_n2373_;
  assign new_n2375_ = new_n1852_ & new_n2361_;
  assign new_n2376_ = new_n49_ & new_n1514_;
  assign new_n2377_ = new_n1867_ & new_n2376_;
  assign new_n2378_ = ~new_n2375_ & ~new_n2377_;
  assign new_n2379_ = new_n2374_ & new_n2378_;
  assign new_n2380_ = new_n1870_ & new_n2376_;
  assign new_n2381_ = new_n631_ & new_n1514_;
  assign new_n2382_ = new_n1746_ & new_n2381_;
  assign new_n2383_ = ~new_n2380_ & ~new_n2382_;
  assign new_n2384_ = new_n1749_ & new_n2381_;
  assign new_n2385_ = new_n1349_ & new_n1514_;
  assign new_n2386_ = new_n1751_ & new_n2385_;
  assign new_n2387_ = ~new_n2384_ & ~new_n2386_;
  assign new_n2388_ = new_n2383_ & new_n2387_;
  assign new_n2389_ = new_n2379_ & new_n2388_;
  assign new_n2390_ = new_n1757_ & new_n2385_;
  assign new_n2391_ = new_n1514_ & new_n1880_;
  assign new_n2392_ = new_n1755_ & new_n2391_;
  assign new_n2393_ = ~new_n2390_ & ~new_n2392_;
  assign new_n2394_ = new_n1755_ & new_n2381_;
  assign new_n2395_ = new_n205_ & new_n562_;
  assign new_n2396_ = new_n2108_ & new_n2395_;
  assign new_n2397_ = ~new_n2394_ & ~new_n2396_;
  assign new_n2398_ = new_n2393_ & new_n2397_;
  assign new_n2399_ = new_n216_ & new_n1052_;
  assign new_n2400_ = new_n2108_ & new_n2399_;
  assign new_n2401_ = new_n2139_ & new_n2395_;
  assign new_n2402_ = ~new_n2400_ & ~new_n2401_;
  assign new_n2403_ = new_n2139_ & new_n2399_;
  assign new_n2404_ = new_n2151_ & new_n2395_;
  assign new_n2405_ = ~new_n2403_ & ~new_n2404_;
  assign new_n2406_ = new_n2402_ & new_n2405_;
  assign new_n2407_ = new_n2398_ & new_n2406_;
  assign new_n2408_ = new_n2389_ & new_n2407_;
  assign new_n2409_ = new_n2151_ & new_n2399_;
  assign new_n2410_ = ~A298 & A268;
  assign new_n2411_ = new_n92_ & new_n2410_;
  assign new_n2412_ = new_n2163_ & new_n2411_;
  assign new_n2413_ = ~new_n2409_ & ~new_n2412_;
  assign new_n2414_ = ~A300 & A268;
  assign new_n2415_ = new_n99_ & new_n2414_;
  assign new_n2416_ = new_n2163_ & new_n2415_;
  assign new_n2417_ = new_n2172_ & new_n2411_;
  assign new_n2418_ = ~new_n2416_ & ~new_n2417_;
  assign new_n2419_ = new_n2413_ & new_n2418_;
  assign new_n2420_ = new_n2172_ & new_n2415_;
  assign new_n2421_ = new_n256_ & new_n2199_;
  assign new_n2422_ = ~new_n2420_ & ~new_n2421_;
  assign new_n2423_ = new_n264_ & new_n2199_;
  assign new_n2424_ = new_n256_ & new_n2189_;
  assign new_n2425_ = ~new_n2423_ & ~new_n2424_;
  assign new_n2426_ = new_n2422_ & new_n2425_;
  assign new_n2427_ = new_n2419_ & new_n2426_;
  assign new_n2428_ = new_n264_ & new_n2189_;
  assign new_n2429_ = new_n1793_ & new_n2238_;
  assign new_n2430_ = new_n29_ & new_n2429_;
  assign new_n2431_ = ~new_n2428_ & ~new_n2430_;
  assign new_n2432_ = new_n256_ & new_n2208_;
  assign new_n2433_ = new_n264_ & new_n2208_;
  assign new_n2434_ = ~new_n2432_ & ~new_n2433_;
  assign new_n2435_ = new_n2431_ & new_n2434_;
  assign new_n2436_ = new_n256_ & new_n2203_;
  assign new_n2437_ = new_n264_ & new_n2203_;
  assign new_n2438_ = ~new_n2436_ & ~new_n2437_;
  assign new_n2439_ = new_n1218_ & new_n2238_;
  assign new_n2440_ = new_n29_ & new_n2439_;
  assign new_n2441_ = new_n2220_ & new_n2395_;
  assign new_n2442_ = ~new_n2440_ & ~new_n2441_;
  assign new_n2443_ = new_n2438_ & new_n2442_;
  assign new_n2444_ = new_n2435_ & new_n2443_;
  assign new_n2445_ = new_n2427_ & new_n2444_;
  assign new_n2446_ = new_n2408_ & new_n2445_;
  assign new_n2447_ = new_n2220_ & new_n2399_;
  assign new_n2448_ = new_n94_ & new_n2231_;
  assign new_n2449_ = ~new_n2447_ & ~new_n2448_;
  assign new_n2450_ = new_n101_ & new_n2231_;
  assign new_n2451_ = new_n94_ & new_n2233_;
  assign new_n2452_ = ~new_n2450_ & ~new_n2451_;
  assign new_n2453_ = new_n2449_ & new_n2452_;
  assign new_n2454_ = new_n101_ & new_n2233_;
  assign new_n2455_ = new_n113_ & new_n2230_;
  assign new_n2456_ = new_n29_ & new_n2455_;
  assign new_n2457_ = ~new_n2454_ & ~new_n2456_;
  assign new_n2458_ = new_n117_ & new_n2230_;
  assign new_n2459_ = new_n29_ & new_n2458_;
  assign new_n2460_ = new_n2250_ & new_n2411_;
  assign new_n2461_ = ~new_n2459_ & ~new_n2460_;
  assign new_n2462_ = new_n2457_ & new_n2461_;
  assign new_n2463_ = new_n2453_ & new_n2462_;
  assign new_n2464_ = new_n2250_ & new_n2415_;
  assign new_n2465_ = new_n2270_ & new_n2411_;
  assign new_n2466_ = ~new_n2464_ & ~new_n2465_;
  assign new_n2467_ = new_n2270_ & new_n2415_;
  assign new_n2468_ = new_n2298_ & new_n2411_;
  assign new_n2469_ = ~new_n2467_ & ~new_n2468_;
  assign new_n2470_ = new_n2466_ & new_n2469_;
  assign new_n2471_ = new_n2298_ & new_n2415_;
  assign new_n2472_ = new_n2307_ & new_n2411_;
  assign new_n2473_ = ~new_n2471_ & ~new_n2472_;
  assign new_n2474_ = new_n2307_ & new_n2415_;
  assign new_n2475_ = new_n256_ & new_n2334_;
  assign new_n2476_ = ~new_n2474_ & ~new_n2475_;
  assign new_n2477_ = new_n2473_ & new_n2476_;
  assign new_n2478_ = new_n2470_ & new_n2477_;
  assign new_n2479_ = new_n2463_ & new_n2478_;
  assign new_n2480_ = new_n264_ & new_n2334_;
  assign new_n2481_ = new_n256_ & new_n2323_;
  assign new_n2482_ = ~new_n2480_ & ~new_n2481_;
  assign new_n2483_ = new_n264_ & new_n2323_;
  assign new_n2484_ = A268 & A202;
  assign new_n2485_ = new_n1434_ & new_n2484_;
  assign new_n2486_ = new_n29_ & new_n2485_;
  assign new_n2487_ = ~new_n2483_ & ~new_n2486_;
  assign new_n2488_ = new_n2482_ & new_n2487_;
  assign new_n2489_ = new_n2353_ & new_n2411_;
  assign new_n2490_ = new_n2353_ & new_n2415_;
  assign new_n2491_ = ~new_n2489_ & ~new_n2490_;
  assign new_n2492_ = new_n2361_ & new_n2411_;
  assign new_n2493_ = new_n2361_ & new_n2415_;
  assign new_n2494_ = ~new_n2492_ & ~new_n2493_;
  assign new_n2495_ = new_n2491_ & new_n2494_;
  assign new_n2496_ = new_n2488_ & new_n2495_;
  assign new_n2497_ = new_n256_ & new_n2391_;
  assign new_n2498_ = new_n264_ & new_n2391_;
  assign new_n2499_ = ~new_n2497_ & ~new_n2498_;
  assign new_n2500_ = new_n256_ & new_n2381_;
  assign new_n2501_ = new_n264_ & new_n2381_;
  assign new_n2502_ = ~new_n2500_ & ~new_n2501_;
  assign new_n2503_ = new_n2499_ & new_n2502_;
  assign new_n2504_ = A169 & new_n279_;
  assign new_n2505_ = new_n2415_ & new_n2504_;
  assign new_n2506_ = new_n1514_ & new_n2484_;
  assign new_n2507_ = new_n29_ & new_n2506_;
  assign new_n2508_ = new_n2411_ & new_n2504_;
  assign new_n2509_ = ~new_n2507_ & ~new_n2508_;
  assign new_n2510_ = ~new_n2505_ & new_n2509_;
  assign new_n2511_ = new_n2503_ & new_n2510_;
  assign new_n2512_ = new_n2496_ & new_n2511_;
  assign new_n2513_ = new_n2479_ & new_n2512_;
  assign new_n2514_ = new_n2446_ & new_n2513_;
  assign new_n2515_ = A169 & new_n285_;
  assign new_n2516_ = new_n2411_ & new_n2515_;
  assign new_n2517_ = new_n2415_ & new_n2515_;
  assign new_n2518_ = ~new_n2516_ & ~new_n2517_;
  assign new_n2519_ = A169 & new_n1880_;
  assign new_n2520_ = new_n256_ & new_n2519_;
  assign new_n2521_ = new_n264_ & new_n2519_;
  assign new_n2522_ = ~new_n2520_ & ~new_n2521_;
  assign new_n2523_ = new_n2518_ & new_n2522_;
  assign new_n2524_ = A169 & new_n631_;
  assign new_n2525_ = new_n256_ & new_n2524_;
  assign new_n2526_ = new_n264_ & new_n2524_;
  assign new_n2527_ = ~new_n2525_ & ~new_n2526_;
  assign new_n2528_ = A169 & new_n2484_;
  assign new_n2529_ = new_n29_ & new_n2528_;
  assign new_n2530_ = A202 & A167;
  assign new_n2531_ = A168 & new_n2530_;
  assign new_n2532_ = new_n2411_ & new_n2531_;
  assign new_n2533_ = ~new_n2529_ & ~new_n2532_;
  assign new_n2534_ = new_n2527_ & new_n2533_;
  assign new_n2535_ = new_n2523_ & new_n2534_;
  assign new_n2536_ = new_n2415_ & new_n2531_;
  assign new_n2537_ = A168 & new_n1106_;
  assign new_n2538_ = new_n2411_ & new_n2537_;
  assign new_n2539_ = ~new_n2536_ & ~new_n2538_;
  assign new_n2540_ = new_n2415_ & new_n2537_;
  assign new_n2541_ = new_n439_ & new_n2528_;
  assign new_n2542_ = ~new_n2540_ & ~new_n2541_;
  assign new_n2543_ = new_n2539_ & new_n2542_;
  assign new_n2544_ = new_n443_ & new_n2528_;
  assign new_n2545_ = A236 & ~A233;
  assign new_n2546_ = A232 & new_n2545_;
  assign new_n2547_ = new_n140_ & new_n2546_;
  assign new_n2548_ = ~new_n2544_ & ~new_n2547_;
  assign new_n2549_ = A236 & A233;
  assign new_n2550_ = ~A232 & new_n2549_;
  assign new_n2551_ = new_n140_ & new_n2550_;
  assign new_n2552_ = new_n146_ & new_n2546_;
  assign new_n2553_ = ~new_n2551_ & ~new_n2552_;
  assign new_n2554_ = new_n2548_ & new_n2553_;
  assign new_n2555_ = new_n2543_ & new_n2554_;
  assign new_n2556_ = new_n2535_ & new_n2555_;
  assign new_n2557_ = new_n146_ & new_n2550_;
  assign new_n2558_ = new_n158_ & new_n2546_;
  assign new_n2559_ = ~new_n2557_ & ~new_n2558_;
  assign new_n2560_ = new_n158_ & new_n2550_;
  assign new_n2561_ = new_n164_ & new_n2546_;
  assign new_n2562_ = ~new_n2560_ & ~new_n2561_;
  assign new_n2563_ = new_n2559_ & new_n2562_;
  assign new_n2564_ = new_n164_ & new_n2550_;
  assign new_n2565_ = A234 & A233;
  assign new_n2566_ = A166 & new_n2565_;
  assign new_n2567_ = new_n1248_ & new_n2566_;
  assign new_n2568_ = ~new_n2564_ & ~new_n2567_;
  assign new_n2569_ = A234 & A232;
  assign new_n2570_ = A166 & new_n2569_;
  assign new_n2571_ = new_n1248_ & new_n2570_;
  assign new_n2572_ = ~A166 & new_n2565_;
  assign new_n2573_ = new_n1353_ & new_n2572_;
  assign new_n2574_ = ~new_n2571_ & ~new_n2573_;
  assign new_n2575_ = new_n2568_ & new_n2574_;
  assign new_n2576_ = new_n2563_ & new_n2575_;
  assign new_n2577_ = ~A166 & new_n2569_;
  assign new_n2578_ = new_n1353_ & new_n2577_;
  assign new_n2579_ = new_n1434_ & new_n2546_;
  assign new_n2580_ = ~new_n2578_ & ~new_n2579_;
  assign new_n2581_ = new_n1434_ & new_n2550_;
  assign new_n2582_ = new_n1514_ & new_n2546_;
  assign new_n2583_ = ~new_n2581_ & ~new_n2582_;
  assign new_n2584_ = new_n2580_ & new_n2583_;
  assign new_n2585_ = new_n1514_ & new_n2550_;
  assign new_n2586_ = A203 & new_n2565_;
  assign new_n2587_ = new_n208_ & new_n2586_;
  assign new_n2588_ = ~new_n2585_ & ~new_n2587_;
  assign new_n2589_ = A203 & new_n2569_;
  assign new_n2590_ = new_n208_ & new_n2589_;
  assign new_n2591_ = new_n240_ & new_n2586_;
  assign new_n2592_ = ~new_n2590_ & ~new_n2591_;
  assign new_n2593_ = new_n2588_ & new_n2592_;
  assign new_n2594_ = new_n2584_ & new_n2593_;
  assign new_n2595_ = new_n2576_ & new_n2594_;
  assign new_n2596_ = new_n2556_ & new_n2595_;
  assign new_n2597_ = new_n240_ & new_n2589_;
  assign new_n2598_ = new_n279_ & new_n2546_;
  assign new_n2599_ = ~new_n2597_ & ~new_n2598_;
  assign new_n2600_ = new_n279_ & new_n2550_;
  assign new_n2601_ = new_n285_ & new_n2546_;
  assign new_n2602_ = ~new_n2600_ & ~new_n2601_;
  assign new_n2603_ = new_n2599_ & new_n2602_;
  assign new_n2604_ = new_n285_ & new_n2550_;
  assign new_n2605_ = A232 & A169;
  assign new_n2606_ = new_n2545_ & new_n2605_;
  assign new_n2607_ = ~new_n2604_ & ~new_n2606_;
  assign new_n2608_ = ~A232 & A169;
  assign new_n2609_ = new_n2549_ & new_n2608_;
  assign new_n2610_ = A235 & A166;
  assign new_n2611_ = new_n1248_ & new_n2610_;
  assign new_n2612_ = ~new_n2609_ & ~new_n2611_;
  assign new_n2613_ = new_n2607_ & new_n2612_;
  assign new_n2614_ = new_n2603_ & new_n2613_;
  assign new_n2615_ = A235 & ~A166;
  assign new_n2616_ = new_n1353_ & new_n2615_;
  assign new_n2617_ = new_n1434_ & new_n2565_;
  assign new_n2618_ = ~new_n2616_ & ~new_n2617_;
  assign new_n2619_ = new_n1434_ & new_n2569_;
  assign new_n2620_ = new_n1514_ & new_n2565_;
  assign new_n2621_ = ~new_n2619_ & ~new_n2620_;
  assign new_n2622_ = new_n2618_ & new_n2621_;
  assign new_n2623_ = new_n1514_ & new_n2569_;
  assign new_n2624_ = A235 & A203;
  assign new_n2625_ = new_n208_ & new_n2624_;
  assign new_n2626_ = ~new_n2623_ & ~new_n2625_;
  assign new_n2627_ = new_n240_ & new_n2624_;
  assign new_n2628_ = new_n279_ & new_n2565_;
  assign new_n2629_ = ~new_n2627_ & ~new_n2628_;
  assign new_n2630_ = new_n2626_ & new_n2629_;
  assign new_n2631_ = new_n2622_ & new_n2630_;
  assign new_n2632_ = new_n2614_ & new_n2631_;
  assign new_n2633_ = new_n279_ & new_n2569_;
  assign new_n2634_ = new_n285_ & new_n2565_;
  assign new_n2635_ = ~new_n2633_ & ~new_n2634_;
  assign new_n2636_ = new_n285_ & new_n2569_;
  assign new_n2637_ = A232 & A202;
  assign new_n2638_ = new_n2545_ & new_n2637_;
  assign new_n2639_ = ~new_n2636_ & ~new_n2638_;
  assign new_n2640_ = new_n2635_ & new_n2639_;
  assign new_n2641_ = ~A232 & A202;
  assign new_n2642_ = new_n2549_ & new_n2641_;
  assign new_n2643_ = A169 & new_n2565_;
  assign new_n2644_ = ~new_n2642_ & ~new_n2643_;
  assign new_n2645_ = A169 & new_n2569_;
  assign new_n2646_ = A235 & A167;
  assign new_n2647_ = A168 & new_n2646_;
  assign new_n2648_ = ~new_n2645_ & ~new_n2647_;
  assign new_n2649_ = new_n2644_ & new_n2648_;
  assign new_n2650_ = new_n2640_ & new_n2649_;
  assign new_n2651_ = A168 & new_n2610_;
  assign new_n2652_ = A235 & A201;
  assign new_n2653_ = A200 & new_n2652_;
  assign new_n2654_ = ~new_n2651_ & ~new_n2653_;
  assign new_n2655_ = A199 & new_n2652_;
  assign new_n2656_ = A202 & new_n2565_;
  assign new_n2657_ = ~new_n2655_ & ~new_n2656_;
  assign new_n2658_ = new_n2654_ & new_n2657_;
  assign new_n2659_ = A235 & A202;
  assign new_n2660_ = A202 & new_n2569_;
  assign new_n2661_ = A235 & A169;
  assign new_n2662_ = ~new_n2660_ & ~new_n2661_;
  assign new_n2663_ = ~new_n2659_ & new_n2662_;
  assign new_n2664_ = new_n2658_ & new_n2663_;
  assign new_n2665_ = new_n2650_ & new_n2664_;
  assign new_n2666_ = new_n2632_ & new_n2665_;
  assign new_n2667_ = new_n2596_ & new_n2666_;
  assign new_n2668_ = new_n2514_ & new_n2667_;
  assign new_n2669_ = new_n2371_ & new_n2668_;
  assign new_n2670_ = new_n2063_ & new_n2669_;
  assign A73 = ~new_n1459_ | ~new_n2670_;
endmodule


