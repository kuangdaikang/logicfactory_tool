// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:40 2022

module intb  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    \v15.0 , \v15.1 , \v15.2 , \v15.3 , \v15.4 , \v15.5 , \v15.6   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14;
  output \v15.0 , \v15.1 , \v15.2 , \v15.3 , \v15.4 , \v15.5 , \v15.6 ;
  wire new_n23_, new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_,
    new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_,
    new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_,
    new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_,
    new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_,
    new_n58_, new_n59_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_;
  assign new_n23_ = v7 & ~v11;
  assign new_n24_ = v6 & ~v10;
  assign new_n25_ = v5 & ~v9;
  assign new_n26_ = v8 & ~new_n25_;
  assign new_n27_ = ~v4 & v9;
  assign new_n28_ = ~new_n26_ & ~new_n27_;
  assign new_n29_ = ~new_n24_ & ~new_n28_;
  assign new_n30_ = ~v5 & v10;
  assign new_n31_ = ~v4 & new_n30_;
  assign new_n32_ = ~new_n29_ & ~new_n31_;
  assign new_n33_ = ~new_n23_ & ~new_n32_;
  assign new_n34_ = ~v4 & ~v5;
  assign new_n35_ = ~v6 & v11;
  assign new_n36_ = new_n34_ & new_n35_;
  assign new_n37_ = v2 & ~new_n36_;
  assign new_n38_ = ~new_n33_ & new_n37_;
  assign new_n39_ = ~v3 & ~new_n38_;
  assign new_n40_ = ~v2 & ~v11;
  assign new_n41_ = v7 & ~new_n40_;
  assign new_n42_ = ~v6 & ~new_n41_;
  assign new_n43_ = v7 & v11;
  assign new_n44_ = ~v10 & ~new_n43_;
  assign new_n45_ = ~v2 & new_n44_;
  assign new_n46_ = ~new_n42_ & ~new_n45_;
  assign new_n47_ = ~v5 & ~new_n46_;
  assign new_n48_ = v6 & v10;
  assign new_n49_ = ~new_n43_ & ~new_n48_;
  assign new_n50_ = ~v9 & new_n49_;
  assign new_n51_ = ~v2 & new_n50_;
  assign new_n52_ = ~new_n47_ & ~new_n51_;
  assign new_n53_ = ~v4 & ~new_n52_;
  assign new_n54_ = v5 & v9;
  assign new_n55_ = ~new_n48_ & ~new_n54_;
  assign new_n56_ = ~new_n43_ & new_n55_;
  assign new_n57_ = ~v8 & new_n56_;
  assign new_n58_ = ~v2 & new_n57_;
  assign new_n59_ = ~new_n53_ & ~new_n58_;
  assign \v15.0  = new_n39_ | ~new_n59_;
  assign new_n61_ = ~v9 & v10;
  assign new_n62_ = v5 & new_n61_;
  assign new_n63_ = ~new_n24_ & ~new_n62_;
  assign new_n64_ = v2 & ~new_n63_;
  assign new_n65_ = ~v6 & ~v10;
  assign new_n66_ = ~v5 & ~v9;
  assign new_n67_ = ~v4 & ~v8;
  assign new_n68_ = ~new_n66_ & ~new_n67_;
  assign new_n69_ = v3 & new_n54_;
  assign new_n70_ = ~new_n68_ & ~new_n69_;
  assign new_n71_ = ~new_n65_ & ~new_n70_;
  assign new_n72_ = v3 & new_n48_;
  assign new_n73_ = ~new_n71_ & ~new_n72_;
  assign new_n74_ = ~new_n64_ & new_n73_;
  assign new_n75_ = v11 & ~new_n74_;
  assign new_n76_ = v8 & ~new_n66_;
  assign new_n77_ = v4 & v9;
  assign new_n78_ = ~new_n76_ & ~new_n77_;
  assign new_n79_ = ~new_n65_ & ~new_n78_;
  assign new_n80_ = v3 & v9;
  assign new_n81_ = ~v4 & ~new_n80_;
  assign new_n82_ = v10 & ~new_n81_;
  assign new_n83_ = v5 & new_n82_;
  assign new_n84_ = ~new_n79_ & ~new_n83_;
  assign new_n85_ = v7 & ~new_n84_;
  assign new_n86_ = ~v1 & ~new_n85_;
  assign new_n87_ = ~new_n75_ & new_n86_;
  assign new_n88_ = v0 & ~new_n87_;
  assign new_n89_ = v6 & v7;
  assign new_n90_ = ~v10 & ~v11;
  assign new_n91_ = v1 & new_n90_;
  assign new_n92_ = ~new_n89_ & ~new_n91_;
  assign new_n93_ = v2 & ~v9;
  assign new_n94_ = ~new_n80_ & ~new_n93_;
  assign new_n95_ = ~v4 & new_n94_;
  assign new_n96_ = ~new_n92_ & ~new_n95_;
  assign new_n97_ = v7 & ~v10;
  assign new_n98_ = v6 & ~v11;
  assign new_n99_ = ~new_n97_ & ~new_n98_;
  assign new_n100_ = v8 & ~new_n93_;
  assign new_n101_ = ~v4 & new_n100_;
  assign new_n102_ = ~new_n99_ & ~new_n101_;
  assign new_n103_ = ~new_n89_ & ~new_n90_;
  assign new_n104_ = ~v8 & ~new_n103_;
  assign new_n105_ = ~new_n102_ & ~new_n104_;
  assign new_n106_ = v1 & ~new_n105_;
  assign new_n107_ = ~new_n96_ & ~new_n106_;
  assign new_n108_ = v5 & ~new_n107_;
  assign new_n109_ = v1 & ~v11;
  assign new_n110_ = ~v7 & ~new_n109_;
  assign new_n111_ = v3 & v10;
  assign new_n112_ = v2 & ~v10;
  assign new_n113_ = ~new_n111_ & ~new_n112_;
  assign new_n114_ = ~new_n110_ & ~new_n113_;
  assign new_n115_ = ~v7 & v11;
  assign new_n116_ = ~v4 & v8;
  assign new_n117_ = ~new_n115_ & ~new_n116_;
  assign new_n118_ = ~v9 & new_n117_;
  assign new_n119_ = v1 & new_n118_;
  assign new_n120_ = ~new_n114_ & ~new_n119_;
  assign new_n121_ = v6 & ~new_n120_;
  assign new_n122_ = ~v10 & new_n117_;
  assign new_n123_ = ~v9 & new_n122_;
  assign new_n124_ = v1 & new_n123_;
  assign new_n125_ = v3 & v11;
  assign new_n126_ = v2 & ~v11;
  assign new_n127_ = ~new_n125_ & ~new_n126_;
  assign new_n128_ = v7 & ~new_n127_;
  assign new_n129_ = ~new_n124_ & ~new_n128_;
  assign new_n130_ = ~new_n121_ & new_n129_;
  assign new_n131_ = ~new_n108_ & new_n130_;
  assign \v15.1  = new_n88_ | ~new_n131_;
  assign new_n133_ = v9 & v10;
  assign new_n134_ = v8 & new_n133_;
  assign new_n135_ = ~v1 & ~new_n134_;
  assign new_n136_ = v0 & ~new_n135_;
  assign new_n137_ = v5 & v6;
  assign new_n138_ = v4 & new_n137_;
  assign new_n139_ = v1 & ~v8;
  assign new_n140_ = ~v9 & ~v10;
  assign new_n141_ = new_n139_ & new_n140_;
  assign new_n142_ = ~new_n138_ & ~new_n141_;
  assign new_n143_ = ~new_n136_ & new_n142_;
  assign new_n144_ = ~v13 & ~new_n143_;
  assign new_n145_ = ~v12 & ~new_n144_;
  assign new_n146_ = ~new_n127_ & ~new_n145_;
  assign new_n147_ = v10 & v11;
  assign new_n148_ = v9 & new_n147_;
  assign new_n149_ = v2 & ~new_n148_;
  assign new_n150_ = ~v0 & v8;
  assign new_n151_ = ~v1 & ~v8;
  assign new_n152_ = ~new_n150_ & ~new_n151_;
  assign new_n153_ = ~new_n149_ & ~new_n152_;
  assign new_n154_ = ~v13 & ~new_n150_;
  assign new_n155_ = ~v5 & ~new_n154_;
  assign new_n156_ = v9 & v13;
  assign new_n157_ = ~new_n155_ & ~new_n156_;
  assign new_n158_ = ~new_n24_ & ~new_n157_;
  assign new_n159_ = ~v0 & ~v6;
  assign new_n160_ = v8 & v9;
  assign new_n161_ = new_n159_ & new_n160_;
  assign new_n162_ = ~new_n158_ & ~new_n161_;
  assign new_n163_ = v11 & ~new_n162_;
  assign new_n164_ = ~new_n153_ & ~new_n163_;
  assign new_n165_ = ~v3 & ~new_n164_;
  assign new_n166_ = ~v13 & ~new_n151_;
  assign new_n167_ = ~new_n54_ & ~new_n166_;
  assign new_n168_ = ~new_n48_ & new_n167_;
  assign new_n169_ = new_n140_ & new_n150_;
  assign new_n170_ = ~new_n168_ & ~new_n169_;
  assign new_n171_ = ~v11 & ~new_n170_;
  assign new_n172_ = ~v2 & new_n171_;
  assign new_n173_ = ~new_n165_ & ~new_n172_;
  assign new_n174_ = ~v4 & ~new_n173_;
  assign new_n175_ = v2 & ~new_n147_;
  assign new_n176_ = ~v0 & v9;
  assign new_n177_ = ~v1 & ~v9;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign new_n179_ = ~new_n175_ & ~new_n178_;
  assign new_n180_ = v8 & v13;
  assign new_n181_ = ~new_n176_ & ~new_n180_;
  assign new_n182_ = ~v6 & ~new_n181_;
  assign new_n183_ = v10 & v13;
  assign new_n184_ = v8 & new_n183_;
  assign new_n185_ = ~new_n182_ & ~new_n184_;
  assign new_n186_ = v11 & ~new_n185_;
  assign new_n187_ = ~new_n179_ & ~new_n186_;
  assign new_n188_ = ~v5 & ~new_n187_;
  assign new_n189_ = v13 & ~new_n24_;
  assign new_n190_ = v9 & new_n189_;
  assign new_n191_ = v8 & new_n190_;
  assign new_n192_ = ~v0 & v10;
  assign new_n193_ = ~v1 & ~v10;
  assign new_n194_ = ~new_n192_ & ~new_n193_;
  assign new_n195_ = ~v6 & ~new_n194_;
  assign new_n196_ = ~new_n191_ & ~new_n195_;
  assign new_n197_ = v11 & ~new_n196_;
  assign new_n198_ = ~v2 & v13;
  assign new_n199_ = ~new_n197_ & ~new_n198_;
  assign new_n200_ = ~new_n188_ & new_n199_;
  assign new_n201_ = ~v3 & ~new_n200_;
  assign new_n202_ = ~v6 & v10;
  assign new_n203_ = v9 & ~v10;
  assign new_n204_ = ~v5 & new_n203_;
  assign new_n205_ = ~new_n202_ & ~new_n204_;
  assign new_n206_ = ~v0 & ~new_n205_;
  assign new_n207_ = ~v8 & v13;
  assign new_n208_ = ~new_n177_ & ~new_n207_;
  assign new_n209_ = ~v5 & ~new_n208_;
  assign new_n210_ = ~v9 & v13;
  assign new_n211_ = ~v8 & new_n210_;
  assign new_n212_ = ~new_n209_ & ~new_n211_;
  assign new_n213_ = ~new_n48_ & ~new_n212_;
  assign new_n214_ = ~v1 & new_n65_;
  assign new_n215_ = ~new_n213_ & ~new_n214_;
  assign new_n216_ = ~new_n206_ & new_n215_;
  assign new_n217_ = ~v11 & ~new_n216_;
  assign new_n218_ = ~v2 & new_n217_;
  assign new_n219_ = ~new_n201_ & ~new_n218_;
  assign new_n220_ = ~new_n174_ & new_n219_;
  assign new_n221_ = ~v12 & ~new_n220_;
  assign new_n222_ = v8 & v11;
  assign new_n223_ = ~v2 & ~new_n222_;
  assign new_n224_ = ~v1 & ~new_n133_;
  assign new_n225_ = v0 & ~new_n224_;
  assign new_n226_ = v1 & new_n140_;
  assign new_n227_ = ~new_n225_ & ~new_n226_;
  assign new_n228_ = ~new_n223_ & ~new_n227_;
  assign new_n229_ = v6 & v9;
  assign new_n230_ = v5 & v10;
  assign new_n231_ = ~new_n229_ & ~new_n230_;
  assign new_n232_ = ~new_n207_ & ~new_n231_;
  assign new_n233_ = v10 & ~v13;
  assign new_n234_ = v9 & new_n233_;
  assign new_n235_ = ~new_n232_ & ~new_n234_;
  assign new_n236_ = v0 & ~new_n235_;
  assign new_n237_ = v6 & v8;
  assign new_n238_ = v5 & new_n237_;
  assign new_n239_ = ~new_n236_ & ~new_n238_;
  assign new_n240_ = v11 & ~new_n239_;
  assign new_n241_ = ~new_n228_ & ~new_n240_;
  assign new_n242_ = v3 & ~new_n241_;
  assign new_n243_ = v1 & ~v10;
  assign new_n244_ = ~v6 & ~new_n243_;
  assign new_n245_ = v5 & ~new_n244_;
  assign new_n246_ = ~v9 & ~new_n202_;
  assign new_n247_ = v1 & new_n246_;
  assign new_n248_ = ~new_n245_ & ~new_n247_;
  assign new_n249_ = ~new_n225_ & new_n248_;
  assign new_n250_ = ~v8 & ~new_n249_;
  assign new_n251_ = v5 & ~v10;
  assign new_n252_ = ~new_n246_ & ~new_n251_;
  assign new_n253_ = ~v13 & ~new_n252_;
  assign new_n254_ = v1 & new_n253_;
  assign new_n255_ = ~new_n250_ & ~new_n254_;
  assign new_n256_ = ~v11 & ~new_n255_;
  assign new_n257_ = v2 & new_n256_;
  assign new_n258_ = ~new_n242_ & ~new_n257_;
  assign new_n259_ = v4 & ~new_n258_;
  assign new_n260_ = v9 & v11;
  assign new_n261_ = ~v2 & ~new_n260_;
  assign new_n262_ = v0 & v10;
  assign new_n263_ = ~new_n243_ & ~new_n262_;
  assign new_n264_ = ~new_n261_ & ~new_n263_;
  assign new_n265_ = ~v13 & ~new_n65_;
  assign new_n266_ = v8 & new_n265_;
  assign new_n267_ = v0 & new_n266_;
  assign new_n268_ = ~new_n229_ & ~new_n267_;
  assign new_n269_ = v11 & ~new_n268_;
  assign new_n270_ = ~new_n264_ & ~new_n269_;
  assign new_n271_ = v3 & ~new_n270_;
  assign new_n272_ = ~v8 & ~v13;
  assign new_n273_ = v1 & new_n272_;
  assign new_n274_ = v9 & ~new_n273_;
  assign new_n275_ = v6 & ~new_n274_;
  assign new_n276_ = v9 & ~new_n272_;
  assign new_n277_ = ~v10 & ~new_n276_;
  assign new_n278_ = v1 & new_n277_;
  assign new_n279_ = v0 & new_n61_;
  assign new_n280_ = ~new_n278_ & ~new_n279_;
  assign new_n281_ = ~new_n275_ & new_n280_;
  assign new_n282_ = ~v11 & ~new_n281_;
  assign new_n283_ = v2 & new_n282_;
  assign new_n284_ = ~new_n271_ & ~new_n283_;
  assign new_n285_ = v5 & ~new_n284_;
  assign new_n286_ = v0 & v8;
  assign new_n287_ = v9 & ~v13;
  assign new_n288_ = new_n286_ & new_n287_;
  assign new_n289_ = ~v10 & ~new_n288_;
  assign new_n290_ = v11 & ~new_n289_;
  assign new_n291_ = ~v2 & ~new_n290_;
  assign new_n292_ = v3 & ~new_n291_;
  assign new_n293_ = ~v9 & ~v13;
  assign new_n294_ = new_n139_ & new_n293_;
  assign new_n295_ = v10 & ~new_n294_;
  assign new_n296_ = ~v11 & ~new_n295_;
  assign new_n297_ = v2 & new_n296_;
  assign new_n298_ = ~new_n292_ & ~new_n297_;
  assign new_n299_ = v6 & ~new_n298_;
  assign new_n300_ = ~new_n285_ & ~new_n299_;
  assign new_n301_ = ~new_n259_ & new_n300_;
  assign new_n302_ = ~new_n221_ & new_n301_;
  assign new_n303_ = ~new_n146_ & new_n302_;
  assign new_n304_ = v7 & ~new_n303_;
  assign new_n305_ = ~v0 & v11;
  assign new_n306_ = ~v1 & ~v11;
  assign new_n307_ = ~new_n305_ & ~new_n306_;
  assign new_n308_ = v4 & v5;
  assign new_n309_ = v6 & ~v13;
  assign new_n310_ = new_n308_ & new_n309_;
  assign new_n311_ = ~v12 & ~new_n310_;
  assign new_n312_ = ~new_n307_ & ~new_n311_;
  assign new_n313_ = ~v2 & ~v10;
  assign new_n314_ = v6 & ~new_n313_;
  assign new_n315_ = v9 & ~new_n67_;
  assign new_n316_ = ~v1 & ~new_n315_;
  assign new_n317_ = ~v4 & v13;
  assign new_n318_ = ~new_n316_ & ~new_n317_;
  assign new_n319_ = ~new_n314_ & ~new_n318_;
  assign new_n320_ = v13 & ~new_n48_;
  assign new_n321_ = ~v8 & new_n320_;
  assign new_n322_ = ~v2 & new_n321_;
  assign new_n323_ = ~new_n319_ & ~new_n322_;
  assign new_n324_ = ~v5 & ~new_n323_;
  assign new_n325_ = ~v4 & ~new_n166_;
  assign new_n326_ = ~new_n207_ & ~new_n325_;
  assign new_n327_ = ~new_n48_ & ~new_n326_;
  assign new_n328_ = ~v9 & new_n327_;
  assign new_n329_ = ~v2 & new_n328_;
  assign new_n330_ = ~new_n214_ & ~new_n329_;
  assign new_n331_ = ~new_n324_ & new_n330_;
  assign new_n332_ = ~v12 & ~new_n331_;
  assign new_n333_ = v0 & new_n332_;
  assign new_n334_ = v4 & ~v8;
  assign new_n335_ = v9 & ~new_n334_;
  assign new_n336_ = ~new_n244_ & ~new_n335_;
  assign new_n337_ = v5 & new_n336_;
  assign new_n338_ = ~v8 & new_n246_;
  assign new_n339_ = v4 & new_n338_;
  assign new_n340_ = v1 & new_n339_;
  assign new_n341_ = ~new_n24_ & ~new_n340_;
  assign new_n342_ = ~new_n337_ & new_n341_;
  assign new_n343_ = v2 & ~new_n342_;
  assign new_n344_ = ~v5 & v9;
  assign new_n345_ = ~v8 & ~new_n344_;
  assign new_n346_ = v4 & ~v9;
  assign new_n347_ = ~new_n345_ & ~new_n346_;
  assign new_n348_ = ~new_n202_ & ~new_n347_;
  assign new_n349_ = v4 & new_n251_;
  assign new_n350_ = ~new_n348_ & ~new_n349_;
  assign new_n351_ = ~v13 & ~new_n350_;
  assign new_n352_ = v1 & new_n351_;
  assign new_n353_ = ~new_n343_ & ~new_n352_;
  assign new_n354_ = ~v0 & ~new_n353_;
  assign new_n355_ = ~new_n333_ & ~new_n354_;
  assign new_n356_ = v11 & ~new_n355_;
  assign new_n357_ = ~v3 & v10;
  assign new_n358_ = v6 & ~new_n357_;
  assign new_n359_ = ~v9 & ~new_n116_;
  assign new_n360_ = ~v0 & ~new_n359_;
  assign new_n361_ = ~new_n317_ & ~new_n360_;
  assign new_n362_ = ~new_n358_ & ~new_n361_;
  assign new_n363_ = v8 & new_n189_;
  assign new_n364_ = ~v3 & new_n363_;
  assign new_n365_ = ~new_n362_ & ~new_n364_;
  assign new_n366_ = ~v5 & ~new_n365_;
  assign new_n367_ = ~v4 & ~new_n154_;
  assign new_n368_ = ~new_n180_ & ~new_n367_;
  assign new_n369_ = ~new_n24_ & ~new_n368_;
  assign new_n370_ = v9 & new_n369_;
  assign new_n371_ = ~v3 & new_n370_;
  assign new_n372_ = ~v0 & new_n202_;
  assign new_n373_ = ~new_n371_ & ~new_n372_;
  assign new_n374_ = ~new_n366_ & new_n373_;
  assign new_n375_ = ~v12 & ~new_n374_;
  assign new_n376_ = v1 & new_n375_;
  assign new_n377_ = v4 & v8;
  assign new_n378_ = ~v9 & ~new_n377_;
  assign new_n379_ = ~v6 & ~new_n262_;
  assign new_n380_ = ~new_n378_ & ~new_n379_;
  assign new_n381_ = v5 & new_n380_;
  assign new_n382_ = v9 & ~new_n65_;
  assign new_n383_ = v8 & new_n382_;
  assign new_n384_ = v4 & new_n383_;
  assign new_n385_ = v0 & new_n384_;
  assign new_n386_ = ~new_n48_ & ~new_n385_;
  assign new_n387_ = ~new_n381_ & new_n386_;
  assign new_n388_ = v3 & ~new_n387_;
  assign new_n389_ = v4 & new_n230_;
  assign new_n390_ = ~new_n79_ & ~new_n389_;
  assign new_n391_ = ~v13 & ~new_n390_;
  assign new_n392_ = v0 & new_n391_;
  assign new_n393_ = ~new_n388_ & ~new_n392_;
  assign new_n394_ = ~v1 & ~new_n393_;
  assign new_n395_ = ~new_n376_ & ~new_n394_;
  assign new_n396_ = ~v11 & ~new_n395_;
  assign new_n397_ = ~new_n356_ & ~new_n396_;
  assign new_n398_ = ~new_n312_ & new_n397_;
  assign new_n399_ = ~v7 & ~new_n398_;
  assign new_n400_ = v8 & ~v9;
  assign new_n401_ = v4 & new_n400_;
  assign new_n402_ = ~new_n54_ & ~new_n401_;
  assign new_n403_ = ~v10 & ~new_n402_;
  assign new_n404_ = v1 & new_n403_;
  assign new_n405_ = v5 & ~new_n378_;
  assign new_n406_ = ~v10 & ~new_n405_;
  assign new_n407_ = v6 & ~new_n406_;
  assign new_n408_ = ~new_n404_ & ~new_n407_;
  assign new_n409_ = v3 & ~new_n408_;
  assign new_n410_ = ~v0 & new_n409_;
  assign new_n411_ = ~v1 & new_n67_;
  assign new_n412_ = ~v13 & ~new_n411_;
  assign new_n413_ = ~v2 & ~new_n412_;
  assign new_n414_ = ~v8 & v9;
  assign new_n415_ = ~v4 & new_n414_;
  assign new_n416_ = ~new_n66_ & ~new_n415_;
  assign new_n417_ = ~v1 & ~new_n416_;
  assign new_n418_ = ~new_n25_ & ~new_n334_;
  assign new_n419_ = v13 & new_n418_;
  assign new_n420_ = ~new_n417_ & ~new_n419_;
  assign new_n421_ = v10 & ~new_n420_;
  assign new_n422_ = v13 & ~new_n28_;
  assign new_n423_ = ~v6 & new_n422_;
  assign new_n424_ = ~new_n421_ & ~new_n423_;
  assign new_n425_ = ~new_n413_ & new_n424_;
  assign new_n426_ = ~v12 & ~new_n425_;
  assign new_n427_ = ~v3 & new_n426_;
  assign new_n428_ = v0 & new_n427_;
  assign new_n429_ = ~new_n410_ & ~new_n428_;
  assign new_n430_ = v11 & ~new_n429_;
  assign new_n431_ = v4 & new_n414_;
  assign new_n432_ = ~new_n25_ & ~new_n431_;
  assign new_n433_ = v10 & ~new_n432_;
  assign new_n434_ = v0 & new_n433_;
  assign new_n435_ = v5 & ~new_n335_;
  assign new_n436_ = v10 & ~new_n435_;
  assign new_n437_ = v6 & ~new_n436_;
  assign new_n438_ = ~new_n434_ & ~new_n437_;
  assign new_n439_ = v2 & ~new_n438_;
  assign new_n440_ = ~v1 & new_n439_;
  assign new_n441_ = ~v0 & new_n116_;
  assign new_n442_ = ~v13 & ~new_n441_;
  assign new_n443_ = ~v3 & ~new_n442_;
  assign new_n444_ = ~v4 & new_n400_;
  assign new_n445_ = ~new_n344_ & ~new_n444_;
  assign new_n446_ = ~v0 & ~new_n445_;
  assign new_n447_ = ~new_n54_ & ~new_n377_;
  assign new_n448_ = v13 & new_n447_;
  assign new_n449_ = ~new_n446_ & ~new_n448_;
  assign new_n450_ = ~v10 & ~new_n449_;
  assign new_n451_ = ~v8 & ~new_n54_;
  assign new_n452_ = ~v4 & ~v9;
  assign new_n453_ = ~new_n451_ & ~new_n452_;
  assign new_n454_ = v13 & ~new_n453_;
  assign new_n455_ = ~v6 & new_n454_;
  assign new_n456_ = ~new_n450_ & ~new_n455_;
  assign new_n457_ = ~new_n443_ & new_n456_;
  assign new_n458_ = ~v12 & ~new_n457_;
  assign new_n459_ = ~v2 & new_n458_;
  assign new_n460_ = v1 & new_n459_;
  assign new_n461_ = ~new_n440_ & ~new_n460_;
  assign new_n462_ = ~v11 & ~new_n461_;
  assign new_n463_ = ~new_n430_ & ~new_n462_;
  assign new_n464_ = ~new_n399_ & new_n463_;
  assign \v15.2  = new_n304_ | ~new_n464_;
  assign new_n466_ = ~v1 & ~new_n160_;
  assign new_n467_ = v0 & ~new_n466_;
  assign new_n468_ = ~v8 & ~v9;
  assign new_n469_ = v1 & new_n468_;
  assign new_n470_ = ~new_n308_ & ~new_n469_;
  assign new_n471_ = ~new_n467_ & new_n470_;
  assign new_n472_ = ~v13 & ~new_n471_;
  assign new_n473_ = ~v12 & ~new_n472_;
  assign new_n474_ = ~new_n113_ & ~new_n473_;
  assign new_n475_ = ~new_n25_ & ~new_n368_;
  assign new_n476_ = ~v0 & new_n344_;
  assign new_n477_ = ~new_n475_ & ~new_n476_;
  assign new_n478_ = ~new_n417_ & new_n477_;
  assign new_n479_ = ~v12 & ~new_n478_;
  assign new_n480_ = ~v3 & new_n479_;
  assign new_n481_ = v9 & ~new_n207_;
  assign new_n482_ = v4 & new_n481_;
  assign new_n483_ = v8 & ~v13;
  assign new_n484_ = v5 & new_n483_;
  assign new_n485_ = ~new_n482_ & ~new_n484_;
  assign new_n486_ = v0 & ~new_n485_;
  assign new_n487_ = v1 & ~v9;
  assign new_n488_ = ~v5 & ~new_n487_;
  assign new_n489_ = v8 & ~new_n488_;
  assign new_n490_ = v4 & new_n489_;
  assign new_n491_ = ~new_n54_ & ~new_n490_;
  assign new_n492_ = ~new_n486_ & new_n491_;
  assign new_n493_ = v3 & ~new_n492_;
  assign new_n494_ = ~new_n480_ & ~new_n493_;
  assign new_n495_ = v10 & ~new_n494_;
  assign new_n496_ = ~v8 & ~v10;
  assign new_n497_ = ~v3 & ~new_n496_;
  assign new_n498_ = v0 & v9;
  assign new_n499_ = ~new_n487_ & ~new_n498_;
  assign new_n500_ = ~new_n497_ & ~new_n499_;
  assign new_n501_ = v5 & ~v8;
  assign new_n502_ = v1 & new_n293_;
  assign new_n503_ = ~new_n501_ & ~new_n502_;
  assign new_n504_ = ~v10 & ~new_n503_;
  assign new_n505_ = ~new_n500_ & ~new_n504_;
  assign new_n506_ = v4 & ~new_n505_;
  assign new_n507_ = ~v10 & ~new_n274_;
  assign new_n508_ = ~v3 & ~new_n507_;
  assign new_n509_ = v5 & ~new_n508_;
  assign new_n510_ = ~new_n506_ & ~new_n509_;
  assign new_n511_ = v2 & ~new_n510_;
  assign new_n512_ = v3 & ~new_n140_;
  assign new_n513_ = ~new_n152_ & ~new_n512_;
  assign new_n514_ = ~v5 & ~new_n166_;
  assign new_n515_ = ~new_n210_ & ~new_n514_;
  assign new_n516_ = ~v10 & ~new_n515_;
  assign new_n517_ = ~new_n513_ & ~new_n516_;
  assign new_n518_ = ~v4 & ~new_n517_;
  assign new_n519_ = v13 & ~new_n54_;
  assign new_n520_ = ~v8 & new_n519_;
  assign new_n521_ = ~v5 & ~new_n178_;
  assign new_n522_ = ~new_n520_ & ~new_n521_;
  assign new_n523_ = ~v10 & ~new_n522_;
  assign new_n524_ = ~v3 & v13;
  assign new_n525_ = ~new_n523_ & ~new_n524_;
  assign new_n526_ = ~new_n518_ & new_n525_;
  assign new_n527_ = ~v12 & ~new_n526_;
  assign new_n528_ = ~v2 & new_n527_;
  assign new_n529_ = ~new_n511_ & ~new_n528_;
  assign new_n530_ = ~new_n495_ & new_n529_;
  assign new_n531_ = ~new_n474_ & new_n530_;
  assign new_n532_ = v6 & ~new_n531_;
  assign new_n533_ = v5 & ~v13;
  assign new_n534_ = v4 & new_n533_;
  assign new_n535_ = ~v12 & ~new_n534_;
  assign new_n536_ = ~new_n194_ & ~new_n535_;
  assign new_n537_ = ~v2 & ~v9;
  assign new_n538_ = v5 & ~new_n537_;
  assign new_n539_ = ~new_n166_ & ~new_n538_;
  assign new_n540_ = ~v4 & new_n539_;
  assign new_n541_ = ~v2 & new_n520_;
  assign new_n542_ = ~v1 & new_n66_;
  assign new_n543_ = ~new_n541_ & ~new_n542_;
  assign new_n544_ = ~new_n540_ & new_n543_;
  assign new_n545_ = ~v12 & ~new_n544_;
  assign new_n546_ = v0 & new_n545_;
  assign new_n547_ = v4 & ~new_n488_;
  assign new_n548_ = v2 & new_n547_;
  assign new_n549_ = ~v13 & ~new_n344_;
  assign new_n550_ = v1 & new_n549_;
  assign new_n551_ = ~new_n548_ & ~new_n550_;
  assign new_n552_ = ~v8 & ~new_n551_;
  assign new_n553_ = v2 & v5;
  assign new_n554_ = v4 & ~v13;
  assign new_n555_ = v1 & new_n554_;
  assign new_n556_ = ~new_n553_ & ~new_n555_;
  assign new_n557_ = ~v9 & ~new_n556_;
  assign new_n558_ = ~new_n552_ & ~new_n557_;
  assign new_n559_ = ~v0 & ~new_n558_;
  assign new_n560_ = ~new_n546_ & ~new_n559_;
  assign new_n561_ = v10 & ~new_n560_;
  assign new_n562_ = ~v3 & v9;
  assign new_n563_ = v5 & ~new_n562_;
  assign new_n564_ = ~new_n154_ & ~new_n563_;
  assign new_n565_ = ~v4 & new_n564_;
  assign new_n566_ = v13 & ~new_n25_;
  assign new_n567_ = v8 & new_n566_;
  assign new_n568_ = ~v3 & new_n567_;
  assign new_n569_ = ~new_n476_ & ~new_n568_;
  assign new_n570_ = ~new_n565_ & new_n569_;
  assign new_n571_ = ~v12 & ~new_n570_;
  assign new_n572_ = v1 & new_n571_;
  assign new_n573_ = ~v5 & ~new_n498_;
  assign new_n574_ = v4 & ~new_n573_;
  assign new_n575_ = v3 & new_n574_;
  assign new_n576_ = ~v13 & ~new_n66_;
  assign new_n577_ = v0 & new_n576_;
  assign new_n578_ = ~new_n575_ & ~new_n577_;
  assign new_n579_ = v8 & ~new_n578_;
  assign new_n580_ = v3 & v5;
  assign new_n581_ = v0 & new_n554_;
  assign new_n582_ = ~new_n580_ & ~new_n581_;
  assign new_n583_ = v9 & ~new_n582_;
  assign new_n584_ = ~new_n579_ & ~new_n583_;
  assign new_n585_ = ~v1 & ~new_n584_;
  assign new_n586_ = ~new_n572_ & ~new_n585_;
  assign new_n587_ = ~v10 & ~new_n586_;
  assign new_n588_ = ~new_n561_ & ~new_n587_;
  assign new_n589_ = ~new_n536_ & new_n588_;
  assign new_n590_ = ~v6 & ~new_n589_;
  assign new_n591_ = v0 & ~v3;
  assign new_n592_ = new_n133_ & new_n591_;
  assign new_n593_ = v1 & ~v2;
  assign new_n594_ = new_n140_ & new_n593_;
  assign new_n595_ = ~new_n592_ & ~new_n594_;
  assign new_n596_ = ~v4 & ~new_n595_;
  assign new_n597_ = v8 & v10;
  assign new_n598_ = new_n591_ & new_n597_;
  assign new_n599_ = new_n496_ & new_n593_;
  assign new_n600_ = ~new_n598_ & ~new_n599_;
  assign new_n601_ = ~v5 & ~new_n600_;
  assign new_n602_ = v2 & ~new_n160_;
  assign new_n603_ = v10 & ~new_n602_;
  assign new_n604_ = v0 & new_n603_;
  assign new_n605_ = v1 & new_n313_;
  assign new_n606_ = ~new_n604_ & ~new_n605_;
  assign new_n607_ = ~v3 & ~new_n606_;
  assign new_n608_ = ~v8 & new_n140_;
  assign new_n609_ = new_n593_ & new_n608_;
  assign new_n610_ = ~new_n607_ & ~new_n609_;
  assign new_n611_ = ~new_n601_ & new_n610_;
  assign new_n612_ = ~new_n596_ & new_n611_;
  assign new_n613_ = v13 & ~new_n612_;
  assign new_n614_ = ~v1 & ~v3;
  assign new_n615_ = v0 & new_n614_;
  assign new_n616_ = ~v8 & new_n133_;
  assign new_n617_ = new_n615_ & new_n616_;
  assign new_n618_ = ~v0 & new_n593_;
  assign new_n619_ = v8 & new_n140_;
  assign new_n620_ = new_n618_ & new_n619_;
  assign new_n621_ = ~new_n617_ & ~new_n620_;
  assign new_n622_ = ~v4 & ~new_n621_;
  assign new_n623_ = ~new_n613_ & ~new_n622_;
  assign new_n624_ = ~v12 & ~new_n623_;
  assign new_n625_ = v10 & ~new_n488_;
  assign new_n626_ = v8 & new_n625_;
  assign new_n627_ = v3 & new_n626_;
  assign new_n628_ = ~v0 & new_n627_;
  assign new_n629_ = ~v10 & ~new_n573_;
  assign new_n630_ = ~v8 & new_n629_;
  assign new_n631_ = v2 & new_n630_;
  assign new_n632_ = ~v1 & new_n631_;
  assign new_n633_ = ~new_n628_ & ~new_n632_;
  assign new_n634_ = v4 & ~new_n633_;
  assign new_n635_ = ~v0 & v3;
  assign new_n636_ = new_n133_ & new_n635_;
  assign new_n637_ = ~v1 & v2;
  assign new_n638_ = new_n140_ & new_n637_;
  assign new_n639_ = ~new_n636_ & ~new_n638_;
  assign new_n640_ = v5 & ~new_n639_;
  assign new_n641_ = ~new_n634_ & ~new_n640_;
  assign new_n642_ = ~new_n624_ & new_n641_;
  assign new_n643_ = ~new_n590_ & new_n642_;
  assign \v15.3  = new_n532_ | ~new_n643_;
  assign new_n645_ = ~new_n139_ & ~new_n286_;
  assign new_n646_ = ~v4 & new_n645_;
  assign new_n647_ = ~v13 & ~new_n646_;
  assign new_n648_ = ~v12 & ~new_n647_;
  assign new_n649_ = ~new_n94_ & ~new_n648_;
  assign new_n650_ = ~new_n537_ & ~new_n562_;
  assign new_n651_ = ~new_n150_ & new_n166_;
  assign new_n652_ = ~new_n650_ & ~new_n651_;
  assign new_n653_ = ~v4 & new_n652_;
  assign new_n654_ = v3 & ~new_n468_;
  assign new_n655_ = ~v2 & ~new_n654_;
  assign new_n656_ = ~v3 & new_n160_;
  assign new_n657_ = ~new_n655_ & ~new_n656_;
  assign new_n658_ = v13 & ~new_n657_;
  assign new_n659_ = ~new_n653_ & ~new_n658_;
  assign new_n660_ = ~v12 & ~new_n659_;
  assign new_n661_ = ~v3 & ~new_n468_;
  assign new_n662_ = v2 & ~new_n661_;
  assign new_n663_ = v3 & new_n160_;
  assign new_n664_ = ~new_n662_ & ~new_n663_;
  assign new_n665_ = v4 & ~new_n664_;
  assign new_n666_ = ~new_n660_ & ~new_n665_;
  assign new_n667_ = ~new_n649_ & new_n666_;
  assign new_n668_ = v5 & ~new_n667_;
  assign new_n669_ = ~new_n177_ & ~new_n476_;
  assign new_n670_ = ~v8 & ~new_n669_;
  assign new_n671_ = v2 & new_n670_;
  assign new_n672_ = ~v5 & ~v13;
  assign new_n673_ = v3 & v8;
  assign new_n674_ = ~new_n672_ & ~new_n673_;
  assign new_n675_ = v9 & ~new_n674_;
  assign new_n676_ = ~v0 & new_n675_;
  assign new_n677_ = v13 & ~new_n673_;
  assign new_n678_ = ~v9 & ~new_n677_;
  assign new_n679_ = ~v5 & new_n678_;
  assign new_n680_ = ~v1 & new_n679_;
  assign new_n681_ = ~new_n676_ & ~new_n680_;
  assign new_n682_ = ~new_n671_ & new_n681_;
  assign new_n683_ = v4 & ~new_n682_;
  assign new_n684_ = v0 & new_n344_;
  assign new_n685_ = ~new_n487_ & ~new_n684_;
  assign new_n686_ = ~v8 & ~new_n685_;
  assign new_n687_ = ~v2 & new_n686_;
  assign new_n688_ = ~v3 & v8;
  assign new_n689_ = ~new_n34_ & ~new_n688_;
  assign new_n690_ = v9 & ~new_n689_;
  assign new_n691_ = v0 & new_n690_;
  assign new_n692_ = v4 & ~new_n688_;
  assign new_n693_ = ~v9 & ~new_n692_;
  assign new_n694_ = ~v5 & new_n693_;
  assign new_n695_ = v1 & new_n694_;
  assign new_n696_ = ~new_n691_ & ~new_n695_;
  assign new_n697_ = ~new_n687_ & new_n696_;
  assign new_n698_ = v13 & ~new_n697_;
  assign new_n699_ = v0 & ~v1;
  assign new_n700_ = new_n414_ & new_n699_;
  assign new_n701_ = ~v0 & v1;
  assign new_n702_ = new_n400_ & new_n701_;
  assign new_n703_ = ~new_n700_ & ~new_n702_;
  assign new_n704_ = ~v5 & ~new_n703_;
  assign new_n705_ = ~v4 & new_n704_;
  assign new_n706_ = ~new_n698_ & ~new_n705_;
  assign new_n707_ = ~v12 & ~new_n706_;
  assign new_n708_ = ~v12 & ~new_n273_;
  assign new_n709_ = v9 & ~new_n708_;
  assign new_n710_ = ~v0 & new_n709_;
  assign new_n711_ = v0 & new_n483_;
  assign new_n712_ = ~v12 & ~new_n711_;
  assign new_n713_ = ~v9 & ~new_n712_;
  assign new_n714_ = ~v1 & new_n713_;
  assign new_n715_ = ~new_n710_ & ~new_n714_;
  assign new_n716_ = ~v5 & ~new_n715_;
  assign new_n717_ = ~new_n707_ & ~new_n716_;
  assign new_n718_ = ~new_n683_ & new_n717_;
  assign \v15.4  = new_n668_ | ~new_n718_;
  assign new_n720_ = ~v12 & v13;
  assign new_n721_ = v2 & ~v8;
  assign new_n722_ = ~new_n673_ & ~new_n721_;
  assign new_n723_ = v4 & ~new_n722_;
  assign new_n724_ = ~v4 & ~new_n152_;
  assign new_n725_ = ~new_n723_ & ~new_n724_;
  assign new_n726_ = ~new_n720_ & ~new_n725_;
  assign new_n727_ = ~v2 & ~v8;
  assign new_n728_ = ~new_n688_ & ~new_n727_;
  assign new_n729_ = v4 & ~new_n728_;
  assign new_n730_ = ~v4 & ~new_n645_;
  assign new_n731_ = ~new_n729_ & ~new_n730_;
  assign new_n732_ = v13 & ~new_n731_;
  assign new_n733_ = ~v12 & new_n732_;
  assign \v15.5  = new_n726_ | new_n733_;
  assign new_n735_ = ~new_n23_ & ~new_n115_;
  assign new_n736_ = v4 & ~v5;
  assign new_n737_ = new_n414_ & new_n736_;
  assign new_n738_ = ~v4 & v5;
  assign new_n739_ = new_n400_ & new_n738_;
  assign new_n740_ = ~new_n737_ & ~new_n739_;
  assign new_n741_ = ~v12 & new_n320_;
  assign new_n742_ = ~v2 & new_n741_;
  assign new_n743_ = v0 & new_n742_;
  assign new_n744_ = v2 & v12;
  assign new_n745_ = ~v0 & new_n744_;
  assign new_n746_ = ~new_n743_ & ~new_n745_;
  assign new_n747_ = ~new_n740_ & ~new_n746_;
  assign new_n748_ = ~v1 & new_n272_;
  assign new_n749_ = ~new_n180_ & ~new_n748_;
  assign new_n750_ = ~v12 & ~new_n749_;
  assign new_n751_ = ~v4 & new_n750_;
  assign new_n752_ = ~v2 & new_n751_;
  assign new_n753_ = v0 & new_n752_;
  assign new_n754_ = v2 & v4;
  assign new_n755_ = ~v0 & new_n754_;
  assign new_n756_ = v6 & new_n272_;
  assign new_n757_ = new_n755_ & new_n756_;
  assign new_n758_ = ~new_n753_ & ~new_n757_;
  assign new_n759_ = ~v10 & ~new_n758_;
  assign new_n760_ = v9 & new_n759_;
  assign new_n761_ = ~v5 & new_n760_;
  assign new_n762_ = ~new_n747_ & ~new_n761_;
  assign new_n763_ = ~new_n735_ & ~new_n762_;
  assign new_n764_ = ~v7 & ~v11;
  assign new_n765_ = ~new_n43_ & ~new_n764_;
  assign new_n766_ = new_n414_ & new_n738_;
  assign new_n767_ = new_n400_ & new_n736_;
  assign new_n768_ = ~new_n766_ & ~new_n767_;
  assign new_n769_ = ~v12 & new_n189_;
  assign new_n770_ = ~v3 & new_n769_;
  assign new_n771_ = v1 & new_n770_;
  assign new_n772_ = v3 & v12;
  assign new_n773_ = ~v1 & new_n772_;
  assign new_n774_ = ~new_n771_ & ~new_n773_;
  assign new_n775_ = ~new_n768_ & ~new_n774_;
  assign new_n776_ = ~v0 & new_n483_;
  assign new_n777_ = ~new_n207_ & ~new_n776_;
  assign new_n778_ = ~v12 & ~new_n777_;
  assign new_n779_ = ~v4 & new_n778_;
  assign new_n780_ = ~v3 & new_n779_;
  assign new_n781_ = v1 & new_n780_;
  assign new_n782_ = v3 & v4;
  assign new_n783_ = ~v1 & new_n782_;
  assign new_n784_ = v6 & new_n483_;
  assign new_n785_ = new_n783_ & new_n784_;
  assign new_n786_ = ~new_n781_ & ~new_n785_;
  assign new_n787_ = v10 & ~new_n786_;
  assign new_n788_ = ~v9 & new_n787_;
  assign new_n789_ = ~v5 & new_n788_;
  assign new_n790_ = ~new_n775_ & ~new_n789_;
  assign new_n791_ = ~new_n765_ & ~new_n790_;
  assign new_n792_ = v2 & v3;
  assign new_n793_ = ~new_n147_ & ~new_n792_;
  assign new_n794_ = v6 & ~new_n793_;
  assign new_n795_ = ~v6 & ~v11;
  assign new_n796_ = ~v2 & new_n795_;
  assign new_n797_ = ~new_n794_ & ~new_n796_;
  assign new_n798_ = v7 & ~new_n797_;
  assign new_n799_ = ~v6 & new_n115_;
  assign new_n800_ = ~new_n798_ & ~new_n799_;
  assign new_n801_ = ~new_n749_ & ~new_n800_;
  assign new_n802_ = v3 & new_n180_;
  assign new_n803_ = ~v10 & ~v13;
  assign new_n804_ = ~v8 & new_n803_;
  assign new_n805_ = ~new_n802_ & ~new_n804_;
  assign new_n806_ = v2 & ~new_n805_;
  assign new_n807_ = ~new_n180_ & ~new_n272_;
  assign new_n808_ = v10 & ~new_n807_;
  assign new_n809_ = ~v7 & new_n808_;
  assign new_n810_ = v3 & new_n809_;
  assign new_n811_ = v7 & ~v8;
  assign new_n812_ = new_n803_ & new_n811_;
  assign new_n813_ = ~new_n810_ & ~new_n812_;
  assign new_n814_ = ~new_n806_ & new_n813_;
  assign new_n815_ = ~v11 & ~new_n814_;
  assign new_n816_ = ~v1 & new_n815_;
  assign new_n817_ = v1 & v7;
  assign new_n818_ = v11 & v13;
  assign new_n819_ = v10 & new_n818_;
  assign new_n820_ = new_n817_ & new_n819_;
  assign new_n821_ = ~new_n816_ & ~new_n820_;
  assign new_n822_ = v6 & ~new_n821_;
  assign new_n823_ = ~new_n801_ & ~new_n822_;
  assign new_n824_ = v9 & ~new_n823_;
  assign new_n825_ = ~v3 & ~v7;
  assign new_n826_ = new_n89_ & new_n222_;
  assign new_n827_ = ~new_n825_ & ~new_n826_;
  assign new_n828_ = v10 & ~new_n827_;
  assign new_n829_ = ~v7 & ~new_n314_;
  assign new_n830_ = ~v11 & ~new_n160_;
  assign new_n831_ = ~v10 & new_n830_;
  assign new_n832_ = ~new_n792_ & ~new_n831_;
  assign new_n833_ = v7 & ~new_n832_;
  assign new_n834_ = v6 & new_n833_;
  assign new_n835_ = ~new_n829_ & ~new_n834_;
  assign new_n836_ = ~new_n828_ & new_n835_;
  assign new_n837_ = v13 & ~new_n836_;
  assign new_n838_ = v1 & new_n837_;
  assign new_n839_ = ~new_n824_ & ~new_n838_;
  assign new_n840_ = v0 & ~new_n839_;
  assign new_n841_ = ~new_n90_ & ~new_n792_;
  assign new_n842_ = v6 & ~new_n841_;
  assign new_n843_ = ~v3 & new_n35_;
  assign new_n844_ = ~new_n842_ & ~new_n843_;
  assign new_n845_ = v7 & ~new_n844_;
  assign new_n846_ = ~v6 & new_n764_;
  assign new_n847_ = ~new_n845_ & ~new_n846_;
  assign new_n848_ = ~new_n777_ & ~new_n847_;
  assign new_n849_ = v2 & new_n207_;
  assign new_n850_ = v8 & new_n233_;
  assign new_n851_ = ~new_n849_ & ~new_n850_;
  assign new_n852_ = v3 & ~new_n851_;
  assign new_n853_ = ~new_n207_ & ~new_n483_;
  assign new_n854_ = ~v10 & ~new_n853_;
  assign new_n855_ = ~v7 & new_n854_;
  assign new_n856_ = v2 & new_n855_;
  assign new_n857_ = v7 & v8;
  assign new_n858_ = new_n233_ & new_n857_;
  assign new_n859_ = ~new_n856_ & ~new_n858_;
  assign new_n860_ = ~new_n852_ & new_n859_;
  assign new_n861_ = v11 & ~new_n860_;
  assign new_n862_ = v6 & new_n861_;
  assign new_n863_ = ~v0 & new_n862_;
  assign new_n864_ = ~new_n848_ & ~new_n863_;
  assign new_n865_ = ~v9 & ~new_n864_;
  assign new_n866_ = v1 & new_n865_;
  assign new_n867_ = ~new_n840_ & ~new_n866_;
  assign new_n868_ = ~v12 & ~new_n867_;
  assign new_n869_ = v7 & new_n160_;
  assign new_n870_ = ~new_n177_ & ~new_n869_;
  assign new_n871_ = ~v11 & ~new_n870_;
  assign new_n872_ = v2 & new_n871_;
  assign new_n873_ = v3 & new_n260_;
  assign new_n874_ = v7 & ~new_n873_;
  assign new_n875_ = ~v1 & ~new_n874_;
  assign new_n876_ = ~v7 & v8;
  assign new_n877_ = new_n260_ & new_n876_;
  assign new_n878_ = ~new_n875_ & ~new_n877_;
  assign new_n879_ = ~new_n872_ & new_n878_;
  assign new_n880_ = ~v0 & ~new_n879_;
  assign new_n881_ = v3 & new_n43_;
  assign new_n882_ = ~new_n764_ & ~new_n881_;
  assign new_n883_ = ~v9 & ~new_n882_;
  assign new_n884_ = ~v8 & new_n883_;
  assign new_n885_ = ~v1 & new_n884_;
  assign new_n886_ = ~new_n880_ & ~new_n885_;
  assign new_n887_ = v12 & ~new_n886_;
  assign new_n888_ = ~new_n868_ & ~new_n887_;
  assign new_n889_ = ~v5 & ~new_n888_;
  assign new_n890_ = ~v9 & v12;
  assign new_n891_ = ~v3 & new_n137_;
  assign new_n892_ = ~v12 & ~v13;
  assign new_n893_ = new_n203_ & new_n892_;
  assign new_n894_ = new_n891_ & new_n893_;
  assign new_n895_ = ~new_n890_ & ~new_n894_;
  assign new_n896_ = v2 & ~new_n895_;
  assign new_n897_ = v9 & v12;
  assign new_n898_ = ~v2 & new_n137_;
  assign new_n899_ = new_n61_ & new_n892_;
  assign new_n900_ = new_n898_ & new_n899_;
  assign new_n901_ = ~new_n897_ & ~new_n900_;
  assign new_n902_ = v3 & ~new_n901_;
  assign new_n903_ = ~new_n896_ & ~new_n902_;
  assign new_n904_ = ~v1 & ~new_n903_;
  assign new_n905_ = v1 & new_n207_;
  assign new_n906_ = ~new_n483_ & ~new_n905_;
  assign new_n907_ = v11 & ~new_n906_;
  assign new_n908_ = ~v10 & new_n907_;
  assign new_n909_ = v6 & new_n908_;
  assign new_n910_ = v2 & new_n909_;
  assign new_n911_ = ~v13 & ~new_n24_;
  assign new_n912_ = ~v11 & new_n911_;
  assign new_n913_ = v8 & new_n912_;
  assign new_n914_ = v1 & new_n913_;
  assign new_n915_ = ~new_n910_ & ~new_n914_;
  assign new_n916_ = ~v12 & ~new_n915_;
  assign new_n917_ = v9 & new_n916_;
  assign new_n918_ = v5 & new_n917_;
  assign new_n919_ = ~v3 & new_n918_;
  assign new_n920_ = ~new_n904_ & ~new_n919_;
  assign new_n921_ = ~v7 & ~new_n920_;
  assign new_n922_ = ~v2 & v3;
  assign new_n923_ = ~v9 & new_n147_;
  assign new_n924_ = new_n922_ & new_n923_;
  assign new_n925_ = ~v3 & v7;
  assign new_n926_ = v9 & new_n90_;
  assign new_n927_ = new_n925_ & new_n926_;
  assign new_n928_ = ~new_n924_ & ~new_n927_;
  assign new_n929_ = v6 & ~new_n928_;
  assign new_n930_ = ~v3 & new_n260_;
  assign new_n931_ = ~v9 & ~v11;
  assign new_n932_ = ~v2 & new_n931_;
  assign new_n933_ = ~new_n930_ & ~new_n932_;
  assign new_n934_ = ~v6 & ~new_n933_;
  assign new_n935_ = ~v9 & new_n90_;
  assign new_n936_ = v3 & ~new_n935_;
  assign new_n937_ = ~v2 & ~new_n936_;
  assign new_n938_ = new_n147_ & new_n562_;
  assign new_n939_ = ~new_n937_ & ~new_n938_;
  assign new_n940_ = ~new_n934_ & new_n939_;
  assign new_n941_ = v7 & ~new_n940_;
  assign new_n942_ = ~v3 & ~v11;
  assign new_n943_ = new_n593_ & new_n942_;
  assign new_n944_ = ~new_n941_ & ~new_n943_;
  assign new_n945_ = ~new_n929_ & new_n944_;
  assign new_n946_ = v5 & ~new_n945_;
  assign new_n947_ = ~v11 & ~new_n48_;
  assign new_n948_ = ~new_n925_ & ~new_n947_;
  assign new_n949_ = ~v9 & ~new_n948_;
  assign new_n950_ = ~v2 & new_n949_;
  assign new_n951_ = v1 & new_n950_;
  assign new_n952_ = ~new_n946_ & ~new_n951_;
  assign new_n953_ = ~v13 & ~new_n952_;
  assign new_n954_ = ~v12 & new_n953_;
  assign new_n955_ = v8 & new_n954_;
  assign new_n956_ = ~new_n921_ & ~new_n955_;
  assign new_n957_ = ~v0 & ~new_n956_;
  assign new_n958_ = v0 & new_n180_;
  assign new_n959_ = ~new_n272_ & ~new_n958_;
  assign new_n960_ = ~v11 & ~new_n959_;
  assign new_n961_ = v10 & new_n960_;
  assign new_n962_ = v6 & new_n961_;
  assign new_n963_ = v3 & new_n962_;
  assign new_n964_ = ~v13 & ~new_n48_;
  assign new_n965_ = v11 & new_n964_;
  assign new_n966_ = ~v8 & new_n965_;
  assign new_n967_ = v0 & new_n966_;
  assign new_n968_ = ~new_n963_ & ~new_n967_;
  assign new_n969_ = ~v7 & ~new_n968_;
  assign new_n970_ = v6 & new_n147_;
  assign new_n971_ = ~new_n947_ & ~new_n970_;
  assign new_n972_ = ~v13 & ~new_n971_;
  assign new_n973_ = ~v8 & new_n972_;
  assign new_n974_ = v7 & new_n973_;
  assign new_n975_ = ~new_n969_ & ~new_n974_;
  assign new_n976_ = ~v1 & ~new_n975_;
  assign new_n977_ = v0 & new_n89_;
  assign new_n978_ = new_n597_ & new_n818_;
  assign new_n979_ = new_n977_ & new_n978_;
  assign new_n980_ = ~new_n976_ & ~new_n979_;
  assign new_n981_ = v5 & ~new_n980_;
  assign new_n982_ = ~v7 & ~v8;
  assign new_n983_ = v11 & ~new_n982_;
  assign new_n984_ = ~new_n48_ & ~new_n983_;
  assign new_n985_ = ~v3 & ~v8;
  assign new_n986_ = ~new_n984_ & ~new_n985_;
  assign new_n987_ = v13 & ~new_n986_;
  assign new_n988_ = v1 & new_n987_;
  assign new_n989_ = v0 & new_n988_;
  assign new_n990_ = ~new_n981_ & ~new_n989_;
  assign new_n991_ = ~v9 & ~new_n990_;
  assign new_n992_ = v7 & v9;
  assign new_n993_ = v5 & v11;
  assign new_n994_ = ~new_n992_ & ~new_n993_;
  assign new_n995_ = ~v13 & ~new_n994_;
  assign new_n996_ = ~v1 & new_n995_;
  assign new_n997_ = ~v11 & v13;
  assign new_n998_ = v1 & new_n997_;
  assign new_n999_ = ~new_n996_ & ~new_n998_;
  assign new_n1000_ = ~v8 & ~new_n999_;
  assign new_n1001_ = v8 & ~new_n931_;
  assign new_n1002_ = ~v5 & ~v7;
  assign new_n1003_ = ~new_n1001_ & new_n1002_;
  assign new_n1004_ = v13 & ~new_n1003_;
  assign new_n1005_ = v1 & new_n1004_;
  assign new_n1006_ = ~new_n1000_ & ~new_n1005_;
  assign new_n1007_ = v0 & ~new_n1006_;
  assign new_n1008_ = ~v1 & v5;
  assign new_n1009_ = v7 & new_n272_;
  assign new_n1010_ = new_n1008_ & new_n1009_;
  assign new_n1011_ = ~new_n1007_ & ~new_n1010_;
  assign new_n1012_ = ~v3 & ~new_n1011_;
  assign new_n1013_ = ~new_n991_ & ~new_n1012_;
  assign new_n1014_ = ~v2 & ~new_n1013_;
  assign new_n1015_ = v5 & v7;
  assign new_n1016_ = ~v0 & ~new_n1015_;
  assign new_n1017_ = ~new_n24_ & ~new_n1016_;
  assign new_n1018_ = v11 & new_n1017_;
  assign new_n1019_ = v6 & new_n90_;
  assign new_n1020_ = new_n553_ & new_n1019_;
  assign new_n1021_ = ~new_n1018_ & ~new_n1020_;
  assign new_n1022_ = ~v13 & ~new_n1021_;
  assign new_n1023_ = ~v1 & new_n1022_;
  assign new_n1024_ = v1 & new_n137_;
  assign new_n1025_ = new_n97_ & new_n997_;
  assign new_n1026_ = new_n1024_ & new_n1025_;
  assign new_n1027_ = ~new_n1023_ & ~new_n1026_;
  assign new_n1028_ = ~v8 & ~new_n1027_;
  assign new_n1029_ = ~v11 & ~new_n876_;
  assign new_n1030_ = ~new_n24_ & ~new_n1029_;
  assign new_n1031_ = v13 & new_n1030_;
  assign new_n1032_ = v1 & new_n1031_;
  assign new_n1033_ = v0 & new_n1032_;
  assign new_n1034_ = ~new_n1028_ & ~new_n1033_;
  assign new_n1035_ = v9 & ~new_n1034_;
  assign new_n1036_ = ~v3 & new_n1035_;
  assign new_n1037_ = ~new_n1014_ & ~new_n1036_;
  assign new_n1038_ = ~v12 & ~new_n1037_;
  assign new_n1039_ = ~new_n957_ & ~new_n1038_;
  assign new_n1040_ = ~new_n889_ & new_n1039_;
  assign new_n1041_ = ~v4 & ~new_n1040_;
  assign new_n1042_ = v7 & v12;
  assign new_n1043_ = v2 & new_n1042_;
  assign new_n1044_ = v6 & ~v7;
  assign new_n1045_ = ~v2 & v5;
  assign new_n1046_ = new_n1044_ & new_n1045_;
  assign new_n1047_ = v10 & ~v11;
  assign new_n1048_ = new_n720_ & new_n1047_;
  assign new_n1049_ = new_n1046_ & new_n1048_;
  assign new_n1050_ = ~new_n1043_ & ~new_n1049_;
  assign new_n1051_ = v3 & ~new_n1050_;
  assign new_n1052_ = ~v6 & ~v7;
  assign new_n1053_ = ~new_n357_ & ~new_n1052_;
  assign new_n1054_ = v0 & ~new_n1053_;
  assign new_n1055_ = v7 & ~new_n24_;
  assign new_n1056_ = ~v3 & new_n1055_;
  assign new_n1057_ = ~new_n1054_ & ~new_n1056_;
  assign new_n1058_ = ~v12 & ~new_n1057_;
  assign new_n1059_ = v11 & new_n1058_;
  assign new_n1060_ = ~v0 & v6;
  assign new_n1061_ = ~v7 & ~v10;
  assign new_n1062_ = new_n1060_ & new_n1061_;
  assign new_n1063_ = ~new_n1059_ & ~new_n1062_;
  assign new_n1064_ = ~v5 & ~new_n1063_;
  assign new_n1065_ = ~v3 & ~v6;
  assign new_n1066_ = v11 & ~v12;
  assign new_n1067_ = ~v10 & new_n1066_;
  assign new_n1068_ = new_n1065_ & new_n1067_;
  assign new_n1069_ = ~new_n1047_ & ~new_n1068_;
  assign new_n1070_ = v0 & ~new_n1069_;
  assign new_n1071_ = ~new_n98_ & ~new_n1070_;
  assign new_n1072_ = v5 & ~new_n1071_;
  assign new_n1073_ = v7 & new_n1066_;
  assign new_n1074_ = new_n1065_ & new_n1073_;
  assign new_n1075_ = ~new_n98_ & ~new_n1074_;
  assign new_n1076_ = ~v10 & ~new_n1075_;
  assign new_n1077_ = ~new_n1072_ & ~new_n1076_;
  assign new_n1078_ = ~new_n1064_ & new_n1077_;
  assign new_n1079_ = ~v13 & ~new_n1078_;
  assign new_n1080_ = v2 & new_n1079_;
  assign new_n1081_ = ~new_n1051_ & ~new_n1080_;
  assign new_n1082_ = ~v1 & ~new_n1081_;
  assign new_n1083_ = ~v0 & new_n115_;
  assign new_n1084_ = ~new_n23_ & ~new_n1083_;
  assign new_n1085_ = ~v13 & ~new_n244_;
  assign new_n1086_ = ~v12 & ~new_n1085_;
  assign new_n1087_ = ~new_n1084_ & ~new_n1086_;
  assign new_n1088_ = v1 & new_n764_;
  assign new_n1089_ = ~v3 & new_n43_;
  assign new_n1090_ = ~new_n1088_ & ~new_n1089_;
  assign new_n1091_ = ~v12 & ~new_n1090_;
  assign new_n1092_ = v10 & new_n1091_;
  assign new_n1093_ = ~v6 & new_n1092_;
  assign new_n1094_ = ~v0 & new_n1093_;
  assign new_n1095_ = v0 & v1;
  assign new_n1096_ = new_n23_ & new_n1095_;
  assign new_n1097_ = ~new_n1094_ & ~new_n1096_;
  assign new_n1098_ = ~v13 & ~new_n1097_;
  assign new_n1099_ = ~new_n1087_ & ~new_n1098_;
  assign new_n1100_ = v2 & ~new_n1099_;
  assign new_n1101_ = v0 & new_n115_;
  assign new_n1102_ = ~new_n23_ & ~new_n1101_;
  assign new_n1103_ = ~new_n48_ & ~new_n1102_;
  assign new_n1104_ = ~v7 & ~new_n635_;
  assign new_n1105_ = v11 & ~new_n1104_;
  assign new_n1106_ = v10 & new_n1105_;
  assign new_n1107_ = v6 & new_n1106_;
  assign new_n1108_ = ~new_n1103_ & ~new_n1107_;
  assign new_n1109_ = v13 & ~new_n1108_;
  assign new_n1110_ = ~v12 & new_n1109_;
  assign new_n1111_ = ~v2 & new_n1110_;
  assign new_n1112_ = ~new_n1100_ & ~new_n1111_;
  assign new_n1113_ = v5 & ~new_n1112_;
  assign new_n1114_ = ~new_n1082_ & ~new_n1113_;
  assign new_n1115_ = ~v9 & ~new_n1114_;
  assign new_n1116_ = ~v1 & v3;
  assign new_n1117_ = new_n764_ & new_n1116_;
  assign new_n1118_ = ~new_n43_ & ~new_n1117_;
  assign new_n1119_ = v13 & ~new_n1118_;
  assign new_n1120_ = ~v2 & new_n1119_;
  assign new_n1121_ = v0 & new_n1120_;
  assign new_n1122_ = ~v0 & v2;
  assign new_n1123_ = v11 & ~v13;
  assign new_n1124_ = v7 & new_n1123_;
  assign new_n1125_ = new_n1122_ & new_n1124_;
  assign new_n1126_ = ~new_n1121_ & ~new_n1125_;
  assign new_n1127_ = v6 & ~new_n1126_;
  assign new_n1128_ = v1 & v2;
  assign new_n1129_ = ~v0 & new_n1128_;
  assign new_n1130_ = ~v11 & ~v13;
  assign new_n1131_ = new_n825_ & new_n1130_;
  assign new_n1132_ = new_n1129_ & new_n1131_;
  assign new_n1133_ = ~new_n1127_ & ~new_n1132_;
  assign new_n1134_ = v10 & ~new_n1133_;
  assign new_n1135_ = ~v13 & ~new_n1090_;
  assign new_n1136_ = ~v6 & new_n1135_;
  assign new_n1137_ = v2 & new_n1136_;
  assign new_n1138_ = ~v0 & new_n1137_;
  assign new_n1139_ = ~new_n1134_ & ~new_n1138_;
  assign new_n1140_ = ~v12 & ~new_n1139_;
  assign new_n1141_ = v9 & new_n1140_;
  assign new_n1142_ = ~v0 & new_n637_;
  assign new_n1143_ = new_n24_ & new_n1130_;
  assign new_n1144_ = new_n1142_ & new_n1143_;
  assign new_n1145_ = ~new_n1141_ & ~new_n1144_;
  assign new_n1146_ = ~v5 & ~new_n1145_;
  assign new_n1147_ = v1 & new_n792_;
  assign new_n1148_ = new_n803_ & new_n1015_;
  assign new_n1149_ = new_n1147_ & new_n1148_;
  assign new_n1150_ = ~new_n1146_ & ~new_n1149_;
  assign new_n1151_ = ~new_n1115_ & new_n1150_;
  assign new_n1152_ = v4 & ~new_n1151_;
  assign new_n1153_ = v5 & new_n1042_;
  assign new_n1154_ = new_n637_ & new_n1153_;
  assign new_n1155_ = ~v2 & v6;
  assign new_n1156_ = new_n701_ & new_n1155_;
  assign new_n1157_ = v11 & new_n720_;
  assign new_n1158_ = new_n61_ & new_n1157_;
  assign new_n1159_ = new_n1156_ & new_n1158_;
  assign new_n1160_ = ~new_n1154_ & ~new_n1159_;
  assign new_n1161_ = v3 & ~new_n1160_;
  assign new_n1162_ = ~v7 & ~v9;
  assign new_n1163_ = v11 & ~new_n1162_;
  assign new_n1164_ = v1 & new_n742_;
  assign new_n1165_ = v0 & new_n1164_;
  assign new_n1166_ = ~v0 & ~v1;
  assign new_n1167_ = new_n744_ & new_n1166_;
  assign new_n1168_ = ~new_n1165_ & ~new_n1167_;
  assign new_n1169_ = ~new_n1163_ & ~new_n1168_;
  assign new_n1170_ = ~v5 & new_n1169_;
  assign new_n1171_ = ~new_n115_ & ~new_n344_;
  assign new_n1172_ = ~v3 & new_n1171_;
  assign new_n1173_ = new_n89_ & new_n147_;
  assign new_n1174_ = ~new_n947_ & ~new_n1173_;
  assign new_n1175_ = ~v9 & ~new_n1174_;
  assign new_n1176_ = ~new_n1172_ & ~new_n1175_;
  assign new_n1177_ = v13 & ~new_n1176_;
  assign new_n1178_ = ~v12 & new_n1177_;
  assign new_n1179_ = ~v2 & new_n1178_;
  assign new_n1180_ = v1 & new_n1179_;
  assign new_n1181_ = ~v11 & v12;
  assign new_n1182_ = ~v9 & new_n1181_;
  assign new_n1183_ = new_n637_ & new_n1182_;
  assign new_n1184_ = ~new_n1180_ & ~new_n1183_;
  assign new_n1185_ = ~new_n1170_ & new_n1184_;
  assign new_n1186_ = ~new_n1161_ & new_n1185_;
  assign new_n1187_ = ~new_n1152_ & new_n1186_;
  assign new_n1188_ = ~v8 & ~new_n1187_;
  assign new_n1189_ = v5 & new_n202_;
  assign new_n1190_ = ~v5 & ~v10;
  assign new_n1191_ = ~new_n1189_ & ~new_n1190_;
  assign new_n1192_ = v1 & ~new_n1191_;
  assign new_n1193_ = ~v5 & ~new_n48_;
  assign new_n1194_ = ~new_n202_ & ~new_n1193_;
  assign new_n1195_ = v7 & ~new_n1194_;
  assign new_n1196_ = ~new_n1192_ & ~new_n1195_;
  assign new_n1197_ = ~v0 & ~new_n1196_;
  assign new_n1198_ = ~v6 & new_n97_;
  assign new_n1199_ = new_n1008_ & new_n1198_;
  assign new_n1200_ = ~new_n1197_ & ~new_n1199_;
  assign new_n1201_ = v9 & ~new_n1200_;
  assign new_n1202_ = ~v1 & ~v5;
  assign new_n1203_ = v7 & ~v9;
  assign new_n1204_ = ~v6 & new_n1203_;
  assign new_n1205_ = new_n1202_ & new_n1204_;
  assign new_n1206_ = ~new_n1201_ & ~new_n1205_;
  assign new_n1207_ = ~v2 & ~new_n1206_;
  assign new_n1208_ = ~v7 & v9;
  assign new_n1209_ = ~v6 & new_n1208_;
  assign new_n1210_ = new_n701_ & new_n1209_;
  assign new_n1211_ = ~v1 & v6;
  assign new_n1212_ = v7 & new_n140_;
  assign new_n1213_ = new_n1211_ & new_n1212_;
  assign new_n1214_ = ~new_n1210_ & ~new_n1213_;
  assign new_n1215_ = ~v5 & ~new_n1214_;
  assign new_n1216_ = ~new_n1207_ & ~new_n1215_;
  assign new_n1217_ = ~v11 & ~new_n1216_;
  assign new_n1218_ = ~v9 & ~new_n314_;
  assign new_n1219_ = ~v5 & new_n1218_;
  assign new_n1220_ = v5 & ~v6;
  assign new_n1221_ = new_n203_ & new_n1220_;
  assign new_n1222_ = ~new_n1219_ & ~new_n1221_;
  assign new_n1223_ = v11 & ~new_n1222_;
  assign new_n1224_ = ~v7 & new_n1223_;
  assign new_n1225_ = ~v1 & new_n1224_;
  assign new_n1226_ = v0 & new_n1225_;
  assign new_n1227_ = ~new_n1217_ & ~new_n1226_;
  assign new_n1228_ = ~v12 & ~new_n1227_;
  assign new_n1229_ = v0 & ~new_n193_;
  assign new_n1230_ = ~v6 & ~new_n1229_;
  assign new_n1231_ = v7 & ~new_n1230_;
  assign new_n1232_ = ~v0 & ~new_n244_;
  assign new_n1233_ = ~new_n1231_ & ~new_n1232_;
  assign new_n1234_ = v11 & ~new_n1233_;
  assign new_n1235_ = ~v11 & ~new_n379_;
  assign new_n1236_ = ~v7 & new_n1235_;
  assign new_n1237_ = ~v1 & new_n1236_;
  assign new_n1238_ = ~new_n1234_ & ~new_n1237_;
  assign new_n1239_ = v5 & ~new_n1238_;
  assign new_n1240_ = ~v1 & new_n1002_;
  assign new_n1241_ = ~v11 & ~new_n1240_;
  assign new_n1242_ = v10 & ~new_n1241_;
  assign new_n1243_ = v6 & new_n1242_;
  assign new_n1244_ = ~v0 & new_n1243_;
  assign new_n1245_ = ~new_n1239_ & ~new_n1244_;
  assign new_n1246_ = v9 & ~new_n1245_;
  assign new_n1247_ = v0 & v2;
  assign new_n1248_ = new_n1015_ & new_n1247_;
  assign new_n1249_ = v6 & v11;
  assign new_n1250_ = ~v5 & new_n1249_;
  assign new_n1251_ = new_n1166_ & new_n1250_;
  assign new_n1252_ = ~new_n1248_ & ~new_n1251_;
  assign new_n1253_ = v10 & ~new_n1252_;
  assign new_n1254_ = ~new_n1246_ & ~new_n1253_;
  assign new_n1255_ = ~new_n1228_ & new_n1254_;
  assign new_n1256_ = v8 & ~new_n1255_;
  assign new_n1257_ = ~v10 & v11;
  assign new_n1258_ = new_n699_ & new_n1257_;
  assign new_n1259_ = new_n701_ & new_n1047_;
  assign new_n1260_ = ~new_n1258_ & ~new_n1259_;
  assign new_n1261_ = ~v12 & ~new_n1260_;
  assign new_n1262_ = ~v7 & new_n1261_;
  assign new_n1263_ = ~v6 & new_n1262_;
  assign new_n1264_ = v7 & v10;
  assign new_n1265_ = v0 & new_n1264_;
  assign new_n1266_ = ~new_n1232_ & ~new_n1265_;
  assign new_n1267_ = v11 & ~new_n1266_;
  assign new_n1268_ = ~v1 & new_n1047_;
  assign new_n1269_ = ~new_n817_ & ~new_n1268_;
  assign new_n1270_ = v0 & ~new_n1269_;
  assign new_n1271_ = ~v7 & ~new_n306_;
  assign new_n1272_ = v6 & ~new_n1271_;
  assign new_n1273_ = new_n90_ & new_n817_;
  assign new_n1274_ = ~new_n1272_ & ~new_n1273_;
  assign new_n1275_ = ~new_n1270_ & new_n1274_;
  assign new_n1276_ = ~new_n1267_ & new_n1275_;
  assign new_n1277_ = ~new_n1263_ & new_n1276_;
  assign new_n1278_ = v5 & ~new_n1277_;
  assign new_n1279_ = v7 & ~new_n178_;
  assign new_n1280_ = ~new_n260_ & ~new_n1202_;
  assign new_n1281_ = ~v0 & ~new_n1280_;
  assign new_n1282_ = ~v1 & new_n931_;
  assign new_n1283_ = ~new_n1281_ & ~new_n1282_;
  assign new_n1284_ = ~new_n1279_ & new_n1283_;
  assign new_n1285_ = v6 & ~new_n1284_;
  assign new_n1286_ = ~new_n1278_ & ~new_n1285_;
  assign new_n1287_ = v2 & ~new_n1286_;
  assign new_n1288_ = ~new_n1256_ & ~new_n1287_;
  assign new_n1289_ = ~v13 & ~new_n1288_;
  assign new_n1290_ = ~v11 & ~new_n344_;
  assign new_n1291_ = ~v1 & new_n1290_;
  assign new_n1292_ = ~v7 & ~new_n305_;
  assign new_n1293_ = v5 & ~new_n1292_;
  assign new_n1294_ = ~v11 & ~new_n857_;
  assign new_n1295_ = v9 & ~new_n1294_;
  assign new_n1296_ = ~v0 & new_n1295_;
  assign new_n1297_ = ~new_n1293_ & ~new_n1296_;
  assign new_n1298_ = ~new_n1291_ & new_n1297_;
  assign new_n1299_ = v2 & ~new_n1298_;
  assign new_n1300_ = ~v1 & new_n764_;
  assign new_n1301_ = ~new_n43_ & ~new_n1300_;
  assign new_n1302_ = v9 & ~new_n1301_;
  assign new_n1303_ = v8 & new_n1302_;
  assign new_n1304_ = v5 & new_n1303_;
  assign new_n1305_ = ~new_n1299_ & ~new_n1304_;
  assign new_n1306_ = v12 & ~new_n1305_;
  assign new_n1307_ = ~new_n1289_ & ~new_n1306_;
  assign new_n1308_ = v3 & ~new_n1307_;
  assign new_n1309_ = v1 & new_n66_;
  assign new_n1310_ = ~new_n54_ & ~new_n1309_;
  assign new_n1311_ = new_n115_ & new_n1122_;
  assign new_n1312_ = ~new_n23_ & ~new_n1311_;
  assign new_n1313_ = ~new_n1310_ & ~new_n1312_;
  assign new_n1314_ = v9 & ~v11;
  assign new_n1315_ = v5 & new_n1314_;
  assign new_n1316_ = new_n637_ & new_n1315_;
  assign new_n1317_ = ~new_n1313_ & ~new_n1316_;
  assign new_n1318_ = ~v10 & ~new_n1317_;
  assign new_n1319_ = v6 & new_n1318_;
  assign new_n1320_ = ~new_n43_ & ~new_n1088_;
  assign new_n1321_ = ~new_n24_ & ~new_n1320_;
  assign new_n1322_ = v9 & new_n1321_;
  assign new_n1323_ = v5 & new_n1322_;
  assign new_n1324_ = ~new_n1319_ & ~new_n1323_;
  assign new_n1325_ = v8 & ~new_n1324_;
  assign new_n1326_ = v9 & ~new_n764_;
  assign new_n1327_ = v1 & ~v5;
  assign new_n1328_ = ~new_n993_ & ~new_n1327_;
  assign new_n1329_ = ~new_n1326_ & new_n1328_;
  assign new_n1330_ = v0 & ~new_n1329_;
  assign new_n1331_ = v5 & ~new_n110_;
  assign new_n1332_ = ~v9 & ~new_n115_;
  assign new_n1333_ = v1 & new_n1332_;
  assign new_n1334_ = ~new_n1331_ & ~new_n1333_;
  assign new_n1335_ = ~new_n1330_ & new_n1334_;
  assign new_n1336_ = ~v2 & ~new_n1335_;
  assign new_n1337_ = ~new_n1325_ & ~new_n1336_;
  assign new_n1338_ = v13 & ~new_n1337_;
  assign new_n1339_ = ~v12 & new_n1338_;
  assign new_n1340_ = ~v3 & new_n1339_;
  assign new_n1341_ = ~new_n1308_ & ~new_n1340_;
  assign new_n1342_ = v4 & ~new_n1341_;
  assign new_n1343_ = new_n635_ & new_n1153_;
  assign new_n1344_ = ~v3 & v6;
  assign new_n1345_ = new_n699_ & new_n1344_;
  assign new_n1346_ = ~v11 & new_n720_;
  assign new_n1347_ = new_n203_ & new_n1346_;
  assign new_n1348_ = new_n1345_ & new_n1347_;
  assign new_n1349_ = ~new_n1343_ & ~new_n1348_;
  assign new_n1350_ = v2 & ~new_n1349_;
  assign new_n1351_ = ~v11 & ~new_n1208_;
  assign new_n1352_ = v0 & new_n771_;
  assign new_n1353_ = new_n772_ & new_n1166_;
  assign new_n1354_ = ~new_n1352_ & ~new_n1353_;
  assign new_n1355_ = ~new_n1351_ & ~new_n1354_;
  assign new_n1356_ = ~v5 & new_n1355_;
  assign new_n1357_ = ~new_n66_ & ~new_n764_;
  assign new_n1358_ = ~v2 & new_n1357_;
  assign new_n1359_ = v11 & ~new_n24_;
  assign new_n1360_ = new_n89_ & new_n90_;
  assign new_n1361_ = ~new_n1359_ & ~new_n1360_;
  assign new_n1362_ = v9 & ~new_n1361_;
  assign new_n1363_ = ~new_n1358_ & ~new_n1362_;
  assign new_n1364_ = v13 & ~new_n1363_;
  assign new_n1365_ = ~v12 & new_n1364_;
  assign new_n1366_ = ~v3 & new_n1365_;
  assign new_n1367_ = v0 & new_n1366_;
  assign new_n1368_ = v11 & v12;
  assign new_n1369_ = v9 & new_n1368_;
  assign new_n1370_ = new_n635_ & new_n1369_;
  assign new_n1371_ = ~new_n1367_ & ~new_n1370_;
  assign new_n1372_ = ~new_n1356_ & new_n1371_;
  assign new_n1373_ = ~new_n1350_ & new_n1372_;
  assign new_n1374_ = v8 & ~new_n1373_;
  assign new_n1375_ = ~new_n1342_ & ~new_n1374_;
  assign new_n1376_ = ~new_n1188_ & new_n1375_;
  assign new_n1377_ = ~new_n1041_ & new_n1376_;
  assign new_n1378_ = ~new_n791_ & new_n1377_;
  assign new_n1379_ = ~new_n763_ & new_n1378_;
  assign \v15.6  = v14 & ~new_n1379_;
endmodule


