// Benchmark "multiplier" written by ABC on Fri Sep 15 11:23:43 2023

module multiplier ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257_, new_n258_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_,
    new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_,
    new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_,
    new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_,
    new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_,
    new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_,
    new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_,
    new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_,
    new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_,
    new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_,
    new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_,
    new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_,
    new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_,
    new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_,
    new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2304_, new_n2305_, new_n2306_, new_n2307_,
    new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_,
    new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_,
    new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_,
    new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_,
    new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_,
    new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_,
    new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_,
    new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_,
    new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_,
    new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_,
    new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_,
    new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_,
    new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_,
    new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_,
    new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_,
    new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_,
    new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_,
    new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_,
    new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_,
    new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_,
    new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_,
    new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_,
    new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_,
    new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_,
    new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_,
    new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_,
    new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_,
    new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_,
    new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_,
    new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_,
    new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_,
    new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_,
    new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_,
    new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_,
    new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_,
    new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_,
    new_n3031_, new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_,
    new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_,
    new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_,
    new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_,
    new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_,
    new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_,
    new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_,
    new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_,
    new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_,
    new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_,
    new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_,
    new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_,
    new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_,
    new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_,
    new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_,
    new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_,
    new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_,
    new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_,
    new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_,
    new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_,
    new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_,
    new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_,
    new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_,
    new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_,
    new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_,
    new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_,
    new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_,
    new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_,
    new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_,
    new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_,
    new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_,
    new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_,
    new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_,
    new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_,
    new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_,
    new_n3399_, new_n3400_, new_n3401_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_,
    new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_,
    new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_,
    new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_,
    new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_,
    new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_,
    new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_,
    new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_,
    new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_,
    new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_,
    new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_,
    new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3616_,
    new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_,
    new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_,
    new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_,
    new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_,
    new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_,
    new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_,
    new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_,
    new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_,
    new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_,
    new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_,
    new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_,
    new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_,
    new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_,
    new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_,
    new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_,
    new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_,
    new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_,
    new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_,
    new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_,
    new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_,
    new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_,
    new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_,
    new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_,
    new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_,
    new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_,
    new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_,
    new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_,
    new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4020_,
    new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_,
    new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_,
    new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_,
    new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_,
    new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_,
    new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_,
    new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_,
    new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_,
    new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_,
    new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_,
    new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_,
    new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_,
    new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_,
    new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_,
    new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_,
    new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_,
    new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_,
    new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_,
    new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_,
    new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_,
    new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4210_, new_n4211_, new_n4212_, new_n4213_,
    new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_,
    new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_,
    new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_,
    new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_,
    new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_,
    new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_,
    new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_,
    new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_,
    new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_,
    new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_,
    new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_,
    new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_,
    new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_,
    new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4399_, new_n4400_,
    new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4406_,
    new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_, new_n4412_,
    new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_, new_n4418_,
    new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_, new_n4424_,
    new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_, new_n4430_,
    new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_,
    new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_,
    new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_,
    new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_,
    new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_,
    new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_,
    new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_,
    new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_,
    new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_,
    new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_,
    new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_,
    new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_,
    new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_,
    new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_,
    new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_,
    new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_,
    new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_,
    new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_,
    new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_,
    new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_,
    new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_,
    new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_,
    new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_,
    new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_,
    new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_,
    new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_,
    new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_,
    new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_,
    new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_,
    new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_,
    new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_,
    new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4664_, new_n4665_,
    new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_,
    new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_,
    new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_,
    new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_,
    new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_,
    new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_,
    new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_,
    new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_,
    new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_,
    new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_,
    new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_,
    new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_,
    new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_,
    new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_,
    new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_,
    new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_,
    new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_,
    new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_,
    new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_,
    new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_,
    new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_,
    new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_,
    new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_,
    new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_,
    new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_,
    new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_,
    new_n4876_, new_n4877_, new_n4878_, new_n4880_, new_n4881_, new_n4882_,
    new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_,
    new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_,
    new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_,
    new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_,
    new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_,
    new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_,
    new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_,
    new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_,
    new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_,
    new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_,
    new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_,
    new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_,
    new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_,
    new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_,
    new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_,
    new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_,
    new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_,
    new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_,
    new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_,
    new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_,
    new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_,
    new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_,
    new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_,
    new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_,
    new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_,
    new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_,
    new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_,
    new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_,
    new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_,
    new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_,
    new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_,
    new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_,
    new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_,
    new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_,
    new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5338_, new_n5339_, new_n5340_,
    new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_,
    new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_,
    new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_,
    new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_,
    new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_,
    new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_,
    new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_,
    new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_,
    new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_,
    new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_,
    new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_,
    new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_,
    new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_,
    new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_,
    new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_,
    new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_,
    new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_,
    new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_,
    new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_,
    new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_,
    new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_,
    new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_,
    new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_,
    new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_,
    new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_,
    new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_,
    new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_,
    new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_,
    new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_,
    new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_,
    new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_,
    new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_,
    new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_,
    new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_,
    new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_,
    new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_,
    new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_,
    new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_,
    new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_,
    new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_,
    new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_,
    new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_,
    new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_,
    new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_,
    new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_,
    new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_,
    new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_,
    new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_,
    new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_,
    new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_,
    new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_,
    new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_,
    new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_,
    new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_,
    new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_,
    new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_,
    new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_,
    new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_,
    new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_,
    new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_,
    new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_,
    new_n5774_, new_n5775_, new_n5776_, new_n5778_, new_n5779_, new_n5780_,
    new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_,
    new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_,
    new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_,
    new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_, new_n5804_,
    new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_,
    new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_,
    new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_,
    new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_,
    new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_,
    new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_,
    new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_,
    new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_,
    new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_,
    new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_,
    new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_,
    new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_,
    new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_,
    new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_,
    new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_,
    new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_,
    new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_,
    new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_,
    new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_,
    new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_,
    new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_,
    new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_,
    new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_,
    new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_,
    new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_,
    new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_,
    new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_,
    new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_,
    new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_,
    new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_,
    new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_,
    new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_,
    new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_,
    new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_,
    new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_,
    new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_,
    new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_,
    new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_,
    new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_,
    new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6045_,
    new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_,
    new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_,
    new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_,
    new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_,
    new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_,
    new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_,
    new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_,
    new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_,
    new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_,
    new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_,
    new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_,
    new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_,
    new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_,
    new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_,
    new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_,
    new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_,
    new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_,
    new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_,
    new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_,
    new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_,
    new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_,
    new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_,
    new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_,
    new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_,
    new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_,
    new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_,
    new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_,
    new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_,
    new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_,
    new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_,
    new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_,
    new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_,
    new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_,
    new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_,
    new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_,
    new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_,
    new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_,
    new_n6292_, new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_,
    new_n6298_, new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_,
    new_n6304_, new_n6305_, new_n6307_, new_n6308_, new_n6309_, new_n6310_,
    new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_,
    new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_,
    new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_,
    new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_,
    new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_,
    new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_,
    new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_,
    new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_,
    new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_,
    new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_,
    new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_,
    new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_,
    new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_,
    new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_,
    new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_,
    new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_,
    new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_,
    new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_,
    new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_,
    new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_,
    new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_,
    new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_,
    new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_,
    new_n6455_, new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_,
    new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_,
    new_n6467_, new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_,
    new_n6473_, new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_,
    new_n6479_, new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_,
    new_n6485_, new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_,
    new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_,
    new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_,
    new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_,
    new_n6509_, new_n6510_, new_n6512_, new_n6513_, new_n6514_, new_n6515_,
    new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_,
    new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_,
    new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_,
    new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_,
    new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_,
    new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_,
    new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_,
    new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_,
    new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_,
    new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_,
    new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_,
    new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_,
    new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_,
    new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_,
    new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_,
    new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_,
    new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_,
    new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_,
    new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_,
    new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_,
    new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_,
    new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_,
    new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_,
    new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_,
    new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_,
    new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_,
    new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_,
    new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_,
    new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_,
    new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_,
    new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_,
    new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_,
    new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_,
    new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_,
    new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_,
    new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_,
    new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_,
    new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_,
    new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_,
    new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_,
    new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_,
    new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_,
    new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_,
    new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_,
    new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_,
    new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_,
    new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_,
    new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_,
    new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_,
    new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_,
    new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_,
    new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_,
    new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_,
    new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_,
    new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_,
    new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_,
    new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_,
    new_n7087_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_,
    new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_,
    new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_,
    new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_,
    new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_,
    new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_,
    new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_,
    new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_,
    new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_,
    new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_,
    new_n7322_, new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_,
    new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_,
    new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_,
    new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_,
    new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_,
    new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_,
    new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_,
    new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_,
    new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_,
    new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_,
    new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_,
    new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_,
    new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_,
    new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_,
    new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_,
    new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_,
    new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_,
    new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_,
    new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_,
    new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_,
    new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_,
    new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_,
    new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_,
    new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_,
    new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_,
    new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_,
    new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_,
    new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_,
    new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_,
    new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_,
    new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_,
    new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_,
    new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_,
    new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_,
    new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_,
    new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_,
    new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_,
    new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_,
    new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_,
    new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_,
    new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_,
    new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_,
    new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_,
    new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_,
    new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_,
    new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_,
    new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_,
    new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_,
    new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_,
    new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_,
    new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_,
    new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_,
    new_n7635_, new_n7636_, new_n7637_, new_n7639_, new_n7640_, new_n7641_,
    new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_,
    new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_,
    new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_,
    new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_,
    new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_,
    new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_,
    new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_,
    new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_,
    new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_,
    new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_,
    new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_,
    new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_,
    new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_,
    new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_,
    new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_,
    new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_,
    new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_,
    new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_,
    new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_,
    new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_,
    new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_,
    new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_,
    new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_,
    new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_,
    new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_,
    new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_,
    new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_,
    new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_,
    new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_,
    new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_,
    new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_,
    new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_,
    new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_,
    new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_,
    new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_,
    new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_,
    new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_,
    new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_,
    new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_,
    new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_,
    new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_,
    new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_,
    new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_,
    new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_,
    new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_,
    new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_,
    new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_,
    new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_,
    new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_,
    new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_,
    new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_,
    new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_,
    new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_,
    new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_,
    new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_,
    new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_,
    new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_,
    new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_,
    new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_,
    new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_,
    new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_,
    new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_,
    new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_,
    new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_,
    new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_,
    new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_,
    new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_,
    new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_,
    new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_,
    new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_,
    new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_,
    new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8489_, new_n8490_,
    new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_,
    new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_,
    new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_,
    new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_,
    new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_,
    new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_,
    new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_,
    new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_,
    new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_,
    new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_,
    new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_,
    new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_,
    new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_,
    new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_,
    new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_,
    new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_,
    new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_,
    new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_,
    new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_,
    new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_,
    new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_,
    new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_,
    new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_,
    new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_,
    new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_,
    new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_,
    new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_,
    new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_,
    new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_,
    new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_,
    new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_,
    new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_,
    new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_,
    new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_,
    new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_,
    new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_,
    new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_,
    new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_,
    new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_,
    new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_,
    new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_,
    new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_,
    new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_,
    new_n8767_, new_n8768_, new_n8769_, new_n8771_, new_n8772_, new_n8773_,
    new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_,
    new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_,
    new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_,
    new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_,
    new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_,
    new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_,
    new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_, new_n8821_,
    new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_,
    new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_,
    new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_,
    new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_,
    new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_,
    new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_,
    new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_,
    new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_,
    new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_,
    new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_,
    new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_,
    new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_,
    new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_,
    new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_,
    new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_,
    new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_,
    new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_,
    new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_,
    new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_,
    new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_,
    new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_,
    new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_,
    new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_,
    new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_,
    new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_,
    new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_,
    new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_,
    new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_,
    new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_,
    new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_,
    new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_,
    new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_,
    new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_,
    new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_,
    new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_,
    new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_,
    new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_,
    new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_,
    new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_,
    new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_,
    new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_,
    new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_,
    new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_,
    new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_,
    new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_,
    new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_,
    new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_,
    new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_,
    new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_,
    new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_,
    new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_,
    new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_,
    new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_,
    new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_,
    new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_,
    new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_,
    new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_,
    new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9374_, new_n9375_,
    new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_,
    new_n9382_, new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_,
    new_n9388_, new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_,
    new_n9394_, new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_,
    new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_,
    new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_,
    new_n9412_, new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_,
    new_n9418_, new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_,
    new_n9424_, new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_,
    new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_,
    new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_,
    new_n9442_, new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_,
    new_n9448_, new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_,
    new_n9454_, new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_,
    new_n9460_, new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_,
    new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_,
    new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_,
    new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_,
    new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_,
    new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_,
    new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_,
    new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_,
    new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_, new_n9513_,
    new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_,
    new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_, new_n9525_,
    new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_, new_n9531_,
    new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_,
    new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_, new_n9543_,
    new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_, new_n9549_,
    new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_, new_n9555_,
    new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_, new_n9561_,
    new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_, new_n9567_,
    new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_, new_n9573_,
    new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_, new_n9579_,
    new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_, new_n9585_,
    new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_, new_n9591_,
    new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_, new_n9597_,
    new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_, new_n9603_,
    new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_,
    new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_,
    new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_,
    new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_,
    new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_,
    new_n9634_, new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_,
    new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_,
    new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_,
    new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_,
    new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_,
    new_n9664_, new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_,
    new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_,
    new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_,
    new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_,
    new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_,
    new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_,
    new_n9700_, new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_,
    new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_,
    new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_,
    new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_,
    new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_,
    new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_,
    new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_,
    new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_,
    new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_, new_n9754_,
    new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_,
    new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_,
    new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_,
    new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_,
    new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_,
    new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_,
    new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_, new_n9796_,
    new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_,
    new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_,
    new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_,
    new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_,
    new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_,
    new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_,
    new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_,
    new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_,
    new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_,
    new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_,
    new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_,
    new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_,
    new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_,
    new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_,
    new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_,
    new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_,
    new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_,
    new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_,
    new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_,
    new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_,
    new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_,
    new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_,
    new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_,
    new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_,
    new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_,
    new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_,
    new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_,
    new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_,
    new_n9965_, new_n9966_, new_n9967_, new_n9969_, new_n9970_, new_n9971_,
    new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_,
    new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10068_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10078_, new_n10079_, new_n10080_,
    new_n10081_, new_n10082_, new_n10083_, new_n10084_, new_n10085_,
    new_n10086_, new_n10087_, new_n10088_, new_n10089_, new_n10090_,
    new_n10091_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10202_, new_n10203_, new_n10204_, new_n10205_,
    new_n10206_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10294_, new_n10295_, new_n10296_,
    new_n10297_, new_n10298_, new_n10299_, new_n10300_, new_n10301_,
    new_n10302_, new_n10303_, new_n10304_, new_n10305_, new_n10306_,
    new_n10307_, new_n10308_, new_n10309_, new_n10310_, new_n10311_,
    new_n10312_, new_n10313_, new_n10314_, new_n10315_, new_n10316_,
    new_n10317_, new_n10318_, new_n10319_, new_n10320_, new_n10321_,
    new_n10322_, new_n10323_, new_n10324_, new_n10325_, new_n10326_,
    new_n10327_, new_n10328_, new_n10329_, new_n10330_, new_n10331_,
    new_n10332_, new_n10333_, new_n10334_, new_n10335_, new_n10336_,
    new_n10337_, new_n10338_, new_n10339_, new_n10340_, new_n10341_,
    new_n10342_, new_n10343_, new_n10344_, new_n10345_, new_n10346_,
    new_n10347_, new_n10348_, new_n10349_, new_n10350_, new_n10351_,
    new_n10352_, new_n10353_, new_n10354_, new_n10355_, new_n10356_,
    new_n10357_, new_n10358_, new_n10359_, new_n10360_, new_n10361_,
    new_n10362_, new_n10363_, new_n10364_, new_n10365_, new_n10366_,
    new_n10367_, new_n10368_, new_n10369_, new_n10370_, new_n10371_,
    new_n10372_, new_n10373_, new_n10374_, new_n10375_, new_n10376_,
    new_n10377_, new_n10378_, new_n10379_, new_n10380_, new_n10381_,
    new_n10382_, new_n10383_, new_n10384_, new_n10385_, new_n10386_,
    new_n10387_, new_n10388_, new_n10389_, new_n10390_, new_n10391_,
    new_n10392_, new_n10393_, new_n10394_, new_n10395_, new_n10396_,
    new_n10397_, new_n10398_, new_n10399_, new_n10400_, new_n10401_,
    new_n10402_, new_n10403_, new_n10404_, new_n10405_, new_n10406_,
    new_n10407_, new_n10408_, new_n10409_, new_n10410_, new_n10411_,
    new_n10412_, new_n10413_, new_n10414_, new_n10415_, new_n10416_,
    new_n10417_, new_n10418_, new_n10419_, new_n10420_, new_n10421_,
    new_n10422_, new_n10423_, new_n10424_, new_n10425_, new_n10426_,
    new_n10427_, new_n10428_, new_n10429_, new_n10430_, new_n10431_,
    new_n10432_, new_n10433_, new_n10434_, new_n10435_, new_n10436_,
    new_n10437_, new_n10438_, new_n10439_, new_n10440_, new_n10441_,
    new_n10442_, new_n10443_, new_n10444_, new_n10445_, new_n10446_,
    new_n10447_, new_n10448_, new_n10449_, new_n10450_, new_n10451_,
    new_n10452_, new_n10453_, new_n10454_, new_n10455_, new_n10456_,
    new_n10457_, new_n10458_, new_n10459_, new_n10460_, new_n10461_,
    new_n10462_, new_n10463_, new_n10464_, new_n10465_, new_n10466_,
    new_n10467_, new_n10468_, new_n10469_, new_n10470_, new_n10471_,
    new_n10472_, new_n10473_, new_n10474_, new_n10475_, new_n10476_,
    new_n10477_, new_n10478_, new_n10479_, new_n10480_, new_n10481_,
    new_n10482_, new_n10483_, new_n10484_, new_n10485_, new_n10486_,
    new_n10487_, new_n10488_, new_n10489_, new_n10490_, new_n10491_,
    new_n10492_, new_n10493_, new_n10494_, new_n10495_, new_n10496_,
    new_n10497_, new_n10498_, new_n10499_, new_n10500_, new_n10501_,
    new_n10502_, new_n10503_, new_n10504_, new_n10505_, new_n10506_,
    new_n10507_, new_n10508_, new_n10509_, new_n10510_, new_n10511_,
    new_n10512_, new_n10513_, new_n10514_, new_n10515_, new_n10516_,
    new_n10517_, new_n10518_, new_n10519_, new_n10520_, new_n10521_,
    new_n10522_, new_n10523_, new_n10524_, new_n10525_, new_n10526_,
    new_n10527_, new_n10528_, new_n10529_, new_n10530_, new_n10531_,
    new_n10532_, new_n10533_, new_n10534_, new_n10535_, new_n10536_,
    new_n10537_, new_n10538_, new_n10539_, new_n10540_, new_n10541_,
    new_n10542_, new_n10543_, new_n10544_, new_n10545_, new_n10546_,
    new_n10547_, new_n10548_, new_n10549_, new_n10550_, new_n10551_,
    new_n10552_, new_n10553_, new_n10554_, new_n10555_, new_n10556_,
    new_n10557_, new_n10558_, new_n10559_, new_n10560_, new_n10561_,
    new_n10562_, new_n10563_, new_n10564_, new_n10565_, new_n10566_,
    new_n10567_, new_n10568_, new_n10569_, new_n10570_, new_n10571_,
    new_n10572_, new_n10573_, new_n10574_, new_n10575_, new_n10576_,
    new_n10577_, new_n10578_, new_n10579_, new_n10580_, new_n10581_,
    new_n10582_, new_n10583_, new_n10584_, new_n10585_, new_n10586_,
    new_n10587_, new_n10588_, new_n10589_, new_n10590_, new_n10591_,
    new_n10592_, new_n10593_, new_n10594_, new_n10595_, new_n10596_,
    new_n10597_, new_n10598_, new_n10599_, new_n10600_, new_n10601_,
    new_n10602_, new_n10603_, new_n10604_, new_n10605_, new_n10606_,
    new_n10607_, new_n10608_, new_n10609_, new_n10610_, new_n10611_,
    new_n10612_, new_n10613_, new_n10614_, new_n10616_, new_n10617_,
    new_n10618_, new_n10619_, new_n10620_, new_n10621_, new_n10622_,
    new_n10623_, new_n10624_, new_n10625_, new_n10626_, new_n10627_,
    new_n10628_, new_n10629_, new_n10630_, new_n10631_, new_n10632_,
    new_n10633_, new_n10634_, new_n10635_, new_n10636_, new_n10637_,
    new_n10638_, new_n10639_, new_n10640_, new_n10641_, new_n10642_,
    new_n10643_, new_n10644_, new_n10645_, new_n10646_, new_n10647_,
    new_n10648_, new_n10649_, new_n10650_, new_n10651_, new_n10652_,
    new_n10653_, new_n10654_, new_n10655_, new_n10656_, new_n10657_,
    new_n10658_, new_n10659_, new_n10660_, new_n10661_, new_n10662_,
    new_n10663_, new_n10664_, new_n10665_, new_n10666_, new_n10667_,
    new_n10668_, new_n10669_, new_n10670_, new_n10671_, new_n10672_,
    new_n10673_, new_n10674_, new_n10675_, new_n10676_, new_n10677_,
    new_n10678_, new_n10679_, new_n10680_, new_n10681_, new_n10682_,
    new_n10683_, new_n10684_, new_n10685_, new_n10686_, new_n10687_,
    new_n10688_, new_n10689_, new_n10690_, new_n10691_, new_n10692_,
    new_n10693_, new_n10694_, new_n10695_, new_n10696_, new_n10697_,
    new_n10698_, new_n10699_, new_n10700_, new_n10701_, new_n10702_,
    new_n10703_, new_n10704_, new_n10705_, new_n10706_, new_n10707_,
    new_n10708_, new_n10709_, new_n10710_, new_n10711_, new_n10712_,
    new_n10713_, new_n10714_, new_n10715_, new_n10716_, new_n10717_,
    new_n10718_, new_n10719_, new_n10720_, new_n10721_, new_n10722_,
    new_n10723_, new_n10724_, new_n10725_, new_n10726_, new_n10727_,
    new_n10728_, new_n10729_, new_n10730_, new_n10731_, new_n10732_,
    new_n10733_, new_n10734_, new_n10735_, new_n10736_, new_n10737_,
    new_n10738_, new_n10739_, new_n10740_, new_n10741_, new_n10742_,
    new_n10743_, new_n10744_, new_n10745_, new_n10746_, new_n10747_,
    new_n10748_, new_n10749_, new_n10750_, new_n10751_, new_n10752_,
    new_n10753_, new_n10754_, new_n10755_, new_n10756_, new_n10757_,
    new_n10758_, new_n10759_, new_n10760_, new_n10761_, new_n10762_,
    new_n10763_, new_n10764_, new_n10765_, new_n10766_, new_n10767_,
    new_n10768_, new_n10769_, new_n10770_, new_n10771_, new_n10772_,
    new_n10773_, new_n10774_, new_n10775_, new_n10776_, new_n10777_,
    new_n10778_, new_n10779_, new_n10780_, new_n10781_, new_n10782_,
    new_n10783_, new_n10784_, new_n10785_, new_n10786_, new_n10787_,
    new_n10788_, new_n10789_, new_n10790_, new_n10791_, new_n10792_,
    new_n10793_, new_n10794_, new_n10795_, new_n10796_, new_n10797_,
    new_n10798_, new_n10799_, new_n10800_, new_n10801_, new_n10802_,
    new_n10803_, new_n10804_, new_n10805_, new_n10806_, new_n10807_,
    new_n10808_, new_n10809_, new_n10810_, new_n10811_, new_n10812_,
    new_n10813_, new_n10814_, new_n10815_, new_n10816_, new_n10817_,
    new_n10818_, new_n10819_, new_n10820_, new_n10821_, new_n10822_,
    new_n10823_, new_n10824_, new_n10825_, new_n10826_, new_n10827_,
    new_n10828_, new_n10829_, new_n10830_, new_n10831_, new_n10832_,
    new_n10833_, new_n10834_, new_n10835_, new_n10836_, new_n10837_,
    new_n10838_, new_n10839_, new_n10840_, new_n10841_, new_n10842_,
    new_n10843_, new_n10844_, new_n10845_, new_n10846_, new_n10847_,
    new_n10848_, new_n10849_, new_n10850_, new_n10851_, new_n10852_,
    new_n10853_, new_n10854_, new_n10855_, new_n10856_, new_n10857_,
    new_n10858_, new_n10859_, new_n10860_, new_n10861_, new_n10862_,
    new_n10863_, new_n10864_, new_n10865_, new_n10866_, new_n10867_,
    new_n10868_, new_n10869_, new_n10870_, new_n10871_, new_n10872_,
    new_n10873_, new_n10874_, new_n10875_, new_n10876_, new_n10877_,
    new_n10878_, new_n10879_, new_n10880_, new_n10881_, new_n10882_,
    new_n10883_, new_n10884_, new_n10885_, new_n10886_, new_n10887_,
    new_n10888_, new_n10889_, new_n10890_, new_n10891_, new_n10892_,
    new_n10893_, new_n10894_, new_n10895_, new_n10896_, new_n10897_,
    new_n10898_, new_n10899_, new_n10900_, new_n10901_, new_n10902_,
    new_n10903_, new_n10904_, new_n10905_, new_n10906_, new_n10907_,
    new_n10909_, new_n10910_, new_n10911_, new_n10912_, new_n10913_,
    new_n10914_, new_n10915_, new_n10916_, new_n10917_, new_n10918_,
    new_n10919_, new_n10920_, new_n10921_, new_n10922_, new_n10923_,
    new_n10924_, new_n10925_, new_n10926_, new_n10927_, new_n10928_,
    new_n10929_, new_n10930_, new_n10931_, new_n10932_, new_n10933_,
    new_n10934_, new_n10935_, new_n10936_, new_n10937_, new_n10938_,
    new_n10939_, new_n10940_, new_n10941_, new_n10942_, new_n10943_,
    new_n10944_, new_n10945_, new_n10946_, new_n10947_, new_n10948_,
    new_n10949_, new_n10950_, new_n10951_, new_n10952_, new_n10953_,
    new_n10954_, new_n10955_, new_n10956_, new_n10957_, new_n10958_,
    new_n10959_, new_n10960_, new_n10961_, new_n10962_, new_n10963_,
    new_n10964_, new_n10965_, new_n10966_, new_n10967_, new_n10968_,
    new_n10969_, new_n10970_, new_n10971_, new_n10972_, new_n10973_,
    new_n10974_, new_n10975_, new_n10976_, new_n10977_, new_n10978_,
    new_n10979_, new_n10980_, new_n10981_, new_n10982_, new_n10983_,
    new_n10984_, new_n10985_, new_n10986_, new_n10987_, new_n10988_,
    new_n10989_, new_n10990_, new_n10991_, new_n10992_, new_n10993_,
    new_n10994_, new_n10995_, new_n10996_, new_n10997_, new_n10998_,
    new_n10999_, new_n11000_, new_n11001_, new_n11002_, new_n11003_,
    new_n11004_, new_n11005_, new_n11006_, new_n11007_, new_n11008_,
    new_n11009_, new_n11010_, new_n11011_, new_n11012_, new_n11013_,
    new_n11014_, new_n11015_, new_n11016_, new_n11017_, new_n11018_,
    new_n11019_, new_n11020_, new_n11021_, new_n11022_, new_n11023_,
    new_n11024_, new_n11025_, new_n11026_, new_n11027_, new_n11028_,
    new_n11029_, new_n11030_, new_n11031_, new_n11032_, new_n11033_,
    new_n11034_, new_n11035_, new_n11036_, new_n11037_, new_n11038_,
    new_n11039_, new_n11040_, new_n11041_, new_n11042_, new_n11043_,
    new_n11044_, new_n11045_, new_n11046_, new_n11047_, new_n11048_,
    new_n11049_, new_n11050_, new_n11051_, new_n11052_, new_n11053_,
    new_n11054_, new_n11055_, new_n11056_, new_n11057_, new_n11058_,
    new_n11059_, new_n11060_, new_n11061_, new_n11062_, new_n11063_,
    new_n11064_, new_n11065_, new_n11066_, new_n11067_, new_n11068_,
    new_n11069_, new_n11070_, new_n11071_, new_n11072_, new_n11073_,
    new_n11074_, new_n11075_, new_n11076_, new_n11077_, new_n11078_,
    new_n11079_, new_n11080_, new_n11081_, new_n11082_, new_n11083_,
    new_n11084_, new_n11085_, new_n11086_, new_n11087_, new_n11088_,
    new_n11089_, new_n11090_, new_n11091_, new_n11092_, new_n11093_,
    new_n11094_, new_n11095_, new_n11096_, new_n11097_, new_n11098_,
    new_n11099_, new_n11100_, new_n11101_, new_n11102_, new_n11103_,
    new_n11104_, new_n11105_, new_n11106_, new_n11107_, new_n11108_,
    new_n11109_, new_n11110_, new_n11111_, new_n11112_, new_n11113_,
    new_n11114_, new_n11115_, new_n11116_, new_n11117_, new_n11118_,
    new_n11119_, new_n11120_, new_n11121_, new_n11122_, new_n11123_,
    new_n11124_, new_n11125_, new_n11126_, new_n11127_, new_n11128_,
    new_n11129_, new_n11130_, new_n11131_, new_n11132_, new_n11133_,
    new_n11134_, new_n11135_, new_n11136_, new_n11137_, new_n11138_,
    new_n11139_, new_n11140_, new_n11141_, new_n11142_, new_n11143_,
    new_n11144_, new_n11145_, new_n11146_, new_n11147_, new_n11148_,
    new_n11149_, new_n11150_, new_n11151_, new_n11152_, new_n11153_,
    new_n11154_, new_n11155_, new_n11156_, new_n11157_, new_n11158_,
    new_n11159_, new_n11160_, new_n11161_, new_n11162_, new_n11163_,
    new_n11164_, new_n11165_, new_n11166_, new_n11167_, new_n11168_,
    new_n11169_, new_n11170_, new_n11171_, new_n11172_, new_n11173_,
    new_n11174_, new_n11175_, new_n11176_, new_n11177_, new_n11178_,
    new_n11179_, new_n11180_, new_n11181_, new_n11182_, new_n11183_,
    new_n11184_, new_n11185_, new_n11186_, new_n11187_, new_n11188_,
    new_n11189_, new_n11190_, new_n11191_, new_n11192_, new_n11193_,
    new_n11194_, new_n11195_, new_n11196_, new_n11197_, new_n11198_,
    new_n11199_, new_n11200_, new_n11201_, new_n11202_, new_n11203_,
    new_n11204_, new_n11205_, new_n11206_, new_n11207_, new_n11208_,
    new_n11209_, new_n11210_, new_n11211_, new_n11212_, new_n11213_,
    new_n11214_, new_n11215_, new_n11216_, new_n11217_, new_n11218_,
    new_n11219_, new_n11220_, new_n11221_, new_n11223_, new_n11224_,
    new_n11225_, new_n11226_, new_n11227_, new_n11228_, new_n11229_,
    new_n11230_, new_n11231_, new_n11232_, new_n11233_, new_n11234_,
    new_n11235_, new_n11236_, new_n11237_, new_n11238_, new_n11239_,
    new_n11240_, new_n11241_, new_n11242_, new_n11243_, new_n11244_,
    new_n11245_, new_n11246_, new_n11247_, new_n11248_, new_n11249_,
    new_n11250_, new_n11251_, new_n11252_, new_n11253_, new_n11254_,
    new_n11255_, new_n11256_, new_n11257_, new_n11258_, new_n11259_,
    new_n11260_, new_n11261_, new_n11262_, new_n11263_, new_n11264_,
    new_n11265_, new_n11266_, new_n11267_, new_n11268_, new_n11269_,
    new_n11270_, new_n11271_, new_n11272_, new_n11273_, new_n11274_,
    new_n11275_, new_n11276_, new_n11277_, new_n11278_, new_n11279_,
    new_n11280_, new_n11281_, new_n11282_, new_n11283_, new_n11284_,
    new_n11285_, new_n11286_, new_n11287_, new_n11288_, new_n11289_,
    new_n11290_, new_n11291_, new_n11292_, new_n11293_, new_n11294_,
    new_n11295_, new_n11296_, new_n11297_, new_n11298_, new_n11299_,
    new_n11300_, new_n11301_, new_n11302_, new_n11303_, new_n11304_,
    new_n11305_, new_n11306_, new_n11307_, new_n11308_, new_n11309_,
    new_n11310_, new_n11311_, new_n11312_, new_n11313_, new_n11314_,
    new_n11315_, new_n11316_, new_n11317_, new_n11318_, new_n11319_,
    new_n11320_, new_n11321_, new_n11322_, new_n11323_, new_n11324_,
    new_n11325_, new_n11326_, new_n11327_, new_n11328_, new_n11329_,
    new_n11330_, new_n11331_, new_n11332_, new_n11333_, new_n11334_,
    new_n11335_, new_n11336_, new_n11337_, new_n11338_, new_n11339_,
    new_n11340_, new_n11341_, new_n11342_, new_n11343_, new_n11344_,
    new_n11345_, new_n11346_, new_n11347_, new_n11348_, new_n11349_,
    new_n11350_, new_n11351_, new_n11352_, new_n11353_, new_n11354_,
    new_n11355_, new_n11356_, new_n11357_, new_n11358_, new_n11359_,
    new_n11360_, new_n11361_, new_n11362_, new_n11363_, new_n11364_,
    new_n11365_, new_n11366_, new_n11367_, new_n11368_, new_n11369_,
    new_n11370_, new_n11371_, new_n11372_, new_n11373_, new_n11374_,
    new_n11375_, new_n11376_, new_n11377_, new_n11378_, new_n11379_,
    new_n11380_, new_n11381_, new_n11382_, new_n11383_, new_n11384_,
    new_n11385_, new_n11386_, new_n11387_, new_n11388_, new_n11389_,
    new_n11390_, new_n11391_, new_n11392_, new_n11393_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11399_,
    new_n11400_, new_n11401_, new_n11402_, new_n11403_, new_n11404_,
    new_n11405_, new_n11406_, new_n11407_, new_n11408_, new_n11409_,
    new_n11410_, new_n11411_, new_n11412_, new_n11413_, new_n11414_,
    new_n11415_, new_n11416_, new_n11417_, new_n11418_, new_n11419_,
    new_n11420_, new_n11421_, new_n11422_, new_n11423_, new_n11424_,
    new_n11425_, new_n11426_, new_n11427_, new_n11428_, new_n11429_,
    new_n11430_, new_n11431_, new_n11432_, new_n11433_, new_n11434_,
    new_n11435_, new_n11436_, new_n11437_, new_n11438_, new_n11439_,
    new_n11440_, new_n11441_, new_n11442_, new_n11443_, new_n11444_,
    new_n11445_, new_n11446_, new_n11447_, new_n11448_, new_n11449_,
    new_n11450_, new_n11451_, new_n11452_, new_n11453_, new_n11454_,
    new_n11455_, new_n11456_, new_n11457_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11496_, new_n11497_, new_n11498_, new_n11499_,
    new_n11500_, new_n11501_, new_n11502_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11507_, new_n11508_, new_n11509_,
    new_n11510_, new_n11511_, new_n11512_, new_n11513_, new_n11514_,
    new_n11515_, new_n11516_, new_n11517_, new_n11518_, new_n11519_,
    new_n11520_, new_n11521_, new_n11522_, new_n11523_, new_n11524_,
    new_n11525_, new_n11526_, new_n11527_, new_n11528_, new_n11529_,
    new_n11530_, new_n11531_, new_n11532_, new_n11533_, new_n11534_,
    new_n11535_, new_n11536_, new_n11537_, new_n11538_, new_n11539_,
    new_n11540_, new_n11541_, new_n11542_, new_n11543_, new_n11544_,
    new_n11545_, new_n11546_, new_n11547_, new_n11548_, new_n11549_,
    new_n11550_, new_n11551_, new_n11552_, new_n11553_, new_n11554_,
    new_n11555_, new_n11556_, new_n11557_, new_n11558_, new_n11559_,
    new_n11560_, new_n11561_, new_n11562_, new_n11563_, new_n11564_,
    new_n11565_, new_n11566_, new_n11567_, new_n11568_, new_n11569_,
    new_n11570_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11622_, new_n11623_, new_n11624_, new_n11625_,
    new_n11626_, new_n11627_, new_n11628_, new_n11629_, new_n11630_,
    new_n11631_, new_n11632_, new_n11633_, new_n11634_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11654_, new_n11655_,
    new_n11656_, new_n11657_, new_n11658_, new_n11659_, new_n11660_,
    new_n11661_, new_n11662_, new_n11663_, new_n11664_, new_n11665_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11693_, new_n11694_, new_n11695_,
    new_n11696_, new_n11697_, new_n11698_, new_n11699_, new_n11700_,
    new_n11701_, new_n11702_, new_n11703_, new_n11704_, new_n11705_,
    new_n11706_, new_n11707_, new_n11708_, new_n11709_, new_n11710_,
    new_n11711_, new_n11712_, new_n11713_, new_n11714_, new_n11715_,
    new_n11716_, new_n11717_, new_n11718_, new_n11719_, new_n11720_,
    new_n11721_, new_n11722_, new_n11723_, new_n11724_, new_n11725_,
    new_n11726_, new_n11727_, new_n11728_, new_n11729_, new_n11730_,
    new_n11731_, new_n11732_, new_n11733_, new_n11734_, new_n11735_,
    new_n11736_, new_n11737_, new_n11738_, new_n11739_, new_n11740_,
    new_n11741_, new_n11742_, new_n11743_, new_n11744_, new_n11745_,
    new_n11746_, new_n11747_, new_n11748_, new_n11749_, new_n11750_,
    new_n11751_, new_n11752_, new_n11753_, new_n11754_, new_n11755_,
    new_n11756_, new_n11757_, new_n11758_, new_n11759_, new_n11760_,
    new_n11761_, new_n11762_, new_n11763_, new_n11764_, new_n11765_,
    new_n11766_, new_n11767_, new_n11768_, new_n11769_, new_n11770_,
    new_n11771_, new_n11772_, new_n11773_, new_n11774_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11780_,
    new_n11781_, new_n11782_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11804_, new_n11805_,
    new_n11806_, new_n11807_, new_n11808_, new_n11809_, new_n11810_,
    new_n11811_, new_n11812_, new_n11813_, new_n11814_, new_n11815_,
    new_n11816_, new_n11817_, new_n11818_, new_n11819_, new_n11820_,
    new_n11821_, new_n11822_, new_n11823_, new_n11824_, new_n11825_,
    new_n11826_, new_n11827_, new_n11828_, new_n11829_, new_n11830_,
    new_n11831_, new_n11832_, new_n11833_, new_n11834_, new_n11835_,
    new_n11836_, new_n11837_, new_n11838_, new_n11839_, new_n11840_,
    new_n11841_, new_n11842_, new_n11843_, new_n11844_, new_n11845_,
    new_n11846_, new_n11847_, new_n11848_, new_n11849_, new_n11850_,
    new_n11851_, new_n11852_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11858_, new_n11859_, new_n11860_,
    new_n11861_, new_n11862_, new_n11863_, new_n11864_, new_n11865_,
    new_n11866_, new_n11867_, new_n11868_, new_n11869_, new_n11870_,
    new_n11871_, new_n11873_, new_n11874_, new_n11875_, new_n11876_,
    new_n11877_, new_n11878_, new_n11879_, new_n11880_, new_n11881_,
    new_n11882_, new_n11883_, new_n11884_, new_n11885_, new_n11886_,
    new_n11887_, new_n11888_, new_n11889_, new_n11890_, new_n11891_,
    new_n11892_, new_n11893_, new_n11894_, new_n11895_, new_n11896_,
    new_n11897_, new_n11898_, new_n11899_, new_n11900_, new_n11901_,
    new_n11902_, new_n11903_, new_n11904_, new_n11905_, new_n11906_,
    new_n11907_, new_n11908_, new_n11909_, new_n11910_, new_n11911_,
    new_n11912_, new_n11913_, new_n11914_, new_n11915_, new_n11916_,
    new_n11917_, new_n11918_, new_n11919_, new_n11920_, new_n11921_,
    new_n11922_, new_n11923_, new_n11924_, new_n11925_, new_n11926_,
    new_n11927_, new_n11928_, new_n11929_, new_n11930_, new_n11931_,
    new_n11932_, new_n11933_, new_n11934_, new_n11935_, new_n11936_,
    new_n11937_, new_n11938_, new_n11939_, new_n11940_, new_n11941_,
    new_n11942_, new_n11943_, new_n11944_, new_n11945_, new_n11946_,
    new_n11947_, new_n11948_, new_n11949_, new_n11950_, new_n11951_,
    new_n11952_, new_n11953_, new_n11954_, new_n11955_, new_n11956_,
    new_n11957_, new_n11958_, new_n11959_, new_n11960_, new_n11961_,
    new_n11962_, new_n11963_, new_n11964_, new_n11965_, new_n11966_,
    new_n11967_, new_n11968_, new_n11969_, new_n11970_, new_n11971_,
    new_n11972_, new_n11973_, new_n11974_, new_n11975_, new_n11976_,
    new_n11977_, new_n11978_, new_n11979_, new_n11980_, new_n11981_,
    new_n11982_, new_n11983_, new_n11984_, new_n11985_, new_n11986_,
    new_n11987_, new_n11988_, new_n11989_, new_n11990_, new_n11991_,
    new_n11992_, new_n11993_, new_n11994_, new_n11995_, new_n11996_,
    new_n11997_, new_n11998_, new_n11999_, new_n12000_, new_n12001_,
    new_n12002_, new_n12003_, new_n12004_, new_n12005_, new_n12006_,
    new_n12007_, new_n12008_, new_n12009_, new_n12010_, new_n12011_,
    new_n12012_, new_n12013_, new_n12014_, new_n12015_, new_n12016_,
    new_n12017_, new_n12018_, new_n12019_, new_n12020_, new_n12021_,
    new_n12022_, new_n12023_, new_n12024_, new_n12025_, new_n12026_,
    new_n12027_, new_n12028_, new_n12029_, new_n12030_, new_n12031_,
    new_n12032_, new_n12033_, new_n12034_, new_n12035_, new_n12036_,
    new_n12037_, new_n12038_, new_n12039_, new_n12040_, new_n12041_,
    new_n12042_, new_n12043_, new_n12044_, new_n12045_, new_n12046_,
    new_n12047_, new_n12048_, new_n12049_, new_n12050_, new_n12051_,
    new_n12052_, new_n12053_, new_n12054_, new_n12055_, new_n12056_,
    new_n12057_, new_n12058_, new_n12059_, new_n12060_, new_n12061_,
    new_n12062_, new_n12063_, new_n12064_, new_n12065_, new_n12066_,
    new_n12067_, new_n12068_, new_n12069_, new_n12070_, new_n12071_,
    new_n12072_, new_n12073_, new_n12074_, new_n12075_, new_n12076_,
    new_n12077_, new_n12078_, new_n12079_, new_n12080_, new_n12081_,
    new_n12082_, new_n12083_, new_n12084_, new_n12085_, new_n12086_,
    new_n12087_, new_n12088_, new_n12089_, new_n12090_, new_n12091_,
    new_n12092_, new_n12093_, new_n12094_, new_n12095_, new_n12096_,
    new_n12097_, new_n12098_, new_n12099_, new_n12100_, new_n12101_,
    new_n12102_, new_n12103_, new_n12104_, new_n12105_, new_n12106_,
    new_n12107_, new_n12108_, new_n12109_, new_n12110_, new_n12111_,
    new_n12112_, new_n12113_, new_n12114_, new_n12115_, new_n12116_,
    new_n12117_, new_n12118_, new_n12119_, new_n12120_, new_n12121_,
    new_n12122_, new_n12123_, new_n12124_, new_n12125_, new_n12126_,
    new_n12127_, new_n12128_, new_n12129_, new_n12130_, new_n12131_,
    new_n12132_, new_n12133_, new_n12134_, new_n12135_, new_n12136_,
    new_n12137_, new_n12138_, new_n12139_, new_n12140_, new_n12141_,
    new_n12142_, new_n12143_, new_n12144_, new_n12145_, new_n12146_,
    new_n12147_, new_n12148_, new_n12149_, new_n12150_, new_n12151_,
    new_n12152_, new_n12153_, new_n12154_, new_n12155_, new_n12156_,
    new_n12157_, new_n12158_, new_n12159_, new_n12160_, new_n12161_,
    new_n12162_, new_n12163_, new_n12164_, new_n12165_, new_n12166_,
    new_n12167_, new_n12168_, new_n12169_, new_n12170_, new_n12171_,
    new_n12172_, new_n12173_, new_n12174_, new_n12175_, new_n12176_,
    new_n12177_, new_n12178_, new_n12179_, new_n12180_, new_n12181_,
    new_n12182_, new_n12183_, new_n12184_, new_n12185_, new_n12186_,
    new_n12187_, new_n12188_, new_n12189_, new_n12190_, new_n12192_,
    new_n12193_, new_n12194_, new_n12195_, new_n12196_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12203_, new_n12204_, new_n12205_, new_n12206_, new_n12207_,
    new_n12208_, new_n12209_, new_n12210_, new_n12211_, new_n12212_,
    new_n12213_, new_n12214_, new_n12215_, new_n12216_, new_n12217_,
    new_n12218_, new_n12219_, new_n12220_, new_n12221_, new_n12222_,
    new_n12223_, new_n12224_, new_n12225_, new_n12226_, new_n12227_,
    new_n12228_, new_n12229_, new_n12230_, new_n12231_, new_n12232_,
    new_n12233_, new_n12234_, new_n12235_, new_n12236_, new_n12237_,
    new_n12238_, new_n12239_, new_n12240_, new_n12241_, new_n12242_,
    new_n12243_, new_n12244_, new_n12245_, new_n12246_, new_n12247_,
    new_n12248_, new_n12249_, new_n12250_, new_n12251_, new_n12252_,
    new_n12253_, new_n12254_, new_n12255_, new_n12256_, new_n12257_,
    new_n12258_, new_n12259_, new_n12260_, new_n12261_, new_n12262_,
    new_n12263_, new_n12264_, new_n12265_, new_n12266_, new_n12267_,
    new_n12268_, new_n12269_, new_n12270_, new_n12271_, new_n12272_,
    new_n12273_, new_n12274_, new_n12275_, new_n12276_, new_n12277_,
    new_n12278_, new_n12279_, new_n12280_, new_n12281_, new_n12282_,
    new_n12283_, new_n12284_, new_n12285_, new_n12286_, new_n12287_,
    new_n12288_, new_n12289_, new_n12290_, new_n12291_, new_n12292_,
    new_n12293_, new_n12294_, new_n12295_, new_n12296_, new_n12297_,
    new_n12298_, new_n12299_, new_n12300_, new_n12301_, new_n12302_,
    new_n12303_, new_n12304_, new_n12305_, new_n12306_, new_n12307_,
    new_n12308_, new_n12309_, new_n12310_, new_n12311_, new_n12312_,
    new_n12313_, new_n12314_, new_n12315_, new_n12316_, new_n12317_,
    new_n12318_, new_n12319_, new_n12320_, new_n12321_, new_n12322_,
    new_n12323_, new_n12324_, new_n12325_, new_n12326_, new_n12327_,
    new_n12328_, new_n12329_, new_n12330_, new_n12331_, new_n12332_,
    new_n12333_, new_n12334_, new_n12335_, new_n12336_, new_n12337_,
    new_n12338_, new_n12339_, new_n12340_, new_n12341_, new_n12342_,
    new_n12343_, new_n12344_, new_n12345_, new_n12346_, new_n12347_,
    new_n12348_, new_n12349_, new_n12350_, new_n12351_, new_n12352_,
    new_n12353_, new_n12354_, new_n12355_, new_n12356_, new_n12357_,
    new_n12358_, new_n12359_, new_n12360_, new_n12361_, new_n12362_,
    new_n12363_, new_n12364_, new_n12365_, new_n12366_, new_n12367_,
    new_n12368_, new_n12369_, new_n12370_, new_n12371_, new_n12372_,
    new_n12373_, new_n12374_, new_n12375_, new_n12376_, new_n12377_,
    new_n12378_, new_n12379_, new_n12380_, new_n12381_, new_n12382_,
    new_n12383_, new_n12384_, new_n12385_, new_n12386_, new_n12387_,
    new_n12388_, new_n12389_, new_n12390_, new_n12391_, new_n12392_,
    new_n12393_, new_n12394_, new_n12395_, new_n12396_, new_n12397_,
    new_n12398_, new_n12399_, new_n12400_, new_n12401_, new_n12402_,
    new_n12403_, new_n12404_, new_n12405_, new_n12406_, new_n12407_,
    new_n12408_, new_n12409_, new_n12410_, new_n12411_, new_n12412_,
    new_n12413_, new_n12414_, new_n12415_, new_n12416_, new_n12417_,
    new_n12418_, new_n12419_, new_n12420_, new_n12421_, new_n12422_,
    new_n12423_, new_n12424_, new_n12425_, new_n12426_, new_n12427_,
    new_n12428_, new_n12429_, new_n12430_, new_n12431_, new_n12432_,
    new_n12433_, new_n12434_, new_n12435_, new_n12436_, new_n12437_,
    new_n12438_, new_n12439_, new_n12440_, new_n12441_, new_n12442_,
    new_n12443_, new_n12444_, new_n12445_, new_n12446_, new_n12447_,
    new_n12448_, new_n12449_, new_n12450_, new_n12451_, new_n12452_,
    new_n12453_, new_n12454_, new_n12455_, new_n12456_, new_n12457_,
    new_n12458_, new_n12459_, new_n12460_, new_n12461_, new_n12462_,
    new_n12463_, new_n12464_, new_n12465_, new_n12466_, new_n12467_,
    new_n12468_, new_n12469_, new_n12470_, new_n12471_, new_n12472_,
    new_n12473_, new_n12474_, new_n12475_, new_n12476_, new_n12477_,
    new_n12478_, new_n12479_, new_n12480_, new_n12481_, new_n12482_,
    new_n12483_, new_n12484_, new_n12485_, new_n12486_, new_n12487_,
    new_n12488_, new_n12489_, new_n12490_, new_n12491_, new_n12492_,
    new_n12493_, new_n12494_, new_n12495_, new_n12496_, new_n12497_,
    new_n12498_, new_n12499_, new_n12500_, new_n12501_, new_n12502_,
    new_n12503_, new_n12504_, new_n12505_, new_n12506_, new_n12507_,
    new_n12508_, new_n12509_, new_n12510_, new_n12511_, new_n12512_,
    new_n12513_, new_n12514_, new_n12515_, new_n12516_, new_n12517_,
    new_n12518_, new_n12519_, new_n12520_, new_n12521_, new_n12522_,
    new_n12523_, new_n12524_, new_n12525_, new_n12526_, new_n12527_,
    new_n12528_, new_n12529_, new_n12530_, new_n12531_, new_n12532_,
    new_n12533_, new_n12534_, new_n12535_, new_n12536_, new_n12537_,
    new_n12538_, new_n12539_, new_n12541_, new_n12542_, new_n12543_,
    new_n12544_, new_n12545_, new_n12546_, new_n12547_, new_n12548_,
    new_n12549_, new_n12550_, new_n12551_, new_n12552_, new_n12553_,
    new_n12554_, new_n12555_, new_n12556_, new_n12557_, new_n12558_,
    new_n12559_, new_n12560_, new_n12561_, new_n12562_, new_n12563_,
    new_n12564_, new_n12565_, new_n12566_, new_n12567_, new_n12568_,
    new_n12569_, new_n12570_, new_n12571_, new_n12572_, new_n12573_,
    new_n12574_, new_n12575_, new_n12576_, new_n12577_, new_n12578_,
    new_n12579_, new_n12580_, new_n12581_, new_n12582_, new_n12583_,
    new_n12584_, new_n12585_, new_n12586_, new_n12587_, new_n12588_,
    new_n12589_, new_n12590_, new_n12591_, new_n12592_, new_n12593_,
    new_n12594_, new_n12595_, new_n12596_, new_n12597_, new_n12598_,
    new_n12599_, new_n12600_, new_n12601_, new_n12602_, new_n12603_,
    new_n12604_, new_n12605_, new_n12606_, new_n12607_, new_n12608_,
    new_n12609_, new_n12610_, new_n12611_, new_n12612_, new_n12613_,
    new_n12614_, new_n12615_, new_n12616_, new_n12617_, new_n12618_,
    new_n12619_, new_n12620_, new_n12621_, new_n12622_, new_n12623_,
    new_n12624_, new_n12625_, new_n12626_, new_n12627_, new_n12628_,
    new_n12629_, new_n12630_, new_n12631_, new_n12632_, new_n12633_,
    new_n12634_, new_n12635_, new_n12636_, new_n12637_, new_n12638_,
    new_n12639_, new_n12640_, new_n12641_, new_n12642_, new_n12643_,
    new_n12644_, new_n12645_, new_n12646_, new_n12647_, new_n12648_,
    new_n12649_, new_n12650_, new_n12651_, new_n12652_, new_n12653_,
    new_n12654_, new_n12655_, new_n12656_, new_n12657_, new_n12658_,
    new_n12659_, new_n12660_, new_n12661_, new_n12662_, new_n12663_,
    new_n12664_, new_n12665_, new_n12666_, new_n12667_, new_n12668_,
    new_n12669_, new_n12670_, new_n12671_, new_n12672_, new_n12673_,
    new_n12674_, new_n12675_, new_n12676_, new_n12677_, new_n12678_,
    new_n12679_, new_n12680_, new_n12681_, new_n12682_, new_n12683_,
    new_n12684_, new_n12685_, new_n12686_, new_n12687_, new_n12688_,
    new_n12689_, new_n12690_, new_n12691_, new_n12692_, new_n12693_,
    new_n12694_, new_n12695_, new_n12696_, new_n12697_, new_n12698_,
    new_n12699_, new_n12700_, new_n12701_, new_n12702_, new_n12703_,
    new_n12704_, new_n12705_, new_n12706_, new_n12707_, new_n12708_,
    new_n12709_, new_n12710_, new_n12711_, new_n12712_, new_n12713_,
    new_n12714_, new_n12715_, new_n12716_, new_n12717_, new_n12718_,
    new_n12719_, new_n12720_, new_n12721_, new_n12722_, new_n12723_,
    new_n12724_, new_n12725_, new_n12726_, new_n12727_, new_n12728_,
    new_n12729_, new_n12730_, new_n12731_, new_n12732_, new_n12733_,
    new_n12734_, new_n12735_, new_n12736_, new_n12737_, new_n12738_,
    new_n12739_, new_n12740_, new_n12741_, new_n12742_, new_n12743_,
    new_n12744_, new_n12745_, new_n12746_, new_n12747_, new_n12748_,
    new_n12749_, new_n12750_, new_n12751_, new_n12752_, new_n12753_,
    new_n12754_, new_n12755_, new_n12756_, new_n12757_, new_n12758_,
    new_n12759_, new_n12760_, new_n12761_, new_n12762_, new_n12763_,
    new_n12764_, new_n12765_, new_n12766_, new_n12767_, new_n12768_,
    new_n12769_, new_n12770_, new_n12771_, new_n12772_, new_n12773_,
    new_n12774_, new_n12775_, new_n12776_, new_n12777_, new_n12778_,
    new_n12779_, new_n12780_, new_n12781_, new_n12782_, new_n12783_,
    new_n12784_, new_n12785_, new_n12786_, new_n12787_, new_n12788_,
    new_n12789_, new_n12790_, new_n12791_, new_n12792_, new_n12793_,
    new_n12794_, new_n12795_, new_n12796_, new_n12797_, new_n12798_,
    new_n12799_, new_n12800_, new_n12801_, new_n12802_, new_n12803_,
    new_n12804_, new_n12805_, new_n12806_, new_n12807_, new_n12808_,
    new_n12809_, new_n12810_, new_n12811_, new_n12812_, new_n12813_,
    new_n12814_, new_n12815_, new_n12816_, new_n12817_, new_n12818_,
    new_n12819_, new_n12820_, new_n12821_, new_n12822_, new_n12823_,
    new_n12824_, new_n12825_, new_n12826_, new_n12827_, new_n12828_,
    new_n12829_, new_n12830_, new_n12831_, new_n12832_, new_n12833_,
    new_n12834_, new_n12835_, new_n12836_, new_n12837_, new_n12838_,
    new_n12839_, new_n12841_, new_n12842_, new_n12843_, new_n12844_,
    new_n12845_, new_n12846_, new_n12847_, new_n12848_, new_n12849_,
    new_n12850_, new_n12851_, new_n12852_, new_n12853_, new_n12854_,
    new_n12855_, new_n12856_, new_n12857_, new_n12858_, new_n12859_,
    new_n12860_, new_n12861_, new_n12862_, new_n12863_, new_n12864_,
    new_n12865_, new_n12866_, new_n12867_, new_n12868_, new_n12869_,
    new_n12870_, new_n12871_, new_n12872_, new_n12873_, new_n12874_,
    new_n12875_, new_n12876_, new_n12877_, new_n12878_, new_n12879_,
    new_n12880_, new_n12881_, new_n12882_, new_n12883_, new_n12884_,
    new_n12885_, new_n12886_, new_n12887_, new_n12888_, new_n12889_,
    new_n12890_, new_n12891_, new_n12892_, new_n12893_, new_n12894_,
    new_n12895_, new_n12896_, new_n12897_, new_n12898_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13006_, new_n13007_, new_n13008_, new_n13009_,
    new_n13010_, new_n13011_, new_n13012_, new_n13013_, new_n13014_,
    new_n13015_, new_n13016_, new_n13017_, new_n13018_, new_n13019_,
    new_n13020_, new_n13021_, new_n13022_, new_n13023_, new_n13024_,
    new_n13025_, new_n13026_, new_n13027_, new_n13028_, new_n13029_,
    new_n13030_, new_n13031_, new_n13032_, new_n13033_, new_n13034_,
    new_n13035_, new_n13036_, new_n13037_, new_n13038_, new_n13039_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13046_, new_n13047_, new_n13048_, new_n13049_,
    new_n13050_, new_n13051_, new_n13052_, new_n13053_, new_n13054_,
    new_n13055_, new_n13056_, new_n13057_, new_n13058_, new_n13059_,
    new_n13060_, new_n13061_, new_n13062_, new_n13063_, new_n13064_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13069_,
    new_n13070_, new_n13071_, new_n13072_, new_n13073_, new_n13074_,
    new_n13075_, new_n13076_, new_n13077_, new_n13078_, new_n13079_,
    new_n13080_, new_n13081_, new_n13082_, new_n13083_, new_n13084_,
    new_n13085_, new_n13086_, new_n13087_, new_n13088_, new_n13089_,
    new_n13090_, new_n13091_, new_n13092_, new_n13093_, new_n13094_,
    new_n13095_, new_n13096_, new_n13097_, new_n13098_, new_n13099_,
    new_n13100_, new_n13101_, new_n13102_, new_n13103_, new_n13104_,
    new_n13105_, new_n13106_, new_n13107_, new_n13108_, new_n13109_,
    new_n13110_, new_n13111_, new_n13112_, new_n13113_, new_n13114_,
    new_n13115_, new_n13116_, new_n13117_, new_n13118_, new_n13119_,
    new_n13120_, new_n13121_, new_n13122_, new_n13123_, new_n13124_,
    new_n13125_, new_n13126_, new_n13127_, new_n13128_, new_n13129_,
    new_n13130_, new_n13131_, new_n13132_, new_n13133_, new_n13134_,
    new_n13135_, new_n13136_, new_n13137_, new_n13138_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13479_, new_n13480_, new_n13481_,
    new_n13482_, new_n13483_, new_n13484_, new_n13485_, new_n13486_,
    new_n13487_, new_n13488_, new_n13489_, new_n13490_, new_n13491_,
    new_n13492_, new_n13493_, new_n13494_, new_n13495_, new_n13496_,
    new_n13497_, new_n13498_, new_n13499_, new_n13500_, new_n13501_,
    new_n13502_, new_n13503_, new_n13504_, new_n13505_, new_n13506_,
    new_n13507_, new_n13508_, new_n13509_, new_n13510_, new_n13511_,
    new_n13512_, new_n13513_, new_n13514_, new_n13515_, new_n13516_,
    new_n13517_, new_n13518_, new_n13519_, new_n13520_, new_n13521_,
    new_n13522_, new_n13523_, new_n13524_, new_n13525_, new_n13526_,
    new_n13527_, new_n13528_, new_n13529_, new_n13530_, new_n13531_,
    new_n13532_, new_n13533_, new_n13534_, new_n13535_, new_n13536_,
    new_n13537_, new_n13538_, new_n13539_, new_n13540_, new_n13541_,
    new_n13542_, new_n13543_, new_n13544_, new_n13545_, new_n13546_,
    new_n13547_, new_n13548_, new_n13549_, new_n13550_, new_n13551_,
    new_n13552_, new_n13553_, new_n13554_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13596_,
    new_n13597_, new_n13598_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13605_, new_n13606_,
    new_n13607_, new_n13608_, new_n13609_, new_n13610_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13637_, new_n13638_, new_n13639_, new_n13640_, new_n13641_,
    new_n13642_, new_n13643_, new_n13644_, new_n13645_, new_n13646_,
    new_n13647_, new_n13648_, new_n13649_, new_n13650_, new_n13651_,
    new_n13652_, new_n13653_, new_n13654_, new_n13655_, new_n13656_,
    new_n13657_, new_n13658_, new_n13659_, new_n13660_, new_n13661_,
    new_n13662_, new_n13663_, new_n13664_, new_n13665_, new_n13666_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13738_, new_n13739_, new_n13740_, new_n13741_, new_n13742_,
    new_n13743_, new_n13744_, new_n13745_, new_n13746_, new_n13747_,
    new_n13748_, new_n13749_, new_n13750_, new_n13751_, new_n13752_,
    new_n13753_, new_n13754_, new_n13755_, new_n13756_, new_n13757_,
    new_n13758_, new_n13759_, new_n13760_, new_n13761_, new_n13762_,
    new_n13763_, new_n13764_, new_n13765_, new_n13766_, new_n13767_,
    new_n13768_, new_n13769_, new_n13770_, new_n13771_, new_n13772_,
    new_n13773_, new_n13774_, new_n13775_, new_n13776_, new_n13777_,
    new_n13778_, new_n13779_, new_n13780_, new_n13781_, new_n13782_,
    new_n13783_, new_n13784_, new_n13785_, new_n13786_, new_n13787_,
    new_n13788_, new_n13789_, new_n13790_, new_n13791_, new_n13792_,
    new_n13793_, new_n13794_, new_n13795_, new_n13796_, new_n13797_,
    new_n13798_, new_n13799_, new_n13800_, new_n13801_, new_n13802_,
    new_n13803_, new_n13804_, new_n13805_, new_n13806_, new_n13807_,
    new_n13808_, new_n13809_, new_n13810_, new_n13811_, new_n13812_,
    new_n13813_, new_n13814_, new_n13815_, new_n13816_, new_n13817_,
    new_n13818_, new_n13819_, new_n13820_, new_n13821_, new_n13822_,
    new_n13823_, new_n13824_, new_n13825_, new_n13826_, new_n13827_,
    new_n13828_, new_n13829_, new_n13830_, new_n13831_, new_n13832_,
    new_n13833_, new_n13834_, new_n13835_, new_n13836_, new_n13837_,
    new_n13838_, new_n13839_, new_n13840_, new_n13841_, new_n13842_,
    new_n13843_, new_n13844_, new_n13845_, new_n13846_, new_n13847_,
    new_n13848_, new_n13849_, new_n13850_, new_n13851_, new_n13852_,
    new_n13853_, new_n13854_, new_n13855_, new_n13856_, new_n13857_,
    new_n13858_, new_n13859_, new_n13860_, new_n13861_, new_n13862_,
    new_n13863_, new_n13864_, new_n13865_, new_n13866_, new_n13867_,
    new_n13868_, new_n13869_, new_n13870_, new_n13871_, new_n13872_,
    new_n13873_, new_n13874_, new_n13875_, new_n13876_, new_n13877_,
    new_n13878_, new_n13879_, new_n13880_, new_n13881_, new_n13882_,
    new_n13883_, new_n13884_, new_n13885_, new_n13886_, new_n13887_,
    new_n13888_, new_n13889_, new_n13890_, new_n13891_, new_n13892_,
    new_n13893_, new_n13894_, new_n13895_, new_n13896_, new_n13897_,
    new_n13898_, new_n13899_, new_n13900_, new_n13901_, new_n13902_,
    new_n13903_, new_n13904_, new_n13905_, new_n13906_, new_n13907_,
    new_n13908_, new_n13909_, new_n13910_, new_n13911_, new_n13912_,
    new_n13913_, new_n13914_, new_n13915_, new_n13916_, new_n13917_,
    new_n13918_, new_n13919_, new_n13920_, new_n13921_, new_n13922_,
    new_n13923_, new_n13924_, new_n13925_, new_n13926_, new_n13927_,
    new_n13928_, new_n13929_, new_n13930_, new_n13931_, new_n13932_,
    new_n13933_, new_n13934_, new_n13935_, new_n13936_, new_n13937_,
    new_n13938_, new_n13939_, new_n13940_, new_n13941_, new_n13942_,
    new_n13943_, new_n13944_, new_n13945_, new_n13946_, new_n13947_,
    new_n13948_, new_n13949_, new_n13950_, new_n13951_, new_n13952_,
    new_n13953_, new_n13954_, new_n13955_, new_n13956_, new_n13957_,
    new_n13958_, new_n13959_, new_n13960_, new_n13961_, new_n13962_,
    new_n13963_, new_n13964_, new_n13965_, new_n13966_, new_n13967_,
    new_n13968_, new_n13969_, new_n13970_, new_n13971_, new_n13972_,
    new_n13973_, new_n13974_, new_n13975_, new_n13976_, new_n13977_,
    new_n13978_, new_n13979_, new_n13980_, new_n13981_, new_n13982_,
    new_n13983_, new_n13984_, new_n13985_, new_n13986_, new_n13987_,
    new_n13988_, new_n13989_, new_n13990_, new_n13991_, new_n13992_,
    new_n13993_, new_n13994_, new_n13995_, new_n13996_, new_n13997_,
    new_n13999_, new_n14000_, new_n14001_, new_n14002_, new_n14003_,
    new_n14004_, new_n14005_, new_n14006_, new_n14007_, new_n14008_,
    new_n14009_, new_n14010_, new_n14011_, new_n14012_, new_n14013_,
    new_n14014_, new_n14015_, new_n14016_, new_n14017_, new_n14018_,
    new_n14019_, new_n14020_, new_n14021_, new_n14022_, new_n14023_,
    new_n14024_, new_n14025_, new_n14026_, new_n14027_, new_n14028_,
    new_n14029_, new_n14030_, new_n14031_, new_n14032_, new_n14033_,
    new_n14034_, new_n14035_, new_n14036_, new_n14037_, new_n14038_,
    new_n14039_, new_n14040_, new_n14041_, new_n14042_, new_n14043_,
    new_n14044_, new_n14045_, new_n14046_, new_n14047_, new_n14048_,
    new_n14049_, new_n14050_, new_n14051_, new_n14052_, new_n14053_,
    new_n14054_, new_n14055_, new_n14056_, new_n14057_, new_n14058_,
    new_n14059_, new_n14060_, new_n14061_, new_n14062_, new_n14063_,
    new_n14064_, new_n14065_, new_n14066_, new_n14067_, new_n14068_,
    new_n14069_, new_n14070_, new_n14071_, new_n14072_, new_n14073_,
    new_n14074_, new_n14075_, new_n14076_, new_n14077_, new_n14078_,
    new_n14079_, new_n14080_, new_n14081_, new_n14082_, new_n14083_,
    new_n14084_, new_n14085_, new_n14086_, new_n14087_, new_n14088_,
    new_n14089_, new_n14090_, new_n14091_, new_n14092_, new_n14093_,
    new_n14094_, new_n14095_, new_n14096_, new_n14097_, new_n14098_,
    new_n14099_, new_n14100_, new_n14101_, new_n14102_, new_n14103_,
    new_n14104_, new_n14105_, new_n14106_, new_n14107_, new_n14108_,
    new_n14109_, new_n14110_, new_n14111_, new_n14112_, new_n14113_,
    new_n14114_, new_n14115_, new_n14116_, new_n14117_, new_n14118_,
    new_n14119_, new_n14120_, new_n14121_, new_n14122_, new_n14123_,
    new_n14124_, new_n14125_, new_n14126_, new_n14127_, new_n14128_,
    new_n14129_, new_n14130_, new_n14131_, new_n14132_, new_n14133_,
    new_n14134_, new_n14135_, new_n14136_, new_n14137_, new_n14138_,
    new_n14139_, new_n14140_, new_n14141_, new_n14142_, new_n14143_,
    new_n14144_, new_n14145_, new_n14146_, new_n14147_, new_n14148_,
    new_n14149_, new_n14150_, new_n14151_, new_n14152_, new_n14153_,
    new_n14154_, new_n14155_, new_n14156_, new_n14157_, new_n14158_,
    new_n14159_, new_n14160_, new_n14161_, new_n14162_, new_n14163_,
    new_n14164_, new_n14165_, new_n14166_, new_n14167_, new_n14168_,
    new_n14169_, new_n14170_, new_n14171_, new_n14172_, new_n14173_,
    new_n14174_, new_n14175_, new_n14176_, new_n14177_, new_n14178_,
    new_n14179_, new_n14180_, new_n14181_, new_n14182_, new_n14183_,
    new_n14184_, new_n14185_, new_n14186_, new_n14187_, new_n14188_,
    new_n14189_, new_n14190_, new_n14191_, new_n14192_, new_n14193_,
    new_n14194_, new_n14195_, new_n14196_, new_n14197_, new_n14198_,
    new_n14199_, new_n14200_, new_n14201_, new_n14202_, new_n14203_,
    new_n14204_, new_n14205_, new_n14206_, new_n14207_, new_n14208_,
    new_n14209_, new_n14210_, new_n14211_, new_n14212_, new_n14213_,
    new_n14214_, new_n14215_, new_n14216_, new_n14217_, new_n14218_,
    new_n14219_, new_n14220_, new_n14221_, new_n14222_, new_n14223_,
    new_n14224_, new_n14225_, new_n14226_, new_n14227_, new_n14228_,
    new_n14229_, new_n14230_, new_n14231_, new_n14232_, new_n14233_,
    new_n14234_, new_n14235_, new_n14236_, new_n14237_, new_n14238_,
    new_n14239_, new_n14240_, new_n14241_, new_n14242_, new_n14243_,
    new_n14244_, new_n14245_, new_n14246_, new_n14247_, new_n14248_,
    new_n14249_, new_n14250_, new_n14251_, new_n14252_, new_n14253_,
    new_n14254_, new_n14255_, new_n14256_, new_n14257_, new_n14258_,
    new_n14259_, new_n14260_, new_n14261_, new_n14262_, new_n14263_,
    new_n14264_, new_n14265_, new_n14266_, new_n14267_, new_n14268_,
    new_n14269_, new_n14271_, new_n14272_, new_n14273_, new_n14274_,
    new_n14275_, new_n14276_, new_n14277_, new_n14278_, new_n14279_,
    new_n14280_, new_n14281_, new_n14282_, new_n14283_, new_n14284_,
    new_n14285_, new_n14286_, new_n14287_, new_n14288_, new_n14289_,
    new_n14290_, new_n14291_, new_n14292_, new_n14293_, new_n14294_,
    new_n14295_, new_n14296_, new_n14297_, new_n14298_, new_n14299_,
    new_n14300_, new_n14301_, new_n14302_, new_n14303_, new_n14304_,
    new_n14305_, new_n14306_, new_n14307_, new_n14308_, new_n14309_,
    new_n14310_, new_n14311_, new_n14312_, new_n14313_, new_n14314_,
    new_n14315_, new_n14316_, new_n14317_, new_n14318_, new_n14319_,
    new_n14320_, new_n14321_, new_n14322_, new_n14323_, new_n14324_,
    new_n14325_, new_n14326_, new_n14327_, new_n14328_, new_n14329_,
    new_n14330_, new_n14331_, new_n14332_, new_n14333_, new_n14334_,
    new_n14335_, new_n14336_, new_n14337_, new_n14338_, new_n14339_,
    new_n14340_, new_n14341_, new_n14342_, new_n14343_, new_n14344_,
    new_n14345_, new_n14346_, new_n14347_, new_n14348_, new_n14349_,
    new_n14350_, new_n14351_, new_n14352_, new_n14353_, new_n14354_,
    new_n14355_, new_n14356_, new_n14357_, new_n14358_, new_n14359_,
    new_n14360_, new_n14361_, new_n14362_, new_n14363_, new_n14364_,
    new_n14365_, new_n14366_, new_n14367_, new_n14368_, new_n14369_,
    new_n14370_, new_n14371_, new_n14372_, new_n14373_, new_n14374_,
    new_n14375_, new_n14376_, new_n14377_, new_n14378_, new_n14379_,
    new_n14380_, new_n14381_, new_n14382_, new_n14383_, new_n14384_,
    new_n14385_, new_n14386_, new_n14387_, new_n14388_, new_n14389_,
    new_n14390_, new_n14391_, new_n14392_, new_n14393_, new_n14394_,
    new_n14395_, new_n14396_, new_n14397_, new_n14398_, new_n14399_,
    new_n14400_, new_n14401_, new_n14402_, new_n14403_, new_n14404_,
    new_n14405_, new_n14406_, new_n14407_, new_n14408_, new_n14409_,
    new_n14410_, new_n14411_, new_n14412_, new_n14413_, new_n14414_,
    new_n14415_, new_n14416_, new_n14417_, new_n14418_, new_n14419_,
    new_n14420_, new_n14421_, new_n14422_, new_n14423_, new_n14424_,
    new_n14425_, new_n14426_, new_n14427_, new_n14428_, new_n14429_,
    new_n14430_, new_n14431_, new_n14432_, new_n14433_, new_n14434_,
    new_n14435_, new_n14436_, new_n14437_, new_n14438_, new_n14439_,
    new_n14440_, new_n14441_, new_n14442_, new_n14443_, new_n14444_,
    new_n14445_, new_n14446_, new_n14447_, new_n14448_, new_n14449_,
    new_n14450_, new_n14451_, new_n14452_, new_n14453_, new_n14454_,
    new_n14455_, new_n14456_, new_n14457_, new_n14458_, new_n14459_,
    new_n14460_, new_n14461_, new_n14462_, new_n14463_, new_n14464_,
    new_n14465_, new_n14466_, new_n14467_, new_n14468_, new_n14469_,
    new_n14470_, new_n14471_, new_n14472_, new_n14473_, new_n14474_,
    new_n14475_, new_n14476_, new_n14477_, new_n14478_, new_n14479_,
    new_n14480_, new_n14481_, new_n14482_, new_n14483_, new_n14484_,
    new_n14485_, new_n14486_, new_n14487_, new_n14488_, new_n14489_,
    new_n14490_, new_n14491_, new_n14492_, new_n14493_, new_n14494_,
    new_n14495_, new_n14496_, new_n14497_, new_n14498_, new_n14499_,
    new_n14501_, new_n14502_, new_n14503_, new_n14504_, new_n14505_,
    new_n14506_, new_n14507_, new_n14508_, new_n14509_, new_n14510_,
    new_n14511_, new_n14512_, new_n14513_, new_n14514_, new_n14515_,
    new_n14516_, new_n14517_, new_n14518_, new_n14519_, new_n14520_,
    new_n14521_, new_n14522_, new_n14523_, new_n14524_, new_n14525_,
    new_n14526_, new_n14527_, new_n14528_, new_n14529_, new_n14530_,
    new_n14531_, new_n14532_, new_n14533_, new_n14534_, new_n14535_,
    new_n14536_, new_n14537_, new_n14538_, new_n14539_, new_n14540_,
    new_n14541_, new_n14542_, new_n14543_, new_n14544_, new_n14545_,
    new_n14546_, new_n14547_, new_n14548_, new_n14549_, new_n14550_,
    new_n14551_, new_n14552_, new_n14553_, new_n14554_, new_n14555_,
    new_n14556_, new_n14557_, new_n14558_, new_n14559_, new_n14560_,
    new_n14561_, new_n14562_, new_n14563_, new_n14564_, new_n14565_,
    new_n14566_, new_n14567_, new_n14568_, new_n14569_, new_n14570_,
    new_n14571_, new_n14572_, new_n14573_, new_n14574_, new_n14575_,
    new_n14576_, new_n14577_, new_n14578_, new_n14579_, new_n14580_,
    new_n14581_, new_n14582_, new_n14583_, new_n14584_, new_n14585_,
    new_n14586_, new_n14587_, new_n14588_, new_n14589_, new_n14590_,
    new_n14591_, new_n14592_, new_n14593_, new_n14594_, new_n14595_,
    new_n14596_, new_n14597_, new_n14598_, new_n14599_, new_n14600_,
    new_n14601_, new_n14602_, new_n14603_, new_n14604_, new_n14605_,
    new_n14606_, new_n14607_, new_n14608_, new_n14609_, new_n14610_,
    new_n14611_, new_n14612_, new_n14613_, new_n14614_, new_n14615_,
    new_n14616_, new_n14617_, new_n14618_, new_n14619_, new_n14620_,
    new_n14621_, new_n14622_, new_n14623_, new_n14624_, new_n14625_,
    new_n14626_, new_n14627_, new_n14628_, new_n14629_, new_n14630_,
    new_n14631_, new_n14632_, new_n14633_, new_n14634_, new_n14635_,
    new_n14636_, new_n14637_, new_n14638_, new_n14639_, new_n14640_,
    new_n14641_, new_n14642_, new_n14643_, new_n14644_, new_n14645_,
    new_n14646_, new_n14647_, new_n14648_, new_n14649_, new_n14650_,
    new_n14651_, new_n14652_, new_n14653_, new_n14654_, new_n14655_,
    new_n14656_, new_n14657_, new_n14658_, new_n14659_, new_n14660_,
    new_n14661_, new_n14662_, new_n14663_, new_n14664_, new_n14665_,
    new_n14666_, new_n14667_, new_n14668_, new_n14669_, new_n14670_,
    new_n14671_, new_n14672_, new_n14673_, new_n14674_, new_n14675_,
    new_n14676_, new_n14677_, new_n14678_, new_n14679_, new_n14680_,
    new_n14681_, new_n14682_, new_n14683_, new_n14684_, new_n14685_,
    new_n14686_, new_n14687_, new_n14688_, new_n14689_, new_n14690_,
    new_n14691_, new_n14692_, new_n14693_, new_n14694_, new_n14695_,
    new_n14696_, new_n14697_, new_n14698_, new_n14699_, new_n14700_,
    new_n14701_, new_n14702_, new_n14703_, new_n14704_, new_n14705_,
    new_n14706_, new_n14707_, new_n14708_, new_n14709_, new_n14710_,
    new_n14711_, new_n14712_, new_n14713_, new_n14714_, new_n14715_,
    new_n14716_, new_n14717_, new_n14718_, new_n14719_, new_n14720_,
    new_n14721_, new_n14722_, new_n14723_, new_n14724_, new_n14725_,
    new_n14726_, new_n14727_, new_n14728_, new_n14729_, new_n14730_,
    new_n14731_, new_n14732_, new_n14733_, new_n14734_, new_n14735_,
    new_n14736_, new_n14737_, new_n14738_, new_n14739_, new_n14740_,
    new_n14741_, new_n14742_, new_n14743_, new_n14745_, new_n14746_,
    new_n14747_, new_n14748_, new_n14749_, new_n14750_, new_n14751_,
    new_n14752_, new_n14753_, new_n14754_, new_n14755_, new_n14756_,
    new_n14757_, new_n14758_, new_n14759_, new_n14760_, new_n14761_,
    new_n14762_, new_n14763_, new_n14764_, new_n14765_, new_n14766_,
    new_n14767_, new_n14768_, new_n14769_, new_n14770_, new_n14771_,
    new_n14772_, new_n14773_, new_n14774_, new_n14775_, new_n14776_,
    new_n14777_, new_n14778_, new_n14779_, new_n14780_, new_n14781_,
    new_n14782_, new_n14783_, new_n14784_, new_n14785_, new_n14786_,
    new_n14787_, new_n14788_, new_n14789_, new_n14790_, new_n14791_,
    new_n14792_, new_n14793_, new_n14794_, new_n14795_, new_n14796_,
    new_n14797_, new_n14798_, new_n14799_, new_n14800_, new_n14801_,
    new_n14802_, new_n14803_, new_n14804_, new_n14805_, new_n14806_,
    new_n14807_, new_n14808_, new_n14809_, new_n14810_, new_n14811_,
    new_n14812_, new_n14813_, new_n14814_, new_n14815_, new_n14816_,
    new_n14817_, new_n14818_, new_n14819_, new_n14820_, new_n14821_,
    new_n14822_, new_n14823_, new_n14824_, new_n14825_, new_n14826_,
    new_n14827_, new_n14828_, new_n14829_, new_n14830_, new_n14831_,
    new_n14832_, new_n14833_, new_n14834_, new_n14835_, new_n14836_,
    new_n14837_, new_n14838_, new_n14839_, new_n14840_, new_n14841_,
    new_n14842_, new_n14843_, new_n14844_, new_n14845_, new_n14846_,
    new_n14847_, new_n14848_, new_n14849_, new_n14850_, new_n14851_,
    new_n14852_, new_n14853_, new_n14854_, new_n14855_, new_n14856_,
    new_n14857_, new_n14858_, new_n14859_, new_n14860_, new_n14861_,
    new_n14862_, new_n14863_, new_n14864_, new_n14865_, new_n14866_,
    new_n14867_, new_n14868_, new_n14869_, new_n14870_, new_n14871_,
    new_n14872_, new_n14873_, new_n14874_, new_n14875_, new_n14876_,
    new_n14877_, new_n14878_, new_n14879_, new_n14880_, new_n14881_,
    new_n14882_, new_n14883_, new_n14884_, new_n14885_, new_n14886_,
    new_n14887_, new_n14888_, new_n14889_, new_n14890_, new_n14891_,
    new_n14892_, new_n14893_, new_n14894_, new_n14895_, new_n14896_,
    new_n14897_, new_n14898_, new_n14899_, new_n14900_, new_n14901_,
    new_n14902_, new_n14903_, new_n14904_, new_n14905_, new_n14906_,
    new_n14907_, new_n14908_, new_n14909_, new_n14910_, new_n14911_,
    new_n14912_, new_n14913_, new_n14914_, new_n14915_, new_n14916_,
    new_n14917_, new_n14918_, new_n14919_, new_n14920_, new_n14921_,
    new_n14922_, new_n14923_, new_n14924_, new_n14925_, new_n14926_,
    new_n14927_, new_n14928_, new_n14929_, new_n14930_, new_n14931_,
    new_n14932_, new_n14933_, new_n14934_, new_n14935_, new_n14936_,
    new_n14937_, new_n14938_, new_n14939_, new_n14940_, new_n14941_,
    new_n14942_, new_n14943_, new_n14944_, new_n14945_, new_n14946_,
    new_n14947_, new_n14948_, new_n14949_, new_n14950_, new_n14951_,
    new_n14952_, new_n14953_, new_n14954_, new_n14955_, new_n14956_,
    new_n14957_, new_n14958_, new_n14959_, new_n14960_, new_n14961_,
    new_n14962_, new_n14963_, new_n14964_, new_n14965_, new_n14966_,
    new_n14967_, new_n14968_, new_n14969_, new_n14970_, new_n14971_,
    new_n14972_, new_n14973_, new_n14974_, new_n14975_, new_n14977_,
    new_n14978_, new_n14979_, new_n14980_, new_n14981_, new_n14982_,
    new_n14983_, new_n14984_, new_n14985_, new_n14986_, new_n14987_,
    new_n14988_, new_n14989_, new_n14990_, new_n14991_, new_n14992_,
    new_n14993_, new_n14994_, new_n14995_, new_n14996_, new_n14997_,
    new_n14998_, new_n14999_, new_n15000_, new_n15001_, new_n15002_,
    new_n15003_, new_n15004_, new_n15005_, new_n15006_, new_n15007_,
    new_n15008_, new_n15009_, new_n15010_, new_n15011_, new_n15012_,
    new_n15013_, new_n15014_, new_n15015_, new_n15016_, new_n15017_,
    new_n15018_, new_n15019_, new_n15020_, new_n15021_, new_n15022_,
    new_n15023_, new_n15024_, new_n15025_, new_n15026_, new_n15027_,
    new_n15028_, new_n15029_, new_n15030_, new_n15031_, new_n15032_,
    new_n15033_, new_n15034_, new_n15035_, new_n15036_, new_n15037_,
    new_n15038_, new_n15039_, new_n15040_, new_n15041_, new_n15042_,
    new_n15043_, new_n15044_, new_n15045_, new_n15046_, new_n15047_,
    new_n15048_, new_n15049_, new_n15050_, new_n15051_, new_n15052_,
    new_n15053_, new_n15054_, new_n15055_, new_n15056_, new_n15057_,
    new_n15058_, new_n15059_, new_n15060_, new_n15061_, new_n15062_,
    new_n15063_, new_n15064_, new_n15065_, new_n15066_, new_n15067_,
    new_n15068_, new_n15069_, new_n15070_, new_n15071_, new_n15072_,
    new_n15073_, new_n15074_, new_n15075_, new_n15076_, new_n15077_,
    new_n15078_, new_n15079_, new_n15080_, new_n15081_, new_n15082_,
    new_n15083_, new_n15084_, new_n15085_, new_n15086_, new_n15087_,
    new_n15088_, new_n15089_, new_n15090_, new_n15091_, new_n15092_,
    new_n15093_, new_n15094_, new_n15095_, new_n15096_, new_n15097_,
    new_n15098_, new_n15099_, new_n15100_, new_n15101_, new_n15102_,
    new_n15103_, new_n15104_, new_n15105_, new_n15106_, new_n15107_,
    new_n15108_, new_n15109_, new_n15110_, new_n15111_, new_n15112_,
    new_n15113_, new_n15114_, new_n15115_, new_n15116_, new_n15117_,
    new_n15118_, new_n15119_, new_n15120_, new_n15121_, new_n15122_,
    new_n15123_, new_n15124_, new_n15125_, new_n15126_, new_n15127_,
    new_n15128_, new_n15129_, new_n15130_, new_n15131_, new_n15132_,
    new_n15133_, new_n15134_, new_n15135_, new_n15136_, new_n15137_,
    new_n15138_, new_n15139_, new_n15140_, new_n15141_, new_n15142_,
    new_n15143_, new_n15144_, new_n15145_, new_n15146_, new_n15147_,
    new_n15148_, new_n15149_, new_n15150_, new_n15151_, new_n15152_,
    new_n15153_, new_n15154_, new_n15155_, new_n15156_, new_n15157_,
    new_n15158_, new_n15159_, new_n15160_, new_n15161_, new_n15162_,
    new_n15163_, new_n15164_, new_n15165_, new_n15166_, new_n15167_,
    new_n15168_, new_n15169_, new_n15170_, new_n15171_, new_n15172_,
    new_n15173_, new_n15174_, new_n15175_, new_n15176_, new_n15177_,
    new_n15178_, new_n15179_, new_n15180_, new_n15181_, new_n15182_,
    new_n15183_, new_n15184_, new_n15185_, new_n15186_, new_n15187_,
    new_n15188_, new_n15189_, new_n15190_, new_n15191_, new_n15192_,
    new_n15193_, new_n15194_, new_n15195_, new_n15196_, new_n15197_,
    new_n15198_, new_n15199_, new_n15200_, new_n15201_, new_n15202_,
    new_n15203_, new_n15204_, new_n15205_, new_n15206_, new_n15207_,
    new_n15208_, new_n15209_, new_n15210_, new_n15211_, new_n15212_,
    new_n15213_, new_n15214_, new_n15216_, new_n15217_, new_n15218_,
    new_n15219_, new_n15220_, new_n15221_, new_n15222_, new_n15223_,
    new_n15224_, new_n15225_, new_n15226_, new_n15227_, new_n15228_,
    new_n15229_, new_n15230_, new_n15231_, new_n15232_, new_n15233_,
    new_n15234_, new_n15235_, new_n15236_, new_n15237_, new_n15238_,
    new_n15239_, new_n15240_, new_n15241_, new_n15242_, new_n15243_,
    new_n15244_, new_n15245_, new_n15246_, new_n15247_, new_n15248_,
    new_n15249_, new_n15250_, new_n15251_, new_n15252_, new_n15253_,
    new_n15254_, new_n15255_, new_n15256_, new_n15257_, new_n15258_,
    new_n15259_, new_n15260_, new_n15261_, new_n15262_, new_n15263_,
    new_n15264_, new_n15265_, new_n15266_, new_n15267_, new_n15268_,
    new_n15269_, new_n15270_, new_n15271_, new_n15272_, new_n15273_,
    new_n15274_, new_n15275_, new_n15276_, new_n15277_, new_n15278_,
    new_n15279_, new_n15280_, new_n15281_, new_n15282_, new_n15283_,
    new_n15284_, new_n15285_, new_n15286_, new_n15287_, new_n15288_,
    new_n15289_, new_n15290_, new_n15291_, new_n15292_, new_n15293_,
    new_n15294_, new_n15295_, new_n15296_, new_n15297_, new_n15298_,
    new_n15299_, new_n15300_, new_n15301_, new_n15302_, new_n15303_,
    new_n15304_, new_n15305_, new_n15306_, new_n15307_, new_n15308_,
    new_n15309_, new_n15310_, new_n15311_, new_n15312_, new_n15313_,
    new_n15314_, new_n15315_, new_n15316_, new_n15317_, new_n15318_,
    new_n15319_, new_n15320_, new_n15321_, new_n15322_, new_n15323_,
    new_n15324_, new_n15325_, new_n15326_, new_n15327_, new_n15328_,
    new_n15329_, new_n15330_, new_n15331_, new_n15332_, new_n15333_,
    new_n15334_, new_n15335_, new_n15336_, new_n15337_, new_n15338_,
    new_n15339_, new_n15340_, new_n15341_, new_n15342_, new_n15343_,
    new_n15344_, new_n15345_, new_n15346_, new_n15347_, new_n15348_,
    new_n15349_, new_n15350_, new_n15351_, new_n15352_, new_n15353_,
    new_n15354_, new_n15355_, new_n15356_, new_n15357_, new_n15358_,
    new_n15359_, new_n15360_, new_n15361_, new_n15362_, new_n15363_,
    new_n15364_, new_n15365_, new_n15366_, new_n15367_, new_n15368_,
    new_n15369_, new_n15370_, new_n15371_, new_n15372_, new_n15373_,
    new_n15374_, new_n15375_, new_n15376_, new_n15377_, new_n15378_,
    new_n15379_, new_n15380_, new_n15381_, new_n15382_, new_n15383_,
    new_n15384_, new_n15385_, new_n15386_, new_n15387_, new_n15388_,
    new_n15389_, new_n15390_, new_n15391_, new_n15392_, new_n15393_,
    new_n15394_, new_n15395_, new_n15396_, new_n15397_, new_n15398_,
    new_n15399_, new_n15400_, new_n15401_, new_n15402_, new_n15403_,
    new_n15404_, new_n15405_, new_n15406_, new_n15407_, new_n15408_,
    new_n15409_, new_n15410_, new_n15411_, new_n15412_, new_n15413_,
    new_n15415_, new_n15416_, new_n15417_, new_n15418_, new_n15419_,
    new_n15420_, new_n15421_, new_n15422_, new_n15423_, new_n15424_,
    new_n15425_, new_n15426_, new_n15427_, new_n15428_, new_n15429_,
    new_n15430_, new_n15431_, new_n15432_, new_n15433_, new_n15434_,
    new_n15435_, new_n15436_, new_n15437_, new_n15438_, new_n15439_,
    new_n15440_, new_n15441_, new_n15442_, new_n15443_, new_n15444_,
    new_n15445_, new_n15446_, new_n15447_, new_n15448_, new_n15449_,
    new_n15450_, new_n15451_, new_n15452_, new_n15453_, new_n15454_,
    new_n15455_, new_n15456_, new_n15457_, new_n15458_, new_n15459_,
    new_n15460_, new_n15461_, new_n15462_, new_n15463_, new_n15464_,
    new_n15465_, new_n15466_, new_n15467_, new_n15468_, new_n15469_,
    new_n15470_, new_n15471_, new_n15472_, new_n15473_, new_n15474_,
    new_n15475_, new_n15476_, new_n15477_, new_n15478_, new_n15479_,
    new_n15480_, new_n15481_, new_n15482_, new_n15483_, new_n15484_,
    new_n15485_, new_n15486_, new_n15487_, new_n15488_, new_n15489_,
    new_n15490_, new_n15491_, new_n15492_, new_n15493_, new_n15494_,
    new_n15495_, new_n15496_, new_n15497_, new_n15498_, new_n15499_,
    new_n15500_, new_n15501_, new_n15502_, new_n15503_, new_n15504_,
    new_n15505_, new_n15506_, new_n15507_, new_n15508_, new_n15509_,
    new_n15510_, new_n15511_, new_n15512_, new_n15513_, new_n15514_,
    new_n15515_, new_n15516_, new_n15517_, new_n15518_, new_n15519_,
    new_n15520_, new_n15521_, new_n15522_, new_n15523_, new_n15524_,
    new_n15525_, new_n15526_, new_n15527_, new_n15528_, new_n15529_,
    new_n15530_, new_n15531_, new_n15532_, new_n15533_, new_n15534_,
    new_n15535_, new_n15536_, new_n15537_, new_n15538_, new_n15539_,
    new_n15540_, new_n15541_, new_n15542_, new_n15543_, new_n15544_,
    new_n15545_, new_n15546_, new_n15547_, new_n15548_, new_n15549_,
    new_n15550_, new_n15551_, new_n15552_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15558_, new_n15559_,
    new_n15560_, new_n15561_, new_n15562_, new_n15563_, new_n15564_,
    new_n15565_, new_n15566_, new_n15567_, new_n15568_, new_n15569_,
    new_n15570_, new_n15571_, new_n15572_, new_n15573_, new_n15574_,
    new_n15575_, new_n15576_, new_n15577_, new_n15578_, new_n15579_,
    new_n15580_, new_n15581_, new_n15582_, new_n15583_, new_n15584_,
    new_n15585_, new_n15586_, new_n15587_, new_n15588_, new_n15589_,
    new_n15590_, new_n15591_, new_n15592_, new_n15593_, new_n15594_,
    new_n15595_, new_n15596_, new_n15597_, new_n15598_, new_n15599_,
    new_n15600_, new_n15601_, new_n15602_, new_n15603_, new_n15604_,
    new_n15605_, new_n15606_, new_n15607_, new_n15608_, new_n15609_,
    new_n15610_, new_n15611_, new_n15612_, new_n15613_, new_n15614_,
    new_n15615_, new_n15616_, new_n15617_, new_n15618_, new_n15619_,
    new_n15620_, new_n15621_, new_n15622_, new_n15623_, new_n15624_,
    new_n15625_, new_n15626_, new_n15627_, new_n15628_, new_n15629_,
    new_n15630_, new_n15631_, new_n15632_, new_n15634_, new_n15635_,
    new_n15636_, new_n15637_, new_n15638_, new_n15639_, new_n15640_,
    new_n15641_, new_n15642_, new_n15643_, new_n15644_, new_n15645_,
    new_n15646_, new_n15647_, new_n15648_, new_n15649_, new_n15650_,
    new_n15651_, new_n15652_, new_n15653_, new_n15654_, new_n15655_,
    new_n15656_, new_n15657_, new_n15658_, new_n15659_, new_n15660_,
    new_n15661_, new_n15662_, new_n15663_, new_n15664_, new_n15665_,
    new_n15666_, new_n15667_, new_n15668_, new_n15669_, new_n15670_,
    new_n15671_, new_n15672_, new_n15673_, new_n15674_, new_n15675_,
    new_n15676_, new_n15677_, new_n15678_, new_n15679_, new_n15680_,
    new_n15681_, new_n15682_, new_n15683_, new_n15684_, new_n15685_,
    new_n15686_, new_n15687_, new_n15688_, new_n15689_, new_n15690_,
    new_n15691_, new_n15692_, new_n15693_, new_n15694_, new_n15695_,
    new_n15696_, new_n15697_, new_n15698_, new_n15699_, new_n15700_,
    new_n15701_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15741_, new_n15742_, new_n15743_, new_n15744_, new_n15745_,
    new_n15746_, new_n15747_, new_n15748_, new_n15749_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15781_, new_n15782_, new_n15783_, new_n15784_, new_n15785_,
    new_n15786_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15797_, new_n15798_, new_n15799_, new_n15800_,
    new_n15801_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15841_,
    new_n15842_, new_n15843_, new_n15844_, new_n15845_, new_n15846_,
    new_n15847_, new_n15848_, new_n15849_, new_n15850_, new_n15851_,
    new_n15852_, new_n15853_, new_n15854_, new_n15855_, new_n15856_,
    new_n15857_, new_n15858_, new_n15859_, new_n15860_, new_n15861_,
    new_n15862_, new_n15863_, new_n15864_, new_n15865_, new_n15866_,
    new_n15867_, new_n15868_, new_n15869_, new_n15870_, new_n15871_,
    new_n15872_, new_n15873_, new_n15874_, new_n15875_, new_n15876_,
    new_n15877_, new_n15878_, new_n15879_, new_n15880_, new_n15881_,
    new_n15882_, new_n15883_, new_n15884_, new_n15885_, new_n15886_,
    new_n15887_, new_n15888_, new_n15889_, new_n15890_, new_n15891_,
    new_n15892_, new_n15893_, new_n15894_, new_n15895_, new_n15896_,
    new_n15897_, new_n15898_, new_n15899_, new_n15900_, new_n15901_,
    new_n15902_, new_n15903_, new_n15904_, new_n15905_, new_n15906_,
    new_n15907_, new_n15908_, new_n15909_, new_n15910_, new_n15911_,
    new_n15912_, new_n15913_, new_n15914_, new_n15915_, new_n15916_,
    new_n15917_, new_n15918_, new_n15919_, new_n15920_, new_n15921_,
    new_n15922_, new_n15923_, new_n15924_, new_n15925_, new_n15926_,
    new_n15927_, new_n15928_, new_n15929_, new_n15930_, new_n15931_,
    new_n15932_, new_n15933_, new_n15934_, new_n15935_, new_n15936_,
    new_n15937_, new_n15938_, new_n15939_, new_n15940_, new_n15941_,
    new_n15942_, new_n15943_, new_n15944_, new_n15945_, new_n15946_,
    new_n15947_, new_n15948_, new_n15949_, new_n15950_, new_n15951_,
    new_n15952_, new_n15953_, new_n15954_, new_n15955_, new_n15956_,
    new_n15957_, new_n15958_, new_n15959_, new_n15960_, new_n15961_,
    new_n15962_, new_n15963_, new_n15964_, new_n15965_, new_n15966_,
    new_n15967_, new_n15968_, new_n15969_, new_n15970_, new_n15971_,
    new_n15972_, new_n15973_, new_n15974_, new_n15975_, new_n15976_,
    new_n15977_, new_n15978_, new_n15979_, new_n15980_, new_n15981_,
    new_n15982_, new_n15983_, new_n15984_, new_n15985_, new_n15986_,
    new_n15987_, new_n15988_, new_n15989_, new_n15990_, new_n15991_,
    new_n15992_, new_n15993_, new_n15994_, new_n15995_, new_n15996_,
    new_n15997_, new_n15998_, new_n15999_, new_n16000_, new_n16001_,
    new_n16002_, new_n16003_, new_n16004_, new_n16005_, new_n16006_,
    new_n16007_, new_n16008_, new_n16009_, new_n16010_, new_n16011_,
    new_n16012_, new_n16013_, new_n16014_, new_n16015_, new_n16016_,
    new_n16017_, new_n16018_, new_n16019_, new_n16020_, new_n16021_,
    new_n16022_, new_n16023_, new_n16024_, new_n16025_, new_n16026_,
    new_n16027_, new_n16028_, new_n16029_, new_n16030_, new_n16031_,
    new_n16032_, new_n16033_, new_n16034_, new_n16035_, new_n16037_,
    new_n16038_, new_n16039_, new_n16040_, new_n16041_, new_n16042_,
    new_n16043_, new_n16044_, new_n16045_, new_n16046_, new_n16047_,
    new_n16048_, new_n16049_, new_n16050_, new_n16051_, new_n16052_,
    new_n16053_, new_n16054_, new_n16055_, new_n16056_, new_n16057_,
    new_n16058_, new_n16059_, new_n16060_, new_n16061_, new_n16062_,
    new_n16063_, new_n16064_, new_n16065_, new_n16066_, new_n16067_,
    new_n16068_, new_n16069_, new_n16070_, new_n16071_, new_n16072_,
    new_n16073_, new_n16074_, new_n16075_, new_n16076_, new_n16077_,
    new_n16078_, new_n16079_, new_n16080_, new_n16081_, new_n16082_,
    new_n16083_, new_n16084_, new_n16085_, new_n16086_, new_n16087_,
    new_n16088_, new_n16089_, new_n16090_, new_n16091_, new_n16092_,
    new_n16093_, new_n16094_, new_n16095_, new_n16096_, new_n16097_,
    new_n16098_, new_n16099_, new_n16100_, new_n16101_, new_n16102_,
    new_n16103_, new_n16104_, new_n16105_, new_n16106_, new_n16107_,
    new_n16108_, new_n16109_, new_n16110_, new_n16111_, new_n16112_,
    new_n16113_, new_n16114_, new_n16115_, new_n16116_, new_n16117_,
    new_n16118_, new_n16119_, new_n16120_, new_n16121_, new_n16122_,
    new_n16123_, new_n16124_, new_n16125_, new_n16126_, new_n16127_,
    new_n16128_, new_n16129_, new_n16130_, new_n16131_, new_n16132_,
    new_n16133_, new_n16134_, new_n16135_, new_n16136_, new_n16137_,
    new_n16138_, new_n16139_, new_n16140_, new_n16141_, new_n16142_,
    new_n16143_, new_n16144_, new_n16145_, new_n16146_, new_n16147_,
    new_n16148_, new_n16149_, new_n16150_, new_n16151_, new_n16152_,
    new_n16153_, new_n16154_, new_n16155_, new_n16156_, new_n16157_,
    new_n16158_, new_n16159_, new_n16160_, new_n16161_, new_n16162_,
    new_n16163_, new_n16164_, new_n16165_, new_n16166_, new_n16167_,
    new_n16168_, new_n16169_, new_n16170_, new_n16171_, new_n16172_,
    new_n16173_, new_n16174_, new_n16175_, new_n16176_, new_n16177_,
    new_n16178_, new_n16179_, new_n16180_, new_n16181_, new_n16182_,
    new_n16183_, new_n16184_, new_n16185_, new_n16186_, new_n16187_,
    new_n16188_, new_n16189_, new_n16190_, new_n16191_, new_n16192_,
    new_n16193_, new_n16194_, new_n16195_, new_n16196_, new_n16197_,
    new_n16198_, new_n16199_, new_n16200_, new_n16201_, new_n16202_,
    new_n16203_, new_n16204_, new_n16205_, new_n16206_, new_n16207_,
    new_n16208_, new_n16209_, new_n16210_, new_n16211_, new_n16212_,
    new_n16213_, new_n16214_, new_n16215_, new_n16216_, new_n16217_,
    new_n16218_, new_n16219_, new_n16220_, new_n16221_, new_n16222_,
    new_n16223_, new_n16224_, new_n16225_, new_n16226_, new_n16227_,
    new_n16228_, new_n16229_, new_n16230_, new_n16231_, new_n16232_,
    new_n16234_, new_n16235_, new_n16236_, new_n16237_, new_n16238_,
    new_n16239_, new_n16240_, new_n16241_, new_n16242_, new_n16243_,
    new_n16244_, new_n16245_, new_n16246_, new_n16247_, new_n16248_,
    new_n16249_, new_n16250_, new_n16251_, new_n16252_, new_n16253_,
    new_n16254_, new_n16255_, new_n16256_, new_n16257_, new_n16258_,
    new_n16259_, new_n16260_, new_n16261_, new_n16262_, new_n16263_,
    new_n16264_, new_n16265_, new_n16266_, new_n16267_, new_n16268_,
    new_n16269_, new_n16270_, new_n16271_, new_n16272_, new_n16273_,
    new_n16274_, new_n16275_, new_n16276_, new_n16277_, new_n16278_,
    new_n16279_, new_n16280_, new_n16281_, new_n16282_, new_n16283_,
    new_n16284_, new_n16285_, new_n16286_, new_n16287_, new_n16288_,
    new_n16289_, new_n16290_, new_n16291_, new_n16292_, new_n16293_,
    new_n16294_, new_n16295_, new_n16296_, new_n16297_, new_n16298_,
    new_n16299_, new_n16300_, new_n16301_, new_n16302_, new_n16303_,
    new_n16304_, new_n16305_, new_n16306_, new_n16307_, new_n16308_,
    new_n16309_, new_n16310_, new_n16311_, new_n16312_, new_n16313_,
    new_n16314_, new_n16315_, new_n16316_, new_n16317_, new_n16318_,
    new_n16319_, new_n16320_, new_n16321_, new_n16322_, new_n16323_,
    new_n16324_, new_n16325_, new_n16326_, new_n16327_, new_n16328_,
    new_n16329_, new_n16330_, new_n16331_, new_n16332_, new_n16333_,
    new_n16334_, new_n16335_, new_n16336_, new_n16337_, new_n16338_,
    new_n16339_, new_n16340_, new_n16341_, new_n16342_, new_n16343_,
    new_n16344_, new_n16345_, new_n16346_, new_n16347_, new_n16348_,
    new_n16349_, new_n16350_, new_n16351_, new_n16352_, new_n16353_,
    new_n16354_, new_n16355_, new_n16356_, new_n16357_, new_n16358_,
    new_n16359_, new_n16360_, new_n16361_, new_n16362_, new_n16363_,
    new_n16364_, new_n16365_, new_n16366_, new_n16367_, new_n16368_,
    new_n16369_, new_n16370_, new_n16371_, new_n16372_, new_n16373_,
    new_n16374_, new_n16375_, new_n16376_, new_n16377_, new_n16378_,
    new_n16379_, new_n16380_, new_n16381_, new_n16382_, new_n16383_,
    new_n16384_, new_n16385_, new_n16386_, new_n16387_, new_n16388_,
    new_n16389_, new_n16390_, new_n16391_, new_n16392_, new_n16393_,
    new_n16394_, new_n16395_, new_n16396_, new_n16397_, new_n16398_,
    new_n16399_, new_n16400_, new_n16401_, new_n16402_, new_n16403_,
    new_n16404_, new_n16405_, new_n16406_, new_n16407_, new_n16408_,
    new_n16409_, new_n16410_, new_n16411_, new_n16412_, new_n16413_,
    new_n16414_, new_n16415_, new_n16416_, new_n16417_, new_n16418_,
    new_n16419_, new_n16420_, new_n16421_, new_n16422_, new_n16423_,
    new_n16424_, new_n16425_, new_n16426_, new_n16427_, new_n16429_,
    new_n16430_, new_n16431_, new_n16432_, new_n16433_, new_n16434_,
    new_n16435_, new_n16436_, new_n16437_, new_n16438_, new_n16439_,
    new_n16440_, new_n16441_, new_n16442_, new_n16443_, new_n16444_,
    new_n16445_, new_n16446_, new_n16447_, new_n16448_, new_n16449_,
    new_n16450_, new_n16451_, new_n16452_, new_n16453_, new_n16454_,
    new_n16455_, new_n16456_, new_n16457_, new_n16458_, new_n16459_,
    new_n16460_, new_n16461_, new_n16462_, new_n16463_, new_n16464_,
    new_n16465_, new_n16466_, new_n16467_, new_n16468_, new_n16469_,
    new_n16470_, new_n16471_, new_n16472_, new_n16473_, new_n16474_,
    new_n16475_, new_n16476_, new_n16477_, new_n16478_, new_n16479_,
    new_n16480_, new_n16481_, new_n16482_, new_n16483_, new_n16484_,
    new_n16485_, new_n16486_, new_n16487_, new_n16488_, new_n16489_,
    new_n16490_, new_n16491_, new_n16492_, new_n16493_, new_n16494_,
    new_n16495_, new_n16496_, new_n16497_, new_n16498_, new_n16499_,
    new_n16500_, new_n16501_, new_n16502_, new_n16503_, new_n16504_,
    new_n16505_, new_n16506_, new_n16507_, new_n16508_, new_n16509_,
    new_n16510_, new_n16511_, new_n16512_, new_n16513_, new_n16514_,
    new_n16515_, new_n16516_, new_n16517_, new_n16518_, new_n16519_,
    new_n16520_, new_n16521_, new_n16522_, new_n16523_, new_n16524_,
    new_n16525_, new_n16526_, new_n16527_, new_n16528_, new_n16529_,
    new_n16530_, new_n16531_, new_n16532_, new_n16533_, new_n16534_,
    new_n16535_, new_n16536_, new_n16537_, new_n16538_, new_n16539_,
    new_n16540_, new_n16541_, new_n16542_, new_n16543_, new_n16544_,
    new_n16545_, new_n16546_, new_n16547_, new_n16548_, new_n16549_,
    new_n16550_, new_n16551_, new_n16552_, new_n16553_, new_n16554_,
    new_n16555_, new_n16556_, new_n16557_, new_n16558_, new_n16559_,
    new_n16560_, new_n16561_, new_n16562_, new_n16563_, new_n16564_,
    new_n16565_, new_n16566_, new_n16567_, new_n16568_, new_n16569_,
    new_n16570_, new_n16571_, new_n16572_, new_n16573_, new_n16574_,
    new_n16575_, new_n16576_, new_n16577_, new_n16578_, new_n16579_,
    new_n16580_, new_n16581_, new_n16582_, new_n16583_, new_n16584_,
    new_n16585_, new_n16586_, new_n16587_, new_n16588_, new_n16589_,
    new_n16590_, new_n16591_, new_n16592_, new_n16593_, new_n16594_,
    new_n16595_, new_n16596_, new_n16597_, new_n16598_, new_n16599_,
    new_n16600_, new_n16601_, new_n16602_, new_n16603_, new_n16604_,
    new_n16605_, new_n16606_, new_n16607_, new_n16608_, new_n16609_,
    new_n16610_, new_n16611_, new_n16612_, new_n16613_, new_n16614_,
    new_n16615_, new_n16616_, new_n16617_, new_n16618_, new_n16619_,
    new_n16620_, new_n16621_, new_n16622_, new_n16623_, new_n16624_,
    new_n16625_, new_n16627_, new_n16628_, new_n16629_, new_n16630_,
    new_n16631_, new_n16632_, new_n16633_, new_n16634_, new_n16635_,
    new_n16636_, new_n16637_, new_n16638_, new_n16639_, new_n16640_,
    new_n16641_, new_n16642_, new_n16643_, new_n16644_, new_n16645_,
    new_n16646_, new_n16647_, new_n16648_, new_n16649_, new_n16650_,
    new_n16651_, new_n16652_, new_n16653_, new_n16654_, new_n16655_,
    new_n16656_, new_n16657_, new_n16658_, new_n16659_, new_n16660_,
    new_n16661_, new_n16662_, new_n16663_, new_n16664_, new_n16665_,
    new_n16666_, new_n16667_, new_n16668_, new_n16669_, new_n16670_,
    new_n16671_, new_n16672_, new_n16673_, new_n16674_, new_n16675_,
    new_n16676_, new_n16677_, new_n16678_, new_n16679_, new_n16680_,
    new_n16681_, new_n16682_, new_n16683_, new_n16684_, new_n16685_,
    new_n16686_, new_n16687_, new_n16688_, new_n16689_, new_n16690_,
    new_n16691_, new_n16692_, new_n16693_, new_n16694_, new_n16695_,
    new_n16696_, new_n16697_, new_n16698_, new_n16699_, new_n16700_,
    new_n16701_, new_n16702_, new_n16703_, new_n16704_, new_n16705_,
    new_n16706_, new_n16707_, new_n16708_, new_n16709_, new_n16710_,
    new_n16711_, new_n16712_, new_n16713_, new_n16714_, new_n16715_,
    new_n16716_, new_n16717_, new_n16718_, new_n16719_, new_n16720_,
    new_n16721_, new_n16722_, new_n16723_, new_n16724_, new_n16725_,
    new_n16726_, new_n16727_, new_n16728_, new_n16729_, new_n16730_,
    new_n16731_, new_n16732_, new_n16733_, new_n16734_, new_n16735_,
    new_n16736_, new_n16737_, new_n16738_, new_n16739_, new_n16740_,
    new_n16741_, new_n16742_, new_n16743_, new_n16744_, new_n16745_,
    new_n16746_, new_n16747_, new_n16748_, new_n16749_, new_n16750_,
    new_n16751_, new_n16752_, new_n16753_, new_n16754_, new_n16755_,
    new_n16756_, new_n16757_, new_n16758_, new_n16759_, new_n16760_,
    new_n16761_, new_n16762_, new_n16763_, new_n16764_, new_n16765_,
    new_n16766_, new_n16767_, new_n16768_, new_n16769_, new_n16770_,
    new_n16771_, new_n16772_, new_n16773_, new_n16774_, new_n16775_,
    new_n16776_, new_n16777_, new_n16778_, new_n16779_, new_n16780_,
    new_n16781_, new_n16782_, new_n16783_, new_n16784_, new_n16785_,
    new_n16786_, new_n16787_, new_n16788_, new_n16789_, new_n16790_,
    new_n16791_, new_n16792_, new_n16794_, new_n16795_, new_n16796_,
    new_n16797_, new_n16798_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16804_, new_n16805_, new_n16806_,
    new_n16807_, new_n16808_, new_n16809_, new_n16810_, new_n16811_,
    new_n16812_, new_n16813_, new_n16814_, new_n16815_, new_n16816_,
    new_n16817_, new_n16818_, new_n16819_, new_n16820_, new_n16821_,
    new_n16822_, new_n16823_, new_n16824_, new_n16825_, new_n16826_,
    new_n16827_, new_n16828_, new_n16829_, new_n16830_, new_n16831_,
    new_n16832_, new_n16833_, new_n16834_, new_n16835_, new_n16836_,
    new_n16837_, new_n16838_, new_n16839_, new_n16840_, new_n16841_,
    new_n16842_, new_n16843_, new_n16844_, new_n16845_, new_n16846_,
    new_n16847_, new_n16848_, new_n16849_, new_n16850_, new_n16851_,
    new_n16852_, new_n16853_, new_n16854_, new_n16855_, new_n16856_,
    new_n16857_, new_n16858_, new_n16859_, new_n16860_, new_n16861_,
    new_n16862_, new_n16863_, new_n16864_, new_n16865_, new_n16866_,
    new_n16867_, new_n16868_, new_n16869_, new_n16870_, new_n16871_,
    new_n16872_, new_n16873_, new_n16874_, new_n16875_, new_n16876_,
    new_n16877_, new_n16878_, new_n16879_, new_n16880_, new_n16881_,
    new_n16882_, new_n16883_, new_n16884_, new_n16885_, new_n16886_,
    new_n16887_, new_n16888_, new_n16889_, new_n16890_, new_n16891_,
    new_n16892_, new_n16893_, new_n16894_, new_n16895_, new_n16896_,
    new_n16897_, new_n16898_, new_n16899_, new_n16900_, new_n16901_,
    new_n16902_, new_n16903_, new_n16904_, new_n16905_, new_n16906_,
    new_n16907_, new_n16908_, new_n16909_, new_n16910_, new_n16911_,
    new_n16912_, new_n16913_, new_n16914_, new_n16915_, new_n16916_,
    new_n16917_, new_n16918_, new_n16919_, new_n16920_, new_n16921_,
    new_n16922_, new_n16923_, new_n16924_, new_n16925_, new_n16926_,
    new_n16927_, new_n16928_, new_n16929_, new_n16930_, new_n16931_,
    new_n16932_, new_n16933_, new_n16934_, new_n16935_, new_n16936_,
    new_n16937_, new_n16938_, new_n16939_, new_n16940_, new_n16941_,
    new_n16942_, new_n16943_, new_n16944_, new_n16945_, new_n16946_,
    new_n16947_, new_n16948_, new_n16949_, new_n16950_, new_n16951_,
    new_n16952_, new_n16953_, new_n16954_, new_n16955_, new_n16956_,
    new_n16957_, new_n16958_, new_n16959_, new_n16960_, new_n16961_,
    new_n16962_, new_n16963_, new_n16964_, new_n16965_, new_n16966_,
    new_n16967_, new_n16968_, new_n16969_, new_n16970_, new_n16971_,
    new_n16972_, new_n16973_, new_n16974_, new_n16975_, new_n16976_,
    new_n16977_, new_n16978_, new_n16979_, new_n16981_, new_n16982_,
    new_n16983_, new_n16984_, new_n16985_, new_n16986_, new_n16987_,
    new_n16988_, new_n16989_, new_n16990_, new_n16991_, new_n16992_,
    new_n16993_, new_n16994_, new_n16995_, new_n16996_, new_n16997_,
    new_n16998_, new_n16999_, new_n17000_, new_n17001_, new_n17002_,
    new_n17003_, new_n17004_, new_n17005_, new_n17006_, new_n17007_,
    new_n17008_, new_n17009_, new_n17010_, new_n17011_, new_n17012_,
    new_n17013_, new_n17014_, new_n17015_, new_n17016_, new_n17017_,
    new_n17018_, new_n17019_, new_n17020_, new_n17021_, new_n17022_,
    new_n17023_, new_n17024_, new_n17025_, new_n17026_, new_n17027_,
    new_n17028_, new_n17029_, new_n17030_, new_n17031_, new_n17032_,
    new_n17033_, new_n17034_, new_n17035_, new_n17036_, new_n17037_,
    new_n17038_, new_n17039_, new_n17040_, new_n17041_, new_n17042_,
    new_n17043_, new_n17044_, new_n17045_, new_n17046_, new_n17047_,
    new_n17048_, new_n17049_, new_n17050_, new_n17051_, new_n17052_,
    new_n17053_, new_n17054_, new_n17055_, new_n17056_, new_n17057_,
    new_n17058_, new_n17059_, new_n17060_, new_n17061_, new_n17062_,
    new_n17063_, new_n17064_, new_n17065_, new_n17066_, new_n17067_,
    new_n17068_, new_n17069_, new_n17070_, new_n17071_, new_n17072_,
    new_n17073_, new_n17074_, new_n17075_, new_n17076_, new_n17077_,
    new_n17078_, new_n17079_, new_n17080_, new_n17081_, new_n17082_,
    new_n17083_, new_n17084_, new_n17085_, new_n17086_, new_n17087_,
    new_n17088_, new_n17089_, new_n17090_, new_n17091_, new_n17092_,
    new_n17093_, new_n17094_, new_n17095_, new_n17096_, new_n17097_,
    new_n17098_, new_n17099_, new_n17100_, new_n17101_, new_n17102_,
    new_n17103_, new_n17104_, new_n17105_, new_n17106_, new_n17107_,
    new_n17108_, new_n17109_, new_n17110_, new_n17111_, new_n17112_,
    new_n17113_, new_n17114_, new_n17115_, new_n17116_, new_n17117_,
    new_n17118_, new_n17119_, new_n17120_, new_n17121_, new_n17122_,
    new_n17123_, new_n17124_, new_n17125_, new_n17126_, new_n17127_,
    new_n17128_, new_n17129_, new_n17130_, new_n17131_, new_n17132_,
    new_n17133_, new_n17134_, new_n17135_, new_n17136_, new_n17137_,
    new_n17138_, new_n17139_, new_n17140_, new_n17141_, new_n17142_,
    new_n17143_, new_n17144_, new_n17145_, new_n17146_, new_n17147_,
    new_n17148_, new_n17149_, new_n17150_, new_n17151_, new_n17152_,
    new_n17153_, new_n17154_, new_n17155_, new_n17156_, new_n17157_,
    new_n17159_, new_n17160_, new_n17161_, new_n17162_, new_n17163_,
    new_n17164_, new_n17165_, new_n17166_, new_n17167_, new_n17168_,
    new_n17169_, new_n17170_, new_n17171_, new_n17172_, new_n17173_,
    new_n17174_, new_n17175_, new_n17176_, new_n17177_, new_n17178_,
    new_n17179_, new_n17180_, new_n17181_, new_n17182_, new_n17183_,
    new_n17184_, new_n17185_, new_n17186_, new_n17187_, new_n17188_,
    new_n17189_, new_n17190_, new_n17191_, new_n17192_, new_n17193_,
    new_n17194_, new_n17195_, new_n17196_, new_n17197_, new_n17198_,
    new_n17199_, new_n17200_, new_n17201_, new_n17202_, new_n17203_,
    new_n17204_, new_n17205_, new_n17206_, new_n17207_, new_n17208_,
    new_n17209_, new_n17210_, new_n17211_, new_n17212_, new_n17213_,
    new_n17214_, new_n17215_, new_n17216_, new_n17217_, new_n17218_,
    new_n17219_, new_n17220_, new_n17221_, new_n17222_, new_n17223_,
    new_n17224_, new_n17225_, new_n17226_, new_n17227_, new_n17228_,
    new_n17229_, new_n17230_, new_n17231_, new_n17232_, new_n17233_,
    new_n17234_, new_n17235_, new_n17236_, new_n17237_, new_n17238_,
    new_n17239_, new_n17240_, new_n17241_, new_n17242_, new_n17243_,
    new_n17244_, new_n17245_, new_n17246_, new_n17247_, new_n17248_,
    new_n17249_, new_n17250_, new_n17251_, new_n17252_, new_n17253_,
    new_n17254_, new_n17255_, new_n17256_, new_n17257_, new_n17258_,
    new_n17259_, new_n17260_, new_n17261_, new_n17262_, new_n17263_,
    new_n17264_, new_n17265_, new_n17266_, new_n17267_, new_n17268_,
    new_n17269_, new_n17270_, new_n17271_, new_n17272_, new_n17273_,
    new_n17274_, new_n17275_, new_n17276_, new_n17277_, new_n17278_,
    new_n17279_, new_n17280_, new_n17281_, new_n17282_, new_n17283_,
    new_n17284_, new_n17285_, new_n17286_, new_n17287_, new_n17288_,
    new_n17289_, new_n17290_, new_n17291_, new_n17292_, new_n17293_,
    new_n17294_, new_n17295_, new_n17296_, new_n17297_, new_n17298_,
    new_n17299_, new_n17300_, new_n17301_, new_n17302_, new_n17303_,
    new_n17304_, new_n17305_, new_n17306_, new_n17307_, new_n17308_,
    new_n17309_, new_n17310_, new_n17311_, new_n17312_, new_n17313_,
    new_n17314_, new_n17315_, new_n17316_, new_n17317_, new_n17318_,
    new_n17319_, new_n17320_, new_n17321_, new_n17323_, new_n17324_,
    new_n17325_, new_n17326_, new_n17327_, new_n17328_, new_n17329_,
    new_n17330_, new_n17331_, new_n17332_, new_n17333_, new_n17334_,
    new_n17335_, new_n17336_, new_n17337_, new_n17338_, new_n17339_,
    new_n17340_, new_n17341_, new_n17342_, new_n17343_, new_n17344_,
    new_n17345_, new_n17346_, new_n17347_, new_n17348_, new_n17349_,
    new_n17350_, new_n17351_, new_n17352_, new_n17353_, new_n17354_,
    new_n17355_, new_n17356_, new_n17357_, new_n17358_, new_n17359_,
    new_n17360_, new_n17361_, new_n17362_, new_n17363_, new_n17364_,
    new_n17365_, new_n17366_, new_n17367_, new_n17368_, new_n17369_,
    new_n17370_, new_n17371_, new_n17372_, new_n17373_, new_n17374_,
    new_n17375_, new_n17376_, new_n17377_, new_n17378_, new_n17379_,
    new_n17380_, new_n17381_, new_n17382_, new_n17383_, new_n17384_,
    new_n17385_, new_n17386_, new_n17387_, new_n17388_, new_n17389_,
    new_n17390_, new_n17391_, new_n17392_, new_n17393_, new_n17394_,
    new_n17395_, new_n17396_, new_n17397_, new_n17398_, new_n17399_,
    new_n17400_, new_n17401_, new_n17402_, new_n17403_, new_n17404_,
    new_n17405_, new_n17406_, new_n17407_, new_n17408_, new_n17409_,
    new_n17410_, new_n17411_, new_n17412_, new_n17413_, new_n17414_,
    new_n17415_, new_n17416_, new_n17417_, new_n17418_, new_n17419_,
    new_n17420_, new_n17421_, new_n17422_, new_n17423_, new_n17424_,
    new_n17425_, new_n17426_, new_n17427_, new_n17428_, new_n17429_,
    new_n17430_, new_n17431_, new_n17432_, new_n17433_, new_n17434_,
    new_n17435_, new_n17436_, new_n17437_, new_n17438_, new_n17439_,
    new_n17440_, new_n17441_, new_n17442_, new_n17443_, new_n17444_,
    new_n17445_, new_n17446_, new_n17447_, new_n17448_, new_n17449_,
    new_n17450_, new_n17451_, new_n17452_, new_n17453_, new_n17454_,
    new_n17455_, new_n17456_, new_n17457_, new_n17458_, new_n17459_,
    new_n17460_, new_n17461_, new_n17462_, new_n17463_, new_n17464_,
    new_n17465_, new_n17466_, new_n17467_, new_n17468_, new_n17469_,
    new_n17470_, new_n17471_, new_n17472_, new_n17473_, new_n17474_,
    new_n17475_, new_n17476_, new_n17477_, new_n17478_, new_n17479_,
    new_n17480_, new_n17481_, new_n17482_, new_n17483_, new_n17484_,
    new_n17485_, new_n17486_, new_n17487_, new_n17488_, new_n17489_,
    new_n17490_, new_n17491_, new_n17492_, new_n17493_, new_n17494_,
    new_n17495_, new_n17496_, new_n17497_, new_n17498_, new_n17499_,
    new_n17500_, new_n17501_, new_n17502_, new_n17504_, new_n17505_,
    new_n17506_, new_n17507_, new_n17508_, new_n17509_, new_n17510_,
    new_n17511_, new_n17512_, new_n17513_, new_n17514_, new_n17515_,
    new_n17516_, new_n17517_, new_n17518_, new_n17519_, new_n17520_,
    new_n17521_, new_n17522_, new_n17523_, new_n17524_, new_n17525_,
    new_n17526_, new_n17527_, new_n17528_, new_n17529_, new_n17530_,
    new_n17531_, new_n17532_, new_n17533_, new_n17534_, new_n17535_,
    new_n17536_, new_n17537_, new_n17538_, new_n17539_, new_n17540_,
    new_n17541_, new_n17542_, new_n17543_, new_n17544_, new_n17545_,
    new_n17546_, new_n17547_, new_n17548_, new_n17549_, new_n17550_,
    new_n17551_, new_n17552_, new_n17553_, new_n17554_, new_n17555_,
    new_n17556_, new_n17557_, new_n17558_, new_n17559_, new_n17560_,
    new_n17561_, new_n17562_, new_n17563_, new_n17564_, new_n17565_,
    new_n17566_, new_n17567_, new_n17568_, new_n17569_, new_n17570_,
    new_n17571_, new_n17572_, new_n17573_, new_n17574_, new_n17575_,
    new_n17576_, new_n17577_, new_n17578_, new_n17579_, new_n17580_,
    new_n17581_, new_n17582_, new_n17583_, new_n17584_, new_n17585_,
    new_n17586_, new_n17587_, new_n17588_, new_n17589_, new_n17590_,
    new_n17591_, new_n17592_, new_n17593_, new_n17594_, new_n17595_,
    new_n17596_, new_n17597_, new_n17598_, new_n17599_, new_n17600_,
    new_n17601_, new_n17602_, new_n17603_, new_n17604_, new_n17605_,
    new_n17606_, new_n17607_, new_n17608_, new_n17609_, new_n17610_,
    new_n17611_, new_n17612_, new_n17613_, new_n17614_, new_n17615_,
    new_n17616_, new_n17617_, new_n17618_, new_n17619_, new_n17620_,
    new_n17621_, new_n17622_, new_n17623_, new_n17624_, new_n17625_,
    new_n17626_, new_n17627_, new_n17628_, new_n17629_, new_n17630_,
    new_n17631_, new_n17632_, new_n17633_, new_n17634_, new_n17635_,
    new_n17636_, new_n17637_, new_n17638_, new_n17639_, new_n17640_,
    new_n17641_, new_n17642_, new_n17643_, new_n17644_, new_n17645_,
    new_n17646_, new_n17647_, new_n17648_, new_n17649_, new_n17650_,
    new_n17651_, new_n17652_, new_n17653_, new_n17654_, new_n17655_,
    new_n17656_, new_n17657_, new_n17658_, new_n17659_, new_n17660_,
    new_n17661_, new_n17662_, new_n17663_, new_n17664_, new_n17665_,
    new_n17666_, new_n17668_, new_n17669_, new_n17670_, new_n17671_,
    new_n17672_, new_n17673_, new_n17674_, new_n17675_, new_n17676_,
    new_n17677_, new_n17678_, new_n17679_, new_n17680_, new_n17681_,
    new_n17682_, new_n17683_, new_n17684_, new_n17685_, new_n17686_,
    new_n17687_, new_n17688_, new_n17689_, new_n17690_, new_n17691_,
    new_n17692_, new_n17693_, new_n17694_, new_n17695_, new_n17696_,
    new_n17697_, new_n17698_, new_n17699_, new_n17700_, new_n17701_,
    new_n17702_, new_n17703_, new_n17704_, new_n17705_, new_n17706_,
    new_n17707_, new_n17708_, new_n17709_, new_n17710_, new_n17711_,
    new_n17712_, new_n17713_, new_n17714_, new_n17715_, new_n17716_,
    new_n17717_, new_n17718_, new_n17719_, new_n17720_, new_n17721_,
    new_n17722_, new_n17723_, new_n17724_, new_n17725_, new_n17726_,
    new_n17727_, new_n17728_, new_n17729_, new_n17730_, new_n17731_,
    new_n17732_, new_n17733_, new_n17734_, new_n17735_, new_n17736_,
    new_n17737_, new_n17738_, new_n17739_, new_n17740_, new_n17741_,
    new_n17742_, new_n17743_, new_n17744_, new_n17745_, new_n17746_,
    new_n17747_, new_n17748_, new_n17749_, new_n17750_, new_n17751_,
    new_n17752_, new_n17753_, new_n17754_, new_n17755_, new_n17756_,
    new_n17757_, new_n17758_, new_n17759_, new_n17760_, new_n17761_,
    new_n17762_, new_n17763_, new_n17764_, new_n17765_, new_n17766_,
    new_n17767_, new_n17768_, new_n17769_, new_n17770_, new_n17771_,
    new_n17772_, new_n17773_, new_n17774_, new_n17775_, new_n17776_,
    new_n17777_, new_n17778_, new_n17779_, new_n17780_, new_n17781_,
    new_n17782_, new_n17783_, new_n17784_, new_n17785_, new_n17786_,
    new_n17787_, new_n17788_, new_n17789_, new_n17790_, new_n17791_,
    new_n17792_, new_n17793_, new_n17794_, new_n17795_, new_n17796_,
    new_n17797_, new_n17798_, new_n17799_, new_n17800_, new_n17801_,
    new_n17802_, new_n17803_, new_n17804_, new_n17805_, new_n17806_,
    new_n17807_, new_n17808_, new_n17809_, new_n17810_, new_n17811_,
    new_n17812_, new_n17813_, new_n17814_, new_n17815_, new_n17816_,
    new_n17817_, new_n17818_, new_n17820_, new_n17821_, new_n17822_,
    new_n17823_, new_n17824_, new_n17825_, new_n17826_, new_n17827_,
    new_n17828_, new_n17829_, new_n17830_, new_n17831_, new_n17832_,
    new_n17833_, new_n17834_, new_n17835_, new_n17836_, new_n17837_,
    new_n17838_, new_n17839_, new_n17840_, new_n17841_, new_n17842_,
    new_n17843_, new_n17844_, new_n17845_, new_n17846_, new_n17847_,
    new_n17848_, new_n17849_, new_n17850_, new_n17851_, new_n17852_,
    new_n17853_, new_n17854_, new_n17855_, new_n17856_, new_n17857_,
    new_n17858_, new_n17859_, new_n17860_, new_n17861_, new_n17862_,
    new_n17863_, new_n17864_, new_n17865_, new_n17866_, new_n17867_,
    new_n17868_, new_n17869_, new_n17870_, new_n17871_, new_n17872_,
    new_n17873_, new_n17874_, new_n17875_, new_n17876_, new_n17877_,
    new_n17878_, new_n17879_, new_n17880_, new_n17881_, new_n17882_,
    new_n17883_, new_n17884_, new_n17885_, new_n17886_, new_n17887_,
    new_n17888_, new_n17889_, new_n17890_, new_n17891_, new_n17892_,
    new_n17893_, new_n17894_, new_n17895_, new_n17896_, new_n17897_,
    new_n17898_, new_n17899_, new_n17900_, new_n17901_, new_n17902_,
    new_n17903_, new_n17904_, new_n17905_, new_n17906_, new_n17907_,
    new_n17908_, new_n17909_, new_n17910_, new_n17911_, new_n17912_,
    new_n17913_, new_n17914_, new_n17915_, new_n17916_, new_n17917_,
    new_n17918_, new_n17919_, new_n17920_, new_n17921_, new_n17922_,
    new_n17923_, new_n17924_, new_n17925_, new_n17926_, new_n17927_,
    new_n17928_, new_n17929_, new_n17930_, new_n17931_, new_n17932_,
    new_n17933_, new_n17934_, new_n17935_, new_n17936_, new_n17937_,
    new_n17938_, new_n17939_, new_n17940_, new_n17941_, new_n17942_,
    new_n17943_, new_n17944_, new_n17945_, new_n17946_, new_n17947_,
    new_n17948_, new_n17949_, new_n17950_, new_n17951_, new_n17952_,
    new_n17953_, new_n17954_, new_n17955_, new_n17956_, new_n17957_,
    new_n17958_, new_n17959_, new_n17960_, new_n17961_, new_n17962_,
    new_n17963_, new_n17964_, new_n17965_, new_n17966_, new_n17967_,
    new_n17968_, new_n17969_, new_n17970_, new_n17971_, new_n17972_,
    new_n17973_, new_n17974_, new_n17975_, new_n17976_, new_n17977_,
    new_n17978_, new_n17979_, new_n17980_, new_n17981_, new_n17982_,
    new_n17983_, new_n17984_, new_n17985_, new_n17987_, new_n17988_,
    new_n17989_, new_n17990_, new_n17991_, new_n17992_, new_n17993_,
    new_n17994_, new_n17995_, new_n17996_, new_n17997_, new_n17998_,
    new_n17999_, new_n18000_, new_n18001_, new_n18002_, new_n18003_,
    new_n18004_, new_n18005_, new_n18006_, new_n18007_, new_n18008_,
    new_n18009_, new_n18010_, new_n18011_, new_n18012_, new_n18013_,
    new_n18014_, new_n18015_, new_n18016_, new_n18017_, new_n18018_,
    new_n18019_, new_n18020_, new_n18021_, new_n18022_, new_n18023_,
    new_n18024_, new_n18025_, new_n18026_, new_n18027_, new_n18028_,
    new_n18029_, new_n18030_, new_n18031_, new_n18032_, new_n18033_,
    new_n18034_, new_n18035_, new_n18036_, new_n18037_, new_n18038_,
    new_n18039_, new_n18040_, new_n18041_, new_n18042_, new_n18043_,
    new_n18044_, new_n18045_, new_n18046_, new_n18047_, new_n18048_,
    new_n18049_, new_n18050_, new_n18051_, new_n18052_, new_n18053_,
    new_n18054_, new_n18055_, new_n18056_, new_n18057_, new_n18058_,
    new_n18059_, new_n18060_, new_n18061_, new_n18062_, new_n18063_,
    new_n18064_, new_n18065_, new_n18066_, new_n18067_, new_n18068_,
    new_n18069_, new_n18070_, new_n18071_, new_n18072_, new_n18073_,
    new_n18074_, new_n18075_, new_n18076_, new_n18077_, new_n18078_,
    new_n18079_, new_n18080_, new_n18081_, new_n18082_, new_n18083_,
    new_n18084_, new_n18085_, new_n18086_, new_n18087_, new_n18088_,
    new_n18089_, new_n18090_, new_n18091_, new_n18092_, new_n18093_,
    new_n18094_, new_n18095_, new_n18096_, new_n18097_, new_n18098_,
    new_n18099_, new_n18100_, new_n18101_, new_n18102_, new_n18103_,
    new_n18104_, new_n18105_, new_n18106_, new_n18107_, new_n18108_,
    new_n18109_, new_n18110_, new_n18111_, new_n18112_, new_n18113_,
    new_n18114_, new_n18115_, new_n18116_, new_n18117_, new_n18118_,
    new_n18119_, new_n18120_, new_n18121_, new_n18122_, new_n18123_,
    new_n18124_, new_n18125_, new_n18126_, new_n18127_, new_n18128_,
    new_n18129_, new_n18130_, new_n18131_, new_n18132_, new_n18133_,
    new_n18134_, new_n18135_, new_n18136_, new_n18138_, new_n18139_,
    new_n18140_, new_n18141_, new_n18142_, new_n18143_, new_n18144_,
    new_n18145_, new_n18146_, new_n18147_, new_n18148_, new_n18149_,
    new_n18150_, new_n18151_, new_n18152_, new_n18153_, new_n18154_,
    new_n18155_, new_n18156_, new_n18157_, new_n18158_, new_n18159_,
    new_n18160_, new_n18161_, new_n18162_, new_n18163_, new_n18164_,
    new_n18165_, new_n18166_, new_n18167_, new_n18168_, new_n18169_,
    new_n18170_, new_n18171_, new_n18172_, new_n18173_, new_n18174_,
    new_n18175_, new_n18176_, new_n18177_, new_n18178_, new_n18179_,
    new_n18180_, new_n18181_, new_n18182_, new_n18183_, new_n18184_,
    new_n18185_, new_n18186_, new_n18187_, new_n18188_, new_n18189_,
    new_n18190_, new_n18191_, new_n18192_, new_n18193_, new_n18194_,
    new_n18195_, new_n18196_, new_n18197_, new_n18198_, new_n18199_,
    new_n18200_, new_n18201_, new_n18202_, new_n18203_, new_n18204_,
    new_n18205_, new_n18206_, new_n18207_, new_n18208_, new_n18209_,
    new_n18210_, new_n18211_, new_n18212_, new_n18213_, new_n18214_,
    new_n18215_, new_n18216_, new_n18217_, new_n18218_, new_n18219_,
    new_n18220_, new_n18221_, new_n18222_, new_n18223_, new_n18224_,
    new_n18225_, new_n18226_, new_n18227_, new_n18228_, new_n18229_,
    new_n18230_, new_n18231_, new_n18232_, new_n18233_, new_n18234_,
    new_n18235_, new_n18236_, new_n18237_, new_n18238_, new_n18239_,
    new_n18240_, new_n18241_, new_n18242_, new_n18243_, new_n18244_,
    new_n18245_, new_n18246_, new_n18247_, new_n18248_, new_n18249_,
    new_n18250_, new_n18251_, new_n18252_, new_n18253_, new_n18254_,
    new_n18255_, new_n18256_, new_n18257_, new_n18258_, new_n18259_,
    new_n18260_, new_n18261_, new_n18262_, new_n18263_, new_n18264_,
    new_n18265_, new_n18266_, new_n18267_, new_n18268_, new_n18269_,
    new_n18270_, new_n18271_, new_n18272_, new_n18273_, new_n18274_,
    new_n18275_, new_n18276_, new_n18277_, new_n18278_, new_n18279_,
    new_n18280_, new_n18281_, new_n18283_, new_n18284_, new_n18285_,
    new_n18286_, new_n18287_, new_n18288_, new_n18289_, new_n18290_,
    new_n18291_, new_n18292_, new_n18293_, new_n18294_, new_n18295_,
    new_n18296_, new_n18297_, new_n18298_, new_n18299_, new_n18300_,
    new_n18301_, new_n18302_, new_n18303_, new_n18304_, new_n18305_,
    new_n18306_, new_n18307_, new_n18308_, new_n18309_, new_n18310_,
    new_n18311_, new_n18312_, new_n18313_, new_n18314_, new_n18315_,
    new_n18316_, new_n18317_, new_n18318_, new_n18319_, new_n18320_,
    new_n18321_, new_n18322_, new_n18323_, new_n18324_, new_n18325_,
    new_n18326_, new_n18327_, new_n18328_, new_n18329_, new_n18330_,
    new_n18331_, new_n18332_, new_n18333_, new_n18334_, new_n18335_,
    new_n18336_, new_n18337_, new_n18338_, new_n18339_, new_n18340_,
    new_n18341_, new_n18342_, new_n18343_, new_n18344_, new_n18345_,
    new_n18346_, new_n18347_, new_n18348_, new_n18349_, new_n18350_,
    new_n18351_, new_n18352_, new_n18353_, new_n18354_, new_n18355_,
    new_n18356_, new_n18357_, new_n18358_, new_n18359_, new_n18360_,
    new_n18361_, new_n18362_, new_n18363_, new_n18364_, new_n18365_,
    new_n18366_, new_n18367_, new_n18368_, new_n18369_, new_n18370_,
    new_n18371_, new_n18372_, new_n18373_, new_n18374_, new_n18375_,
    new_n18376_, new_n18377_, new_n18378_, new_n18379_, new_n18380_,
    new_n18381_, new_n18382_, new_n18383_, new_n18384_, new_n18385_,
    new_n18386_, new_n18387_, new_n18388_, new_n18389_, new_n18390_,
    new_n18391_, new_n18392_, new_n18393_, new_n18394_, new_n18395_,
    new_n18396_, new_n18397_, new_n18398_, new_n18399_, new_n18400_,
    new_n18401_, new_n18402_, new_n18403_, new_n18404_, new_n18405_,
    new_n18406_, new_n18407_, new_n18408_, new_n18409_, new_n18410_,
    new_n18411_, new_n18412_, new_n18413_, new_n18414_, new_n18415_,
    new_n18416_, new_n18417_, new_n18418_, new_n18419_, new_n18420_,
    new_n18421_, new_n18422_, new_n18423_, new_n18424_, new_n18425_,
    new_n18426_, new_n18427_, new_n18428_, new_n18429_, new_n18430_,
    new_n18431_, new_n18432_, new_n18433_, new_n18434_, new_n18435_,
    new_n18436_, new_n18437_, new_n18438_, new_n18439_, new_n18440_,
    new_n18442_, new_n18443_, new_n18444_, new_n18445_, new_n18446_,
    new_n18447_, new_n18448_, new_n18449_, new_n18450_, new_n18451_,
    new_n18452_, new_n18453_, new_n18454_, new_n18455_, new_n18456_,
    new_n18457_, new_n18458_, new_n18459_, new_n18460_, new_n18461_,
    new_n18462_, new_n18463_, new_n18464_, new_n18465_, new_n18466_,
    new_n18467_, new_n18468_, new_n18469_, new_n18470_, new_n18471_,
    new_n18472_, new_n18473_, new_n18474_, new_n18475_, new_n18476_,
    new_n18477_, new_n18478_, new_n18479_, new_n18480_, new_n18481_,
    new_n18482_, new_n18483_, new_n18484_, new_n18485_, new_n18486_,
    new_n18487_, new_n18488_, new_n18489_, new_n18490_, new_n18491_,
    new_n18492_, new_n18493_, new_n18494_, new_n18495_, new_n18496_,
    new_n18497_, new_n18498_, new_n18499_, new_n18500_, new_n18501_,
    new_n18502_, new_n18503_, new_n18504_, new_n18505_, new_n18506_,
    new_n18507_, new_n18508_, new_n18509_, new_n18510_, new_n18511_,
    new_n18512_, new_n18513_, new_n18514_, new_n18515_, new_n18516_,
    new_n18517_, new_n18518_, new_n18519_, new_n18520_, new_n18521_,
    new_n18522_, new_n18523_, new_n18524_, new_n18525_, new_n18526_,
    new_n18527_, new_n18528_, new_n18529_, new_n18530_, new_n18531_,
    new_n18532_, new_n18533_, new_n18534_, new_n18535_, new_n18536_,
    new_n18537_, new_n18538_, new_n18539_, new_n18540_, new_n18541_,
    new_n18542_, new_n18543_, new_n18544_, new_n18545_, new_n18546_,
    new_n18547_, new_n18548_, new_n18549_, new_n18550_, new_n18551_,
    new_n18552_, new_n18553_, new_n18554_, new_n18555_, new_n18556_,
    new_n18557_, new_n18558_, new_n18559_, new_n18560_, new_n18561_,
    new_n18562_, new_n18563_, new_n18564_, new_n18565_, new_n18566_,
    new_n18567_, new_n18568_, new_n18569_, new_n18570_, new_n18571_,
    new_n18572_, new_n18573_, new_n18574_, new_n18575_, new_n18576_,
    new_n18578_, new_n18579_, new_n18580_, new_n18581_, new_n18582_,
    new_n18583_, new_n18584_, new_n18585_, new_n18586_, new_n18587_,
    new_n18588_, new_n18589_, new_n18590_, new_n18591_, new_n18592_,
    new_n18593_, new_n18594_, new_n18595_, new_n18596_, new_n18597_,
    new_n18598_, new_n18599_, new_n18600_, new_n18601_, new_n18602_,
    new_n18603_, new_n18604_, new_n18605_, new_n18606_, new_n18607_,
    new_n18608_, new_n18609_, new_n18610_, new_n18611_, new_n18612_,
    new_n18613_, new_n18614_, new_n18615_, new_n18616_, new_n18617_,
    new_n18618_, new_n18619_, new_n18620_, new_n18621_, new_n18622_,
    new_n18623_, new_n18624_, new_n18625_, new_n18626_, new_n18627_,
    new_n18628_, new_n18629_, new_n18630_, new_n18631_, new_n18632_,
    new_n18633_, new_n18634_, new_n18635_, new_n18636_, new_n18637_,
    new_n18638_, new_n18639_, new_n18640_, new_n18641_, new_n18642_,
    new_n18643_, new_n18644_, new_n18645_, new_n18646_, new_n18647_,
    new_n18648_, new_n18649_, new_n18650_, new_n18651_, new_n18652_,
    new_n18653_, new_n18654_, new_n18655_, new_n18656_, new_n18657_,
    new_n18658_, new_n18659_, new_n18660_, new_n18661_, new_n18662_,
    new_n18663_, new_n18664_, new_n18665_, new_n18666_, new_n18667_,
    new_n18668_, new_n18669_, new_n18670_, new_n18671_, new_n18672_,
    new_n18673_, new_n18674_, new_n18675_, new_n18676_, new_n18677_,
    new_n18678_, new_n18679_, new_n18680_, new_n18681_, new_n18682_,
    new_n18683_, new_n18684_, new_n18685_, new_n18686_, new_n18687_,
    new_n18688_, new_n18689_, new_n18690_, new_n18691_, new_n18692_,
    new_n18693_, new_n18694_, new_n18695_, new_n18696_, new_n18697_,
    new_n18698_, new_n18699_, new_n18700_, new_n18701_, new_n18702_,
    new_n18703_, new_n18704_, new_n18705_, new_n18706_, new_n18707_,
    new_n18708_, new_n18709_, new_n18710_, new_n18711_, new_n18712_,
    new_n18713_, new_n18715_, new_n18716_, new_n18717_, new_n18718_,
    new_n18719_, new_n18720_, new_n18721_, new_n18722_, new_n18723_,
    new_n18724_, new_n18725_, new_n18726_, new_n18727_, new_n18728_,
    new_n18729_, new_n18730_, new_n18731_, new_n18732_, new_n18733_,
    new_n18734_, new_n18735_, new_n18736_, new_n18737_, new_n18738_,
    new_n18739_, new_n18740_, new_n18741_, new_n18742_, new_n18743_,
    new_n18744_, new_n18745_, new_n18746_, new_n18747_, new_n18748_,
    new_n18749_, new_n18750_, new_n18751_, new_n18752_, new_n18753_,
    new_n18754_, new_n18755_, new_n18756_, new_n18757_, new_n18758_,
    new_n18759_, new_n18760_, new_n18761_, new_n18762_, new_n18763_,
    new_n18764_, new_n18765_, new_n18766_, new_n18767_, new_n18768_,
    new_n18769_, new_n18770_, new_n18771_, new_n18772_, new_n18773_,
    new_n18774_, new_n18775_, new_n18776_, new_n18777_, new_n18778_,
    new_n18779_, new_n18780_, new_n18781_, new_n18782_, new_n18783_,
    new_n18784_, new_n18785_, new_n18786_, new_n18787_, new_n18788_,
    new_n18789_, new_n18790_, new_n18791_, new_n18792_, new_n18793_,
    new_n18794_, new_n18795_, new_n18796_, new_n18797_, new_n18798_,
    new_n18799_, new_n18800_, new_n18801_, new_n18802_, new_n18803_,
    new_n18804_, new_n18805_, new_n18806_, new_n18807_, new_n18808_,
    new_n18809_, new_n18810_, new_n18811_, new_n18812_, new_n18813_,
    new_n18814_, new_n18815_, new_n18816_, new_n18817_, new_n18818_,
    new_n18819_, new_n18820_, new_n18821_, new_n18822_, new_n18823_,
    new_n18824_, new_n18825_, new_n18826_, new_n18827_, new_n18828_,
    new_n18829_, new_n18830_, new_n18831_, new_n18832_, new_n18833_,
    new_n18834_, new_n18835_, new_n18836_, new_n18837_, new_n18838_,
    new_n18839_, new_n18840_, new_n18841_, new_n18842_, new_n18843_,
    new_n18844_, new_n18845_, new_n18846_, new_n18847_, new_n18848_,
    new_n18850_, new_n18851_, new_n18852_, new_n18853_, new_n18854_,
    new_n18855_, new_n18856_, new_n18857_, new_n18858_, new_n18859_,
    new_n18860_, new_n18861_, new_n18862_, new_n18863_, new_n18864_,
    new_n18865_, new_n18866_, new_n18867_, new_n18868_, new_n18869_,
    new_n18870_, new_n18871_, new_n18872_, new_n18873_, new_n18874_,
    new_n18875_, new_n18876_, new_n18877_, new_n18878_, new_n18879_,
    new_n18880_, new_n18881_, new_n18882_, new_n18883_, new_n18884_,
    new_n18885_, new_n18886_, new_n18887_, new_n18888_, new_n18889_,
    new_n18890_, new_n18891_, new_n18892_, new_n18893_, new_n18894_,
    new_n18895_, new_n18896_, new_n18897_, new_n18898_, new_n18899_,
    new_n18900_, new_n18901_, new_n18902_, new_n18903_, new_n18904_,
    new_n18905_, new_n18906_, new_n18907_, new_n18908_, new_n18909_,
    new_n18910_, new_n18911_, new_n18912_, new_n18913_, new_n18914_,
    new_n18915_, new_n18916_, new_n18917_, new_n18918_, new_n18919_,
    new_n18920_, new_n18921_, new_n18922_, new_n18923_, new_n18924_,
    new_n18925_, new_n18926_, new_n18927_, new_n18928_, new_n18929_,
    new_n18930_, new_n18931_, new_n18932_, new_n18933_, new_n18934_,
    new_n18935_, new_n18936_, new_n18937_, new_n18938_, new_n18939_,
    new_n18940_, new_n18941_, new_n18942_, new_n18943_, new_n18944_,
    new_n18945_, new_n18946_, new_n18947_, new_n18948_, new_n18949_,
    new_n18950_, new_n18951_, new_n18952_, new_n18953_, new_n18954_,
    new_n18955_, new_n18956_, new_n18957_, new_n18958_, new_n18959_,
    new_n18960_, new_n18961_, new_n18962_, new_n18963_, new_n18964_,
    new_n18965_, new_n18966_, new_n18967_, new_n18968_, new_n18969_,
    new_n18970_, new_n18971_, new_n18972_, new_n18973_, new_n18974_,
    new_n18975_, new_n18976_, new_n18977_, new_n18978_, new_n18979_,
    new_n18980_, new_n18982_, new_n18983_, new_n18984_, new_n18985_,
    new_n18986_, new_n18987_, new_n18988_, new_n18989_, new_n18990_,
    new_n18991_, new_n18992_, new_n18993_, new_n18994_, new_n18995_,
    new_n18996_, new_n18997_, new_n18998_, new_n18999_, new_n19000_,
    new_n19001_, new_n19002_, new_n19003_, new_n19004_, new_n19005_,
    new_n19006_, new_n19007_, new_n19008_, new_n19009_, new_n19010_,
    new_n19011_, new_n19012_, new_n19013_, new_n19014_, new_n19015_,
    new_n19016_, new_n19017_, new_n19018_, new_n19019_, new_n19020_,
    new_n19021_, new_n19022_, new_n19023_, new_n19024_, new_n19025_,
    new_n19026_, new_n19027_, new_n19028_, new_n19029_, new_n19030_,
    new_n19031_, new_n19032_, new_n19033_, new_n19034_, new_n19035_,
    new_n19036_, new_n19037_, new_n19038_, new_n19039_, new_n19040_,
    new_n19041_, new_n19042_, new_n19043_, new_n19044_, new_n19045_,
    new_n19046_, new_n19047_, new_n19048_, new_n19049_, new_n19050_,
    new_n19051_, new_n19052_, new_n19053_, new_n19054_, new_n19055_,
    new_n19056_, new_n19057_, new_n19058_, new_n19059_, new_n19060_,
    new_n19061_, new_n19062_, new_n19063_, new_n19064_, new_n19065_,
    new_n19066_, new_n19067_, new_n19068_, new_n19069_, new_n19070_,
    new_n19071_, new_n19072_, new_n19073_, new_n19074_, new_n19075_,
    new_n19076_, new_n19077_, new_n19078_, new_n19079_, new_n19080_,
    new_n19081_, new_n19082_, new_n19083_, new_n19084_, new_n19085_,
    new_n19086_, new_n19087_, new_n19088_, new_n19089_, new_n19090_,
    new_n19091_, new_n19092_, new_n19093_, new_n19094_, new_n19095_,
    new_n19096_, new_n19097_, new_n19098_, new_n19099_, new_n19100_,
    new_n19101_, new_n19102_, new_n19103_, new_n19104_, new_n19105_,
    new_n19106_, new_n19108_, new_n19109_, new_n19110_, new_n19111_,
    new_n19112_, new_n19113_, new_n19114_, new_n19115_, new_n19116_,
    new_n19117_, new_n19118_, new_n19119_, new_n19120_, new_n19121_,
    new_n19122_, new_n19123_, new_n19124_, new_n19125_, new_n19126_,
    new_n19127_, new_n19128_, new_n19129_, new_n19130_, new_n19131_,
    new_n19132_, new_n19133_, new_n19134_, new_n19135_, new_n19136_,
    new_n19137_, new_n19138_, new_n19139_, new_n19140_, new_n19141_,
    new_n19142_, new_n19143_, new_n19144_, new_n19145_, new_n19146_,
    new_n19147_, new_n19148_, new_n19149_, new_n19150_, new_n19151_,
    new_n19152_, new_n19153_, new_n19154_, new_n19155_, new_n19156_,
    new_n19157_, new_n19158_, new_n19159_, new_n19160_, new_n19161_,
    new_n19162_, new_n19163_, new_n19164_, new_n19165_, new_n19166_,
    new_n19167_, new_n19168_, new_n19169_, new_n19170_, new_n19171_,
    new_n19172_, new_n19173_, new_n19174_, new_n19175_, new_n19176_,
    new_n19177_, new_n19178_, new_n19179_, new_n19180_, new_n19181_,
    new_n19182_, new_n19183_, new_n19184_, new_n19185_, new_n19186_,
    new_n19187_, new_n19188_, new_n19189_, new_n19190_, new_n19191_,
    new_n19192_, new_n19193_, new_n19194_, new_n19195_, new_n19196_,
    new_n19197_, new_n19198_, new_n19199_, new_n19200_, new_n19201_,
    new_n19202_, new_n19203_, new_n19204_, new_n19205_, new_n19206_,
    new_n19207_, new_n19208_, new_n19209_, new_n19210_, new_n19211_,
    new_n19212_, new_n19213_, new_n19214_, new_n19215_, new_n19216_,
    new_n19217_, new_n19218_, new_n19219_, new_n19220_, new_n19221_,
    new_n19222_, new_n19223_, new_n19224_, new_n19225_, new_n19226_,
    new_n19227_, new_n19228_, new_n19229_, new_n19230_, new_n19231_,
    new_n19232_, new_n19233_, new_n19235_, new_n19236_, new_n19237_,
    new_n19238_, new_n19239_, new_n19240_, new_n19241_, new_n19242_,
    new_n19243_, new_n19244_, new_n19245_, new_n19246_, new_n19247_,
    new_n19248_, new_n19249_, new_n19250_, new_n19251_, new_n19252_,
    new_n19253_, new_n19254_, new_n19255_, new_n19256_, new_n19257_,
    new_n19258_, new_n19259_, new_n19260_, new_n19261_, new_n19262_,
    new_n19263_, new_n19264_, new_n19265_, new_n19266_, new_n19267_,
    new_n19268_, new_n19269_, new_n19270_, new_n19271_, new_n19272_,
    new_n19273_, new_n19274_, new_n19275_, new_n19276_, new_n19277_,
    new_n19278_, new_n19279_, new_n19280_, new_n19281_, new_n19282_,
    new_n19283_, new_n19284_, new_n19285_, new_n19286_, new_n19287_,
    new_n19288_, new_n19289_, new_n19290_, new_n19291_, new_n19292_,
    new_n19293_, new_n19294_, new_n19295_, new_n19296_, new_n19297_,
    new_n19298_, new_n19299_, new_n19300_, new_n19301_, new_n19302_,
    new_n19303_, new_n19304_, new_n19305_, new_n19306_, new_n19307_,
    new_n19308_, new_n19309_, new_n19310_, new_n19311_, new_n19312_,
    new_n19313_, new_n19314_, new_n19315_, new_n19316_, new_n19317_,
    new_n19318_, new_n19319_, new_n19320_, new_n19321_, new_n19322_,
    new_n19323_, new_n19324_, new_n19325_, new_n19326_, new_n19327_,
    new_n19328_, new_n19329_, new_n19330_, new_n19331_, new_n19332_,
    new_n19333_, new_n19334_, new_n19335_, new_n19336_, new_n19337_,
    new_n19338_, new_n19339_, new_n19340_, new_n19341_, new_n19342_,
    new_n19343_, new_n19344_, new_n19345_, new_n19346_, new_n19347_,
    new_n19348_, new_n19349_, new_n19350_, new_n19351_, new_n19352_,
    new_n19353_, new_n19355_, new_n19356_, new_n19357_, new_n19358_,
    new_n19359_, new_n19360_, new_n19361_, new_n19362_, new_n19363_,
    new_n19364_, new_n19365_, new_n19366_, new_n19367_, new_n19368_,
    new_n19369_, new_n19370_, new_n19371_, new_n19372_, new_n19373_,
    new_n19374_, new_n19375_, new_n19376_, new_n19377_, new_n19378_,
    new_n19379_, new_n19380_, new_n19381_, new_n19382_, new_n19383_,
    new_n19384_, new_n19385_, new_n19386_, new_n19387_, new_n19388_,
    new_n19389_, new_n19390_, new_n19391_, new_n19392_, new_n19393_,
    new_n19394_, new_n19395_, new_n19396_, new_n19397_, new_n19398_,
    new_n19399_, new_n19400_, new_n19401_, new_n19402_, new_n19403_,
    new_n19404_, new_n19405_, new_n19406_, new_n19407_, new_n19408_,
    new_n19409_, new_n19410_, new_n19411_, new_n19412_, new_n19413_,
    new_n19414_, new_n19415_, new_n19416_, new_n19417_, new_n19418_,
    new_n19419_, new_n19420_, new_n19421_, new_n19422_, new_n19423_,
    new_n19424_, new_n19425_, new_n19426_, new_n19427_, new_n19428_,
    new_n19429_, new_n19430_, new_n19431_, new_n19432_, new_n19433_,
    new_n19434_, new_n19435_, new_n19436_, new_n19437_, new_n19438_,
    new_n19439_, new_n19440_, new_n19441_, new_n19442_, new_n19443_,
    new_n19444_, new_n19445_, new_n19446_, new_n19447_, new_n19448_,
    new_n19449_, new_n19450_, new_n19451_, new_n19452_, new_n19453_,
    new_n19454_, new_n19455_, new_n19456_, new_n19457_, new_n19458_,
    new_n19459_, new_n19460_, new_n19461_, new_n19462_, new_n19463_,
    new_n19464_, new_n19465_, new_n19466_, new_n19467_, new_n19468_,
    new_n19469_, new_n19470_, new_n19472_, new_n19473_, new_n19474_,
    new_n19475_, new_n19476_, new_n19477_, new_n19478_, new_n19479_,
    new_n19480_, new_n19481_, new_n19482_, new_n19483_, new_n19484_,
    new_n19485_, new_n19486_, new_n19487_, new_n19488_, new_n19489_,
    new_n19490_, new_n19491_, new_n19492_, new_n19493_, new_n19494_,
    new_n19495_, new_n19496_, new_n19497_, new_n19498_, new_n19499_,
    new_n19500_, new_n19501_, new_n19502_, new_n19503_, new_n19504_,
    new_n19505_, new_n19506_, new_n19507_, new_n19508_, new_n19509_,
    new_n19510_, new_n19511_, new_n19512_, new_n19513_, new_n19514_,
    new_n19515_, new_n19516_, new_n19517_, new_n19518_, new_n19519_,
    new_n19520_, new_n19521_, new_n19522_, new_n19523_, new_n19524_,
    new_n19525_, new_n19526_, new_n19527_, new_n19528_, new_n19529_,
    new_n19530_, new_n19531_, new_n19532_, new_n19533_, new_n19534_,
    new_n19535_, new_n19536_, new_n19537_, new_n19538_, new_n19539_,
    new_n19540_, new_n19541_, new_n19542_, new_n19543_, new_n19544_,
    new_n19545_, new_n19546_, new_n19547_, new_n19548_, new_n19549_,
    new_n19550_, new_n19551_, new_n19552_, new_n19553_, new_n19554_,
    new_n19555_, new_n19556_, new_n19557_, new_n19558_, new_n19559_,
    new_n19560_, new_n19561_, new_n19562_, new_n19563_, new_n19564_,
    new_n19565_, new_n19566_, new_n19567_, new_n19568_, new_n19569_,
    new_n19570_, new_n19571_, new_n19572_, new_n19573_, new_n19574_,
    new_n19575_, new_n19576_, new_n19577_, new_n19578_, new_n19579_,
    new_n19580_, new_n19581_, new_n19582_, new_n19583_, new_n19584_,
    new_n19585_, new_n19587_, new_n19588_, new_n19589_, new_n19590_,
    new_n19591_, new_n19592_, new_n19593_, new_n19594_, new_n19595_,
    new_n19596_, new_n19597_, new_n19598_, new_n19599_, new_n19600_,
    new_n19601_, new_n19602_, new_n19603_, new_n19604_, new_n19605_,
    new_n19606_, new_n19607_, new_n19608_, new_n19609_, new_n19610_,
    new_n19611_, new_n19612_, new_n19613_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19636_, new_n19637_, new_n19638_, new_n19639_, new_n19640_,
    new_n19641_, new_n19642_, new_n19643_, new_n19644_, new_n19645_,
    new_n19646_, new_n19647_, new_n19648_, new_n19649_, new_n19650_,
    new_n19651_, new_n19652_, new_n19653_, new_n19654_, new_n19655_,
    new_n19656_, new_n19657_, new_n19658_, new_n19659_, new_n19660_,
    new_n19661_, new_n19662_, new_n19663_, new_n19664_, new_n19665_,
    new_n19666_, new_n19667_, new_n19668_, new_n19669_, new_n19670_,
    new_n19671_, new_n19672_, new_n19673_, new_n19674_, new_n19675_,
    new_n19676_, new_n19677_, new_n19678_, new_n19679_, new_n19680_,
    new_n19681_, new_n19682_, new_n19683_, new_n19684_, new_n19685_,
    new_n19686_, new_n19687_, new_n19688_, new_n19689_, new_n19690_,
    new_n19691_, new_n19692_, new_n19693_, new_n19694_, new_n19695_,
    new_n19696_, new_n19697_, new_n19699_, new_n19700_, new_n19701_,
    new_n19702_, new_n19703_, new_n19704_, new_n19705_, new_n19706_,
    new_n19707_, new_n19708_, new_n19709_, new_n19710_, new_n19711_,
    new_n19712_, new_n19713_, new_n19714_, new_n19715_, new_n19716_,
    new_n19717_, new_n19718_, new_n19719_, new_n19720_, new_n19721_,
    new_n19722_, new_n19723_, new_n19724_, new_n19725_, new_n19726_,
    new_n19727_, new_n19728_, new_n19729_, new_n19730_, new_n19731_,
    new_n19732_, new_n19733_, new_n19734_, new_n19735_, new_n19736_,
    new_n19737_, new_n19738_, new_n19739_, new_n19740_, new_n19741_,
    new_n19742_, new_n19743_, new_n19744_, new_n19745_, new_n19746_,
    new_n19747_, new_n19748_, new_n19749_, new_n19750_, new_n19751_,
    new_n19752_, new_n19753_, new_n19754_, new_n19755_, new_n19756_,
    new_n19757_, new_n19758_, new_n19759_, new_n19760_, new_n19761_,
    new_n19762_, new_n19763_, new_n19764_, new_n19765_, new_n19766_,
    new_n19767_, new_n19768_, new_n19769_, new_n19770_, new_n19771_,
    new_n19772_, new_n19773_, new_n19774_, new_n19775_, new_n19776_,
    new_n19777_, new_n19778_, new_n19779_, new_n19780_, new_n19781_,
    new_n19782_, new_n19783_, new_n19784_, new_n19785_, new_n19786_,
    new_n19787_, new_n19788_, new_n19789_, new_n19790_, new_n19791_,
    new_n19792_, new_n19793_, new_n19794_, new_n19795_, new_n19796_,
    new_n19797_, new_n19798_, new_n19799_, new_n19800_, new_n19801_,
    new_n19802_, new_n19803_, new_n19805_, new_n19806_, new_n19807_,
    new_n19808_, new_n19809_, new_n19810_, new_n19811_, new_n19812_,
    new_n19813_, new_n19814_, new_n19815_, new_n19816_, new_n19817_,
    new_n19818_, new_n19819_, new_n19820_, new_n19821_, new_n19822_,
    new_n19823_, new_n19824_, new_n19825_, new_n19826_, new_n19827_,
    new_n19828_, new_n19829_, new_n19830_, new_n19831_, new_n19832_,
    new_n19833_, new_n19834_, new_n19835_, new_n19836_, new_n19837_,
    new_n19838_, new_n19839_, new_n19840_, new_n19841_, new_n19842_,
    new_n19843_, new_n19844_, new_n19845_, new_n19846_, new_n19847_,
    new_n19848_, new_n19849_, new_n19850_, new_n19851_, new_n19852_,
    new_n19853_, new_n19854_, new_n19855_, new_n19856_, new_n19857_,
    new_n19858_, new_n19859_, new_n19860_, new_n19861_, new_n19862_,
    new_n19863_, new_n19864_, new_n19865_, new_n19866_, new_n19867_,
    new_n19868_, new_n19869_, new_n19870_, new_n19871_, new_n19872_,
    new_n19873_, new_n19874_, new_n19875_, new_n19876_, new_n19877_,
    new_n19878_, new_n19879_, new_n19880_, new_n19881_, new_n19882_,
    new_n19883_, new_n19884_, new_n19885_, new_n19886_, new_n19887_,
    new_n19888_, new_n19889_, new_n19890_, new_n19891_, new_n19892_,
    new_n19893_, new_n19894_, new_n19895_, new_n19896_, new_n19897_,
    new_n19898_, new_n19899_, new_n19900_, new_n19901_, new_n19902_,
    new_n19903_, new_n19904_, new_n19905_, new_n19906_, new_n19907_,
    new_n19908_, new_n19909_, new_n19910_, new_n19911_, new_n19912_,
    new_n19913_, new_n19914_, new_n19916_, new_n19917_, new_n19918_,
    new_n19919_, new_n19920_, new_n19921_, new_n19922_, new_n19923_,
    new_n19924_, new_n19925_, new_n19926_, new_n19927_, new_n19928_,
    new_n19929_, new_n19930_, new_n19931_, new_n19932_, new_n19933_,
    new_n19934_, new_n19935_, new_n19936_, new_n19937_, new_n19938_,
    new_n19939_, new_n19940_, new_n19941_, new_n19942_, new_n19943_,
    new_n19944_, new_n19945_, new_n19946_, new_n19947_, new_n19948_,
    new_n19949_, new_n19950_, new_n19951_, new_n19952_, new_n19953_,
    new_n19954_, new_n19955_, new_n19956_, new_n19957_, new_n19958_,
    new_n19959_, new_n19960_, new_n19961_, new_n19962_, new_n19963_,
    new_n19964_, new_n19965_, new_n19966_, new_n19967_, new_n19968_,
    new_n19969_, new_n19970_, new_n19971_, new_n19972_, new_n19973_,
    new_n19974_, new_n19975_, new_n19976_, new_n19977_, new_n19978_,
    new_n19979_, new_n19980_, new_n19981_, new_n19982_, new_n19983_,
    new_n19984_, new_n19985_, new_n19986_, new_n19987_, new_n19988_,
    new_n19989_, new_n19990_, new_n19991_, new_n19992_, new_n19993_,
    new_n19994_, new_n19995_, new_n19996_, new_n19997_, new_n19998_,
    new_n19999_, new_n20000_, new_n20001_, new_n20002_, new_n20003_,
    new_n20004_, new_n20005_, new_n20006_, new_n20007_, new_n20008_,
    new_n20009_, new_n20010_, new_n20011_, new_n20012_, new_n20014_,
    new_n20015_, new_n20016_, new_n20017_, new_n20018_, new_n20019_,
    new_n20020_, new_n20021_, new_n20022_, new_n20023_, new_n20024_,
    new_n20025_, new_n20026_, new_n20027_, new_n20028_, new_n20029_,
    new_n20030_, new_n20031_, new_n20032_, new_n20033_, new_n20034_,
    new_n20035_, new_n20036_, new_n20037_, new_n20038_, new_n20039_,
    new_n20040_, new_n20041_, new_n20042_, new_n20043_, new_n20044_,
    new_n20045_, new_n20046_, new_n20047_, new_n20048_, new_n20049_,
    new_n20050_, new_n20051_, new_n20052_, new_n20053_, new_n20054_,
    new_n20055_, new_n20056_, new_n20057_, new_n20058_, new_n20059_,
    new_n20060_, new_n20061_, new_n20062_, new_n20063_, new_n20064_,
    new_n20065_, new_n20066_, new_n20067_, new_n20068_, new_n20069_,
    new_n20070_, new_n20071_, new_n20072_, new_n20073_, new_n20074_,
    new_n20075_, new_n20076_, new_n20077_, new_n20078_, new_n20079_,
    new_n20080_, new_n20081_, new_n20082_, new_n20083_, new_n20084_,
    new_n20085_, new_n20086_, new_n20087_, new_n20088_, new_n20089_,
    new_n20090_, new_n20091_, new_n20092_, new_n20093_, new_n20094_,
    new_n20095_, new_n20096_, new_n20097_, new_n20098_, new_n20099_,
    new_n20100_, new_n20101_, new_n20102_, new_n20103_, new_n20104_,
    new_n20105_, new_n20106_, new_n20107_, new_n20109_, new_n20110_,
    new_n20111_, new_n20112_, new_n20113_, new_n20114_, new_n20115_,
    new_n20116_, new_n20117_, new_n20118_, new_n20119_, new_n20120_,
    new_n20121_, new_n20122_, new_n20123_, new_n20124_, new_n20125_,
    new_n20126_, new_n20127_, new_n20128_, new_n20129_, new_n20130_,
    new_n20131_, new_n20132_, new_n20133_, new_n20134_, new_n20135_,
    new_n20136_, new_n20137_, new_n20138_, new_n20139_, new_n20140_,
    new_n20141_, new_n20142_, new_n20143_, new_n20144_, new_n20145_,
    new_n20146_, new_n20147_, new_n20148_, new_n20149_, new_n20150_,
    new_n20151_, new_n20152_, new_n20153_, new_n20154_, new_n20155_,
    new_n20156_, new_n20157_, new_n20158_, new_n20159_, new_n20160_,
    new_n20161_, new_n20162_, new_n20163_, new_n20164_, new_n20165_,
    new_n20166_, new_n20167_, new_n20168_, new_n20169_, new_n20170_,
    new_n20171_, new_n20172_, new_n20173_, new_n20174_, new_n20175_,
    new_n20176_, new_n20177_, new_n20178_, new_n20179_, new_n20180_,
    new_n20181_, new_n20182_, new_n20183_, new_n20184_, new_n20185_,
    new_n20186_, new_n20187_, new_n20188_, new_n20189_, new_n20190_,
    new_n20191_, new_n20192_, new_n20193_, new_n20194_, new_n20195_,
    new_n20196_, new_n20197_, new_n20198_, new_n20199_, new_n20200_,
    new_n20201_, new_n20203_, new_n20204_, new_n20205_, new_n20206_,
    new_n20207_, new_n20208_, new_n20209_, new_n20210_, new_n20211_,
    new_n20212_, new_n20213_, new_n20214_, new_n20215_, new_n20216_,
    new_n20217_, new_n20218_, new_n20219_, new_n20220_, new_n20221_,
    new_n20222_, new_n20223_, new_n20224_, new_n20225_, new_n20226_,
    new_n20227_, new_n20228_, new_n20229_, new_n20230_, new_n20231_,
    new_n20232_, new_n20233_, new_n20234_, new_n20235_, new_n20236_,
    new_n20237_, new_n20238_, new_n20239_, new_n20240_, new_n20241_,
    new_n20242_, new_n20243_, new_n20244_, new_n20245_, new_n20246_,
    new_n20247_, new_n20248_, new_n20249_, new_n20250_, new_n20251_,
    new_n20252_, new_n20253_, new_n20254_, new_n20255_, new_n20256_,
    new_n20257_, new_n20258_, new_n20259_, new_n20260_, new_n20261_,
    new_n20262_, new_n20263_, new_n20264_, new_n20265_, new_n20266_,
    new_n20267_, new_n20268_, new_n20269_, new_n20270_, new_n20271_,
    new_n20272_, new_n20273_, new_n20274_, new_n20275_, new_n20276_,
    new_n20277_, new_n20278_, new_n20279_, new_n20280_, new_n20281_,
    new_n20282_, new_n20283_, new_n20284_, new_n20285_, new_n20286_,
    new_n20287_, new_n20288_, new_n20289_, new_n20290_, new_n20291_,
    new_n20292_, new_n20293_, new_n20294_, new_n20295_, new_n20297_,
    new_n20298_, new_n20299_, new_n20300_, new_n20301_, new_n20302_,
    new_n20303_, new_n20304_, new_n20305_, new_n20306_, new_n20307_,
    new_n20308_, new_n20309_, new_n20310_, new_n20311_, new_n20312_,
    new_n20313_, new_n20314_, new_n20315_, new_n20316_, new_n20317_,
    new_n20318_, new_n20319_, new_n20320_, new_n20321_, new_n20322_,
    new_n20323_, new_n20324_, new_n20325_, new_n20326_, new_n20327_,
    new_n20328_, new_n20329_, new_n20330_, new_n20331_, new_n20332_,
    new_n20333_, new_n20334_, new_n20335_, new_n20336_, new_n20337_,
    new_n20338_, new_n20339_, new_n20340_, new_n20341_, new_n20342_,
    new_n20343_, new_n20344_, new_n20345_, new_n20346_, new_n20347_,
    new_n20348_, new_n20349_, new_n20350_, new_n20351_, new_n20352_,
    new_n20353_, new_n20354_, new_n20355_, new_n20356_, new_n20357_,
    new_n20358_, new_n20359_, new_n20360_, new_n20361_, new_n20362_,
    new_n20363_, new_n20364_, new_n20365_, new_n20366_, new_n20367_,
    new_n20368_, new_n20369_, new_n20370_, new_n20371_, new_n20372_,
    new_n20373_, new_n20374_, new_n20375_, new_n20377_, new_n20378_,
    new_n20379_, new_n20380_, new_n20381_, new_n20382_, new_n20383_,
    new_n20384_, new_n20385_, new_n20386_, new_n20387_, new_n20388_,
    new_n20389_, new_n20390_, new_n20391_, new_n20392_, new_n20393_,
    new_n20394_, new_n20395_, new_n20396_, new_n20397_, new_n20398_,
    new_n20399_, new_n20400_, new_n20401_, new_n20402_, new_n20403_,
    new_n20404_, new_n20405_, new_n20406_, new_n20407_, new_n20408_,
    new_n20409_, new_n20410_, new_n20411_, new_n20412_, new_n20413_,
    new_n20414_, new_n20415_, new_n20416_, new_n20417_, new_n20418_,
    new_n20419_, new_n20420_, new_n20421_, new_n20422_, new_n20423_,
    new_n20424_, new_n20425_, new_n20426_, new_n20427_, new_n20428_,
    new_n20429_, new_n20430_, new_n20431_, new_n20432_, new_n20433_,
    new_n20434_, new_n20435_, new_n20436_, new_n20437_, new_n20438_,
    new_n20439_, new_n20440_, new_n20441_, new_n20442_, new_n20443_,
    new_n20444_, new_n20445_, new_n20446_, new_n20447_, new_n20448_,
    new_n20449_, new_n20450_, new_n20451_, new_n20452_, new_n20453_,
    new_n20454_, new_n20455_, new_n20456_, new_n20457_, new_n20458_,
    new_n20459_, new_n20460_, new_n20461_, new_n20462_, new_n20464_,
    new_n20465_, new_n20466_, new_n20467_, new_n20468_, new_n20469_,
    new_n20470_, new_n20471_, new_n20472_, new_n20473_, new_n20474_,
    new_n20475_, new_n20476_, new_n20477_, new_n20478_, new_n20479_,
    new_n20480_, new_n20481_, new_n20482_, new_n20483_, new_n20484_,
    new_n20485_, new_n20486_, new_n20487_, new_n20488_, new_n20489_,
    new_n20490_, new_n20491_, new_n20492_, new_n20493_, new_n20494_,
    new_n20495_, new_n20496_, new_n20497_, new_n20498_, new_n20499_,
    new_n20500_, new_n20501_, new_n20502_, new_n20503_, new_n20504_,
    new_n20505_, new_n20506_, new_n20507_, new_n20508_, new_n20509_,
    new_n20510_, new_n20511_, new_n20512_, new_n20513_, new_n20514_,
    new_n20515_, new_n20516_, new_n20517_, new_n20518_, new_n20519_,
    new_n20520_, new_n20521_, new_n20522_, new_n20523_, new_n20524_,
    new_n20525_, new_n20526_, new_n20527_, new_n20528_, new_n20529_,
    new_n20530_, new_n20531_, new_n20532_, new_n20533_, new_n20534_,
    new_n20536_, new_n20537_, new_n20538_, new_n20539_, new_n20540_,
    new_n20541_, new_n20542_, new_n20543_, new_n20544_, new_n20545_,
    new_n20546_, new_n20547_, new_n20548_, new_n20549_, new_n20550_,
    new_n20551_, new_n20552_, new_n20553_, new_n20554_, new_n20555_,
    new_n20556_, new_n20557_, new_n20558_, new_n20559_, new_n20560_,
    new_n20561_, new_n20562_, new_n20563_, new_n20564_, new_n20565_,
    new_n20566_, new_n20567_, new_n20568_, new_n20569_, new_n20570_,
    new_n20571_, new_n20572_, new_n20573_, new_n20574_, new_n20575_,
    new_n20576_, new_n20577_, new_n20578_, new_n20579_, new_n20580_,
    new_n20581_, new_n20582_, new_n20583_, new_n20584_, new_n20585_,
    new_n20586_, new_n20587_, new_n20588_, new_n20589_, new_n20590_,
    new_n20591_, new_n20592_, new_n20593_, new_n20594_, new_n20595_,
    new_n20596_, new_n20597_, new_n20598_, new_n20599_, new_n20600_,
    new_n20601_, new_n20602_, new_n20604_, new_n20605_, new_n20606_,
    new_n20607_, new_n20608_, new_n20609_, new_n20610_, new_n20611_,
    new_n20612_, new_n20613_, new_n20614_, new_n20615_, new_n20616_,
    new_n20617_, new_n20618_, new_n20619_, new_n20620_, new_n20621_,
    new_n20622_, new_n20623_, new_n20624_, new_n20625_, new_n20626_,
    new_n20627_, new_n20628_, new_n20629_, new_n20630_, new_n20631_,
    new_n20632_, new_n20633_, new_n20634_, new_n20635_, new_n20636_,
    new_n20637_, new_n20638_, new_n20639_, new_n20640_, new_n20641_,
    new_n20642_, new_n20643_, new_n20644_, new_n20645_, new_n20646_,
    new_n20647_, new_n20648_, new_n20649_, new_n20650_, new_n20651_,
    new_n20652_, new_n20653_, new_n20654_, new_n20655_, new_n20656_,
    new_n20657_, new_n20658_, new_n20659_, new_n20660_, new_n20661_,
    new_n20662_, new_n20663_, new_n20664_, new_n20665_, new_n20666_,
    new_n20667_, new_n20668_, new_n20669_, new_n20670_, new_n20671_,
    new_n20672_, new_n20673_, new_n20674_, new_n20675_, new_n20676_,
    new_n20677_, new_n20678_, new_n20680_, new_n20681_, new_n20682_,
    new_n20683_, new_n20684_, new_n20685_, new_n20686_, new_n20687_,
    new_n20688_, new_n20689_, new_n20690_, new_n20691_, new_n20692_,
    new_n20693_, new_n20694_, new_n20695_, new_n20696_, new_n20697_,
    new_n20698_, new_n20699_, new_n20700_, new_n20701_, new_n20702_,
    new_n20703_, new_n20704_, new_n20705_, new_n20706_, new_n20707_,
    new_n20708_, new_n20709_, new_n20710_, new_n20711_, new_n20712_,
    new_n20713_, new_n20714_, new_n20715_, new_n20716_, new_n20717_,
    new_n20718_, new_n20719_, new_n20720_, new_n20721_, new_n20722_,
    new_n20723_, new_n20724_, new_n20725_, new_n20726_, new_n20727_,
    new_n20728_, new_n20729_, new_n20730_, new_n20731_, new_n20732_,
    new_n20733_, new_n20734_, new_n20735_, new_n20736_, new_n20737_,
    new_n20738_, new_n20739_, new_n20740_, new_n20741_, new_n20742_,
    new_n20743_, new_n20744_, new_n20745_, new_n20747_, new_n20748_,
    new_n20749_, new_n20750_, new_n20751_, new_n20752_, new_n20753_,
    new_n20754_, new_n20755_, new_n20756_, new_n20757_, new_n20758_,
    new_n20759_, new_n20760_, new_n20761_, new_n20762_, new_n20763_,
    new_n20764_, new_n20765_, new_n20766_, new_n20767_, new_n20768_,
    new_n20769_, new_n20770_, new_n20771_, new_n20772_, new_n20773_,
    new_n20774_, new_n20775_, new_n20776_, new_n20777_, new_n20778_,
    new_n20779_, new_n20780_, new_n20781_, new_n20782_, new_n20783_,
    new_n20784_, new_n20785_, new_n20786_, new_n20787_, new_n20788_,
    new_n20789_, new_n20790_, new_n20791_, new_n20792_, new_n20793_,
    new_n20794_, new_n20795_, new_n20796_, new_n20797_, new_n20798_,
    new_n20799_, new_n20800_, new_n20801_, new_n20803_, new_n20804_,
    new_n20805_, new_n20806_, new_n20807_, new_n20808_, new_n20809_,
    new_n20810_, new_n20811_, new_n20812_, new_n20813_, new_n20814_,
    new_n20815_, new_n20816_, new_n20817_, new_n20818_, new_n20819_,
    new_n20820_, new_n20821_, new_n20822_, new_n20823_, new_n20824_,
    new_n20825_, new_n20826_, new_n20827_, new_n20828_, new_n20829_,
    new_n20830_, new_n20831_, new_n20832_, new_n20833_, new_n20834_,
    new_n20835_, new_n20836_, new_n20837_, new_n20838_, new_n20839_,
    new_n20840_, new_n20841_, new_n20842_, new_n20843_, new_n20844_,
    new_n20845_, new_n20846_, new_n20847_, new_n20848_, new_n20849_,
    new_n20850_, new_n20851_, new_n20852_, new_n20853_, new_n20854_,
    new_n20855_, new_n20856_, new_n20857_, new_n20858_, new_n20859_,
    new_n20860_, new_n20861_, new_n20862_, new_n20863_, new_n20864_,
    new_n20865_, new_n20866_, new_n20867_, new_n20868_, new_n20869_,
    new_n20870_, new_n20871_, new_n20872_, new_n20873_, new_n20875_,
    new_n20876_, new_n20877_, new_n20878_, new_n20879_, new_n20880_,
    new_n20881_, new_n20882_, new_n20883_, new_n20884_, new_n20885_,
    new_n20886_, new_n20887_, new_n20888_, new_n20889_, new_n20890_,
    new_n20891_, new_n20892_, new_n20893_, new_n20894_, new_n20895_,
    new_n20896_, new_n20897_, new_n20898_, new_n20899_, new_n20900_,
    new_n20901_, new_n20902_, new_n20903_, new_n20904_, new_n20905_,
    new_n20906_, new_n20907_, new_n20908_, new_n20909_, new_n20910_,
    new_n20911_, new_n20912_, new_n20913_, new_n20914_, new_n20915_,
    new_n20916_, new_n20917_, new_n20918_, new_n20919_, new_n20920_,
    new_n20921_, new_n20923_, new_n20924_, new_n20925_, new_n20926_,
    new_n20927_, new_n20928_, new_n20929_, new_n20930_, new_n20931_,
    new_n20932_, new_n20933_, new_n20934_, new_n20935_, new_n20936_,
    new_n20937_, new_n20938_, new_n20939_, new_n20940_, new_n20941_,
    new_n20942_, new_n20943_, new_n20944_, new_n20945_, new_n20946_,
    new_n20947_, new_n20948_, new_n20949_, new_n20950_, new_n20951_,
    new_n20952_, new_n20953_, new_n20954_, new_n20955_, new_n20956_,
    new_n20957_, new_n20958_, new_n20959_, new_n20960_, new_n20961_,
    new_n20962_, new_n20963_, new_n20964_, new_n20965_, new_n20966_,
    new_n20967_, new_n20968_, new_n20970_, new_n20971_, new_n20972_,
    new_n20973_, new_n20974_, new_n20975_, new_n20976_, new_n20977_,
    new_n20978_, new_n20979_, new_n20980_, new_n20981_, new_n20982_,
    new_n20983_, new_n20984_, new_n20985_, new_n20986_, new_n20987_,
    new_n20988_, new_n20989_, new_n20990_, new_n20991_, new_n20992_,
    new_n20993_, new_n20994_, new_n20995_, new_n20996_, new_n20997_,
    new_n20998_, new_n20999_, new_n21000_, new_n21001_, new_n21002_,
    new_n21003_, new_n21004_, new_n21005_, new_n21006_, new_n21007_,
    new_n21008_, new_n21009_, new_n21010_, new_n21011_, new_n21012_,
    new_n21013_, new_n21014_, new_n21015_, new_n21016_, new_n21017_,
    new_n21018_, new_n21020_, new_n21021_, new_n21022_, new_n21023_,
    new_n21024_, new_n21025_, new_n21026_, new_n21027_, new_n21028_,
    new_n21029_, new_n21030_, new_n21031_, new_n21032_, new_n21033_,
    new_n21034_, new_n21035_, new_n21036_, new_n21037_, new_n21038_,
    new_n21039_, new_n21040_, new_n21041_, new_n21042_, new_n21043_,
    new_n21044_, new_n21045_, new_n21046_, new_n21047_, new_n21048_,
    new_n21049_, new_n21050_, new_n21051_, new_n21052_, new_n21053_,
    new_n21054_, new_n21055_, new_n21056_, new_n21057_, new_n21058_,
    new_n21059_, new_n21060_, new_n21061_, new_n21062_, new_n21063_,
    new_n21065_, new_n21066_, new_n21067_, new_n21068_, new_n21069_,
    new_n21070_, new_n21071_, new_n21072_, new_n21073_, new_n21074_,
    new_n21075_, new_n21076_, new_n21077_, new_n21078_, new_n21079_,
    new_n21080_, new_n21081_, new_n21082_, new_n21083_, new_n21084_,
    new_n21085_, new_n21086_, new_n21087_, new_n21088_, new_n21089_,
    new_n21090_, new_n21091_, new_n21092_, new_n21093_, new_n21094_,
    new_n21095_, new_n21096_, new_n21097_, new_n21098_, new_n21099_,
    new_n21100_, new_n21101_, new_n21103_, new_n21104_, new_n21105_,
    new_n21106_, new_n21107_, new_n21108_, new_n21109_, new_n21110_,
    new_n21111_, new_n21112_, new_n21113_, new_n21114_, new_n21115_,
    new_n21116_, new_n21117_, new_n21118_, new_n21119_, new_n21120_,
    new_n21121_, new_n21122_, new_n21123_, new_n21124_, new_n21125_,
    new_n21126_, new_n21127_, new_n21128_, new_n21129_, new_n21130_,
    new_n21131_, new_n21132_, new_n21133_, new_n21134_, new_n21135_,
    new_n21136_, new_n21137_, new_n21138_, new_n21139_, new_n21140_,
    new_n21141_, new_n21143_, new_n21144_, new_n21145_, new_n21146_,
    new_n21147_, new_n21148_, new_n21149_, new_n21150_, new_n21151_,
    new_n21152_, new_n21153_, new_n21154_, new_n21155_, new_n21156_,
    new_n21157_, new_n21158_, new_n21159_, new_n21160_, new_n21161_,
    new_n21162_, new_n21163_, new_n21164_, new_n21165_, new_n21166_,
    new_n21167_, new_n21168_, new_n21169_, new_n21170_, new_n21171_,
    new_n21172_, new_n21173_, new_n21174_, new_n21175_, new_n21176_,
    new_n21177_, new_n21179_, new_n21180_, new_n21181_, new_n21182_,
    new_n21183_, new_n21184_, new_n21185_, new_n21186_, new_n21187_,
    new_n21188_, new_n21189_, new_n21190_, new_n21191_, new_n21192_,
    new_n21193_, new_n21194_, new_n21195_, new_n21196_, new_n21197_,
    new_n21198_, new_n21199_, new_n21200_, new_n21201_, new_n21202_,
    new_n21203_, new_n21205_, new_n21206_, new_n21207_, new_n21208_,
    new_n21209_, new_n21210_, new_n21211_, new_n21212_, new_n21213_,
    new_n21214_, new_n21215_, new_n21216_, new_n21217_, new_n21218_,
    new_n21219_, new_n21220_, new_n21221_, new_n21222_, new_n21223_,
    new_n21224_, new_n21225_, new_n21226_, new_n21227_, new_n21228_,
    new_n21229_, new_n21230_, new_n21231_, new_n21232_, new_n21233_,
    new_n21235_, new_n21236_, new_n21237_, new_n21238_, new_n21239_,
    new_n21240_, new_n21241_, new_n21242_, new_n21243_, new_n21244_,
    new_n21245_, new_n21246_, new_n21247_, new_n21248_, new_n21249_,
    new_n21250_, new_n21251_, new_n21252_, new_n21253_, new_n21254_,
    new_n21255_, new_n21256_, new_n21258_, new_n21259_, new_n21260_,
    new_n21261_, new_n21262_, new_n21263_, new_n21264_, new_n21265_,
    new_n21266_, new_n21267_, new_n21268_, new_n21269_, new_n21270_,
    new_n21271_, new_n21272_, new_n21273_, new_n21274_, new_n21276_,
    new_n21277_, new_n21278_, new_n21279_, new_n21280_, new_n21281_,
    new_n21282_, new_n21283_, new_n21284_, new_n21285_, new_n21286_,
    new_n21287_, new_n21288_, new_n21289_, new_n21290_, new_n21291_,
    new_n21292_, new_n21293_, new_n21294_, new_n21295_, new_n21296_,
    new_n21298_, new_n21299_, new_n21300_, new_n21301_, new_n21302_,
    new_n21303_, new_n21304_, new_n21305_, new_n21306_, new_n21307_,
    new_n21308_;
  INV_X1     g00000(.I(\a[0] ), .ZN(new_n257_));
  INV_X1     g00001(.I(\b[0] ), .ZN(new_n258_));
  NOR2_X1    g00002(.A1(new_n257_), .A2(new_n258_), .ZN(\f[0] ));
  INV_X1     g00003(.I(\a[1] ), .ZN(new_n260_));
  NOR2_X1    g00004(.A1(new_n260_), .A2(\a[0] ), .ZN(new_n261_));
  INV_X1     g00005(.I(new_n261_), .ZN(new_n262_));
  XOR2_X1    g00006(.A1(\b[0] ), .A2(\b[1] ), .Z(new_n263_));
  XNOR2_X1   g00007(.A1(\a[1] ), .A2(\a[2] ), .ZN(new_n264_));
  NOR2_X1    g00008(.A1(new_n264_), .A2(new_n257_), .ZN(new_n265_));
  XOR2_X1    g00009(.A1(\a[1] ), .A2(\a[2] ), .Z(new_n266_));
  NOR2_X1    g00010(.A1(new_n266_), .A2(new_n257_), .ZN(new_n267_));
  AOI22_X1   g00011(.A1(new_n265_), .A2(new_n263_), .B1(new_n267_), .B2(\b[1] ), .ZN(new_n268_));
  OAI21_X1   g00012(.A1(new_n258_), .A2(new_n262_), .B(new_n268_), .ZN(new_n269_));
  INV_X1     g00013(.I(\a[2] ), .ZN(new_n270_));
  NOR3_X1    g00014(.A1(new_n257_), .A2(new_n270_), .A3(new_n258_), .ZN(new_n271_));
  XOR2_X1    g00015(.A1(new_n269_), .A2(new_n271_), .Z(\f[1] ));
  NOR2_X1    g00016(.A1(new_n269_), .A2(\f[0] ), .ZN(new_n273_));
  NAND2_X1   g00017(.A1(new_n273_), .A2(\a[2] ), .ZN(new_n274_));
  INV_X1     g00018(.I(\b[1] ), .ZN(new_n275_));
  INV_X1     g00019(.I(\b[2] ), .ZN(new_n276_));
  INV_X1     g00020(.I(new_n267_), .ZN(new_n277_));
  OAI22_X1   g00021(.A1(new_n277_), .A2(new_n276_), .B1(new_n275_), .B2(new_n262_), .ZN(new_n278_));
  INV_X1     g00022(.I(new_n265_), .ZN(new_n279_));
  AOI21_X1   g00023(.A1(new_n258_), .A2(\b[1] ), .B(new_n276_), .ZN(new_n280_));
  NOR3_X1    g00024(.A1(new_n275_), .A2(\b[0] ), .A3(\b[2] ), .ZN(new_n281_));
  NOR2_X1    g00025(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NOR3_X1    g00026(.A1(new_n270_), .A2(\a[0] ), .A3(\a[1] ), .ZN(new_n283_));
  INV_X1     g00027(.I(new_n283_), .ZN(new_n284_));
  OAI22_X1   g00028(.A1(new_n279_), .A2(new_n282_), .B1(new_n258_), .B2(new_n284_), .ZN(new_n285_));
  NOR2_X1    g00029(.A1(new_n285_), .A2(new_n278_), .ZN(new_n286_));
  XOR2_X1    g00030(.A1(new_n286_), .A2(\a[2] ), .Z(new_n287_));
  XOR2_X1    g00031(.A1(new_n287_), .A2(new_n274_), .Z(\f[2] ));
  NAND3_X1   g00032(.A1(new_n273_), .A2(\a[2] ), .A3(new_n286_), .ZN(new_n289_));
  INV_X1     g00033(.I(\b[3] ), .ZN(new_n290_));
  OAI22_X1   g00034(.A1(new_n277_), .A2(new_n290_), .B1(new_n275_), .B2(new_n284_), .ZN(new_n291_));
  AOI21_X1   g00035(.A1(\b[2] ), .A2(new_n261_), .B(new_n291_), .ZN(new_n292_));
  NAND3_X1   g00036(.A1(new_n276_), .A2(\b[0] ), .A3(\b[1] ), .ZN(new_n293_));
  NAND2_X1   g00037(.A1(new_n275_), .A2(\b[2] ), .ZN(new_n294_));
  AOI21_X1   g00038(.A1(new_n293_), .A2(new_n294_), .B(new_n290_), .ZN(new_n295_));
  NOR3_X1    g00039(.A1(new_n258_), .A2(new_n275_), .A3(\b[2] ), .ZN(new_n296_));
  NOR2_X1    g00040(.A1(new_n276_), .A2(\b[1] ), .ZN(new_n297_));
  NOR3_X1    g00041(.A1(new_n296_), .A2(\b[3] ), .A3(new_n297_), .ZN(new_n298_));
  NOR2_X1    g00042(.A1(new_n298_), .A2(new_n295_), .ZN(new_n299_));
  NAND2_X1   g00043(.A1(new_n299_), .A2(new_n265_), .ZN(new_n300_));
  AOI21_X1   g00044(.A1(new_n292_), .A2(new_n300_), .B(new_n270_), .ZN(new_n301_));
  NAND3_X1   g00045(.A1(new_n292_), .A2(new_n270_), .A3(new_n300_), .ZN(new_n302_));
  INV_X1     g00046(.I(new_n302_), .ZN(new_n303_));
  XNOR2_X1   g00047(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n304_));
  NOR2_X1    g00048(.A1(new_n304_), .A2(new_n258_), .ZN(new_n305_));
  INV_X1     g00049(.I(new_n305_), .ZN(new_n306_));
  OAI21_X1   g00050(.A1(new_n303_), .A2(new_n301_), .B(new_n306_), .ZN(new_n307_));
  INV_X1     g00051(.I(new_n301_), .ZN(new_n308_));
  NAND3_X1   g00052(.A1(new_n308_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n309_));
  NAND2_X1   g00053(.A1(new_n309_), .A2(new_n307_), .ZN(new_n310_));
  XOR2_X1    g00054(.A1(new_n310_), .A2(new_n289_), .Z(\f[3] ));
  INV_X1     g00055(.I(\a[5] ), .ZN(new_n312_));
  XNOR2_X1   g00056(.A1(\b[0] ), .A2(\b[1] ), .ZN(new_n313_));
  XOR2_X1    g00057(.A1(\a[2] ), .A2(\a[3] ), .Z(new_n314_));
  NOR2_X1    g00058(.A1(new_n312_), .A2(\a[4] ), .ZN(new_n315_));
  INV_X1     g00059(.I(\a[4] ), .ZN(new_n316_));
  NOR2_X1    g00060(.A1(new_n316_), .A2(\a[5] ), .ZN(new_n317_));
  OAI21_X1   g00061(.A1(new_n315_), .A2(new_n317_), .B(new_n314_), .ZN(new_n318_));
  NOR2_X1    g00062(.A1(new_n318_), .A2(new_n313_), .ZN(new_n319_));
  XNOR2_X1   g00063(.A1(\a[4] ), .A2(\a[5] ), .ZN(new_n320_));
  NAND2_X1   g00064(.A1(new_n320_), .A2(new_n314_), .ZN(new_n321_));
  NOR2_X1    g00065(.A1(new_n321_), .A2(new_n275_), .ZN(new_n322_));
  NOR3_X1    g00066(.A1(new_n316_), .A2(\a[2] ), .A3(\a[3] ), .ZN(new_n323_));
  AND3_X2    g00067(.A1(new_n316_), .A2(\a[2] ), .A3(\a[3] ), .Z(new_n324_));
  NOR2_X1    g00068(.A1(new_n324_), .A2(new_n323_), .ZN(new_n325_));
  NOR2_X1    g00069(.A1(new_n325_), .A2(new_n258_), .ZN(new_n326_));
  NOR3_X1    g00070(.A1(new_n319_), .A2(new_n322_), .A3(new_n326_), .ZN(new_n327_));
  NOR2_X1    g00071(.A1(new_n327_), .A2(new_n312_), .ZN(new_n328_));
  NOR2_X1    g00072(.A1(new_n315_), .A2(new_n317_), .ZN(new_n329_));
  NOR2_X1    g00073(.A1(new_n329_), .A2(new_n304_), .ZN(new_n330_));
  NAND2_X1   g00074(.A1(new_n330_), .A2(new_n263_), .ZN(new_n331_));
  XOR2_X1    g00075(.A1(\a[4] ), .A2(\a[5] ), .Z(new_n332_));
  NOR2_X1    g00076(.A1(new_n304_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1   g00077(.A1(new_n333_), .A2(\b[1] ), .ZN(new_n334_));
  INV_X1     g00078(.I(new_n326_), .ZN(new_n335_));
  NAND3_X1   g00079(.A1(new_n335_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n336_));
  NOR2_X1    g00080(.A1(new_n336_), .A2(\a[5] ), .ZN(new_n337_));
  NOR2_X1    g00081(.A1(new_n284_), .A2(new_n276_), .ZN(new_n338_));
  INV_X1     g00082(.I(\b[4] ), .ZN(new_n339_));
  OAI22_X1   g00083(.A1(new_n277_), .A2(new_n339_), .B1(new_n290_), .B2(new_n262_), .ZN(new_n340_));
  NAND2_X1   g00084(.A1(\b[3] ), .A2(\b[4] ), .ZN(new_n341_));
  NOR2_X1    g00085(.A1(\b[3] ), .A2(\b[4] ), .ZN(new_n342_));
  INV_X1     g00086(.I(new_n342_), .ZN(new_n343_));
  OAI21_X1   g00087(.A1(\b[1] ), .A2(\b[3] ), .B(\b[2] ), .ZN(new_n344_));
  NAND3_X1   g00088(.A1(\b[0] ), .A2(\b[1] ), .A3(\b[3] ), .ZN(new_n345_));
  AOI22_X1   g00089(.A1(new_n343_), .A2(new_n341_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1     g00090(.I(new_n341_), .ZN(new_n347_));
  NOR2_X1    g00091(.A1(\b[1] ), .A2(\b[3] ), .ZN(new_n348_));
  NOR2_X1    g00092(.A1(new_n348_), .A2(new_n276_), .ZN(new_n349_));
  AND3_X2    g00093(.A1(\b[0] ), .A2(\b[1] ), .A3(\b[3] ), .Z(new_n350_));
  NOR4_X1    g00094(.A1(new_n349_), .A2(new_n350_), .A3(new_n347_), .A4(new_n342_), .ZN(new_n351_));
  NOR2_X1    g00095(.A1(new_n351_), .A2(new_n346_), .ZN(new_n352_));
  NOR2_X1    g00096(.A1(new_n352_), .A2(new_n279_), .ZN(new_n353_));
  NOR3_X1    g00097(.A1(new_n340_), .A2(new_n353_), .A3(new_n338_), .ZN(new_n354_));
  INV_X1     g00098(.I(new_n354_), .ZN(new_n355_));
  NOR3_X1    g00099(.A1(new_n355_), .A2(new_n337_), .A3(new_n328_), .ZN(new_n356_));
  INV_X1     g00100(.I(new_n356_), .ZN(new_n357_));
  OAI21_X1   g00101(.A1(new_n328_), .A2(new_n337_), .B(new_n355_), .ZN(new_n358_));
  NOR2_X1    g00102(.A1(new_n305_), .A2(new_n312_), .ZN(new_n359_));
  XOR2_X1    g00103(.A1(new_n359_), .A2(new_n270_), .Z(new_n360_));
  AOI21_X1   g00104(.A1(new_n357_), .A2(new_n358_), .B(new_n360_), .ZN(new_n361_));
  NOR2_X1    g00105(.A1(new_n337_), .A2(new_n328_), .ZN(new_n362_));
  NOR2_X1    g00106(.A1(new_n362_), .A2(new_n354_), .ZN(new_n363_));
  INV_X1     g00107(.I(new_n360_), .ZN(new_n364_));
  NOR3_X1    g00108(.A1(new_n363_), .A2(new_n356_), .A3(new_n364_), .ZN(new_n365_));
  NOR2_X1    g00109(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  AOI21_X1   g00110(.A1(new_n308_), .A2(new_n302_), .B(new_n305_), .ZN(new_n367_));
  AOI21_X1   g00111(.A1(new_n289_), .A2(new_n309_), .B(new_n367_), .ZN(new_n368_));
  XOR2_X1    g00112(.A1(new_n366_), .A2(new_n368_), .Z(\f[4] ));
  NAND2_X1   g00113(.A1(new_n261_), .A2(\b[4] ), .ZN(new_n370_));
  AOI22_X1   g00114(.A1(new_n267_), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n283_), .ZN(new_n371_));
  NAND2_X1   g00115(.A1(new_n371_), .A2(new_n370_), .ZN(new_n372_));
  NAND2_X1   g00116(.A1(new_n344_), .A2(new_n345_), .ZN(new_n373_));
  AOI21_X1   g00117(.A1(new_n373_), .A2(\b[4] ), .B(new_n290_), .ZN(new_n374_));
  NOR2_X1    g00118(.A1(new_n373_), .A2(\b[4] ), .ZN(new_n375_));
  NOR3_X1    g00119(.A1(new_n349_), .A2(new_n350_), .A3(\b[5] ), .ZN(new_n376_));
  INV_X1     g00120(.I(\b[5] ), .ZN(new_n377_));
  AOI21_X1   g00121(.A1(new_n344_), .A2(new_n345_), .B(new_n377_), .ZN(new_n378_));
  OAI22_X1   g00122(.A1(new_n374_), .A2(new_n375_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1     g00123(.I(new_n379_), .ZN(new_n380_));
  NOR4_X1    g00124(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .A4(new_n378_), .ZN(new_n381_));
  NOR2_X1    g00125(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1   g00126(.A1(new_n382_), .A2(new_n265_), .B(new_n372_), .ZN(new_n383_));
  NOR2_X1    g00127(.A1(new_n383_), .A2(new_n270_), .ZN(new_n384_));
  NAND2_X1   g00128(.A1(new_n383_), .A2(new_n270_), .ZN(new_n385_));
  INV_X1     g00129(.I(new_n385_), .ZN(new_n386_));
  OAI21_X1   g00130(.A1(new_n386_), .A2(new_n384_), .B(new_n312_), .ZN(new_n387_));
  INV_X1     g00131(.I(new_n384_), .ZN(new_n388_));
  NAND3_X1   g00132(.A1(new_n388_), .A2(new_n385_), .A3(\a[5] ), .ZN(new_n389_));
  OAI21_X1   g00133(.A1(\a[4] ), .A2(new_n312_), .B(new_n270_), .ZN(new_n390_));
  OAI21_X1   g00134(.A1(new_n316_), .A2(\a[5] ), .B(\a[2] ), .ZN(new_n391_));
  NAND3_X1   g00135(.A1(new_n304_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NOR2_X1    g00136(.A1(new_n392_), .A2(new_n258_), .ZN(new_n393_));
  OAI22_X1   g00137(.A1(new_n321_), .A2(new_n276_), .B1(new_n325_), .B2(new_n275_), .ZN(new_n394_));
  NOR2_X1    g00138(.A1(new_n318_), .A2(new_n282_), .ZN(new_n395_));
  OR3_X2     g00139(.A1(new_n394_), .A2(new_n393_), .A3(new_n395_), .Z(new_n396_));
  NAND2_X1   g00140(.A1(new_n327_), .A2(new_n359_), .ZN(new_n397_));
  NAND2_X1   g00141(.A1(new_n397_), .A2(new_n396_), .ZN(new_n398_));
  NOR2_X1    g00142(.A1(new_n397_), .A2(new_n396_), .ZN(new_n399_));
  INV_X1     g00143(.I(new_n399_), .ZN(new_n400_));
  NAND2_X1   g00144(.A1(new_n400_), .A2(new_n398_), .ZN(new_n401_));
  NAND3_X1   g00145(.A1(new_n387_), .A2(new_n389_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1   g00146(.A1(new_n388_), .A2(new_n385_), .B(\a[5] ), .ZN(new_n403_));
  NOR3_X1    g00147(.A1(new_n386_), .A2(new_n384_), .A3(new_n312_), .ZN(new_n404_));
  INV_X1     g00148(.I(new_n401_), .ZN(new_n405_));
  OAI21_X1   g00149(.A1(new_n403_), .A2(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NAND2_X1   g00150(.A1(new_n406_), .A2(new_n402_), .ZN(new_n407_));
  NAND3_X1   g00151(.A1(new_n336_), .A2(\a[5] ), .A3(new_n306_), .ZN(new_n408_));
  INV_X1     g00152(.I(new_n408_), .ZN(new_n409_));
  NOR3_X1    g00153(.A1(new_n337_), .A2(new_n328_), .A3(new_n359_), .ZN(new_n410_));
  NOR2_X1    g00154(.A1(new_n410_), .A2(new_n409_), .ZN(new_n411_));
  XOR2_X1    g00155(.A1(new_n354_), .A2(\a[2] ), .Z(new_n412_));
  NOR2_X1    g00156(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1   g00157(.A1(new_n366_), .A2(new_n368_), .B(new_n413_), .ZN(new_n414_));
  XOR2_X1    g00158(.A1(new_n407_), .A2(new_n414_), .Z(\f[5] ));
  INV_X1     g00159(.I(\a[6] ), .ZN(new_n416_));
  NOR2_X1    g00160(.A1(new_n312_), .A2(new_n416_), .ZN(new_n417_));
  NOR2_X1    g00161(.A1(\a[5] ), .A2(\a[6] ), .ZN(new_n418_));
  NOR3_X1    g00162(.A1(new_n417_), .A2(new_n258_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1     g00163(.I(new_n419_), .ZN(new_n420_));
  OAI21_X1   g00164(.A1(new_n397_), .A2(new_n396_), .B(new_n420_), .ZN(new_n421_));
  NOR3_X1    g00165(.A1(new_n397_), .A2(new_n396_), .A3(new_n420_), .ZN(new_n422_));
  INV_X1     g00166(.I(new_n422_), .ZN(new_n423_));
  NAND2_X1   g00167(.A1(new_n423_), .A2(new_n421_), .ZN(new_n424_));
  OAI22_X1   g00168(.A1(new_n321_), .A2(new_n290_), .B1(new_n325_), .B2(new_n276_), .ZN(new_n425_));
  NOR2_X1    g00169(.A1(new_n392_), .A2(new_n275_), .ZN(new_n426_));
  OAI21_X1   g00170(.A1(new_n296_), .A2(new_n297_), .B(\b[3] ), .ZN(new_n427_));
  NAND3_X1   g00171(.A1(new_n293_), .A2(new_n294_), .A3(new_n290_), .ZN(new_n428_));
  NAND2_X1   g00172(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1    g00173(.A1(new_n429_), .A2(new_n318_), .ZN(new_n430_));
  NOR3_X1    g00174(.A1(new_n425_), .A2(new_n430_), .A3(new_n426_), .ZN(new_n431_));
  NOR2_X1    g00175(.A1(new_n431_), .A2(new_n312_), .ZN(new_n432_));
  NOR4_X1    g00176(.A1(new_n425_), .A2(new_n430_), .A3(\a[5] ), .A4(new_n426_), .ZN(new_n433_));
  NOR2_X1    g00177(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1     g00178(.I(new_n434_), .ZN(new_n435_));
  XOR2_X1    g00179(.A1(new_n424_), .A2(new_n435_), .Z(new_n436_));
  INV_X1     g00180(.I(new_n436_), .ZN(new_n437_));
  INV_X1     g00181(.I(\b[6] ), .ZN(new_n438_));
  OAI22_X1   g00182(.A1(new_n277_), .A2(new_n438_), .B1(new_n377_), .B2(new_n262_), .ZN(new_n439_));
  AOI21_X1   g00183(.A1(\b[4] ), .A2(new_n283_), .B(new_n439_), .ZN(new_n440_));
  NAND3_X1   g00184(.A1(new_n344_), .A2(new_n345_), .A3(new_n377_), .ZN(new_n441_));
  AOI21_X1   g00185(.A1(new_n441_), .A2(\b[4] ), .B(\b[3] ), .ZN(new_n442_));
  AOI21_X1   g00186(.A1(new_n373_), .A2(\b[5] ), .B(\b[4] ), .ZN(new_n443_));
  XNOR2_X1   g00187(.A1(\b[5] ), .A2(\b[6] ), .ZN(new_n444_));
  INV_X1     g00188(.I(new_n444_), .ZN(new_n445_));
  OAI21_X1   g00189(.A1(new_n442_), .A2(new_n443_), .B(new_n445_), .ZN(new_n446_));
  INV_X1     g00190(.I(new_n446_), .ZN(new_n447_));
  XOR2_X1    g00191(.A1(\b[5] ), .A2(\b[6] ), .Z(new_n448_));
  NOR3_X1    g00192(.A1(new_n442_), .A2(new_n443_), .A3(new_n448_), .ZN(new_n449_));
  NOR2_X1    g00193(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1   g00194(.A1(new_n450_), .A2(new_n279_), .B(new_n440_), .ZN(new_n451_));
  XOR2_X1    g00195(.A1(new_n451_), .A2(new_n270_), .Z(new_n452_));
  INV_X1     g00196(.I(new_n452_), .ZN(new_n453_));
  XOR2_X1    g00197(.A1(new_n396_), .A2(new_n312_), .Z(new_n454_));
  NAND2_X1   g00198(.A1(new_n454_), .A2(new_n397_), .ZN(new_n455_));
  NAND4_X1   g00199(.A1(new_n455_), .A2(new_n388_), .A3(new_n385_), .A4(new_n400_), .ZN(new_n456_));
  OAI21_X1   g00200(.A1(new_n407_), .A2(new_n414_), .B(new_n456_), .ZN(new_n457_));
  NAND2_X1   g00201(.A1(new_n457_), .A2(new_n453_), .ZN(new_n458_));
  OAI21_X1   g00202(.A1(new_n363_), .A2(new_n356_), .B(new_n364_), .ZN(new_n459_));
  NAND3_X1   g00203(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n460_));
  NAND2_X1   g00204(.A1(new_n460_), .A2(new_n459_), .ZN(new_n461_));
  NAND2_X1   g00205(.A1(new_n309_), .A2(new_n289_), .ZN(new_n462_));
  NAND2_X1   g00206(.A1(new_n462_), .A2(new_n307_), .ZN(new_n463_));
  OAI22_X1   g00207(.A1(new_n463_), .A2(new_n461_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n464_));
  NAND3_X1   g00208(.A1(new_n464_), .A2(new_n402_), .A3(new_n406_), .ZN(new_n465_));
  NAND3_X1   g00209(.A1(new_n465_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n466_));
  NAND2_X1   g00210(.A1(new_n466_), .A2(new_n458_), .ZN(new_n467_));
  XOR2_X1    g00211(.A1(new_n467_), .A2(new_n437_), .Z(\f[6] ));
  NOR2_X1    g00212(.A1(new_n457_), .A2(new_n453_), .ZN(new_n469_));
  AOI21_X1   g00213(.A1(new_n437_), .A2(new_n458_), .B(new_n469_), .ZN(new_n470_));
  INV_X1     g00214(.I(\b[7] ), .ZN(new_n471_));
  OAI22_X1   g00215(.A1(new_n277_), .A2(new_n471_), .B1(new_n438_), .B2(new_n262_), .ZN(new_n472_));
  AOI21_X1   g00216(.A1(\b[5] ), .A2(new_n283_), .B(new_n472_), .ZN(new_n473_));
  NOR2_X1    g00217(.A1(new_n442_), .A2(new_n443_), .ZN(new_n474_));
  NOR3_X1    g00218(.A1(new_n474_), .A2(\b[5] ), .A3(new_n438_), .ZN(new_n475_));
  NOR4_X1    g00219(.A1(new_n442_), .A2(new_n443_), .A3(new_n377_), .A4(\b[6] ), .ZN(new_n476_));
  OAI21_X1   g00220(.A1(new_n475_), .A2(new_n476_), .B(\b[7] ), .ZN(new_n477_));
  OAI21_X1   g00221(.A1(new_n376_), .A2(new_n339_), .B(new_n290_), .ZN(new_n478_));
  NOR2_X1    g00222(.A1(new_n349_), .A2(new_n350_), .ZN(new_n479_));
  OAI21_X1   g00223(.A1(new_n479_), .A2(new_n377_), .B(new_n339_), .ZN(new_n480_));
  NAND2_X1   g00224(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1   g00225(.A1(new_n481_), .A2(new_n377_), .A3(\b[6] ), .ZN(new_n482_));
  INV_X1     g00226(.I(new_n476_), .ZN(new_n483_));
  NAND3_X1   g00227(.A1(new_n482_), .A2(new_n471_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1   g00228(.A1(new_n484_), .A2(new_n477_), .ZN(new_n485_));
  OAI21_X1   g00229(.A1(new_n485_), .A2(new_n279_), .B(new_n473_), .ZN(new_n486_));
  XOR2_X1    g00230(.A1(new_n486_), .A2(\a[2] ), .Z(new_n487_));
  INV_X1     g00231(.I(\a[8] ), .ZN(new_n488_));
  XNOR2_X1   g00232(.A1(\a[5] ), .A2(\a[6] ), .ZN(new_n489_));
  XOR2_X1    g00233(.A1(\a[7] ), .A2(\a[8] ), .Z(new_n490_));
  NOR3_X1    g00234(.A1(new_n489_), .A2(new_n490_), .A3(new_n275_), .ZN(new_n491_));
  NAND3_X1   g00235(.A1(new_n312_), .A2(new_n416_), .A3(\a[7] ), .ZN(new_n492_));
  INV_X1     g00236(.I(\a[7] ), .ZN(new_n493_));
  NAND3_X1   g00237(.A1(new_n493_), .A2(\a[5] ), .A3(\a[6] ), .ZN(new_n494_));
  AOI21_X1   g00238(.A1(new_n492_), .A2(new_n494_), .B(new_n258_), .ZN(new_n495_));
  XNOR2_X1   g00239(.A1(\a[7] ), .A2(\a[8] ), .ZN(new_n496_));
  NOR3_X1    g00240(.A1(new_n313_), .A2(new_n489_), .A3(new_n496_), .ZN(new_n497_));
  NOR3_X1    g00241(.A1(new_n497_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n498_));
  NOR2_X1    g00242(.A1(new_n498_), .A2(new_n488_), .ZN(new_n499_));
  XOR2_X1    g00243(.A1(\a[5] ), .A2(\a[6] ), .Z(new_n500_));
  NAND2_X1   g00244(.A1(\a[7] ), .A2(\a[8] ), .ZN(new_n501_));
  NOR2_X1    g00245(.A1(\a[7] ), .A2(\a[8] ), .ZN(new_n502_));
  INV_X1     g00246(.I(new_n502_), .ZN(new_n503_));
  NAND2_X1   g00247(.A1(new_n503_), .A2(new_n501_), .ZN(new_n504_));
  NAND3_X1   g00248(.A1(new_n504_), .A2(new_n500_), .A3(\b[1] ), .ZN(new_n505_));
  NOR3_X1    g00249(.A1(new_n493_), .A2(\a[5] ), .A3(\a[6] ), .ZN(new_n506_));
  NOR3_X1    g00250(.A1(new_n312_), .A2(new_n416_), .A3(\a[7] ), .ZN(new_n507_));
  OAI21_X1   g00251(.A1(new_n507_), .A2(new_n506_), .B(\b[0] ), .ZN(new_n508_));
  NAND2_X1   g00252(.A1(new_n493_), .A2(\a[8] ), .ZN(new_n509_));
  NAND2_X1   g00253(.A1(new_n488_), .A2(\a[7] ), .ZN(new_n510_));
  NAND2_X1   g00254(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1   g00255(.A1(new_n511_), .A2(new_n263_), .A3(new_n500_), .ZN(new_n512_));
  NAND3_X1   g00256(.A1(new_n512_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n513_));
  NOR2_X1    g00257(.A1(new_n513_), .A2(\a[8] ), .ZN(new_n514_));
  OAI22_X1   g00258(.A1(new_n499_), .A2(new_n514_), .B1(new_n488_), .B2(new_n419_), .ZN(new_n515_));
  NAND2_X1   g00259(.A1(new_n312_), .A2(\a[6] ), .ZN(new_n516_));
  NAND2_X1   g00260(.A1(new_n416_), .A2(\a[5] ), .ZN(new_n517_));
  AOI22_X1   g00261(.A1(new_n501_), .A2(new_n503_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  AOI21_X1   g00262(.A1(new_n518_), .A2(\b[1] ), .B(new_n495_), .ZN(new_n519_));
  NAND4_X1   g00263(.A1(new_n519_), .A2(\a[8] ), .A3(new_n420_), .A4(new_n512_), .ZN(new_n520_));
  NOR2_X1    g00264(.A1(new_n392_), .A2(new_n276_), .ZN(new_n521_));
  OAI22_X1   g00265(.A1(new_n321_), .A2(new_n339_), .B1(new_n325_), .B2(new_n290_), .ZN(new_n522_));
  NOR2_X1    g00266(.A1(new_n352_), .A2(new_n318_), .ZN(new_n523_));
  NOR3_X1    g00267(.A1(new_n523_), .A2(new_n522_), .A3(new_n521_), .ZN(new_n524_));
  NAND2_X1   g00268(.A1(new_n524_), .A2(new_n312_), .ZN(new_n525_));
  NOR2_X1    g00269(.A1(new_n524_), .A2(new_n312_), .ZN(new_n526_));
  INV_X1     g00270(.I(new_n526_), .ZN(new_n527_));
  AOI22_X1   g00271(.A1(new_n527_), .A2(new_n525_), .B1(new_n515_), .B2(new_n520_), .ZN(new_n528_));
  NAND4_X1   g00272(.A1(new_n527_), .A2(new_n525_), .A3(new_n515_), .A4(new_n520_), .ZN(new_n529_));
  INV_X1     g00273(.I(new_n529_), .ZN(new_n530_));
  NOR2_X1    g00274(.A1(new_n530_), .A2(new_n528_), .ZN(new_n531_));
  OAI21_X1   g00275(.A1(new_n434_), .A2(new_n422_), .B(new_n421_), .ZN(new_n532_));
  INV_X1     g00276(.I(new_n532_), .ZN(new_n533_));
  XOR2_X1    g00277(.A1(new_n531_), .A2(new_n533_), .Z(new_n534_));
  NOR2_X1    g00278(.A1(new_n534_), .A2(new_n487_), .ZN(new_n535_));
  NAND2_X1   g00279(.A1(new_n534_), .A2(new_n487_), .ZN(new_n536_));
  INV_X1     g00280(.I(new_n536_), .ZN(new_n537_));
  NOR2_X1    g00281(.A1(new_n537_), .A2(new_n535_), .ZN(new_n538_));
  XOR2_X1    g00282(.A1(new_n470_), .A2(new_n538_), .Z(\f[7] ));
  OAI21_X1   g00283(.A1(new_n532_), .A2(new_n528_), .B(new_n529_), .ZN(new_n540_));
  INV_X1     g00284(.I(new_n540_), .ZN(new_n541_));
  NAND2_X1   g00285(.A1(new_n505_), .A2(new_n508_), .ZN(new_n542_));
  NOR4_X1    g00286(.A1(new_n542_), .A2(new_n488_), .A3(new_n419_), .A4(new_n497_), .ZN(new_n543_));
  NOR3_X1    g00287(.A1(new_n282_), .A2(new_n489_), .A3(new_n496_), .ZN(new_n544_));
  NAND3_X1   g00288(.A1(new_n504_), .A2(new_n500_), .A3(\b[2] ), .ZN(new_n545_));
  OAI21_X1   g00289(.A1(new_n507_), .A2(new_n506_), .B(\b[1] ), .ZN(new_n546_));
  NOR4_X1    g00290(.A1(new_n312_), .A2(new_n416_), .A3(new_n493_), .A4(\a[8] ), .ZN(new_n547_));
  NOR4_X1    g00291(.A1(new_n488_), .A2(\a[5] ), .A3(\a[6] ), .A4(\a[7] ), .ZN(new_n548_));
  OAI21_X1   g00292(.A1(new_n547_), .A2(new_n548_), .B(\b[0] ), .ZN(new_n549_));
  NAND3_X1   g00293(.A1(new_n545_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  OAI21_X1   g00294(.A1(new_n550_), .A2(new_n544_), .B(\a[8] ), .ZN(new_n551_));
  OAI21_X1   g00295(.A1(new_n275_), .A2(\b[0] ), .B(\b[2] ), .ZN(new_n552_));
  NAND3_X1   g00296(.A1(new_n258_), .A2(new_n276_), .A3(\b[1] ), .ZN(new_n553_));
  NAND2_X1   g00297(.A1(new_n553_), .A2(new_n552_), .ZN(new_n554_));
  NAND3_X1   g00298(.A1(new_n554_), .A2(new_n511_), .A3(new_n500_), .ZN(new_n555_));
  AOI21_X1   g00299(.A1(new_n492_), .A2(new_n494_), .B(new_n275_), .ZN(new_n556_));
  AOI21_X1   g00300(.A1(new_n518_), .A2(\b[2] ), .B(new_n556_), .ZN(new_n557_));
  NAND4_X1   g00301(.A1(new_n557_), .A2(new_n488_), .A3(new_n555_), .A4(new_n549_), .ZN(new_n558_));
  AOI21_X1   g00302(.A1(new_n551_), .A2(new_n558_), .B(new_n543_), .ZN(new_n559_));
  NAND4_X1   g00303(.A1(new_n555_), .A2(new_n545_), .A3(new_n546_), .A4(new_n549_), .ZN(new_n560_));
  NOR4_X1    g00304(.A1(new_n560_), .A2(new_n513_), .A3(new_n488_), .A4(new_n419_), .ZN(new_n561_));
  OAI21_X1   g00305(.A1(new_n479_), .A2(new_n339_), .B(\b[3] ), .ZN(new_n562_));
  NAND2_X1   g00306(.A1(new_n479_), .A2(new_n339_), .ZN(new_n563_));
  INV_X1     g00307(.I(new_n378_), .ZN(new_n564_));
  NAND4_X1   g00308(.A1(new_n562_), .A2(new_n563_), .A3(new_n441_), .A4(new_n564_), .ZN(new_n565_));
  NAND2_X1   g00309(.A1(new_n565_), .A2(new_n379_), .ZN(new_n566_));
  OAI22_X1   g00310(.A1(new_n321_), .A2(new_n377_), .B1(new_n325_), .B2(new_n339_), .ZN(new_n567_));
  NOR2_X1    g00311(.A1(new_n392_), .A2(new_n290_), .ZN(new_n568_));
  NOR2_X1    g00312(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1   g00313(.A1(new_n566_), .A2(new_n318_), .B(new_n569_), .ZN(new_n570_));
  NOR2_X1    g00314(.A1(new_n570_), .A2(\a[5] ), .ZN(new_n571_));
  AND2_X2    g00315(.A1(new_n570_), .A2(\a[5] ), .Z(new_n572_));
  OAI22_X1   g00316(.A1(new_n572_), .A2(new_n571_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n573_));
  INV_X1     g00317(.I(new_n573_), .ZN(new_n574_));
  NOR4_X1    g00318(.A1(new_n572_), .A2(new_n571_), .A3(new_n559_), .A4(new_n561_), .ZN(new_n575_));
  NOR2_X1    g00319(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1     g00320(.I(\b[8] ), .ZN(new_n577_));
  OAI22_X1   g00321(.A1(new_n277_), .A2(new_n577_), .B1(new_n471_), .B2(new_n262_), .ZN(new_n578_));
  AOI21_X1   g00322(.A1(\b[6] ), .A2(new_n283_), .B(new_n578_), .ZN(new_n579_));
  XOR2_X1    g00323(.A1(\b[7] ), .A2(\b[8] ), .Z(new_n580_));
  NOR3_X1    g00324(.A1(new_n442_), .A2(new_n443_), .A3(new_n377_), .ZN(new_n581_));
  OAI21_X1   g00325(.A1(new_n581_), .A2(\b[6] ), .B(\b[7] ), .ZN(new_n582_));
  OAI21_X1   g00326(.A1(new_n474_), .A2(\b[5] ), .B(\b[6] ), .ZN(new_n583_));
  AOI21_X1   g00327(.A1(new_n582_), .A2(new_n583_), .B(new_n580_), .ZN(new_n584_));
  NAND3_X1   g00328(.A1(new_n582_), .A2(new_n583_), .A3(new_n580_), .ZN(new_n585_));
  INV_X1     g00329(.I(new_n585_), .ZN(new_n586_));
  NOR2_X1    g00330(.A1(new_n586_), .A2(new_n584_), .ZN(new_n587_));
  OAI21_X1   g00331(.A1(new_n587_), .A2(new_n279_), .B(new_n579_), .ZN(new_n588_));
  XOR2_X1    g00332(.A1(new_n588_), .A2(\a[2] ), .Z(new_n589_));
  NOR2_X1    g00333(.A1(new_n589_), .A2(new_n576_), .ZN(new_n590_));
  INV_X1     g00334(.I(new_n576_), .ZN(new_n591_));
  INV_X1     g00335(.I(new_n589_), .ZN(new_n592_));
  NOR2_X1    g00336(.A1(new_n592_), .A2(new_n591_), .ZN(new_n593_));
  NOR3_X1    g00337(.A1(new_n593_), .A2(new_n541_), .A3(new_n590_), .ZN(new_n594_));
  INV_X1     g00338(.I(new_n590_), .ZN(new_n595_));
  INV_X1     g00339(.I(new_n593_), .ZN(new_n596_));
  AOI21_X1   g00340(.A1(new_n596_), .A2(new_n595_), .B(new_n540_), .ZN(new_n597_));
  NOR2_X1    g00341(.A1(new_n597_), .A2(new_n594_), .ZN(new_n598_));
  INV_X1     g00342(.I(new_n535_), .ZN(new_n599_));
  AOI21_X1   g00343(.A1(new_n470_), .A2(new_n599_), .B(new_n537_), .ZN(new_n600_));
  XNOR2_X1   g00344(.A1(new_n600_), .A2(new_n598_), .ZN(\f[8] ));
  INV_X1     g00345(.I(new_n392_), .ZN(new_n602_));
  OAI22_X1   g00346(.A1(new_n321_), .A2(new_n438_), .B1(new_n325_), .B2(new_n377_), .ZN(new_n603_));
  AOI21_X1   g00347(.A1(\b[4] ), .A2(new_n602_), .B(new_n603_), .ZN(new_n604_));
  OAI21_X1   g00348(.A1(new_n450_), .A2(new_n318_), .B(new_n604_), .ZN(new_n605_));
  XOR2_X1    g00349(.A1(new_n605_), .A2(new_n312_), .Z(new_n606_));
  NOR2_X1    g00350(.A1(new_n416_), .A2(\a[5] ), .ZN(new_n607_));
  NOR2_X1    g00351(.A1(new_n312_), .A2(\a[6] ), .ZN(new_n608_));
  INV_X1     g00352(.I(new_n501_), .ZN(new_n609_));
  OAI22_X1   g00353(.A1(new_n609_), .A2(new_n502_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n610_));
  NOR2_X1    g00354(.A1(new_n610_), .A2(new_n290_), .ZN(new_n611_));
  NOR2_X1    g00355(.A1(new_n507_), .A2(new_n506_), .ZN(new_n612_));
  NOR2_X1    g00356(.A1(new_n612_), .A2(new_n276_), .ZN(new_n613_));
  NAND4_X1   g00357(.A1(new_n488_), .A2(\a[5] ), .A3(\a[6] ), .A4(\a[7] ), .ZN(new_n614_));
  NAND3_X1   g00358(.A1(new_n418_), .A2(new_n493_), .A3(\a[8] ), .ZN(new_n615_));
  AOI21_X1   g00359(.A1(new_n615_), .A2(new_n614_), .B(new_n275_), .ZN(new_n616_));
  NOR3_X1    g00360(.A1(new_n611_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n617_));
  AOI22_X1   g00361(.A1(new_n516_), .A2(new_n517_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n618_));
  NAND2_X1   g00362(.A1(new_n299_), .A2(new_n618_), .ZN(new_n619_));
  AOI21_X1   g00363(.A1(new_n617_), .A2(new_n619_), .B(new_n488_), .ZN(new_n620_));
  OAI22_X1   g00364(.A1(new_n610_), .A2(new_n290_), .B1(new_n276_), .B2(new_n612_), .ZN(new_n621_));
  NOR2_X1    g00365(.A1(new_n488_), .A2(\a[7] ), .ZN(new_n622_));
  NOR2_X1    g00366(.A1(new_n493_), .A2(\a[8] ), .ZN(new_n623_));
  OAI22_X1   g00367(.A1(new_n607_), .A2(new_n608_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NOR3_X1    g00368(.A1(new_n624_), .A2(new_n298_), .A3(new_n295_), .ZN(new_n625_));
  NOR4_X1    g00369(.A1(new_n621_), .A2(new_n625_), .A3(\a[8] ), .A4(new_n616_), .ZN(new_n626_));
  NOR2_X1    g00370(.A1(new_n620_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1     g00371(.I(\a[9] ), .ZN(new_n628_));
  NOR2_X1    g00372(.A1(new_n628_), .A2(\a[8] ), .ZN(new_n629_));
  NOR2_X1    g00373(.A1(new_n488_), .A2(\a[9] ), .ZN(new_n630_));
  NOR2_X1    g00374(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1    g00375(.A1(new_n631_), .A2(new_n258_), .ZN(new_n632_));
  INV_X1     g00376(.I(new_n632_), .ZN(new_n633_));
  NOR2_X1    g00377(.A1(new_n627_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1   g00378(.A1(new_n518_), .A2(\b[3] ), .ZN(new_n635_));
  NAND2_X1   g00379(.A1(new_n492_), .A2(new_n494_), .ZN(new_n636_));
  NAND2_X1   g00380(.A1(new_n636_), .A2(\b[2] ), .ZN(new_n637_));
  INV_X1     g00381(.I(new_n616_), .ZN(new_n638_));
  NAND3_X1   g00382(.A1(new_n635_), .A2(new_n638_), .A3(new_n637_), .ZN(new_n639_));
  OAI21_X1   g00383(.A1(new_n639_), .A2(new_n625_), .B(\a[8] ), .ZN(new_n640_));
  AOI22_X1   g00384(.A1(new_n518_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n636_), .ZN(new_n641_));
  NAND4_X1   g00385(.A1(new_n619_), .A2(new_n488_), .A3(new_n641_), .A4(new_n638_), .ZN(new_n642_));
  NAND2_X1   g00386(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1    g00387(.A1(new_n643_), .A2(new_n632_), .ZN(new_n644_));
  NOR2_X1    g00388(.A1(new_n634_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1    g00389(.A1(new_n645_), .A2(new_n561_), .ZN(new_n646_));
  NOR3_X1    g00390(.A1(new_n489_), .A2(new_n490_), .A3(new_n276_), .ZN(new_n647_));
  AOI21_X1   g00391(.A1(new_n615_), .A2(new_n614_), .B(new_n258_), .ZN(new_n648_));
  NOR4_X1    g00392(.A1(new_n544_), .A2(new_n647_), .A3(new_n556_), .A4(new_n648_), .ZN(new_n649_));
  NAND4_X1   g00393(.A1(new_n649_), .A2(\a[8] ), .A3(new_n420_), .A4(new_n498_), .ZN(new_n650_));
  NOR3_X1    g00394(.A1(new_n634_), .A2(new_n644_), .A3(new_n650_), .ZN(new_n651_));
  NOR2_X1    g00395(.A1(new_n646_), .A2(new_n651_), .ZN(new_n652_));
  XOR2_X1    g00396(.A1(new_n652_), .A2(new_n606_), .Z(new_n653_));
  OAI21_X1   g00397(.A1(new_n540_), .A2(new_n575_), .B(new_n573_), .ZN(new_n654_));
  XOR2_X1    g00398(.A1(new_n653_), .A2(new_n654_), .Z(new_n655_));
  INV_X1     g00399(.I(new_n655_), .ZN(new_n656_));
  NAND2_X1   g00400(.A1(new_n283_), .A2(\b[7] ), .ZN(new_n657_));
  AOI22_X1   g00401(.A1(new_n267_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n261_), .ZN(new_n658_));
  NAND2_X1   g00402(.A1(new_n582_), .A2(new_n583_), .ZN(new_n659_));
  AOI21_X1   g00403(.A1(new_n659_), .A2(\b[8] ), .B(new_n471_), .ZN(new_n660_));
  NOR2_X1    g00404(.A1(new_n659_), .A2(\b[8] ), .ZN(new_n661_));
  NOR2_X1    g00405(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1   g00406(.A1(new_n478_), .A2(new_n480_), .A3(\b[5] ), .ZN(new_n663_));
  AOI21_X1   g00407(.A1(new_n663_), .A2(new_n438_), .B(new_n471_), .ZN(new_n664_));
  AOI21_X1   g00408(.A1(new_n481_), .A2(new_n377_), .B(new_n438_), .ZN(new_n665_));
  NOR3_X1    g00409(.A1(new_n664_), .A2(new_n665_), .A3(\b[9] ), .ZN(new_n666_));
  INV_X1     g00410(.I(\b[9] ), .ZN(new_n667_));
  NOR2_X1    g00411(.A1(new_n664_), .A2(new_n665_), .ZN(new_n668_));
  NOR2_X1    g00412(.A1(new_n668_), .A2(new_n667_), .ZN(new_n669_));
  NOR2_X1    g00413(.A1(new_n669_), .A2(new_n666_), .ZN(new_n670_));
  NOR2_X1    g00414(.A1(new_n670_), .A2(new_n662_), .ZN(new_n671_));
  NAND3_X1   g00415(.A1(new_n582_), .A2(new_n583_), .A3(new_n667_), .ZN(new_n672_));
  NAND2_X1   g00416(.A1(new_n659_), .A2(\b[9] ), .ZN(new_n673_));
  NAND2_X1   g00417(.A1(new_n673_), .A2(new_n672_), .ZN(new_n674_));
  NOR3_X1    g00418(.A1(new_n674_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n675_));
  NOR2_X1    g00419(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1   g00420(.A1(new_n676_), .A2(new_n265_), .ZN(new_n677_));
  NAND4_X1   g00421(.A1(new_n677_), .A2(\a[2] ), .A3(new_n657_), .A4(new_n658_), .ZN(new_n678_));
  NAND3_X1   g00422(.A1(new_n677_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n679_));
  NAND2_X1   g00423(.A1(new_n679_), .A2(new_n270_), .ZN(new_n680_));
  NAND2_X1   g00424(.A1(new_n680_), .A2(new_n678_), .ZN(new_n681_));
  NAND2_X1   g00425(.A1(new_n656_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1   g00426(.A1(new_n655_), .A2(new_n678_), .A3(new_n680_), .ZN(new_n683_));
  NAND2_X1   g00427(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1   g00428(.A1(new_n465_), .A2(new_n456_), .B(new_n452_), .ZN(new_n685_));
  OAI21_X1   g00429(.A1(new_n436_), .A2(new_n685_), .B(new_n466_), .ZN(new_n686_));
  OAI21_X1   g00430(.A1(new_n686_), .A2(new_n535_), .B(new_n536_), .ZN(new_n687_));
  XOR2_X1    g00431(.A1(new_n576_), .A2(new_n541_), .Z(new_n688_));
  NOR2_X1    g00432(.A1(new_n688_), .A2(new_n592_), .ZN(new_n689_));
  AOI21_X1   g00433(.A1(new_n687_), .A2(new_n598_), .B(new_n689_), .ZN(new_n690_));
  XOR2_X1    g00434(.A1(new_n690_), .A2(new_n684_), .Z(\f[9] ));
  OAI21_X1   g00435(.A1(new_n690_), .A2(new_n684_), .B(new_n682_), .ZN(new_n692_));
  NAND2_X1   g00436(.A1(new_n654_), .A2(new_n606_), .ZN(new_n693_));
  OAI21_X1   g00437(.A1(new_n654_), .A2(new_n606_), .B(new_n652_), .ZN(new_n694_));
  NAND2_X1   g00438(.A1(new_n694_), .A2(new_n693_), .ZN(new_n695_));
  OAI22_X1   g00439(.A1(new_n321_), .A2(new_n471_), .B1(new_n325_), .B2(new_n438_), .ZN(new_n696_));
  NOR2_X1    g00440(.A1(new_n392_), .A2(new_n377_), .ZN(new_n697_));
  NOR2_X1    g00441(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI21_X1   g00442(.A1(new_n485_), .A2(new_n318_), .B(new_n698_), .ZN(new_n699_));
  NAND2_X1   g00443(.A1(new_n699_), .A2(\a[5] ), .ZN(new_n700_));
  OR2_X2     g00444(.A1(new_n699_), .A2(\a[5] ), .Z(new_n701_));
  NAND2_X1   g00445(.A1(new_n701_), .A2(new_n700_), .ZN(new_n702_));
  NAND2_X1   g00446(.A1(new_n650_), .A2(new_n633_), .ZN(new_n703_));
  NOR3_X1    g00447(.A1(new_n647_), .A2(new_n556_), .A3(new_n648_), .ZN(new_n704_));
  AOI21_X1   g00448(.A1(new_n704_), .A2(new_n555_), .B(new_n488_), .ZN(new_n705_));
  OAI21_X1   g00449(.A1(new_n610_), .A2(new_n276_), .B(new_n546_), .ZN(new_n706_));
  NOR4_X1    g00450(.A1(new_n706_), .A2(\a[8] ), .A3(new_n544_), .A4(new_n648_), .ZN(new_n707_));
  NOR4_X1    g00451(.A1(new_n705_), .A2(new_n707_), .A3(new_n520_), .A4(new_n633_), .ZN(new_n708_));
  AOI21_X1   g00452(.A1(new_n703_), .A2(new_n627_), .B(new_n708_), .ZN(new_n709_));
  NAND2_X1   g00453(.A1(\a[10] ), .A2(\a[11] ), .ZN(new_n710_));
  INV_X1     g00454(.I(new_n710_), .ZN(new_n711_));
  NOR2_X1    g00455(.A1(\a[10] ), .A2(\a[11] ), .ZN(new_n712_));
  OAI22_X1   g00456(.A1(new_n711_), .A2(new_n712_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n713_));
  INV_X1     g00457(.I(\a[10] ), .ZN(new_n714_));
  NOR3_X1    g00458(.A1(new_n714_), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n715_));
  NOR3_X1    g00459(.A1(new_n488_), .A2(new_n628_), .A3(\a[10] ), .ZN(new_n716_));
  NOR2_X1    g00460(.A1(new_n716_), .A2(new_n715_), .ZN(new_n717_));
  OAI22_X1   g00461(.A1(new_n713_), .A2(new_n275_), .B1(new_n258_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1   g00462(.A1(new_n488_), .A2(\a[9] ), .ZN(new_n719_));
  NAND2_X1   g00463(.A1(new_n628_), .A2(\a[8] ), .ZN(new_n720_));
  NAND2_X1   g00464(.A1(new_n714_), .A2(\a[11] ), .ZN(new_n721_));
  INV_X1     g00465(.I(\a[11] ), .ZN(new_n722_));
  NAND2_X1   g00466(.A1(new_n722_), .A2(\a[10] ), .ZN(new_n723_));
  AOI22_X1   g00467(.A1(new_n719_), .A2(new_n720_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1   g00468(.A1(new_n724_), .A2(new_n263_), .ZN(new_n725_));
  INV_X1     g00469(.I(new_n725_), .ZN(new_n726_));
  OAI21_X1   g00470(.A1(new_n726_), .A2(new_n718_), .B(\a[11] ), .ZN(new_n727_));
  INV_X1     g00471(.I(new_n712_), .ZN(new_n728_));
  AOI22_X1   g00472(.A1(new_n710_), .A2(new_n728_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n729_));
  NAND3_X1   g00473(.A1(new_n488_), .A2(new_n628_), .A3(\a[10] ), .ZN(new_n730_));
  NAND3_X1   g00474(.A1(new_n714_), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n731_));
  NAND2_X1   g00475(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  AOI22_X1   g00476(.A1(new_n729_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n732_), .ZN(new_n733_));
  NAND3_X1   g00477(.A1(new_n733_), .A2(new_n722_), .A3(new_n725_), .ZN(new_n734_));
  NOR2_X1    g00478(.A1(new_n632_), .A2(new_n722_), .ZN(new_n735_));
  INV_X1     g00479(.I(new_n735_), .ZN(new_n736_));
  NAND3_X1   g00480(.A1(new_n727_), .A2(new_n734_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1   g00481(.A1(new_n733_), .A2(new_n725_), .B(new_n722_), .ZN(new_n738_));
  NAND2_X1   g00482(.A1(new_n738_), .A2(new_n633_), .ZN(new_n739_));
  NAND3_X1   g00483(.A1(new_n504_), .A2(new_n500_), .A3(\b[4] ), .ZN(new_n740_));
  AOI21_X1   g00484(.A1(new_n492_), .A2(new_n494_), .B(new_n290_), .ZN(new_n741_));
  INV_X1     g00485(.I(new_n741_), .ZN(new_n742_));
  OAI21_X1   g00486(.A1(new_n547_), .A2(new_n548_), .B(\b[2] ), .ZN(new_n743_));
  NAND3_X1   g00487(.A1(new_n742_), .A2(new_n740_), .A3(new_n743_), .ZN(new_n744_));
  OAI22_X1   g00488(.A1(new_n349_), .A2(new_n350_), .B1(new_n347_), .B2(new_n342_), .ZN(new_n745_));
  NAND4_X1   g00489(.A1(new_n343_), .A2(new_n341_), .A3(new_n344_), .A4(new_n345_), .ZN(new_n746_));
  AOI21_X1   g00490(.A1(new_n745_), .A2(new_n746_), .B(new_n624_), .ZN(new_n747_));
  OAI21_X1   g00491(.A1(new_n744_), .A2(new_n747_), .B(\a[8] ), .ZN(new_n748_));
  NOR3_X1    g00492(.A1(new_n489_), .A2(new_n490_), .A3(new_n339_), .ZN(new_n749_));
  AOI21_X1   g00493(.A1(new_n615_), .A2(new_n614_), .B(new_n276_), .ZN(new_n750_));
  NOR3_X1    g00494(.A1(new_n749_), .A2(new_n741_), .A3(new_n750_), .ZN(new_n751_));
  OAI21_X1   g00495(.A1(new_n346_), .A2(new_n351_), .B(new_n618_), .ZN(new_n752_));
  NAND3_X1   g00496(.A1(new_n751_), .A2(new_n752_), .A3(new_n488_), .ZN(new_n753_));
  NAND2_X1   g00497(.A1(new_n748_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1   g00498(.A1(new_n737_), .A2(new_n754_), .A3(new_n739_), .ZN(new_n755_));
  NOR3_X1    g00499(.A1(new_n726_), .A2(new_n718_), .A3(\a[11] ), .ZN(new_n756_));
  NOR3_X1    g00500(.A1(new_n756_), .A2(new_n738_), .A3(new_n735_), .ZN(new_n757_));
  NOR2_X1    g00501(.A1(new_n727_), .A2(new_n632_), .ZN(new_n758_));
  AOI21_X1   g00502(.A1(new_n751_), .A2(new_n752_), .B(new_n488_), .ZN(new_n759_));
  NOR3_X1    g00503(.A1(new_n744_), .A2(new_n747_), .A3(\a[8] ), .ZN(new_n760_));
  NOR2_X1    g00504(.A1(new_n760_), .A2(new_n759_), .ZN(new_n761_));
  OAI21_X1   g00505(.A1(new_n757_), .A2(new_n758_), .B(new_n761_), .ZN(new_n762_));
  NAND3_X1   g00506(.A1(new_n709_), .A2(new_n755_), .A3(new_n762_), .ZN(new_n763_));
  NOR2_X1    g00507(.A1(new_n561_), .A2(new_n632_), .ZN(new_n764_));
  NAND4_X1   g00508(.A1(new_n543_), .A2(new_n551_), .A3(new_n558_), .A4(new_n632_), .ZN(new_n765_));
  OAI21_X1   g00509(.A1(new_n764_), .A2(new_n643_), .B(new_n765_), .ZN(new_n766_));
  NOR3_X1    g00510(.A1(new_n757_), .A2(new_n761_), .A3(new_n758_), .ZN(new_n767_));
  AOI21_X1   g00511(.A1(new_n737_), .A2(new_n739_), .B(new_n754_), .ZN(new_n768_));
  OAI21_X1   g00512(.A1(new_n767_), .A2(new_n768_), .B(new_n766_), .ZN(new_n769_));
  NAND2_X1   g00513(.A1(new_n769_), .A2(new_n763_), .ZN(new_n770_));
  NOR2_X1    g00514(.A1(new_n702_), .A2(new_n770_), .ZN(new_n771_));
  AOI22_X1   g00515(.A1(new_n701_), .A2(new_n700_), .B1(new_n769_), .B2(new_n763_), .ZN(new_n772_));
  NOR2_X1    g00516(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  XNOR2_X1   g00517(.A1(new_n695_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1     g00518(.I(new_n774_), .ZN(new_n775_));
  INV_X1     g00519(.I(\b[10] ), .ZN(new_n776_));
  OAI22_X1   g00520(.A1(new_n277_), .A2(new_n776_), .B1(new_n667_), .B2(new_n262_), .ZN(new_n777_));
  AOI21_X1   g00521(.A1(\b[8] ), .A2(new_n283_), .B(new_n777_), .ZN(new_n778_));
  AOI21_X1   g00522(.A1(new_n672_), .A2(\b[8] ), .B(\b[7] ), .ZN(new_n779_));
  AOI21_X1   g00523(.A1(new_n659_), .A2(\b[9] ), .B(\b[8] ), .ZN(new_n780_));
  NOR2_X1    g00524(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1   g00525(.A1(\b[9] ), .A2(\b[10] ), .ZN(new_n782_));
  NOR2_X1    g00526(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  XOR2_X1    g00527(.A1(\b[9] ), .A2(\b[10] ), .Z(new_n784_));
  INV_X1     g00528(.I(new_n784_), .ZN(new_n785_));
  AOI21_X1   g00529(.A1(new_n781_), .A2(new_n785_), .B(new_n783_), .ZN(new_n786_));
  OAI21_X1   g00530(.A1(new_n786_), .A2(new_n279_), .B(new_n778_), .ZN(new_n787_));
  XOR2_X1    g00531(.A1(new_n787_), .A2(\a[2] ), .Z(new_n788_));
  NOR2_X1    g00532(.A1(new_n775_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1   g00533(.A1(new_n775_), .A2(new_n788_), .ZN(new_n790_));
  INV_X1     g00534(.I(new_n790_), .ZN(new_n791_));
  NOR2_X1    g00535(.A1(new_n791_), .A2(new_n789_), .ZN(new_n792_));
  XOR2_X1    g00536(.A1(new_n692_), .A2(new_n792_), .Z(\f[10] ));
  NAND3_X1   g00537(.A1(new_n770_), .A2(new_n701_), .A3(new_n700_), .ZN(new_n794_));
  OAI21_X1   g00538(.A1(new_n695_), .A2(new_n773_), .B(new_n794_), .ZN(new_n795_));
  INV_X1     g00539(.I(new_n795_), .ZN(new_n796_));
  INV_X1     g00540(.I(new_n580_), .ZN(new_n797_));
  NAND2_X1   g00541(.A1(new_n659_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1   g00542(.A1(new_n798_), .A2(new_n585_), .ZN(new_n799_));
  INV_X1     g00543(.I(new_n325_), .ZN(new_n800_));
  AOI22_X1   g00544(.A1(new_n800_), .A2(\b[7] ), .B1(\b[8] ), .B2(new_n333_), .ZN(new_n801_));
  OAI21_X1   g00545(.A1(new_n438_), .A2(new_n392_), .B(new_n801_), .ZN(new_n802_));
  AOI21_X1   g00546(.A1(new_n799_), .A2(new_n330_), .B(new_n802_), .ZN(new_n803_));
  XOR2_X1    g00547(.A1(new_n803_), .A2(new_n312_), .Z(new_n804_));
  NAND2_X1   g00548(.A1(new_n724_), .A2(new_n554_), .ZN(new_n805_));
  NAND2_X1   g00549(.A1(new_n729_), .A2(\b[2] ), .ZN(new_n806_));
  NAND2_X1   g00550(.A1(new_n732_), .A2(\b[1] ), .ZN(new_n807_));
  AOI21_X1   g00551(.A1(new_n714_), .A2(\a[11] ), .B(\a[8] ), .ZN(new_n808_));
  INV_X1     g00552(.I(new_n808_), .ZN(new_n809_));
  OAI21_X1   g00553(.A1(new_n714_), .A2(\a[11] ), .B(\a[8] ), .ZN(new_n810_));
  NAND4_X1   g00554(.A1(new_n631_), .A2(new_n809_), .A3(\b[0] ), .A4(new_n810_), .ZN(new_n811_));
  NAND4_X1   g00555(.A1(new_n805_), .A2(new_n806_), .A3(new_n811_), .A4(new_n807_), .ZN(new_n812_));
  NAND2_X1   g00556(.A1(new_n812_), .A2(\a[11] ), .ZN(new_n813_));
  NOR2_X1    g00557(.A1(new_n713_), .A2(new_n276_), .ZN(new_n814_));
  NOR2_X1    g00558(.A1(new_n717_), .A2(new_n275_), .ZN(new_n815_));
  NAND2_X1   g00559(.A1(new_n719_), .A2(new_n720_), .ZN(new_n816_));
  INV_X1     g00560(.I(new_n810_), .ZN(new_n817_));
  NOR4_X1    g00561(.A1(new_n816_), .A2(new_n817_), .A3(new_n258_), .A4(new_n808_), .ZN(new_n818_));
  NOR3_X1    g00562(.A1(new_n814_), .A2(new_n818_), .A3(new_n815_), .ZN(new_n819_));
  NAND3_X1   g00563(.A1(new_n819_), .A2(new_n722_), .A3(new_n805_), .ZN(new_n820_));
  NAND4_X1   g00564(.A1(new_n733_), .A2(new_n633_), .A3(\a[11] ), .A4(new_n725_), .ZN(new_n821_));
  INV_X1     g00565(.I(new_n821_), .ZN(new_n822_));
  AOI21_X1   g00566(.A1(new_n813_), .A2(new_n820_), .B(new_n822_), .ZN(new_n823_));
  NAND2_X1   g00567(.A1(new_n733_), .A2(new_n725_), .ZN(new_n824_));
  NOR4_X1    g00568(.A1(new_n812_), .A2(new_n824_), .A3(new_n722_), .A4(new_n632_), .ZN(new_n825_));
  NAND2_X1   g00569(.A1(new_n615_), .A2(new_n614_), .ZN(new_n826_));
  OAI22_X1   g00570(.A1(new_n610_), .A2(new_n377_), .B1(new_n339_), .B2(new_n612_), .ZN(new_n827_));
  AOI21_X1   g00571(.A1(\b[3] ), .A2(new_n826_), .B(new_n827_), .ZN(new_n828_));
  NAND3_X1   g00572(.A1(new_n565_), .A2(new_n379_), .A3(new_n618_), .ZN(new_n829_));
  NAND3_X1   g00573(.A1(new_n829_), .A2(new_n488_), .A3(new_n828_), .ZN(new_n830_));
  INV_X1     g00574(.I(new_n830_), .ZN(new_n831_));
  AOI21_X1   g00575(.A1(new_n829_), .A2(new_n828_), .B(new_n488_), .ZN(new_n832_));
  OAI22_X1   g00576(.A1(new_n831_), .A2(new_n832_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n833_));
  AOI21_X1   g00577(.A1(new_n819_), .A2(new_n805_), .B(new_n722_), .ZN(new_n834_));
  NOR2_X1    g00578(.A1(new_n812_), .A2(\a[11] ), .ZN(new_n835_));
  OAI21_X1   g00579(.A1(new_n835_), .A2(new_n834_), .B(new_n821_), .ZN(new_n836_));
  INV_X1     g00580(.I(new_n825_), .ZN(new_n837_));
  INV_X1     g00581(.I(new_n832_), .ZN(new_n838_));
  NAND4_X1   g00582(.A1(new_n838_), .A2(new_n836_), .A3(new_n837_), .A4(new_n830_), .ZN(new_n839_));
  NAND2_X1   g00583(.A1(new_n833_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1   g00584(.A1(new_n766_), .A2(new_n755_), .B(new_n768_), .ZN(new_n841_));
  XOR2_X1    g00585(.A1(new_n840_), .A2(new_n841_), .Z(new_n842_));
  NOR2_X1    g00586(.A1(new_n842_), .A2(new_n804_), .ZN(new_n843_));
  INV_X1     g00587(.I(new_n843_), .ZN(new_n844_));
  NAND2_X1   g00588(.A1(new_n842_), .A2(new_n804_), .ZN(new_n845_));
  AOI22_X1   g00589(.A1(new_n267_), .A2(\b[11] ), .B1(\b[10] ), .B2(new_n261_), .ZN(new_n846_));
  OAI21_X1   g00590(.A1(new_n667_), .A2(new_n284_), .B(new_n846_), .ZN(new_n847_));
  INV_X1     g00591(.I(new_n847_), .ZN(new_n848_));
  NOR3_X1    g00592(.A1(new_n781_), .A2(\b[9] ), .A3(new_n776_), .ZN(new_n849_));
  NOR4_X1    g00593(.A1(new_n779_), .A2(new_n780_), .A3(new_n667_), .A4(\b[10] ), .ZN(new_n850_));
  OAI21_X1   g00594(.A1(new_n849_), .A2(new_n850_), .B(\b[11] ), .ZN(new_n851_));
  INV_X1     g00595(.I(\b[11] ), .ZN(new_n852_));
  OAI21_X1   g00596(.A1(new_n666_), .A2(new_n577_), .B(new_n471_), .ZN(new_n853_));
  OAI21_X1   g00597(.A1(new_n668_), .A2(new_n667_), .B(new_n577_), .ZN(new_n854_));
  NAND2_X1   g00598(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1   g00599(.A1(new_n855_), .A2(new_n667_), .A3(\b[10] ), .ZN(new_n856_));
  INV_X1     g00600(.I(new_n850_), .ZN(new_n857_));
  NAND3_X1   g00601(.A1(new_n856_), .A2(new_n852_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1   g00602(.A1(new_n858_), .A2(new_n851_), .ZN(new_n859_));
  OAI21_X1   g00603(.A1(new_n859_), .A2(new_n279_), .B(new_n848_), .ZN(new_n860_));
  AND2_X2    g00604(.A1(new_n860_), .A2(\a[2] ), .Z(new_n861_));
  NOR2_X1    g00605(.A1(new_n860_), .A2(\a[2] ), .ZN(new_n862_));
  NOR2_X1    g00606(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1   g00607(.A1(new_n844_), .A2(new_n845_), .B(new_n863_), .ZN(new_n864_));
  NAND3_X1   g00608(.A1(new_n863_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n865_));
  INV_X1     g00609(.I(new_n865_), .ZN(new_n866_));
  NOR3_X1    g00610(.A1(new_n866_), .A2(new_n864_), .A3(new_n796_), .ZN(new_n867_));
  NAND2_X1   g00611(.A1(new_n844_), .A2(new_n845_), .ZN(new_n868_));
  INV_X1     g00612(.I(new_n863_), .ZN(new_n869_));
  NAND2_X1   g00613(.A1(new_n869_), .A2(new_n868_), .ZN(new_n870_));
  AOI21_X1   g00614(.A1(new_n870_), .A2(new_n865_), .B(new_n795_), .ZN(new_n871_));
  NOR2_X1    g00615(.A1(new_n867_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1     g00616(.I(new_n682_), .ZN(new_n873_));
  OR2_X2     g00617(.A1(new_n597_), .A2(new_n594_), .Z(new_n874_));
  INV_X1     g00618(.I(new_n689_), .ZN(new_n875_));
  OAI21_X1   g00619(.A1(new_n874_), .A2(new_n600_), .B(new_n875_), .ZN(new_n876_));
  AOI21_X1   g00620(.A1(new_n876_), .A2(new_n683_), .B(new_n873_), .ZN(new_n877_));
  OAI21_X1   g00621(.A1(new_n877_), .A2(new_n789_), .B(new_n790_), .ZN(new_n878_));
  XOR2_X1    g00622(.A1(new_n878_), .A2(new_n872_), .Z(\f[11] ));
  AOI22_X1   g00623(.A1(new_n800_), .A2(\b[8] ), .B1(\b[9] ), .B2(new_n333_), .ZN(new_n880_));
  OAI21_X1   g00624(.A1(new_n471_), .A2(new_n392_), .B(new_n880_), .ZN(new_n881_));
  INV_X1     g00625(.I(new_n881_), .ZN(new_n882_));
  NAND2_X1   g00626(.A1(new_n676_), .A2(new_n330_), .ZN(new_n883_));
  AOI21_X1   g00627(.A1(new_n883_), .A2(new_n882_), .B(new_n312_), .ZN(new_n884_));
  AND3_X2    g00628(.A1(new_n883_), .A2(new_n312_), .A3(new_n882_), .Z(new_n885_));
  NOR2_X1    g00629(.A1(new_n885_), .A2(new_n884_), .ZN(new_n886_));
  NOR4_X1    g00630(.A1(new_n816_), .A2(new_n817_), .A3(new_n275_), .A4(new_n808_), .ZN(new_n887_));
  OAI21_X1   g00631(.A1(new_n716_), .A2(new_n715_), .B(\b[2] ), .ZN(new_n888_));
  OAI21_X1   g00632(.A1(new_n713_), .A2(new_n290_), .B(new_n888_), .ZN(new_n889_));
  XNOR2_X1   g00633(.A1(\a[10] ), .A2(\a[11] ), .ZN(new_n890_));
  NOR4_X1    g00634(.A1(new_n298_), .A2(new_n295_), .A3(new_n631_), .A4(new_n890_), .ZN(new_n891_));
  NOR3_X1    g00635(.A1(new_n889_), .A2(new_n891_), .A3(new_n887_), .ZN(new_n892_));
  NOR2_X1    g00636(.A1(new_n892_), .A2(new_n722_), .ZN(new_n893_));
  NOR4_X1    g00637(.A1(new_n889_), .A2(new_n891_), .A3(\a[11] ), .A4(new_n887_), .ZN(new_n894_));
  INV_X1     g00638(.I(\a[12] ), .ZN(new_n895_));
  NOR2_X1    g00639(.A1(new_n895_), .A2(\a[11] ), .ZN(new_n896_));
  NOR2_X1    g00640(.A1(new_n722_), .A2(\a[12] ), .ZN(new_n897_));
  NOR2_X1    g00641(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1    g00642(.A1(new_n898_), .A2(new_n258_), .ZN(new_n899_));
  INV_X1     g00643(.I(new_n899_), .ZN(new_n900_));
  OAI21_X1   g00644(.A1(new_n893_), .A2(new_n894_), .B(new_n900_), .ZN(new_n901_));
  NAND4_X1   g00645(.A1(new_n631_), .A2(new_n809_), .A3(\b[1] ), .A4(new_n810_), .ZN(new_n902_));
  AOI21_X1   g00646(.A1(new_n730_), .A2(new_n731_), .B(new_n276_), .ZN(new_n903_));
  AOI21_X1   g00647(.A1(new_n729_), .A2(\b[3] ), .B(new_n903_), .ZN(new_n904_));
  NAND3_X1   g00648(.A1(new_n724_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n905_));
  NAND3_X1   g00649(.A1(new_n904_), .A2(new_n905_), .A3(new_n902_), .ZN(new_n906_));
  NAND2_X1   g00650(.A1(new_n906_), .A2(\a[11] ), .ZN(new_n907_));
  NAND4_X1   g00651(.A1(new_n904_), .A2(new_n905_), .A3(new_n722_), .A4(new_n902_), .ZN(new_n908_));
  NAND3_X1   g00652(.A1(new_n907_), .A2(new_n908_), .A3(new_n899_), .ZN(new_n909_));
  NAND3_X1   g00653(.A1(new_n837_), .A2(new_n901_), .A3(new_n909_), .ZN(new_n910_));
  AOI21_X1   g00654(.A1(new_n907_), .A2(new_n908_), .B(new_n899_), .ZN(new_n911_));
  NOR3_X1    g00655(.A1(new_n893_), .A2(new_n894_), .A3(new_n900_), .ZN(new_n912_));
  OAI21_X1   g00656(.A1(new_n912_), .A2(new_n911_), .B(new_n825_), .ZN(new_n913_));
  AND2_X2    g00657(.A1(new_n910_), .A2(new_n913_), .Z(new_n914_));
  OR3_X2     g00658(.A1(new_n442_), .A2(new_n443_), .A3(new_n448_), .Z(new_n915_));
  NAND2_X1   g00659(.A1(new_n915_), .A2(new_n446_), .ZN(new_n916_));
  INV_X1     g00660(.I(new_n826_), .ZN(new_n917_));
  AOI22_X1   g00661(.A1(new_n518_), .A2(\b[6] ), .B1(\b[5] ), .B2(new_n636_), .ZN(new_n918_));
  OAI21_X1   g00662(.A1(new_n339_), .A2(new_n917_), .B(new_n918_), .ZN(new_n919_));
  AOI21_X1   g00663(.A1(new_n916_), .A2(new_n618_), .B(new_n919_), .ZN(new_n920_));
  XOR2_X1    g00664(.A1(new_n920_), .A2(new_n488_), .Z(new_n921_));
  AOI22_X1   g00665(.A1(new_n838_), .A2(new_n830_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n922_));
  OAI21_X1   g00666(.A1(new_n841_), .A2(new_n922_), .B(new_n839_), .ZN(new_n923_));
  NAND2_X1   g00667(.A1(new_n923_), .A2(new_n921_), .ZN(new_n924_));
  INV_X1     g00668(.I(new_n921_), .ZN(new_n925_));
  NOR4_X1    g00669(.A1(new_n831_), .A2(new_n823_), .A3(new_n825_), .A4(new_n832_), .ZN(new_n926_));
  OAI21_X1   g00670(.A1(new_n709_), .A2(new_n767_), .B(new_n762_), .ZN(new_n927_));
  AOI21_X1   g00671(.A1(new_n927_), .A2(new_n833_), .B(new_n926_), .ZN(new_n928_));
  NAND2_X1   g00672(.A1(new_n928_), .A2(new_n925_), .ZN(new_n929_));
  NAND3_X1   g00673(.A1(new_n929_), .A2(new_n924_), .A3(new_n914_), .ZN(new_n930_));
  AOI21_X1   g00674(.A1(new_n929_), .A2(new_n924_), .B(new_n914_), .ZN(new_n931_));
  INV_X1     g00675(.I(new_n931_), .ZN(new_n932_));
  NAND2_X1   g00676(.A1(new_n932_), .A2(new_n930_), .ZN(new_n933_));
  NOR2_X1    g00677(.A1(new_n933_), .A2(new_n886_), .ZN(new_n934_));
  NAND2_X1   g00678(.A1(new_n933_), .A2(new_n886_), .ZN(new_n935_));
  INV_X1     g00679(.I(new_n935_), .ZN(new_n936_));
  NOR2_X1    g00680(.A1(new_n936_), .A2(new_n934_), .ZN(new_n937_));
  INV_X1     g00681(.I(new_n845_), .ZN(new_n938_));
  OAI21_X1   g00682(.A1(new_n795_), .A2(new_n938_), .B(new_n844_), .ZN(new_n939_));
  XOR2_X1    g00683(.A1(new_n937_), .A2(new_n939_), .Z(new_n940_));
  INV_X1     g00684(.I(\b[12] ), .ZN(new_n941_));
  OAI22_X1   g00685(.A1(new_n277_), .A2(new_n941_), .B1(new_n852_), .B2(new_n262_), .ZN(new_n942_));
  AOI21_X1   g00686(.A1(\b[10] ), .A2(new_n283_), .B(new_n942_), .ZN(new_n943_));
  XOR2_X1    g00687(.A1(\b[11] ), .A2(\b[12] ), .Z(new_n944_));
  NOR3_X1    g00688(.A1(new_n779_), .A2(new_n780_), .A3(new_n667_), .ZN(new_n945_));
  OAI21_X1   g00689(.A1(new_n945_), .A2(\b[10] ), .B(\b[11] ), .ZN(new_n946_));
  OAI21_X1   g00690(.A1(new_n781_), .A2(\b[9] ), .B(\b[10] ), .ZN(new_n947_));
  AND2_X2    g00691(.A1(new_n946_), .A2(new_n947_), .Z(new_n948_));
  NOR2_X1    g00692(.A1(new_n948_), .A2(new_n944_), .ZN(new_n949_));
  INV_X1     g00693(.I(new_n944_), .ZN(new_n950_));
  NAND2_X1   g00694(.A1(new_n946_), .A2(new_n947_), .ZN(new_n951_));
  NOR2_X1    g00695(.A1(new_n951_), .A2(new_n950_), .ZN(new_n952_));
  NOR2_X1    g00696(.A1(new_n949_), .A2(new_n952_), .ZN(new_n953_));
  OAI21_X1   g00697(.A1(new_n953_), .A2(new_n279_), .B(new_n943_), .ZN(new_n954_));
  XOR2_X1    g00698(.A1(new_n954_), .A2(\a[2] ), .Z(new_n955_));
  NAND3_X1   g00699(.A1(new_n870_), .A2(new_n865_), .A3(new_n795_), .ZN(new_n956_));
  OAI21_X1   g00700(.A1(new_n866_), .A2(new_n864_), .B(new_n796_), .ZN(new_n957_));
  NAND2_X1   g00701(.A1(new_n957_), .A2(new_n956_), .ZN(new_n958_));
  INV_X1     g00702(.I(new_n789_), .ZN(new_n959_));
  AOI21_X1   g00703(.A1(new_n692_), .A2(new_n959_), .B(new_n791_), .ZN(new_n960_));
  XOR2_X1    g00704(.A1(new_n868_), .A2(new_n795_), .Z(new_n961_));
  NOR2_X1    g00705(.A1(new_n961_), .A2(new_n869_), .ZN(new_n962_));
  INV_X1     g00706(.I(new_n962_), .ZN(new_n963_));
  OAI21_X1   g00707(.A1(new_n960_), .A2(new_n958_), .B(new_n963_), .ZN(new_n964_));
  NAND2_X1   g00708(.A1(new_n964_), .A2(new_n955_), .ZN(new_n965_));
  INV_X1     g00709(.I(new_n955_), .ZN(new_n966_));
  AOI21_X1   g00710(.A1(new_n878_), .A2(new_n872_), .B(new_n962_), .ZN(new_n967_));
  NAND2_X1   g00711(.A1(new_n967_), .A2(new_n966_), .ZN(new_n968_));
  NAND2_X1   g00712(.A1(new_n965_), .A2(new_n968_), .ZN(new_n969_));
  XOR2_X1    g00713(.A1(new_n969_), .A2(new_n940_), .Z(\f[12] ));
  OAI21_X1   g00714(.A1(new_n967_), .A2(new_n966_), .B(new_n940_), .ZN(new_n971_));
  NAND2_X1   g00715(.A1(new_n971_), .A2(new_n968_), .ZN(new_n972_));
  OAI21_X1   g00716(.A1(new_n939_), .A2(new_n934_), .B(new_n935_), .ZN(new_n973_));
  INV_X1     g00717(.I(new_n973_), .ZN(new_n974_));
  OAI22_X1   g00718(.A1(new_n713_), .A2(new_n339_), .B1(new_n290_), .B2(new_n717_), .ZN(new_n975_));
  NOR4_X1    g00719(.A1(new_n816_), .A2(new_n817_), .A3(new_n276_), .A4(new_n808_), .ZN(new_n976_));
  NOR2_X1    g00720(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  OAI21_X1   g00721(.A1(new_n346_), .A2(new_n351_), .B(new_n724_), .ZN(new_n978_));
  AOI21_X1   g00722(.A1(new_n977_), .A2(new_n978_), .B(new_n722_), .ZN(new_n979_));
  NAND2_X1   g00723(.A1(new_n728_), .A2(new_n710_), .ZN(new_n980_));
  NAND3_X1   g00724(.A1(new_n980_), .A2(new_n816_), .A3(\b[4] ), .ZN(new_n981_));
  NAND2_X1   g00725(.A1(new_n732_), .A2(\b[3] ), .ZN(new_n982_));
  NAND4_X1   g00726(.A1(new_n631_), .A2(new_n809_), .A3(\b[2] ), .A4(new_n810_), .ZN(new_n983_));
  NAND3_X1   g00727(.A1(new_n983_), .A2(new_n981_), .A3(new_n982_), .ZN(new_n984_));
  NAND2_X1   g00728(.A1(new_n721_), .A2(new_n723_), .ZN(new_n985_));
  NAND2_X1   g00729(.A1(new_n816_), .A2(new_n985_), .ZN(new_n986_));
  NOR2_X1    g00730(.A1(new_n352_), .A2(new_n986_), .ZN(new_n987_));
  NOR3_X1    g00731(.A1(new_n987_), .A2(new_n984_), .A3(\a[11] ), .ZN(new_n988_));
  NOR2_X1    g00732(.A1(new_n979_), .A2(new_n988_), .ZN(new_n989_));
  NAND2_X1   g00733(.A1(\a[13] ), .A2(\a[14] ), .ZN(new_n990_));
  INV_X1     g00734(.I(new_n990_), .ZN(new_n991_));
  NOR2_X1    g00735(.A1(\a[13] ), .A2(\a[14] ), .ZN(new_n992_));
  OAI22_X1   g00736(.A1(new_n991_), .A2(new_n992_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n993_));
  INV_X1     g00737(.I(\a[13] ), .ZN(new_n994_));
  NOR3_X1    g00738(.A1(new_n994_), .A2(\a[11] ), .A3(\a[12] ), .ZN(new_n995_));
  NOR3_X1    g00739(.A1(new_n722_), .A2(new_n895_), .A3(\a[13] ), .ZN(new_n996_));
  NOR2_X1    g00740(.A1(new_n996_), .A2(new_n995_), .ZN(new_n997_));
  OAI22_X1   g00741(.A1(new_n993_), .A2(new_n275_), .B1(new_n258_), .B2(new_n997_), .ZN(new_n998_));
  XNOR2_X1   g00742(.A1(\a[13] ), .A2(\a[14] ), .ZN(new_n999_));
  NOR3_X1    g00743(.A1(new_n898_), .A2(new_n999_), .A3(new_n313_), .ZN(new_n1000_));
  OAI21_X1   g00744(.A1(new_n998_), .A2(new_n1000_), .B(\a[14] ), .ZN(new_n1001_));
  INV_X1     g00745(.I(\a[14] ), .ZN(new_n1002_));
  NAND2_X1   g00746(.A1(new_n722_), .A2(\a[12] ), .ZN(new_n1003_));
  NAND2_X1   g00747(.A1(new_n895_), .A2(\a[11] ), .ZN(new_n1004_));
  INV_X1     g00748(.I(new_n992_), .ZN(new_n1005_));
  AOI22_X1   g00749(.A1(new_n990_), .A2(new_n1005_), .B1(new_n1003_), .B2(new_n1004_), .ZN(new_n1006_));
  NAND3_X1   g00750(.A1(new_n722_), .A2(new_n895_), .A3(\a[13] ), .ZN(new_n1007_));
  NAND3_X1   g00751(.A1(new_n994_), .A2(\a[11] ), .A3(\a[12] ), .ZN(new_n1008_));
  NAND2_X1   g00752(.A1(new_n1007_), .A2(new_n1008_), .ZN(new_n1009_));
  AOI22_X1   g00753(.A1(new_n1006_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n1009_), .ZN(new_n1010_));
  NAND2_X1   g00754(.A1(new_n994_), .A2(\a[14] ), .ZN(new_n1011_));
  NAND2_X1   g00755(.A1(new_n1002_), .A2(\a[13] ), .ZN(new_n1012_));
  AOI22_X1   g00756(.A1(new_n1003_), .A2(new_n1004_), .B1(new_n1011_), .B2(new_n1012_), .ZN(new_n1013_));
  NAND2_X1   g00757(.A1(new_n1013_), .A2(new_n263_), .ZN(new_n1014_));
  NAND3_X1   g00758(.A1(new_n1010_), .A2(new_n1002_), .A3(new_n1014_), .ZN(new_n1015_));
  NAND2_X1   g00759(.A1(new_n900_), .A2(\a[14] ), .ZN(new_n1016_));
  NAND3_X1   g00760(.A1(new_n1001_), .A2(new_n1015_), .A3(new_n1016_), .ZN(new_n1017_));
  NAND2_X1   g00761(.A1(new_n1010_), .A2(new_n1014_), .ZN(new_n1018_));
  NAND3_X1   g00762(.A1(new_n1018_), .A2(\a[14] ), .A3(new_n900_), .ZN(new_n1019_));
  NAND2_X1   g00763(.A1(new_n1017_), .A2(new_n1019_), .ZN(new_n1020_));
  NAND2_X1   g00764(.A1(new_n1020_), .A2(new_n989_), .ZN(new_n1021_));
  OAI21_X1   g00765(.A1(new_n987_), .A2(new_n984_), .B(\a[11] ), .ZN(new_n1022_));
  AOI22_X1   g00766(.A1(new_n729_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n732_), .ZN(new_n1023_));
  NAND4_X1   g00767(.A1(new_n978_), .A2(new_n1023_), .A3(new_n722_), .A4(new_n983_), .ZN(new_n1024_));
  NAND2_X1   g00768(.A1(new_n1022_), .A2(new_n1024_), .ZN(new_n1025_));
  NAND3_X1   g00769(.A1(new_n1025_), .A2(new_n1017_), .A3(new_n1019_), .ZN(new_n1026_));
  OAI21_X1   g00770(.A1(new_n825_), .A2(new_n912_), .B(new_n901_), .ZN(new_n1027_));
  AOI21_X1   g00771(.A1(new_n1021_), .A2(new_n1026_), .B(new_n1027_), .ZN(new_n1028_));
  AOI21_X1   g00772(.A1(new_n1017_), .A2(new_n1019_), .B(new_n1025_), .ZN(new_n1029_));
  NOR2_X1    g00773(.A1(new_n1020_), .A2(new_n989_), .ZN(new_n1030_));
  AOI21_X1   g00774(.A1(new_n837_), .A2(new_n909_), .B(new_n911_), .ZN(new_n1031_));
  NOR3_X1    g00775(.A1(new_n1031_), .A2(new_n1030_), .A3(new_n1029_), .ZN(new_n1032_));
  OAI22_X1   g00776(.A1(new_n610_), .A2(new_n471_), .B1(new_n438_), .B2(new_n612_), .ZN(new_n1033_));
  NOR2_X1    g00777(.A1(new_n917_), .A2(new_n377_), .ZN(new_n1034_));
  NOR2_X1    g00778(.A1(new_n1034_), .A2(new_n1033_), .ZN(new_n1035_));
  INV_X1     g00779(.I(new_n1035_), .ZN(new_n1036_));
  AOI21_X1   g00780(.A1(new_n482_), .A2(new_n483_), .B(new_n471_), .ZN(new_n1037_));
  NOR3_X1    g00781(.A1(new_n475_), .A2(\b[7] ), .A3(new_n476_), .ZN(new_n1038_));
  NOR3_X1    g00782(.A1(new_n1037_), .A2(new_n1038_), .A3(new_n624_), .ZN(new_n1039_));
  OAI21_X1   g00783(.A1(new_n1039_), .A2(new_n1036_), .B(\a[8] ), .ZN(new_n1040_));
  NAND3_X1   g00784(.A1(new_n484_), .A2(new_n477_), .A3(new_n618_), .ZN(new_n1041_));
  NAND3_X1   g00785(.A1(new_n1041_), .A2(new_n488_), .A3(new_n1035_), .ZN(new_n1042_));
  NAND2_X1   g00786(.A1(new_n1040_), .A2(new_n1042_), .ZN(new_n1043_));
  INV_X1     g00787(.I(new_n1043_), .ZN(new_n1044_));
  NOR3_X1    g00788(.A1(new_n1044_), .A2(new_n1028_), .A3(new_n1032_), .ZN(new_n1045_));
  NOR2_X1    g00789(.A1(new_n1028_), .A2(new_n1032_), .ZN(new_n1046_));
  NOR2_X1    g00790(.A1(new_n1046_), .A2(new_n1043_), .ZN(new_n1047_));
  NOR2_X1    g00791(.A1(new_n1045_), .A2(new_n1047_), .ZN(new_n1048_));
  OAI21_X1   g00792(.A1(new_n928_), .A2(new_n925_), .B(new_n914_), .ZN(new_n1049_));
  NAND2_X1   g00793(.A1(new_n1049_), .A2(new_n929_), .ZN(new_n1050_));
  NAND2_X1   g00794(.A1(new_n1048_), .A2(new_n1050_), .ZN(new_n1051_));
  NOR2_X1    g00795(.A1(new_n923_), .A2(new_n921_), .ZN(new_n1052_));
  NAND2_X1   g00796(.A1(new_n910_), .A2(new_n913_), .ZN(new_n1053_));
  AOI21_X1   g00797(.A1(new_n923_), .A2(new_n921_), .B(new_n1053_), .ZN(new_n1054_));
  NOR2_X1    g00798(.A1(new_n1054_), .A2(new_n1052_), .ZN(new_n1055_));
  OAI21_X1   g00799(.A1(new_n1045_), .A2(new_n1047_), .B(new_n1055_), .ZN(new_n1056_));
  NAND2_X1   g00800(.A1(new_n1056_), .A2(new_n1051_), .ZN(new_n1057_));
  NAND2_X1   g00801(.A1(new_n781_), .A2(new_n785_), .ZN(new_n1058_));
  OAI21_X1   g00802(.A1(new_n781_), .A2(new_n782_), .B(new_n1058_), .ZN(new_n1059_));
  AOI22_X1   g00803(.A1(new_n800_), .A2(\b[9] ), .B1(\b[10] ), .B2(new_n333_), .ZN(new_n1060_));
  OAI21_X1   g00804(.A1(new_n577_), .A2(new_n392_), .B(new_n1060_), .ZN(new_n1061_));
  AOI21_X1   g00805(.A1(new_n1059_), .A2(new_n330_), .B(new_n1061_), .ZN(new_n1062_));
  XOR2_X1    g00806(.A1(new_n1062_), .A2(new_n312_), .Z(new_n1063_));
  NAND2_X1   g00807(.A1(new_n1057_), .A2(new_n1063_), .ZN(new_n1064_));
  OR2_X2     g00808(.A1(new_n1057_), .A2(new_n1063_), .Z(new_n1065_));
  NAND2_X1   g00809(.A1(new_n1065_), .A2(new_n1064_), .ZN(new_n1066_));
  NAND2_X1   g00810(.A1(new_n974_), .A2(new_n1066_), .ZN(new_n1067_));
  NAND3_X1   g00811(.A1(new_n973_), .A2(new_n1064_), .A3(new_n1065_), .ZN(new_n1068_));
  NAND2_X1   g00812(.A1(new_n1067_), .A2(new_n1068_), .ZN(new_n1069_));
  INV_X1     g00813(.I(\b[13] ), .ZN(new_n1070_));
  OAI22_X1   g00814(.A1(new_n277_), .A2(new_n1070_), .B1(new_n941_), .B2(new_n262_), .ZN(new_n1071_));
  AOI21_X1   g00815(.A1(\b[11] ), .A2(new_n283_), .B(new_n1071_), .ZN(new_n1072_));
  AOI21_X1   g00816(.A1(new_n951_), .A2(\b[12] ), .B(new_n852_), .ZN(new_n1073_));
  NOR2_X1    g00817(.A1(new_n951_), .A2(\b[12] ), .ZN(new_n1074_));
  NAND3_X1   g00818(.A1(new_n946_), .A2(new_n947_), .A3(new_n1070_), .ZN(new_n1075_));
  INV_X1     g00819(.I(new_n1075_), .ZN(new_n1076_));
  NOR2_X1    g00820(.A1(new_n948_), .A2(new_n1070_), .ZN(new_n1077_));
  OAI22_X1   g00821(.A1(new_n1077_), .A2(new_n1076_), .B1(new_n1073_), .B2(new_n1074_), .ZN(new_n1078_));
  NOR2_X1    g00822(.A1(new_n1073_), .A2(new_n1074_), .ZN(new_n1079_));
  NOR2_X1    g00823(.A1(new_n1077_), .A2(new_n1076_), .ZN(new_n1080_));
  NAND2_X1   g00824(.A1(new_n1080_), .A2(new_n1079_), .ZN(new_n1081_));
  NAND2_X1   g00825(.A1(new_n1081_), .A2(new_n1078_), .ZN(new_n1082_));
  OAI21_X1   g00826(.A1(new_n1082_), .A2(new_n279_), .B(new_n1072_), .ZN(new_n1083_));
  XOR2_X1    g00827(.A1(new_n1083_), .A2(\a[2] ), .Z(new_n1084_));
  INV_X1     g00828(.I(new_n1084_), .ZN(new_n1085_));
  NAND2_X1   g00829(.A1(new_n1069_), .A2(new_n1085_), .ZN(new_n1086_));
  NOR2_X1    g00830(.A1(new_n1069_), .A2(new_n1085_), .ZN(new_n1087_));
  INV_X1     g00831(.I(new_n1087_), .ZN(new_n1088_));
  NAND2_X1   g00832(.A1(new_n1088_), .A2(new_n1086_), .ZN(new_n1089_));
  XOR2_X1    g00833(.A1(new_n972_), .A2(new_n1089_), .Z(\f[13] ));
  NAND3_X1   g00834(.A1(new_n971_), .A2(new_n968_), .A3(new_n1086_), .ZN(new_n1091_));
  NAND2_X1   g00835(.A1(new_n1091_), .A2(new_n1088_), .ZN(new_n1092_));
  INV_X1     g00836(.I(\b[14] ), .ZN(new_n1093_));
  OAI22_X1   g00837(.A1(new_n277_), .A2(new_n1093_), .B1(new_n1070_), .B2(new_n262_), .ZN(new_n1094_));
  AOI21_X1   g00838(.A1(\b[12] ), .A2(new_n283_), .B(new_n1094_), .ZN(new_n1095_));
  AOI21_X1   g00839(.A1(new_n1075_), .A2(\b[12] ), .B(\b[11] ), .ZN(new_n1096_));
  AOI21_X1   g00840(.A1(new_n951_), .A2(\b[13] ), .B(\b[12] ), .ZN(new_n1097_));
  NOR2_X1    g00841(.A1(new_n1096_), .A2(new_n1097_), .ZN(new_n1098_));
  XNOR2_X1   g00842(.A1(\b[13] ), .A2(\b[14] ), .ZN(new_n1099_));
  NOR2_X1    g00843(.A1(new_n1098_), .A2(new_n1099_), .ZN(new_n1100_));
  XOR2_X1    g00844(.A1(\b[13] ), .A2(\b[14] ), .Z(new_n1101_));
  NOR3_X1    g00845(.A1(new_n1096_), .A2(new_n1097_), .A3(new_n1101_), .ZN(new_n1102_));
  NOR2_X1    g00846(.A1(new_n1100_), .A2(new_n1102_), .ZN(new_n1103_));
  OAI21_X1   g00847(.A1(new_n1103_), .A2(new_n279_), .B(new_n1095_), .ZN(new_n1104_));
  XOR2_X1    g00848(.A1(new_n1104_), .A2(\a[2] ), .Z(new_n1105_));
  OAI22_X1   g00849(.A1(new_n321_), .A2(new_n852_), .B1(new_n325_), .B2(new_n776_), .ZN(new_n1106_));
  AOI21_X1   g00850(.A1(\b[9] ), .A2(new_n602_), .B(new_n1106_), .ZN(new_n1107_));
  OAI21_X1   g00851(.A1(new_n859_), .A2(new_n318_), .B(new_n1107_), .ZN(new_n1108_));
  XOR2_X1    g00852(.A1(new_n1108_), .A2(\a[5] ), .Z(new_n1109_));
  NAND2_X1   g00853(.A1(new_n1046_), .A2(new_n1043_), .ZN(new_n1110_));
  OAI22_X1   g00854(.A1(new_n1054_), .A2(new_n1052_), .B1(new_n1046_), .B2(new_n1043_), .ZN(new_n1111_));
  OAI22_X1   g00855(.A1(new_n610_), .A2(new_n577_), .B1(new_n471_), .B2(new_n612_), .ZN(new_n1112_));
  NOR2_X1    g00856(.A1(new_n917_), .A2(new_n438_), .ZN(new_n1113_));
  NOR2_X1    g00857(.A1(new_n1113_), .A2(new_n1112_), .ZN(new_n1114_));
  INV_X1     g00858(.I(new_n1114_), .ZN(new_n1115_));
  AOI21_X1   g00859(.A1(new_n798_), .A2(new_n585_), .B(new_n624_), .ZN(new_n1116_));
  OAI21_X1   g00860(.A1(new_n1116_), .A2(new_n1115_), .B(\a[8] ), .ZN(new_n1117_));
  OAI21_X1   g00861(.A1(new_n586_), .A2(new_n584_), .B(new_n618_), .ZN(new_n1118_));
  NAND3_X1   g00862(.A1(new_n1118_), .A2(new_n488_), .A3(new_n1114_), .ZN(new_n1119_));
  OAI21_X1   g00863(.A1(new_n1027_), .A2(new_n1030_), .B(new_n1021_), .ZN(new_n1120_));
  NAND3_X1   g00864(.A1(new_n1120_), .A2(new_n1117_), .A3(new_n1119_), .ZN(new_n1121_));
  AOI21_X1   g00865(.A1(new_n1118_), .A2(new_n1114_), .B(new_n488_), .ZN(new_n1122_));
  NOR3_X1    g00866(.A1(new_n1116_), .A2(\a[8] ), .A3(new_n1115_), .ZN(new_n1123_));
  AOI21_X1   g00867(.A1(new_n1031_), .A2(new_n1026_), .B(new_n1029_), .ZN(new_n1124_));
  OAI21_X1   g00868(.A1(new_n1122_), .A2(new_n1123_), .B(new_n1124_), .ZN(new_n1125_));
  NOR3_X1    g00869(.A1(new_n816_), .A2(new_n817_), .A3(new_n808_), .ZN(new_n1126_));
  INV_X1     g00870(.I(new_n1126_), .ZN(new_n1127_));
  AOI22_X1   g00871(.A1(new_n729_), .A2(\b[5] ), .B1(\b[4] ), .B2(new_n732_), .ZN(new_n1128_));
  OAI21_X1   g00872(.A1(new_n290_), .A2(new_n1127_), .B(new_n1128_), .ZN(new_n1129_));
  NOR3_X1    g00873(.A1(new_n380_), .A2(new_n381_), .A3(new_n986_), .ZN(new_n1130_));
  OAI21_X1   g00874(.A1(new_n1130_), .A2(new_n1129_), .B(\a[11] ), .ZN(new_n1131_));
  NAND2_X1   g00875(.A1(new_n1126_), .A2(\b[3] ), .ZN(new_n1132_));
  AND2_X2    g00876(.A1(new_n1132_), .A2(new_n1128_), .Z(new_n1133_));
  NAND3_X1   g00877(.A1(new_n565_), .A2(new_n379_), .A3(new_n724_), .ZN(new_n1134_));
  NAND3_X1   g00878(.A1(new_n1134_), .A2(new_n1133_), .A3(new_n722_), .ZN(new_n1135_));
  NAND2_X1   g00879(.A1(new_n1013_), .A2(new_n554_), .ZN(new_n1136_));
  NOR2_X1    g00880(.A1(new_n991_), .A2(new_n992_), .ZN(new_n1137_));
  NOR3_X1    g00881(.A1(new_n898_), .A2(new_n1137_), .A3(new_n276_), .ZN(new_n1138_));
  NOR2_X1    g00882(.A1(new_n997_), .A2(new_n275_), .ZN(new_n1139_));
  NAND2_X1   g00883(.A1(new_n1003_), .A2(new_n1004_), .ZN(new_n1140_));
  AOI21_X1   g00884(.A1(new_n994_), .A2(\a[14] ), .B(\a[11] ), .ZN(new_n1141_));
  OAI21_X1   g00885(.A1(new_n994_), .A2(\a[14] ), .B(\a[11] ), .ZN(new_n1142_));
  INV_X1     g00886(.I(new_n1142_), .ZN(new_n1143_));
  NOR4_X1    g00887(.A1(new_n1140_), .A2(new_n1143_), .A3(new_n258_), .A4(new_n1141_), .ZN(new_n1144_));
  NOR3_X1    g00888(.A1(new_n1144_), .A2(new_n1138_), .A3(new_n1139_), .ZN(new_n1145_));
  AOI21_X1   g00889(.A1(new_n1145_), .A2(new_n1136_), .B(new_n1002_), .ZN(new_n1146_));
  INV_X1     g00890(.I(new_n1136_), .ZN(new_n1147_));
  OAI22_X1   g00891(.A1(new_n993_), .A2(new_n276_), .B1(new_n275_), .B2(new_n997_), .ZN(new_n1148_));
  NOR4_X1    g00892(.A1(new_n1147_), .A2(new_n1148_), .A3(\a[14] ), .A4(new_n1144_), .ZN(new_n1149_));
  NAND4_X1   g00893(.A1(new_n1010_), .A2(new_n900_), .A3(\a[14] ), .A4(new_n1014_), .ZN(new_n1150_));
  OAI21_X1   g00894(.A1(new_n1146_), .A2(new_n1149_), .B(new_n1150_), .ZN(new_n1151_));
  NOR2_X1    g00895(.A1(new_n998_), .A2(new_n1000_), .ZN(new_n1152_));
  NAND2_X1   g00896(.A1(new_n1006_), .A2(\b[2] ), .ZN(new_n1153_));
  NAND2_X1   g00897(.A1(new_n1009_), .A2(\b[1] ), .ZN(new_n1154_));
  INV_X1     g00898(.I(new_n1141_), .ZN(new_n1155_));
  NAND4_X1   g00899(.A1(new_n898_), .A2(new_n1155_), .A3(\b[0] ), .A4(new_n1142_), .ZN(new_n1156_));
  NAND3_X1   g00900(.A1(new_n1153_), .A2(new_n1156_), .A3(new_n1154_), .ZN(new_n1157_));
  NOR2_X1    g00901(.A1(new_n1157_), .A2(new_n1147_), .ZN(new_n1158_));
  NAND4_X1   g00902(.A1(new_n1158_), .A2(\a[14] ), .A3(new_n1152_), .A4(new_n900_), .ZN(new_n1159_));
  NAND4_X1   g00903(.A1(new_n1131_), .A2(new_n1135_), .A3(new_n1151_), .A4(new_n1159_), .ZN(new_n1160_));
  AOI21_X1   g00904(.A1(new_n1134_), .A2(new_n1133_), .B(new_n722_), .ZN(new_n1161_));
  NOR3_X1    g00905(.A1(new_n1130_), .A2(\a[11] ), .A3(new_n1129_), .ZN(new_n1162_));
  OAI21_X1   g00906(.A1(new_n1157_), .A2(new_n1147_), .B(\a[14] ), .ZN(new_n1163_));
  NAND3_X1   g00907(.A1(new_n1145_), .A2(new_n1002_), .A3(new_n1136_), .ZN(new_n1164_));
  NOR4_X1    g00908(.A1(new_n998_), .A2(new_n1002_), .A3(new_n899_), .A4(new_n1000_), .ZN(new_n1165_));
  AOI21_X1   g00909(.A1(new_n1163_), .A2(new_n1164_), .B(new_n1165_), .ZN(new_n1166_));
  NOR3_X1    g00910(.A1(new_n1146_), .A2(new_n1149_), .A3(new_n1150_), .ZN(new_n1167_));
  OAI22_X1   g00911(.A1(new_n1162_), .A2(new_n1161_), .B1(new_n1166_), .B2(new_n1167_), .ZN(new_n1168_));
  NAND2_X1   g00912(.A1(new_n1168_), .A2(new_n1160_), .ZN(new_n1169_));
  INV_X1     g00913(.I(new_n1169_), .ZN(new_n1170_));
  NAND3_X1   g00914(.A1(new_n1125_), .A2(new_n1121_), .A3(new_n1170_), .ZN(new_n1171_));
  NOR3_X1    g00915(.A1(new_n1124_), .A2(new_n1123_), .A3(new_n1122_), .ZN(new_n1172_));
  AOI21_X1   g00916(.A1(new_n1117_), .A2(new_n1119_), .B(new_n1120_), .ZN(new_n1173_));
  OAI21_X1   g00917(.A1(new_n1173_), .A2(new_n1172_), .B(new_n1169_), .ZN(new_n1174_));
  NAND4_X1   g00918(.A1(new_n1111_), .A2(new_n1110_), .A3(new_n1171_), .A4(new_n1174_), .ZN(new_n1175_));
  OAI21_X1   g00919(.A1(new_n1055_), .A2(new_n1047_), .B(new_n1110_), .ZN(new_n1176_));
  NAND2_X1   g00920(.A1(new_n1174_), .A2(new_n1171_), .ZN(new_n1177_));
  NAND2_X1   g00921(.A1(new_n1176_), .A2(new_n1177_), .ZN(new_n1178_));
  NAND2_X1   g00922(.A1(new_n1178_), .A2(new_n1175_), .ZN(new_n1179_));
  XOR2_X1    g00923(.A1(new_n1109_), .A2(new_n1179_), .Z(new_n1180_));
  INV_X1     g00924(.I(new_n1064_), .ZN(new_n1181_));
  AOI21_X1   g00925(.A1(new_n973_), .A2(new_n1065_), .B(new_n1181_), .ZN(new_n1182_));
  INV_X1     g00926(.I(new_n1182_), .ZN(new_n1183_));
  NAND2_X1   g00927(.A1(new_n1183_), .A2(new_n1180_), .ZN(new_n1184_));
  INV_X1     g00928(.I(new_n1180_), .ZN(new_n1185_));
  NAND2_X1   g00929(.A1(new_n1185_), .A2(new_n1182_), .ZN(new_n1186_));
  NAND2_X1   g00930(.A1(new_n1184_), .A2(new_n1186_), .ZN(new_n1187_));
  XOR2_X1    g00931(.A1(new_n1187_), .A2(new_n1105_), .Z(new_n1188_));
  XOR2_X1    g00932(.A1(new_n1092_), .A2(new_n1188_), .Z(\f[14] ));
  INV_X1     g00933(.I(new_n1109_), .ZN(new_n1190_));
  OAI21_X1   g00934(.A1(new_n1182_), .A2(new_n1190_), .B(new_n1179_), .ZN(new_n1191_));
  NAND2_X1   g00935(.A1(new_n1182_), .A2(new_n1190_), .ZN(new_n1192_));
  NAND2_X1   g00936(.A1(new_n1191_), .A2(new_n1192_), .ZN(new_n1193_));
  INV_X1     g00937(.I(new_n953_), .ZN(new_n1194_));
  AOI22_X1   g00938(.A1(new_n800_), .A2(\b[11] ), .B1(\b[12] ), .B2(new_n333_), .ZN(new_n1195_));
  OAI21_X1   g00939(.A1(new_n776_), .A2(new_n392_), .B(new_n1195_), .ZN(new_n1196_));
  AOI21_X1   g00940(.A1(new_n1194_), .A2(new_n330_), .B(new_n1196_), .ZN(new_n1197_));
  XOR2_X1    g00941(.A1(new_n1197_), .A2(new_n312_), .Z(new_n1198_));
  NAND4_X1   g00942(.A1(new_n898_), .A2(new_n1155_), .A3(\b[1] ), .A4(new_n1142_), .ZN(new_n1199_));
  AOI21_X1   g00943(.A1(new_n1007_), .A2(new_n1008_), .B(new_n276_), .ZN(new_n1200_));
  AOI21_X1   g00944(.A1(new_n1006_), .A2(\b[3] ), .B(new_n1200_), .ZN(new_n1201_));
  NAND3_X1   g00945(.A1(new_n1013_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n1202_));
  NAND3_X1   g00946(.A1(new_n1201_), .A2(new_n1202_), .A3(new_n1199_), .ZN(new_n1203_));
  NAND2_X1   g00947(.A1(new_n1203_), .A2(\a[14] ), .ZN(new_n1204_));
  NAND4_X1   g00948(.A1(new_n1201_), .A2(new_n1202_), .A3(new_n1002_), .A4(new_n1199_), .ZN(new_n1205_));
  XNOR2_X1   g00949(.A1(\a[14] ), .A2(\a[15] ), .ZN(new_n1206_));
  NOR2_X1    g00950(.A1(new_n1206_), .A2(new_n258_), .ZN(new_n1207_));
  AOI21_X1   g00951(.A1(new_n1204_), .A2(new_n1205_), .B(new_n1207_), .ZN(new_n1208_));
  NOR2_X1    g00952(.A1(new_n993_), .A2(new_n290_), .ZN(new_n1209_));
  NOR4_X1    g00953(.A1(new_n298_), .A2(new_n295_), .A3(new_n898_), .A4(new_n999_), .ZN(new_n1210_));
  NOR3_X1    g00954(.A1(new_n1210_), .A2(new_n1209_), .A3(new_n1200_), .ZN(new_n1211_));
  AOI21_X1   g00955(.A1(new_n1211_), .A2(new_n1199_), .B(new_n1002_), .ZN(new_n1212_));
  INV_X1     g00956(.I(new_n1205_), .ZN(new_n1213_));
  INV_X1     g00957(.I(new_n1207_), .ZN(new_n1214_));
  NOR3_X1    g00958(.A1(new_n1212_), .A2(new_n1213_), .A3(new_n1214_), .ZN(new_n1215_));
  NOR3_X1    g00959(.A1(new_n1215_), .A2(new_n1208_), .A3(new_n1167_), .ZN(new_n1216_));
  OAI21_X1   g00960(.A1(new_n1212_), .A2(new_n1213_), .B(new_n1214_), .ZN(new_n1217_));
  NAND3_X1   g00961(.A1(new_n1204_), .A2(new_n1205_), .A3(new_n1207_), .ZN(new_n1218_));
  AOI21_X1   g00962(.A1(new_n1217_), .A2(new_n1218_), .B(new_n1159_), .ZN(new_n1219_));
  NOR2_X1    g00963(.A1(new_n1216_), .A2(new_n1219_), .ZN(new_n1220_));
  INV_X1     g00964(.I(new_n1220_), .ZN(new_n1221_));
  OAI22_X1   g00965(.A1(new_n713_), .A2(new_n438_), .B1(new_n377_), .B2(new_n717_), .ZN(new_n1222_));
  AOI21_X1   g00966(.A1(\b[4] ), .A2(new_n1126_), .B(new_n1222_), .ZN(new_n1223_));
  OAI21_X1   g00967(.A1(new_n450_), .A2(new_n986_), .B(new_n1223_), .ZN(new_n1224_));
  XOR2_X1    g00968(.A1(new_n1224_), .A2(\a[11] ), .Z(new_n1225_));
  INV_X1     g00969(.I(new_n1225_), .ZN(new_n1226_));
  INV_X1     g00970(.I(new_n1160_), .ZN(new_n1227_));
  AOI21_X1   g00971(.A1(new_n1120_), .A2(new_n1168_), .B(new_n1227_), .ZN(new_n1228_));
  NOR2_X1    g00972(.A1(new_n1228_), .A2(new_n1226_), .ZN(new_n1229_));
  INV_X1     g00973(.I(new_n1168_), .ZN(new_n1230_));
  OAI21_X1   g00974(.A1(new_n1124_), .A2(new_n1230_), .B(new_n1160_), .ZN(new_n1231_));
  NOR2_X1    g00975(.A1(new_n1231_), .A2(new_n1225_), .ZN(new_n1232_));
  NOR3_X1    g00976(.A1(new_n1229_), .A2(new_n1232_), .A3(new_n1221_), .ZN(new_n1233_));
  NAND2_X1   g00977(.A1(new_n1231_), .A2(new_n1225_), .ZN(new_n1234_));
  NAND2_X1   g00978(.A1(new_n1228_), .A2(new_n1226_), .ZN(new_n1235_));
  AOI21_X1   g00979(.A1(new_n1235_), .A2(new_n1234_), .B(new_n1220_), .ZN(new_n1236_));
  NOR2_X1    g00980(.A1(new_n1236_), .A2(new_n1233_), .ZN(new_n1237_));
  OAI21_X1   g00981(.A1(new_n660_), .A2(new_n661_), .B(new_n674_), .ZN(new_n1238_));
  NAND2_X1   g00982(.A1(new_n670_), .A2(new_n662_), .ZN(new_n1239_));
  NAND2_X1   g00983(.A1(new_n1239_), .A2(new_n1238_), .ZN(new_n1240_));
  AOI22_X1   g00984(.A1(new_n518_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n636_), .ZN(new_n1241_));
  OAI21_X1   g00985(.A1(new_n471_), .A2(new_n917_), .B(new_n1241_), .ZN(new_n1242_));
  INV_X1     g00986(.I(new_n1242_), .ZN(new_n1243_));
  OAI21_X1   g00987(.A1(new_n1240_), .A2(new_n624_), .B(new_n1243_), .ZN(new_n1244_));
  NAND2_X1   g00988(.A1(new_n1244_), .A2(\a[8] ), .ZN(new_n1245_));
  NAND2_X1   g00989(.A1(new_n676_), .A2(new_n618_), .ZN(new_n1246_));
  NAND3_X1   g00990(.A1(new_n1246_), .A2(new_n488_), .A3(new_n1243_), .ZN(new_n1247_));
  NAND2_X1   g00991(.A1(new_n1245_), .A2(new_n1247_), .ZN(new_n1248_));
  XOR2_X1    g00992(.A1(new_n1169_), .A2(new_n1124_), .Z(new_n1249_));
  NAND3_X1   g00993(.A1(new_n1249_), .A2(new_n1117_), .A3(new_n1119_), .ZN(new_n1250_));
  AOI21_X1   g00994(.A1(new_n1175_), .A2(new_n1250_), .B(new_n1248_), .ZN(new_n1251_));
  INV_X1     g00995(.I(new_n1251_), .ZN(new_n1252_));
  NAND3_X1   g00996(.A1(new_n1175_), .A2(new_n1248_), .A3(new_n1250_), .ZN(new_n1253_));
  NAND3_X1   g00997(.A1(new_n1252_), .A2(new_n1253_), .A3(new_n1237_), .ZN(new_n1254_));
  NAND3_X1   g00998(.A1(new_n1235_), .A2(new_n1234_), .A3(new_n1220_), .ZN(new_n1255_));
  OAI21_X1   g00999(.A1(new_n1229_), .A2(new_n1232_), .B(new_n1221_), .ZN(new_n1256_));
  NAND2_X1   g01000(.A1(new_n1256_), .A2(new_n1255_), .ZN(new_n1257_));
  INV_X1     g01001(.I(new_n1248_), .ZN(new_n1258_));
  OAI21_X1   g01002(.A1(new_n1176_), .A2(new_n1177_), .B(new_n1250_), .ZN(new_n1259_));
  NOR2_X1    g01003(.A1(new_n1259_), .A2(new_n1258_), .ZN(new_n1260_));
  OAI21_X1   g01004(.A1(new_n1260_), .A2(new_n1251_), .B(new_n1257_), .ZN(new_n1261_));
  NAND2_X1   g01005(.A1(new_n1254_), .A2(new_n1261_), .ZN(new_n1262_));
  NOR2_X1    g01006(.A1(new_n1262_), .A2(new_n1198_), .ZN(new_n1263_));
  INV_X1     g01007(.I(new_n1263_), .ZN(new_n1264_));
  NAND2_X1   g01008(.A1(new_n1262_), .A2(new_n1198_), .ZN(new_n1265_));
  NAND2_X1   g01009(.A1(new_n1264_), .A2(new_n1265_), .ZN(new_n1266_));
  XNOR2_X1   g01010(.A1(new_n1266_), .A2(new_n1193_), .ZN(new_n1267_));
  INV_X1     g01011(.I(\b[15] ), .ZN(new_n1268_));
  OAI22_X1   g01012(.A1(new_n277_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n262_), .ZN(new_n1269_));
  AOI21_X1   g01013(.A1(\b[13] ), .A2(new_n283_), .B(new_n1269_), .ZN(new_n1270_));
  OAI21_X1   g01014(.A1(new_n1096_), .A2(new_n1097_), .B(new_n1070_), .ZN(new_n1271_));
  NOR3_X1    g01015(.A1(new_n1096_), .A2(new_n1097_), .A3(new_n1070_), .ZN(new_n1272_));
  NAND2_X1   g01016(.A1(new_n1272_), .A2(new_n1093_), .ZN(new_n1273_));
  OAI21_X1   g01017(.A1(new_n1093_), .A2(new_n1271_), .B(new_n1273_), .ZN(new_n1274_));
  XOR2_X1    g01018(.A1(new_n1274_), .A2(new_n1268_), .Z(new_n1275_));
  OAI21_X1   g01019(.A1(new_n1275_), .A2(new_n279_), .B(new_n1270_), .ZN(new_n1276_));
  XOR2_X1    g01020(.A1(new_n1276_), .A2(\a[2] ), .Z(new_n1277_));
  INV_X1     g01021(.I(new_n1105_), .ZN(new_n1278_));
  XOR2_X1    g01022(.A1(new_n1187_), .A2(new_n1278_), .Z(new_n1279_));
  AOI21_X1   g01023(.A1(new_n1091_), .A2(new_n1088_), .B(new_n1279_), .ZN(new_n1280_));
  AOI21_X1   g01024(.A1(new_n1184_), .A2(new_n1186_), .B(new_n1278_), .ZN(new_n1281_));
  OAI21_X1   g01025(.A1(new_n1280_), .A2(new_n1281_), .B(new_n1277_), .ZN(new_n1282_));
  INV_X1     g01026(.I(new_n1277_), .ZN(new_n1283_));
  NOR2_X1    g01027(.A1(new_n964_), .A2(new_n955_), .ZN(new_n1284_));
  INV_X1     g01028(.I(new_n940_), .ZN(new_n1285_));
  AOI21_X1   g01029(.A1(new_n964_), .A2(new_n955_), .B(new_n1285_), .ZN(new_n1286_));
  INV_X1     g01030(.I(new_n1086_), .ZN(new_n1287_));
  NOR3_X1    g01031(.A1(new_n1286_), .A2(new_n1284_), .A3(new_n1287_), .ZN(new_n1288_));
  OAI21_X1   g01032(.A1(new_n1288_), .A2(new_n1087_), .B(new_n1188_), .ZN(new_n1289_));
  INV_X1     g01033(.I(new_n1281_), .ZN(new_n1290_));
  NAND3_X1   g01034(.A1(new_n1289_), .A2(new_n1283_), .A3(new_n1290_), .ZN(new_n1291_));
  NAND2_X1   g01035(.A1(new_n1291_), .A2(new_n1282_), .ZN(new_n1292_));
  XOR2_X1    g01036(.A1(new_n1292_), .A2(new_n1267_), .Z(\f[15] ));
  NOR3_X1    g01037(.A1(new_n1280_), .A2(new_n1277_), .A3(new_n1281_), .ZN(new_n1294_));
  AOI21_X1   g01038(.A1(new_n1267_), .A2(new_n1282_), .B(new_n1294_), .ZN(new_n1295_));
  INV_X1     g01039(.I(\b[16] ), .ZN(new_n1296_));
  OAI22_X1   g01040(.A1(new_n277_), .A2(new_n1296_), .B1(new_n1268_), .B2(new_n262_), .ZN(new_n1297_));
  AOI21_X1   g01041(.A1(\b[14] ), .A2(new_n283_), .B(new_n1297_), .ZN(new_n1298_));
  XOR2_X1    g01042(.A1(\b[15] ), .A2(\b[16] ), .Z(new_n1299_));
  OAI21_X1   g01043(.A1(new_n1272_), .A2(\b[14] ), .B(\b[15] ), .ZN(new_n1300_));
  NAND2_X1   g01044(.A1(new_n1271_), .A2(\b[14] ), .ZN(new_n1301_));
  AOI21_X1   g01045(.A1(new_n1300_), .A2(new_n1301_), .B(new_n1299_), .ZN(new_n1302_));
  INV_X1     g01046(.I(new_n1299_), .ZN(new_n1303_));
  NAND2_X1   g01047(.A1(new_n1300_), .A2(new_n1301_), .ZN(new_n1304_));
  NOR2_X1    g01048(.A1(new_n1304_), .A2(new_n1303_), .ZN(new_n1305_));
  NOR2_X1    g01049(.A1(new_n1305_), .A2(new_n1302_), .ZN(new_n1306_));
  OAI21_X1   g01050(.A1(new_n1306_), .A2(new_n279_), .B(new_n1298_), .ZN(new_n1307_));
  XOR2_X1    g01051(.A1(new_n1307_), .A2(\a[2] ), .Z(new_n1308_));
  AOI22_X1   g01052(.A1(new_n1191_), .A2(new_n1192_), .B1(new_n1198_), .B2(new_n1262_), .ZN(new_n1309_));
  AOI22_X1   g01053(.A1(new_n800_), .A2(\b[12] ), .B1(\b[13] ), .B2(new_n333_), .ZN(new_n1310_));
  OAI21_X1   g01054(.A1(new_n852_), .A2(new_n392_), .B(new_n1310_), .ZN(new_n1311_));
  INV_X1     g01055(.I(new_n1311_), .ZN(new_n1312_));
  OAI21_X1   g01056(.A1(new_n1082_), .A2(new_n318_), .B(new_n1312_), .ZN(new_n1313_));
  XOR2_X1    g01057(.A1(new_n1313_), .A2(new_n312_), .Z(new_n1314_));
  OAI21_X1   g01058(.A1(new_n1257_), .A2(new_n1251_), .B(new_n1253_), .ZN(new_n1315_));
  OAI21_X1   g01059(.A1(new_n1228_), .A2(new_n1226_), .B(new_n1220_), .ZN(new_n1316_));
  NAND2_X1   g01060(.A1(new_n1316_), .A2(new_n1235_), .ZN(new_n1317_));
  NAND2_X1   g01061(.A1(new_n1005_), .A2(new_n990_), .ZN(new_n1318_));
  NAND3_X1   g01062(.A1(new_n1318_), .A2(new_n1140_), .A3(\b[4] ), .ZN(new_n1319_));
  NAND2_X1   g01063(.A1(new_n1009_), .A2(\b[3] ), .ZN(new_n1320_));
  NAND4_X1   g01064(.A1(new_n898_), .A2(new_n1155_), .A3(\b[2] ), .A4(new_n1142_), .ZN(new_n1321_));
  NAND3_X1   g01065(.A1(new_n1321_), .A2(new_n1319_), .A3(new_n1320_), .ZN(new_n1322_));
  INV_X1     g01066(.I(new_n1013_), .ZN(new_n1323_));
  NOR2_X1    g01067(.A1(new_n352_), .A2(new_n1323_), .ZN(new_n1324_));
  OAI21_X1   g01068(.A1(new_n1324_), .A2(new_n1322_), .B(\a[14] ), .ZN(new_n1325_));
  AOI22_X1   g01069(.A1(new_n1006_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n1009_), .ZN(new_n1326_));
  OAI21_X1   g01070(.A1(new_n346_), .A2(new_n351_), .B(new_n1013_), .ZN(new_n1327_));
  NAND4_X1   g01071(.A1(new_n1327_), .A2(new_n1326_), .A3(new_n1002_), .A4(new_n1321_), .ZN(new_n1328_));
  NAND2_X1   g01072(.A1(new_n1325_), .A2(new_n1328_), .ZN(new_n1329_));
  NAND2_X1   g01073(.A1(new_n1002_), .A2(\a[15] ), .ZN(new_n1330_));
  INV_X1     g01074(.I(\a[15] ), .ZN(new_n1331_));
  NAND2_X1   g01075(.A1(new_n1331_), .A2(\a[14] ), .ZN(new_n1332_));
  NAND2_X1   g01076(.A1(new_n1330_), .A2(new_n1332_), .ZN(new_n1333_));
  XNOR2_X1   g01077(.A1(\a[16] ), .A2(\a[17] ), .ZN(new_n1334_));
  NAND3_X1   g01078(.A1(new_n1333_), .A2(new_n1334_), .A3(\b[1] ), .ZN(new_n1335_));
  INV_X1     g01079(.I(\a[16] ), .ZN(new_n1336_));
  NOR3_X1    g01080(.A1(new_n1336_), .A2(\a[14] ), .A3(\a[15] ), .ZN(new_n1337_));
  NOR3_X1    g01081(.A1(new_n1002_), .A2(new_n1331_), .A3(\a[16] ), .ZN(new_n1338_));
  OAI21_X1   g01082(.A1(new_n1338_), .A2(new_n1337_), .B(\b[0] ), .ZN(new_n1339_));
  NAND2_X1   g01083(.A1(new_n1335_), .A2(new_n1339_), .ZN(new_n1340_));
  XNOR2_X1   g01084(.A1(\a[16] ), .A2(\a[17] ), .ZN(new_n1341_));
  NOR3_X1    g01085(.A1(new_n1206_), .A2(new_n1341_), .A3(new_n313_), .ZN(new_n1342_));
  OAI21_X1   g01086(.A1(new_n1340_), .A2(new_n1342_), .B(\a[17] ), .ZN(new_n1343_));
  INV_X1     g01087(.I(\a[17] ), .ZN(new_n1344_));
  XOR2_X1    g01088(.A1(\a[16] ), .A2(\a[17] ), .Z(new_n1345_));
  NOR3_X1    g01089(.A1(new_n1206_), .A2(new_n1345_), .A3(new_n275_), .ZN(new_n1346_));
  INV_X1     g01090(.I(new_n1339_), .ZN(new_n1347_));
  NOR3_X1    g01091(.A1(new_n1342_), .A2(new_n1347_), .A3(new_n1346_), .ZN(new_n1348_));
  NAND2_X1   g01092(.A1(new_n1348_), .A2(new_n1344_), .ZN(new_n1349_));
  NAND2_X1   g01093(.A1(new_n1214_), .A2(\a[17] ), .ZN(new_n1350_));
  NAND3_X1   g01094(.A1(new_n1349_), .A2(new_n1343_), .A3(new_n1350_), .ZN(new_n1351_));
  NAND2_X1   g01095(.A1(new_n1336_), .A2(\a[17] ), .ZN(new_n1352_));
  NAND2_X1   g01096(.A1(new_n1344_), .A2(\a[16] ), .ZN(new_n1353_));
  AOI22_X1   g01097(.A1(new_n1330_), .A2(new_n1332_), .B1(new_n1352_), .B2(new_n1353_), .ZN(new_n1354_));
  NAND2_X1   g01098(.A1(new_n1354_), .A2(new_n263_), .ZN(new_n1355_));
  NAND3_X1   g01099(.A1(new_n1355_), .A2(new_n1335_), .A3(new_n1339_), .ZN(new_n1356_));
  NAND3_X1   g01100(.A1(new_n1356_), .A2(\a[17] ), .A3(new_n1214_), .ZN(new_n1357_));
  AOI21_X1   g01101(.A1(new_n1351_), .A2(new_n1357_), .B(new_n1329_), .ZN(new_n1358_));
  AND3_X2    g01102(.A1(new_n1321_), .A2(new_n1319_), .A3(new_n1320_), .Z(new_n1359_));
  AOI21_X1   g01103(.A1(new_n1359_), .A2(new_n1327_), .B(new_n1002_), .ZN(new_n1360_));
  INV_X1     g01104(.I(new_n1328_), .ZN(new_n1361_));
  NOR2_X1    g01105(.A1(new_n1360_), .A2(new_n1361_), .ZN(new_n1362_));
  NAND2_X1   g01106(.A1(new_n1351_), .A2(new_n1357_), .ZN(new_n1363_));
  NOR2_X1    g01107(.A1(new_n1363_), .A2(new_n1362_), .ZN(new_n1364_));
  NOR2_X1    g01108(.A1(new_n1364_), .A2(new_n1358_), .ZN(new_n1365_));
  OAI21_X1   g01109(.A1(new_n1167_), .A2(new_n1215_), .B(new_n1217_), .ZN(new_n1366_));
  NOR2_X1    g01110(.A1(new_n1365_), .A2(new_n1366_), .ZN(new_n1367_));
  NAND2_X1   g01111(.A1(new_n1363_), .A2(new_n1362_), .ZN(new_n1368_));
  NAND3_X1   g01112(.A1(new_n1329_), .A2(new_n1351_), .A3(new_n1357_), .ZN(new_n1369_));
  NAND2_X1   g01113(.A1(new_n1368_), .A2(new_n1369_), .ZN(new_n1370_));
  AOI21_X1   g01114(.A1(new_n1159_), .A2(new_n1218_), .B(new_n1208_), .ZN(new_n1371_));
  NOR2_X1    g01115(.A1(new_n1370_), .A2(new_n1371_), .ZN(new_n1372_));
  OAI22_X1   g01116(.A1(new_n713_), .A2(new_n471_), .B1(new_n438_), .B2(new_n717_), .ZN(new_n1373_));
  NOR2_X1    g01117(.A1(new_n1127_), .A2(new_n377_), .ZN(new_n1374_));
  NOR2_X1    g01118(.A1(new_n1374_), .A2(new_n1373_), .ZN(new_n1375_));
  NAND3_X1   g01119(.A1(new_n484_), .A2(new_n477_), .A3(new_n724_), .ZN(new_n1376_));
  AOI21_X1   g01120(.A1(new_n1376_), .A2(new_n1375_), .B(new_n722_), .ZN(new_n1377_));
  INV_X1     g01121(.I(new_n1375_), .ZN(new_n1378_));
  NOR3_X1    g01122(.A1(new_n1037_), .A2(new_n1038_), .A3(new_n986_), .ZN(new_n1379_));
  NOR3_X1    g01123(.A1(new_n1379_), .A2(\a[11] ), .A3(new_n1378_), .ZN(new_n1380_));
  NOR2_X1    g01124(.A1(new_n1380_), .A2(new_n1377_), .ZN(new_n1381_));
  NOR3_X1    g01125(.A1(new_n1367_), .A2(new_n1372_), .A3(new_n1381_), .ZN(new_n1382_));
  NAND2_X1   g01126(.A1(new_n1370_), .A2(new_n1371_), .ZN(new_n1383_));
  NAND2_X1   g01127(.A1(new_n1365_), .A2(new_n1366_), .ZN(new_n1384_));
  OAI21_X1   g01128(.A1(new_n1379_), .A2(new_n1378_), .B(\a[11] ), .ZN(new_n1385_));
  NAND3_X1   g01129(.A1(new_n1376_), .A2(new_n722_), .A3(new_n1375_), .ZN(new_n1386_));
  NAND2_X1   g01130(.A1(new_n1385_), .A2(new_n1386_), .ZN(new_n1387_));
  AOI21_X1   g01131(.A1(new_n1384_), .A2(new_n1383_), .B(new_n1387_), .ZN(new_n1388_));
  NOR2_X1    g01132(.A1(new_n1388_), .A2(new_n1382_), .ZN(new_n1389_));
  NAND2_X1   g01133(.A1(new_n1317_), .A2(new_n1389_), .ZN(new_n1390_));
  AOI21_X1   g01134(.A1(new_n1231_), .A2(new_n1225_), .B(new_n1221_), .ZN(new_n1391_));
  NOR2_X1    g01135(.A1(new_n1391_), .A2(new_n1232_), .ZN(new_n1392_));
  NAND3_X1   g01136(.A1(new_n1384_), .A2(new_n1383_), .A3(new_n1387_), .ZN(new_n1393_));
  OAI21_X1   g01137(.A1(new_n1367_), .A2(new_n1372_), .B(new_n1381_), .ZN(new_n1394_));
  NAND2_X1   g01138(.A1(new_n1394_), .A2(new_n1393_), .ZN(new_n1395_));
  NAND2_X1   g01139(.A1(new_n1392_), .A2(new_n1395_), .ZN(new_n1396_));
  AOI22_X1   g01140(.A1(new_n518_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n636_), .ZN(new_n1397_));
  OAI21_X1   g01141(.A1(new_n577_), .A2(new_n917_), .B(new_n1397_), .ZN(new_n1398_));
  INV_X1     g01142(.I(new_n1398_), .ZN(new_n1399_));
  OAI21_X1   g01143(.A1(new_n786_), .A2(new_n624_), .B(new_n1399_), .ZN(new_n1400_));
  NAND2_X1   g01144(.A1(new_n1400_), .A2(\a[8] ), .ZN(new_n1401_));
  AOI21_X1   g01145(.A1(new_n1059_), .A2(new_n618_), .B(new_n1398_), .ZN(new_n1402_));
  NAND2_X1   g01146(.A1(new_n1402_), .A2(new_n488_), .ZN(new_n1403_));
  NAND2_X1   g01147(.A1(new_n1401_), .A2(new_n1403_), .ZN(new_n1404_));
  AOI21_X1   g01148(.A1(new_n1390_), .A2(new_n1396_), .B(new_n1404_), .ZN(new_n1405_));
  NOR2_X1    g01149(.A1(new_n1392_), .A2(new_n1395_), .ZN(new_n1406_));
  NOR2_X1    g01150(.A1(new_n1317_), .A2(new_n1389_), .ZN(new_n1407_));
  NOR2_X1    g01151(.A1(new_n1402_), .A2(new_n488_), .ZN(new_n1408_));
  NOR2_X1    g01152(.A1(new_n1400_), .A2(\a[8] ), .ZN(new_n1409_));
  NOR2_X1    g01153(.A1(new_n1409_), .A2(new_n1408_), .ZN(new_n1410_));
  NOR3_X1    g01154(.A1(new_n1410_), .A2(new_n1407_), .A3(new_n1406_), .ZN(new_n1411_));
  NOR2_X1    g01155(.A1(new_n1405_), .A2(new_n1411_), .ZN(new_n1412_));
  XOR2_X1    g01156(.A1(new_n1315_), .A2(new_n1412_), .Z(new_n1413_));
  NOR2_X1    g01157(.A1(new_n1413_), .A2(new_n1314_), .ZN(new_n1414_));
  XOR2_X1    g01158(.A1(new_n1313_), .A2(\a[5] ), .Z(new_n1415_));
  NAND2_X1   g01159(.A1(new_n1315_), .A2(new_n1412_), .ZN(new_n1416_));
  INV_X1     g01160(.I(new_n1416_), .ZN(new_n1417_));
  NOR2_X1    g01161(.A1(new_n1315_), .A2(new_n1412_), .ZN(new_n1418_));
  NOR3_X1    g01162(.A1(new_n1415_), .A2(new_n1417_), .A3(new_n1418_), .ZN(new_n1419_));
  NOR4_X1    g01163(.A1(new_n1309_), .A2(new_n1263_), .A3(new_n1414_), .A4(new_n1419_), .ZN(new_n1420_));
  INV_X1     g01164(.I(new_n1420_), .ZN(new_n1421_));
  OAI22_X1   g01165(.A1(new_n1309_), .A2(new_n1263_), .B1(new_n1414_), .B2(new_n1419_), .ZN(new_n1422_));
  NAND2_X1   g01166(.A1(new_n1421_), .A2(new_n1422_), .ZN(new_n1423_));
  INV_X1     g01167(.I(new_n1423_), .ZN(new_n1424_));
  NOR2_X1    g01168(.A1(new_n1424_), .A2(new_n1308_), .ZN(new_n1425_));
  NAND2_X1   g01169(.A1(new_n1424_), .A2(new_n1308_), .ZN(new_n1426_));
  INV_X1     g01170(.I(new_n1426_), .ZN(new_n1427_));
  NOR2_X1    g01171(.A1(new_n1427_), .A2(new_n1425_), .ZN(new_n1428_));
  XOR2_X1    g01172(.A1(new_n1295_), .A2(new_n1428_), .Z(\f[16] ));
  INV_X1     g01173(.I(new_n1425_), .ZN(new_n1430_));
  AOI21_X1   g01174(.A1(new_n1295_), .A2(new_n1430_), .B(new_n1427_), .ZN(new_n1431_));
  INV_X1     g01175(.I(\b[17] ), .ZN(new_n1432_));
  OAI22_X1   g01176(.A1(new_n277_), .A2(new_n1432_), .B1(new_n1296_), .B2(new_n262_), .ZN(new_n1433_));
  AOI21_X1   g01177(.A1(\b[15] ), .A2(new_n283_), .B(new_n1433_), .ZN(new_n1434_));
  AOI21_X1   g01178(.A1(new_n1304_), .A2(\b[16] ), .B(new_n1268_), .ZN(new_n1435_));
  NOR2_X1    g01179(.A1(new_n1304_), .A2(\b[16] ), .ZN(new_n1436_));
  NAND3_X1   g01180(.A1(new_n1300_), .A2(new_n1301_), .A3(new_n1432_), .ZN(new_n1437_));
  INV_X1     g01181(.I(new_n1437_), .ZN(new_n1438_));
  AOI21_X1   g01182(.A1(new_n1300_), .A2(new_n1301_), .B(new_n1432_), .ZN(new_n1439_));
  OAI22_X1   g01183(.A1(new_n1435_), .A2(new_n1436_), .B1(new_n1438_), .B2(new_n1439_), .ZN(new_n1440_));
  NOR2_X1    g01184(.A1(new_n1435_), .A2(new_n1436_), .ZN(new_n1441_));
  NOR2_X1    g01185(.A1(new_n1438_), .A2(new_n1439_), .ZN(new_n1442_));
  NAND2_X1   g01186(.A1(new_n1441_), .A2(new_n1442_), .ZN(new_n1443_));
  NAND2_X1   g01187(.A1(new_n1443_), .A2(new_n1440_), .ZN(new_n1444_));
  OAI21_X1   g01188(.A1(new_n1444_), .A2(new_n279_), .B(new_n1434_), .ZN(new_n1445_));
  XOR2_X1    g01189(.A1(new_n1445_), .A2(\a[2] ), .Z(new_n1446_));
  OR2_X2     g01190(.A1(new_n1098_), .A2(new_n1099_), .Z(new_n1447_));
  INV_X1     g01191(.I(new_n1102_), .ZN(new_n1448_));
  NAND2_X1   g01192(.A1(new_n1447_), .A2(new_n1448_), .ZN(new_n1449_));
  AOI22_X1   g01193(.A1(new_n800_), .A2(\b[13] ), .B1(\b[14] ), .B2(new_n333_), .ZN(new_n1450_));
  OAI21_X1   g01194(.A1(new_n941_), .A2(new_n392_), .B(new_n1450_), .ZN(new_n1451_));
  AOI21_X1   g01195(.A1(new_n1449_), .A2(new_n330_), .B(new_n1451_), .ZN(new_n1452_));
  XOR2_X1    g01196(.A1(new_n1452_), .A2(new_n312_), .Z(new_n1453_));
  INV_X1     g01197(.I(new_n1453_), .ZN(new_n1454_));
  OAI21_X1   g01198(.A1(new_n1406_), .A2(new_n1407_), .B(new_n1410_), .ZN(new_n1455_));
  AOI21_X1   g01199(.A1(new_n1315_), .A2(new_n1455_), .B(new_n1411_), .ZN(new_n1456_));
  AOI22_X1   g01200(.A1(new_n518_), .A2(\b[11] ), .B1(\b[10] ), .B2(new_n636_), .ZN(new_n1457_));
  OAI21_X1   g01201(.A1(new_n667_), .A2(new_n917_), .B(new_n1457_), .ZN(new_n1458_));
  AOI21_X1   g01202(.A1(new_n856_), .A2(new_n857_), .B(new_n852_), .ZN(new_n1459_));
  NOR3_X1    g01203(.A1(new_n849_), .A2(\b[11] ), .A3(new_n850_), .ZN(new_n1460_));
  NOR3_X1    g01204(.A1(new_n1459_), .A2(new_n624_), .A3(new_n1460_), .ZN(new_n1461_));
  OAI21_X1   g01205(.A1(new_n1461_), .A2(new_n1458_), .B(\a[8] ), .ZN(new_n1462_));
  INV_X1     g01206(.I(new_n1458_), .ZN(new_n1463_));
  NAND3_X1   g01207(.A1(new_n858_), .A2(new_n618_), .A3(new_n851_), .ZN(new_n1464_));
  NAND3_X1   g01208(.A1(new_n1464_), .A2(new_n488_), .A3(new_n1463_), .ZN(new_n1465_));
  OAI21_X1   g01209(.A1(new_n1391_), .A2(new_n1232_), .B(new_n1394_), .ZN(new_n1466_));
  OAI22_X1   g01210(.A1(new_n713_), .A2(new_n577_), .B1(new_n471_), .B2(new_n717_), .ZN(new_n1467_));
  NOR2_X1    g01211(.A1(new_n1127_), .A2(new_n438_), .ZN(new_n1468_));
  NOR2_X1    g01212(.A1(new_n1468_), .A2(new_n1467_), .ZN(new_n1469_));
  INV_X1     g01213(.I(new_n1469_), .ZN(new_n1470_));
  AOI21_X1   g01214(.A1(new_n798_), .A2(new_n585_), .B(new_n986_), .ZN(new_n1471_));
  OAI21_X1   g01215(.A1(new_n1471_), .A2(new_n1470_), .B(\a[11] ), .ZN(new_n1472_));
  OAI21_X1   g01216(.A1(new_n586_), .A2(new_n584_), .B(new_n724_), .ZN(new_n1473_));
  NAND3_X1   g01217(.A1(new_n1473_), .A2(new_n722_), .A3(new_n1469_), .ZN(new_n1474_));
  OAI21_X1   g01218(.A1(new_n1366_), .A2(new_n1364_), .B(new_n1368_), .ZN(new_n1475_));
  NAND3_X1   g01219(.A1(new_n1475_), .A2(new_n1472_), .A3(new_n1474_), .ZN(new_n1476_));
  AOI21_X1   g01220(.A1(new_n1473_), .A2(new_n1469_), .B(new_n722_), .ZN(new_n1477_));
  NOR3_X1    g01221(.A1(new_n1471_), .A2(\a[11] ), .A3(new_n1470_), .ZN(new_n1478_));
  AOI21_X1   g01222(.A1(new_n1371_), .A2(new_n1369_), .B(new_n1358_), .ZN(new_n1479_));
  OAI21_X1   g01223(.A1(new_n1477_), .A2(new_n1478_), .B(new_n1479_), .ZN(new_n1480_));
  NAND3_X1   g01224(.A1(new_n898_), .A2(new_n1155_), .A3(new_n1142_), .ZN(new_n1481_));
  AOI22_X1   g01225(.A1(new_n1006_), .A2(\b[5] ), .B1(\b[4] ), .B2(new_n1009_), .ZN(new_n1482_));
  OAI21_X1   g01226(.A1(new_n290_), .A2(new_n1481_), .B(new_n1482_), .ZN(new_n1483_));
  AOI21_X1   g01227(.A1(new_n382_), .A2(new_n1013_), .B(new_n1483_), .ZN(new_n1484_));
  NOR2_X1    g01228(.A1(new_n1484_), .A2(new_n1002_), .ZN(new_n1485_));
  INV_X1     g01229(.I(new_n1481_), .ZN(new_n1486_));
  OAI22_X1   g01230(.A1(new_n993_), .A2(new_n377_), .B1(new_n339_), .B2(new_n997_), .ZN(new_n1487_));
  AOI21_X1   g01231(.A1(\b[3] ), .A2(new_n1486_), .B(new_n1487_), .ZN(new_n1488_));
  OAI21_X1   g01232(.A1(new_n566_), .A2(new_n1323_), .B(new_n1488_), .ZN(new_n1489_));
  NOR2_X1    g01233(.A1(new_n1489_), .A2(\a[14] ), .ZN(new_n1490_));
  NAND2_X1   g01234(.A1(new_n1354_), .A2(new_n554_), .ZN(new_n1491_));
  NAND3_X1   g01235(.A1(new_n1333_), .A2(new_n1334_), .A3(\b[2] ), .ZN(new_n1492_));
  NAND3_X1   g01236(.A1(new_n1002_), .A2(new_n1331_), .A3(\a[16] ), .ZN(new_n1493_));
  NAND3_X1   g01237(.A1(new_n1336_), .A2(\a[14] ), .A3(\a[15] ), .ZN(new_n1494_));
  NAND2_X1   g01238(.A1(new_n1493_), .A2(new_n1494_), .ZN(new_n1495_));
  NAND2_X1   g01239(.A1(new_n1495_), .A2(\b[1] ), .ZN(new_n1496_));
  AOI21_X1   g01240(.A1(new_n1336_), .A2(\a[17] ), .B(\a[14] ), .ZN(new_n1497_));
  INV_X1     g01241(.I(new_n1497_), .ZN(new_n1498_));
  NAND2_X1   g01242(.A1(new_n1353_), .A2(\a[14] ), .ZN(new_n1499_));
  NAND4_X1   g01243(.A1(new_n1206_), .A2(new_n1498_), .A3(new_n1499_), .A4(\b[0] ), .ZN(new_n1500_));
  NAND4_X1   g01244(.A1(new_n1491_), .A2(new_n1500_), .A3(new_n1492_), .A4(new_n1496_), .ZN(new_n1501_));
  NAND2_X1   g01245(.A1(new_n1501_), .A2(\a[17] ), .ZN(new_n1502_));
  NOR3_X1    g01246(.A1(new_n282_), .A2(new_n1206_), .A3(new_n1341_), .ZN(new_n1503_));
  NOR3_X1    g01247(.A1(new_n1206_), .A2(new_n1345_), .A3(new_n276_), .ZN(new_n1504_));
  NOR2_X1    g01248(.A1(new_n1338_), .A2(new_n1337_), .ZN(new_n1505_));
  NOR2_X1    g01249(.A1(new_n1505_), .A2(new_n275_), .ZN(new_n1506_));
  AOI21_X1   g01250(.A1(\a[16] ), .A2(new_n1344_), .B(new_n1002_), .ZN(new_n1507_));
  NOR4_X1    g01251(.A1(new_n1333_), .A2(new_n258_), .A3(new_n1497_), .A4(new_n1507_), .ZN(new_n1508_));
  NOR4_X1    g01252(.A1(new_n1503_), .A2(new_n1508_), .A3(new_n1506_), .A4(new_n1504_), .ZN(new_n1509_));
  NAND2_X1   g01253(.A1(new_n1509_), .A2(new_n1344_), .ZN(new_n1510_));
  NOR3_X1    g01254(.A1(new_n1356_), .A2(new_n1344_), .A3(new_n1207_), .ZN(new_n1511_));
  AOI21_X1   g01255(.A1(new_n1502_), .A2(new_n1510_), .B(new_n1511_), .ZN(new_n1512_));
  NOR4_X1    g01256(.A1(new_n1501_), .A2(new_n1356_), .A3(new_n1344_), .A4(new_n1207_), .ZN(new_n1513_));
  NOR4_X1    g01257(.A1(new_n1485_), .A2(new_n1490_), .A3(new_n1512_), .A4(new_n1513_), .ZN(new_n1514_));
  NAND2_X1   g01258(.A1(new_n1489_), .A2(\a[14] ), .ZN(new_n1515_));
  NAND2_X1   g01259(.A1(new_n1484_), .A2(new_n1002_), .ZN(new_n1516_));
  NAND2_X1   g01260(.A1(new_n1502_), .A2(new_n1510_), .ZN(new_n1517_));
  INV_X1     g01261(.I(new_n1511_), .ZN(new_n1518_));
  NAND2_X1   g01262(.A1(new_n1517_), .A2(new_n1518_), .ZN(new_n1519_));
  NAND4_X1   g01263(.A1(new_n1509_), .A2(\a[17] ), .A3(new_n1348_), .A4(new_n1214_), .ZN(new_n1520_));
  AOI22_X1   g01264(.A1(new_n1516_), .A2(new_n1515_), .B1(new_n1519_), .B2(new_n1520_), .ZN(new_n1521_));
  NOR2_X1    g01265(.A1(new_n1521_), .A2(new_n1514_), .ZN(new_n1522_));
  NAND3_X1   g01266(.A1(new_n1480_), .A2(new_n1476_), .A3(new_n1522_), .ZN(new_n1523_));
  NOR3_X1    g01267(.A1(new_n1479_), .A2(new_n1478_), .A3(new_n1477_), .ZN(new_n1524_));
  AOI21_X1   g01268(.A1(new_n1472_), .A2(new_n1474_), .B(new_n1475_), .ZN(new_n1525_));
  NAND4_X1   g01269(.A1(new_n1516_), .A2(new_n1519_), .A3(new_n1515_), .A4(new_n1520_), .ZN(new_n1526_));
  OAI22_X1   g01270(.A1(new_n1485_), .A2(new_n1490_), .B1(new_n1512_), .B2(new_n1513_), .ZN(new_n1527_));
  NAND2_X1   g01271(.A1(new_n1527_), .A2(new_n1526_), .ZN(new_n1528_));
  OAI21_X1   g01272(.A1(new_n1525_), .A2(new_n1524_), .B(new_n1528_), .ZN(new_n1529_));
  NAND4_X1   g01273(.A1(new_n1466_), .A2(new_n1393_), .A3(new_n1523_), .A4(new_n1529_), .ZN(new_n1530_));
  AOI21_X1   g01274(.A1(new_n1316_), .A2(new_n1235_), .B(new_n1388_), .ZN(new_n1531_));
  NOR3_X1    g01275(.A1(new_n1525_), .A2(new_n1524_), .A3(new_n1528_), .ZN(new_n1532_));
  AOI21_X1   g01276(.A1(new_n1480_), .A2(new_n1476_), .B(new_n1522_), .ZN(new_n1533_));
  OAI22_X1   g01277(.A1(new_n1531_), .A2(new_n1382_), .B1(new_n1532_), .B2(new_n1533_), .ZN(new_n1534_));
  NAND4_X1   g01278(.A1(new_n1534_), .A2(new_n1530_), .A3(new_n1462_), .A4(new_n1465_), .ZN(new_n1535_));
  AOI21_X1   g01279(.A1(new_n1464_), .A2(new_n1463_), .B(new_n488_), .ZN(new_n1536_));
  NOR3_X1    g01280(.A1(new_n1461_), .A2(\a[8] ), .A3(new_n1458_), .ZN(new_n1537_));
  NAND2_X1   g01281(.A1(new_n1529_), .A2(new_n1523_), .ZN(new_n1538_));
  NOR3_X1    g01282(.A1(new_n1538_), .A2(new_n1531_), .A3(new_n1382_), .ZN(new_n1539_));
  AOI22_X1   g01283(.A1(new_n1466_), .A2(new_n1393_), .B1(new_n1523_), .B2(new_n1529_), .ZN(new_n1540_));
  OAI22_X1   g01284(.A1(new_n1539_), .A2(new_n1540_), .B1(new_n1536_), .B2(new_n1537_), .ZN(new_n1541_));
  NAND2_X1   g01285(.A1(new_n1541_), .A2(new_n1535_), .ZN(new_n1542_));
  XOR2_X1    g01286(.A1(new_n1456_), .A2(new_n1542_), .Z(new_n1543_));
  XOR2_X1    g01287(.A1(new_n1543_), .A2(new_n1454_), .Z(new_n1544_));
  NOR2_X1    g01288(.A1(new_n1420_), .A2(new_n1414_), .ZN(new_n1545_));
  XOR2_X1    g01289(.A1(new_n1545_), .A2(new_n1544_), .Z(new_n1546_));
  XOR2_X1    g01290(.A1(new_n1546_), .A2(new_n1446_), .Z(new_n1547_));
  XOR2_X1    g01291(.A1(new_n1431_), .A2(new_n1547_), .Z(\f[17] ));
  INV_X1     g01292(.I(new_n1446_), .ZN(new_n1549_));
  NOR2_X1    g01293(.A1(new_n1546_), .A2(new_n1549_), .ZN(new_n1550_));
  INV_X1     g01294(.I(new_n1550_), .ZN(new_n1551_));
  OAI21_X1   g01295(.A1(new_n1431_), .A2(new_n1547_), .B(new_n1551_), .ZN(new_n1552_));
  INV_X1     g01296(.I(\b[18] ), .ZN(new_n1553_));
  OAI22_X1   g01297(.A1(new_n277_), .A2(new_n1553_), .B1(new_n1432_), .B2(new_n262_), .ZN(new_n1554_));
  AOI21_X1   g01298(.A1(\b[16] ), .A2(new_n283_), .B(new_n1554_), .ZN(new_n1555_));
  AOI21_X1   g01299(.A1(new_n1437_), .A2(\b[16] ), .B(\b[15] ), .ZN(new_n1556_));
  NOR2_X1    g01300(.A1(new_n1439_), .A2(\b[16] ), .ZN(new_n1557_));
  NOR2_X1    g01301(.A1(new_n1556_), .A2(new_n1557_), .ZN(new_n1558_));
  XNOR2_X1   g01302(.A1(\b[17] ), .A2(\b[18] ), .ZN(new_n1559_));
  NOR2_X1    g01303(.A1(new_n1558_), .A2(new_n1559_), .ZN(new_n1560_));
  XOR2_X1    g01304(.A1(\b[17] ), .A2(\b[18] ), .Z(new_n1561_));
  INV_X1     g01305(.I(new_n1561_), .ZN(new_n1562_));
  AOI21_X1   g01306(.A1(new_n1558_), .A2(new_n1562_), .B(new_n1560_), .ZN(new_n1563_));
  OAI21_X1   g01307(.A1(new_n1563_), .A2(new_n279_), .B(new_n1555_), .ZN(new_n1564_));
  XOR2_X1    g01308(.A1(new_n1564_), .A2(\a[2] ), .Z(new_n1565_));
  INV_X1     g01309(.I(new_n1565_), .ZN(new_n1566_));
  OAI21_X1   g01310(.A1(new_n1420_), .A2(new_n1414_), .B(new_n1453_), .ZN(new_n1567_));
  NOR3_X1    g01311(.A1(new_n1420_), .A2(new_n1414_), .A3(new_n1453_), .ZN(new_n1568_));
  AOI21_X1   g01312(.A1(new_n1543_), .A2(new_n1567_), .B(new_n1568_), .ZN(new_n1569_));
  OAI22_X1   g01313(.A1(new_n321_), .A2(new_n1268_), .B1(new_n325_), .B2(new_n1093_), .ZN(new_n1570_));
  AOI21_X1   g01314(.A1(\b[13] ), .A2(new_n602_), .B(new_n1570_), .ZN(new_n1571_));
  OAI21_X1   g01315(.A1(new_n1275_), .A2(new_n318_), .B(new_n1571_), .ZN(new_n1572_));
  XOR2_X1    g01316(.A1(new_n1572_), .A2(\a[5] ), .Z(new_n1573_));
  OAI21_X1   g01317(.A1(new_n1479_), .A2(new_n1521_), .B(new_n1526_), .ZN(new_n1574_));
  OAI22_X1   g01318(.A1(new_n993_), .A2(new_n438_), .B1(new_n377_), .B2(new_n997_), .ZN(new_n1575_));
  NOR2_X1    g01319(.A1(new_n1481_), .A2(new_n339_), .ZN(new_n1576_));
  NOR2_X1    g01320(.A1(new_n1576_), .A2(new_n1575_), .ZN(new_n1577_));
  OAI21_X1   g01321(.A1(new_n447_), .A2(new_n449_), .B(new_n1013_), .ZN(new_n1578_));
  AOI21_X1   g01322(.A1(new_n1578_), .A2(new_n1577_), .B(new_n1002_), .ZN(new_n1579_));
  INV_X1     g01323(.I(new_n1577_), .ZN(new_n1580_));
  AOI21_X1   g01324(.A1(new_n915_), .A2(new_n446_), .B(new_n1323_), .ZN(new_n1581_));
  NOR3_X1    g01325(.A1(new_n1581_), .A2(new_n1580_), .A3(\a[14] ), .ZN(new_n1582_));
  NOR2_X1    g01326(.A1(new_n1579_), .A2(new_n1582_), .ZN(new_n1583_));
  NOR3_X1    g01327(.A1(new_n1333_), .A2(new_n1497_), .A3(new_n1507_), .ZN(new_n1584_));
  NAND2_X1   g01328(.A1(new_n1584_), .A2(\b[1] ), .ZN(new_n1585_));
  NOR2_X1    g01329(.A1(new_n1206_), .A2(new_n1345_), .ZN(new_n1586_));
  AOI21_X1   g01330(.A1(new_n1493_), .A2(new_n1494_), .B(new_n276_), .ZN(new_n1587_));
  AOI21_X1   g01331(.A1(new_n1586_), .A2(\b[3] ), .B(new_n1587_), .ZN(new_n1588_));
  NAND3_X1   g01332(.A1(new_n1354_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n1589_));
  NAND3_X1   g01333(.A1(new_n1585_), .A2(new_n1588_), .A3(new_n1589_), .ZN(new_n1590_));
  NAND2_X1   g01334(.A1(new_n1590_), .A2(\a[17] ), .ZN(new_n1591_));
  NAND2_X1   g01335(.A1(new_n1333_), .A2(new_n1334_), .ZN(new_n1592_));
  NOR2_X1    g01336(.A1(new_n1592_), .A2(new_n290_), .ZN(new_n1593_));
  NOR4_X1    g01337(.A1(new_n298_), .A2(new_n295_), .A3(new_n1206_), .A4(new_n1341_), .ZN(new_n1594_));
  NOR3_X1    g01338(.A1(new_n1593_), .A2(new_n1594_), .A3(new_n1587_), .ZN(new_n1595_));
  NAND3_X1   g01339(.A1(new_n1595_), .A2(new_n1344_), .A3(new_n1585_), .ZN(new_n1596_));
  XNOR2_X1   g01340(.A1(\a[17] ), .A2(\a[18] ), .ZN(new_n1597_));
  NOR2_X1    g01341(.A1(new_n1597_), .A2(new_n258_), .ZN(new_n1598_));
  INV_X1     g01342(.I(new_n1598_), .ZN(new_n1599_));
  AOI21_X1   g01343(.A1(new_n1591_), .A2(new_n1596_), .B(new_n1599_), .ZN(new_n1600_));
  AOI21_X1   g01344(.A1(new_n1595_), .A2(new_n1585_), .B(new_n1344_), .ZN(new_n1601_));
  NOR2_X1    g01345(.A1(new_n1590_), .A2(\a[17] ), .ZN(new_n1602_));
  NOR3_X1    g01346(.A1(new_n1602_), .A2(new_n1601_), .A3(new_n1598_), .ZN(new_n1603_));
  OAI21_X1   g01347(.A1(new_n1603_), .A2(new_n1600_), .B(new_n1520_), .ZN(new_n1604_));
  OAI21_X1   g01348(.A1(new_n1602_), .A2(new_n1601_), .B(new_n1598_), .ZN(new_n1605_));
  NAND3_X1   g01349(.A1(new_n1591_), .A2(new_n1596_), .A3(new_n1599_), .ZN(new_n1606_));
  NAND3_X1   g01350(.A1(new_n1605_), .A2(new_n1606_), .A3(new_n1513_), .ZN(new_n1607_));
  NAND3_X1   g01351(.A1(new_n1604_), .A2(new_n1607_), .A3(new_n1583_), .ZN(new_n1608_));
  OAI21_X1   g01352(.A1(new_n1581_), .A2(new_n1580_), .B(\a[14] ), .ZN(new_n1609_));
  NAND3_X1   g01353(.A1(new_n1578_), .A2(new_n1002_), .A3(new_n1577_), .ZN(new_n1610_));
  NAND2_X1   g01354(.A1(new_n1609_), .A2(new_n1610_), .ZN(new_n1611_));
  AOI21_X1   g01355(.A1(new_n1605_), .A2(new_n1606_), .B(new_n1513_), .ZN(new_n1612_));
  NOR3_X1    g01356(.A1(new_n1603_), .A2(new_n1600_), .A3(new_n1520_), .ZN(new_n1613_));
  OAI21_X1   g01357(.A1(new_n1613_), .A2(new_n1612_), .B(new_n1611_), .ZN(new_n1614_));
  NAND2_X1   g01358(.A1(new_n1614_), .A2(new_n1608_), .ZN(new_n1615_));
  XOR2_X1    g01359(.A1(new_n1615_), .A2(new_n1574_), .Z(new_n1616_));
  INV_X1     g01360(.I(new_n1616_), .ZN(new_n1617_));
  AOI22_X1   g01361(.A1(new_n729_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n732_), .ZN(new_n1618_));
  OAI21_X1   g01362(.A1(new_n471_), .A2(new_n1127_), .B(new_n1618_), .ZN(new_n1619_));
  INV_X1     g01363(.I(new_n1619_), .ZN(new_n1620_));
  OAI21_X1   g01364(.A1(new_n1240_), .A2(new_n986_), .B(new_n1620_), .ZN(new_n1621_));
  XOR2_X1    g01365(.A1(new_n1621_), .A2(new_n722_), .Z(new_n1622_));
  NAND2_X1   g01366(.A1(new_n1472_), .A2(new_n1474_), .ZN(new_n1623_));
  NOR2_X1    g01367(.A1(new_n1528_), .A2(new_n1479_), .ZN(new_n1624_));
  NOR2_X1    g01368(.A1(new_n1522_), .A2(new_n1475_), .ZN(new_n1625_));
  NOR3_X1    g01369(.A1(new_n1625_), .A2(new_n1624_), .A3(new_n1623_), .ZN(new_n1626_));
  INV_X1     g01370(.I(new_n1626_), .ZN(new_n1627_));
  AOI21_X1   g01371(.A1(new_n1530_), .A2(new_n1627_), .B(new_n1622_), .ZN(new_n1628_));
  XOR2_X1    g01372(.A1(new_n1621_), .A2(\a[11] ), .Z(new_n1629_));
  NOR3_X1    g01373(.A1(new_n1539_), .A2(new_n1629_), .A3(new_n1626_), .ZN(new_n1630_));
  NOR3_X1    g01374(.A1(new_n1630_), .A2(new_n1628_), .A3(new_n1617_), .ZN(new_n1631_));
  OAI21_X1   g01375(.A1(new_n1539_), .A2(new_n1626_), .B(new_n1629_), .ZN(new_n1632_));
  NAND3_X1   g01376(.A1(new_n1530_), .A2(new_n1622_), .A3(new_n1627_), .ZN(new_n1633_));
  AOI21_X1   g01377(.A1(new_n1632_), .A2(new_n1633_), .B(new_n1616_), .ZN(new_n1634_));
  NOR2_X1    g01378(.A1(new_n1631_), .A2(new_n1634_), .ZN(new_n1635_));
  INV_X1     g01379(.I(new_n1411_), .ZN(new_n1636_));
  AOI21_X1   g01380(.A1(new_n1259_), .A2(new_n1258_), .B(new_n1257_), .ZN(new_n1637_));
  OAI21_X1   g01381(.A1(new_n1637_), .A2(new_n1260_), .B(new_n1455_), .ZN(new_n1638_));
  NAND2_X1   g01382(.A1(new_n1462_), .A2(new_n1465_), .ZN(new_n1639_));
  NOR3_X1    g01383(.A1(new_n1639_), .A2(new_n1539_), .A3(new_n1540_), .ZN(new_n1640_));
  AOI22_X1   g01384(.A1(new_n1534_), .A2(new_n1530_), .B1(new_n1462_), .B2(new_n1465_), .ZN(new_n1641_));
  NOR2_X1    g01385(.A1(new_n1641_), .A2(new_n1640_), .ZN(new_n1642_));
  NAND3_X1   g01386(.A1(new_n1638_), .A2(new_n1642_), .A3(new_n1636_), .ZN(new_n1643_));
  AOI22_X1   g01387(.A1(new_n518_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n636_), .ZN(new_n1644_));
  OAI21_X1   g01388(.A1(new_n776_), .A2(new_n917_), .B(new_n1644_), .ZN(new_n1645_));
  AOI21_X1   g01389(.A1(new_n1194_), .A2(new_n618_), .B(new_n1645_), .ZN(new_n1646_));
  XOR2_X1    g01390(.A1(new_n1646_), .A2(\a[8] ), .Z(new_n1647_));
  AOI21_X1   g01391(.A1(new_n1643_), .A2(new_n1535_), .B(new_n1647_), .ZN(new_n1648_));
  OAI21_X1   g01392(.A1(new_n1028_), .A2(new_n1032_), .B(new_n1044_), .ZN(new_n1649_));
  AOI21_X1   g01393(.A1(new_n1050_), .A2(new_n1649_), .B(new_n1045_), .ZN(new_n1650_));
  NOR3_X1    g01394(.A1(new_n1173_), .A2(new_n1172_), .A3(new_n1169_), .ZN(new_n1651_));
  AOI21_X1   g01395(.A1(new_n1125_), .A2(new_n1121_), .B(new_n1170_), .ZN(new_n1652_));
  NOR2_X1    g01396(.A1(new_n1651_), .A2(new_n1652_), .ZN(new_n1653_));
  XOR2_X1    g01397(.A1(new_n1169_), .A2(new_n1120_), .Z(new_n1654_));
  NOR3_X1    g01398(.A1(new_n1654_), .A2(new_n1122_), .A3(new_n1123_), .ZN(new_n1655_));
  AOI21_X1   g01399(.A1(new_n1650_), .A2(new_n1653_), .B(new_n1655_), .ZN(new_n1656_));
  OAI21_X1   g01400(.A1(new_n1656_), .A2(new_n1248_), .B(new_n1237_), .ZN(new_n1657_));
  AOI21_X1   g01401(.A1(new_n1657_), .A2(new_n1253_), .B(new_n1405_), .ZN(new_n1658_));
  NOR3_X1    g01402(.A1(new_n1658_), .A2(new_n1411_), .A3(new_n1542_), .ZN(new_n1659_));
  XOR2_X1    g01403(.A1(new_n1646_), .A2(new_n488_), .Z(new_n1660_));
  NOR3_X1    g01404(.A1(new_n1659_), .A2(new_n1640_), .A3(new_n1660_), .ZN(new_n1661_));
  NOR2_X1    g01405(.A1(new_n1661_), .A2(new_n1648_), .ZN(new_n1662_));
  NAND2_X1   g01406(.A1(new_n1662_), .A2(new_n1635_), .ZN(new_n1663_));
  NOR2_X1    g01407(.A1(new_n1662_), .A2(new_n1635_), .ZN(new_n1664_));
  INV_X1     g01408(.I(new_n1664_), .ZN(new_n1665_));
  AOI21_X1   g01409(.A1(new_n1665_), .A2(new_n1663_), .B(new_n1573_), .ZN(new_n1666_));
  INV_X1     g01410(.I(new_n1573_), .ZN(new_n1667_));
  INV_X1     g01411(.I(new_n1663_), .ZN(new_n1668_));
  NOR3_X1    g01412(.A1(new_n1667_), .A2(new_n1668_), .A3(new_n1664_), .ZN(new_n1669_));
  NOR2_X1    g01413(.A1(new_n1669_), .A2(new_n1666_), .ZN(new_n1670_));
  XOR2_X1    g01414(.A1(new_n1569_), .A2(new_n1670_), .Z(new_n1671_));
  NOR2_X1    g01415(.A1(new_n1671_), .A2(new_n1566_), .ZN(new_n1672_));
  OAI21_X1   g01416(.A1(new_n1668_), .A2(new_n1664_), .B(new_n1667_), .ZN(new_n1673_));
  NAND3_X1   g01417(.A1(new_n1665_), .A2(new_n1573_), .A3(new_n1663_), .ZN(new_n1674_));
  NAND2_X1   g01418(.A1(new_n1673_), .A2(new_n1674_), .ZN(new_n1675_));
  NOR2_X1    g01419(.A1(new_n1569_), .A2(new_n1675_), .ZN(new_n1676_));
  NAND2_X1   g01420(.A1(new_n1567_), .A2(new_n1543_), .ZN(new_n1677_));
  INV_X1     g01421(.I(new_n1568_), .ZN(new_n1678_));
  NAND2_X1   g01422(.A1(new_n1677_), .A2(new_n1678_), .ZN(new_n1679_));
  NOR2_X1    g01423(.A1(new_n1679_), .A2(new_n1670_), .ZN(new_n1680_));
  NOR2_X1    g01424(.A1(new_n1680_), .A2(new_n1676_), .ZN(new_n1681_));
  NOR2_X1    g01425(.A1(new_n1681_), .A2(new_n1565_), .ZN(new_n1682_));
  OR2_X2     g01426(.A1(new_n1672_), .A2(new_n1682_), .Z(new_n1683_));
  XOR2_X1    g01427(.A1(new_n1552_), .A2(new_n1683_), .Z(\f[18] ));
  NOR2_X1    g01428(.A1(new_n284_), .A2(new_n1432_), .ZN(new_n1685_));
  INV_X1     g01429(.I(new_n1685_), .ZN(new_n1686_));
  AOI22_X1   g01430(.A1(new_n267_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n261_), .ZN(new_n1687_));
  INV_X1     g01431(.I(new_n1687_), .ZN(new_n1688_));
  OAI21_X1   g01432(.A1(new_n1556_), .A2(new_n1557_), .B(new_n1432_), .ZN(new_n1689_));
  NOR2_X1    g01433(.A1(new_n1689_), .A2(new_n1553_), .ZN(new_n1690_));
  NOR4_X1    g01434(.A1(new_n1556_), .A2(new_n1557_), .A3(new_n1432_), .A4(\b[18] ), .ZN(new_n1691_));
  OAI21_X1   g01435(.A1(new_n1690_), .A2(new_n1691_), .B(\b[19] ), .ZN(new_n1692_));
  INV_X1     g01436(.I(new_n1692_), .ZN(new_n1693_));
  NOR3_X1    g01437(.A1(new_n1690_), .A2(\b[19] ), .A3(new_n1691_), .ZN(new_n1694_));
  NOR2_X1    g01438(.A1(new_n1693_), .A2(new_n1694_), .ZN(new_n1695_));
  AOI21_X1   g01439(.A1(new_n1695_), .A2(new_n265_), .B(new_n1688_), .ZN(new_n1696_));
  AOI21_X1   g01440(.A1(new_n1696_), .A2(new_n1686_), .B(new_n270_), .ZN(new_n1697_));
  AND3_X2    g01441(.A1(new_n1696_), .A2(new_n270_), .A3(new_n1686_), .Z(new_n1698_));
  NOR2_X1    g01442(.A1(new_n1698_), .A2(new_n1697_), .ZN(new_n1699_));
  AOI21_X1   g01443(.A1(new_n1569_), .A2(new_n1673_), .B(new_n1669_), .ZN(new_n1700_));
  INV_X1     g01444(.I(new_n1306_), .ZN(new_n1701_));
  AOI22_X1   g01445(.A1(new_n800_), .A2(\b[15] ), .B1(\b[16] ), .B2(new_n333_), .ZN(new_n1702_));
  OAI21_X1   g01446(.A1(new_n1093_), .A2(new_n392_), .B(new_n1702_), .ZN(new_n1703_));
  AOI21_X1   g01447(.A1(new_n1701_), .A2(new_n330_), .B(new_n1703_), .ZN(new_n1704_));
  XOR2_X1    g01448(.A1(new_n1704_), .A2(new_n312_), .Z(new_n1705_));
  INV_X1     g01449(.I(new_n1705_), .ZN(new_n1706_));
  NAND3_X1   g01450(.A1(new_n1643_), .A2(new_n1535_), .A3(new_n1647_), .ZN(new_n1707_));
  OAI21_X1   g01451(.A1(new_n1635_), .A2(new_n1648_), .B(new_n1707_), .ZN(new_n1708_));
  AOI21_X1   g01452(.A1(new_n1617_), .A2(new_n1632_), .B(new_n1630_), .ZN(new_n1709_));
  AOI21_X1   g01453(.A1(new_n1475_), .A2(new_n1527_), .B(new_n1514_), .ZN(new_n1710_));
  NOR3_X1    g01454(.A1(new_n1613_), .A2(new_n1612_), .A3(new_n1611_), .ZN(new_n1711_));
  AOI21_X1   g01455(.A1(new_n1604_), .A2(new_n1607_), .B(new_n1583_), .ZN(new_n1712_));
  NOR2_X1    g01456(.A1(new_n1711_), .A2(new_n1712_), .ZN(new_n1713_));
  AOI21_X1   g01457(.A1(new_n1604_), .A2(new_n1607_), .B(new_n1611_), .ZN(new_n1714_));
  INV_X1     g01458(.I(new_n1714_), .ZN(new_n1715_));
  OAI21_X1   g01459(.A1(new_n1713_), .A2(new_n1710_), .B(new_n1715_), .ZN(new_n1716_));
  NOR2_X1    g01460(.A1(new_n1602_), .A2(new_n1601_), .ZN(new_n1717_));
  NAND2_X1   g01461(.A1(new_n1520_), .A2(new_n1599_), .ZN(new_n1718_));
  NOR2_X1    g01462(.A1(new_n1520_), .A2(new_n1599_), .ZN(new_n1719_));
  AOI21_X1   g01463(.A1(new_n1717_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n1720_));
  NOR3_X1    g01464(.A1(new_n1206_), .A2(new_n1345_), .A3(new_n339_), .ZN(new_n1721_));
  NOR2_X1    g01465(.A1(new_n1505_), .A2(new_n290_), .ZN(new_n1722_));
  NOR4_X1    g01466(.A1(new_n1333_), .A2(new_n276_), .A3(new_n1497_), .A4(new_n1507_), .ZN(new_n1723_));
  NOR3_X1    g01467(.A1(new_n1723_), .A2(new_n1722_), .A3(new_n1721_), .ZN(new_n1724_));
  NAND2_X1   g01468(.A1(new_n745_), .A2(new_n746_), .ZN(new_n1725_));
  NAND2_X1   g01469(.A1(new_n1725_), .A2(new_n1354_), .ZN(new_n1726_));
  AOI21_X1   g01470(.A1(new_n1726_), .A2(new_n1724_), .B(new_n1344_), .ZN(new_n1727_));
  NAND3_X1   g01471(.A1(new_n1333_), .A2(new_n1334_), .A3(\b[4] ), .ZN(new_n1728_));
  NAND2_X1   g01472(.A1(new_n1495_), .A2(\b[3] ), .ZN(new_n1729_));
  NAND4_X1   g01473(.A1(new_n1206_), .A2(new_n1498_), .A3(new_n1499_), .A4(\b[2] ), .ZN(new_n1730_));
  NAND3_X1   g01474(.A1(new_n1730_), .A2(new_n1728_), .A3(new_n1729_), .ZN(new_n1731_));
  INV_X1     g01475(.I(new_n1354_), .ZN(new_n1732_));
  NOR2_X1    g01476(.A1(new_n352_), .A2(new_n1732_), .ZN(new_n1733_));
  NOR3_X1    g01477(.A1(new_n1733_), .A2(new_n1731_), .A3(\a[17] ), .ZN(new_n1734_));
  NOR2_X1    g01478(.A1(new_n1727_), .A2(new_n1734_), .ZN(new_n1735_));
  INV_X1     g01479(.I(\a[20] ), .ZN(new_n1736_));
  XOR2_X1    g01480(.A1(\a[19] ), .A2(\a[20] ), .Z(new_n1737_));
  NOR2_X1    g01481(.A1(new_n1597_), .A2(new_n1737_), .ZN(new_n1738_));
  INV_X1     g01482(.I(\a[18] ), .ZN(new_n1739_));
  NAND3_X1   g01483(.A1(new_n1344_), .A2(new_n1739_), .A3(\a[19] ), .ZN(new_n1740_));
  INV_X1     g01484(.I(\a[19] ), .ZN(new_n1741_));
  NAND3_X1   g01485(.A1(new_n1741_), .A2(\a[17] ), .A3(\a[18] ), .ZN(new_n1742_));
  NAND2_X1   g01486(.A1(new_n1740_), .A2(new_n1742_), .ZN(new_n1743_));
  AOI22_X1   g01487(.A1(new_n1738_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n1743_), .ZN(new_n1744_));
  XNOR2_X1   g01488(.A1(\a[19] ), .A2(\a[20] ), .ZN(new_n1745_));
  NOR2_X1    g01489(.A1(new_n1597_), .A2(new_n1745_), .ZN(new_n1746_));
  NAND2_X1   g01490(.A1(new_n1746_), .A2(new_n263_), .ZN(new_n1747_));
  AOI21_X1   g01491(.A1(new_n1744_), .A2(new_n1747_), .B(new_n1736_), .ZN(new_n1748_));
  XOR2_X1    g01492(.A1(\a[17] ), .A2(\a[18] ), .Z(new_n1749_));
  XNOR2_X1   g01493(.A1(\a[19] ), .A2(\a[20] ), .ZN(new_n1750_));
  NAND2_X1   g01494(.A1(new_n1750_), .A2(new_n1749_), .ZN(new_n1751_));
  NOR3_X1    g01495(.A1(new_n1741_), .A2(\a[17] ), .A3(\a[18] ), .ZN(new_n1752_));
  NOR3_X1    g01496(.A1(new_n1344_), .A2(new_n1739_), .A3(\a[19] ), .ZN(new_n1753_));
  NOR2_X1    g01497(.A1(new_n1753_), .A2(new_n1752_), .ZN(new_n1754_));
  OAI22_X1   g01498(.A1(new_n1751_), .A2(new_n275_), .B1(new_n258_), .B2(new_n1754_), .ZN(new_n1755_));
  XOR2_X1    g01499(.A1(\a[19] ), .A2(\a[20] ), .Z(new_n1756_));
  NAND2_X1   g01500(.A1(new_n1749_), .A2(new_n1756_), .ZN(new_n1757_));
  NOR2_X1    g01501(.A1(new_n1757_), .A2(new_n313_), .ZN(new_n1758_));
  NOR3_X1    g01502(.A1(new_n1755_), .A2(new_n1758_), .A3(\a[20] ), .ZN(new_n1759_));
  NOR2_X1    g01503(.A1(new_n1598_), .A2(new_n1736_), .ZN(new_n1760_));
  NOR3_X1    g01504(.A1(new_n1748_), .A2(new_n1759_), .A3(new_n1760_), .ZN(new_n1761_));
  OAI21_X1   g01505(.A1(new_n1755_), .A2(new_n1758_), .B(\a[20] ), .ZN(new_n1762_));
  NOR2_X1    g01506(.A1(new_n1762_), .A2(new_n1598_), .ZN(new_n1763_));
  OAI21_X1   g01507(.A1(new_n1761_), .A2(new_n1763_), .B(new_n1735_), .ZN(new_n1764_));
  OAI21_X1   g01508(.A1(new_n1733_), .A2(new_n1731_), .B(\a[17] ), .ZN(new_n1765_));
  NAND3_X1   g01509(.A1(new_n1726_), .A2(new_n1724_), .A3(new_n1344_), .ZN(new_n1766_));
  NAND2_X1   g01510(.A1(new_n1765_), .A2(new_n1766_), .ZN(new_n1767_));
  NAND3_X1   g01511(.A1(new_n1744_), .A2(new_n1736_), .A3(new_n1747_), .ZN(new_n1768_));
  INV_X1     g01512(.I(new_n1760_), .ZN(new_n1769_));
  NAND3_X1   g01513(.A1(new_n1762_), .A2(new_n1768_), .A3(new_n1769_), .ZN(new_n1770_));
  NAND2_X1   g01514(.A1(new_n1748_), .A2(new_n1599_), .ZN(new_n1771_));
  NAND3_X1   g01515(.A1(new_n1767_), .A2(new_n1770_), .A3(new_n1771_), .ZN(new_n1772_));
  AOI21_X1   g01516(.A1(new_n1764_), .A2(new_n1772_), .B(new_n1720_), .ZN(new_n1773_));
  NAND2_X1   g01517(.A1(new_n1591_), .A2(new_n1596_), .ZN(new_n1774_));
  NOR2_X1    g01518(.A1(new_n1513_), .A2(new_n1598_), .ZN(new_n1775_));
  NAND2_X1   g01519(.A1(new_n1513_), .A2(new_n1598_), .ZN(new_n1776_));
  OAI21_X1   g01520(.A1(new_n1774_), .A2(new_n1775_), .B(new_n1776_), .ZN(new_n1777_));
  AOI21_X1   g01521(.A1(new_n1770_), .A2(new_n1771_), .B(new_n1767_), .ZN(new_n1778_));
  NOR3_X1    g01522(.A1(new_n1735_), .A2(new_n1761_), .A3(new_n1763_), .ZN(new_n1779_));
  NOR3_X1    g01523(.A1(new_n1777_), .A2(new_n1778_), .A3(new_n1779_), .ZN(new_n1780_));
  NOR2_X1    g01524(.A1(new_n1773_), .A2(new_n1780_), .ZN(new_n1781_));
  OAI22_X1   g01525(.A1(new_n993_), .A2(new_n471_), .B1(new_n438_), .B2(new_n997_), .ZN(new_n1782_));
  AOI21_X1   g01526(.A1(\b[5] ), .A2(new_n1486_), .B(new_n1782_), .ZN(new_n1783_));
  NAND3_X1   g01527(.A1(new_n484_), .A2(new_n477_), .A3(new_n1013_), .ZN(new_n1784_));
  AOI21_X1   g01528(.A1(new_n1784_), .A2(new_n1783_), .B(new_n1002_), .ZN(new_n1785_));
  INV_X1     g01529(.I(new_n1785_), .ZN(new_n1786_));
  NAND3_X1   g01530(.A1(new_n1784_), .A2(new_n1002_), .A3(new_n1783_), .ZN(new_n1787_));
  NAND2_X1   g01531(.A1(new_n1786_), .A2(new_n1787_), .ZN(new_n1788_));
  NAND2_X1   g01532(.A1(new_n1781_), .A2(new_n1788_), .ZN(new_n1789_));
  OAI21_X1   g01533(.A1(new_n1778_), .A2(new_n1779_), .B(new_n1777_), .ZN(new_n1790_));
  NAND3_X1   g01534(.A1(new_n1720_), .A2(new_n1764_), .A3(new_n1772_), .ZN(new_n1791_));
  NAND2_X1   g01535(.A1(new_n1790_), .A2(new_n1791_), .ZN(new_n1792_));
  INV_X1     g01536(.I(new_n1787_), .ZN(new_n1793_));
  NOR2_X1    g01537(.A1(new_n1793_), .A2(new_n1785_), .ZN(new_n1794_));
  NAND2_X1   g01538(.A1(new_n1792_), .A2(new_n1794_), .ZN(new_n1795_));
  NAND2_X1   g01539(.A1(new_n1789_), .A2(new_n1795_), .ZN(new_n1796_));
  NAND2_X1   g01540(.A1(new_n1796_), .A2(new_n1716_), .ZN(new_n1797_));
  NOR2_X1    g01541(.A1(new_n1796_), .A2(new_n1716_), .ZN(new_n1798_));
  INV_X1     g01542(.I(new_n1798_), .ZN(new_n1799_));
  OAI22_X1   g01543(.A1(new_n713_), .A2(new_n776_), .B1(new_n667_), .B2(new_n717_), .ZN(new_n1800_));
  AOI21_X1   g01544(.A1(\b[8] ), .A2(new_n1126_), .B(new_n1800_), .ZN(new_n1801_));
  OAI21_X1   g01545(.A1(new_n786_), .A2(new_n986_), .B(new_n1801_), .ZN(new_n1802_));
  XOR2_X1    g01546(.A1(new_n1802_), .A2(new_n722_), .Z(new_n1803_));
  NAND3_X1   g01547(.A1(new_n1799_), .A2(new_n1803_), .A3(new_n1797_), .ZN(new_n1804_));
  INV_X1     g01548(.I(new_n1797_), .ZN(new_n1805_));
  XOR2_X1    g01549(.A1(new_n1802_), .A2(\a[11] ), .Z(new_n1806_));
  OAI21_X1   g01550(.A1(new_n1805_), .A2(new_n1798_), .B(new_n1806_), .ZN(new_n1807_));
  NAND2_X1   g01551(.A1(new_n1807_), .A2(new_n1804_), .ZN(new_n1808_));
  NAND2_X1   g01552(.A1(new_n1709_), .A2(new_n1808_), .ZN(new_n1809_));
  OAI21_X1   g01553(.A1(new_n1628_), .A2(new_n1616_), .B(new_n1633_), .ZN(new_n1810_));
  NAND3_X1   g01554(.A1(new_n1810_), .A2(new_n1804_), .A3(new_n1807_), .ZN(new_n1811_));
  OAI22_X1   g01555(.A1(new_n610_), .A2(new_n1070_), .B1(new_n941_), .B2(new_n612_), .ZN(new_n1812_));
  AOI21_X1   g01556(.A1(\b[11] ), .A2(new_n826_), .B(new_n1812_), .ZN(new_n1813_));
  OAI21_X1   g01557(.A1(new_n1082_), .A2(new_n624_), .B(new_n1813_), .ZN(new_n1814_));
  NAND2_X1   g01558(.A1(new_n1814_), .A2(\a[8] ), .ZN(new_n1815_));
  INV_X1     g01559(.I(new_n1078_), .ZN(new_n1816_));
  NOR4_X1    g01560(.A1(new_n1077_), .A2(new_n1073_), .A3(new_n1074_), .A4(new_n1076_), .ZN(new_n1817_));
  NOR2_X1    g01561(.A1(new_n1816_), .A2(new_n1817_), .ZN(new_n1818_));
  NAND2_X1   g01562(.A1(new_n1818_), .A2(new_n618_), .ZN(new_n1819_));
  NAND3_X1   g01563(.A1(new_n1819_), .A2(new_n488_), .A3(new_n1813_), .ZN(new_n1820_));
  NAND2_X1   g01564(.A1(new_n1820_), .A2(new_n1815_), .ZN(new_n1821_));
  NAND3_X1   g01565(.A1(new_n1821_), .A2(new_n1809_), .A3(new_n1811_), .ZN(new_n1822_));
  INV_X1     g01566(.I(new_n1822_), .ZN(new_n1823_));
  AOI21_X1   g01567(.A1(new_n1809_), .A2(new_n1811_), .B(new_n1821_), .ZN(new_n1824_));
  NOR2_X1    g01568(.A1(new_n1823_), .A2(new_n1824_), .ZN(new_n1825_));
  NAND2_X1   g01569(.A1(new_n1825_), .A2(new_n1708_), .ZN(new_n1826_));
  INV_X1     g01570(.I(new_n1635_), .ZN(new_n1827_));
  OAI21_X1   g01571(.A1(new_n1659_), .A2(new_n1640_), .B(new_n1660_), .ZN(new_n1828_));
  AOI21_X1   g01572(.A1(new_n1827_), .A2(new_n1828_), .B(new_n1661_), .ZN(new_n1829_));
  NAND2_X1   g01573(.A1(new_n1809_), .A2(new_n1811_), .ZN(new_n1830_));
  NAND3_X1   g01574(.A1(new_n1830_), .A2(new_n1815_), .A3(new_n1820_), .ZN(new_n1831_));
  NAND2_X1   g01575(.A1(new_n1831_), .A2(new_n1822_), .ZN(new_n1832_));
  NAND2_X1   g01576(.A1(new_n1832_), .A2(new_n1829_), .ZN(new_n1833_));
  NAND2_X1   g01577(.A1(new_n1826_), .A2(new_n1833_), .ZN(new_n1834_));
  NOR2_X1    g01578(.A1(new_n1834_), .A2(new_n1706_), .ZN(new_n1835_));
  NOR2_X1    g01579(.A1(new_n1832_), .A2(new_n1829_), .ZN(new_n1836_));
  NOR2_X1    g01580(.A1(new_n1825_), .A2(new_n1708_), .ZN(new_n1837_));
  NOR2_X1    g01581(.A1(new_n1837_), .A2(new_n1836_), .ZN(new_n1838_));
  NOR2_X1    g01582(.A1(new_n1838_), .A2(new_n1705_), .ZN(new_n1839_));
  NOR2_X1    g01583(.A1(new_n1839_), .A2(new_n1835_), .ZN(new_n1840_));
  XOR2_X1    g01584(.A1(new_n1700_), .A2(new_n1840_), .Z(new_n1841_));
  NOR2_X1    g01585(.A1(new_n1841_), .A2(new_n1699_), .ZN(new_n1842_));
  NAND2_X1   g01586(.A1(new_n1841_), .A2(new_n1699_), .ZN(new_n1843_));
  INV_X1     g01587(.I(new_n1843_), .ZN(new_n1844_));
  NOR2_X1    g01588(.A1(new_n1844_), .A2(new_n1842_), .ZN(new_n1845_));
  INV_X1     g01589(.I(new_n1267_), .ZN(new_n1846_));
  AOI21_X1   g01590(.A1(new_n1289_), .A2(new_n1290_), .B(new_n1283_), .ZN(new_n1847_));
  OAI21_X1   g01591(.A1(new_n1846_), .A2(new_n1847_), .B(new_n1291_), .ZN(new_n1848_));
  OAI21_X1   g01592(.A1(new_n1848_), .A2(new_n1425_), .B(new_n1426_), .ZN(new_n1849_));
  INV_X1     g01593(.I(new_n1547_), .ZN(new_n1850_));
  AOI21_X1   g01594(.A1(new_n1849_), .A2(new_n1850_), .B(new_n1550_), .ZN(new_n1851_));
  NOR2_X1    g01595(.A1(new_n1672_), .A2(new_n1682_), .ZN(new_n1852_));
  NOR2_X1    g01596(.A1(new_n1681_), .A2(new_n1566_), .ZN(new_n1853_));
  INV_X1     g01597(.I(new_n1853_), .ZN(new_n1854_));
  OAI21_X1   g01598(.A1(new_n1851_), .A2(new_n1852_), .B(new_n1854_), .ZN(new_n1855_));
  XOR2_X1    g01599(.A1(new_n1855_), .A2(new_n1845_), .Z(\f[19] ));
  AOI21_X1   g01600(.A1(new_n1552_), .A2(new_n1683_), .B(new_n1853_), .ZN(new_n1857_));
  OAI21_X1   g01601(.A1(new_n1857_), .A2(new_n1842_), .B(new_n1843_), .ZN(new_n1858_));
  INV_X1     g01602(.I(\b[19] ), .ZN(new_n1859_));
  INV_X1     g01603(.I(\b[20] ), .ZN(new_n1860_));
  OAI22_X1   g01604(.A1(new_n277_), .A2(new_n1860_), .B1(new_n1859_), .B2(new_n262_), .ZN(new_n1861_));
  AOI21_X1   g01605(.A1(\b[18] ), .A2(new_n283_), .B(new_n1861_), .ZN(new_n1862_));
  XOR2_X1    g01606(.A1(\b[19] ), .A2(\b[20] ), .Z(new_n1863_));
  NOR3_X1    g01607(.A1(new_n1556_), .A2(new_n1557_), .A3(new_n1432_), .ZN(new_n1864_));
  OAI21_X1   g01608(.A1(new_n1864_), .A2(\b[18] ), .B(\b[19] ), .ZN(new_n1865_));
  NAND2_X1   g01609(.A1(new_n1689_), .A2(\b[18] ), .ZN(new_n1866_));
  AOI21_X1   g01610(.A1(new_n1865_), .A2(new_n1866_), .B(new_n1863_), .ZN(new_n1867_));
  INV_X1     g01611(.I(new_n1863_), .ZN(new_n1868_));
  NAND2_X1   g01612(.A1(new_n1865_), .A2(new_n1866_), .ZN(new_n1869_));
  NOR2_X1    g01613(.A1(new_n1869_), .A2(new_n1868_), .ZN(new_n1870_));
  NOR2_X1    g01614(.A1(new_n1870_), .A2(new_n1867_), .ZN(new_n1871_));
  OAI21_X1   g01615(.A1(new_n1871_), .A2(new_n279_), .B(new_n1862_), .ZN(new_n1872_));
  XOR2_X1    g01616(.A1(new_n1872_), .A2(\a[2] ), .Z(new_n1873_));
  INV_X1     g01617(.I(new_n1873_), .ZN(new_n1874_));
  OAI22_X1   g01618(.A1(new_n321_), .A2(new_n1432_), .B1(new_n325_), .B2(new_n1296_), .ZN(new_n1875_));
  AOI21_X1   g01619(.A1(\b[15] ), .A2(new_n602_), .B(new_n1875_), .ZN(new_n1876_));
  OAI21_X1   g01620(.A1(new_n1444_), .A2(new_n318_), .B(new_n1876_), .ZN(new_n1877_));
  XOR2_X1    g01621(.A1(new_n1877_), .A2(\a[5] ), .Z(new_n1878_));
  AOI22_X1   g01622(.A1(new_n518_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n636_), .ZN(new_n1879_));
  OAI21_X1   g01623(.A1(new_n941_), .A2(new_n917_), .B(new_n1879_), .ZN(new_n1880_));
  INV_X1     g01624(.I(new_n1880_), .ZN(new_n1881_));
  OAI21_X1   g01625(.A1(new_n1100_), .A2(new_n1102_), .B(new_n618_), .ZN(new_n1882_));
  AOI21_X1   g01626(.A1(new_n1882_), .A2(new_n1881_), .B(new_n488_), .ZN(new_n1883_));
  INV_X1     g01627(.I(new_n1883_), .ZN(new_n1884_));
  NAND3_X1   g01628(.A1(new_n1882_), .A2(new_n488_), .A3(new_n1881_), .ZN(new_n1885_));
  NAND2_X1   g01629(.A1(new_n1884_), .A2(new_n1885_), .ZN(new_n1886_));
  NOR3_X1    g01630(.A1(new_n1805_), .A2(new_n1806_), .A3(new_n1798_), .ZN(new_n1887_));
  NOR2_X1    g01631(.A1(new_n1531_), .A2(new_n1382_), .ZN(new_n1888_));
  NOR2_X1    g01632(.A1(new_n1532_), .A2(new_n1533_), .ZN(new_n1889_));
  AOI21_X1   g01633(.A1(new_n1888_), .A2(new_n1889_), .B(new_n1626_), .ZN(new_n1890_));
  OAI21_X1   g01634(.A1(new_n1890_), .A2(new_n1622_), .B(new_n1617_), .ZN(new_n1891_));
  AOI21_X1   g01635(.A1(new_n1799_), .A2(new_n1797_), .B(new_n1803_), .ZN(new_n1892_));
  AOI21_X1   g01636(.A1(new_n1891_), .A2(new_n1633_), .B(new_n1892_), .ZN(new_n1893_));
  AOI22_X1   g01637(.A1(new_n729_), .A2(\b[11] ), .B1(\b[10] ), .B2(new_n732_), .ZN(new_n1894_));
  OAI21_X1   g01638(.A1(new_n667_), .A2(new_n1127_), .B(new_n1894_), .ZN(new_n1895_));
  NOR3_X1    g01639(.A1(new_n1459_), .A2(new_n986_), .A3(new_n1460_), .ZN(new_n1896_));
  OAI21_X1   g01640(.A1(new_n1896_), .A2(new_n1895_), .B(\a[11] ), .ZN(new_n1897_));
  NOR3_X1    g01641(.A1(new_n1896_), .A2(\a[11] ), .A3(new_n1895_), .ZN(new_n1898_));
  INV_X1     g01642(.I(new_n1898_), .ZN(new_n1899_));
  AOI21_X1   g01643(.A1(new_n1615_), .A2(new_n1574_), .B(new_n1714_), .ZN(new_n1900_));
  NOR2_X1    g01644(.A1(new_n1792_), .A2(new_n1794_), .ZN(new_n1901_));
  AOI21_X1   g01645(.A1(new_n1900_), .A2(new_n1795_), .B(new_n1901_), .ZN(new_n1902_));
  OAI22_X1   g01646(.A1(new_n993_), .A2(new_n577_), .B1(new_n471_), .B2(new_n997_), .ZN(new_n1903_));
  AOI21_X1   g01647(.A1(\b[6] ), .A2(new_n1486_), .B(new_n1903_), .ZN(new_n1904_));
  OAI21_X1   g01648(.A1(new_n586_), .A2(new_n584_), .B(new_n1013_), .ZN(new_n1905_));
  AOI21_X1   g01649(.A1(new_n1905_), .A2(new_n1904_), .B(new_n1002_), .ZN(new_n1906_));
  INV_X1     g01650(.I(new_n1904_), .ZN(new_n1907_));
  AOI21_X1   g01651(.A1(new_n798_), .A2(new_n585_), .B(new_n1323_), .ZN(new_n1908_));
  NOR3_X1    g01652(.A1(new_n1908_), .A2(\a[14] ), .A3(new_n1907_), .ZN(new_n1909_));
  AOI21_X1   g01653(.A1(new_n1777_), .A2(new_n1772_), .B(new_n1778_), .ZN(new_n1910_));
  NOR3_X1    g01654(.A1(new_n1910_), .A2(new_n1909_), .A3(new_n1906_), .ZN(new_n1911_));
  OAI21_X1   g01655(.A1(new_n1908_), .A2(new_n1907_), .B(\a[14] ), .ZN(new_n1912_));
  NAND3_X1   g01656(.A1(new_n1905_), .A2(new_n1002_), .A3(new_n1904_), .ZN(new_n1913_));
  OAI21_X1   g01657(.A1(new_n1720_), .A2(new_n1779_), .B(new_n1764_), .ZN(new_n1914_));
  AOI21_X1   g01658(.A1(new_n1912_), .A2(new_n1913_), .B(new_n1914_), .ZN(new_n1915_));
  OAI22_X1   g01659(.A1(new_n1592_), .A2(new_n377_), .B1(new_n339_), .B2(new_n1505_), .ZN(new_n1916_));
  NAND3_X1   g01660(.A1(new_n1206_), .A2(new_n1498_), .A3(new_n1499_), .ZN(new_n1917_));
  NOR2_X1    g01661(.A1(new_n1917_), .A2(new_n290_), .ZN(new_n1918_));
  NOR2_X1    g01662(.A1(new_n1916_), .A2(new_n1918_), .ZN(new_n1919_));
  OAI21_X1   g01663(.A1(new_n566_), .A2(new_n1732_), .B(new_n1919_), .ZN(new_n1920_));
  NAND2_X1   g01664(.A1(new_n1920_), .A2(\a[17] ), .ZN(new_n1921_));
  NAND2_X1   g01665(.A1(new_n382_), .A2(new_n1354_), .ZN(new_n1922_));
  NAND3_X1   g01666(.A1(new_n1922_), .A2(new_n1344_), .A3(new_n1919_), .ZN(new_n1923_));
  NAND2_X1   g01667(.A1(new_n1762_), .A2(new_n1768_), .ZN(new_n1924_));
  NOR2_X1    g01668(.A1(new_n1757_), .A2(new_n282_), .ZN(new_n1925_));
  NOR2_X1    g01669(.A1(new_n1751_), .A2(new_n276_), .ZN(new_n1926_));
  NOR2_X1    g01670(.A1(new_n1754_), .A2(new_n275_), .ZN(new_n1927_));
  AOI21_X1   g01671(.A1(new_n1741_), .A2(\a[20] ), .B(\a[17] ), .ZN(new_n1928_));
  INV_X1     g01672(.I(new_n1928_), .ZN(new_n1929_));
  OAI21_X1   g01673(.A1(new_n1741_), .A2(\a[20] ), .B(\a[17] ), .ZN(new_n1930_));
  NAND3_X1   g01674(.A1(new_n1929_), .A2(new_n1597_), .A3(new_n1930_), .ZN(new_n1931_));
  NOR2_X1    g01675(.A1(new_n1931_), .A2(new_n258_), .ZN(new_n1932_));
  NOR4_X1    g01676(.A1(new_n1932_), .A2(new_n1925_), .A3(new_n1926_), .A4(new_n1927_), .ZN(new_n1933_));
  NOR2_X1    g01677(.A1(new_n1933_), .A2(new_n1736_), .ZN(new_n1934_));
  NAND2_X1   g01678(.A1(new_n1746_), .A2(new_n554_), .ZN(new_n1935_));
  NAND2_X1   g01679(.A1(new_n1738_), .A2(\b[2] ), .ZN(new_n1936_));
  NAND2_X1   g01680(.A1(new_n1743_), .A2(\b[1] ), .ZN(new_n1937_));
  AOI21_X1   g01681(.A1(\a[19] ), .A2(new_n1736_), .B(new_n1344_), .ZN(new_n1938_));
  NOR3_X1    g01682(.A1(new_n1749_), .A2(new_n1928_), .A3(new_n1938_), .ZN(new_n1939_));
  NAND2_X1   g01683(.A1(new_n1939_), .A2(\b[0] ), .ZN(new_n1940_));
  NAND4_X1   g01684(.A1(new_n1935_), .A2(new_n1940_), .A3(new_n1936_), .A4(new_n1937_), .ZN(new_n1941_));
  NOR2_X1    g01685(.A1(new_n1941_), .A2(\a[20] ), .ZN(new_n1942_));
  OAI22_X1   g01686(.A1(new_n1924_), .A2(new_n1769_), .B1(new_n1934_), .B2(new_n1942_), .ZN(new_n1943_));
  NOR2_X1    g01687(.A1(new_n1755_), .A2(new_n1758_), .ZN(new_n1944_));
  NAND4_X1   g01688(.A1(new_n1933_), .A2(\a[20] ), .A3(new_n1944_), .A4(new_n1599_), .ZN(new_n1945_));
  NAND4_X1   g01689(.A1(new_n1943_), .A2(new_n1923_), .A3(new_n1921_), .A4(new_n1945_), .ZN(new_n1946_));
  INV_X1     g01690(.I(new_n1921_), .ZN(new_n1947_));
  NOR2_X1    g01691(.A1(new_n1920_), .A2(\a[17] ), .ZN(new_n1948_));
  NOR2_X1    g01692(.A1(new_n1748_), .A2(new_n1759_), .ZN(new_n1949_));
  NAND2_X1   g01693(.A1(new_n1941_), .A2(\a[20] ), .ZN(new_n1950_));
  NAND2_X1   g01694(.A1(new_n1933_), .A2(new_n1736_), .ZN(new_n1951_));
  AOI22_X1   g01695(.A1(new_n1949_), .A2(new_n1760_), .B1(new_n1951_), .B2(new_n1950_), .ZN(new_n1952_));
  NAND2_X1   g01696(.A1(new_n1744_), .A2(new_n1747_), .ZN(new_n1953_));
  NOR4_X1    g01697(.A1(new_n1941_), .A2(new_n1953_), .A3(new_n1736_), .A4(new_n1598_), .ZN(new_n1954_));
  OAI22_X1   g01698(.A1(new_n1947_), .A2(new_n1948_), .B1(new_n1952_), .B2(new_n1954_), .ZN(new_n1955_));
  NAND2_X1   g01699(.A1(new_n1955_), .A2(new_n1946_), .ZN(new_n1956_));
  NOR3_X1    g01700(.A1(new_n1915_), .A2(new_n1911_), .A3(new_n1956_), .ZN(new_n1957_));
  NAND3_X1   g01701(.A1(new_n1914_), .A2(new_n1912_), .A3(new_n1913_), .ZN(new_n1958_));
  OAI21_X1   g01702(.A1(new_n1906_), .A2(new_n1909_), .B(new_n1910_), .ZN(new_n1959_));
  NOR4_X1    g01703(.A1(new_n1947_), .A2(new_n1948_), .A3(new_n1952_), .A4(new_n1954_), .ZN(new_n1960_));
  AOI22_X1   g01704(.A1(new_n1943_), .A2(new_n1945_), .B1(new_n1923_), .B2(new_n1921_), .ZN(new_n1961_));
  NOR2_X1    g01705(.A1(new_n1960_), .A2(new_n1961_), .ZN(new_n1962_));
  AOI21_X1   g01706(.A1(new_n1959_), .A2(new_n1958_), .B(new_n1962_), .ZN(new_n1963_));
  NOR2_X1    g01707(.A1(new_n1957_), .A2(new_n1963_), .ZN(new_n1964_));
  NAND2_X1   g01708(.A1(new_n1964_), .A2(new_n1902_), .ZN(new_n1965_));
  NOR2_X1    g01709(.A1(new_n1781_), .A2(new_n1788_), .ZN(new_n1966_));
  OAI21_X1   g01710(.A1(new_n1716_), .A2(new_n1966_), .B(new_n1789_), .ZN(new_n1967_));
  NAND3_X1   g01711(.A1(new_n1959_), .A2(new_n1958_), .A3(new_n1962_), .ZN(new_n1968_));
  OAI21_X1   g01712(.A1(new_n1915_), .A2(new_n1911_), .B(new_n1956_), .ZN(new_n1969_));
  NAND2_X1   g01713(.A1(new_n1969_), .A2(new_n1968_), .ZN(new_n1970_));
  NAND2_X1   g01714(.A1(new_n1967_), .A2(new_n1970_), .ZN(new_n1971_));
  NAND4_X1   g01715(.A1(new_n1965_), .A2(new_n1971_), .A3(new_n1899_), .A4(new_n1897_), .ZN(new_n1972_));
  INV_X1     g01716(.I(new_n1897_), .ZN(new_n1973_));
  NOR2_X1    g01717(.A1(new_n1967_), .A2(new_n1970_), .ZN(new_n1974_));
  NOR2_X1    g01718(.A1(new_n1964_), .A2(new_n1902_), .ZN(new_n1975_));
  OAI22_X1   g01719(.A1(new_n1974_), .A2(new_n1975_), .B1(new_n1973_), .B2(new_n1898_), .ZN(new_n1976_));
  NAND2_X1   g01720(.A1(new_n1976_), .A2(new_n1972_), .ZN(new_n1977_));
  NOR3_X1    g01721(.A1(new_n1893_), .A2(new_n1887_), .A3(new_n1977_), .ZN(new_n1978_));
  NAND2_X1   g01722(.A1(new_n1466_), .A2(new_n1393_), .ZN(new_n1979_));
  OAI21_X1   g01723(.A1(new_n1979_), .A2(new_n1538_), .B(new_n1627_), .ZN(new_n1980_));
  AOI21_X1   g01724(.A1(new_n1980_), .A2(new_n1629_), .B(new_n1616_), .ZN(new_n1981_));
  OAI21_X1   g01725(.A1(new_n1981_), .A2(new_n1630_), .B(new_n1807_), .ZN(new_n1982_));
  NOR4_X1    g01726(.A1(new_n1974_), .A2(new_n1975_), .A3(new_n1973_), .A4(new_n1898_), .ZN(new_n1983_));
  AOI22_X1   g01727(.A1(new_n1971_), .A2(new_n1965_), .B1(new_n1899_), .B2(new_n1897_), .ZN(new_n1984_));
  NOR2_X1    g01728(.A1(new_n1984_), .A2(new_n1983_), .ZN(new_n1985_));
  AOI21_X1   g01729(.A1(new_n1982_), .A2(new_n1804_), .B(new_n1985_), .ZN(new_n1986_));
  OAI21_X1   g01730(.A1(new_n1978_), .A2(new_n1986_), .B(new_n1886_), .ZN(new_n1987_));
  INV_X1     g01731(.I(new_n1885_), .ZN(new_n1988_));
  NOR2_X1    g01732(.A1(new_n1988_), .A2(new_n1883_), .ZN(new_n1989_));
  NAND3_X1   g01733(.A1(new_n1982_), .A2(new_n1804_), .A3(new_n1985_), .ZN(new_n1990_));
  OAI21_X1   g01734(.A1(new_n1893_), .A2(new_n1887_), .B(new_n1977_), .ZN(new_n1991_));
  NAND3_X1   g01735(.A1(new_n1991_), .A2(new_n1990_), .A3(new_n1989_), .ZN(new_n1992_));
  NAND2_X1   g01736(.A1(new_n1987_), .A2(new_n1992_), .ZN(new_n1993_));
  AOI21_X1   g01737(.A1(new_n1456_), .A2(new_n1642_), .B(new_n1640_), .ZN(new_n1994_));
  OAI21_X1   g01738(.A1(new_n1994_), .A2(new_n1647_), .B(new_n1827_), .ZN(new_n1995_));
  NAND3_X1   g01739(.A1(new_n1995_), .A2(new_n1707_), .A3(new_n1822_), .ZN(new_n1996_));
  AOI21_X1   g01740(.A1(new_n1996_), .A2(new_n1831_), .B(new_n1993_), .ZN(new_n1997_));
  INV_X1     g01741(.I(new_n1997_), .ZN(new_n1998_));
  AOI21_X1   g01742(.A1(new_n1829_), .A2(new_n1822_), .B(new_n1824_), .ZN(new_n1999_));
  NAND2_X1   g01743(.A1(new_n1999_), .A2(new_n1993_), .ZN(new_n2000_));
  NAND2_X1   g01744(.A1(new_n1998_), .A2(new_n2000_), .ZN(new_n2001_));
  INV_X1     g01745(.I(new_n2001_), .ZN(new_n2002_));
  NOR2_X1    g01746(.A1(new_n2002_), .A2(new_n1878_), .ZN(new_n2003_));
  NAND2_X1   g01747(.A1(new_n2002_), .A2(new_n1878_), .ZN(new_n2004_));
  INV_X1     g01748(.I(new_n2004_), .ZN(new_n2005_));
  OAI21_X1   g01749(.A1(new_n1679_), .A2(new_n1666_), .B(new_n1674_), .ZN(new_n2006_));
  INV_X1     g01750(.I(new_n1840_), .ZN(new_n2007_));
  NOR2_X1    g01751(.A1(new_n1838_), .A2(new_n1706_), .ZN(new_n2008_));
  AOI21_X1   g01752(.A1(new_n2006_), .A2(new_n2007_), .B(new_n2008_), .ZN(new_n2009_));
  NOR3_X1    g01753(.A1(new_n2009_), .A2(new_n2003_), .A3(new_n2005_), .ZN(new_n2010_));
  INV_X1     g01754(.I(new_n2003_), .ZN(new_n2011_));
  INV_X1     g01755(.I(new_n2008_), .ZN(new_n2012_));
  OAI21_X1   g01756(.A1(new_n1700_), .A2(new_n1840_), .B(new_n2012_), .ZN(new_n2013_));
  AOI21_X1   g01757(.A1(new_n2011_), .A2(new_n2004_), .B(new_n2013_), .ZN(new_n2014_));
  NOR3_X1    g01758(.A1(new_n2010_), .A2(new_n2014_), .A3(new_n1874_), .ZN(new_n2015_));
  NOR2_X1    g01759(.A1(new_n2010_), .A2(new_n2014_), .ZN(new_n2016_));
  NOR2_X1    g01760(.A1(new_n2016_), .A2(new_n1873_), .ZN(new_n2017_));
  NOR2_X1    g01761(.A1(new_n2017_), .A2(new_n2015_), .ZN(new_n2018_));
  XOR2_X1    g01762(.A1(new_n1858_), .A2(new_n2018_), .Z(\f[20] ));
  AOI21_X1   g01763(.A1(new_n1858_), .A2(new_n2018_), .B(new_n2015_), .ZN(new_n2020_));
  NAND2_X1   g01764(.A1(new_n283_), .A2(\b[19] ), .ZN(new_n2021_));
  AOI22_X1   g01765(.A1(new_n267_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n261_), .ZN(new_n2022_));
  INV_X1     g01766(.I(new_n2022_), .ZN(new_n2023_));
  AOI21_X1   g01767(.A1(new_n1869_), .A2(\b[20] ), .B(new_n1859_), .ZN(new_n2024_));
  NOR2_X1    g01768(.A1(new_n1869_), .A2(\b[20] ), .ZN(new_n2025_));
  NOR2_X1    g01769(.A1(new_n2024_), .A2(new_n2025_), .ZN(new_n2026_));
  INV_X1     g01770(.I(\b[21] ), .ZN(new_n2027_));
  NAND3_X1   g01771(.A1(new_n1865_), .A2(new_n1866_), .A3(new_n2027_), .ZN(new_n2028_));
  NAND2_X1   g01772(.A1(new_n1869_), .A2(\b[21] ), .ZN(new_n2029_));
  AOI21_X1   g01773(.A1(new_n2028_), .A2(new_n2029_), .B(new_n2026_), .ZN(new_n2030_));
  AND3_X2    g01774(.A1(new_n2026_), .A2(new_n2028_), .A3(new_n2029_), .Z(new_n2031_));
  NOR2_X1    g01775(.A1(new_n2031_), .A2(new_n2030_), .ZN(new_n2032_));
  AOI21_X1   g01776(.A1(new_n2032_), .A2(new_n265_), .B(new_n2023_), .ZN(new_n2033_));
  AOI21_X1   g01777(.A1(new_n2033_), .A2(new_n2021_), .B(new_n270_), .ZN(new_n2034_));
  NAND2_X1   g01778(.A1(new_n2033_), .A2(new_n2021_), .ZN(new_n2035_));
  NOR2_X1    g01779(.A1(new_n2035_), .A2(\a[2] ), .ZN(new_n2036_));
  NOR2_X1    g01780(.A1(new_n2036_), .A2(new_n2034_), .ZN(new_n2037_));
  INV_X1     g01781(.I(new_n1563_), .ZN(new_n2038_));
  AOI22_X1   g01782(.A1(new_n800_), .A2(\b[17] ), .B1(\b[18] ), .B2(new_n333_), .ZN(new_n2039_));
  OAI21_X1   g01783(.A1(new_n1296_), .A2(new_n392_), .B(new_n2039_), .ZN(new_n2040_));
  AOI21_X1   g01784(.A1(new_n2038_), .A2(new_n330_), .B(new_n2040_), .ZN(new_n2041_));
  XOR2_X1    g01785(.A1(new_n2041_), .A2(new_n312_), .Z(new_n2042_));
  OAI21_X1   g01786(.A1(new_n1910_), .A2(new_n1961_), .B(new_n1946_), .ZN(new_n2043_));
  AOI22_X1   g01787(.A1(new_n1586_), .A2(\b[6] ), .B1(\b[5] ), .B2(new_n1495_), .ZN(new_n2044_));
  OAI21_X1   g01788(.A1(new_n339_), .A2(new_n1917_), .B(new_n2044_), .ZN(new_n2045_));
  AOI21_X1   g01789(.A1(new_n916_), .A2(new_n1354_), .B(new_n2045_), .ZN(new_n2046_));
  NOR2_X1    g01790(.A1(new_n2046_), .A2(new_n1344_), .ZN(new_n2047_));
  NOR2_X1    g01791(.A1(new_n450_), .A2(new_n1732_), .ZN(new_n2048_));
  NOR3_X1    g01792(.A1(new_n2048_), .A2(\a[17] ), .A3(new_n2045_), .ZN(new_n2049_));
  NOR2_X1    g01793(.A1(new_n2047_), .A2(new_n2049_), .ZN(new_n2050_));
  NAND2_X1   g01794(.A1(new_n1939_), .A2(\b[1] ), .ZN(new_n2051_));
  AOI22_X1   g01795(.A1(new_n1738_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n1743_), .ZN(new_n2052_));
  NAND2_X1   g01796(.A1(new_n299_), .A2(new_n1746_), .ZN(new_n2053_));
  NAND3_X1   g01797(.A1(new_n2053_), .A2(new_n2052_), .A3(new_n2051_), .ZN(new_n2054_));
  NAND2_X1   g01798(.A1(new_n2054_), .A2(\a[20] ), .ZN(new_n2055_));
  NOR2_X1    g01799(.A1(new_n1931_), .A2(new_n275_), .ZN(new_n2056_));
  OAI22_X1   g01800(.A1(new_n1751_), .A2(new_n290_), .B1(new_n276_), .B2(new_n1754_), .ZN(new_n2057_));
  NOR2_X1    g01801(.A1(new_n429_), .A2(new_n1757_), .ZN(new_n2058_));
  NOR3_X1    g01802(.A1(new_n2058_), .A2(new_n2057_), .A3(new_n2056_), .ZN(new_n2059_));
  NAND2_X1   g01803(.A1(new_n2059_), .A2(new_n1736_), .ZN(new_n2060_));
  XNOR2_X1   g01804(.A1(\a[20] ), .A2(\a[21] ), .ZN(new_n2061_));
  NOR2_X1    g01805(.A1(new_n2061_), .A2(new_n258_), .ZN(new_n2062_));
  INV_X1     g01806(.I(new_n2062_), .ZN(new_n2063_));
  AOI21_X1   g01807(.A1(new_n2060_), .A2(new_n2055_), .B(new_n2063_), .ZN(new_n2064_));
  NOR2_X1    g01808(.A1(new_n2059_), .A2(new_n1736_), .ZN(new_n2065_));
  NOR2_X1    g01809(.A1(new_n2054_), .A2(\a[20] ), .ZN(new_n2066_));
  NOR3_X1    g01810(.A1(new_n2065_), .A2(new_n2066_), .A3(new_n2062_), .ZN(new_n2067_));
  OAI21_X1   g01811(.A1(new_n2064_), .A2(new_n2067_), .B(new_n1945_), .ZN(new_n2068_));
  OAI21_X1   g01812(.A1(new_n2065_), .A2(new_n2066_), .B(new_n2062_), .ZN(new_n2069_));
  NAND3_X1   g01813(.A1(new_n2060_), .A2(new_n2055_), .A3(new_n2063_), .ZN(new_n2070_));
  NAND3_X1   g01814(.A1(new_n2069_), .A2(new_n2070_), .A3(new_n1954_), .ZN(new_n2071_));
  NAND3_X1   g01815(.A1(new_n2050_), .A2(new_n2068_), .A3(new_n2071_), .ZN(new_n2072_));
  OAI21_X1   g01816(.A1(new_n2048_), .A2(new_n2045_), .B(\a[17] ), .ZN(new_n2073_));
  NAND2_X1   g01817(.A1(new_n2046_), .A2(new_n1344_), .ZN(new_n2074_));
  NAND2_X1   g01818(.A1(new_n2074_), .A2(new_n2073_), .ZN(new_n2075_));
  AOI21_X1   g01819(.A1(new_n2069_), .A2(new_n2070_), .B(new_n1954_), .ZN(new_n2076_));
  NOR3_X1    g01820(.A1(new_n2064_), .A2(new_n2067_), .A3(new_n1945_), .ZN(new_n2077_));
  OAI21_X1   g01821(.A1(new_n2076_), .A2(new_n2077_), .B(new_n2075_), .ZN(new_n2078_));
  NAND2_X1   g01822(.A1(new_n2078_), .A2(new_n2072_), .ZN(new_n2079_));
  XOR2_X1    g01823(.A1(new_n2079_), .A2(new_n2043_), .Z(new_n2080_));
  INV_X1     g01824(.I(new_n2080_), .ZN(new_n2081_));
  OAI22_X1   g01825(.A1(new_n993_), .A2(new_n667_), .B1(new_n577_), .B2(new_n997_), .ZN(new_n2082_));
  AOI21_X1   g01826(.A1(\b[7] ), .A2(new_n1486_), .B(new_n2082_), .ZN(new_n2083_));
  OAI21_X1   g01827(.A1(new_n1240_), .A2(new_n1323_), .B(new_n2083_), .ZN(new_n2084_));
  XOR2_X1    g01828(.A1(new_n2084_), .A2(new_n1002_), .Z(new_n2085_));
  NOR2_X1    g01829(.A1(new_n1909_), .A2(new_n1906_), .ZN(new_n2086_));
  NAND2_X1   g01830(.A1(new_n1962_), .A2(new_n1914_), .ZN(new_n2087_));
  NAND2_X1   g01831(.A1(new_n1956_), .A2(new_n1910_), .ZN(new_n2088_));
  AND3_X2    g01832(.A1(new_n2087_), .A2(new_n2088_), .A3(new_n2086_), .Z(new_n2089_));
  AOI21_X1   g01833(.A1(new_n1902_), .A2(new_n1964_), .B(new_n2089_), .ZN(new_n2090_));
  NOR2_X1    g01834(.A1(new_n2090_), .A2(new_n2085_), .ZN(new_n2091_));
  XOR2_X1    g01835(.A1(new_n2084_), .A2(\a[14] ), .Z(new_n2092_));
  NAND3_X1   g01836(.A1(new_n2087_), .A2(new_n2088_), .A3(new_n2086_), .ZN(new_n2093_));
  OAI21_X1   g01837(.A1(new_n1967_), .A2(new_n1970_), .B(new_n2093_), .ZN(new_n2094_));
  NOR2_X1    g01838(.A1(new_n2094_), .A2(new_n2092_), .ZN(new_n2095_));
  NOR3_X1    g01839(.A1(new_n2091_), .A2(new_n2081_), .A3(new_n2095_), .ZN(new_n2096_));
  NAND2_X1   g01840(.A1(new_n2094_), .A2(new_n2092_), .ZN(new_n2097_));
  NAND2_X1   g01841(.A1(new_n2090_), .A2(new_n2085_), .ZN(new_n2098_));
  AOI21_X1   g01842(.A1(new_n2098_), .A2(new_n2097_), .B(new_n2080_), .ZN(new_n2099_));
  OR2_X2     g01843(.A1(new_n2096_), .A2(new_n2099_), .Z(new_n2100_));
  OAI22_X1   g01844(.A1(new_n713_), .A2(new_n941_), .B1(new_n852_), .B2(new_n717_), .ZN(new_n2101_));
  AOI21_X1   g01845(.A1(\b[10] ), .A2(new_n1126_), .B(new_n2101_), .ZN(new_n2102_));
  OAI21_X1   g01846(.A1(new_n953_), .A2(new_n986_), .B(new_n2102_), .ZN(new_n2103_));
  XOR2_X1    g01847(.A1(new_n2103_), .A2(\a[11] ), .Z(new_n2104_));
  INV_X1     g01848(.I(new_n2104_), .ZN(new_n2105_));
  AOI21_X1   g01849(.A1(new_n1990_), .A2(new_n1972_), .B(new_n2105_), .ZN(new_n2106_));
  NOR3_X1    g01850(.A1(new_n1978_), .A2(new_n1983_), .A3(new_n2104_), .ZN(new_n2107_));
  NOR3_X1    g01851(.A1(new_n2107_), .A2(new_n2106_), .A3(new_n2100_), .ZN(new_n2108_));
  NOR2_X1    g01852(.A1(new_n2096_), .A2(new_n2099_), .ZN(new_n2109_));
  OAI21_X1   g01853(.A1(new_n1978_), .A2(new_n1983_), .B(new_n2104_), .ZN(new_n2110_));
  NAND3_X1   g01854(.A1(new_n1990_), .A2(new_n1972_), .A3(new_n2105_), .ZN(new_n2111_));
  AOI21_X1   g01855(.A1(new_n2110_), .A2(new_n2111_), .B(new_n2109_), .ZN(new_n2112_));
  NOR2_X1    g01856(.A1(new_n2108_), .A2(new_n2112_), .ZN(new_n2113_));
  INV_X1     g01857(.I(new_n1992_), .ZN(new_n2114_));
  AOI22_X1   g01858(.A1(new_n518_), .A2(\b[15] ), .B1(\b[14] ), .B2(new_n636_), .ZN(new_n2115_));
  OAI21_X1   g01859(.A1(new_n1070_), .A2(new_n917_), .B(new_n2115_), .ZN(new_n2116_));
  INV_X1     g01860(.I(new_n2116_), .ZN(new_n2117_));
  OAI21_X1   g01861(.A1(new_n1275_), .A2(new_n624_), .B(new_n2117_), .ZN(new_n2118_));
  XOR2_X1    g01862(.A1(new_n2118_), .A2(\a[8] ), .Z(new_n2119_));
  OAI21_X1   g01863(.A1(new_n1997_), .A2(new_n2114_), .B(new_n2119_), .ZN(new_n2120_));
  INV_X1     g01864(.I(new_n2120_), .ZN(new_n2121_));
  NOR3_X1    g01865(.A1(new_n1997_), .A2(new_n2114_), .A3(new_n2119_), .ZN(new_n2122_));
  NOR2_X1    g01866(.A1(new_n2121_), .A2(new_n2122_), .ZN(new_n2123_));
  NAND2_X1   g01867(.A1(new_n2123_), .A2(new_n2113_), .ZN(new_n2124_));
  OR2_X2     g01868(.A1(new_n2108_), .A2(new_n2112_), .Z(new_n2125_));
  OAI21_X1   g01869(.A1(new_n2121_), .A2(new_n2122_), .B(new_n2125_), .ZN(new_n2126_));
  AOI21_X1   g01870(.A1(new_n2124_), .A2(new_n2126_), .B(new_n2042_), .ZN(new_n2127_));
  NAND3_X1   g01871(.A1(new_n2124_), .A2(new_n2042_), .A3(new_n2126_), .ZN(new_n2128_));
  INV_X1     g01872(.I(new_n2128_), .ZN(new_n2129_));
  AOI21_X1   g01873(.A1(new_n2009_), .A2(new_n2004_), .B(new_n2003_), .ZN(new_n2130_));
  NOR3_X1    g01874(.A1(new_n2130_), .A2(new_n2127_), .A3(new_n2129_), .ZN(new_n2131_));
  INV_X1     g01875(.I(new_n2127_), .ZN(new_n2132_));
  OAI21_X1   g01876(.A1(new_n2013_), .A2(new_n2005_), .B(new_n2011_), .ZN(new_n2133_));
  AOI21_X1   g01877(.A1(new_n2132_), .A2(new_n2128_), .B(new_n2133_), .ZN(new_n2134_));
  NOR2_X1    g01878(.A1(new_n2131_), .A2(new_n2134_), .ZN(new_n2135_));
  XOR2_X1    g01879(.A1(new_n2135_), .A2(new_n2037_), .Z(new_n2136_));
  XOR2_X1    g01880(.A1(new_n2020_), .A2(new_n2136_), .Z(\f[21] ));
  INV_X1     g01881(.I(new_n2037_), .ZN(new_n2138_));
  NOR2_X1    g01882(.A1(new_n2135_), .A2(new_n2138_), .ZN(new_n2139_));
  INV_X1     g01883(.I(new_n2139_), .ZN(new_n2140_));
  OAI21_X1   g01884(.A1(new_n2020_), .A2(new_n2136_), .B(new_n2140_), .ZN(new_n2141_));
  INV_X1     g01885(.I(\b[22] ), .ZN(new_n2142_));
  OAI22_X1   g01886(.A1(new_n277_), .A2(new_n2142_), .B1(new_n2027_), .B2(new_n262_), .ZN(new_n2143_));
  AOI21_X1   g01887(.A1(\b[20] ), .A2(new_n283_), .B(new_n2143_), .ZN(new_n2144_));
  AOI21_X1   g01888(.A1(new_n2028_), .A2(\b[20] ), .B(\b[19] ), .ZN(new_n2145_));
  AOI21_X1   g01889(.A1(new_n1869_), .A2(\b[21] ), .B(\b[20] ), .ZN(new_n2146_));
  NOR2_X1    g01890(.A1(new_n2145_), .A2(new_n2146_), .ZN(new_n2147_));
  XNOR2_X1   g01891(.A1(\b[21] ), .A2(\b[22] ), .ZN(new_n2148_));
  NOR2_X1    g01892(.A1(new_n2147_), .A2(new_n2148_), .ZN(new_n2149_));
  INV_X1     g01893(.I(new_n2147_), .ZN(new_n2150_));
  XOR2_X1    g01894(.A1(\b[21] ), .A2(\b[22] ), .Z(new_n2151_));
  NOR2_X1    g01895(.A1(new_n2150_), .A2(new_n2151_), .ZN(new_n2152_));
  NOR2_X1    g01896(.A1(new_n2152_), .A2(new_n2149_), .ZN(new_n2153_));
  OAI21_X1   g01897(.A1(new_n2153_), .A2(new_n279_), .B(new_n2144_), .ZN(new_n2154_));
  XOR2_X1    g01898(.A1(new_n2154_), .A2(\a[2] ), .Z(new_n2155_));
  OAI21_X1   g01899(.A1(new_n2133_), .A2(new_n2127_), .B(new_n2128_), .ZN(new_n2156_));
  AOI22_X1   g01900(.A1(new_n800_), .A2(\b[18] ), .B1(\b[19] ), .B2(new_n333_), .ZN(new_n2157_));
  OAI21_X1   g01901(.A1(new_n1432_), .A2(new_n392_), .B(new_n2157_), .ZN(new_n2158_));
  INV_X1     g01902(.I(new_n2158_), .ZN(new_n2159_));
  NAND2_X1   g01903(.A1(new_n1695_), .A2(new_n330_), .ZN(new_n2160_));
  AOI21_X1   g01904(.A1(new_n2160_), .A2(new_n2159_), .B(new_n312_), .ZN(new_n2161_));
  AND3_X2    g01905(.A1(new_n2160_), .A2(new_n312_), .A3(new_n2159_), .Z(new_n2162_));
  NOR2_X1    g01906(.A1(new_n2162_), .A2(new_n2161_), .ZN(new_n2163_));
  AOI21_X1   g01907(.A1(new_n2125_), .A2(new_n2120_), .B(new_n2122_), .ZN(new_n2164_));
  INV_X1     g01908(.I(new_n2164_), .ZN(new_n2165_));
  OAI21_X1   g01909(.A1(new_n2109_), .A2(new_n2106_), .B(new_n2111_), .ZN(new_n2166_));
  AOI21_X1   g01910(.A1(new_n2094_), .A2(new_n2092_), .B(new_n2080_), .ZN(new_n2167_));
  NOR2_X1    g01911(.A1(new_n2167_), .A2(new_n2095_), .ZN(new_n2168_));
  INV_X1     g01912(.I(new_n2168_), .ZN(new_n2169_));
  AOI21_X1   g01913(.A1(new_n2068_), .A2(new_n2071_), .B(new_n2075_), .ZN(new_n2170_));
  AOI21_X1   g01914(.A1(new_n2079_), .A2(new_n2043_), .B(new_n2170_), .ZN(new_n2171_));
  NOR2_X1    g01915(.A1(new_n2065_), .A2(new_n2066_), .ZN(new_n2172_));
  NAND2_X1   g01916(.A1(new_n1945_), .A2(new_n2063_), .ZN(new_n2173_));
  NOR2_X1    g01917(.A1(new_n1945_), .A2(new_n2063_), .ZN(new_n2174_));
  AOI21_X1   g01918(.A1(new_n2172_), .A2(new_n2173_), .B(new_n2174_), .ZN(new_n2175_));
  OAI22_X1   g01919(.A1(new_n1751_), .A2(new_n339_), .B1(new_n290_), .B2(new_n1754_), .ZN(new_n2176_));
  NOR2_X1    g01920(.A1(new_n1931_), .A2(new_n276_), .ZN(new_n2177_));
  NOR2_X1    g01921(.A1(new_n2176_), .A2(new_n2177_), .ZN(new_n2178_));
  NAND2_X1   g01922(.A1(new_n1725_), .A2(new_n1746_), .ZN(new_n2179_));
  AOI21_X1   g01923(.A1(new_n2178_), .A2(new_n2179_), .B(new_n1736_), .ZN(new_n2180_));
  AOI22_X1   g01924(.A1(new_n1738_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n1743_), .ZN(new_n2181_));
  NAND2_X1   g01925(.A1(new_n1939_), .A2(\b[2] ), .ZN(new_n2182_));
  NAND2_X1   g01926(.A1(new_n2181_), .A2(new_n2182_), .ZN(new_n2183_));
  NOR2_X1    g01927(.A1(new_n352_), .A2(new_n1757_), .ZN(new_n2184_));
  NOR3_X1    g01928(.A1(new_n2183_), .A2(\a[20] ), .A3(new_n2184_), .ZN(new_n2185_));
  NOR2_X1    g01929(.A1(new_n2185_), .A2(new_n2180_), .ZN(new_n2186_));
  XOR2_X1    g01930(.A1(\a[20] ), .A2(\a[21] ), .Z(new_n2187_));
  XNOR2_X1   g01931(.A1(\a[22] ), .A2(\a[23] ), .ZN(new_n2188_));
  NAND2_X1   g01932(.A1(new_n2188_), .A2(new_n2187_), .ZN(new_n2189_));
  INV_X1     g01933(.I(\a[22] ), .ZN(new_n2190_));
  NOR3_X1    g01934(.A1(new_n2190_), .A2(\a[20] ), .A3(\a[21] ), .ZN(new_n2191_));
  INV_X1     g01935(.I(\a[21] ), .ZN(new_n2192_));
  NOR3_X1    g01936(.A1(new_n1736_), .A2(new_n2192_), .A3(\a[22] ), .ZN(new_n2193_));
  NOR2_X1    g01937(.A1(new_n2193_), .A2(new_n2191_), .ZN(new_n2194_));
  OAI22_X1   g01938(.A1(new_n2189_), .A2(new_n275_), .B1(new_n258_), .B2(new_n2194_), .ZN(new_n2195_));
  XOR2_X1    g01939(.A1(\a[22] ), .A2(\a[23] ), .Z(new_n2196_));
  NAND2_X1   g01940(.A1(new_n2187_), .A2(new_n2196_), .ZN(new_n2197_));
  NOR2_X1    g01941(.A1(new_n2197_), .A2(new_n313_), .ZN(new_n2198_));
  OAI21_X1   g01942(.A1(new_n2195_), .A2(new_n2198_), .B(\a[23] ), .ZN(new_n2199_));
  INV_X1     g01943(.I(\a[23] ), .ZN(new_n2200_));
  XOR2_X1    g01944(.A1(\a[22] ), .A2(\a[23] ), .Z(new_n2201_));
  NOR2_X1    g01945(.A1(new_n2061_), .A2(new_n2201_), .ZN(new_n2202_));
  NAND3_X1   g01946(.A1(new_n1736_), .A2(new_n2192_), .A3(\a[22] ), .ZN(new_n2203_));
  NAND3_X1   g01947(.A1(new_n2190_), .A2(\a[20] ), .A3(\a[21] ), .ZN(new_n2204_));
  NAND2_X1   g01948(.A1(new_n2203_), .A2(new_n2204_), .ZN(new_n2205_));
  AOI22_X1   g01949(.A1(new_n2202_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n2205_), .ZN(new_n2206_));
  XNOR2_X1   g01950(.A1(\a[22] ), .A2(\a[23] ), .ZN(new_n2207_));
  NOR2_X1    g01951(.A1(new_n2061_), .A2(new_n2207_), .ZN(new_n2208_));
  NAND2_X1   g01952(.A1(new_n2208_), .A2(new_n263_), .ZN(new_n2209_));
  NAND3_X1   g01953(.A1(new_n2206_), .A2(new_n2209_), .A3(new_n2200_), .ZN(new_n2210_));
  NAND2_X1   g01954(.A1(new_n2063_), .A2(\a[23] ), .ZN(new_n2211_));
  NAND3_X1   g01955(.A1(new_n2199_), .A2(new_n2210_), .A3(new_n2211_), .ZN(new_n2212_));
  NAND2_X1   g01956(.A1(new_n2206_), .A2(new_n2209_), .ZN(new_n2213_));
  NAND3_X1   g01957(.A1(new_n2213_), .A2(\a[23] ), .A3(new_n2063_), .ZN(new_n2214_));
  NAND2_X1   g01958(.A1(new_n2212_), .A2(new_n2214_), .ZN(new_n2215_));
  NAND2_X1   g01959(.A1(new_n2215_), .A2(new_n2186_), .ZN(new_n2216_));
  OAI21_X1   g01960(.A1(new_n2183_), .A2(new_n2184_), .B(\a[20] ), .ZN(new_n2217_));
  NAND3_X1   g01961(.A1(new_n2178_), .A2(new_n1736_), .A3(new_n2179_), .ZN(new_n2218_));
  NAND2_X1   g01962(.A1(new_n2217_), .A2(new_n2218_), .ZN(new_n2219_));
  NAND3_X1   g01963(.A1(new_n2219_), .A2(new_n2212_), .A3(new_n2214_), .ZN(new_n2220_));
  AOI21_X1   g01964(.A1(new_n2216_), .A2(new_n2220_), .B(new_n2175_), .ZN(new_n2221_));
  NAND2_X1   g01965(.A1(new_n2060_), .A2(new_n2055_), .ZN(new_n2222_));
  NOR2_X1    g01966(.A1(new_n1954_), .A2(new_n2062_), .ZN(new_n2223_));
  NAND2_X1   g01967(.A1(new_n1954_), .A2(new_n2062_), .ZN(new_n2224_));
  OAI21_X1   g01968(.A1(new_n2223_), .A2(new_n2222_), .B(new_n2224_), .ZN(new_n2225_));
  AOI21_X1   g01969(.A1(new_n2212_), .A2(new_n2214_), .B(new_n2219_), .ZN(new_n2226_));
  NOR2_X1    g01970(.A1(new_n2215_), .A2(new_n2186_), .ZN(new_n2227_));
  NOR3_X1    g01971(.A1(new_n2225_), .A2(new_n2226_), .A3(new_n2227_), .ZN(new_n2228_));
  NOR2_X1    g01972(.A1(new_n2221_), .A2(new_n2228_), .ZN(new_n2229_));
  OAI22_X1   g01973(.A1(new_n1592_), .A2(new_n471_), .B1(new_n438_), .B2(new_n1505_), .ZN(new_n2230_));
  AOI21_X1   g01974(.A1(\b[5] ), .A2(new_n1584_), .B(new_n2230_), .ZN(new_n2231_));
  OAI21_X1   g01975(.A1(new_n485_), .A2(new_n1732_), .B(new_n2231_), .ZN(new_n2232_));
  XOR2_X1    g01976(.A1(new_n2232_), .A2(new_n1344_), .Z(new_n2233_));
  NAND2_X1   g01977(.A1(new_n2229_), .A2(new_n2233_), .ZN(new_n2234_));
  OAI21_X1   g01978(.A1(new_n2226_), .A2(new_n2227_), .B(new_n2225_), .ZN(new_n2235_));
  NAND3_X1   g01979(.A1(new_n2175_), .A2(new_n2216_), .A3(new_n2220_), .ZN(new_n2236_));
  NAND2_X1   g01980(.A1(new_n2235_), .A2(new_n2236_), .ZN(new_n2237_));
  XOR2_X1    g01981(.A1(new_n2232_), .A2(\a[17] ), .Z(new_n2238_));
  NAND2_X1   g01982(.A1(new_n2237_), .A2(new_n2238_), .ZN(new_n2239_));
  AOI21_X1   g01983(.A1(new_n2234_), .A2(new_n2239_), .B(new_n2171_), .ZN(new_n2240_));
  AOI21_X1   g01984(.A1(new_n1914_), .A2(new_n1955_), .B(new_n1960_), .ZN(new_n2241_));
  NOR3_X1    g01985(.A1(new_n2075_), .A2(new_n2077_), .A3(new_n2076_), .ZN(new_n2242_));
  AOI21_X1   g01986(.A1(new_n2068_), .A2(new_n2071_), .B(new_n2050_), .ZN(new_n2243_));
  NOR2_X1    g01987(.A1(new_n2243_), .A2(new_n2242_), .ZN(new_n2244_));
  INV_X1     g01988(.I(new_n2170_), .ZN(new_n2245_));
  OAI21_X1   g01989(.A1(new_n2244_), .A2(new_n2241_), .B(new_n2245_), .ZN(new_n2246_));
  NOR2_X1    g01990(.A1(new_n2237_), .A2(new_n2238_), .ZN(new_n2247_));
  NOR2_X1    g01991(.A1(new_n2229_), .A2(new_n2233_), .ZN(new_n2248_));
  NOR3_X1    g01992(.A1(new_n2246_), .A2(new_n2247_), .A3(new_n2248_), .ZN(new_n2249_));
  OAI22_X1   g01993(.A1(new_n993_), .A2(new_n776_), .B1(new_n667_), .B2(new_n997_), .ZN(new_n2250_));
  AOI21_X1   g01994(.A1(\b[8] ), .A2(new_n1486_), .B(new_n2250_), .ZN(new_n2251_));
  OAI21_X1   g01995(.A1(new_n786_), .A2(new_n1323_), .B(new_n2251_), .ZN(new_n2252_));
  XOR2_X1    g01996(.A1(new_n2252_), .A2(\a[14] ), .Z(new_n2253_));
  NOR3_X1    g01997(.A1(new_n2253_), .A2(new_n2249_), .A3(new_n2240_), .ZN(new_n2254_));
  NOR2_X1    g01998(.A1(new_n2240_), .A2(new_n2249_), .ZN(new_n2255_));
  XOR2_X1    g01999(.A1(new_n2252_), .A2(new_n1002_), .Z(new_n2256_));
  NOR2_X1    g02000(.A1(new_n2255_), .A2(new_n2256_), .ZN(new_n2257_));
  NOR2_X1    g02001(.A1(new_n2257_), .A2(new_n2254_), .ZN(new_n2258_));
  NOR2_X1    g02002(.A1(new_n2169_), .A2(new_n2258_), .ZN(new_n2259_));
  INV_X1     g02003(.I(new_n2258_), .ZN(new_n2260_));
  NOR2_X1    g02004(.A1(new_n2260_), .A2(new_n2168_), .ZN(new_n2261_));
  AOI22_X1   g02005(.A1(new_n729_), .A2(\b[13] ), .B1(\b[12] ), .B2(new_n732_), .ZN(new_n2262_));
  OAI21_X1   g02006(.A1(new_n852_), .A2(new_n1127_), .B(new_n2262_), .ZN(new_n2263_));
  INV_X1     g02007(.I(new_n2263_), .ZN(new_n2264_));
  OAI21_X1   g02008(.A1(new_n1082_), .A2(new_n986_), .B(new_n2264_), .ZN(new_n2265_));
  XOR2_X1    g02009(.A1(new_n2265_), .A2(\a[11] ), .Z(new_n2266_));
  NOR3_X1    g02010(.A1(new_n2266_), .A2(new_n2261_), .A3(new_n2259_), .ZN(new_n2267_));
  NAND2_X1   g02011(.A1(new_n2260_), .A2(new_n2168_), .ZN(new_n2268_));
  NAND2_X1   g02012(.A1(new_n2169_), .A2(new_n2258_), .ZN(new_n2269_));
  XOR2_X1    g02013(.A1(new_n2265_), .A2(new_n722_), .Z(new_n2270_));
  AOI21_X1   g02014(.A1(new_n2268_), .A2(new_n2269_), .B(new_n2270_), .ZN(new_n2271_));
  NOR2_X1    g02015(.A1(new_n2271_), .A2(new_n2267_), .ZN(new_n2272_));
  NAND2_X1   g02016(.A1(new_n2272_), .A2(new_n2166_), .ZN(new_n2273_));
  AOI21_X1   g02017(.A1(new_n2100_), .A2(new_n2110_), .B(new_n2107_), .ZN(new_n2274_));
  NAND3_X1   g02018(.A1(new_n2270_), .A2(new_n2268_), .A3(new_n2269_), .ZN(new_n2275_));
  OAI21_X1   g02019(.A1(new_n2259_), .A2(new_n2261_), .B(new_n2266_), .ZN(new_n2276_));
  NAND2_X1   g02020(.A1(new_n2276_), .A2(new_n2275_), .ZN(new_n2277_));
  NAND2_X1   g02021(.A1(new_n2274_), .A2(new_n2277_), .ZN(new_n2278_));
  AOI22_X1   g02022(.A1(new_n518_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n636_), .ZN(new_n2279_));
  OAI21_X1   g02023(.A1(new_n1093_), .A2(new_n917_), .B(new_n2279_), .ZN(new_n2280_));
  AOI21_X1   g02024(.A1(new_n1701_), .A2(new_n618_), .B(new_n2280_), .ZN(new_n2281_));
  XOR2_X1    g02025(.A1(new_n2281_), .A2(new_n488_), .Z(new_n2282_));
  INV_X1     g02026(.I(new_n2282_), .ZN(new_n2283_));
  AOI21_X1   g02027(.A1(new_n2278_), .A2(new_n2273_), .B(new_n2283_), .ZN(new_n2284_));
  NOR2_X1    g02028(.A1(new_n2274_), .A2(new_n2277_), .ZN(new_n2285_));
  NOR2_X1    g02029(.A1(new_n2272_), .A2(new_n2166_), .ZN(new_n2286_));
  NOR3_X1    g02030(.A1(new_n2285_), .A2(new_n2286_), .A3(new_n2282_), .ZN(new_n2287_));
  NOR2_X1    g02031(.A1(new_n2284_), .A2(new_n2287_), .ZN(new_n2288_));
  NAND2_X1   g02032(.A1(new_n2165_), .A2(new_n2288_), .ZN(new_n2289_));
  INV_X1     g02033(.I(new_n2288_), .ZN(new_n2290_));
  NAND2_X1   g02034(.A1(new_n2290_), .A2(new_n2164_), .ZN(new_n2291_));
  NAND3_X1   g02035(.A1(new_n2289_), .A2(new_n2291_), .A3(new_n2163_), .ZN(new_n2292_));
  INV_X1     g02036(.I(new_n2163_), .ZN(new_n2293_));
  NOR2_X1    g02037(.A1(new_n2290_), .A2(new_n2164_), .ZN(new_n2294_));
  NOR2_X1    g02038(.A1(new_n2165_), .A2(new_n2288_), .ZN(new_n2295_));
  OAI21_X1   g02039(.A1(new_n2295_), .A2(new_n2294_), .B(new_n2293_), .ZN(new_n2296_));
  NAND2_X1   g02040(.A1(new_n2296_), .A2(new_n2292_), .ZN(new_n2297_));
  XOR2_X1    g02041(.A1(new_n2156_), .A2(new_n2297_), .Z(new_n2298_));
  NOR2_X1    g02042(.A1(new_n2298_), .A2(new_n2155_), .ZN(new_n2299_));
  NAND2_X1   g02043(.A1(new_n2298_), .A2(new_n2155_), .ZN(new_n2300_));
  INV_X1     g02044(.I(new_n2300_), .ZN(new_n2301_));
  NOR2_X1    g02045(.A1(new_n2301_), .A2(new_n2299_), .ZN(new_n2302_));
  XOR2_X1    g02046(.A1(new_n2141_), .A2(new_n2302_), .Z(\f[22] ));
  AOI21_X1   g02047(.A1(new_n2289_), .A2(new_n2291_), .B(new_n2293_), .ZN(new_n2304_));
  AOI21_X1   g02048(.A1(new_n2156_), .A2(new_n2297_), .B(new_n2304_), .ZN(new_n2305_));
  INV_X1     g02049(.I(new_n2287_), .ZN(new_n2306_));
  AOI22_X1   g02050(.A1(new_n518_), .A2(\b[17] ), .B1(\b[16] ), .B2(new_n636_), .ZN(new_n2307_));
  OAI21_X1   g02051(.A1(new_n1268_), .A2(new_n917_), .B(new_n2307_), .ZN(new_n2308_));
  INV_X1     g02052(.I(new_n2308_), .ZN(new_n2309_));
  NAND3_X1   g02053(.A1(new_n1443_), .A2(new_n618_), .A3(new_n1440_), .ZN(new_n2310_));
  AOI21_X1   g02054(.A1(new_n2310_), .A2(new_n2309_), .B(new_n488_), .ZN(new_n2311_));
  NAND3_X1   g02055(.A1(new_n2310_), .A2(new_n488_), .A3(new_n2309_), .ZN(new_n2312_));
  INV_X1     g02056(.I(new_n2312_), .ZN(new_n2313_));
  NOR2_X1    g02057(.A1(new_n2313_), .A2(new_n2311_), .ZN(new_n2314_));
  AOI22_X1   g02058(.A1(new_n729_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n732_), .ZN(new_n2315_));
  OAI21_X1   g02059(.A1(new_n941_), .A2(new_n1127_), .B(new_n2315_), .ZN(new_n2316_));
  INV_X1     g02060(.I(new_n2316_), .ZN(new_n2317_));
  OAI21_X1   g02061(.A1(new_n1100_), .A2(new_n1102_), .B(new_n724_), .ZN(new_n2318_));
  AOI21_X1   g02062(.A1(new_n2318_), .A2(new_n2317_), .B(new_n722_), .ZN(new_n2319_));
  NAND3_X1   g02063(.A1(new_n2318_), .A2(new_n722_), .A3(new_n2317_), .ZN(new_n2320_));
  INV_X1     g02064(.I(new_n2320_), .ZN(new_n2321_));
  NOR2_X1    g02065(.A1(new_n2321_), .A2(new_n2319_), .ZN(new_n2322_));
  INV_X1     g02066(.I(new_n2254_), .ZN(new_n2323_));
  OAI22_X1   g02067(.A1(new_n2167_), .A2(new_n2095_), .B1(new_n2255_), .B2(new_n2256_), .ZN(new_n2324_));
  NOR2_X1    g02068(.A1(new_n1459_), .A2(new_n1460_), .ZN(new_n2325_));
  AOI22_X1   g02069(.A1(new_n1006_), .A2(\b[11] ), .B1(\b[10] ), .B2(new_n1009_), .ZN(new_n2326_));
  OAI21_X1   g02070(.A1(new_n667_), .A2(new_n1481_), .B(new_n2326_), .ZN(new_n2327_));
  AOI21_X1   g02071(.A1(new_n2325_), .A2(new_n1013_), .B(new_n2327_), .ZN(new_n2328_));
  NOR2_X1    g02072(.A1(new_n2328_), .A2(new_n1002_), .ZN(new_n2329_));
  INV_X1     g02073(.I(new_n2327_), .ZN(new_n2330_));
  OAI21_X1   g02074(.A1(new_n859_), .A2(new_n1323_), .B(new_n2330_), .ZN(new_n2331_));
  NOR2_X1    g02075(.A1(new_n2331_), .A2(\a[14] ), .ZN(new_n2332_));
  OAI21_X1   g02076(.A1(new_n2246_), .A2(new_n2248_), .B(new_n2234_), .ZN(new_n2333_));
  OAI22_X1   g02077(.A1(new_n1592_), .A2(new_n577_), .B1(new_n471_), .B2(new_n1505_), .ZN(new_n2334_));
  NOR2_X1    g02078(.A1(new_n1917_), .A2(new_n438_), .ZN(new_n2335_));
  NOR2_X1    g02079(.A1(new_n2334_), .A2(new_n2335_), .ZN(new_n2336_));
  OAI21_X1   g02080(.A1(new_n587_), .A2(new_n1732_), .B(new_n2336_), .ZN(new_n2337_));
  NAND2_X1   g02081(.A1(new_n2337_), .A2(\a[17] ), .ZN(new_n2338_));
  INV_X1     g02082(.I(new_n2336_), .ZN(new_n2339_));
  AOI21_X1   g02083(.A1(new_n799_), .A2(new_n1354_), .B(new_n2339_), .ZN(new_n2340_));
  NAND2_X1   g02084(.A1(new_n2340_), .A2(new_n1344_), .ZN(new_n2341_));
  OAI21_X1   g02085(.A1(new_n2175_), .A2(new_n2227_), .B(new_n2216_), .ZN(new_n2342_));
  NAND3_X1   g02086(.A1(new_n2341_), .A2(new_n2342_), .A3(new_n2338_), .ZN(new_n2343_));
  NOR2_X1    g02087(.A1(new_n2340_), .A2(new_n1344_), .ZN(new_n2344_));
  NOR2_X1    g02088(.A1(new_n2337_), .A2(\a[17] ), .ZN(new_n2345_));
  AOI21_X1   g02089(.A1(new_n2225_), .A2(new_n2220_), .B(new_n2226_), .ZN(new_n2346_));
  OAI21_X1   g02090(.A1(new_n2344_), .A2(new_n2345_), .B(new_n2346_), .ZN(new_n2347_));
  AOI22_X1   g02091(.A1(new_n1738_), .A2(\b[5] ), .B1(\b[4] ), .B2(new_n1743_), .ZN(new_n2348_));
  NAND2_X1   g02092(.A1(new_n1939_), .A2(\b[3] ), .ZN(new_n2349_));
  NAND2_X1   g02093(.A1(new_n2348_), .A2(new_n2349_), .ZN(new_n2350_));
  AOI21_X1   g02094(.A1(new_n382_), .A2(new_n1746_), .B(new_n2350_), .ZN(new_n2351_));
  NOR2_X1    g02095(.A1(new_n2351_), .A2(new_n1736_), .ZN(new_n2352_));
  INV_X1     g02096(.I(new_n2350_), .ZN(new_n2353_));
  OAI21_X1   g02097(.A1(new_n566_), .A2(new_n1757_), .B(new_n2353_), .ZN(new_n2354_));
  NOR2_X1    g02098(.A1(new_n2354_), .A2(\a[20] ), .ZN(new_n2355_));
  NAND2_X1   g02099(.A1(new_n2208_), .A2(new_n554_), .ZN(new_n2356_));
  NAND2_X1   g02100(.A1(new_n2202_), .A2(\b[2] ), .ZN(new_n2357_));
  NAND2_X1   g02101(.A1(new_n2205_), .A2(\b[1] ), .ZN(new_n2358_));
  AOI21_X1   g02102(.A1(new_n2190_), .A2(\a[23] ), .B(\a[20] ), .ZN(new_n2359_));
  AOI21_X1   g02103(.A1(\a[22] ), .A2(new_n2200_), .B(new_n1736_), .ZN(new_n2360_));
  NOR3_X1    g02104(.A1(new_n2187_), .A2(new_n2359_), .A3(new_n2360_), .ZN(new_n2361_));
  NAND2_X1   g02105(.A1(new_n2361_), .A2(\b[0] ), .ZN(new_n2362_));
  NAND4_X1   g02106(.A1(new_n2356_), .A2(new_n2362_), .A3(new_n2357_), .A4(new_n2358_), .ZN(new_n2363_));
  NAND2_X1   g02107(.A1(new_n2363_), .A2(\a[23] ), .ZN(new_n2364_));
  NOR2_X1    g02108(.A1(new_n2197_), .A2(new_n282_), .ZN(new_n2365_));
  NOR2_X1    g02109(.A1(new_n2189_), .A2(new_n276_), .ZN(new_n2366_));
  NOR2_X1    g02110(.A1(new_n2194_), .A2(new_n275_), .ZN(new_n2367_));
  INV_X1     g02111(.I(new_n2359_), .ZN(new_n2368_));
  OAI21_X1   g02112(.A1(new_n2190_), .A2(\a[23] ), .B(\a[20] ), .ZN(new_n2369_));
  NAND3_X1   g02113(.A1(new_n2368_), .A2(new_n2061_), .A3(new_n2369_), .ZN(new_n2370_));
  NOR2_X1    g02114(.A1(new_n2370_), .A2(new_n258_), .ZN(new_n2371_));
  NOR4_X1    g02115(.A1(new_n2371_), .A2(new_n2365_), .A3(new_n2366_), .A4(new_n2367_), .ZN(new_n2372_));
  NAND2_X1   g02116(.A1(new_n2372_), .A2(new_n2200_), .ZN(new_n2373_));
  NOR3_X1    g02117(.A1(new_n2213_), .A2(new_n2200_), .A3(new_n2062_), .ZN(new_n2374_));
  AOI21_X1   g02118(.A1(new_n2364_), .A2(new_n2373_), .B(new_n2374_), .ZN(new_n2375_));
  NOR4_X1    g02119(.A1(new_n2363_), .A2(new_n2213_), .A3(new_n2200_), .A4(new_n2062_), .ZN(new_n2376_));
  NOR4_X1    g02120(.A1(new_n2355_), .A2(new_n2352_), .A3(new_n2375_), .A4(new_n2376_), .ZN(new_n2377_));
  NAND2_X1   g02121(.A1(new_n2354_), .A2(\a[20] ), .ZN(new_n2378_));
  NAND2_X1   g02122(.A1(new_n2351_), .A2(new_n1736_), .ZN(new_n2379_));
  NAND2_X1   g02123(.A1(new_n2373_), .A2(new_n2364_), .ZN(new_n2380_));
  NOR2_X1    g02124(.A1(new_n2195_), .A2(new_n2198_), .ZN(new_n2381_));
  NAND3_X1   g02125(.A1(new_n2381_), .A2(\a[23] ), .A3(new_n2063_), .ZN(new_n2382_));
  NAND2_X1   g02126(.A1(new_n2380_), .A2(new_n2382_), .ZN(new_n2383_));
  NAND4_X1   g02127(.A1(new_n2372_), .A2(\a[23] ), .A3(new_n2381_), .A4(new_n2063_), .ZN(new_n2384_));
  AOI22_X1   g02128(.A1(new_n2383_), .A2(new_n2384_), .B1(new_n2378_), .B2(new_n2379_), .ZN(new_n2385_));
  NOR2_X1    g02129(.A1(new_n2385_), .A2(new_n2377_), .ZN(new_n2386_));
  NAND3_X1   g02130(.A1(new_n2347_), .A2(new_n2343_), .A3(new_n2386_), .ZN(new_n2387_));
  NOR3_X1    g02131(.A1(new_n2344_), .A2(new_n2346_), .A3(new_n2345_), .ZN(new_n2388_));
  AOI21_X1   g02132(.A1(new_n2338_), .A2(new_n2341_), .B(new_n2342_), .ZN(new_n2389_));
  NAND4_X1   g02133(.A1(new_n2383_), .A2(new_n2378_), .A3(new_n2379_), .A4(new_n2384_), .ZN(new_n2390_));
  OAI22_X1   g02134(.A1(new_n2355_), .A2(new_n2352_), .B1(new_n2375_), .B2(new_n2376_), .ZN(new_n2391_));
  NAND2_X1   g02135(.A1(new_n2390_), .A2(new_n2391_), .ZN(new_n2392_));
  OAI21_X1   g02136(.A1(new_n2389_), .A2(new_n2388_), .B(new_n2392_), .ZN(new_n2393_));
  NAND2_X1   g02137(.A1(new_n2393_), .A2(new_n2387_), .ZN(new_n2394_));
  NOR2_X1    g02138(.A1(new_n2394_), .A2(new_n2333_), .ZN(new_n2395_));
  AOI21_X1   g02139(.A1(new_n2171_), .A2(new_n2239_), .B(new_n2247_), .ZN(new_n2396_));
  NOR3_X1    g02140(.A1(new_n2389_), .A2(new_n2388_), .A3(new_n2392_), .ZN(new_n2397_));
  AOI21_X1   g02141(.A1(new_n2347_), .A2(new_n2343_), .B(new_n2386_), .ZN(new_n2398_));
  NOR2_X1    g02142(.A1(new_n2397_), .A2(new_n2398_), .ZN(new_n2399_));
  NOR2_X1    g02143(.A1(new_n2399_), .A2(new_n2396_), .ZN(new_n2400_));
  NOR4_X1    g02144(.A1(new_n2400_), .A2(new_n2395_), .A3(new_n2329_), .A4(new_n2332_), .ZN(new_n2401_));
  NAND2_X1   g02145(.A1(new_n2331_), .A2(\a[14] ), .ZN(new_n2402_));
  NAND2_X1   g02146(.A1(new_n2328_), .A2(new_n1002_), .ZN(new_n2403_));
  NAND3_X1   g02147(.A1(new_n2396_), .A2(new_n2387_), .A3(new_n2393_), .ZN(new_n2404_));
  NAND2_X1   g02148(.A1(new_n2394_), .A2(new_n2333_), .ZN(new_n2405_));
  AOI22_X1   g02149(.A1(new_n2405_), .A2(new_n2404_), .B1(new_n2402_), .B2(new_n2403_), .ZN(new_n2406_));
  NOR2_X1    g02150(.A1(new_n2401_), .A2(new_n2406_), .ZN(new_n2407_));
  NAND3_X1   g02151(.A1(new_n2407_), .A2(new_n2324_), .A3(new_n2323_), .ZN(new_n2408_));
  OAI21_X1   g02152(.A1(new_n2090_), .A2(new_n2085_), .B(new_n2081_), .ZN(new_n2409_));
  AOI21_X1   g02153(.A1(new_n2409_), .A2(new_n2098_), .B(new_n2257_), .ZN(new_n2410_));
  NAND4_X1   g02154(.A1(new_n2405_), .A2(new_n2404_), .A3(new_n2402_), .A4(new_n2403_), .ZN(new_n2411_));
  OAI22_X1   g02155(.A1(new_n2400_), .A2(new_n2395_), .B1(new_n2329_), .B2(new_n2332_), .ZN(new_n2412_));
  NAND2_X1   g02156(.A1(new_n2412_), .A2(new_n2411_), .ZN(new_n2413_));
  OAI21_X1   g02157(.A1(new_n2254_), .A2(new_n2410_), .B(new_n2413_), .ZN(new_n2414_));
  AOI21_X1   g02158(.A1(new_n2414_), .A2(new_n2408_), .B(new_n2322_), .ZN(new_n2415_));
  INV_X1     g02159(.I(new_n2322_), .ZN(new_n2416_));
  NOR3_X1    g02160(.A1(new_n2413_), .A2(new_n2410_), .A3(new_n2254_), .ZN(new_n2417_));
  AOI21_X1   g02161(.A1(new_n2323_), .A2(new_n2324_), .B(new_n2407_), .ZN(new_n2418_));
  NOR3_X1    g02162(.A1(new_n2418_), .A2(new_n2416_), .A3(new_n2417_), .ZN(new_n2419_));
  NOR2_X1    g02163(.A1(new_n2419_), .A2(new_n2415_), .ZN(new_n2420_));
  OAI21_X1   g02164(.A1(new_n1709_), .A2(new_n1892_), .B(new_n1804_), .ZN(new_n2421_));
  OAI21_X1   g02165(.A1(new_n2421_), .A2(new_n1977_), .B(new_n1972_), .ZN(new_n2422_));
  AOI21_X1   g02166(.A1(new_n2422_), .A2(new_n2104_), .B(new_n2109_), .ZN(new_n2423_));
  NOR3_X1    g02167(.A1(new_n2423_), .A2(new_n2107_), .A3(new_n2267_), .ZN(new_n2424_));
  OAI21_X1   g02168(.A1(new_n2424_), .A2(new_n2271_), .B(new_n2420_), .ZN(new_n2425_));
  OAI21_X1   g02169(.A1(new_n2418_), .A2(new_n2417_), .B(new_n2416_), .ZN(new_n2426_));
  NAND3_X1   g02170(.A1(new_n2414_), .A2(new_n2408_), .A3(new_n2322_), .ZN(new_n2427_));
  NAND2_X1   g02171(.A1(new_n2426_), .A2(new_n2427_), .ZN(new_n2428_));
  AOI21_X1   g02172(.A1(new_n1810_), .A2(new_n1807_), .B(new_n1887_), .ZN(new_n2429_));
  AOI21_X1   g02173(.A1(new_n2429_), .A2(new_n1985_), .B(new_n1983_), .ZN(new_n2430_));
  OAI21_X1   g02174(.A1(new_n2430_), .A2(new_n2105_), .B(new_n2100_), .ZN(new_n2431_));
  NAND3_X1   g02175(.A1(new_n2431_), .A2(new_n2111_), .A3(new_n2275_), .ZN(new_n2432_));
  NAND3_X1   g02176(.A1(new_n2432_), .A2(new_n2428_), .A3(new_n2276_), .ZN(new_n2433_));
  AOI21_X1   g02177(.A1(new_n2425_), .A2(new_n2433_), .B(new_n2314_), .ZN(new_n2434_));
  INV_X1     g02178(.I(new_n2311_), .ZN(new_n2435_));
  NAND2_X1   g02179(.A1(new_n2435_), .A2(new_n2312_), .ZN(new_n2436_));
  AOI21_X1   g02180(.A1(new_n2432_), .A2(new_n2276_), .B(new_n2428_), .ZN(new_n2437_));
  NOR3_X1    g02181(.A1(new_n2424_), .A2(new_n2271_), .A3(new_n2420_), .ZN(new_n2438_));
  NOR3_X1    g02182(.A1(new_n2438_), .A2(new_n2437_), .A3(new_n2436_), .ZN(new_n2439_));
  NOR2_X1    g02183(.A1(new_n2439_), .A2(new_n2434_), .ZN(new_n2440_));
  OAI21_X1   g02184(.A1(new_n1999_), .A2(new_n1993_), .B(new_n1992_), .ZN(new_n2441_));
  AOI21_X1   g02185(.A1(new_n2441_), .A2(new_n2119_), .B(new_n2113_), .ZN(new_n2442_));
  OAI21_X1   g02186(.A1(new_n2285_), .A2(new_n2286_), .B(new_n2282_), .ZN(new_n2443_));
  OAI21_X1   g02187(.A1(new_n2442_), .A2(new_n2122_), .B(new_n2443_), .ZN(new_n2444_));
  NAND3_X1   g02188(.A1(new_n2444_), .A2(new_n2306_), .A3(new_n2440_), .ZN(new_n2445_));
  OAI21_X1   g02189(.A1(new_n2438_), .A2(new_n2437_), .B(new_n2436_), .ZN(new_n2446_));
  NAND3_X1   g02190(.A1(new_n2425_), .A2(new_n2433_), .A3(new_n2314_), .ZN(new_n2447_));
  NAND2_X1   g02191(.A1(new_n2446_), .A2(new_n2447_), .ZN(new_n2448_));
  OAI21_X1   g02192(.A1(new_n2164_), .A2(new_n2284_), .B(new_n2306_), .ZN(new_n2449_));
  NAND2_X1   g02193(.A1(new_n2449_), .A2(new_n2448_), .ZN(new_n2450_));
  NAND2_X1   g02194(.A1(new_n2450_), .A2(new_n2445_), .ZN(new_n2451_));
  INV_X1     g02195(.I(new_n1871_), .ZN(new_n2452_));
  AOI22_X1   g02196(.A1(new_n800_), .A2(\b[19] ), .B1(\b[20] ), .B2(new_n333_), .ZN(new_n2453_));
  OAI21_X1   g02197(.A1(new_n1553_), .A2(new_n392_), .B(new_n2453_), .ZN(new_n2454_));
  AOI21_X1   g02198(.A1(new_n2452_), .A2(new_n330_), .B(new_n2454_), .ZN(new_n2455_));
  XOR2_X1    g02199(.A1(new_n2455_), .A2(new_n312_), .Z(new_n2456_));
  INV_X1     g02200(.I(new_n2456_), .ZN(new_n2457_));
  NAND2_X1   g02201(.A1(new_n2451_), .A2(new_n2457_), .ZN(new_n2458_));
  NOR2_X1    g02202(.A1(new_n2451_), .A2(new_n2457_), .ZN(new_n2459_));
  INV_X1     g02203(.I(new_n2459_), .ZN(new_n2460_));
  NAND2_X1   g02204(.A1(new_n283_), .A2(\b[21] ), .ZN(new_n2461_));
  AOI22_X1   g02205(.A1(new_n267_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n261_), .ZN(new_n2462_));
  INV_X1     g02206(.I(\b[23] ), .ZN(new_n2463_));
  NAND3_X1   g02207(.A1(new_n2150_), .A2(new_n2027_), .A3(\b[22] ), .ZN(new_n2464_));
  NAND3_X1   g02208(.A1(new_n2147_), .A2(\b[21] ), .A3(new_n2142_), .ZN(new_n2465_));
  AOI21_X1   g02209(.A1(new_n2464_), .A2(new_n2465_), .B(new_n2463_), .ZN(new_n2466_));
  NOR3_X1    g02210(.A1(new_n2147_), .A2(\b[21] ), .A3(new_n2142_), .ZN(new_n2467_));
  INV_X1     g02211(.I(new_n2465_), .ZN(new_n2468_));
  NOR3_X1    g02212(.A1(new_n2468_), .A2(\b[23] ), .A3(new_n2467_), .ZN(new_n2469_));
  NOR2_X1    g02213(.A1(new_n2469_), .A2(new_n2466_), .ZN(new_n2470_));
  NAND2_X1   g02214(.A1(new_n2470_), .A2(new_n265_), .ZN(new_n2471_));
  NAND3_X1   g02215(.A1(new_n2471_), .A2(new_n2461_), .A3(new_n2462_), .ZN(new_n2472_));
  XOR2_X1    g02216(.A1(new_n2472_), .A2(\a[2] ), .Z(new_n2473_));
  AOI21_X1   g02217(.A1(new_n2458_), .A2(new_n2460_), .B(new_n2473_), .ZN(new_n2474_));
  NAND2_X1   g02218(.A1(new_n2460_), .A2(new_n2458_), .ZN(new_n2475_));
  INV_X1     g02219(.I(new_n2473_), .ZN(new_n2476_));
  NOR2_X1    g02220(.A1(new_n2476_), .A2(new_n2475_), .ZN(new_n2477_));
  NOR3_X1    g02221(.A1(new_n2477_), .A2(new_n2305_), .A3(new_n2474_), .ZN(new_n2478_));
  NAND2_X1   g02222(.A1(new_n2156_), .A2(new_n2297_), .ZN(new_n2479_));
  INV_X1     g02223(.I(new_n2304_), .ZN(new_n2480_));
  NAND2_X1   g02224(.A1(new_n2479_), .A2(new_n2480_), .ZN(new_n2481_));
  NAND2_X1   g02225(.A1(new_n2476_), .A2(new_n2475_), .ZN(new_n2482_));
  NAND3_X1   g02226(.A1(new_n2473_), .A2(new_n2458_), .A3(new_n2460_), .ZN(new_n2483_));
  AOI21_X1   g02227(.A1(new_n2482_), .A2(new_n2483_), .B(new_n2481_), .ZN(new_n2484_));
  NOR2_X1    g02228(.A1(new_n2478_), .A2(new_n2484_), .ZN(new_n2485_));
  INV_X1     g02229(.I(new_n2485_), .ZN(new_n2486_));
  INV_X1     g02230(.I(new_n2299_), .ZN(new_n2487_));
  AOI21_X1   g02231(.A1(new_n2141_), .A2(new_n2487_), .B(new_n2301_), .ZN(new_n2488_));
  XOR2_X1    g02232(.A1(new_n2488_), .A2(new_n2486_), .Z(\f[23] ));
  NAND2_X1   g02233(.A1(new_n2481_), .A2(new_n2475_), .ZN(new_n2490_));
  NAND3_X1   g02234(.A1(new_n2305_), .A2(new_n2458_), .A3(new_n2460_), .ZN(new_n2491_));
  AOI21_X1   g02235(.A1(new_n2490_), .A2(new_n2491_), .B(new_n2476_), .ZN(new_n2492_));
  INV_X1     g02236(.I(new_n2492_), .ZN(new_n2493_));
  OAI21_X1   g02237(.A1(new_n2488_), .A2(new_n2486_), .B(new_n2493_), .ZN(new_n2494_));
  INV_X1     g02238(.I(\b[24] ), .ZN(new_n2495_));
  OAI22_X1   g02239(.A1(new_n277_), .A2(new_n2495_), .B1(new_n2463_), .B2(new_n262_), .ZN(new_n2496_));
  AOI21_X1   g02240(.A1(\b[22] ), .A2(new_n283_), .B(new_n2496_), .ZN(new_n2497_));
  XOR2_X1    g02241(.A1(\b[23] ), .A2(\b[24] ), .Z(new_n2498_));
  NAND2_X1   g02242(.A1(new_n2147_), .A2(\b[21] ), .ZN(new_n2499_));
  AOI21_X1   g02243(.A1(new_n2499_), .A2(new_n2142_), .B(new_n2463_), .ZN(new_n2500_));
  AOI21_X1   g02244(.A1(new_n2150_), .A2(new_n2027_), .B(new_n2142_), .ZN(new_n2501_));
  NOR2_X1    g02245(.A1(new_n2500_), .A2(new_n2501_), .ZN(new_n2502_));
  NOR2_X1    g02246(.A1(new_n2502_), .A2(new_n2498_), .ZN(new_n2503_));
  NAND2_X1   g02247(.A1(new_n2502_), .A2(new_n2498_), .ZN(new_n2504_));
  INV_X1     g02248(.I(new_n2504_), .ZN(new_n2505_));
  NOR2_X1    g02249(.A1(new_n2505_), .A2(new_n2503_), .ZN(new_n2506_));
  OAI21_X1   g02250(.A1(new_n2506_), .A2(new_n279_), .B(new_n2497_), .ZN(new_n2507_));
  XOR2_X1    g02251(.A1(new_n2507_), .A2(\a[2] ), .Z(new_n2508_));
  INV_X1     g02252(.I(new_n2508_), .ZN(new_n2509_));
  AOI22_X1   g02253(.A1(new_n800_), .A2(\b[20] ), .B1(\b[21] ), .B2(new_n333_), .ZN(new_n2510_));
  OAI21_X1   g02254(.A1(new_n1859_), .A2(new_n392_), .B(new_n2510_), .ZN(new_n2511_));
  AOI21_X1   g02255(.A1(new_n2032_), .A2(new_n330_), .B(new_n2511_), .ZN(new_n2512_));
  XOR2_X1    g02256(.A1(new_n2512_), .A2(new_n312_), .Z(new_n2513_));
  INV_X1     g02257(.I(new_n2513_), .ZN(new_n2514_));
  OAI21_X1   g02258(.A1(new_n2346_), .A2(new_n2385_), .B(new_n2390_), .ZN(new_n2515_));
  OAI22_X1   g02259(.A1(new_n1751_), .A2(new_n438_), .B1(new_n377_), .B2(new_n1754_), .ZN(new_n2516_));
  AOI21_X1   g02260(.A1(\b[4] ), .A2(new_n1939_), .B(new_n2516_), .ZN(new_n2517_));
  NAND2_X1   g02261(.A1(new_n916_), .A2(new_n1746_), .ZN(new_n2518_));
  AOI21_X1   g02262(.A1(new_n2518_), .A2(new_n2517_), .B(new_n1736_), .ZN(new_n2519_));
  OAI21_X1   g02263(.A1(new_n450_), .A2(new_n1757_), .B(new_n2517_), .ZN(new_n2520_));
  NOR2_X1    g02264(.A1(new_n2520_), .A2(\a[20] ), .ZN(new_n2521_));
  NOR2_X1    g02265(.A1(new_n2521_), .A2(new_n2519_), .ZN(new_n2522_));
  NAND2_X1   g02266(.A1(new_n2361_), .A2(\b[1] ), .ZN(new_n2523_));
  AOI22_X1   g02267(.A1(new_n2202_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n2205_), .ZN(new_n2524_));
  NAND2_X1   g02268(.A1(new_n299_), .A2(new_n2208_), .ZN(new_n2525_));
  NAND3_X1   g02269(.A1(new_n2525_), .A2(new_n2524_), .A3(new_n2523_), .ZN(new_n2526_));
  NAND2_X1   g02270(.A1(new_n2526_), .A2(\a[23] ), .ZN(new_n2527_));
  NOR2_X1    g02271(.A1(new_n2370_), .A2(new_n275_), .ZN(new_n2528_));
  OAI22_X1   g02272(.A1(new_n2189_), .A2(new_n290_), .B1(new_n276_), .B2(new_n2194_), .ZN(new_n2529_));
  NOR2_X1    g02273(.A1(new_n429_), .A2(new_n2197_), .ZN(new_n2530_));
  NOR3_X1    g02274(.A1(new_n2530_), .A2(new_n2529_), .A3(new_n2528_), .ZN(new_n2531_));
  NAND2_X1   g02275(.A1(new_n2531_), .A2(new_n2200_), .ZN(new_n2532_));
  XNOR2_X1   g02276(.A1(\a[23] ), .A2(\a[24] ), .ZN(new_n2533_));
  NOR2_X1    g02277(.A1(new_n2533_), .A2(new_n258_), .ZN(new_n2534_));
  INV_X1     g02278(.I(new_n2534_), .ZN(new_n2535_));
  AOI21_X1   g02279(.A1(new_n2532_), .A2(new_n2527_), .B(new_n2535_), .ZN(new_n2536_));
  NOR2_X1    g02280(.A1(new_n2531_), .A2(new_n2200_), .ZN(new_n2537_));
  NOR2_X1    g02281(.A1(new_n2526_), .A2(\a[23] ), .ZN(new_n2538_));
  NOR3_X1    g02282(.A1(new_n2537_), .A2(new_n2538_), .A3(new_n2534_), .ZN(new_n2539_));
  OAI21_X1   g02283(.A1(new_n2536_), .A2(new_n2539_), .B(new_n2384_), .ZN(new_n2540_));
  OAI21_X1   g02284(.A1(new_n2537_), .A2(new_n2538_), .B(new_n2534_), .ZN(new_n2541_));
  NAND3_X1   g02285(.A1(new_n2532_), .A2(new_n2527_), .A3(new_n2535_), .ZN(new_n2542_));
  NAND3_X1   g02286(.A1(new_n2541_), .A2(new_n2542_), .A3(new_n2376_), .ZN(new_n2543_));
  NAND3_X1   g02287(.A1(new_n2522_), .A2(new_n2540_), .A3(new_n2543_), .ZN(new_n2544_));
  XOR2_X1    g02288(.A1(new_n2520_), .A2(new_n1736_), .Z(new_n2545_));
  AOI21_X1   g02289(.A1(new_n2541_), .A2(new_n2542_), .B(new_n2376_), .ZN(new_n2546_));
  NOR3_X1    g02290(.A1(new_n2536_), .A2(new_n2539_), .A3(new_n2384_), .ZN(new_n2547_));
  OAI21_X1   g02291(.A1(new_n2546_), .A2(new_n2547_), .B(new_n2545_), .ZN(new_n2548_));
  NAND2_X1   g02292(.A1(new_n2548_), .A2(new_n2544_), .ZN(new_n2549_));
  NAND2_X1   g02293(.A1(new_n2549_), .A2(new_n2515_), .ZN(new_n2550_));
  AOI21_X1   g02294(.A1(new_n2342_), .A2(new_n2391_), .B(new_n2377_), .ZN(new_n2551_));
  NOR3_X1    g02295(.A1(new_n2545_), .A2(new_n2546_), .A3(new_n2547_), .ZN(new_n2552_));
  AOI21_X1   g02296(.A1(new_n2540_), .A2(new_n2543_), .B(new_n2522_), .ZN(new_n2553_));
  NOR2_X1    g02297(.A1(new_n2552_), .A2(new_n2553_), .ZN(new_n2554_));
  NAND2_X1   g02298(.A1(new_n2554_), .A2(new_n2551_), .ZN(new_n2555_));
  NAND2_X1   g02299(.A1(new_n2550_), .A2(new_n2555_), .ZN(new_n2556_));
  OAI22_X1   g02300(.A1(new_n1592_), .A2(new_n667_), .B1(new_n577_), .B2(new_n1505_), .ZN(new_n2557_));
  AOI21_X1   g02301(.A1(\b[7] ), .A2(new_n1584_), .B(new_n2557_), .ZN(new_n2558_));
  OAI21_X1   g02302(.A1(new_n1240_), .A2(new_n1732_), .B(new_n2558_), .ZN(new_n2559_));
  XOR2_X1    g02303(.A1(new_n2559_), .A2(\a[17] ), .Z(new_n2560_));
  INV_X1     g02304(.I(new_n2560_), .ZN(new_n2561_));
  NAND2_X1   g02305(.A1(new_n2341_), .A2(new_n2338_), .ZN(new_n2562_));
  NOR2_X1    g02306(.A1(new_n2392_), .A2(new_n2346_), .ZN(new_n2563_));
  NOR2_X1    g02307(.A1(new_n2386_), .A2(new_n2342_), .ZN(new_n2564_));
  NOR3_X1    g02308(.A1(new_n2564_), .A2(new_n2563_), .A3(new_n2562_), .ZN(new_n2565_));
  AOI21_X1   g02309(.A1(new_n2399_), .A2(new_n2396_), .B(new_n2565_), .ZN(new_n2566_));
  NOR2_X1    g02310(.A1(new_n2566_), .A2(new_n2561_), .ZN(new_n2567_));
  INV_X1     g02311(.I(new_n2565_), .ZN(new_n2568_));
  OAI21_X1   g02312(.A1(new_n2394_), .A2(new_n2333_), .B(new_n2568_), .ZN(new_n2569_));
  NOR2_X1    g02313(.A1(new_n2569_), .A2(new_n2560_), .ZN(new_n2570_));
  NOR3_X1    g02314(.A1(new_n2567_), .A2(new_n2570_), .A3(new_n2556_), .ZN(new_n2571_));
  INV_X1     g02315(.I(new_n2556_), .ZN(new_n2572_));
  NAND2_X1   g02316(.A1(new_n2569_), .A2(new_n2560_), .ZN(new_n2573_));
  NAND2_X1   g02317(.A1(new_n2566_), .A2(new_n2561_), .ZN(new_n2574_));
  AOI21_X1   g02318(.A1(new_n2574_), .A2(new_n2573_), .B(new_n2572_), .ZN(new_n2575_));
  NOR2_X1    g02319(.A1(new_n2575_), .A2(new_n2571_), .ZN(new_n2576_));
  INV_X1     g02320(.I(new_n2576_), .ZN(new_n2577_));
  OAI22_X1   g02321(.A1(new_n993_), .A2(new_n941_), .B1(new_n852_), .B2(new_n997_), .ZN(new_n2578_));
  AOI21_X1   g02322(.A1(\b[10] ), .A2(new_n1486_), .B(new_n2578_), .ZN(new_n2579_));
  OAI21_X1   g02323(.A1(new_n953_), .A2(new_n1323_), .B(new_n2579_), .ZN(new_n2580_));
  XOR2_X1    g02324(.A1(new_n2580_), .A2(\a[14] ), .Z(new_n2581_));
  INV_X1     g02325(.I(new_n2581_), .ZN(new_n2582_));
  AOI21_X1   g02326(.A1(new_n2408_), .A2(new_n2411_), .B(new_n2582_), .ZN(new_n2583_));
  NOR3_X1    g02327(.A1(new_n2417_), .A2(new_n2401_), .A3(new_n2581_), .ZN(new_n2584_));
  NOR3_X1    g02328(.A1(new_n2584_), .A2(new_n2583_), .A3(new_n2577_), .ZN(new_n2585_));
  OAI21_X1   g02329(.A1(new_n2417_), .A2(new_n2401_), .B(new_n2581_), .ZN(new_n2586_));
  NAND3_X1   g02330(.A1(new_n2408_), .A2(new_n2411_), .A3(new_n2582_), .ZN(new_n2587_));
  AOI21_X1   g02331(.A1(new_n2586_), .A2(new_n2587_), .B(new_n2576_), .ZN(new_n2588_));
  NOR2_X1    g02332(.A1(new_n2585_), .A2(new_n2588_), .ZN(new_n2589_));
  INV_X1     g02333(.I(new_n2589_), .ZN(new_n2590_));
  OAI22_X1   g02334(.A1(new_n713_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n717_), .ZN(new_n2591_));
  AOI21_X1   g02335(.A1(\b[13] ), .A2(new_n1126_), .B(new_n2591_), .ZN(new_n2592_));
  OAI21_X1   g02336(.A1(new_n1275_), .A2(new_n986_), .B(new_n2592_), .ZN(new_n2593_));
  XOR2_X1    g02337(.A1(new_n2593_), .A2(\a[11] ), .Z(new_n2594_));
  INV_X1     g02338(.I(new_n2594_), .ZN(new_n2595_));
  AOI21_X1   g02339(.A1(new_n2425_), .A2(new_n2427_), .B(new_n2595_), .ZN(new_n2596_));
  NOR3_X1    g02340(.A1(new_n2437_), .A2(new_n2419_), .A3(new_n2594_), .ZN(new_n2597_));
  NOR3_X1    g02341(.A1(new_n2596_), .A2(new_n2597_), .A3(new_n2590_), .ZN(new_n2598_));
  OAI21_X1   g02342(.A1(new_n2437_), .A2(new_n2419_), .B(new_n2594_), .ZN(new_n2599_));
  NAND3_X1   g02343(.A1(new_n2425_), .A2(new_n2427_), .A3(new_n2595_), .ZN(new_n2600_));
  AOI21_X1   g02344(.A1(new_n2600_), .A2(new_n2599_), .B(new_n2589_), .ZN(new_n2601_));
  NOR2_X1    g02345(.A1(new_n2598_), .A2(new_n2601_), .ZN(new_n2602_));
  INV_X1     g02346(.I(new_n2602_), .ZN(new_n2603_));
  AOI22_X1   g02347(.A1(new_n518_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n636_), .ZN(new_n2604_));
  OAI21_X1   g02348(.A1(new_n1296_), .A2(new_n917_), .B(new_n2604_), .ZN(new_n2605_));
  AOI21_X1   g02349(.A1(new_n2038_), .A2(new_n618_), .B(new_n2605_), .ZN(new_n2606_));
  XOR2_X1    g02350(.A1(new_n2606_), .A2(new_n488_), .Z(new_n2607_));
  INV_X1     g02351(.I(new_n2607_), .ZN(new_n2608_));
  AOI21_X1   g02352(.A1(new_n2445_), .A2(new_n2447_), .B(new_n2608_), .ZN(new_n2609_));
  INV_X1     g02353(.I(new_n2119_), .ZN(new_n2610_));
  OAI21_X1   g02354(.A1(new_n1708_), .A2(new_n1823_), .B(new_n1831_), .ZN(new_n2611_));
  AOI21_X1   g02355(.A1(new_n2611_), .A2(new_n1987_), .B(new_n2114_), .ZN(new_n2612_));
  NAND2_X1   g02356(.A1(new_n2612_), .A2(new_n2610_), .ZN(new_n2613_));
  OAI21_X1   g02357(.A1(new_n2612_), .A2(new_n2610_), .B(new_n2125_), .ZN(new_n2614_));
  AOI21_X1   g02358(.A1(new_n2614_), .A2(new_n2613_), .B(new_n2284_), .ZN(new_n2615_));
  NOR3_X1    g02359(.A1(new_n2615_), .A2(new_n2287_), .A3(new_n2448_), .ZN(new_n2616_));
  NOR3_X1    g02360(.A1(new_n2616_), .A2(new_n2439_), .A3(new_n2607_), .ZN(new_n2617_));
  NOR3_X1    g02361(.A1(new_n2609_), .A2(new_n2617_), .A3(new_n2603_), .ZN(new_n2618_));
  OAI21_X1   g02362(.A1(new_n2616_), .A2(new_n2439_), .B(new_n2607_), .ZN(new_n2619_));
  NAND3_X1   g02363(.A1(new_n2445_), .A2(new_n2447_), .A3(new_n2608_), .ZN(new_n2620_));
  AOI21_X1   g02364(.A1(new_n2620_), .A2(new_n2619_), .B(new_n2602_), .ZN(new_n2621_));
  OAI21_X1   g02365(.A1(new_n2621_), .A2(new_n2618_), .B(new_n2514_), .ZN(new_n2622_));
  INV_X1     g02366(.I(new_n2622_), .ZN(new_n2623_));
  NOR3_X1    g02367(.A1(new_n2514_), .A2(new_n2621_), .A3(new_n2618_), .ZN(new_n2624_));
  INV_X1     g02368(.I(new_n2458_), .ZN(new_n2625_));
  AOI21_X1   g02369(.A1(new_n2305_), .A2(new_n2460_), .B(new_n2625_), .ZN(new_n2626_));
  OAI21_X1   g02370(.A1(new_n2623_), .A2(new_n2624_), .B(new_n2626_), .ZN(new_n2627_));
  INV_X1     g02371(.I(new_n2627_), .ZN(new_n2628_));
  NOR3_X1    g02372(.A1(new_n2626_), .A2(new_n2623_), .A3(new_n2624_), .ZN(new_n2629_));
  NOR3_X1    g02373(.A1(new_n2628_), .A2(new_n2509_), .A3(new_n2629_), .ZN(new_n2630_));
  INV_X1     g02374(.I(new_n2629_), .ZN(new_n2631_));
  AOI21_X1   g02375(.A1(new_n2631_), .A2(new_n2627_), .B(new_n2508_), .ZN(new_n2632_));
  NOR2_X1    g02376(.A1(new_n2630_), .A2(new_n2632_), .ZN(new_n2633_));
  INV_X1     g02377(.I(new_n2633_), .ZN(new_n2634_));
  XOR2_X1    g02378(.A1(new_n2494_), .A2(new_n2634_), .Z(\f[24] ));
  AOI21_X1   g02379(.A1(new_n1855_), .A2(new_n1845_), .B(new_n1844_), .ZN(new_n2636_));
  INV_X1     g02380(.I(new_n2015_), .ZN(new_n2637_));
  OAI21_X1   g02381(.A1(new_n2636_), .A2(new_n2017_), .B(new_n2637_), .ZN(new_n2638_));
  XOR2_X1    g02382(.A1(new_n2135_), .A2(new_n2138_), .Z(new_n2639_));
  AOI21_X1   g02383(.A1(new_n2638_), .A2(new_n2639_), .B(new_n2139_), .ZN(new_n2640_));
  OAI21_X1   g02384(.A1(new_n2640_), .A2(new_n2299_), .B(new_n2300_), .ZN(new_n2641_));
  AOI21_X1   g02385(.A1(new_n2641_), .A2(new_n2485_), .B(new_n2492_), .ZN(new_n2642_));
  AOI21_X1   g02386(.A1(new_n2631_), .A2(new_n2627_), .B(new_n2509_), .ZN(new_n2643_));
  INV_X1     g02387(.I(new_n2643_), .ZN(new_n2644_));
  OAI21_X1   g02388(.A1(new_n2642_), .A2(new_n2633_), .B(new_n2644_), .ZN(new_n2645_));
  INV_X1     g02389(.I(\b[25] ), .ZN(new_n2646_));
  OAI22_X1   g02390(.A1(new_n277_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n262_), .ZN(new_n2647_));
  AOI21_X1   g02391(.A1(\b[23] ), .A2(new_n283_), .B(new_n2647_), .ZN(new_n2648_));
  OAI21_X1   g02392(.A1(new_n2502_), .A2(new_n2495_), .B(\b[23] ), .ZN(new_n2649_));
  NAND2_X1   g02393(.A1(new_n2502_), .A2(new_n2495_), .ZN(new_n2650_));
  NAND2_X1   g02394(.A1(new_n2649_), .A2(new_n2650_), .ZN(new_n2651_));
  NOR3_X1    g02395(.A1(new_n2500_), .A2(new_n2501_), .A3(\b[25] ), .ZN(new_n2652_));
  NOR2_X1    g02396(.A1(new_n2502_), .A2(new_n2646_), .ZN(new_n2653_));
  NOR2_X1    g02397(.A1(new_n2653_), .A2(new_n2652_), .ZN(new_n2654_));
  XOR2_X1    g02398(.A1(new_n2651_), .A2(new_n2654_), .Z(new_n2655_));
  OAI21_X1   g02399(.A1(new_n2655_), .A2(new_n279_), .B(new_n2648_), .ZN(new_n2656_));
  XOR2_X1    g02400(.A1(new_n2656_), .A2(\a[2] ), .Z(new_n2657_));
  AOI21_X1   g02401(.A1(new_n2626_), .A2(new_n2622_), .B(new_n2624_), .ZN(new_n2658_));
  INV_X1     g02402(.I(new_n2153_), .ZN(new_n2659_));
  AOI22_X1   g02403(.A1(new_n800_), .A2(\b[21] ), .B1(\b[22] ), .B2(new_n333_), .ZN(new_n2660_));
  OAI21_X1   g02404(.A1(new_n1860_), .A2(new_n392_), .B(new_n2660_), .ZN(new_n2661_));
  AOI21_X1   g02405(.A1(new_n2659_), .A2(new_n330_), .B(new_n2661_), .ZN(new_n2662_));
  XOR2_X1    g02406(.A1(new_n2662_), .A2(new_n312_), .Z(new_n2663_));
  INV_X1     g02407(.I(new_n2663_), .ZN(new_n2664_));
  AOI21_X1   g02408(.A1(new_n2603_), .A2(new_n2619_), .B(new_n2617_), .ZN(new_n2665_));
  AOI22_X1   g02409(.A1(new_n518_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n636_), .ZN(new_n2666_));
  OAI21_X1   g02410(.A1(new_n1432_), .A2(new_n917_), .B(new_n2666_), .ZN(new_n2667_));
  INV_X1     g02411(.I(new_n2667_), .ZN(new_n2668_));
  NAND2_X1   g02412(.A1(new_n1695_), .A2(new_n618_), .ZN(new_n2669_));
  AOI21_X1   g02413(.A1(new_n2669_), .A2(new_n2668_), .B(new_n488_), .ZN(new_n2670_));
  NAND3_X1   g02414(.A1(new_n2669_), .A2(new_n488_), .A3(new_n2668_), .ZN(new_n2671_));
  INV_X1     g02415(.I(new_n2671_), .ZN(new_n2672_));
  NOR2_X1    g02416(.A1(new_n2672_), .A2(new_n2670_), .ZN(new_n2673_));
  OAI21_X1   g02417(.A1(new_n2166_), .A2(new_n2267_), .B(new_n2276_), .ZN(new_n2674_));
  AOI21_X1   g02418(.A1(new_n2674_), .A2(new_n2420_), .B(new_n2419_), .ZN(new_n2675_));
  OAI21_X1   g02419(.A1(new_n2675_), .A2(new_n2595_), .B(new_n2590_), .ZN(new_n2676_));
  OAI22_X1   g02420(.A1(new_n713_), .A2(new_n1296_), .B1(new_n1268_), .B2(new_n717_), .ZN(new_n2677_));
  AOI21_X1   g02421(.A1(\b[14] ), .A2(new_n1126_), .B(new_n2677_), .ZN(new_n2678_));
  OAI21_X1   g02422(.A1(new_n1306_), .A2(new_n986_), .B(new_n2678_), .ZN(new_n2679_));
  XOR2_X1    g02423(.A1(new_n2679_), .A2(\a[11] ), .Z(new_n2680_));
  NAND2_X1   g02424(.A1(new_n2324_), .A2(new_n2323_), .ZN(new_n2681_));
  OAI21_X1   g02425(.A1(new_n2681_), .A2(new_n2413_), .B(new_n2411_), .ZN(new_n2682_));
  AOI21_X1   g02426(.A1(new_n2682_), .A2(new_n2581_), .B(new_n2576_), .ZN(new_n2683_));
  AOI21_X1   g02427(.A1(new_n2569_), .A2(new_n2560_), .B(new_n2572_), .ZN(new_n2684_));
  OAI21_X1   g02428(.A1(new_n2546_), .A2(new_n2547_), .B(new_n2522_), .ZN(new_n2685_));
  INV_X1     g02429(.I(new_n2685_), .ZN(new_n2686_));
  AOI21_X1   g02430(.A1(new_n2549_), .A2(new_n2515_), .B(new_n2686_), .ZN(new_n2687_));
  NOR2_X1    g02431(.A1(new_n2537_), .A2(new_n2538_), .ZN(new_n2688_));
  NAND2_X1   g02432(.A1(new_n2384_), .A2(new_n2535_), .ZN(new_n2689_));
  NOR2_X1    g02433(.A1(new_n2384_), .A2(new_n2535_), .ZN(new_n2690_));
  AOI21_X1   g02434(.A1(new_n2688_), .A2(new_n2689_), .B(new_n2690_), .ZN(new_n2691_));
  AOI22_X1   g02435(.A1(new_n2202_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n2205_), .ZN(new_n2692_));
  NAND2_X1   g02436(.A1(new_n2361_), .A2(\b[2] ), .ZN(new_n2693_));
  NAND2_X1   g02437(.A1(new_n2692_), .A2(new_n2693_), .ZN(new_n2694_));
  NOR2_X1    g02438(.A1(new_n352_), .A2(new_n2197_), .ZN(new_n2695_));
  OAI21_X1   g02439(.A1(new_n2694_), .A2(new_n2695_), .B(\a[23] ), .ZN(new_n2696_));
  NAND2_X1   g02440(.A1(new_n1725_), .A2(new_n2208_), .ZN(new_n2697_));
  NAND4_X1   g02441(.A1(new_n2697_), .A2(new_n2200_), .A3(new_n2692_), .A4(new_n2693_), .ZN(new_n2698_));
  NAND2_X1   g02442(.A1(new_n2696_), .A2(new_n2698_), .ZN(new_n2699_));
  INV_X1     g02443(.I(new_n2699_), .ZN(new_n2700_));
  XOR2_X1    g02444(.A1(\a[23] ), .A2(\a[24] ), .Z(new_n2701_));
  XNOR2_X1   g02445(.A1(\a[25] ), .A2(\a[26] ), .ZN(new_n2702_));
  NAND2_X1   g02446(.A1(new_n2702_), .A2(new_n2701_), .ZN(new_n2703_));
  INV_X1     g02447(.I(\a[25] ), .ZN(new_n2704_));
  NOR3_X1    g02448(.A1(new_n2704_), .A2(\a[23] ), .A3(\a[24] ), .ZN(new_n2705_));
  INV_X1     g02449(.I(\a[24] ), .ZN(new_n2706_));
  NOR3_X1    g02450(.A1(new_n2200_), .A2(new_n2706_), .A3(\a[25] ), .ZN(new_n2707_));
  NOR2_X1    g02451(.A1(new_n2707_), .A2(new_n2705_), .ZN(new_n2708_));
  OAI22_X1   g02452(.A1(new_n2703_), .A2(new_n275_), .B1(new_n258_), .B2(new_n2708_), .ZN(new_n2709_));
  XOR2_X1    g02453(.A1(\a[25] ), .A2(\a[26] ), .Z(new_n2710_));
  NAND2_X1   g02454(.A1(new_n2701_), .A2(new_n2710_), .ZN(new_n2711_));
  NOR2_X1    g02455(.A1(new_n2711_), .A2(new_n313_), .ZN(new_n2712_));
  OAI21_X1   g02456(.A1(new_n2709_), .A2(new_n2712_), .B(\a[26] ), .ZN(new_n2713_));
  INV_X1     g02457(.I(\a[26] ), .ZN(new_n2714_));
  XOR2_X1    g02458(.A1(\a[25] ), .A2(\a[26] ), .Z(new_n2715_));
  NOR2_X1    g02459(.A1(new_n2533_), .A2(new_n2715_), .ZN(new_n2716_));
  NAND3_X1   g02460(.A1(new_n2200_), .A2(new_n2706_), .A3(\a[25] ), .ZN(new_n2717_));
  NAND3_X1   g02461(.A1(new_n2704_), .A2(\a[23] ), .A3(\a[24] ), .ZN(new_n2718_));
  NAND2_X1   g02462(.A1(new_n2717_), .A2(new_n2718_), .ZN(new_n2719_));
  AOI22_X1   g02463(.A1(new_n2716_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n2719_), .ZN(new_n2720_));
  XNOR2_X1   g02464(.A1(\a[25] ), .A2(\a[26] ), .ZN(new_n2721_));
  NOR2_X1    g02465(.A1(new_n2533_), .A2(new_n2721_), .ZN(new_n2722_));
  NAND2_X1   g02466(.A1(new_n2722_), .A2(new_n263_), .ZN(new_n2723_));
  NAND3_X1   g02467(.A1(new_n2720_), .A2(new_n2723_), .A3(new_n2714_), .ZN(new_n2724_));
  NAND2_X1   g02468(.A1(new_n2535_), .A2(\a[26] ), .ZN(new_n2725_));
  NAND3_X1   g02469(.A1(new_n2713_), .A2(new_n2724_), .A3(new_n2725_), .ZN(new_n2726_));
  NAND2_X1   g02470(.A1(new_n2720_), .A2(new_n2723_), .ZN(new_n2727_));
  NAND3_X1   g02471(.A1(new_n2727_), .A2(\a[26] ), .A3(new_n2535_), .ZN(new_n2728_));
  NAND2_X1   g02472(.A1(new_n2726_), .A2(new_n2728_), .ZN(new_n2729_));
  NAND2_X1   g02473(.A1(new_n2700_), .A2(new_n2729_), .ZN(new_n2730_));
  NAND3_X1   g02474(.A1(new_n2699_), .A2(new_n2726_), .A3(new_n2728_), .ZN(new_n2731_));
  AOI21_X1   g02475(.A1(new_n2730_), .A2(new_n2731_), .B(new_n2691_), .ZN(new_n2732_));
  NAND2_X1   g02476(.A1(new_n2532_), .A2(new_n2527_), .ZN(new_n2733_));
  NOR2_X1    g02477(.A1(new_n2376_), .A2(new_n2534_), .ZN(new_n2734_));
  NAND2_X1   g02478(.A1(new_n2376_), .A2(new_n2534_), .ZN(new_n2735_));
  OAI21_X1   g02479(.A1(new_n2733_), .A2(new_n2734_), .B(new_n2735_), .ZN(new_n2736_));
  AOI21_X1   g02480(.A1(new_n2726_), .A2(new_n2728_), .B(new_n2699_), .ZN(new_n2737_));
  NOR2_X1    g02481(.A1(new_n2700_), .A2(new_n2729_), .ZN(new_n2738_));
  NOR3_X1    g02482(.A1(new_n2736_), .A2(new_n2738_), .A3(new_n2737_), .ZN(new_n2739_));
  NOR2_X1    g02483(.A1(new_n2732_), .A2(new_n2739_), .ZN(new_n2740_));
  OAI22_X1   g02484(.A1(new_n1751_), .A2(new_n471_), .B1(new_n438_), .B2(new_n1754_), .ZN(new_n2741_));
  AOI21_X1   g02485(.A1(\b[5] ), .A2(new_n1939_), .B(new_n2741_), .ZN(new_n2742_));
  OAI21_X1   g02486(.A1(new_n485_), .A2(new_n1757_), .B(new_n2742_), .ZN(new_n2743_));
  XOR2_X1    g02487(.A1(new_n2743_), .A2(new_n1736_), .Z(new_n2744_));
  NAND2_X1   g02488(.A1(new_n2740_), .A2(new_n2744_), .ZN(new_n2745_));
  OAI21_X1   g02489(.A1(new_n2737_), .A2(new_n2738_), .B(new_n2736_), .ZN(new_n2746_));
  NAND3_X1   g02490(.A1(new_n2691_), .A2(new_n2730_), .A3(new_n2731_), .ZN(new_n2747_));
  NAND2_X1   g02491(.A1(new_n2746_), .A2(new_n2747_), .ZN(new_n2748_));
  XOR2_X1    g02492(.A1(new_n2743_), .A2(\a[20] ), .Z(new_n2749_));
  NAND2_X1   g02493(.A1(new_n2748_), .A2(new_n2749_), .ZN(new_n2750_));
  AOI21_X1   g02494(.A1(new_n2745_), .A2(new_n2750_), .B(new_n2687_), .ZN(new_n2751_));
  OAI21_X1   g02495(.A1(new_n2554_), .A2(new_n2551_), .B(new_n2685_), .ZN(new_n2752_));
  NOR2_X1    g02496(.A1(new_n2748_), .A2(new_n2749_), .ZN(new_n2753_));
  NOR2_X1    g02497(.A1(new_n2740_), .A2(new_n2744_), .ZN(new_n2754_));
  NOR3_X1    g02498(.A1(new_n2752_), .A2(new_n2754_), .A3(new_n2753_), .ZN(new_n2755_));
  AOI22_X1   g02499(.A1(new_n1586_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n1495_), .ZN(new_n2756_));
  OAI21_X1   g02500(.A1(new_n577_), .A2(new_n1917_), .B(new_n2756_), .ZN(new_n2757_));
  INV_X1     g02501(.I(new_n2757_), .ZN(new_n2758_));
  NAND2_X1   g02502(.A1(new_n1059_), .A2(new_n1354_), .ZN(new_n2759_));
  AOI21_X1   g02503(.A1(new_n2759_), .A2(new_n2758_), .B(new_n1344_), .ZN(new_n2760_));
  NOR2_X1    g02504(.A1(new_n786_), .A2(new_n1732_), .ZN(new_n2761_));
  NOR3_X1    g02505(.A1(new_n2761_), .A2(\a[17] ), .A3(new_n2757_), .ZN(new_n2762_));
  NOR2_X1    g02506(.A1(new_n2762_), .A2(new_n2760_), .ZN(new_n2763_));
  NOR3_X1    g02507(.A1(new_n2751_), .A2(new_n2763_), .A3(new_n2755_), .ZN(new_n2764_));
  OAI21_X1   g02508(.A1(new_n2753_), .A2(new_n2754_), .B(new_n2752_), .ZN(new_n2765_));
  NAND3_X1   g02509(.A1(new_n2687_), .A2(new_n2745_), .A3(new_n2750_), .ZN(new_n2766_));
  OAI21_X1   g02510(.A1(new_n2761_), .A2(new_n2757_), .B(\a[17] ), .ZN(new_n2767_));
  NAND3_X1   g02511(.A1(new_n2759_), .A2(new_n1344_), .A3(new_n2758_), .ZN(new_n2768_));
  NAND2_X1   g02512(.A1(new_n2767_), .A2(new_n2768_), .ZN(new_n2769_));
  AOI21_X1   g02513(.A1(new_n2765_), .A2(new_n2766_), .B(new_n2769_), .ZN(new_n2770_));
  NOR2_X1    g02514(.A1(new_n2764_), .A2(new_n2770_), .ZN(new_n2771_));
  NOR3_X1    g02515(.A1(new_n2771_), .A2(new_n2684_), .A3(new_n2570_), .ZN(new_n2772_));
  OAI21_X1   g02516(.A1(new_n2566_), .A2(new_n2561_), .B(new_n2556_), .ZN(new_n2773_));
  NAND3_X1   g02517(.A1(new_n2765_), .A2(new_n2766_), .A3(new_n2769_), .ZN(new_n2774_));
  OAI21_X1   g02518(.A1(new_n2751_), .A2(new_n2755_), .B(new_n2763_), .ZN(new_n2775_));
  NAND2_X1   g02519(.A1(new_n2775_), .A2(new_n2774_), .ZN(new_n2776_));
  AOI21_X1   g02520(.A1(new_n2574_), .A2(new_n2773_), .B(new_n2776_), .ZN(new_n2777_));
  AOI22_X1   g02521(.A1(new_n1006_), .A2(\b[13] ), .B1(\b[12] ), .B2(new_n1009_), .ZN(new_n2778_));
  OAI21_X1   g02522(.A1(new_n852_), .A2(new_n1481_), .B(new_n2778_), .ZN(new_n2779_));
  INV_X1     g02523(.I(new_n2779_), .ZN(new_n2780_));
  NAND3_X1   g02524(.A1(new_n1081_), .A2(new_n1013_), .A3(new_n1078_), .ZN(new_n2781_));
  AOI21_X1   g02525(.A1(new_n2781_), .A2(new_n2780_), .B(new_n1002_), .ZN(new_n2782_));
  NOR3_X1    g02526(.A1(new_n1816_), .A2(new_n1323_), .A3(new_n1817_), .ZN(new_n2783_));
  NOR3_X1    g02527(.A1(new_n2783_), .A2(\a[14] ), .A3(new_n2779_), .ZN(new_n2784_));
  NOR2_X1    g02528(.A1(new_n2784_), .A2(new_n2782_), .ZN(new_n2785_));
  NOR3_X1    g02529(.A1(new_n2777_), .A2(new_n2785_), .A3(new_n2772_), .ZN(new_n2786_));
  NAND3_X1   g02530(.A1(new_n2776_), .A2(new_n2773_), .A3(new_n2574_), .ZN(new_n2787_));
  NAND2_X1   g02531(.A1(new_n2773_), .A2(new_n2574_), .ZN(new_n2788_));
  NAND2_X1   g02532(.A1(new_n2788_), .A2(new_n2771_), .ZN(new_n2789_));
  OAI21_X1   g02533(.A1(new_n2783_), .A2(new_n2779_), .B(\a[14] ), .ZN(new_n2790_));
  NAND3_X1   g02534(.A1(new_n2781_), .A2(new_n1002_), .A3(new_n2780_), .ZN(new_n2791_));
  NAND2_X1   g02535(.A1(new_n2790_), .A2(new_n2791_), .ZN(new_n2792_));
  AOI21_X1   g02536(.A1(new_n2789_), .A2(new_n2787_), .B(new_n2792_), .ZN(new_n2793_));
  NOR2_X1    g02537(.A1(new_n2793_), .A2(new_n2786_), .ZN(new_n2794_));
  OAI21_X1   g02538(.A1(new_n2683_), .A2(new_n2584_), .B(new_n2794_), .ZN(new_n2795_));
  NAND2_X1   g02539(.A1(new_n2586_), .A2(new_n2577_), .ZN(new_n2796_));
  NAND3_X1   g02540(.A1(new_n2789_), .A2(new_n2792_), .A3(new_n2787_), .ZN(new_n2797_));
  OAI21_X1   g02541(.A1(new_n2777_), .A2(new_n2772_), .B(new_n2785_), .ZN(new_n2798_));
  NAND2_X1   g02542(.A1(new_n2797_), .A2(new_n2798_), .ZN(new_n2799_));
  NAND3_X1   g02543(.A1(new_n2796_), .A2(new_n2587_), .A3(new_n2799_), .ZN(new_n2800_));
  NAND3_X1   g02544(.A1(new_n2800_), .A2(new_n2795_), .A3(new_n2680_), .ZN(new_n2801_));
  INV_X1     g02545(.I(new_n2680_), .ZN(new_n2802_));
  AOI21_X1   g02546(.A1(new_n2796_), .A2(new_n2587_), .B(new_n2799_), .ZN(new_n2803_));
  NOR3_X1    g02547(.A1(new_n2683_), .A2(new_n2794_), .A3(new_n2584_), .ZN(new_n2804_));
  OAI21_X1   g02548(.A1(new_n2803_), .A2(new_n2804_), .B(new_n2802_), .ZN(new_n2805_));
  NAND2_X1   g02549(.A1(new_n2805_), .A2(new_n2801_), .ZN(new_n2806_));
  NAND3_X1   g02550(.A1(new_n2676_), .A2(new_n2600_), .A3(new_n2806_), .ZN(new_n2807_));
  AOI21_X1   g02551(.A1(new_n2274_), .A2(new_n2275_), .B(new_n2271_), .ZN(new_n2808_));
  OAI21_X1   g02552(.A1(new_n2808_), .A2(new_n2428_), .B(new_n2427_), .ZN(new_n2809_));
  AOI21_X1   g02553(.A1(new_n2809_), .A2(new_n2594_), .B(new_n2589_), .ZN(new_n2810_));
  NOR3_X1    g02554(.A1(new_n2803_), .A2(new_n2804_), .A3(new_n2802_), .ZN(new_n2811_));
  AOI21_X1   g02555(.A1(new_n2800_), .A2(new_n2795_), .B(new_n2680_), .ZN(new_n2812_));
  NOR2_X1    g02556(.A1(new_n2811_), .A2(new_n2812_), .ZN(new_n2813_));
  OAI21_X1   g02557(.A1(new_n2810_), .A2(new_n2597_), .B(new_n2813_), .ZN(new_n2814_));
  NAND3_X1   g02558(.A1(new_n2814_), .A2(new_n2807_), .A3(new_n2673_), .ZN(new_n2815_));
  INV_X1     g02559(.I(new_n2670_), .ZN(new_n2816_));
  NAND2_X1   g02560(.A1(new_n2816_), .A2(new_n2671_), .ZN(new_n2817_));
  NOR3_X1    g02561(.A1(new_n2810_), .A2(new_n2597_), .A3(new_n2813_), .ZN(new_n2818_));
  AOI21_X1   g02562(.A1(new_n2676_), .A2(new_n2600_), .B(new_n2806_), .ZN(new_n2819_));
  OAI21_X1   g02563(.A1(new_n2818_), .A2(new_n2819_), .B(new_n2817_), .ZN(new_n2820_));
  AND2_X2    g02564(.A1(new_n2820_), .A2(new_n2815_), .Z(new_n2821_));
  NAND2_X1   g02565(.A1(new_n2665_), .A2(new_n2821_), .ZN(new_n2822_));
  OAI21_X1   g02566(.A1(new_n2602_), .A2(new_n2609_), .B(new_n2620_), .ZN(new_n2823_));
  NAND2_X1   g02567(.A1(new_n2820_), .A2(new_n2815_), .ZN(new_n2824_));
  NAND2_X1   g02568(.A1(new_n2823_), .A2(new_n2824_), .ZN(new_n2825_));
  AOI21_X1   g02569(.A1(new_n2825_), .A2(new_n2822_), .B(new_n2664_), .ZN(new_n2826_));
  OAI21_X1   g02570(.A1(new_n2449_), .A2(new_n2448_), .B(new_n2447_), .ZN(new_n2827_));
  AOI21_X1   g02571(.A1(new_n2827_), .A2(new_n2607_), .B(new_n2602_), .ZN(new_n2828_));
  NOR3_X1    g02572(.A1(new_n2828_), .A2(new_n2617_), .A3(new_n2824_), .ZN(new_n2829_));
  NOR2_X1    g02573(.A1(new_n2665_), .A2(new_n2821_), .ZN(new_n2830_));
  NOR3_X1    g02574(.A1(new_n2830_), .A2(new_n2663_), .A3(new_n2829_), .ZN(new_n2831_));
  NOR2_X1    g02575(.A1(new_n2826_), .A2(new_n2831_), .ZN(new_n2832_));
  XNOR2_X1   g02576(.A1(new_n2658_), .A2(new_n2832_), .ZN(new_n2833_));
  INV_X1     g02577(.I(new_n2833_), .ZN(new_n2834_));
  NOR2_X1    g02578(.A1(new_n2834_), .A2(new_n2657_), .ZN(new_n2835_));
  NAND2_X1   g02579(.A1(new_n2834_), .A2(new_n2657_), .ZN(new_n2836_));
  INV_X1     g02580(.I(new_n2836_), .ZN(new_n2837_));
  NOR2_X1    g02581(.A1(new_n2837_), .A2(new_n2835_), .ZN(new_n2838_));
  XOR2_X1    g02582(.A1(new_n2838_), .A2(new_n2645_), .Z(\f[25] ));
  INV_X1     g02583(.I(new_n2624_), .ZN(new_n2840_));
  NAND2_X1   g02584(.A1(new_n2626_), .A2(new_n2622_), .ZN(new_n2841_));
  NAND2_X1   g02585(.A1(new_n2841_), .A2(new_n2840_), .ZN(new_n2842_));
  INV_X1     g02586(.I(new_n2832_), .ZN(new_n2843_));
  NOR3_X1    g02587(.A1(new_n2830_), .A2(new_n2664_), .A3(new_n2829_), .ZN(new_n2844_));
  AOI21_X1   g02588(.A1(new_n2842_), .A2(new_n2843_), .B(new_n2844_), .ZN(new_n2845_));
  AOI22_X1   g02589(.A1(new_n800_), .A2(\b[22] ), .B1(\b[23] ), .B2(new_n333_), .ZN(new_n2846_));
  OAI21_X1   g02590(.A1(new_n2027_), .A2(new_n392_), .B(new_n2846_), .ZN(new_n2847_));
  AOI21_X1   g02591(.A1(new_n2470_), .A2(new_n330_), .B(new_n2847_), .ZN(new_n2848_));
  XOR2_X1    g02592(.A1(new_n2848_), .A2(new_n312_), .Z(new_n2849_));
  INV_X1     g02593(.I(new_n2849_), .ZN(new_n2850_));
  AOI21_X1   g02594(.A1(new_n2800_), .A2(new_n2795_), .B(new_n2802_), .ZN(new_n2851_));
  AOI22_X1   g02595(.A1(new_n729_), .A2(\b[17] ), .B1(\b[16] ), .B2(new_n732_), .ZN(new_n2852_));
  OAI21_X1   g02596(.A1(new_n1268_), .A2(new_n1127_), .B(new_n2852_), .ZN(new_n2853_));
  INV_X1     g02597(.I(new_n2853_), .ZN(new_n2854_));
  NOR2_X1    g02598(.A1(new_n1441_), .A2(new_n1442_), .ZN(new_n2855_));
  NOR4_X1    g02599(.A1(new_n1435_), .A2(new_n1436_), .A3(new_n1438_), .A4(new_n1439_), .ZN(new_n2856_));
  NOR2_X1    g02600(.A1(new_n2855_), .A2(new_n2856_), .ZN(new_n2857_));
  NAND2_X1   g02601(.A1(new_n2857_), .A2(new_n724_), .ZN(new_n2858_));
  AOI21_X1   g02602(.A1(new_n2858_), .A2(new_n2854_), .B(new_n722_), .ZN(new_n2859_));
  OAI21_X1   g02603(.A1(new_n1444_), .A2(new_n986_), .B(new_n2854_), .ZN(new_n2860_));
  NOR2_X1    g02604(.A1(new_n2860_), .A2(\a[11] ), .ZN(new_n2861_));
  NOR2_X1    g02605(.A1(new_n2859_), .A2(new_n2861_), .ZN(new_n2862_));
  AOI22_X1   g02606(.A1(new_n1006_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n1009_), .ZN(new_n2863_));
  OAI21_X1   g02607(.A1(new_n941_), .A2(new_n1481_), .B(new_n2863_), .ZN(new_n2864_));
  INV_X1     g02608(.I(new_n2864_), .ZN(new_n2865_));
  OAI21_X1   g02609(.A1(new_n1103_), .A2(new_n1323_), .B(new_n2865_), .ZN(new_n2866_));
  NAND2_X1   g02610(.A1(new_n2866_), .A2(\a[14] ), .ZN(new_n2867_));
  INV_X1     g02611(.I(new_n2867_), .ZN(new_n2868_));
  NOR2_X1    g02612(.A1(new_n2866_), .A2(\a[14] ), .ZN(new_n2869_));
  NOR2_X1    g02613(.A1(new_n2868_), .A2(new_n2869_), .ZN(new_n2870_));
  OAI21_X1   g02614(.A1(new_n2684_), .A2(new_n2570_), .B(new_n2775_), .ZN(new_n2871_));
  AOI22_X1   g02615(.A1(new_n1586_), .A2(\b[11] ), .B1(\b[10] ), .B2(new_n1495_), .ZN(new_n2872_));
  OAI21_X1   g02616(.A1(new_n667_), .A2(new_n1917_), .B(new_n2872_), .ZN(new_n2873_));
  INV_X1     g02617(.I(new_n2873_), .ZN(new_n2874_));
  OAI21_X1   g02618(.A1(new_n859_), .A2(new_n1732_), .B(new_n2874_), .ZN(new_n2875_));
  NAND2_X1   g02619(.A1(new_n2875_), .A2(\a[17] ), .ZN(new_n2876_));
  INV_X1     g02620(.I(new_n2876_), .ZN(new_n2877_));
  NOR2_X1    g02621(.A1(new_n2875_), .A2(\a[17] ), .ZN(new_n2878_));
  OAI21_X1   g02622(.A1(new_n2752_), .A2(new_n2754_), .B(new_n2745_), .ZN(new_n2879_));
  OAI22_X1   g02623(.A1(new_n1751_), .A2(new_n577_), .B1(new_n471_), .B2(new_n1754_), .ZN(new_n2880_));
  NOR2_X1    g02624(.A1(new_n1931_), .A2(new_n438_), .ZN(new_n2881_));
  NOR2_X1    g02625(.A1(new_n2880_), .A2(new_n2881_), .ZN(new_n2882_));
  OAI21_X1   g02626(.A1(new_n587_), .A2(new_n1757_), .B(new_n2882_), .ZN(new_n2883_));
  NAND2_X1   g02627(.A1(new_n2883_), .A2(\a[20] ), .ZN(new_n2884_));
  INV_X1     g02628(.I(new_n2882_), .ZN(new_n2885_));
  AOI21_X1   g02629(.A1(new_n799_), .A2(new_n1746_), .B(new_n2885_), .ZN(new_n2886_));
  NAND2_X1   g02630(.A1(new_n2886_), .A2(new_n1736_), .ZN(new_n2887_));
  OAI21_X1   g02631(.A1(new_n2691_), .A2(new_n2738_), .B(new_n2730_), .ZN(new_n2888_));
  NAND3_X1   g02632(.A1(new_n2888_), .A2(new_n2887_), .A3(new_n2884_), .ZN(new_n2889_));
  NOR2_X1    g02633(.A1(new_n2886_), .A2(new_n1736_), .ZN(new_n2890_));
  NOR2_X1    g02634(.A1(new_n2883_), .A2(\a[20] ), .ZN(new_n2891_));
  AOI21_X1   g02635(.A1(new_n2736_), .A2(new_n2731_), .B(new_n2737_), .ZN(new_n2892_));
  OAI21_X1   g02636(.A1(new_n2891_), .A2(new_n2890_), .B(new_n2892_), .ZN(new_n2893_));
  OAI22_X1   g02637(.A1(new_n2189_), .A2(new_n377_), .B1(new_n339_), .B2(new_n2194_), .ZN(new_n2894_));
  NOR2_X1    g02638(.A1(new_n2370_), .A2(new_n290_), .ZN(new_n2895_));
  NOR2_X1    g02639(.A1(new_n2894_), .A2(new_n2895_), .ZN(new_n2896_));
  OAI21_X1   g02640(.A1(new_n566_), .A2(new_n2197_), .B(new_n2896_), .ZN(new_n2897_));
  NAND2_X1   g02641(.A1(new_n2897_), .A2(\a[23] ), .ZN(new_n2898_));
  INV_X1     g02642(.I(new_n2898_), .ZN(new_n2899_));
  NOR2_X1    g02643(.A1(new_n2897_), .A2(\a[23] ), .ZN(new_n2900_));
  NAND2_X1   g02644(.A1(new_n2722_), .A2(new_n554_), .ZN(new_n2901_));
  NAND2_X1   g02645(.A1(new_n2716_), .A2(\b[2] ), .ZN(new_n2902_));
  NAND2_X1   g02646(.A1(new_n2719_), .A2(\b[1] ), .ZN(new_n2903_));
  AOI21_X1   g02647(.A1(new_n2704_), .A2(\a[26] ), .B(\a[23] ), .ZN(new_n2904_));
  AOI21_X1   g02648(.A1(\a[25] ), .A2(new_n2714_), .B(new_n2200_), .ZN(new_n2905_));
  NOR3_X1    g02649(.A1(new_n2701_), .A2(new_n2904_), .A3(new_n2905_), .ZN(new_n2906_));
  NAND2_X1   g02650(.A1(new_n2906_), .A2(\b[0] ), .ZN(new_n2907_));
  NAND4_X1   g02651(.A1(new_n2901_), .A2(new_n2907_), .A3(new_n2902_), .A4(new_n2903_), .ZN(new_n2908_));
  XOR2_X1    g02652(.A1(new_n2908_), .A2(\a[26] ), .Z(new_n2909_));
  NOR3_X1    g02653(.A1(new_n2727_), .A2(new_n2714_), .A3(new_n2534_), .ZN(new_n2910_));
  NOR2_X1    g02654(.A1(new_n2909_), .A2(new_n2910_), .ZN(new_n2911_));
  NOR4_X1    g02655(.A1(new_n2908_), .A2(new_n2727_), .A3(new_n2714_), .A4(new_n2534_), .ZN(new_n2912_));
  NOR4_X1    g02656(.A1(new_n2911_), .A2(new_n2899_), .A3(new_n2900_), .A4(new_n2912_), .ZN(new_n2913_));
  INV_X1     g02657(.I(new_n2900_), .ZN(new_n2914_));
  XOR2_X1    g02658(.A1(new_n2908_), .A2(new_n2714_), .Z(new_n2915_));
  INV_X1     g02659(.I(new_n2910_), .ZN(new_n2916_));
  NAND2_X1   g02660(.A1(new_n2915_), .A2(new_n2916_), .ZN(new_n2917_));
  NOR2_X1    g02661(.A1(new_n2709_), .A2(new_n2712_), .ZN(new_n2918_));
  NOR2_X1    g02662(.A1(new_n2711_), .A2(new_n282_), .ZN(new_n2919_));
  NOR2_X1    g02663(.A1(new_n2703_), .A2(new_n276_), .ZN(new_n2920_));
  INV_X1     g02664(.I(new_n2903_), .ZN(new_n2921_));
  INV_X1     g02665(.I(new_n2904_), .ZN(new_n2922_));
  OAI21_X1   g02666(.A1(new_n2704_), .A2(\a[26] ), .B(\a[23] ), .ZN(new_n2923_));
  NAND3_X1   g02667(.A1(new_n2922_), .A2(new_n2533_), .A3(new_n2923_), .ZN(new_n2924_));
  NOR2_X1    g02668(.A1(new_n2924_), .A2(new_n258_), .ZN(new_n2925_));
  NOR4_X1    g02669(.A1(new_n2919_), .A2(new_n2925_), .A3(new_n2921_), .A4(new_n2920_), .ZN(new_n2926_));
  NAND4_X1   g02670(.A1(new_n2926_), .A2(\a[26] ), .A3(new_n2918_), .A4(new_n2535_), .ZN(new_n2927_));
  AOI22_X1   g02671(.A1(new_n2917_), .A2(new_n2927_), .B1(new_n2914_), .B2(new_n2898_), .ZN(new_n2928_));
  NOR2_X1    g02672(.A1(new_n2928_), .A2(new_n2913_), .ZN(new_n2929_));
  NAND3_X1   g02673(.A1(new_n2889_), .A2(new_n2893_), .A3(new_n2929_), .ZN(new_n2930_));
  NOR3_X1    g02674(.A1(new_n2890_), .A2(new_n2891_), .A3(new_n2892_), .ZN(new_n2931_));
  AOI21_X1   g02675(.A1(new_n2884_), .A2(new_n2887_), .B(new_n2888_), .ZN(new_n2932_));
  NAND4_X1   g02676(.A1(new_n2917_), .A2(new_n2914_), .A3(new_n2898_), .A4(new_n2927_), .ZN(new_n2933_));
  OAI22_X1   g02677(.A1(new_n2911_), .A2(new_n2912_), .B1(new_n2899_), .B2(new_n2900_), .ZN(new_n2934_));
  NAND2_X1   g02678(.A1(new_n2934_), .A2(new_n2933_), .ZN(new_n2935_));
  OAI21_X1   g02679(.A1(new_n2932_), .A2(new_n2931_), .B(new_n2935_), .ZN(new_n2936_));
  NAND2_X1   g02680(.A1(new_n2936_), .A2(new_n2930_), .ZN(new_n2937_));
  NOR2_X1    g02681(.A1(new_n2937_), .A2(new_n2879_), .ZN(new_n2938_));
  AOI21_X1   g02682(.A1(new_n2687_), .A2(new_n2750_), .B(new_n2753_), .ZN(new_n2939_));
  NOR3_X1    g02683(.A1(new_n2932_), .A2(new_n2931_), .A3(new_n2935_), .ZN(new_n2940_));
  AOI21_X1   g02684(.A1(new_n2889_), .A2(new_n2893_), .B(new_n2929_), .ZN(new_n2941_));
  NOR2_X1    g02685(.A1(new_n2940_), .A2(new_n2941_), .ZN(new_n2942_));
  NOR2_X1    g02686(.A1(new_n2939_), .A2(new_n2942_), .ZN(new_n2943_));
  NOR4_X1    g02687(.A1(new_n2943_), .A2(new_n2877_), .A3(new_n2938_), .A4(new_n2878_), .ZN(new_n2944_));
  NAND2_X1   g02688(.A1(new_n2325_), .A2(new_n1354_), .ZN(new_n2945_));
  NAND3_X1   g02689(.A1(new_n2945_), .A2(new_n1344_), .A3(new_n2874_), .ZN(new_n2946_));
  NAND2_X1   g02690(.A1(new_n2939_), .A2(new_n2942_), .ZN(new_n2947_));
  NAND2_X1   g02691(.A1(new_n2937_), .A2(new_n2879_), .ZN(new_n2948_));
  AOI22_X1   g02692(.A1(new_n2947_), .A2(new_n2948_), .B1(new_n2876_), .B2(new_n2946_), .ZN(new_n2949_));
  NOR2_X1    g02693(.A1(new_n2944_), .A2(new_n2949_), .ZN(new_n2950_));
  NAND3_X1   g02694(.A1(new_n2950_), .A2(new_n2871_), .A3(new_n2774_), .ZN(new_n2951_));
  NAND2_X1   g02695(.A1(new_n2871_), .A2(new_n2774_), .ZN(new_n2952_));
  NAND4_X1   g02696(.A1(new_n2947_), .A2(new_n2948_), .A3(new_n2876_), .A4(new_n2946_), .ZN(new_n2953_));
  OAI22_X1   g02697(.A1(new_n2943_), .A2(new_n2938_), .B1(new_n2877_), .B2(new_n2878_), .ZN(new_n2954_));
  NAND2_X1   g02698(.A1(new_n2954_), .A2(new_n2953_), .ZN(new_n2955_));
  NAND2_X1   g02699(.A1(new_n2952_), .A2(new_n2955_), .ZN(new_n2956_));
  AOI21_X1   g02700(.A1(new_n2956_), .A2(new_n2951_), .B(new_n2870_), .ZN(new_n2957_));
  INV_X1     g02701(.I(new_n2869_), .ZN(new_n2958_));
  NAND2_X1   g02702(.A1(new_n2958_), .A2(new_n2867_), .ZN(new_n2959_));
  AOI21_X1   g02703(.A1(new_n2773_), .A2(new_n2574_), .B(new_n2770_), .ZN(new_n2960_));
  NOR3_X1    g02704(.A1(new_n2955_), .A2(new_n2960_), .A3(new_n2764_), .ZN(new_n2961_));
  AOI21_X1   g02705(.A1(new_n2774_), .A2(new_n2871_), .B(new_n2950_), .ZN(new_n2962_));
  NOR3_X1    g02706(.A1(new_n2962_), .A2(new_n2959_), .A3(new_n2961_), .ZN(new_n2963_));
  NOR2_X1    g02707(.A1(new_n2957_), .A2(new_n2963_), .ZN(new_n2964_));
  NOR3_X1    g02708(.A1(new_n2683_), .A2(new_n2584_), .A3(new_n2786_), .ZN(new_n2965_));
  OAI21_X1   g02709(.A1(new_n2965_), .A2(new_n2793_), .B(new_n2964_), .ZN(new_n2966_));
  OAI21_X1   g02710(.A1(new_n2962_), .A2(new_n2961_), .B(new_n2959_), .ZN(new_n2967_));
  NAND3_X1   g02711(.A1(new_n2956_), .A2(new_n2951_), .A3(new_n2870_), .ZN(new_n2968_));
  NAND2_X1   g02712(.A1(new_n2968_), .A2(new_n2967_), .ZN(new_n2969_));
  NAND3_X1   g02713(.A1(new_n2796_), .A2(new_n2587_), .A3(new_n2797_), .ZN(new_n2970_));
  NAND3_X1   g02714(.A1(new_n2970_), .A2(new_n2798_), .A3(new_n2969_), .ZN(new_n2971_));
  NAND3_X1   g02715(.A1(new_n2971_), .A2(new_n2966_), .A3(new_n2862_), .ZN(new_n2972_));
  XOR2_X1    g02716(.A1(new_n2860_), .A2(new_n722_), .Z(new_n2973_));
  AOI21_X1   g02717(.A1(new_n2970_), .A2(new_n2798_), .B(new_n2969_), .ZN(new_n2974_));
  NOR3_X1    g02718(.A1(new_n2965_), .A2(new_n2964_), .A3(new_n2793_), .ZN(new_n2975_));
  OAI21_X1   g02719(.A1(new_n2974_), .A2(new_n2975_), .B(new_n2973_), .ZN(new_n2976_));
  NAND2_X1   g02720(.A1(new_n2976_), .A2(new_n2972_), .ZN(new_n2977_));
  OAI21_X1   g02721(.A1(new_n2818_), .A2(new_n2851_), .B(new_n2977_), .ZN(new_n2978_));
  INV_X1     g02722(.I(new_n2851_), .ZN(new_n2979_));
  NOR3_X1    g02723(.A1(new_n2974_), .A2(new_n2973_), .A3(new_n2975_), .ZN(new_n2980_));
  AOI21_X1   g02724(.A1(new_n2971_), .A2(new_n2966_), .B(new_n2862_), .ZN(new_n2981_));
  NOR2_X1    g02725(.A1(new_n2980_), .A2(new_n2981_), .ZN(new_n2982_));
  NAND3_X1   g02726(.A1(new_n2807_), .A2(new_n2982_), .A3(new_n2979_), .ZN(new_n2983_));
  AOI22_X1   g02727(.A1(new_n518_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n636_), .ZN(new_n2984_));
  OAI21_X1   g02728(.A1(new_n1553_), .A2(new_n917_), .B(new_n2984_), .ZN(new_n2985_));
  AOI21_X1   g02729(.A1(new_n2452_), .A2(new_n618_), .B(new_n2985_), .ZN(new_n2986_));
  XOR2_X1    g02730(.A1(new_n2986_), .A2(new_n488_), .Z(new_n2987_));
  INV_X1     g02731(.I(new_n2987_), .ZN(new_n2988_));
  NAND3_X1   g02732(.A1(new_n2978_), .A2(new_n2988_), .A3(new_n2983_), .ZN(new_n2989_));
  AOI21_X1   g02733(.A1(new_n2807_), .A2(new_n2979_), .B(new_n2982_), .ZN(new_n2990_));
  NOR3_X1    g02734(.A1(new_n2818_), .A2(new_n2851_), .A3(new_n2977_), .ZN(new_n2991_));
  OAI21_X1   g02735(.A1(new_n2991_), .A2(new_n2990_), .B(new_n2987_), .ZN(new_n2992_));
  NAND2_X1   g02736(.A1(new_n2992_), .A2(new_n2989_), .ZN(new_n2993_));
  NOR3_X1    g02737(.A1(new_n2818_), .A2(new_n2819_), .A3(new_n2817_), .ZN(new_n2994_));
  AOI21_X1   g02738(.A1(new_n2665_), .A2(new_n2821_), .B(new_n2994_), .ZN(new_n2995_));
  NOR2_X1    g02739(.A1(new_n2995_), .A2(new_n2993_), .ZN(new_n2996_));
  NOR3_X1    g02740(.A1(new_n2991_), .A2(new_n2990_), .A3(new_n2987_), .ZN(new_n2997_));
  AOI21_X1   g02741(.A1(new_n2978_), .A2(new_n2983_), .B(new_n2988_), .ZN(new_n2998_));
  NOR2_X1    g02742(.A1(new_n2998_), .A2(new_n2997_), .ZN(new_n2999_));
  OAI21_X1   g02743(.A1(new_n2823_), .A2(new_n2824_), .B(new_n2815_), .ZN(new_n3000_));
  NOR2_X1    g02744(.A1(new_n3000_), .A2(new_n2999_), .ZN(new_n3001_));
  OAI21_X1   g02745(.A1(new_n2996_), .A2(new_n3001_), .B(new_n2850_), .ZN(new_n3002_));
  INV_X1     g02746(.I(new_n3002_), .ZN(new_n3003_));
  NOR3_X1    g02747(.A1(new_n2996_), .A2(new_n3001_), .A3(new_n2850_), .ZN(new_n3004_));
  NOR2_X1    g02748(.A1(new_n3003_), .A2(new_n3004_), .ZN(new_n3005_));
  INV_X1     g02749(.I(\b[26] ), .ZN(new_n3006_));
  OAI22_X1   g02750(.A1(new_n277_), .A2(new_n3006_), .B1(new_n2646_), .B2(new_n262_), .ZN(new_n3007_));
  AOI21_X1   g02751(.A1(\b[24] ), .A2(new_n283_), .B(new_n3007_), .ZN(new_n3008_));
  OAI21_X1   g02752(.A1(new_n2652_), .A2(new_n2495_), .B(new_n2463_), .ZN(new_n3009_));
  OAI21_X1   g02753(.A1(new_n2502_), .A2(new_n2646_), .B(new_n2495_), .ZN(new_n3010_));
  XNOR2_X1   g02754(.A1(\b[25] ), .A2(\b[26] ), .ZN(new_n3011_));
  AOI21_X1   g02755(.A1(new_n3009_), .A2(new_n3010_), .B(new_n3011_), .ZN(new_n3012_));
  NAND2_X1   g02756(.A1(new_n3009_), .A2(new_n3010_), .ZN(new_n3013_));
  XOR2_X1    g02757(.A1(\b[25] ), .A2(\b[26] ), .Z(new_n3014_));
  NOR2_X1    g02758(.A1(new_n3013_), .A2(new_n3014_), .ZN(new_n3015_));
  NOR2_X1    g02759(.A1(new_n3015_), .A2(new_n3012_), .ZN(new_n3016_));
  OAI21_X1   g02760(.A1(new_n3016_), .A2(new_n279_), .B(new_n3008_), .ZN(new_n3017_));
  XOR2_X1    g02761(.A1(new_n3017_), .A2(\a[2] ), .Z(new_n3018_));
  INV_X1     g02762(.I(new_n3018_), .ZN(new_n3019_));
  NOR2_X1    g02763(.A1(new_n3005_), .A2(new_n3019_), .ZN(new_n3020_));
  NAND2_X1   g02764(.A1(new_n3005_), .A2(new_n3019_), .ZN(new_n3021_));
  INV_X1     g02765(.I(new_n3021_), .ZN(new_n3022_));
  NOR3_X1    g02766(.A1(new_n3022_), .A2(new_n2845_), .A3(new_n3020_), .ZN(new_n3023_));
  INV_X1     g02767(.I(new_n2844_), .ZN(new_n3024_));
  OAI21_X1   g02768(.A1(new_n2658_), .A2(new_n2832_), .B(new_n3024_), .ZN(new_n3025_));
  INV_X1     g02769(.I(new_n3020_), .ZN(new_n3026_));
  AOI21_X1   g02770(.A1(new_n3026_), .A2(new_n3021_), .B(new_n3025_), .ZN(new_n3027_));
  NOR2_X1    g02771(.A1(new_n3027_), .A2(new_n3023_), .ZN(new_n3028_));
  INV_X1     g02772(.I(new_n3028_), .ZN(new_n3029_));
  AOI21_X1   g02773(.A1(new_n2494_), .A2(new_n2634_), .B(new_n2643_), .ZN(new_n3030_));
  AOI21_X1   g02774(.A1(new_n3030_), .A2(new_n2836_), .B(new_n2835_), .ZN(new_n3031_));
  XOR2_X1    g02775(.A1(new_n3031_), .A2(new_n3029_), .Z(\f[26] ));
  INV_X1     g02776(.I(new_n2506_), .ZN(new_n3033_));
  AOI22_X1   g02777(.A1(new_n800_), .A2(\b[23] ), .B1(\b[24] ), .B2(new_n333_), .ZN(new_n3034_));
  OAI21_X1   g02778(.A1(new_n2142_), .A2(new_n392_), .B(new_n3034_), .ZN(new_n3035_));
  AOI21_X1   g02779(.A1(new_n3033_), .A2(new_n330_), .B(new_n3035_), .ZN(new_n3036_));
  XOR2_X1    g02780(.A1(new_n3036_), .A2(new_n312_), .Z(new_n3037_));
  AOI21_X1   g02781(.A1(new_n2888_), .A2(new_n2934_), .B(new_n2913_), .ZN(new_n3038_));
  OAI22_X1   g02782(.A1(new_n2189_), .A2(new_n438_), .B1(new_n377_), .B2(new_n2194_), .ZN(new_n3039_));
  AOI21_X1   g02783(.A1(\b[4] ), .A2(new_n2361_), .B(new_n3039_), .ZN(new_n3040_));
  OAI21_X1   g02784(.A1(new_n450_), .A2(new_n2197_), .B(new_n3040_), .ZN(new_n3041_));
  XOR2_X1    g02785(.A1(new_n3041_), .A2(new_n2200_), .Z(new_n3042_));
  NOR2_X1    g02786(.A1(new_n2924_), .A2(new_n275_), .ZN(new_n3043_));
  OAI22_X1   g02787(.A1(new_n2703_), .A2(new_n290_), .B1(new_n276_), .B2(new_n2708_), .ZN(new_n3044_));
  NOR2_X1    g02788(.A1(new_n429_), .A2(new_n2711_), .ZN(new_n3045_));
  NOR3_X1    g02789(.A1(new_n3045_), .A2(new_n3044_), .A3(new_n3043_), .ZN(new_n3046_));
  NOR2_X1    g02790(.A1(new_n3046_), .A2(new_n2714_), .ZN(new_n3047_));
  NAND2_X1   g02791(.A1(new_n2906_), .A2(\b[1] ), .ZN(new_n3048_));
  AOI22_X1   g02792(.A1(new_n2716_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n2719_), .ZN(new_n3049_));
  NAND2_X1   g02793(.A1(new_n299_), .A2(new_n2722_), .ZN(new_n3050_));
  NAND3_X1   g02794(.A1(new_n3050_), .A2(new_n3049_), .A3(new_n3048_), .ZN(new_n3051_));
  NOR2_X1    g02795(.A1(new_n3051_), .A2(\a[26] ), .ZN(new_n3052_));
  XOR2_X1    g02796(.A1(\a[26] ), .A2(\a[27] ), .Z(new_n3053_));
  NAND2_X1   g02797(.A1(new_n3053_), .A2(\b[0] ), .ZN(new_n3054_));
  INV_X1     g02798(.I(new_n3054_), .ZN(new_n3055_));
  OAI21_X1   g02799(.A1(new_n3047_), .A2(new_n3052_), .B(new_n3055_), .ZN(new_n3056_));
  NAND2_X1   g02800(.A1(new_n3051_), .A2(\a[26] ), .ZN(new_n3057_));
  NAND2_X1   g02801(.A1(new_n3046_), .A2(new_n2714_), .ZN(new_n3058_));
  NAND3_X1   g02802(.A1(new_n3058_), .A2(new_n3057_), .A3(new_n3054_), .ZN(new_n3059_));
  AOI21_X1   g02803(.A1(new_n3056_), .A2(new_n3059_), .B(new_n2912_), .ZN(new_n3060_));
  AOI21_X1   g02804(.A1(new_n3058_), .A2(new_n3057_), .B(new_n3054_), .ZN(new_n3061_));
  NOR3_X1    g02805(.A1(new_n3047_), .A2(new_n3052_), .A3(new_n3055_), .ZN(new_n3062_));
  NOR3_X1    g02806(.A1(new_n3061_), .A2(new_n3062_), .A3(new_n2927_), .ZN(new_n3063_));
  NOR3_X1    g02807(.A1(new_n3042_), .A2(new_n3060_), .A3(new_n3063_), .ZN(new_n3064_));
  NAND2_X1   g02808(.A1(new_n916_), .A2(new_n2208_), .ZN(new_n3065_));
  AOI21_X1   g02809(.A1(new_n3065_), .A2(new_n3040_), .B(new_n2200_), .ZN(new_n3066_));
  NOR2_X1    g02810(.A1(new_n3041_), .A2(\a[23] ), .ZN(new_n3067_));
  NOR2_X1    g02811(.A1(new_n3067_), .A2(new_n3066_), .ZN(new_n3068_));
  OAI21_X1   g02812(.A1(new_n3061_), .A2(new_n3062_), .B(new_n2927_), .ZN(new_n3069_));
  NAND3_X1   g02813(.A1(new_n3056_), .A2(new_n3059_), .A3(new_n2912_), .ZN(new_n3070_));
  AOI21_X1   g02814(.A1(new_n3069_), .A2(new_n3070_), .B(new_n3068_), .ZN(new_n3071_));
  NOR2_X1    g02815(.A1(new_n3064_), .A2(new_n3071_), .ZN(new_n3072_));
  XOR2_X1    g02816(.A1(new_n3072_), .A2(new_n3038_), .Z(new_n3073_));
  AOI22_X1   g02817(.A1(new_n1738_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n1743_), .ZN(new_n3074_));
  OAI21_X1   g02818(.A1(new_n471_), .A2(new_n1931_), .B(new_n3074_), .ZN(new_n3075_));
  AOI21_X1   g02819(.A1(new_n676_), .A2(new_n1746_), .B(new_n3075_), .ZN(new_n3076_));
  XOR2_X1    g02820(.A1(new_n3076_), .A2(new_n1736_), .Z(new_n3077_));
  NOR2_X1    g02821(.A1(new_n2890_), .A2(new_n2891_), .ZN(new_n3078_));
  NAND2_X1   g02822(.A1(new_n2929_), .A2(new_n2888_), .ZN(new_n3079_));
  NAND2_X1   g02823(.A1(new_n2935_), .A2(new_n2892_), .ZN(new_n3080_));
  NAND3_X1   g02824(.A1(new_n3079_), .A2(new_n3080_), .A3(new_n3078_), .ZN(new_n3081_));
  OAI21_X1   g02825(.A1(new_n2937_), .A2(new_n2879_), .B(new_n3081_), .ZN(new_n3082_));
  NAND2_X1   g02826(.A1(new_n3082_), .A2(new_n3077_), .ZN(new_n3083_));
  INV_X1     g02827(.I(new_n3077_), .ZN(new_n3084_));
  AND2_X2    g02828(.A1(new_n3079_), .A2(new_n3080_), .Z(new_n3085_));
  AOI22_X1   g02829(.A1(new_n2939_), .A2(new_n2942_), .B1(new_n3085_), .B2(new_n3078_), .ZN(new_n3086_));
  NAND2_X1   g02830(.A1(new_n3086_), .A2(new_n3084_), .ZN(new_n3087_));
  NAND3_X1   g02831(.A1(new_n3087_), .A2(new_n3073_), .A3(new_n3083_), .ZN(new_n3088_));
  INV_X1     g02832(.I(new_n3073_), .ZN(new_n3089_));
  NOR2_X1    g02833(.A1(new_n3086_), .A2(new_n3084_), .ZN(new_n3090_));
  NOR2_X1    g02834(.A1(new_n3082_), .A2(new_n3077_), .ZN(new_n3091_));
  OAI21_X1   g02835(.A1(new_n3090_), .A2(new_n3091_), .B(new_n3089_), .ZN(new_n3092_));
  NAND2_X1   g02836(.A1(new_n3092_), .A2(new_n3088_), .ZN(new_n3093_));
  INV_X1     g02837(.I(new_n3093_), .ZN(new_n3094_));
  OAI22_X1   g02838(.A1(new_n1592_), .A2(new_n941_), .B1(new_n852_), .B2(new_n1505_), .ZN(new_n3095_));
  AOI21_X1   g02839(.A1(\b[10] ), .A2(new_n1584_), .B(new_n3095_), .ZN(new_n3096_));
  OAI21_X1   g02840(.A1(new_n953_), .A2(new_n1732_), .B(new_n3096_), .ZN(new_n3097_));
  XOR2_X1    g02841(.A1(new_n3097_), .A2(\a[17] ), .Z(new_n3098_));
  OAI21_X1   g02842(.A1(new_n2961_), .A2(new_n2944_), .B(new_n3098_), .ZN(new_n3099_));
  INV_X1     g02843(.I(new_n3098_), .ZN(new_n3100_));
  NAND3_X1   g02844(.A1(new_n2951_), .A2(new_n2953_), .A3(new_n3100_), .ZN(new_n3101_));
  NAND3_X1   g02845(.A1(new_n3099_), .A2(new_n3101_), .A3(new_n3094_), .ZN(new_n3102_));
  NAND2_X1   g02846(.A1(new_n3099_), .A2(new_n3101_), .ZN(new_n3103_));
  NAND2_X1   g02847(.A1(new_n3103_), .A2(new_n3093_), .ZN(new_n3104_));
  NAND2_X1   g02848(.A1(new_n3104_), .A2(new_n3102_), .ZN(new_n3105_));
  OAI22_X1   g02849(.A1(new_n993_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n997_), .ZN(new_n3106_));
  AOI21_X1   g02850(.A1(\b[13] ), .A2(new_n1486_), .B(new_n3106_), .ZN(new_n3107_));
  OAI21_X1   g02851(.A1(new_n1275_), .A2(new_n1323_), .B(new_n3107_), .ZN(new_n3108_));
  XOR2_X1    g02852(.A1(new_n3108_), .A2(\a[14] ), .Z(new_n3109_));
  INV_X1     g02853(.I(new_n3109_), .ZN(new_n3110_));
  AOI21_X1   g02854(.A1(new_n2966_), .A2(new_n2968_), .B(new_n3110_), .ZN(new_n3111_));
  NOR3_X1    g02855(.A1(new_n2974_), .A2(new_n2963_), .A3(new_n3109_), .ZN(new_n3112_));
  NOR3_X1    g02856(.A1(new_n3112_), .A2(new_n3111_), .A3(new_n3105_), .ZN(new_n3113_));
  XOR2_X1    g02857(.A1(new_n3103_), .A2(new_n3093_), .Z(new_n3114_));
  OAI21_X1   g02858(.A1(new_n2974_), .A2(new_n2963_), .B(new_n3109_), .ZN(new_n3115_));
  NAND3_X1   g02859(.A1(new_n2966_), .A2(new_n2968_), .A3(new_n3110_), .ZN(new_n3116_));
  AOI21_X1   g02860(.A1(new_n3115_), .A2(new_n3116_), .B(new_n3114_), .ZN(new_n3117_));
  NOR2_X1    g02861(.A1(new_n3113_), .A2(new_n3117_), .ZN(new_n3118_));
  INV_X1     g02862(.I(new_n3118_), .ZN(new_n3119_));
  OAI22_X1   g02863(.A1(new_n713_), .A2(new_n1553_), .B1(new_n1432_), .B2(new_n717_), .ZN(new_n3120_));
  AOI21_X1   g02864(.A1(\b[16] ), .A2(new_n1126_), .B(new_n3120_), .ZN(new_n3121_));
  OAI21_X1   g02865(.A1(new_n1563_), .A2(new_n986_), .B(new_n3121_), .ZN(new_n3122_));
  XOR2_X1    g02866(.A1(new_n3122_), .A2(\a[11] ), .Z(new_n3123_));
  INV_X1     g02867(.I(new_n3123_), .ZN(new_n3124_));
  OAI21_X1   g02868(.A1(new_n2818_), .A2(new_n2851_), .B(new_n2982_), .ZN(new_n3125_));
  AOI21_X1   g02869(.A1(new_n3125_), .A2(new_n2972_), .B(new_n3124_), .ZN(new_n3126_));
  AOI21_X1   g02870(.A1(new_n2807_), .A2(new_n2979_), .B(new_n2977_), .ZN(new_n3127_));
  NOR3_X1    g02871(.A1(new_n3127_), .A2(new_n2980_), .A3(new_n3123_), .ZN(new_n3128_));
  NOR3_X1    g02872(.A1(new_n3126_), .A2(new_n3128_), .A3(new_n3119_), .ZN(new_n3129_));
  OAI21_X1   g02873(.A1(new_n3127_), .A2(new_n2980_), .B(new_n3123_), .ZN(new_n3130_));
  NAND3_X1   g02874(.A1(new_n3125_), .A2(new_n2972_), .A3(new_n3124_), .ZN(new_n3131_));
  AOI21_X1   g02875(.A1(new_n3131_), .A2(new_n3130_), .B(new_n3118_), .ZN(new_n3132_));
  NOR2_X1    g02876(.A1(new_n3129_), .A2(new_n3132_), .ZN(new_n3133_));
  AOI22_X1   g02877(.A1(new_n518_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n636_), .ZN(new_n3134_));
  OAI21_X1   g02878(.A1(new_n1859_), .A2(new_n917_), .B(new_n3134_), .ZN(new_n3135_));
  AOI21_X1   g02879(.A1(new_n2032_), .A2(new_n618_), .B(new_n3135_), .ZN(new_n3136_));
  XOR2_X1    g02880(.A1(new_n3136_), .A2(new_n488_), .Z(new_n3137_));
  OAI21_X1   g02881(.A1(new_n2995_), .A2(new_n2993_), .B(new_n2992_), .ZN(new_n3138_));
  NAND2_X1   g02882(.A1(new_n3138_), .A2(new_n3137_), .ZN(new_n3139_));
  OAI21_X1   g02883(.A1(new_n2829_), .A2(new_n2994_), .B(new_n2999_), .ZN(new_n3140_));
  INV_X1     g02884(.I(new_n3137_), .ZN(new_n3141_));
  NAND3_X1   g02885(.A1(new_n3140_), .A2(new_n2992_), .A3(new_n3141_), .ZN(new_n3142_));
  NAND3_X1   g02886(.A1(new_n3139_), .A2(new_n3142_), .A3(new_n3133_), .ZN(new_n3143_));
  OR2_X2     g02887(.A1(new_n3129_), .A2(new_n3132_), .Z(new_n3144_));
  AOI21_X1   g02888(.A1(new_n3140_), .A2(new_n2992_), .B(new_n3141_), .ZN(new_n3145_));
  NOR2_X1    g02889(.A1(new_n3138_), .A2(new_n3137_), .ZN(new_n3146_));
  OAI21_X1   g02890(.A1(new_n3146_), .A2(new_n3145_), .B(new_n3144_), .ZN(new_n3147_));
  AOI21_X1   g02891(.A1(new_n3147_), .A2(new_n3143_), .B(new_n3037_), .ZN(new_n3148_));
  INV_X1     g02892(.I(new_n3148_), .ZN(new_n3149_));
  NAND3_X1   g02893(.A1(new_n3147_), .A2(new_n3143_), .A3(new_n3037_), .ZN(new_n3150_));
  OAI21_X1   g02894(.A1(new_n3025_), .A2(new_n3004_), .B(new_n3002_), .ZN(new_n3151_));
  NAND3_X1   g02895(.A1(new_n3149_), .A2(new_n3150_), .A3(new_n3151_), .ZN(new_n3152_));
  INV_X1     g02896(.I(new_n3150_), .ZN(new_n3153_));
  INV_X1     g02897(.I(new_n3004_), .ZN(new_n3154_));
  AOI21_X1   g02898(.A1(new_n2845_), .A2(new_n3154_), .B(new_n3003_), .ZN(new_n3155_));
  OAI21_X1   g02899(.A1(new_n3148_), .A2(new_n3153_), .B(new_n3155_), .ZN(new_n3156_));
  NAND2_X1   g02900(.A1(new_n3156_), .A2(new_n3152_), .ZN(new_n3157_));
  INV_X1     g02901(.I(\b[27] ), .ZN(new_n3158_));
  OAI22_X1   g02902(.A1(new_n277_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n262_), .ZN(new_n3159_));
  AOI21_X1   g02903(.A1(\b[25] ), .A2(new_n283_), .B(new_n3159_), .ZN(new_n3160_));
  NAND2_X1   g02904(.A1(new_n3013_), .A2(new_n2646_), .ZN(new_n3161_));
  NOR2_X1    g02905(.A1(new_n3013_), .A2(new_n2646_), .ZN(new_n3162_));
  NAND2_X1   g02906(.A1(new_n3162_), .A2(new_n3006_), .ZN(new_n3163_));
  OAI21_X1   g02907(.A1(new_n3006_), .A2(new_n3161_), .B(new_n3163_), .ZN(new_n3164_));
  XOR2_X1    g02908(.A1(new_n3164_), .A2(new_n3158_), .Z(new_n3165_));
  OAI21_X1   g02909(.A1(new_n3165_), .A2(new_n279_), .B(new_n3160_), .ZN(new_n3166_));
  XOR2_X1    g02910(.A1(new_n3166_), .A2(\a[2] ), .Z(new_n3167_));
  INV_X1     g02911(.I(new_n3167_), .ZN(new_n3168_));
  OAI21_X1   g02912(.A1(new_n3003_), .A2(new_n3004_), .B(new_n3025_), .ZN(new_n3169_));
  NAND2_X1   g02913(.A1(new_n2845_), .A2(new_n3005_), .ZN(new_n3170_));
  AOI21_X1   g02914(.A1(new_n3170_), .A2(new_n3169_), .B(new_n3019_), .ZN(new_n3171_));
  AOI21_X1   g02915(.A1(new_n3031_), .A2(new_n3029_), .B(new_n3171_), .ZN(new_n3172_));
  NOR2_X1    g02916(.A1(new_n3172_), .A2(new_n3168_), .ZN(new_n3173_));
  INV_X1     g02917(.I(new_n2835_), .ZN(new_n3174_));
  OAI21_X1   g02918(.A1(new_n2645_), .A2(new_n2837_), .B(new_n3174_), .ZN(new_n3175_));
  INV_X1     g02919(.I(new_n3171_), .ZN(new_n3176_));
  OAI21_X1   g02920(.A1(new_n3175_), .A2(new_n3028_), .B(new_n3176_), .ZN(new_n3177_));
  NOR2_X1    g02921(.A1(new_n3177_), .A2(new_n3167_), .ZN(new_n3178_));
  NOR2_X1    g02922(.A1(new_n3178_), .A2(new_n3173_), .ZN(new_n3179_));
  XOR2_X1    g02923(.A1(new_n3179_), .A2(new_n3157_), .Z(\f[27] ));
  NAND2_X1   g02924(.A1(new_n3172_), .A2(new_n3168_), .ZN(new_n3181_));
  INV_X1     g02925(.I(new_n3157_), .ZN(new_n3182_));
  OAI21_X1   g02926(.A1(new_n3172_), .A2(new_n3168_), .B(new_n3182_), .ZN(new_n3183_));
  NAND2_X1   g02927(.A1(new_n3183_), .A2(new_n3181_), .ZN(new_n3184_));
  INV_X1     g02928(.I(\b[28] ), .ZN(new_n3185_));
  OAI22_X1   g02929(.A1(new_n277_), .A2(new_n3185_), .B1(new_n3158_), .B2(new_n262_), .ZN(new_n3186_));
  AOI21_X1   g02930(.A1(\b[26] ), .A2(new_n283_), .B(new_n3186_), .ZN(new_n3187_));
  XOR2_X1    g02931(.A1(\b[27] ), .A2(\b[28] ), .Z(new_n3188_));
  OAI21_X1   g02932(.A1(new_n3162_), .A2(\b[26] ), .B(\b[27] ), .ZN(new_n3189_));
  NAND2_X1   g02933(.A1(new_n3161_), .A2(\b[26] ), .ZN(new_n3190_));
  NAND2_X1   g02934(.A1(new_n3189_), .A2(new_n3190_), .ZN(new_n3191_));
  INV_X1     g02935(.I(new_n3191_), .ZN(new_n3192_));
  NOR2_X1    g02936(.A1(new_n3192_), .A2(new_n3188_), .ZN(new_n3193_));
  INV_X1     g02937(.I(new_n3188_), .ZN(new_n3194_));
  NOR2_X1    g02938(.A1(new_n3191_), .A2(new_n3194_), .ZN(new_n3195_));
  NOR2_X1    g02939(.A1(new_n3193_), .A2(new_n3195_), .ZN(new_n3196_));
  OAI21_X1   g02940(.A1(new_n3196_), .A2(new_n279_), .B(new_n3187_), .ZN(new_n3197_));
  XOR2_X1    g02941(.A1(new_n3197_), .A2(\a[2] ), .Z(new_n3198_));
  OAI21_X1   g02942(.A1(new_n3151_), .A2(new_n3148_), .B(new_n3150_), .ZN(new_n3199_));
  AOI22_X1   g02943(.A1(new_n800_), .A2(\b[24] ), .B1(\b[25] ), .B2(new_n333_), .ZN(new_n3200_));
  OAI21_X1   g02944(.A1(new_n2463_), .A2(new_n392_), .B(new_n3200_), .ZN(new_n3201_));
  INV_X1     g02945(.I(new_n3201_), .ZN(new_n3202_));
  OAI21_X1   g02946(.A1(new_n2655_), .A2(new_n318_), .B(new_n3202_), .ZN(new_n3203_));
  XOR2_X1    g02947(.A1(new_n3203_), .A2(new_n312_), .Z(new_n3204_));
  AOI21_X1   g02948(.A1(new_n3000_), .A2(new_n2999_), .B(new_n2998_), .ZN(new_n3205_));
  OAI21_X1   g02949(.A1(new_n3205_), .A2(new_n3141_), .B(new_n3144_), .ZN(new_n3206_));
  AOI22_X1   g02950(.A1(new_n518_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n636_), .ZN(new_n3207_));
  OAI21_X1   g02951(.A1(new_n1860_), .A2(new_n917_), .B(new_n3207_), .ZN(new_n3208_));
  AOI21_X1   g02952(.A1(new_n2659_), .A2(new_n618_), .B(new_n3208_), .ZN(new_n3209_));
  XOR2_X1    g02953(.A1(new_n3209_), .A2(new_n488_), .Z(new_n3210_));
  INV_X1     g02954(.I(new_n3210_), .ZN(new_n3211_));
  AOI21_X1   g02955(.A1(new_n2590_), .A2(new_n2599_), .B(new_n2597_), .ZN(new_n3212_));
  AOI21_X1   g02956(.A1(new_n3212_), .A2(new_n2806_), .B(new_n2851_), .ZN(new_n3213_));
  OAI21_X1   g02957(.A1(new_n3213_), .A2(new_n2977_), .B(new_n2972_), .ZN(new_n3214_));
  AOI21_X1   g02958(.A1(new_n3214_), .A2(new_n3123_), .B(new_n3118_), .ZN(new_n3215_));
  AOI22_X1   g02959(.A1(new_n729_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n732_), .ZN(new_n3216_));
  OAI21_X1   g02960(.A1(new_n1432_), .A2(new_n1127_), .B(new_n3216_), .ZN(new_n3217_));
  INV_X1     g02961(.I(new_n3217_), .ZN(new_n3218_));
  NAND2_X1   g02962(.A1(new_n1695_), .A2(new_n724_), .ZN(new_n3219_));
  AOI21_X1   g02963(.A1(new_n3219_), .A2(new_n3218_), .B(new_n722_), .ZN(new_n3220_));
  NAND3_X1   g02964(.A1(new_n3219_), .A2(new_n722_), .A3(new_n3218_), .ZN(new_n3221_));
  INV_X1     g02965(.I(new_n3221_), .ZN(new_n3222_));
  NOR2_X1    g02966(.A1(new_n3222_), .A2(new_n3220_), .ZN(new_n3223_));
  OAI21_X1   g02967(.A1(new_n2576_), .A2(new_n2583_), .B(new_n2587_), .ZN(new_n3224_));
  OAI21_X1   g02968(.A1(new_n3224_), .A2(new_n2786_), .B(new_n2798_), .ZN(new_n3225_));
  AOI21_X1   g02969(.A1(new_n3225_), .A2(new_n2964_), .B(new_n2963_), .ZN(new_n3226_));
  OAI21_X1   g02970(.A1(new_n3226_), .A2(new_n3110_), .B(new_n3105_), .ZN(new_n3227_));
  OAI22_X1   g02971(.A1(new_n993_), .A2(new_n1296_), .B1(new_n1268_), .B2(new_n997_), .ZN(new_n3228_));
  AOI21_X1   g02972(.A1(\b[14] ), .A2(new_n1486_), .B(new_n3228_), .ZN(new_n3229_));
  OAI21_X1   g02973(.A1(new_n1306_), .A2(new_n1323_), .B(new_n3229_), .ZN(new_n3230_));
  XOR2_X1    g02974(.A1(new_n3230_), .A2(\a[14] ), .Z(new_n3231_));
  AOI21_X1   g02975(.A1(new_n3082_), .A2(new_n3077_), .B(new_n3073_), .ZN(new_n3232_));
  OAI21_X1   g02976(.A1(new_n2892_), .A2(new_n2928_), .B(new_n2933_), .ZN(new_n3233_));
  NAND3_X1   g02977(.A1(new_n3068_), .A2(new_n3069_), .A3(new_n3070_), .ZN(new_n3234_));
  OAI21_X1   g02978(.A1(new_n3060_), .A2(new_n3063_), .B(new_n3042_), .ZN(new_n3235_));
  NAND2_X1   g02979(.A1(new_n3235_), .A2(new_n3234_), .ZN(new_n3236_));
  OAI21_X1   g02980(.A1(new_n3060_), .A2(new_n3063_), .B(new_n3068_), .ZN(new_n3237_));
  INV_X1     g02981(.I(new_n3237_), .ZN(new_n3238_));
  AOI21_X1   g02982(.A1(new_n3236_), .A2(new_n3233_), .B(new_n3238_), .ZN(new_n3239_));
  NOR2_X1    g02983(.A1(new_n3047_), .A2(new_n3052_), .ZN(new_n3240_));
  NAND2_X1   g02984(.A1(new_n2927_), .A2(new_n3054_), .ZN(new_n3241_));
  NOR2_X1    g02985(.A1(new_n2927_), .A2(new_n3054_), .ZN(new_n3242_));
  AOI21_X1   g02986(.A1(new_n3240_), .A2(new_n3241_), .B(new_n3242_), .ZN(new_n3243_));
  AOI22_X1   g02987(.A1(new_n2716_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n2719_), .ZN(new_n3244_));
  NAND2_X1   g02988(.A1(new_n2906_), .A2(\b[2] ), .ZN(new_n3245_));
  NAND2_X1   g02989(.A1(new_n1725_), .A2(new_n2722_), .ZN(new_n3246_));
  NAND3_X1   g02990(.A1(new_n3246_), .A2(new_n3244_), .A3(new_n3245_), .ZN(new_n3247_));
  NAND2_X1   g02991(.A1(new_n3247_), .A2(\a[26] ), .ZN(new_n3248_));
  NAND4_X1   g02992(.A1(new_n3246_), .A2(new_n2714_), .A3(new_n3244_), .A4(new_n3245_), .ZN(new_n3249_));
  NAND2_X1   g02993(.A1(new_n3248_), .A2(new_n3249_), .ZN(new_n3250_));
  INV_X1     g02994(.I(new_n3250_), .ZN(new_n3251_));
  XNOR2_X1   g02995(.A1(\a[28] ), .A2(\a[29] ), .ZN(new_n3252_));
  NAND2_X1   g02996(.A1(new_n3252_), .A2(new_n3053_), .ZN(new_n3253_));
  INV_X1     g02997(.I(\a[28] ), .ZN(new_n3254_));
  NOR3_X1    g02998(.A1(new_n3254_), .A2(\a[26] ), .A3(\a[27] ), .ZN(new_n3255_));
  NAND3_X1   g02999(.A1(new_n3254_), .A2(\a[26] ), .A3(\a[27] ), .ZN(new_n3256_));
  INV_X1     g03000(.I(new_n3256_), .ZN(new_n3257_));
  NOR2_X1    g03001(.A1(new_n3257_), .A2(new_n3255_), .ZN(new_n3258_));
  OAI22_X1   g03002(.A1(new_n275_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n258_), .ZN(new_n3259_));
  XOR2_X1    g03003(.A1(\a[28] ), .A2(\a[29] ), .Z(new_n3260_));
  NAND2_X1   g03004(.A1(new_n3053_), .A2(new_n3260_), .ZN(new_n3261_));
  NOR2_X1    g03005(.A1(new_n3261_), .A2(new_n313_), .ZN(new_n3262_));
  OAI21_X1   g03006(.A1(new_n3259_), .A2(new_n3262_), .B(\a[29] ), .ZN(new_n3263_));
  INV_X1     g03007(.I(\a[29] ), .ZN(new_n3264_));
  XNOR2_X1   g03008(.A1(\a[26] ), .A2(\a[27] ), .ZN(new_n3265_));
  XOR2_X1    g03009(.A1(\a[28] ), .A2(\a[29] ), .Z(new_n3266_));
  NOR2_X1    g03010(.A1(new_n3265_), .A2(new_n3266_), .ZN(new_n3267_));
  INV_X1     g03011(.I(\a[27] ), .ZN(new_n3268_));
  NAND3_X1   g03012(.A1(new_n2714_), .A2(new_n3268_), .A3(\a[28] ), .ZN(new_n3269_));
  NAND2_X1   g03013(.A1(new_n3269_), .A2(new_n3256_), .ZN(new_n3270_));
  AOI22_X1   g03014(.A1(new_n3267_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n3270_), .ZN(new_n3271_));
  XNOR2_X1   g03015(.A1(\a[28] ), .A2(\a[29] ), .ZN(new_n3272_));
  NOR2_X1    g03016(.A1(new_n3265_), .A2(new_n3272_), .ZN(new_n3273_));
  NAND2_X1   g03017(.A1(new_n3273_), .A2(new_n263_), .ZN(new_n3274_));
  NAND3_X1   g03018(.A1(new_n3271_), .A2(new_n3274_), .A3(new_n3264_), .ZN(new_n3275_));
  NAND2_X1   g03019(.A1(new_n3054_), .A2(\a[29] ), .ZN(new_n3276_));
  NAND3_X1   g03020(.A1(new_n3263_), .A2(new_n3275_), .A3(new_n3276_), .ZN(new_n3277_));
  NAND2_X1   g03021(.A1(new_n3271_), .A2(new_n3274_), .ZN(new_n3278_));
  NAND3_X1   g03022(.A1(new_n3278_), .A2(\a[29] ), .A3(new_n3054_), .ZN(new_n3279_));
  NAND2_X1   g03023(.A1(new_n3277_), .A2(new_n3279_), .ZN(new_n3280_));
  NAND2_X1   g03024(.A1(new_n3251_), .A2(new_n3280_), .ZN(new_n3281_));
  NAND3_X1   g03025(.A1(new_n3250_), .A2(new_n3277_), .A3(new_n3279_), .ZN(new_n3282_));
  AOI21_X1   g03026(.A1(new_n3281_), .A2(new_n3282_), .B(new_n3243_), .ZN(new_n3283_));
  NAND2_X1   g03027(.A1(new_n3058_), .A2(new_n3057_), .ZN(new_n3284_));
  NOR2_X1    g03028(.A1(new_n2912_), .A2(new_n3055_), .ZN(new_n3285_));
  NAND2_X1   g03029(.A1(new_n2912_), .A2(new_n3055_), .ZN(new_n3286_));
  OAI21_X1   g03030(.A1(new_n3284_), .A2(new_n3285_), .B(new_n3286_), .ZN(new_n3287_));
  AOI21_X1   g03031(.A1(new_n3277_), .A2(new_n3279_), .B(new_n3250_), .ZN(new_n3288_));
  NOR2_X1    g03032(.A1(new_n3251_), .A2(new_n3280_), .ZN(new_n3289_));
  NOR3_X1    g03033(.A1(new_n3289_), .A2(new_n3287_), .A3(new_n3288_), .ZN(new_n3290_));
  NOR2_X1    g03034(.A1(new_n3283_), .A2(new_n3290_), .ZN(new_n3291_));
  OAI22_X1   g03035(.A1(new_n2189_), .A2(new_n471_), .B1(new_n438_), .B2(new_n2194_), .ZN(new_n3292_));
  AOI21_X1   g03036(.A1(\b[5] ), .A2(new_n2361_), .B(new_n3292_), .ZN(new_n3293_));
  OAI21_X1   g03037(.A1(new_n485_), .A2(new_n2197_), .B(new_n3293_), .ZN(new_n3294_));
  XOR2_X1    g03038(.A1(new_n3294_), .A2(new_n2200_), .Z(new_n3295_));
  NAND2_X1   g03039(.A1(new_n3291_), .A2(new_n3295_), .ZN(new_n3296_));
  OAI21_X1   g03040(.A1(new_n3289_), .A2(new_n3288_), .B(new_n3287_), .ZN(new_n3297_));
  NAND3_X1   g03041(.A1(new_n3281_), .A2(new_n3243_), .A3(new_n3282_), .ZN(new_n3298_));
  NAND2_X1   g03042(.A1(new_n3298_), .A2(new_n3297_), .ZN(new_n3299_));
  XOR2_X1    g03043(.A1(new_n3294_), .A2(\a[23] ), .Z(new_n3300_));
  NAND2_X1   g03044(.A1(new_n3299_), .A2(new_n3300_), .ZN(new_n3301_));
  AOI21_X1   g03045(.A1(new_n3296_), .A2(new_n3301_), .B(new_n3239_), .ZN(new_n3302_));
  NAND3_X1   g03046(.A1(new_n3239_), .A2(new_n3296_), .A3(new_n3301_), .ZN(new_n3303_));
  INV_X1     g03047(.I(new_n3303_), .ZN(new_n3304_));
  AOI22_X1   g03048(.A1(new_n1738_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n1743_), .ZN(new_n3305_));
  OAI21_X1   g03049(.A1(new_n577_), .A2(new_n1931_), .B(new_n3305_), .ZN(new_n3306_));
  INV_X1     g03050(.I(new_n3306_), .ZN(new_n3307_));
  OAI21_X1   g03051(.A1(new_n786_), .A2(new_n1757_), .B(new_n3307_), .ZN(new_n3308_));
  XOR2_X1    g03052(.A1(new_n3308_), .A2(\a[20] ), .Z(new_n3309_));
  NOR3_X1    g03053(.A1(new_n3304_), .A2(new_n3302_), .A3(new_n3309_), .ZN(new_n3310_));
  OAI21_X1   g03054(.A1(new_n3072_), .A2(new_n3038_), .B(new_n3237_), .ZN(new_n3311_));
  NAND2_X1   g03055(.A1(new_n3296_), .A2(new_n3301_), .ZN(new_n3312_));
  NAND2_X1   g03056(.A1(new_n3312_), .A2(new_n3311_), .ZN(new_n3313_));
  XOR2_X1    g03057(.A1(new_n3308_), .A2(new_n1736_), .Z(new_n3314_));
  AOI21_X1   g03058(.A1(new_n3313_), .A2(new_n3303_), .B(new_n3314_), .ZN(new_n3315_));
  NOR2_X1    g03059(.A1(new_n3310_), .A2(new_n3315_), .ZN(new_n3316_));
  NOR3_X1    g03060(.A1(new_n3316_), .A2(new_n3232_), .A3(new_n3091_), .ZN(new_n3317_));
  OAI21_X1   g03061(.A1(new_n3086_), .A2(new_n3084_), .B(new_n3089_), .ZN(new_n3318_));
  NAND3_X1   g03062(.A1(new_n3313_), .A2(new_n3314_), .A3(new_n3303_), .ZN(new_n3319_));
  OAI21_X1   g03063(.A1(new_n3304_), .A2(new_n3302_), .B(new_n3309_), .ZN(new_n3320_));
  NAND2_X1   g03064(.A1(new_n3320_), .A2(new_n3319_), .ZN(new_n3321_));
  AOI21_X1   g03065(.A1(new_n3318_), .A2(new_n3087_), .B(new_n3321_), .ZN(new_n3322_));
  AOI22_X1   g03066(.A1(new_n1586_), .A2(\b[13] ), .B1(\b[12] ), .B2(new_n1495_), .ZN(new_n3323_));
  OAI21_X1   g03067(.A1(new_n852_), .A2(new_n1917_), .B(new_n3323_), .ZN(new_n3324_));
  INV_X1     g03068(.I(new_n3324_), .ZN(new_n3325_));
  NAND3_X1   g03069(.A1(new_n1081_), .A2(new_n1078_), .A3(new_n1354_), .ZN(new_n3326_));
  AOI21_X1   g03070(.A1(new_n3326_), .A2(new_n3325_), .B(new_n1344_), .ZN(new_n3327_));
  NAND3_X1   g03071(.A1(new_n3326_), .A2(new_n1344_), .A3(new_n3325_), .ZN(new_n3328_));
  INV_X1     g03072(.I(new_n3328_), .ZN(new_n3329_));
  NOR2_X1    g03073(.A1(new_n3329_), .A2(new_n3327_), .ZN(new_n3330_));
  NOR3_X1    g03074(.A1(new_n3322_), .A2(new_n3330_), .A3(new_n3317_), .ZN(new_n3331_));
  NAND3_X1   g03075(.A1(new_n3321_), .A2(new_n3318_), .A3(new_n3087_), .ZN(new_n3332_));
  OAI21_X1   g03076(.A1(new_n3091_), .A2(new_n3232_), .B(new_n3316_), .ZN(new_n3333_));
  NOR3_X1    g03077(.A1(new_n1816_), .A2(new_n1817_), .A3(new_n1732_), .ZN(new_n3334_));
  OAI21_X1   g03078(.A1(new_n3334_), .A2(new_n3324_), .B(\a[17] ), .ZN(new_n3335_));
  NAND2_X1   g03079(.A1(new_n3335_), .A2(new_n3328_), .ZN(new_n3336_));
  AOI21_X1   g03080(.A1(new_n3333_), .A2(new_n3332_), .B(new_n3336_), .ZN(new_n3337_));
  NOR2_X1    g03081(.A1(new_n3331_), .A2(new_n3337_), .ZN(new_n3338_));
  AOI21_X1   g03082(.A1(new_n2951_), .A2(new_n2953_), .B(new_n3100_), .ZN(new_n3339_));
  OAI21_X1   g03083(.A1(new_n3094_), .A2(new_n3339_), .B(new_n3101_), .ZN(new_n3340_));
  NAND2_X1   g03084(.A1(new_n3340_), .A2(new_n3338_), .ZN(new_n3341_));
  NAND3_X1   g03085(.A1(new_n3333_), .A2(new_n3332_), .A3(new_n3336_), .ZN(new_n3342_));
  OAI21_X1   g03086(.A1(new_n3322_), .A2(new_n3317_), .B(new_n3330_), .ZN(new_n3343_));
  NAND2_X1   g03087(.A1(new_n3343_), .A2(new_n3342_), .ZN(new_n3344_));
  NOR2_X1    g03088(.A1(new_n2960_), .A2(new_n2764_), .ZN(new_n3345_));
  AOI21_X1   g03089(.A1(new_n3345_), .A2(new_n2950_), .B(new_n2944_), .ZN(new_n3346_));
  OAI21_X1   g03090(.A1(new_n3346_), .A2(new_n3100_), .B(new_n3093_), .ZN(new_n3347_));
  NAND3_X1   g03091(.A1(new_n3347_), .A2(new_n3344_), .A3(new_n3101_), .ZN(new_n3348_));
  NAND3_X1   g03092(.A1(new_n3341_), .A2(new_n3348_), .A3(new_n3231_), .ZN(new_n3349_));
  INV_X1     g03093(.I(new_n3231_), .ZN(new_n3350_));
  AOI21_X1   g03094(.A1(new_n3347_), .A2(new_n3101_), .B(new_n3344_), .ZN(new_n3351_));
  NOR2_X1    g03095(.A1(new_n3340_), .A2(new_n3338_), .ZN(new_n3352_));
  OAI21_X1   g03096(.A1(new_n3352_), .A2(new_n3351_), .B(new_n3350_), .ZN(new_n3353_));
  NAND2_X1   g03097(.A1(new_n3353_), .A2(new_n3349_), .ZN(new_n3354_));
  NAND3_X1   g03098(.A1(new_n3227_), .A2(new_n3354_), .A3(new_n3116_), .ZN(new_n3355_));
  NOR2_X1    g03099(.A1(new_n2965_), .A2(new_n2793_), .ZN(new_n3356_));
  OAI21_X1   g03100(.A1(new_n3356_), .A2(new_n2969_), .B(new_n2968_), .ZN(new_n3357_));
  AOI21_X1   g03101(.A1(new_n3357_), .A2(new_n3109_), .B(new_n3114_), .ZN(new_n3358_));
  NOR3_X1    g03102(.A1(new_n3352_), .A2(new_n3351_), .A3(new_n3350_), .ZN(new_n3359_));
  AOI21_X1   g03103(.A1(new_n3341_), .A2(new_n3348_), .B(new_n3231_), .ZN(new_n3360_));
  NOR2_X1    g03104(.A1(new_n3359_), .A2(new_n3360_), .ZN(new_n3361_));
  OAI21_X1   g03105(.A1(new_n3358_), .A2(new_n3112_), .B(new_n3361_), .ZN(new_n3362_));
  NAND3_X1   g03106(.A1(new_n3362_), .A2(new_n3355_), .A3(new_n3223_), .ZN(new_n3363_));
  INV_X1     g03107(.I(new_n3220_), .ZN(new_n3364_));
  NAND2_X1   g03108(.A1(new_n3364_), .A2(new_n3221_), .ZN(new_n3365_));
  NOR3_X1    g03109(.A1(new_n3358_), .A2(new_n3112_), .A3(new_n3361_), .ZN(new_n3366_));
  AOI21_X1   g03110(.A1(new_n3227_), .A2(new_n3116_), .B(new_n3354_), .ZN(new_n3367_));
  OAI21_X1   g03111(.A1(new_n3366_), .A2(new_n3367_), .B(new_n3365_), .ZN(new_n3368_));
  NAND2_X1   g03112(.A1(new_n3368_), .A2(new_n3363_), .ZN(new_n3369_));
  NOR3_X1    g03113(.A1(new_n3215_), .A2(new_n3128_), .A3(new_n3369_), .ZN(new_n3370_));
  OAI21_X1   g03114(.A1(new_n3215_), .A2(new_n3128_), .B(new_n3369_), .ZN(new_n3371_));
  INV_X1     g03115(.I(new_n3371_), .ZN(new_n3372_));
  OAI21_X1   g03116(.A1(new_n3372_), .A2(new_n3370_), .B(new_n3211_), .ZN(new_n3373_));
  OAI21_X1   g03117(.A1(new_n2589_), .A2(new_n2596_), .B(new_n2600_), .ZN(new_n3374_));
  OAI21_X1   g03118(.A1(new_n3374_), .A2(new_n2813_), .B(new_n2979_), .ZN(new_n3375_));
  AOI21_X1   g03119(.A1(new_n3375_), .A2(new_n2982_), .B(new_n2980_), .ZN(new_n3376_));
  OAI21_X1   g03120(.A1(new_n3376_), .A2(new_n3124_), .B(new_n3119_), .ZN(new_n3377_));
  NOR3_X1    g03121(.A1(new_n3366_), .A2(new_n3367_), .A3(new_n3365_), .ZN(new_n3378_));
  AOI21_X1   g03122(.A1(new_n3362_), .A2(new_n3355_), .B(new_n3223_), .ZN(new_n3379_));
  NOR2_X1    g03123(.A1(new_n3378_), .A2(new_n3379_), .ZN(new_n3380_));
  NAND3_X1   g03124(.A1(new_n3377_), .A2(new_n3131_), .A3(new_n3380_), .ZN(new_n3381_));
  NAND3_X1   g03125(.A1(new_n3381_), .A2(new_n3371_), .A3(new_n3210_), .ZN(new_n3382_));
  NAND2_X1   g03126(.A1(new_n3373_), .A2(new_n3382_), .ZN(new_n3383_));
  AOI21_X1   g03127(.A1(new_n3206_), .A2(new_n3142_), .B(new_n3383_), .ZN(new_n3384_));
  AOI21_X1   g03128(.A1(new_n3138_), .A2(new_n3137_), .B(new_n3133_), .ZN(new_n3385_));
  AOI21_X1   g03129(.A1(new_n3381_), .A2(new_n3371_), .B(new_n3210_), .ZN(new_n3386_));
  INV_X1     g03130(.I(new_n3382_), .ZN(new_n3387_));
  NOR2_X1    g03131(.A1(new_n3387_), .A2(new_n3386_), .ZN(new_n3388_));
  NOR3_X1    g03132(.A1(new_n3388_), .A2(new_n3385_), .A3(new_n3146_), .ZN(new_n3389_));
  NOR3_X1    g03133(.A1(new_n3384_), .A2(new_n3389_), .A3(new_n3204_), .ZN(new_n3390_));
  XOR2_X1    g03134(.A1(new_n3203_), .A2(\a[5] ), .Z(new_n3391_));
  OAI21_X1   g03135(.A1(new_n3385_), .A2(new_n3146_), .B(new_n3388_), .ZN(new_n3392_));
  NAND3_X1   g03136(.A1(new_n3383_), .A2(new_n3206_), .A3(new_n3142_), .ZN(new_n3393_));
  AOI21_X1   g03137(.A1(new_n3392_), .A2(new_n3393_), .B(new_n3391_), .ZN(new_n3394_));
  NOR2_X1    g03138(.A1(new_n3394_), .A2(new_n3390_), .ZN(new_n3395_));
  XOR2_X1    g03139(.A1(new_n3395_), .A2(new_n3199_), .Z(new_n3396_));
  INV_X1     g03140(.I(new_n3396_), .ZN(new_n3397_));
  NOR2_X1    g03141(.A1(new_n3397_), .A2(new_n3198_), .ZN(new_n3398_));
  INV_X1     g03142(.I(new_n3398_), .ZN(new_n3399_));
  NAND2_X1   g03143(.A1(new_n3397_), .A2(new_n3198_), .ZN(new_n3400_));
  NAND2_X1   g03144(.A1(new_n3399_), .A2(new_n3400_), .ZN(new_n3401_));
  XOR2_X1    g03145(.A1(new_n3184_), .A2(new_n3401_), .Z(\f[28] ));
  AOI21_X1   g03146(.A1(new_n3155_), .A2(new_n3149_), .B(new_n3153_), .ZN(new_n3403_));
  AOI21_X1   g03147(.A1(new_n3392_), .A2(new_n3393_), .B(new_n3204_), .ZN(new_n3404_));
  INV_X1     g03148(.I(new_n3404_), .ZN(new_n3405_));
  OAI21_X1   g03149(.A1(new_n3403_), .A2(new_n3395_), .B(new_n3405_), .ZN(new_n3406_));
  INV_X1     g03150(.I(new_n3016_), .ZN(new_n3407_));
  AOI22_X1   g03151(.A1(new_n800_), .A2(\b[25] ), .B1(\b[26] ), .B2(new_n333_), .ZN(new_n3408_));
  OAI21_X1   g03152(.A1(new_n2495_), .A2(new_n392_), .B(new_n3408_), .ZN(new_n3409_));
  AOI21_X1   g03153(.A1(new_n3407_), .A2(new_n330_), .B(new_n3409_), .ZN(new_n3410_));
  XOR2_X1    g03154(.A1(new_n3410_), .A2(new_n312_), .Z(new_n3411_));
  AOI22_X1   g03155(.A1(new_n1006_), .A2(\b[17] ), .B1(\b[16] ), .B2(new_n1009_), .ZN(new_n3412_));
  OAI21_X1   g03156(.A1(new_n1268_), .A2(new_n1481_), .B(new_n3412_), .ZN(new_n3413_));
  INV_X1     g03157(.I(new_n3413_), .ZN(new_n3414_));
  NAND2_X1   g03158(.A1(new_n2857_), .A2(new_n1013_), .ZN(new_n3415_));
  AOI21_X1   g03159(.A1(new_n3415_), .A2(new_n3414_), .B(new_n1002_), .ZN(new_n3416_));
  OAI21_X1   g03160(.A1(new_n1444_), .A2(new_n1323_), .B(new_n3414_), .ZN(new_n3417_));
  NOR2_X1    g03161(.A1(new_n3417_), .A2(\a[14] ), .ZN(new_n3418_));
  OR2_X2     g03162(.A1(new_n3416_), .A2(new_n3418_), .Z(new_n3419_));
  AOI22_X1   g03163(.A1(new_n1586_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n1495_), .ZN(new_n3420_));
  OAI21_X1   g03164(.A1(new_n941_), .A2(new_n1917_), .B(new_n3420_), .ZN(new_n3421_));
  AOI21_X1   g03165(.A1(new_n1449_), .A2(new_n1354_), .B(new_n3421_), .ZN(new_n3422_));
  XOR2_X1    g03166(.A1(new_n3422_), .A2(\a[17] ), .Z(new_n3423_));
  AOI21_X1   g03167(.A1(new_n3318_), .A2(new_n3087_), .B(new_n3315_), .ZN(new_n3424_));
  AOI22_X1   g03168(.A1(new_n1738_), .A2(\b[11] ), .B1(\b[10] ), .B2(new_n1743_), .ZN(new_n3425_));
  OAI21_X1   g03169(.A1(new_n667_), .A2(new_n1931_), .B(new_n3425_), .ZN(new_n3426_));
  AOI21_X1   g03170(.A1(new_n2325_), .A2(new_n1746_), .B(new_n3426_), .ZN(new_n3427_));
  NOR2_X1    g03171(.A1(new_n3427_), .A2(new_n1736_), .ZN(new_n3428_));
  INV_X1     g03172(.I(new_n3428_), .ZN(new_n3429_));
  NAND2_X1   g03173(.A1(new_n3427_), .A2(new_n1736_), .ZN(new_n3430_));
  NOR2_X1    g03174(.A1(new_n3299_), .A2(new_n3300_), .ZN(new_n3431_));
  AOI21_X1   g03175(.A1(new_n3239_), .A2(new_n3301_), .B(new_n3431_), .ZN(new_n3432_));
  OAI22_X1   g03176(.A1(new_n2189_), .A2(new_n577_), .B1(new_n471_), .B2(new_n2194_), .ZN(new_n3433_));
  NOR2_X1    g03177(.A1(new_n2370_), .A2(new_n438_), .ZN(new_n3434_));
  NOR2_X1    g03178(.A1(new_n3433_), .A2(new_n3434_), .ZN(new_n3435_));
  INV_X1     g03179(.I(new_n3435_), .ZN(new_n3436_));
  AOI21_X1   g03180(.A1(new_n799_), .A2(new_n2208_), .B(new_n3436_), .ZN(new_n3437_));
  NOR2_X1    g03181(.A1(new_n3437_), .A2(new_n2200_), .ZN(new_n3438_));
  OAI21_X1   g03182(.A1(new_n587_), .A2(new_n2197_), .B(new_n3435_), .ZN(new_n3439_));
  NOR2_X1    g03183(.A1(new_n3439_), .A2(\a[23] ), .ZN(new_n3440_));
  AOI21_X1   g03184(.A1(new_n3287_), .A2(new_n3282_), .B(new_n3288_), .ZN(new_n3441_));
  NOR3_X1    g03185(.A1(new_n3441_), .A2(new_n3438_), .A3(new_n3440_), .ZN(new_n3442_));
  NAND2_X1   g03186(.A1(new_n3439_), .A2(\a[23] ), .ZN(new_n3443_));
  NAND2_X1   g03187(.A1(new_n3437_), .A2(new_n2200_), .ZN(new_n3444_));
  OAI21_X1   g03188(.A1(new_n3243_), .A2(new_n3289_), .B(new_n3281_), .ZN(new_n3445_));
  AOI21_X1   g03189(.A1(new_n3443_), .A2(new_n3444_), .B(new_n3445_), .ZN(new_n3446_));
  OAI22_X1   g03190(.A1(new_n2703_), .A2(new_n377_), .B1(new_n339_), .B2(new_n2708_), .ZN(new_n3447_));
  AOI21_X1   g03191(.A1(\b[3] ), .A2(new_n2906_), .B(new_n3447_), .ZN(new_n3448_));
  OAI21_X1   g03192(.A1(new_n566_), .A2(new_n2711_), .B(new_n3448_), .ZN(new_n3449_));
  XOR2_X1    g03193(.A1(new_n3449_), .A2(\a[26] ), .Z(new_n3450_));
  NAND2_X1   g03194(.A1(new_n3273_), .A2(new_n554_), .ZN(new_n3451_));
  NAND2_X1   g03195(.A1(new_n3267_), .A2(\b[2] ), .ZN(new_n3452_));
  NAND2_X1   g03196(.A1(new_n3270_), .A2(\b[1] ), .ZN(new_n3453_));
  AOI21_X1   g03197(.A1(new_n3254_), .A2(\a[29] ), .B(\a[26] ), .ZN(new_n3454_));
  AOI21_X1   g03198(.A1(\a[28] ), .A2(new_n3264_), .B(new_n2714_), .ZN(new_n3455_));
  NOR3_X1    g03199(.A1(new_n3053_), .A2(new_n3454_), .A3(new_n3455_), .ZN(new_n3456_));
  NAND2_X1   g03200(.A1(new_n3456_), .A2(\b[0] ), .ZN(new_n3457_));
  NAND4_X1   g03201(.A1(new_n3451_), .A2(new_n3457_), .A3(new_n3452_), .A4(new_n3453_), .ZN(new_n3458_));
  XOR2_X1    g03202(.A1(new_n3458_), .A2(\a[29] ), .Z(new_n3459_));
  NOR3_X1    g03203(.A1(new_n3278_), .A2(new_n3264_), .A3(new_n3055_), .ZN(new_n3460_));
  NOR2_X1    g03204(.A1(new_n3459_), .A2(new_n3460_), .ZN(new_n3461_));
  NOR4_X1    g03205(.A1(new_n3458_), .A2(new_n3278_), .A3(new_n3264_), .A4(new_n3055_), .ZN(new_n3462_));
  NOR2_X1    g03206(.A1(new_n3461_), .A2(new_n3462_), .ZN(new_n3463_));
  NAND2_X1   g03207(.A1(new_n3463_), .A2(new_n3450_), .ZN(new_n3464_));
  XOR2_X1    g03208(.A1(new_n3449_), .A2(new_n2714_), .Z(new_n3465_));
  XOR2_X1    g03209(.A1(new_n3458_), .A2(new_n3264_), .Z(new_n3466_));
  INV_X1     g03210(.I(new_n3460_), .ZN(new_n3467_));
  NAND2_X1   g03211(.A1(new_n3466_), .A2(new_n3467_), .ZN(new_n3468_));
  NOR2_X1    g03212(.A1(new_n3259_), .A2(new_n3262_), .ZN(new_n3469_));
  NOR2_X1    g03213(.A1(new_n3261_), .A2(new_n282_), .ZN(new_n3470_));
  NOR2_X1    g03214(.A1(new_n3253_), .A2(new_n276_), .ZN(new_n3471_));
  INV_X1     g03215(.I(new_n3453_), .ZN(new_n3472_));
  INV_X1     g03216(.I(new_n3454_), .ZN(new_n3473_));
  OAI21_X1   g03217(.A1(new_n3254_), .A2(\a[29] ), .B(\a[26] ), .ZN(new_n3474_));
  NAND3_X1   g03218(.A1(new_n3473_), .A2(new_n3265_), .A3(new_n3474_), .ZN(new_n3475_));
  NOR2_X1    g03219(.A1(new_n3475_), .A2(new_n258_), .ZN(new_n3476_));
  NOR4_X1    g03220(.A1(new_n3470_), .A2(new_n3476_), .A3(new_n3472_), .A4(new_n3471_), .ZN(new_n3477_));
  NAND4_X1   g03221(.A1(new_n3477_), .A2(new_n3469_), .A3(\a[29] ), .A4(new_n3054_), .ZN(new_n3478_));
  NAND2_X1   g03222(.A1(new_n3468_), .A2(new_n3478_), .ZN(new_n3479_));
  NAND2_X1   g03223(.A1(new_n3479_), .A2(new_n3465_), .ZN(new_n3480_));
  NAND2_X1   g03224(.A1(new_n3464_), .A2(new_n3480_), .ZN(new_n3481_));
  NOR3_X1    g03225(.A1(new_n3446_), .A2(new_n3481_), .A3(new_n3442_), .ZN(new_n3482_));
  NAND3_X1   g03226(.A1(new_n3445_), .A2(new_n3443_), .A3(new_n3444_), .ZN(new_n3483_));
  OAI21_X1   g03227(.A1(new_n3438_), .A2(new_n3440_), .B(new_n3441_), .ZN(new_n3484_));
  NOR2_X1    g03228(.A1(new_n3479_), .A2(new_n3465_), .ZN(new_n3485_));
  NOR2_X1    g03229(.A1(new_n3463_), .A2(new_n3450_), .ZN(new_n3486_));
  NOR2_X1    g03230(.A1(new_n3486_), .A2(new_n3485_), .ZN(new_n3487_));
  AOI21_X1   g03231(.A1(new_n3484_), .A2(new_n3483_), .B(new_n3487_), .ZN(new_n3488_));
  NOR2_X1    g03232(.A1(new_n3482_), .A2(new_n3488_), .ZN(new_n3489_));
  NAND2_X1   g03233(.A1(new_n3489_), .A2(new_n3432_), .ZN(new_n3490_));
  NOR2_X1    g03234(.A1(new_n3291_), .A2(new_n3295_), .ZN(new_n3491_));
  OAI21_X1   g03235(.A1(new_n3311_), .A2(new_n3491_), .B(new_n3296_), .ZN(new_n3492_));
  NAND3_X1   g03236(.A1(new_n3484_), .A2(new_n3487_), .A3(new_n3483_), .ZN(new_n3493_));
  OAI21_X1   g03237(.A1(new_n3446_), .A2(new_n3442_), .B(new_n3481_), .ZN(new_n3494_));
  NAND2_X1   g03238(.A1(new_n3494_), .A2(new_n3493_), .ZN(new_n3495_));
  NAND2_X1   g03239(.A1(new_n3495_), .A2(new_n3492_), .ZN(new_n3496_));
  NAND4_X1   g03240(.A1(new_n3490_), .A2(new_n3496_), .A3(new_n3429_), .A4(new_n3430_), .ZN(new_n3497_));
  NOR2_X1    g03241(.A1(new_n859_), .A2(new_n1757_), .ZN(new_n3498_));
  NOR3_X1    g03242(.A1(new_n3498_), .A2(\a[20] ), .A3(new_n3426_), .ZN(new_n3499_));
  NOR2_X1    g03243(.A1(new_n3495_), .A2(new_n3492_), .ZN(new_n3500_));
  NOR2_X1    g03244(.A1(new_n3489_), .A2(new_n3432_), .ZN(new_n3501_));
  OAI22_X1   g03245(.A1(new_n3501_), .A2(new_n3500_), .B1(new_n3428_), .B2(new_n3499_), .ZN(new_n3502_));
  NAND2_X1   g03246(.A1(new_n3502_), .A2(new_n3497_), .ZN(new_n3503_));
  NOR3_X1    g03247(.A1(new_n3424_), .A2(new_n3503_), .A3(new_n3310_), .ZN(new_n3504_));
  OAI21_X1   g03248(.A1(new_n3232_), .A2(new_n3091_), .B(new_n3320_), .ZN(new_n3505_));
  NOR4_X1    g03249(.A1(new_n3501_), .A2(new_n3500_), .A3(new_n3428_), .A4(new_n3499_), .ZN(new_n3506_));
  AOI22_X1   g03250(.A1(new_n3490_), .A2(new_n3496_), .B1(new_n3429_), .B2(new_n3430_), .ZN(new_n3507_));
  NOR2_X1    g03251(.A1(new_n3507_), .A2(new_n3506_), .ZN(new_n3508_));
  AOI21_X1   g03252(.A1(new_n3319_), .A2(new_n3505_), .B(new_n3508_), .ZN(new_n3509_));
  OAI21_X1   g03253(.A1(new_n3509_), .A2(new_n3504_), .B(new_n3423_), .ZN(new_n3510_));
  NOR2_X1    g03254(.A1(new_n3422_), .A2(new_n1344_), .ZN(new_n3511_));
  NOR2_X1    g03255(.A1(new_n1103_), .A2(new_n1732_), .ZN(new_n3512_));
  NOR3_X1    g03256(.A1(new_n3512_), .A2(\a[17] ), .A3(new_n3421_), .ZN(new_n3513_));
  NOR2_X1    g03257(.A1(new_n3511_), .A2(new_n3513_), .ZN(new_n3514_));
  NAND3_X1   g03258(.A1(new_n3508_), .A2(new_n3319_), .A3(new_n3505_), .ZN(new_n3515_));
  OAI21_X1   g03259(.A1(new_n3424_), .A2(new_n3310_), .B(new_n3503_), .ZN(new_n3516_));
  NAND3_X1   g03260(.A1(new_n3516_), .A2(new_n3515_), .A3(new_n3514_), .ZN(new_n3517_));
  NAND2_X1   g03261(.A1(new_n3510_), .A2(new_n3517_), .ZN(new_n3518_));
  NAND3_X1   g03262(.A1(new_n3347_), .A2(new_n3101_), .A3(new_n3342_), .ZN(new_n3519_));
  AOI21_X1   g03263(.A1(new_n3519_), .A2(new_n3343_), .B(new_n3518_), .ZN(new_n3520_));
  AOI21_X1   g03264(.A1(new_n3516_), .A2(new_n3515_), .B(new_n3514_), .ZN(new_n3521_));
  NOR3_X1    g03265(.A1(new_n3509_), .A2(new_n3423_), .A3(new_n3504_), .ZN(new_n3522_));
  NOR2_X1    g03266(.A1(new_n3522_), .A2(new_n3521_), .ZN(new_n3523_));
  OAI21_X1   g03267(.A1(new_n3340_), .A2(new_n3331_), .B(new_n3343_), .ZN(new_n3524_));
  NOR2_X1    g03268(.A1(new_n3524_), .A2(new_n3523_), .ZN(new_n3525_));
  OAI21_X1   g03269(.A1(new_n3525_), .A2(new_n3520_), .B(new_n3419_), .ZN(new_n3526_));
  NOR2_X1    g03270(.A1(new_n3416_), .A2(new_n3418_), .ZN(new_n3527_));
  NOR3_X1    g03271(.A1(new_n2961_), .A2(new_n2944_), .A3(new_n3098_), .ZN(new_n3528_));
  NOR2_X1    g03272(.A1(new_n3339_), .A2(new_n3094_), .ZN(new_n3529_));
  NOR3_X1    g03273(.A1(new_n3529_), .A2(new_n3528_), .A3(new_n3331_), .ZN(new_n3530_));
  OAI21_X1   g03274(.A1(new_n3530_), .A2(new_n3337_), .B(new_n3523_), .ZN(new_n3531_));
  NAND3_X1   g03275(.A1(new_n3519_), .A2(new_n3518_), .A3(new_n3343_), .ZN(new_n3532_));
  NAND3_X1   g03276(.A1(new_n3531_), .A2(new_n3532_), .A3(new_n3527_), .ZN(new_n3533_));
  NAND2_X1   g03277(.A1(new_n3526_), .A2(new_n3533_), .ZN(new_n3534_));
  AOI21_X1   g03278(.A1(new_n3341_), .A2(new_n3348_), .B(new_n3350_), .ZN(new_n3535_));
  INV_X1     g03279(.I(new_n3535_), .ZN(new_n3536_));
  AOI21_X1   g03280(.A1(new_n3355_), .A2(new_n3536_), .B(new_n3534_), .ZN(new_n3537_));
  AOI21_X1   g03281(.A1(new_n3531_), .A2(new_n3532_), .B(new_n3527_), .ZN(new_n3538_));
  NOR3_X1    g03282(.A1(new_n3525_), .A2(new_n3419_), .A3(new_n3520_), .ZN(new_n3539_));
  NOR2_X1    g03283(.A1(new_n3539_), .A2(new_n3538_), .ZN(new_n3540_));
  NOR3_X1    g03284(.A1(new_n3366_), .A2(new_n3540_), .A3(new_n3535_), .ZN(new_n3541_));
  NOR2_X1    g03285(.A1(new_n3541_), .A2(new_n3537_), .ZN(new_n3542_));
  INV_X1     g03286(.I(new_n3542_), .ZN(new_n3543_));
  AOI21_X1   g03287(.A1(new_n3381_), .A2(new_n3363_), .B(new_n3543_), .ZN(new_n3544_));
  NOR3_X1    g03288(.A1(new_n3370_), .A2(new_n3378_), .A3(new_n3542_), .ZN(new_n3545_));
  AOI22_X1   g03289(.A1(new_n518_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n636_), .ZN(new_n3546_));
  OAI21_X1   g03290(.A1(new_n2027_), .A2(new_n917_), .B(new_n3546_), .ZN(new_n3547_));
  AOI21_X1   g03291(.A1(new_n2470_), .A2(new_n618_), .B(new_n3547_), .ZN(new_n3548_));
  NOR2_X1    g03292(.A1(new_n3548_), .A2(new_n488_), .ZN(new_n3549_));
  OAI21_X1   g03293(.A1(new_n2468_), .A2(new_n2467_), .B(\b[23] ), .ZN(new_n3550_));
  NAND3_X1   g03294(.A1(new_n2464_), .A2(new_n2463_), .A3(new_n2465_), .ZN(new_n3551_));
  NAND2_X1   g03295(.A1(new_n3550_), .A2(new_n3551_), .ZN(new_n3552_));
  INV_X1     g03296(.I(new_n3547_), .ZN(new_n3553_));
  OAI21_X1   g03297(.A1(new_n3552_), .A2(new_n624_), .B(new_n3553_), .ZN(new_n3554_));
  NOR2_X1    g03298(.A1(new_n3554_), .A2(\a[8] ), .ZN(new_n3555_));
  OAI22_X1   g03299(.A1(new_n713_), .A2(new_n1860_), .B1(new_n1859_), .B2(new_n717_), .ZN(new_n3556_));
  AOI21_X1   g03300(.A1(\b[18] ), .A2(new_n1126_), .B(new_n3556_), .ZN(new_n3557_));
  OAI21_X1   g03301(.A1(new_n1871_), .A2(new_n986_), .B(new_n3557_), .ZN(new_n3558_));
  XOR2_X1    g03302(.A1(new_n3558_), .A2(\a[11] ), .Z(new_n3559_));
  INV_X1     g03303(.I(new_n3559_), .ZN(new_n3560_));
  OAI21_X1   g03304(.A1(new_n3549_), .A2(new_n3555_), .B(new_n3560_), .ZN(new_n3561_));
  NAND2_X1   g03305(.A1(new_n3554_), .A2(\a[8] ), .ZN(new_n3562_));
  NAND2_X1   g03306(.A1(new_n3548_), .A2(new_n488_), .ZN(new_n3563_));
  NAND3_X1   g03307(.A1(new_n3563_), .A2(new_n3562_), .A3(new_n3559_), .ZN(new_n3564_));
  NAND2_X1   g03308(.A1(new_n3561_), .A2(new_n3564_), .ZN(new_n3565_));
  NOR3_X1    g03309(.A1(new_n3544_), .A2(new_n3545_), .A3(new_n3565_), .ZN(new_n3566_));
  OAI21_X1   g03310(.A1(new_n3370_), .A2(new_n3378_), .B(new_n3542_), .ZN(new_n3567_));
  NAND3_X1   g03311(.A1(new_n3381_), .A2(new_n3363_), .A3(new_n3543_), .ZN(new_n3568_));
  AOI21_X1   g03312(.A1(new_n3563_), .A2(new_n3562_), .B(new_n3559_), .ZN(new_n3569_));
  NOR3_X1    g03313(.A1(new_n3549_), .A2(new_n3555_), .A3(new_n3560_), .ZN(new_n3570_));
  NOR2_X1    g03314(.A1(new_n3569_), .A2(new_n3570_), .ZN(new_n3571_));
  AOI21_X1   g03315(.A1(new_n3568_), .A2(new_n3567_), .B(new_n3571_), .ZN(new_n3572_));
  NOR2_X1    g03316(.A1(new_n3572_), .A2(new_n3566_), .ZN(new_n3573_));
  NOR3_X1    g03317(.A1(new_n3385_), .A2(new_n3146_), .A3(new_n3386_), .ZN(new_n3574_));
  OAI21_X1   g03318(.A1(new_n3574_), .A2(new_n3387_), .B(new_n3573_), .ZN(new_n3575_));
  NAND3_X1   g03319(.A1(new_n3568_), .A2(new_n3567_), .A3(new_n3571_), .ZN(new_n3576_));
  OAI21_X1   g03320(.A1(new_n3544_), .A2(new_n3545_), .B(new_n3565_), .ZN(new_n3577_));
  NAND2_X1   g03321(.A1(new_n3576_), .A2(new_n3577_), .ZN(new_n3578_));
  NAND3_X1   g03322(.A1(new_n3206_), .A2(new_n3142_), .A3(new_n3373_), .ZN(new_n3579_));
  NAND3_X1   g03323(.A1(new_n3579_), .A2(new_n3382_), .A3(new_n3578_), .ZN(new_n3580_));
  AOI21_X1   g03324(.A1(new_n3575_), .A2(new_n3580_), .B(new_n3411_), .ZN(new_n3581_));
  NAND3_X1   g03325(.A1(new_n3575_), .A2(new_n3580_), .A3(new_n3411_), .ZN(new_n3582_));
  INV_X1     g03326(.I(new_n3582_), .ZN(new_n3583_));
  NOR2_X1    g03327(.A1(new_n3583_), .A2(new_n3581_), .ZN(new_n3584_));
  INV_X1     g03328(.I(new_n3584_), .ZN(new_n3585_));
  NOR2_X1    g03329(.A1(new_n284_), .A2(new_n3158_), .ZN(new_n3586_));
  INV_X1     g03330(.I(new_n3586_), .ZN(new_n3587_));
  AOI22_X1   g03331(.A1(new_n267_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n261_), .ZN(new_n3588_));
  AOI21_X1   g03332(.A1(new_n3191_), .A2(\b[28] ), .B(new_n3158_), .ZN(new_n3589_));
  NOR2_X1    g03333(.A1(new_n3191_), .A2(\b[28] ), .ZN(new_n3590_));
  NOR2_X1    g03334(.A1(new_n3191_), .A2(\b[29] ), .ZN(new_n3591_));
  INV_X1     g03335(.I(\b[29] ), .ZN(new_n3592_));
  AOI21_X1   g03336(.A1(new_n3189_), .A2(new_n3190_), .B(new_n3592_), .ZN(new_n3593_));
  OAI22_X1   g03337(.A1(new_n3589_), .A2(new_n3590_), .B1(new_n3591_), .B2(new_n3593_), .ZN(new_n3594_));
  NOR4_X1    g03338(.A1(new_n3589_), .A2(new_n3590_), .A3(new_n3591_), .A4(new_n3593_), .ZN(new_n3595_));
  INV_X1     g03339(.I(new_n3595_), .ZN(new_n3596_));
  NAND3_X1   g03340(.A1(new_n3596_), .A2(new_n265_), .A3(new_n3594_), .ZN(new_n3597_));
  NAND3_X1   g03341(.A1(new_n3597_), .A2(new_n3587_), .A3(new_n3588_), .ZN(new_n3598_));
  XOR2_X1    g03342(.A1(new_n3598_), .A2(new_n270_), .Z(new_n3599_));
  NAND2_X1   g03343(.A1(new_n3599_), .A2(new_n3585_), .ZN(new_n3600_));
  XOR2_X1    g03344(.A1(new_n3598_), .A2(\a[2] ), .Z(new_n3601_));
  NAND2_X1   g03345(.A1(new_n3601_), .A2(new_n3584_), .ZN(new_n3602_));
  NAND3_X1   g03346(.A1(new_n3600_), .A2(new_n3602_), .A3(new_n3406_), .ZN(new_n3603_));
  NAND3_X1   g03347(.A1(new_n3392_), .A2(new_n3391_), .A3(new_n3393_), .ZN(new_n3604_));
  OAI21_X1   g03348(.A1(new_n3384_), .A2(new_n3389_), .B(new_n3204_), .ZN(new_n3605_));
  NAND2_X1   g03349(.A1(new_n3604_), .A2(new_n3605_), .ZN(new_n3606_));
  AOI21_X1   g03350(.A1(new_n3606_), .A2(new_n3199_), .B(new_n3404_), .ZN(new_n3607_));
  NOR2_X1    g03351(.A1(new_n3601_), .A2(new_n3584_), .ZN(new_n3608_));
  NOR2_X1    g03352(.A1(new_n3599_), .A2(new_n3585_), .ZN(new_n3609_));
  OAI21_X1   g03353(.A1(new_n3609_), .A2(new_n3608_), .B(new_n3607_), .ZN(new_n3610_));
  NAND2_X1   g03354(.A1(new_n3610_), .A2(new_n3603_), .ZN(new_n3611_));
  INV_X1     g03355(.I(new_n3611_), .ZN(new_n3612_));
  NAND3_X1   g03356(.A1(new_n3183_), .A2(new_n3181_), .A3(new_n3399_), .ZN(new_n3613_));
  NAND2_X1   g03357(.A1(new_n3613_), .A2(new_n3400_), .ZN(new_n3614_));
  XOR2_X1    g03358(.A1(new_n3614_), .A2(new_n3612_), .Z(\f[29] ));
  INV_X1     g03359(.I(new_n3400_), .ZN(new_n3616_));
  AOI21_X1   g03360(.A1(new_n3177_), .A2(new_n3167_), .B(new_n3157_), .ZN(new_n3617_));
  NOR3_X1    g03361(.A1(new_n3617_), .A2(new_n3178_), .A3(new_n3398_), .ZN(new_n3618_));
  OAI21_X1   g03362(.A1(new_n3618_), .A2(new_n3616_), .B(new_n3612_), .ZN(new_n3619_));
  NOR2_X1    g03363(.A1(new_n3584_), .A2(new_n3607_), .ZN(new_n3620_));
  NAND2_X1   g03364(.A1(new_n3584_), .A2(new_n3607_), .ZN(new_n3621_));
  INV_X1     g03365(.I(new_n3621_), .ZN(new_n3622_));
  OAI21_X1   g03366(.A1(new_n3622_), .A2(new_n3620_), .B(new_n3601_), .ZN(new_n3623_));
  INV_X1     g03367(.I(\b[30] ), .ZN(new_n3624_));
  OAI22_X1   g03368(.A1(new_n277_), .A2(new_n3624_), .B1(new_n3592_), .B2(new_n262_), .ZN(new_n3625_));
  AOI21_X1   g03369(.A1(\b[28] ), .A2(new_n283_), .B(new_n3625_), .ZN(new_n3626_));
  OAI21_X1   g03370(.A1(new_n3591_), .A2(new_n3185_), .B(new_n3158_), .ZN(new_n3627_));
  OAI21_X1   g03371(.A1(new_n3192_), .A2(new_n3592_), .B(new_n3185_), .ZN(new_n3628_));
  XNOR2_X1   g03372(.A1(\b[29] ), .A2(\b[30] ), .ZN(new_n3629_));
  AOI21_X1   g03373(.A1(new_n3627_), .A2(new_n3628_), .B(new_n3629_), .ZN(new_n3630_));
  NAND2_X1   g03374(.A1(new_n3627_), .A2(new_n3628_), .ZN(new_n3631_));
  XOR2_X1    g03375(.A1(\b[29] ), .A2(\b[30] ), .Z(new_n3632_));
  NOR2_X1    g03376(.A1(new_n3631_), .A2(new_n3632_), .ZN(new_n3633_));
  NOR2_X1    g03377(.A1(new_n3633_), .A2(new_n3630_), .ZN(new_n3634_));
  OAI21_X1   g03378(.A1(new_n3634_), .A2(new_n279_), .B(new_n3626_), .ZN(new_n3635_));
  XOR2_X1    g03379(.A1(new_n3635_), .A2(\a[2] ), .Z(new_n3636_));
  INV_X1     g03380(.I(new_n3636_), .ZN(new_n3637_));
  OAI22_X1   g03381(.A1(new_n321_), .A2(new_n3158_), .B1(new_n325_), .B2(new_n3006_), .ZN(new_n3638_));
  AOI21_X1   g03382(.A1(\b[25] ), .A2(new_n602_), .B(new_n3638_), .ZN(new_n3639_));
  OAI21_X1   g03383(.A1(new_n3165_), .A2(new_n318_), .B(new_n3639_), .ZN(new_n3640_));
  XOR2_X1    g03384(.A1(new_n3640_), .A2(\a[5] ), .Z(new_n3641_));
  OAI21_X1   g03385(.A1(new_n3441_), .A2(new_n3486_), .B(new_n3464_), .ZN(new_n3642_));
  OAI22_X1   g03386(.A1(new_n2703_), .A2(new_n438_), .B1(new_n377_), .B2(new_n2708_), .ZN(new_n3643_));
  AOI21_X1   g03387(.A1(\b[4] ), .A2(new_n2906_), .B(new_n3643_), .ZN(new_n3644_));
  OAI21_X1   g03388(.A1(new_n450_), .A2(new_n2711_), .B(new_n3644_), .ZN(new_n3645_));
  XOR2_X1    g03389(.A1(new_n3645_), .A2(\a[26] ), .Z(new_n3646_));
  NAND2_X1   g03390(.A1(new_n3456_), .A2(\b[1] ), .ZN(new_n3647_));
  AOI22_X1   g03391(.A1(new_n3267_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n3270_), .ZN(new_n3648_));
  NAND2_X1   g03392(.A1(new_n299_), .A2(new_n3273_), .ZN(new_n3649_));
  NAND3_X1   g03393(.A1(new_n3649_), .A2(new_n3648_), .A3(new_n3647_), .ZN(new_n3650_));
  NAND2_X1   g03394(.A1(new_n3650_), .A2(\a[29] ), .ZN(new_n3651_));
  NAND4_X1   g03395(.A1(new_n3649_), .A2(new_n3648_), .A3(new_n3264_), .A4(new_n3647_), .ZN(new_n3652_));
  XNOR2_X1   g03396(.A1(\a[29] ), .A2(\a[30] ), .ZN(new_n3653_));
  NOR2_X1    g03397(.A1(new_n3653_), .A2(new_n258_), .ZN(new_n3654_));
  INV_X1     g03398(.I(new_n3654_), .ZN(new_n3655_));
  AOI21_X1   g03399(.A1(new_n3651_), .A2(new_n3652_), .B(new_n3655_), .ZN(new_n3656_));
  NAND3_X1   g03400(.A1(new_n3651_), .A2(new_n3652_), .A3(new_n3655_), .ZN(new_n3657_));
  INV_X1     g03401(.I(new_n3657_), .ZN(new_n3658_));
  OAI21_X1   g03402(.A1(new_n3658_), .A2(new_n3656_), .B(new_n3478_), .ZN(new_n3659_));
  INV_X1     g03403(.I(new_n3656_), .ZN(new_n3660_));
  NAND3_X1   g03404(.A1(new_n3660_), .A2(new_n3462_), .A3(new_n3657_), .ZN(new_n3661_));
  NAND3_X1   g03405(.A1(new_n3659_), .A2(new_n3661_), .A3(new_n3646_), .ZN(new_n3662_));
  XOR2_X1    g03406(.A1(new_n3645_), .A2(new_n2714_), .Z(new_n3663_));
  AOI21_X1   g03407(.A1(new_n3660_), .A2(new_n3657_), .B(new_n3462_), .ZN(new_n3664_));
  NOR3_X1    g03408(.A1(new_n3658_), .A2(new_n3478_), .A3(new_n3656_), .ZN(new_n3665_));
  OAI21_X1   g03409(.A1(new_n3665_), .A2(new_n3664_), .B(new_n3663_), .ZN(new_n3666_));
  NAND2_X1   g03410(.A1(new_n3666_), .A2(new_n3662_), .ZN(new_n3667_));
  NAND2_X1   g03411(.A1(new_n3642_), .A2(new_n3667_), .ZN(new_n3668_));
  AOI21_X1   g03412(.A1(new_n3445_), .A2(new_n3480_), .B(new_n3485_), .ZN(new_n3669_));
  NOR3_X1    g03413(.A1(new_n3665_), .A2(new_n3664_), .A3(new_n3663_), .ZN(new_n3670_));
  AOI21_X1   g03414(.A1(new_n3659_), .A2(new_n3661_), .B(new_n3646_), .ZN(new_n3671_));
  NOR2_X1    g03415(.A1(new_n3670_), .A2(new_n3671_), .ZN(new_n3672_));
  NAND2_X1   g03416(.A1(new_n3669_), .A2(new_n3672_), .ZN(new_n3673_));
  NAND2_X1   g03417(.A1(new_n3673_), .A2(new_n3668_), .ZN(new_n3674_));
  INV_X1     g03418(.I(new_n3674_), .ZN(new_n3675_));
  AOI22_X1   g03419(.A1(new_n2202_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n2205_), .ZN(new_n3676_));
  OAI21_X1   g03420(.A1(new_n471_), .A2(new_n2370_), .B(new_n3676_), .ZN(new_n3677_));
  AOI21_X1   g03421(.A1(new_n676_), .A2(new_n2208_), .B(new_n3677_), .ZN(new_n3678_));
  XOR2_X1    g03422(.A1(new_n3678_), .A2(new_n2200_), .Z(new_n3679_));
  NAND2_X1   g03423(.A1(new_n3487_), .A2(new_n3445_), .ZN(new_n3680_));
  NAND2_X1   g03424(.A1(new_n3481_), .A2(new_n3441_), .ZN(new_n3681_));
  NAND4_X1   g03425(.A1(new_n3680_), .A2(new_n3681_), .A3(new_n3443_), .A4(new_n3444_), .ZN(new_n3682_));
  OAI21_X1   g03426(.A1(new_n3495_), .A2(new_n3492_), .B(new_n3682_), .ZN(new_n3683_));
  NAND2_X1   g03427(.A1(new_n3683_), .A2(new_n3679_), .ZN(new_n3684_));
  INV_X1     g03428(.I(new_n3679_), .ZN(new_n3685_));
  NOR2_X1    g03429(.A1(new_n3481_), .A2(new_n3441_), .ZN(new_n3686_));
  NOR2_X1    g03430(.A1(new_n3487_), .A2(new_n3445_), .ZN(new_n3687_));
  NOR4_X1    g03431(.A1(new_n3687_), .A2(new_n3686_), .A3(new_n3438_), .A4(new_n3440_), .ZN(new_n3688_));
  AOI21_X1   g03432(.A1(new_n3489_), .A2(new_n3432_), .B(new_n3688_), .ZN(new_n3689_));
  NAND2_X1   g03433(.A1(new_n3689_), .A2(new_n3685_), .ZN(new_n3690_));
  AND3_X2    g03434(.A1(new_n3690_), .A2(new_n3675_), .A3(new_n3684_), .Z(new_n3691_));
  AOI21_X1   g03435(.A1(new_n3690_), .A2(new_n3684_), .B(new_n3675_), .ZN(new_n3692_));
  NOR2_X1    g03436(.A1(new_n3691_), .A2(new_n3692_), .ZN(new_n3693_));
  INV_X1     g03437(.I(new_n3693_), .ZN(new_n3694_));
  AOI22_X1   g03438(.A1(new_n1738_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n1743_), .ZN(new_n3695_));
  OAI21_X1   g03439(.A1(new_n776_), .A2(new_n1931_), .B(new_n3695_), .ZN(new_n3696_));
  AOI21_X1   g03440(.A1(new_n1194_), .A2(new_n1746_), .B(new_n3696_), .ZN(new_n3697_));
  XOR2_X1    g03441(.A1(new_n3697_), .A2(new_n1736_), .Z(new_n3698_));
  INV_X1     g03442(.I(new_n3698_), .ZN(new_n3699_));
  AOI21_X1   g03443(.A1(new_n3515_), .A2(new_n3497_), .B(new_n3699_), .ZN(new_n3700_));
  NOR3_X1    g03444(.A1(new_n3504_), .A2(new_n3506_), .A3(new_n3698_), .ZN(new_n3701_));
  NOR3_X1    g03445(.A1(new_n3701_), .A2(new_n3700_), .A3(new_n3694_), .ZN(new_n3702_));
  OAI21_X1   g03446(.A1(new_n3504_), .A2(new_n3506_), .B(new_n3698_), .ZN(new_n3703_));
  NAND3_X1   g03447(.A1(new_n3515_), .A2(new_n3497_), .A3(new_n3699_), .ZN(new_n3704_));
  AOI21_X1   g03448(.A1(new_n3703_), .A2(new_n3704_), .B(new_n3693_), .ZN(new_n3705_));
  NOR2_X1    g03449(.A1(new_n3702_), .A2(new_n3705_), .ZN(new_n3706_));
  INV_X1     g03450(.I(new_n3706_), .ZN(new_n3707_));
  OAI22_X1   g03451(.A1(new_n1592_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n1505_), .ZN(new_n3708_));
  AOI21_X1   g03452(.A1(\b[13] ), .A2(new_n1584_), .B(new_n3708_), .ZN(new_n3709_));
  OAI21_X1   g03453(.A1(new_n1275_), .A2(new_n1732_), .B(new_n3709_), .ZN(new_n3710_));
  XOR2_X1    g03454(.A1(new_n3710_), .A2(\a[17] ), .Z(new_n3711_));
  OAI21_X1   g03455(.A1(new_n3520_), .A2(new_n3522_), .B(new_n3711_), .ZN(new_n3712_));
  INV_X1     g03456(.I(new_n3711_), .ZN(new_n3713_));
  NAND3_X1   g03457(.A1(new_n3531_), .A2(new_n3517_), .A3(new_n3713_), .ZN(new_n3714_));
  NAND2_X1   g03458(.A1(new_n3714_), .A2(new_n3712_), .ZN(new_n3715_));
  XOR2_X1    g03459(.A1(new_n3715_), .A2(new_n3707_), .Z(new_n3716_));
  OAI22_X1   g03460(.A1(new_n993_), .A2(new_n1553_), .B1(new_n1432_), .B2(new_n997_), .ZN(new_n3717_));
  AOI21_X1   g03461(.A1(\b[16] ), .A2(new_n1486_), .B(new_n3717_), .ZN(new_n3718_));
  OAI21_X1   g03462(.A1(new_n1563_), .A2(new_n1323_), .B(new_n3718_), .ZN(new_n3719_));
  XOR2_X1    g03463(.A1(new_n3719_), .A2(\a[14] ), .Z(new_n3720_));
  OAI21_X1   g03464(.A1(new_n3537_), .A2(new_n3539_), .B(new_n3720_), .ZN(new_n3721_));
  OAI21_X1   g03465(.A1(new_n3366_), .A2(new_n3535_), .B(new_n3540_), .ZN(new_n3722_));
  INV_X1     g03466(.I(new_n3720_), .ZN(new_n3723_));
  NAND3_X1   g03467(.A1(new_n3722_), .A2(new_n3533_), .A3(new_n3723_), .ZN(new_n3724_));
  NAND2_X1   g03468(.A1(new_n3724_), .A2(new_n3721_), .ZN(new_n3725_));
  XOR2_X1    g03469(.A1(new_n3725_), .A2(new_n3716_), .Z(new_n3726_));
  INV_X1     g03470(.I(new_n2032_), .ZN(new_n3727_));
  OAI22_X1   g03471(.A1(new_n713_), .A2(new_n2027_), .B1(new_n1860_), .B2(new_n717_), .ZN(new_n3728_));
  AOI21_X1   g03472(.A1(\b[19] ), .A2(new_n1126_), .B(new_n3728_), .ZN(new_n3729_));
  OAI21_X1   g03473(.A1(new_n3727_), .A2(new_n986_), .B(new_n3729_), .ZN(new_n3730_));
  XOR2_X1    g03474(.A1(new_n3730_), .A2(\a[11] ), .Z(new_n3731_));
  INV_X1     g03475(.I(new_n3731_), .ZN(new_n3732_));
  NAND3_X1   g03476(.A1(new_n3355_), .A2(new_n3534_), .A3(new_n3536_), .ZN(new_n3733_));
  NAND3_X1   g03477(.A1(new_n3722_), .A2(new_n3733_), .A3(new_n3559_), .ZN(new_n3734_));
  NOR3_X1    g03478(.A1(new_n3541_), .A2(new_n3537_), .A3(new_n3560_), .ZN(new_n3735_));
  AOI21_X1   g03479(.A1(new_n3722_), .A2(new_n3733_), .B(new_n3559_), .ZN(new_n3736_));
  NOR2_X1    g03480(.A1(new_n3735_), .A2(new_n3736_), .ZN(new_n3737_));
  OAI21_X1   g03481(.A1(new_n3370_), .A2(new_n3378_), .B(new_n3737_), .ZN(new_n3738_));
  AOI21_X1   g03482(.A1(new_n3738_), .A2(new_n3734_), .B(new_n3732_), .ZN(new_n3739_));
  OAI21_X1   g03483(.A1(new_n3541_), .A2(new_n3537_), .B(new_n3560_), .ZN(new_n3740_));
  NAND2_X1   g03484(.A1(new_n3740_), .A2(new_n3734_), .ZN(new_n3741_));
  AOI21_X1   g03485(.A1(new_n3381_), .A2(new_n3363_), .B(new_n3741_), .ZN(new_n3742_));
  NOR3_X1    g03486(.A1(new_n3742_), .A2(new_n3731_), .A3(new_n3735_), .ZN(new_n3743_));
  NOR3_X1    g03487(.A1(new_n3743_), .A2(new_n3739_), .A3(new_n3726_), .ZN(new_n3744_));
  NAND3_X1   g03488(.A1(new_n3714_), .A2(new_n3712_), .A3(new_n3706_), .ZN(new_n3745_));
  NAND2_X1   g03489(.A1(new_n3715_), .A2(new_n3707_), .ZN(new_n3746_));
  NAND2_X1   g03490(.A1(new_n3746_), .A2(new_n3745_), .ZN(new_n3747_));
  NOR2_X1    g03491(.A1(new_n3725_), .A2(new_n3747_), .ZN(new_n3748_));
  AOI21_X1   g03492(.A1(new_n3724_), .A2(new_n3721_), .B(new_n3716_), .ZN(new_n3749_));
  NOR2_X1    g03493(.A1(new_n3748_), .A2(new_n3749_), .ZN(new_n3750_));
  OAI21_X1   g03494(.A1(new_n3742_), .A2(new_n3735_), .B(new_n3731_), .ZN(new_n3751_));
  NAND3_X1   g03495(.A1(new_n3738_), .A2(new_n3732_), .A3(new_n3734_), .ZN(new_n3752_));
  AOI21_X1   g03496(.A1(new_n3751_), .A2(new_n3752_), .B(new_n3750_), .ZN(new_n3753_));
  NOR2_X1    g03497(.A1(new_n3744_), .A2(new_n3753_), .ZN(new_n3754_));
  AOI21_X1   g03498(.A1(new_n3579_), .A2(new_n3382_), .B(new_n3578_), .ZN(new_n3755_));
  AOI22_X1   g03499(.A1(new_n518_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n636_), .ZN(new_n3756_));
  OAI21_X1   g03500(.A1(new_n2142_), .A2(new_n917_), .B(new_n3756_), .ZN(new_n3757_));
  AOI21_X1   g03501(.A1(new_n3033_), .A2(new_n618_), .B(new_n3757_), .ZN(new_n3758_));
  XOR2_X1    g03502(.A1(new_n3758_), .A2(new_n488_), .Z(new_n3759_));
  NOR2_X1    g03503(.A1(new_n3549_), .A2(new_n3555_), .ZN(new_n3760_));
  AOI21_X1   g03504(.A1(new_n3119_), .A2(new_n3130_), .B(new_n3128_), .ZN(new_n3761_));
  AOI21_X1   g03505(.A1(new_n3761_), .A2(new_n3380_), .B(new_n3378_), .ZN(new_n3762_));
  NAND2_X1   g03506(.A1(new_n3762_), .A2(new_n3741_), .ZN(new_n3763_));
  NAND3_X1   g03507(.A1(new_n3763_), .A2(new_n3760_), .A3(new_n3738_), .ZN(new_n3764_));
  INV_X1     g03508(.I(new_n3764_), .ZN(new_n3765_));
  OAI21_X1   g03509(.A1(new_n3755_), .A2(new_n3765_), .B(new_n3759_), .ZN(new_n3766_));
  INV_X1     g03510(.I(new_n3759_), .ZN(new_n3767_));
  NAND3_X1   g03511(.A1(new_n3575_), .A2(new_n3767_), .A3(new_n3764_), .ZN(new_n3768_));
  NAND3_X1   g03512(.A1(new_n3768_), .A2(new_n3766_), .A3(new_n3754_), .ZN(new_n3769_));
  INV_X1     g03513(.I(new_n3754_), .ZN(new_n3770_));
  AOI21_X1   g03514(.A1(new_n3575_), .A2(new_n3764_), .B(new_n3767_), .ZN(new_n3771_));
  NOR3_X1    g03515(.A1(new_n3755_), .A2(new_n3759_), .A3(new_n3765_), .ZN(new_n3772_));
  OAI21_X1   g03516(.A1(new_n3771_), .A2(new_n3772_), .B(new_n3770_), .ZN(new_n3773_));
  AOI21_X1   g03517(.A1(new_n3773_), .A2(new_n3769_), .B(new_n3641_), .ZN(new_n3774_));
  NAND3_X1   g03518(.A1(new_n3773_), .A2(new_n3769_), .A3(new_n3641_), .ZN(new_n3775_));
  INV_X1     g03519(.I(new_n3775_), .ZN(new_n3776_));
  AOI21_X1   g03520(.A1(new_n3607_), .A2(new_n3582_), .B(new_n3581_), .ZN(new_n3777_));
  NOR3_X1    g03521(.A1(new_n3776_), .A2(new_n3774_), .A3(new_n3777_), .ZN(new_n3778_));
  OAI21_X1   g03522(.A1(new_n3776_), .A2(new_n3774_), .B(new_n3777_), .ZN(new_n3779_));
  INV_X1     g03523(.I(new_n3779_), .ZN(new_n3780_));
  NOR3_X1    g03524(.A1(new_n3780_), .A2(new_n3778_), .A3(new_n3637_), .ZN(new_n3781_));
  INV_X1     g03525(.I(new_n3778_), .ZN(new_n3782_));
  AOI21_X1   g03526(.A1(new_n3782_), .A2(new_n3779_), .B(new_n3636_), .ZN(new_n3783_));
  NOR2_X1    g03527(.A1(new_n3783_), .A2(new_n3781_), .ZN(new_n3784_));
  AOI21_X1   g03528(.A1(new_n3619_), .A2(new_n3623_), .B(new_n3784_), .ZN(new_n3785_));
  AOI21_X1   g03529(.A1(new_n3613_), .A2(new_n3400_), .B(new_n3611_), .ZN(new_n3786_));
  INV_X1     g03530(.I(new_n3623_), .ZN(new_n3787_));
  NOR4_X1    g03531(.A1(new_n3786_), .A2(new_n3787_), .A3(new_n3781_), .A4(new_n3783_), .ZN(new_n3788_));
  NOR2_X1    g03532(.A1(new_n3785_), .A2(new_n3788_), .ZN(\f[30] ));
  NAND2_X1   g03533(.A1(new_n283_), .A2(\b[29] ), .ZN(new_n3790_));
  AOI22_X1   g03534(.A1(new_n267_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n261_), .ZN(new_n3791_));
  NAND2_X1   g03535(.A1(new_n3631_), .A2(new_n3592_), .ZN(new_n3792_));
  NOR2_X1    g03536(.A1(new_n3631_), .A2(new_n3592_), .ZN(new_n3793_));
  NAND2_X1   g03537(.A1(new_n3793_), .A2(new_n3624_), .ZN(new_n3794_));
  OAI21_X1   g03538(.A1(new_n3624_), .A2(new_n3792_), .B(new_n3794_), .ZN(new_n3795_));
  XOR2_X1    g03539(.A1(new_n3795_), .A2(\b[31] ), .Z(new_n3796_));
  NAND2_X1   g03540(.A1(new_n3796_), .A2(new_n265_), .ZN(new_n3797_));
  NAND3_X1   g03541(.A1(new_n3797_), .A2(new_n3790_), .A3(new_n3791_), .ZN(new_n3798_));
  XOR2_X1    g03542(.A1(new_n3798_), .A2(\a[2] ), .Z(new_n3799_));
  INV_X1     g03543(.I(new_n3799_), .ZN(new_n3800_));
  OAI22_X1   g03544(.A1(new_n3786_), .A2(new_n3787_), .B1(new_n3781_), .B2(new_n3783_), .ZN(new_n3801_));
  AOI21_X1   g03545(.A1(new_n3782_), .A2(new_n3779_), .B(new_n3637_), .ZN(new_n3802_));
  INV_X1     g03546(.I(new_n3802_), .ZN(new_n3803_));
  INV_X1     g03547(.I(new_n3581_), .ZN(new_n3804_));
  OAI21_X1   g03548(.A1(new_n3406_), .A2(new_n3583_), .B(new_n3804_), .ZN(new_n3805_));
  OAI21_X1   g03549(.A1(new_n3805_), .A2(new_n3774_), .B(new_n3775_), .ZN(new_n3806_));
  INV_X1     g03550(.I(new_n3196_), .ZN(new_n3807_));
  AOI22_X1   g03551(.A1(new_n800_), .A2(\b[27] ), .B1(\b[28] ), .B2(new_n333_), .ZN(new_n3808_));
  OAI21_X1   g03552(.A1(new_n3006_), .A2(new_n392_), .B(new_n3808_), .ZN(new_n3809_));
  AOI21_X1   g03553(.A1(new_n3807_), .A2(new_n330_), .B(new_n3809_), .ZN(new_n3810_));
  XOR2_X1    g03554(.A1(new_n3810_), .A2(new_n312_), .Z(new_n3811_));
  NOR2_X1    g03555(.A1(new_n3771_), .A2(new_n3754_), .ZN(new_n3812_));
  AOI22_X1   g03556(.A1(new_n518_), .A2(\b[25] ), .B1(\b[24] ), .B2(new_n636_), .ZN(new_n3813_));
  OAI21_X1   g03557(.A1(new_n2463_), .A2(new_n917_), .B(new_n3813_), .ZN(new_n3814_));
  INV_X1     g03558(.I(new_n3814_), .ZN(new_n3815_));
  XNOR2_X1   g03559(.A1(new_n2651_), .A2(new_n2654_), .ZN(new_n3816_));
  NAND2_X1   g03560(.A1(new_n3816_), .A2(new_n618_), .ZN(new_n3817_));
  AOI21_X1   g03561(.A1(new_n3817_), .A2(new_n3815_), .B(new_n488_), .ZN(new_n3818_));
  OAI21_X1   g03562(.A1(new_n2655_), .A2(new_n624_), .B(new_n3815_), .ZN(new_n3819_));
  NOR2_X1    g03563(.A1(new_n3819_), .A2(\a[8] ), .ZN(new_n3820_));
  NOR2_X1    g03564(.A1(new_n3818_), .A2(new_n3820_), .ZN(new_n3821_));
  OAI21_X1   g03565(.A1(new_n3118_), .A2(new_n3126_), .B(new_n3131_), .ZN(new_n3822_));
  OAI21_X1   g03566(.A1(new_n3822_), .A2(new_n3369_), .B(new_n3363_), .ZN(new_n3823_));
  AOI21_X1   g03567(.A1(new_n3823_), .A2(new_n3737_), .B(new_n3735_), .ZN(new_n3824_));
  OAI21_X1   g03568(.A1(new_n3824_), .A2(new_n3732_), .B(new_n3726_), .ZN(new_n3825_));
  OAI22_X1   g03569(.A1(new_n713_), .A2(new_n2142_), .B1(new_n2027_), .B2(new_n717_), .ZN(new_n3826_));
  AOI21_X1   g03570(.A1(\b[20] ), .A2(new_n1126_), .B(new_n3826_), .ZN(new_n3827_));
  OAI21_X1   g03571(.A1(new_n2153_), .A2(new_n986_), .B(new_n3827_), .ZN(new_n3828_));
  XOR2_X1    g03572(.A1(new_n3828_), .A2(\a[11] ), .Z(new_n3829_));
  NOR3_X1    g03573(.A1(new_n3537_), .A2(new_n3539_), .A3(new_n3720_), .ZN(new_n3830_));
  AOI21_X1   g03574(.A1(new_n3105_), .A2(new_n3115_), .B(new_n3112_), .ZN(new_n3831_));
  AOI21_X1   g03575(.A1(new_n3831_), .A2(new_n3354_), .B(new_n3535_), .ZN(new_n3832_));
  OAI21_X1   g03576(.A1(new_n3832_), .A2(new_n3534_), .B(new_n3533_), .ZN(new_n3833_));
  AOI21_X1   g03577(.A1(new_n3833_), .A2(new_n3720_), .B(new_n3716_), .ZN(new_n3834_));
  AOI22_X1   g03578(.A1(new_n1006_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n1009_), .ZN(new_n3835_));
  OAI21_X1   g03579(.A1(new_n1432_), .A2(new_n1481_), .B(new_n3835_), .ZN(new_n3836_));
  INV_X1     g03580(.I(new_n3836_), .ZN(new_n3837_));
  NAND2_X1   g03581(.A1(new_n1695_), .A2(new_n1013_), .ZN(new_n3838_));
  AOI21_X1   g03582(.A1(new_n3838_), .A2(new_n3837_), .B(new_n1002_), .ZN(new_n3839_));
  AND3_X2    g03583(.A1(new_n3838_), .A2(new_n1002_), .A3(new_n3837_), .Z(new_n3840_));
  NOR2_X1    g03584(.A1(new_n3840_), .A2(new_n3839_), .ZN(new_n3841_));
  AOI21_X1   g03585(.A1(new_n3524_), .A2(new_n3523_), .B(new_n3522_), .ZN(new_n3842_));
  OAI21_X1   g03586(.A1(new_n3842_), .A2(new_n3713_), .B(new_n3707_), .ZN(new_n3843_));
  OAI22_X1   g03587(.A1(new_n1592_), .A2(new_n1296_), .B1(new_n1268_), .B2(new_n1505_), .ZN(new_n3844_));
  AOI21_X1   g03588(.A1(\b[14] ), .A2(new_n1584_), .B(new_n3844_), .ZN(new_n3845_));
  OAI21_X1   g03589(.A1(new_n1306_), .A2(new_n1732_), .B(new_n3845_), .ZN(new_n3846_));
  XOR2_X1    g03590(.A1(new_n3846_), .A2(\a[17] ), .Z(new_n3847_));
  OAI21_X1   g03591(.A1(new_n3693_), .A2(new_n3700_), .B(new_n3704_), .ZN(new_n3848_));
  NOR2_X1    g03592(.A1(new_n3683_), .A2(new_n3679_), .ZN(new_n3849_));
  AOI21_X1   g03593(.A1(new_n3683_), .A2(new_n3679_), .B(new_n3675_), .ZN(new_n3850_));
  AOI21_X1   g03594(.A1(new_n3659_), .A2(new_n3661_), .B(new_n3663_), .ZN(new_n3851_));
  AOI21_X1   g03595(.A1(new_n3642_), .A2(new_n3667_), .B(new_n3851_), .ZN(new_n3852_));
  NAND2_X1   g03596(.A1(new_n3651_), .A2(new_n3652_), .ZN(new_n3853_));
  INV_X1     g03597(.I(new_n3853_), .ZN(new_n3854_));
  NAND2_X1   g03598(.A1(new_n3478_), .A2(new_n3655_), .ZN(new_n3855_));
  NOR2_X1    g03599(.A1(new_n3478_), .A2(new_n3655_), .ZN(new_n3856_));
  AOI21_X1   g03600(.A1(new_n3854_), .A2(new_n3855_), .B(new_n3856_), .ZN(new_n3857_));
  AOI22_X1   g03601(.A1(new_n3267_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n3270_), .ZN(new_n3858_));
  NAND2_X1   g03602(.A1(new_n3456_), .A2(\b[2] ), .ZN(new_n3859_));
  NAND2_X1   g03603(.A1(new_n1725_), .A2(new_n3273_), .ZN(new_n3860_));
  NAND3_X1   g03604(.A1(new_n3860_), .A2(new_n3858_), .A3(new_n3859_), .ZN(new_n3861_));
  XOR2_X1    g03605(.A1(new_n3861_), .A2(\a[29] ), .Z(new_n3862_));
  XOR2_X1    g03606(.A1(\a[31] ), .A2(\a[32] ), .Z(new_n3863_));
  NOR2_X1    g03607(.A1(new_n3653_), .A2(new_n3863_), .ZN(new_n3864_));
  INV_X1     g03608(.I(\a[30] ), .ZN(new_n3865_));
  NAND3_X1   g03609(.A1(new_n3264_), .A2(new_n3865_), .A3(\a[31] ), .ZN(new_n3866_));
  INV_X1     g03610(.I(\a[31] ), .ZN(new_n3867_));
  NAND3_X1   g03611(.A1(new_n3867_), .A2(\a[29] ), .A3(\a[30] ), .ZN(new_n3868_));
  NAND2_X1   g03612(.A1(new_n3866_), .A2(new_n3868_), .ZN(new_n3869_));
  AOI22_X1   g03613(.A1(new_n3864_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n3869_), .ZN(new_n3870_));
  XNOR2_X1   g03614(.A1(\a[31] ), .A2(\a[32] ), .ZN(new_n3871_));
  NOR2_X1    g03615(.A1(new_n3653_), .A2(new_n3871_), .ZN(new_n3872_));
  NAND2_X1   g03616(.A1(new_n3872_), .A2(new_n263_), .ZN(new_n3873_));
  NAND2_X1   g03617(.A1(new_n3870_), .A2(new_n3873_), .ZN(new_n3874_));
  NAND2_X1   g03618(.A1(new_n3874_), .A2(\a[32] ), .ZN(new_n3875_));
  INV_X1     g03619(.I(\a[32] ), .ZN(new_n3876_));
  NAND3_X1   g03620(.A1(new_n3870_), .A2(new_n3873_), .A3(new_n3876_), .ZN(new_n3877_));
  NAND2_X1   g03621(.A1(new_n3655_), .A2(\a[32] ), .ZN(new_n3878_));
  NAND3_X1   g03622(.A1(new_n3875_), .A2(new_n3877_), .A3(new_n3878_), .ZN(new_n3879_));
  NAND3_X1   g03623(.A1(new_n3874_), .A2(\a[32] ), .A3(new_n3655_), .ZN(new_n3880_));
  NAND2_X1   g03624(.A1(new_n3879_), .A2(new_n3880_), .ZN(new_n3881_));
  NAND2_X1   g03625(.A1(new_n3881_), .A2(new_n3862_), .ZN(new_n3882_));
  XOR2_X1    g03626(.A1(new_n3861_), .A2(new_n3264_), .Z(new_n3883_));
  NAND3_X1   g03627(.A1(new_n3883_), .A2(new_n3879_), .A3(new_n3880_), .ZN(new_n3884_));
  AOI21_X1   g03628(.A1(new_n3882_), .A2(new_n3884_), .B(new_n3857_), .ZN(new_n3885_));
  NOR2_X1    g03629(.A1(new_n3462_), .A2(new_n3654_), .ZN(new_n3886_));
  NAND2_X1   g03630(.A1(new_n3462_), .A2(new_n3654_), .ZN(new_n3887_));
  OAI21_X1   g03631(.A1(new_n3853_), .A2(new_n3886_), .B(new_n3887_), .ZN(new_n3888_));
  AOI21_X1   g03632(.A1(new_n3879_), .A2(new_n3880_), .B(new_n3883_), .ZN(new_n3889_));
  NOR2_X1    g03633(.A1(new_n3881_), .A2(new_n3862_), .ZN(new_n3890_));
  NOR3_X1    g03634(.A1(new_n3889_), .A2(new_n3888_), .A3(new_n3890_), .ZN(new_n3891_));
  NOR2_X1    g03635(.A1(new_n3885_), .A2(new_n3891_), .ZN(new_n3892_));
  OAI22_X1   g03636(.A1(new_n2703_), .A2(new_n471_), .B1(new_n438_), .B2(new_n2708_), .ZN(new_n3893_));
  AOI21_X1   g03637(.A1(\b[5] ), .A2(new_n2906_), .B(new_n3893_), .ZN(new_n3894_));
  OAI21_X1   g03638(.A1(new_n485_), .A2(new_n2711_), .B(new_n3894_), .ZN(new_n3895_));
  XOR2_X1    g03639(.A1(new_n3895_), .A2(\a[26] ), .Z(new_n3896_));
  INV_X1     g03640(.I(new_n3896_), .ZN(new_n3897_));
  NAND2_X1   g03641(.A1(new_n3897_), .A2(new_n3892_), .ZN(new_n3898_));
  OR2_X2     g03642(.A1(new_n3885_), .A2(new_n3891_), .Z(new_n3899_));
  NAND2_X1   g03643(.A1(new_n3899_), .A2(new_n3896_), .ZN(new_n3900_));
  AOI21_X1   g03644(.A1(new_n3898_), .A2(new_n3900_), .B(new_n3852_), .ZN(new_n3901_));
  INV_X1     g03645(.I(new_n3851_), .ZN(new_n3902_));
  OAI21_X1   g03646(.A1(new_n3669_), .A2(new_n3672_), .B(new_n3902_), .ZN(new_n3903_));
  NOR2_X1    g03647(.A1(new_n3899_), .A2(new_n3896_), .ZN(new_n3904_));
  NOR2_X1    g03648(.A1(new_n3897_), .A2(new_n3892_), .ZN(new_n3905_));
  NOR3_X1    g03649(.A1(new_n3904_), .A2(new_n3903_), .A3(new_n3905_), .ZN(new_n3906_));
  AOI22_X1   g03650(.A1(new_n2202_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n2205_), .ZN(new_n3907_));
  OAI21_X1   g03651(.A1(new_n577_), .A2(new_n2370_), .B(new_n3907_), .ZN(new_n3908_));
  AOI21_X1   g03652(.A1(new_n1059_), .A2(new_n2208_), .B(new_n3908_), .ZN(new_n3909_));
  XOR2_X1    g03653(.A1(new_n3909_), .A2(new_n2200_), .Z(new_n3910_));
  NOR3_X1    g03654(.A1(new_n3901_), .A2(new_n3906_), .A3(new_n3910_), .ZN(new_n3911_));
  OAI21_X1   g03655(.A1(new_n3904_), .A2(new_n3905_), .B(new_n3903_), .ZN(new_n3912_));
  NAND3_X1   g03656(.A1(new_n3900_), .A2(new_n3852_), .A3(new_n3898_), .ZN(new_n3913_));
  XOR2_X1    g03657(.A1(new_n3909_), .A2(\a[23] ), .Z(new_n3914_));
  AOI21_X1   g03658(.A1(new_n3912_), .A2(new_n3913_), .B(new_n3914_), .ZN(new_n3915_));
  NOR2_X1    g03659(.A1(new_n3911_), .A2(new_n3915_), .ZN(new_n3916_));
  NOR3_X1    g03660(.A1(new_n3916_), .A2(new_n3849_), .A3(new_n3850_), .ZN(new_n3917_));
  INV_X1     g03661(.I(new_n3917_), .ZN(new_n3918_));
  OAI21_X1   g03662(.A1(new_n3849_), .A2(new_n3850_), .B(new_n3916_), .ZN(new_n3919_));
  AOI22_X1   g03663(.A1(new_n1738_), .A2(\b[13] ), .B1(\b[12] ), .B2(new_n1743_), .ZN(new_n3920_));
  OAI21_X1   g03664(.A1(new_n852_), .A2(new_n1931_), .B(new_n3920_), .ZN(new_n3921_));
  INV_X1     g03665(.I(new_n3921_), .ZN(new_n3922_));
  OAI21_X1   g03666(.A1(new_n1082_), .A2(new_n1757_), .B(new_n3922_), .ZN(new_n3923_));
  NAND2_X1   g03667(.A1(new_n3923_), .A2(\a[20] ), .ZN(new_n3924_));
  AOI21_X1   g03668(.A1(new_n1818_), .A2(new_n1746_), .B(new_n3921_), .ZN(new_n3925_));
  NAND2_X1   g03669(.A1(new_n3925_), .A2(new_n1736_), .ZN(new_n3926_));
  NAND2_X1   g03670(.A1(new_n3926_), .A2(new_n3924_), .ZN(new_n3927_));
  AOI21_X1   g03671(.A1(new_n3918_), .A2(new_n3919_), .B(new_n3927_), .ZN(new_n3928_));
  NOR2_X1    g03672(.A1(new_n3850_), .A2(new_n3849_), .ZN(new_n3929_));
  NOR3_X1    g03673(.A1(new_n3929_), .A2(new_n3911_), .A3(new_n3915_), .ZN(new_n3930_));
  XOR2_X1    g03674(.A1(new_n3923_), .A2(\a[20] ), .Z(new_n3931_));
  NOR3_X1    g03675(.A1(new_n3931_), .A2(new_n3930_), .A3(new_n3917_), .ZN(new_n3932_));
  NOR2_X1    g03676(.A1(new_n3928_), .A2(new_n3932_), .ZN(new_n3933_));
  NAND2_X1   g03677(.A1(new_n3848_), .A2(new_n3933_), .ZN(new_n3934_));
  NAND2_X1   g03678(.A1(new_n3703_), .A2(new_n3694_), .ZN(new_n3935_));
  OAI21_X1   g03679(.A1(new_n3917_), .A2(new_n3930_), .B(new_n3931_), .ZN(new_n3936_));
  NAND3_X1   g03680(.A1(new_n3918_), .A2(new_n3927_), .A3(new_n3919_), .ZN(new_n3937_));
  NAND2_X1   g03681(.A1(new_n3936_), .A2(new_n3937_), .ZN(new_n3938_));
  NAND3_X1   g03682(.A1(new_n3938_), .A2(new_n3935_), .A3(new_n3704_), .ZN(new_n3939_));
  NAND3_X1   g03683(.A1(new_n3939_), .A2(new_n3934_), .A3(new_n3847_), .ZN(new_n3940_));
  INV_X1     g03684(.I(new_n3847_), .ZN(new_n3941_));
  AOI21_X1   g03685(.A1(new_n3694_), .A2(new_n3703_), .B(new_n3701_), .ZN(new_n3942_));
  NOR2_X1    g03686(.A1(new_n3942_), .A2(new_n3938_), .ZN(new_n3943_));
  NOR2_X1    g03687(.A1(new_n3848_), .A2(new_n3933_), .ZN(new_n3944_));
  OAI21_X1   g03688(.A1(new_n3943_), .A2(new_n3944_), .B(new_n3941_), .ZN(new_n3945_));
  NAND2_X1   g03689(.A1(new_n3945_), .A2(new_n3940_), .ZN(new_n3946_));
  NAND3_X1   g03690(.A1(new_n3946_), .A2(new_n3843_), .A3(new_n3714_), .ZN(new_n3947_));
  NOR3_X1    g03691(.A1(new_n3520_), .A2(new_n3522_), .A3(new_n3711_), .ZN(new_n3948_));
  AOI21_X1   g03692(.A1(new_n3093_), .A2(new_n3099_), .B(new_n3528_), .ZN(new_n3949_));
  AOI21_X1   g03693(.A1(new_n3949_), .A2(new_n3342_), .B(new_n3337_), .ZN(new_n3950_));
  OAI21_X1   g03694(.A1(new_n3950_), .A2(new_n3518_), .B(new_n3517_), .ZN(new_n3951_));
  AOI21_X1   g03695(.A1(new_n3951_), .A2(new_n3711_), .B(new_n3706_), .ZN(new_n3952_));
  NOR3_X1    g03696(.A1(new_n3943_), .A2(new_n3944_), .A3(new_n3941_), .ZN(new_n3953_));
  AOI21_X1   g03697(.A1(new_n3939_), .A2(new_n3934_), .B(new_n3847_), .ZN(new_n3954_));
  NOR2_X1    g03698(.A1(new_n3953_), .A2(new_n3954_), .ZN(new_n3955_));
  OAI21_X1   g03699(.A1(new_n3952_), .A2(new_n3948_), .B(new_n3955_), .ZN(new_n3956_));
  NAND3_X1   g03700(.A1(new_n3956_), .A2(new_n3947_), .A3(new_n3841_), .ZN(new_n3957_));
  INV_X1     g03701(.I(new_n3841_), .ZN(new_n3958_));
  NOR3_X1    g03702(.A1(new_n3955_), .A2(new_n3952_), .A3(new_n3948_), .ZN(new_n3959_));
  AOI21_X1   g03703(.A1(new_n3843_), .A2(new_n3714_), .B(new_n3946_), .ZN(new_n3960_));
  OAI21_X1   g03704(.A1(new_n3959_), .A2(new_n3960_), .B(new_n3958_), .ZN(new_n3961_));
  NAND2_X1   g03705(.A1(new_n3961_), .A2(new_n3957_), .ZN(new_n3962_));
  NOR3_X1    g03706(.A1(new_n3834_), .A2(new_n3830_), .A3(new_n3962_), .ZN(new_n3963_));
  OAI21_X1   g03707(.A1(new_n3114_), .A2(new_n3111_), .B(new_n3116_), .ZN(new_n3964_));
  OAI21_X1   g03708(.A1(new_n3964_), .A2(new_n3361_), .B(new_n3536_), .ZN(new_n3965_));
  AOI21_X1   g03709(.A1(new_n3965_), .A2(new_n3540_), .B(new_n3539_), .ZN(new_n3966_));
  OAI21_X1   g03710(.A1(new_n3966_), .A2(new_n3723_), .B(new_n3747_), .ZN(new_n3967_));
  NOR3_X1    g03711(.A1(new_n3958_), .A2(new_n3960_), .A3(new_n3959_), .ZN(new_n3968_));
  AOI21_X1   g03712(.A1(new_n3956_), .A2(new_n3947_), .B(new_n3841_), .ZN(new_n3969_));
  NOR2_X1    g03713(.A1(new_n3968_), .A2(new_n3969_), .ZN(new_n3970_));
  AOI21_X1   g03714(.A1(new_n3967_), .A2(new_n3724_), .B(new_n3970_), .ZN(new_n3971_));
  OAI21_X1   g03715(.A1(new_n3963_), .A2(new_n3971_), .B(new_n3829_), .ZN(new_n3972_));
  INV_X1     g03716(.I(new_n3829_), .ZN(new_n3973_));
  NAND3_X1   g03717(.A1(new_n3967_), .A2(new_n3970_), .A3(new_n3724_), .ZN(new_n3974_));
  OAI21_X1   g03718(.A1(new_n3834_), .A2(new_n3830_), .B(new_n3962_), .ZN(new_n3975_));
  NAND3_X1   g03719(.A1(new_n3975_), .A2(new_n3973_), .A3(new_n3974_), .ZN(new_n3976_));
  NAND2_X1   g03720(.A1(new_n3972_), .A2(new_n3976_), .ZN(new_n3977_));
  NAND3_X1   g03721(.A1(new_n3825_), .A2(new_n3752_), .A3(new_n3977_), .ZN(new_n3978_));
  OAI21_X1   g03722(.A1(new_n3762_), .A2(new_n3741_), .B(new_n3734_), .ZN(new_n3979_));
  AOI21_X1   g03723(.A1(new_n3979_), .A2(new_n3731_), .B(new_n3750_), .ZN(new_n3980_));
  AOI21_X1   g03724(.A1(new_n3975_), .A2(new_n3974_), .B(new_n3973_), .ZN(new_n3981_));
  NOR3_X1    g03725(.A1(new_n3963_), .A2(new_n3971_), .A3(new_n3829_), .ZN(new_n3982_));
  NOR2_X1    g03726(.A1(new_n3982_), .A2(new_n3981_), .ZN(new_n3983_));
  OAI21_X1   g03727(.A1(new_n3980_), .A2(new_n3743_), .B(new_n3983_), .ZN(new_n3984_));
  NAND3_X1   g03728(.A1(new_n3978_), .A2(new_n3984_), .A3(new_n3821_), .ZN(new_n3985_));
  INV_X1     g03729(.I(new_n3821_), .ZN(new_n3986_));
  NOR3_X1    g03730(.A1(new_n3980_), .A2(new_n3983_), .A3(new_n3743_), .ZN(new_n3987_));
  AOI21_X1   g03731(.A1(new_n3825_), .A2(new_n3752_), .B(new_n3977_), .ZN(new_n3988_));
  OAI21_X1   g03732(.A1(new_n3988_), .A2(new_n3987_), .B(new_n3986_), .ZN(new_n3989_));
  NAND2_X1   g03733(.A1(new_n3989_), .A2(new_n3985_), .ZN(new_n3990_));
  NOR3_X1    g03734(.A1(new_n3812_), .A2(new_n3772_), .A3(new_n3990_), .ZN(new_n3991_));
  OAI21_X1   g03735(.A1(new_n3133_), .A2(new_n3145_), .B(new_n3142_), .ZN(new_n3992_));
  OAI21_X1   g03736(.A1(new_n3992_), .A2(new_n3386_), .B(new_n3382_), .ZN(new_n3993_));
  AOI21_X1   g03737(.A1(new_n3993_), .A2(new_n3573_), .B(new_n3765_), .ZN(new_n3994_));
  OAI21_X1   g03738(.A1(new_n3994_), .A2(new_n3767_), .B(new_n3770_), .ZN(new_n3995_));
  NOR3_X1    g03739(.A1(new_n3988_), .A2(new_n3987_), .A3(new_n3986_), .ZN(new_n3996_));
  AOI21_X1   g03740(.A1(new_n3978_), .A2(new_n3984_), .B(new_n3821_), .ZN(new_n3997_));
  NOR2_X1    g03741(.A1(new_n3996_), .A2(new_n3997_), .ZN(new_n3998_));
  AOI21_X1   g03742(.A1(new_n3995_), .A2(new_n3768_), .B(new_n3998_), .ZN(new_n3999_));
  OAI21_X1   g03743(.A1(new_n3991_), .A2(new_n3999_), .B(new_n3811_), .ZN(new_n4000_));
  XOR2_X1    g03744(.A1(new_n3810_), .A2(\a[5] ), .Z(new_n4001_));
  NAND3_X1   g03745(.A1(new_n3995_), .A2(new_n3768_), .A3(new_n3998_), .ZN(new_n4002_));
  OAI21_X1   g03746(.A1(new_n3754_), .A2(new_n3771_), .B(new_n3768_), .ZN(new_n4003_));
  NAND2_X1   g03747(.A1(new_n4003_), .A2(new_n3990_), .ZN(new_n4004_));
  NAND3_X1   g03748(.A1(new_n4004_), .A2(new_n4001_), .A3(new_n4002_), .ZN(new_n4005_));
  NAND2_X1   g03749(.A1(new_n4005_), .A2(new_n4000_), .ZN(new_n4006_));
  NAND2_X1   g03750(.A1(new_n4006_), .A2(new_n3806_), .ZN(new_n4007_));
  XOR2_X1    g03751(.A1(new_n3640_), .A2(new_n312_), .Z(new_n4008_));
  NOR3_X1    g03752(.A1(new_n3771_), .A2(new_n3772_), .A3(new_n3770_), .ZN(new_n4009_));
  AOI21_X1   g03753(.A1(new_n3768_), .A2(new_n3766_), .B(new_n3754_), .ZN(new_n4010_));
  OAI21_X1   g03754(.A1(new_n4010_), .A2(new_n4009_), .B(new_n4008_), .ZN(new_n4011_));
  NAND2_X1   g03755(.A1(new_n3777_), .A2(new_n4011_), .ZN(new_n4012_));
  NAND4_X1   g03756(.A1(new_n4012_), .A2(new_n4005_), .A3(new_n4000_), .A4(new_n3775_), .ZN(new_n4013_));
  NAND2_X1   g03757(.A1(new_n4007_), .A2(new_n4013_), .ZN(new_n4014_));
  NAND3_X1   g03758(.A1(new_n3801_), .A2(new_n3803_), .A3(new_n4014_), .ZN(new_n4015_));
  INV_X1     g03759(.I(new_n4014_), .ZN(new_n4016_));
  OAI21_X1   g03760(.A1(new_n3785_), .A2(new_n3802_), .B(new_n4016_), .ZN(new_n4017_));
  NAND2_X1   g03761(.A1(new_n4017_), .A2(new_n4015_), .ZN(new_n4018_));
  XOR2_X1    g03762(.A1(new_n4018_), .A2(new_n3800_), .Z(\f[31] ));
  AOI21_X1   g03763(.A1(new_n3801_), .A2(new_n3803_), .B(new_n4014_), .ZN(new_n4020_));
  OAI21_X1   g03764(.A1(new_n3799_), .A2(new_n4020_), .B(new_n4015_), .ZN(new_n4021_));
  INV_X1     g03765(.I(\b[31] ), .ZN(new_n4022_));
  INV_X1     g03766(.I(\b[32] ), .ZN(new_n4023_));
  OAI22_X1   g03767(.A1(new_n277_), .A2(new_n4023_), .B1(new_n4022_), .B2(new_n262_), .ZN(new_n4024_));
  AOI21_X1   g03768(.A1(\b[30] ), .A2(new_n283_), .B(new_n4024_), .ZN(new_n4025_));
  XOR2_X1    g03769(.A1(\b[31] ), .A2(\b[32] ), .Z(new_n4026_));
  OAI21_X1   g03770(.A1(new_n3793_), .A2(\b[30] ), .B(\b[31] ), .ZN(new_n4027_));
  NAND2_X1   g03771(.A1(new_n3792_), .A2(\b[30] ), .ZN(new_n4028_));
  NAND2_X1   g03772(.A1(new_n4027_), .A2(new_n4028_), .ZN(new_n4029_));
  XOR2_X1    g03773(.A1(new_n4029_), .A2(new_n4026_), .Z(new_n4030_));
  INV_X1     g03774(.I(new_n4030_), .ZN(new_n4031_));
  OAI21_X1   g03775(.A1(new_n4031_), .A2(new_n279_), .B(new_n4025_), .ZN(new_n4032_));
  XOR2_X1    g03776(.A1(new_n4032_), .A2(\a[2] ), .Z(new_n4033_));
  NOR3_X1    g03777(.A1(new_n3963_), .A2(new_n3973_), .A3(new_n3971_), .ZN(new_n4034_));
  OAI22_X1   g03778(.A1(new_n713_), .A2(new_n2463_), .B1(new_n2142_), .B2(new_n717_), .ZN(new_n4035_));
  AOI21_X1   g03779(.A1(\b[21] ), .A2(new_n1126_), .B(new_n4035_), .ZN(new_n4036_));
  OAI21_X1   g03780(.A1(new_n3552_), .A2(new_n986_), .B(new_n4036_), .ZN(new_n4037_));
  XOR2_X1    g03781(.A1(new_n4037_), .A2(\a[11] ), .Z(new_n4038_));
  OAI22_X1   g03782(.A1(new_n993_), .A2(new_n1860_), .B1(new_n1859_), .B2(new_n997_), .ZN(new_n4039_));
  AOI21_X1   g03783(.A1(\b[18] ), .A2(new_n1486_), .B(new_n4039_), .ZN(new_n4040_));
  OAI21_X1   g03784(.A1(new_n1871_), .A2(new_n1323_), .B(new_n4040_), .ZN(new_n4041_));
  XOR2_X1    g03785(.A1(new_n4041_), .A2(\a[14] ), .Z(new_n4042_));
  INV_X1     g03786(.I(new_n4042_), .ZN(new_n4043_));
  OAI22_X1   g03787(.A1(new_n1592_), .A2(new_n1432_), .B1(new_n1296_), .B2(new_n1505_), .ZN(new_n4044_));
  AOI21_X1   g03788(.A1(\b[15] ), .A2(new_n1584_), .B(new_n4044_), .ZN(new_n4045_));
  OAI21_X1   g03789(.A1(new_n1444_), .A2(new_n1732_), .B(new_n4045_), .ZN(new_n4046_));
  XOR2_X1    g03790(.A1(new_n4046_), .A2(new_n1344_), .Z(new_n4047_));
  NAND2_X1   g03791(.A1(new_n3872_), .A2(new_n554_), .ZN(new_n4048_));
  AOI22_X1   g03792(.A1(new_n3864_), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n3869_), .ZN(new_n4049_));
  XOR2_X1    g03793(.A1(\a[29] ), .A2(\a[30] ), .Z(new_n4050_));
  AOI21_X1   g03794(.A1(new_n3867_), .A2(\a[32] ), .B(\a[29] ), .ZN(new_n4051_));
  AOI21_X1   g03795(.A1(\a[31] ), .A2(new_n3876_), .B(new_n3264_), .ZN(new_n4052_));
  NOR3_X1    g03796(.A1(new_n4050_), .A2(new_n4051_), .A3(new_n4052_), .ZN(new_n4053_));
  NAND2_X1   g03797(.A1(new_n4053_), .A2(\b[0] ), .ZN(new_n4054_));
  NAND3_X1   g03798(.A1(new_n4049_), .A2(new_n4048_), .A3(new_n4054_), .ZN(new_n4055_));
  XOR2_X1    g03799(.A1(new_n4055_), .A2(new_n3876_), .Z(new_n4056_));
  NAND4_X1   g03800(.A1(new_n3870_), .A2(\a[32] ), .A3(new_n3873_), .A4(new_n3655_), .ZN(new_n4057_));
  XOR2_X1    g03801(.A1(new_n4056_), .A2(new_n4057_), .Z(new_n4058_));
  OAI21_X1   g03802(.A1(new_n3857_), .A2(new_n3890_), .B(new_n3882_), .ZN(new_n4059_));
  NAND2_X1   g03803(.A1(new_n4059_), .A2(new_n4058_), .ZN(new_n4060_));
  NAND2_X1   g03804(.A1(new_n4056_), .A2(new_n4057_), .ZN(new_n4061_));
  NOR4_X1    g03805(.A1(new_n4055_), .A2(new_n3874_), .A3(new_n3876_), .A4(new_n3654_), .ZN(new_n4062_));
  INV_X1     g03806(.I(new_n4062_), .ZN(new_n4063_));
  NAND2_X1   g03807(.A1(new_n4061_), .A2(new_n4063_), .ZN(new_n4064_));
  AOI21_X1   g03808(.A1(new_n3888_), .A2(new_n3884_), .B(new_n3889_), .ZN(new_n4065_));
  NAND2_X1   g03809(.A1(new_n4065_), .A2(new_n4064_), .ZN(new_n4066_));
  OAI22_X1   g03810(.A1(new_n377_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n339_), .ZN(new_n4067_));
  AOI21_X1   g03811(.A1(\b[3] ), .A2(new_n3456_), .B(new_n4067_), .ZN(new_n4068_));
  OAI21_X1   g03812(.A1(new_n566_), .A2(new_n3261_), .B(new_n4068_), .ZN(new_n4069_));
  XOR2_X1    g03813(.A1(new_n4069_), .A2(new_n3264_), .Z(new_n4070_));
  OAI22_X1   g03814(.A1(new_n2703_), .A2(new_n577_), .B1(new_n471_), .B2(new_n2708_), .ZN(new_n4071_));
  NOR2_X1    g03815(.A1(new_n2924_), .A2(new_n438_), .ZN(new_n4072_));
  NOR2_X1    g03816(.A1(new_n4071_), .A2(new_n4072_), .ZN(new_n4073_));
  INV_X1     g03817(.I(new_n4073_), .ZN(new_n4074_));
  AOI21_X1   g03818(.A1(new_n799_), .A2(new_n2722_), .B(new_n4074_), .ZN(new_n4075_));
  NOR2_X1    g03819(.A1(new_n4075_), .A2(new_n2714_), .ZN(new_n4076_));
  OAI21_X1   g03820(.A1(new_n587_), .A2(new_n2711_), .B(new_n4073_), .ZN(new_n4077_));
  NOR2_X1    g03821(.A1(new_n4077_), .A2(\a[26] ), .ZN(new_n4078_));
  OAI21_X1   g03822(.A1(new_n4076_), .A2(new_n4078_), .B(new_n4070_), .ZN(new_n4079_));
  XOR2_X1    g03823(.A1(new_n4069_), .A2(\a[29] ), .Z(new_n4080_));
  NAND2_X1   g03824(.A1(new_n4077_), .A2(\a[26] ), .ZN(new_n4081_));
  NAND2_X1   g03825(.A1(new_n4075_), .A2(new_n2714_), .ZN(new_n4082_));
  NAND3_X1   g03826(.A1(new_n4082_), .A2(new_n4081_), .A3(new_n4080_), .ZN(new_n4083_));
  NAND4_X1   g03827(.A1(new_n4066_), .A2(new_n4060_), .A3(new_n4079_), .A4(new_n4083_), .ZN(new_n4084_));
  NOR2_X1    g03828(.A1(new_n4065_), .A2(new_n4064_), .ZN(new_n4085_));
  NOR2_X1    g03829(.A1(new_n4059_), .A2(new_n4058_), .ZN(new_n4086_));
  AOI21_X1   g03830(.A1(new_n4082_), .A2(new_n4081_), .B(new_n4080_), .ZN(new_n4087_));
  NOR3_X1    g03831(.A1(new_n4076_), .A2(new_n4078_), .A3(new_n4070_), .ZN(new_n4088_));
  OAI22_X1   g03832(.A1(new_n4085_), .A2(new_n4086_), .B1(new_n4087_), .B2(new_n4088_), .ZN(new_n4089_));
  NAND2_X1   g03833(.A1(new_n4089_), .A2(new_n4084_), .ZN(new_n4090_));
  OAI21_X1   g03834(.A1(new_n3852_), .A2(new_n3904_), .B(new_n3900_), .ZN(new_n4091_));
  NOR2_X1    g03835(.A1(new_n4091_), .A2(new_n4090_), .ZN(new_n4092_));
  INV_X1     g03836(.I(new_n4090_), .ZN(new_n4093_));
  AOI21_X1   g03837(.A1(new_n3903_), .A2(new_n3898_), .B(new_n3905_), .ZN(new_n4094_));
  NOR2_X1    g03838(.A1(new_n4093_), .A2(new_n4094_), .ZN(new_n4095_));
  NOR2_X1    g03839(.A1(new_n4095_), .A2(new_n4092_), .ZN(new_n4096_));
  INV_X1     g03840(.I(new_n4096_), .ZN(new_n4097_));
  INV_X1     g03841(.I(new_n3915_), .ZN(new_n4098_));
  OAI21_X1   g03842(.A1(new_n3689_), .A2(new_n3685_), .B(new_n3674_), .ZN(new_n4099_));
  NAND3_X1   g03843(.A1(new_n3912_), .A2(new_n3913_), .A3(new_n3914_), .ZN(new_n4100_));
  NAND3_X1   g03844(.A1(new_n4099_), .A2(new_n3690_), .A3(new_n4100_), .ZN(new_n4101_));
  NAND2_X1   g03845(.A1(new_n4101_), .A2(new_n4098_), .ZN(new_n4102_));
  NAND2_X1   g03846(.A1(new_n4102_), .A2(new_n4097_), .ZN(new_n4103_));
  NAND3_X1   g03847(.A1(new_n4101_), .A2(new_n4098_), .A3(new_n4096_), .ZN(new_n4104_));
  AOI22_X1   g03848(.A1(new_n1738_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n1743_), .ZN(new_n4105_));
  OAI21_X1   g03849(.A1(new_n941_), .A2(new_n1931_), .B(new_n4105_), .ZN(new_n4106_));
  INV_X1     g03850(.I(new_n4106_), .ZN(new_n4107_));
  OAI21_X1   g03851(.A1(new_n1103_), .A2(new_n1757_), .B(new_n4107_), .ZN(new_n4108_));
  NAND2_X1   g03852(.A1(new_n4108_), .A2(\a[20] ), .ZN(new_n4109_));
  INV_X1     g03853(.I(new_n4109_), .ZN(new_n4110_));
  NOR2_X1    g03854(.A1(new_n4108_), .A2(\a[20] ), .ZN(new_n4111_));
  OAI22_X1   g03855(.A1(new_n2189_), .A2(new_n852_), .B1(new_n776_), .B2(new_n2194_), .ZN(new_n4112_));
  AOI21_X1   g03856(.A1(\b[9] ), .A2(new_n2361_), .B(new_n4112_), .ZN(new_n4113_));
  OAI21_X1   g03857(.A1(new_n859_), .A2(new_n2197_), .B(new_n4113_), .ZN(new_n4114_));
  XOR2_X1    g03858(.A1(new_n4114_), .A2(\a[23] ), .Z(new_n4115_));
  OAI21_X1   g03859(.A1(new_n4110_), .A2(new_n4111_), .B(new_n4115_), .ZN(new_n4116_));
  INV_X1     g03860(.I(new_n4111_), .ZN(new_n4117_));
  XOR2_X1    g03861(.A1(new_n4114_), .A2(new_n2200_), .Z(new_n4118_));
  NAND3_X1   g03862(.A1(new_n4117_), .A2(new_n4109_), .A3(new_n4118_), .ZN(new_n4119_));
  AOI22_X1   g03863(.A1(new_n4103_), .A2(new_n4104_), .B1(new_n4116_), .B2(new_n4119_), .ZN(new_n4120_));
  AOI21_X1   g03864(.A1(new_n3929_), .A2(new_n4100_), .B(new_n3915_), .ZN(new_n4121_));
  NOR2_X1    g03865(.A1(new_n4121_), .A2(new_n4096_), .ZN(new_n4122_));
  INV_X1     g03866(.I(new_n4104_), .ZN(new_n4123_));
  AOI21_X1   g03867(.A1(new_n4117_), .A2(new_n4109_), .B(new_n4118_), .ZN(new_n4124_));
  NOR3_X1    g03868(.A1(new_n4110_), .A2(new_n4111_), .A3(new_n4115_), .ZN(new_n4125_));
  NOR4_X1    g03869(.A1(new_n4123_), .A2(new_n4122_), .A3(new_n4124_), .A4(new_n4125_), .ZN(new_n4126_));
  NOR2_X1    g03870(.A1(new_n4126_), .A2(new_n4120_), .ZN(new_n4127_));
  AOI21_X1   g03871(.A1(new_n3935_), .A2(new_n3704_), .B(new_n3928_), .ZN(new_n4128_));
  NOR3_X1    g03872(.A1(new_n4128_), .A2(new_n4127_), .A3(new_n3932_), .ZN(new_n4129_));
  OAI22_X1   g03873(.A1(new_n4123_), .A2(new_n4122_), .B1(new_n4124_), .B2(new_n4125_), .ZN(new_n4130_));
  NAND4_X1   g03874(.A1(new_n4103_), .A2(new_n4104_), .A3(new_n4116_), .A4(new_n4119_), .ZN(new_n4131_));
  NAND2_X1   g03875(.A1(new_n4130_), .A2(new_n4131_), .ZN(new_n4132_));
  AOI21_X1   g03876(.A1(new_n3848_), .A2(new_n3936_), .B(new_n3932_), .ZN(new_n4133_));
  NOR2_X1    g03877(.A1(new_n4133_), .A2(new_n4132_), .ZN(new_n4134_));
  OAI21_X1   g03878(.A1(new_n4134_), .A2(new_n4129_), .B(new_n4047_), .ZN(new_n4135_));
  XOR2_X1    g03879(.A1(new_n4046_), .A2(\a[17] ), .Z(new_n4136_));
  NAND2_X1   g03880(.A1(new_n3848_), .A2(new_n3936_), .ZN(new_n4137_));
  NAND3_X1   g03881(.A1(new_n4137_), .A2(new_n4132_), .A3(new_n3937_), .ZN(new_n4138_));
  OAI21_X1   g03882(.A1(new_n4128_), .A2(new_n3932_), .B(new_n4127_), .ZN(new_n4139_));
  NAND3_X1   g03883(.A1(new_n4139_), .A2(new_n4138_), .A3(new_n4136_), .ZN(new_n4140_));
  NAND2_X1   g03884(.A1(new_n4135_), .A2(new_n4140_), .ZN(new_n4141_));
  AOI21_X1   g03885(.A1(new_n3939_), .A2(new_n3934_), .B(new_n3941_), .ZN(new_n4142_));
  INV_X1     g03886(.I(new_n4142_), .ZN(new_n4143_));
  AOI21_X1   g03887(.A1(new_n3947_), .A2(new_n4143_), .B(new_n4141_), .ZN(new_n4144_));
  AOI21_X1   g03888(.A1(new_n4139_), .A2(new_n4138_), .B(new_n4136_), .ZN(new_n4145_));
  NOR3_X1    g03889(.A1(new_n4134_), .A2(new_n4129_), .A3(new_n4047_), .ZN(new_n4146_));
  NOR2_X1    g03890(.A1(new_n4145_), .A2(new_n4146_), .ZN(new_n4147_));
  NOR3_X1    g03891(.A1(new_n3959_), .A2(new_n4147_), .A3(new_n4142_), .ZN(new_n4148_));
  NOR3_X1    g03892(.A1(new_n4144_), .A2(new_n4148_), .A3(new_n4043_), .ZN(new_n4149_));
  OAI21_X1   g03893(.A1(new_n3959_), .A2(new_n4142_), .B(new_n4147_), .ZN(new_n4150_));
  NAND3_X1   g03894(.A1(new_n3947_), .A2(new_n4141_), .A3(new_n4143_), .ZN(new_n4151_));
  AOI21_X1   g03895(.A1(new_n4150_), .A2(new_n4151_), .B(new_n4042_), .ZN(new_n4152_));
  NOR2_X1    g03896(.A1(new_n4149_), .A2(new_n4152_), .ZN(new_n4153_));
  OAI21_X1   g03897(.A1(new_n3963_), .A2(new_n3968_), .B(new_n4153_), .ZN(new_n4154_));
  NAND3_X1   g03898(.A1(new_n4150_), .A2(new_n4151_), .A3(new_n4042_), .ZN(new_n4155_));
  OAI21_X1   g03899(.A1(new_n4144_), .A2(new_n4148_), .B(new_n4043_), .ZN(new_n4156_));
  NAND2_X1   g03900(.A1(new_n4156_), .A2(new_n4155_), .ZN(new_n4157_));
  NAND3_X1   g03901(.A1(new_n3974_), .A2(new_n3957_), .A3(new_n4157_), .ZN(new_n4158_));
  NAND3_X1   g03902(.A1(new_n4154_), .A2(new_n4038_), .A3(new_n4158_), .ZN(new_n4159_));
  INV_X1     g03903(.I(new_n4038_), .ZN(new_n4160_));
  AOI21_X1   g03904(.A1(new_n3974_), .A2(new_n3957_), .B(new_n4157_), .ZN(new_n4161_));
  NOR3_X1    g03905(.A1(new_n3963_), .A2(new_n3968_), .A3(new_n4153_), .ZN(new_n4162_));
  OAI21_X1   g03906(.A1(new_n4162_), .A2(new_n4161_), .B(new_n4160_), .ZN(new_n4163_));
  NAND2_X1   g03907(.A1(new_n4163_), .A2(new_n4159_), .ZN(new_n4164_));
  OAI21_X1   g03908(.A1(new_n3987_), .A2(new_n4034_), .B(new_n4164_), .ZN(new_n4165_));
  INV_X1     g03909(.I(new_n4034_), .ZN(new_n4166_));
  NOR3_X1    g03910(.A1(new_n4162_), .A2(new_n4160_), .A3(new_n4161_), .ZN(new_n4167_));
  AOI21_X1   g03911(.A1(new_n4154_), .A2(new_n4158_), .B(new_n4038_), .ZN(new_n4168_));
  NOR2_X1    g03912(.A1(new_n4167_), .A2(new_n4168_), .ZN(new_n4169_));
  NAND3_X1   g03913(.A1(new_n3978_), .A2(new_n4166_), .A3(new_n4169_), .ZN(new_n4170_));
  AOI22_X1   g03914(.A1(new_n518_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n636_), .ZN(new_n4171_));
  OAI21_X1   g03915(.A1(new_n2495_), .A2(new_n917_), .B(new_n4171_), .ZN(new_n4172_));
  AOI21_X1   g03916(.A1(new_n3407_), .A2(new_n618_), .B(new_n4172_), .ZN(new_n4173_));
  XOR2_X1    g03917(.A1(new_n4173_), .A2(new_n488_), .Z(new_n4174_));
  INV_X1     g03918(.I(new_n4174_), .ZN(new_n4175_));
  NAND3_X1   g03919(.A1(new_n4170_), .A2(new_n4165_), .A3(new_n4175_), .ZN(new_n4176_));
  AOI21_X1   g03920(.A1(new_n3978_), .A2(new_n4166_), .B(new_n4169_), .ZN(new_n4177_));
  NOR3_X1    g03921(.A1(new_n3987_), .A2(new_n4164_), .A3(new_n4034_), .ZN(new_n4178_));
  OAI21_X1   g03922(.A1(new_n4177_), .A2(new_n4178_), .B(new_n4174_), .ZN(new_n4179_));
  NAND2_X1   g03923(.A1(new_n4179_), .A2(new_n4176_), .ZN(new_n4180_));
  AOI21_X1   g03924(.A1(new_n4002_), .A2(new_n3985_), .B(new_n4180_), .ZN(new_n4181_));
  INV_X1     g03925(.I(new_n4181_), .ZN(new_n4182_));
  AOI21_X1   g03926(.A1(new_n3770_), .A2(new_n3766_), .B(new_n3772_), .ZN(new_n4183_));
  AOI21_X1   g03927(.A1(new_n4183_), .A2(new_n3998_), .B(new_n3996_), .ZN(new_n4184_));
  NAND2_X1   g03928(.A1(new_n4184_), .A2(new_n4180_), .ZN(new_n4185_));
  NAND2_X1   g03929(.A1(new_n4182_), .A2(new_n4185_), .ZN(new_n4186_));
  INV_X1     g03930(.I(new_n3594_), .ZN(new_n4187_));
  NOR2_X1    g03931(.A1(new_n4187_), .A2(new_n3595_), .ZN(new_n4188_));
  AOI22_X1   g03932(.A1(new_n800_), .A2(\b[28] ), .B1(\b[29] ), .B2(new_n333_), .ZN(new_n4189_));
  OAI21_X1   g03933(.A1(new_n3158_), .A2(new_n392_), .B(new_n4189_), .ZN(new_n4190_));
  AOI21_X1   g03934(.A1(new_n4188_), .A2(new_n330_), .B(new_n4190_), .ZN(new_n4191_));
  XOR2_X1    g03935(.A1(new_n4191_), .A2(new_n312_), .Z(new_n4192_));
  INV_X1     g03936(.I(new_n4192_), .ZN(new_n4193_));
  NOR3_X1    g03937(.A1(new_n3991_), .A2(new_n3999_), .A3(new_n4001_), .ZN(new_n4194_));
  INV_X1     g03938(.I(new_n4194_), .ZN(new_n4195_));
  AOI21_X1   g03939(.A1(new_n4007_), .A2(new_n4195_), .B(new_n4193_), .ZN(new_n4196_));
  AOI22_X1   g03940(.A1(new_n4012_), .A2(new_n3775_), .B1(new_n4005_), .B2(new_n4000_), .ZN(new_n4197_));
  NOR3_X1    g03941(.A1(new_n4197_), .A2(new_n4192_), .A3(new_n4194_), .ZN(new_n4198_));
  NOR3_X1    g03942(.A1(new_n4196_), .A2(new_n4198_), .A3(new_n4186_), .ZN(new_n4199_));
  INV_X1     g03943(.I(new_n4186_), .ZN(new_n4200_));
  OAI21_X1   g03944(.A1(new_n4197_), .A2(new_n4194_), .B(new_n4192_), .ZN(new_n4201_));
  NAND3_X1   g03945(.A1(new_n4007_), .A2(new_n4193_), .A3(new_n4195_), .ZN(new_n4202_));
  AOI21_X1   g03946(.A1(new_n4202_), .A2(new_n4201_), .B(new_n4200_), .ZN(new_n4203_));
  NOR2_X1    g03947(.A1(new_n4199_), .A2(new_n4203_), .ZN(new_n4204_));
  NOR2_X1    g03948(.A1(new_n4204_), .A2(new_n4033_), .ZN(new_n4205_));
  INV_X1     g03949(.I(new_n4205_), .ZN(new_n4206_));
  NAND2_X1   g03950(.A1(new_n4204_), .A2(new_n4033_), .ZN(new_n4207_));
  NAND2_X1   g03951(.A1(new_n4206_), .A2(new_n4207_), .ZN(new_n4208_));
  XOR2_X1    g03952(.A1(new_n4021_), .A2(new_n4208_), .Z(\f[32] ));
  AOI21_X1   g03953(.A1(new_n4021_), .A2(new_n4207_), .B(new_n4205_), .ZN(new_n4210_));
  NOR2_X1    g03954(.A1(new_n284_), .A2(new_n4022_), .ZN(new_n4211_));
  INV_X1     g03955(.I(new_n4211_), .ZN(new_n4212_));
  AOI22_X1   g03956(.A1(new_n267_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n261_), .ZN(new_n4213_));
  AOI21_X1   g03957(.A1(new_n4029_), .A2(\b[32] ), .B(new_n4022_), .ZN(new_n4214_));
  NOR2_X1    g03958(.A1(new_n4029_), .A2(\b[32] ), .ZN(new_n4215_));
  NOR2_X1    g03959(.A1(new_n4214_), .A2(new_n4215_), .ZN(new_n4216_));
  NOR2_X1    g03960(.A1(new_n4029_), .A2(\b[33] ), .ZN(new_n4217_));
  INV_X1     g03961(.I(new_n4217_), .ZN(new_n4218_));
  NAND2_X1   g03962(.A1(new_n4029_), .A2(\b[33] ), .ZN(new_n4219_));
  AOI21_X1   g03963(.A1(new_n4218_), .A2(new_n4219_), .B(new_n4216_), .ZN(new_n4220_));
  INV_X1     g03964(.I(new_n4219_), .ZN(new_n4221_));
  NOR4_X1    g03965(.A1(new_n4221_), .A2(new_n4214_), .A3(new_n4215_), .A4(new_n4217_), .ZN(new_n4222_));
  NOR2_X1    g03966(.A1(new_n4220_), .A2(new_n4222_), .ZN(new_n4223_));
  NAND2_X1   g03967(.A1(new_n4223_), .A2(new_n265_), .ZN(new_n4224_));
  NAND3_X1   g03968(.A1(new_n4224_), .A2(new_n4212_), .A3(new_n4213_), .ZN(new_n4225_));
  AND2_X2    g03969(.A1(new_n4225_), .A2(\a[2] ), .Z(new_n4226_));
  NOR2_X1    g03970(.A1(new_n4225_), .A2(\a[2] ), .ZN(new_n4227_));
  NOR2_X1    g03971(.A1(new_n4226_), .A2(new_n4227_), .ZN(new_n4228_));
  AOI21_X1   g03972(.A1(new_n4186_), .A2(new_n4201_), .B(new_n4198_), .ZN(new_n4229_));
  INV_X1     g03973(.I(new_n3634_), .ZN(new_n4230_));
  AOI22_X1   g03974(.A1(new_n800_), .A2(\b[29] ), .B1(\b[30] ), .B2(new_n333_), .ZN(new_n4231_));
  OAI21_X1   g03975(.A1(new_n3185_), .A2(new_n392_), .B(new_n4231_), .ZN(new_n4232_));
  AOI21_X1   g03976(.A1(new_n4230_), .A2(new_n330_), .B(new_n4232_), .ZN(new_n4233_));
  XOR2_X1    g03977(.A1(new_n4233_), .A2(new_n312_), .Z(new_n4234_));
  NAND2_X1   g03978(.A1(new_n4058_), .A2(new_n4080_), .ZN(new_n4235_));
  NOR2_X1    g03979(.A1(new_n4058_), .A2(new_n4080_), .ZN(new_n4236_));
  OAI21_X1   g03980(.A1(new_n4065_), .A2(new_n4236_), .B(new_n4235_), .ZN(new_n4237_));
  OAI22_X1   g03981(.A1(new_n438_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n377_), .ZN(new_n4238_));
  AOI21_X1   g03982(.A1(\b[4] ), .A2(new_n3456_), .B(new_n4238_), .ZN(new_n4239_));
  OAI21_X1   g03983(.A1(new_n450_), .A2(new_n3261_), .B(new_n4239_), .ZN(new_n4240_));
  XOR2_X1    g03984(.A1(new_n4240_), .A2(\a[29] ), .Z(new_n4241_));
  NAND2_X1   g03985(.A1(new_n4053_), .A2(\b[1] ), .ZN(new_n4242_));
  AOI22_X1   g03986(.A1(new_n3864_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n3869_), .ZN(new_n4243_));
  NAND2_X1   g03987(.A1(new_n299_), .A2(new_n3872_), .ZN(new_n4244_));
  NAND3_X1   g03988(.A1(new_n4244_), .A2(new_n4243_), .A3(new_n4242_), .ZN(new_n4245_));
  XOR2_X1    g03989(.A1(new_n4245_), .A2(\a[32] ), .Z(new_n4246_));
  XNOR2_X1   g03990(.A1(\a[32] ), .A2(\a[33] ), .ZN(new_n4247_));
  NOR2_X1    g03991(.A1(new_n4247_), .A2(new_n258_), .ZN(new_n4248_));
  INV_X1     g03992(.I(new_n4248_), .ZN(new_n4249_));
  NOR2_X1    g03993(.A1(new_n4246_), .A2(new_n4249_), .ZN(new_n4250_));
  XOR2_X1    g03994(.A1(new_n4245_), .A2(new_n3876_), .Z(new_n4251_));
  NOR2_X1    g03995(.A1(new_n4251_), .A2(new_n4248_), .ZN(new_n4252_));
  OAI21_X1   g03996(.A1(new_n4250_), .A2(new_n4252_), .B(new_n4063_), .ZN(new_n4253_));
  NAND2_X1   g03997(.A1(new_n4251_), .A2(new_n4248_), .ZN(new_n4254_));
  NAND2_X1   g03998(.A1(new_n4246_), .A2(new_n4249_), .ZN(new_n4255_));
  NAND3_X1   g03999(.A1(new_n4254_), .A2(new_n4255_), .A3(new_n4062_), .ZN(new_n4256_));
  NAND3_X1   g04000(.A1(new_n4253_), .A2(new_n4256_), .A3(new_n4241_), .ZN(new_n4257_));
  XOR2_X1    g04001(.A1(new_n4240_), .A2(new_n3264_), .Z(new_n4258_));
  AOI21_X1   g04002(.A1(new_n4254_), .A2(new_n4255_), .B(new_n4062_), .ZN(new_n4259_));
  NOR3_X1    g04003(.A1(new_n4250_), .A2(new_n4252_), .A3(new_n4063_), .ZN(new_n4260_));
  OAI21_X1   g04004(.A1(new_n4259_), .A2(new_n4260_), .B(new_n4258_), .ZN(new_n4261_));
  NAND2_X1   g04005(.A1(new_n4261_), .A2(new_n4257_), .ZN(new_n4262_));
  NAND2_X1   g04006(.A1(new_n4237_), .A2(new_n4262_), .ZN(new_n4263_));
  NOR2_X1    g04007(.A1(new_n4064_), .A2(new_n4070_), .ZN(new_n4264_));
  NAND2_X1   g04008(.A1(new_n4064_), .A2(new_n4070_), .ZN(new_n4265_));
  AOI21_X1   g04009(.A1(new_n4059_), .A2(new_n4265_), .B(new_n4264_), .ZN(new_n4266_));
  NOR3_X1    g04010(.A1(new_n4259_), .A2(new_n4260_), .A3(new_n4258_), .ZN(new_n4267_));
  AOI21_X1   g04011(.A1(new_n4253_), .A2(new_n4256_), .B(new_n4241_), .ZN(new_n4268_));
  NOR2_X1    g04012(.A1(new_n4267_), .A2(new_n4268_), .ZN(new_n4269_));
  NAND2_X1   g04013(.A1(new_n4269_), .A2(new_n4266_), .ZN(new_n4270_));
  NAND2_X1   g04014(.A1(new_n4263_), .A2(new_n4270_), .ZN(new_n4271_));
  AOI22_X1   g04015(.A1(new_n2716_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n2719_), .ZN(new_n4272_));
  OAI21_X1   g04016(.A1(new_n471_), .A2(new_n2924_), .B(new_n4272_), .ZN(new_n4273_));
  AOI21_X1   g04017(.A1(new_n676_), .A2(new_n2722_), .B(new_n4273_), .ZN(new_n4274_));
  XOR2_X1    g04018(.A1(new_n4274_), .A2(new_n2714_), .Z(new_n4275_));
  NOR2_X1    g04019(.A1(new_n4076_), .A2(new_n4078_), .ZN(new_n4276_));
  NAND3_X1   g04020(.A1(new_n4235_), .A2(new_n4059_), .A3(new_n4265_), .ZN(new_n4277_));
  OAI21_X1   g04021(.A1(new_n4236_), .A2(new_n4264_), .B(new_n4065_), .ZN(new_n4278_));
  NAND3_X1   g04022(.A1(new_n4278_), .A2(new_n4277_), .A3(new_n4276_), .ZN(new_n4279_));
  OAI21_X1   g04023(.A1(new_n4094_), .A2(new_n4090_), .B(new_n4279_), .ZN(new_n4280_));
  NAND2_X1   g04024(.A1(new_n4280_), .A2(new_n4275_), .ZN(new_n4281_));
  INV_X1     g04025(.I(new_n4281_), .ZN(new_n4282_));
  NOR2_X1    g04026(.A1(new_n4280_), .A2(new_n4275_), .ZN(new_n4283_));
  NOR3_X1    g04027(.A1(new_n4282_), .A2(new_n4271_), .A3(new_n4283_), .ZN(new_n4284_));
  INV_X1     g04028(.I(new_n4271_), .ZN(new_n4285_));
  INV_X1     g04029(.I(new_n4275_), .ZN(new_n4286_));
  INV_X1     g04030(.I(new_n4279_), .ZN(new_n4287_));
  AOI21_X1   g04031(.A1(new_n4093_), .A2(new_n4091_), .B(new_n4287_), .ZN(new_n4288_));
  NAND2_X1   g04032(.A1(new_n4288_), .A2(new_n4286_), .ZN(new_n4289_));
  AOI21_X1   g04033(.A1(new_n4289_), .A2(new_n4281_), .B(new_n4285_), .ZN(new_n4290_));
  NOR2_X1    g04034(.A1(new_n4284_), .A2(new_n4290_), .ZN(new_n4291_));
  INV_X1     g04035(.I(new_n4291_), .ZN(new_n4292_));
  AOI22_X1   g04036(.A1(new_n2202_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n2205_), .ZN(new_n4293_));
  OAI21_X1   g04037(.A1(new_n776_), .A2(new_n2370_), .B(new_n4293_), .ZN(new_n4294_));
  AOI21_X1   g04038(.A1(new_n1194_), .A2(new_n2208_), .B(new_n4294_), .ZN(new_n4295_));
  XOR2_X1    g04039(.A1(new_n4295_), .A2(new_n2200_), .Z(new_n4296_));
  INV_X1     g04040(.I(new_n4296_), .ZN(new_n4297_));
  NAND2_X1   g04041(.A1(new_n4097_), .A2(new_n4115_), .ZN(new_n4298_));
  OAI21_X1   g04042(.A1(new_n4095_), .A2(new_n4092_), .B(new_n4118_), .ZN(new_n4299_));
  NAND2_X1   g04043(.A1(new_n4093_), .A2(new_n4094_), .ZN(new_n4300_));
  NAND2_X1   g04044(.A1(new_n4091_), .A2(new_n4090_), .ZN(new_n4301_));
  NAND3_X1   g04045(.A1(new_n4300_), .A2(new_n4115_), .A3(new_n4301_), .ZN(new_n4302_));
  NAND2_X1   g04046(.A1(new_n4299_), .A2(new_n4302_), .ZN(new_n4303_));
  NAND2_X1   g04047(.A1(new_n4102_), .A2(new_n4303_), .ZN(new_n4304_));
  AOI21_X1   g04048(.A1(new_n4304_), .A2(new_n4298_), .B(new_n4297_), .ZN(new_n4305_));
  AND2_X2    g04049(.A1(new_n4299_), .A2(new_n4302_), .Z(new_n4306_));
  OAI21_X1   g04050(.A1(new_n4306_), .A2(new_n4121_), .B(new_n4298_), .ZN(new_n4307_));
  NOR2_X1    g04051(.A1(new_n4307_), .A2(new_n4296_), .ZN(new_n4308_));
  NOR3_X1    g04052(.A1(new_n4308_), .A2(new_n4305_), .A3(new_n4292_), .ZN(new_n4309_));
  NOR2_X1    g04053(.A1(new_n4096_), .A2(new_n4118_), .ZN(new_n4310_));
  AOI22_X1   g04054(.A1(new_n4101_), .A2(new_n4098_), .B1(new_n4299_), .B2(new_n4302_), .ZN(new_n4311_));
  OAI21_X1   g04055(.A1(new_n4311_), .A2(new_n4310_), .B(new_n4296_), .ZN(new_n4312_));
  NAND3_X1   g04056(.A1(new_n4304_), .A2(new_n4297_), .A3(new_n4298_), .ZN(new_n4313_));
  AOI21_X1   g04057(.A1(new_n4313_), .A2(new_n4312_), .B(new_n4291_), .ZN(new_n4314_));
  NOR2_X1    g04058(.A1(new_n4309_), .A2(new_n4314_), .ZN(new_n4315_));
  OAI22_X1   g04059(.A1(new_n1751_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n1754_), .ZN(new_n4316_));
  AOI21_X1   g04060(.A1(\b[13] ), .A2(new_n1939_), .B(new_n4316_), .ZN(new_n4317_));
  OAI21_X1   g04061(.A1(new_n1275_), .A2(new_n1757_), .B(new_n4317_), .ZN(new_n4318_));
  XOR2_X1    g04062(.A1(new_n4318_), .A2(\a[20] ), .Z(new_n4319_));
  NAND2_X1   g04063(.A1(new_n4306_), .A2(new_n4121_), .ZN(new_n4320_));
  NAND4_X1   g04064(.A1(new_n4320_), .A2(new_n4304_), .A3(new_n4109_), .A4(new_n4117_), .ZN(new_n4321_));
  INV_X1     g04065(.I(new_n4321_), .ZN(new_n4322_));
  OAI21_X1   g04066(.A1(new_n4129_), .A2(new_n4322_), .B(new_n4319_), .ZN(new_n4323_));
  INV_X1     g04067(.I(new_n4319_), .ZN(new_n4324_));
  NAND3_X1   g04068(.A1(new_n4138_), .A2(new_n4324_), .A3(new_n4321_), .ZN(new_n4325_));
  NAND3_X1   g04069(.A1(new_n4323_), .A2(new_n4325_), .A3(new_n4315_), .ZN(new_n4326_));
  AOI21_X1   g04070(.A1(new_n4323_), .A2(new_n4325_), .B(new_n4315_), .ZN(new_n4327_));
  INV_X1     g04071(.I(new_n4327_), .ZN(new_n4328_));
  NAND2_X1   g04072(.A1(new_n4328_), .A2(new_n4326_), .ZN(new_n4329_));
  OAI22_X1   g04073(.A1(new_n1592_), .A2(new_n1553_), .B1(new_n1432_), .B2(new_n1505_), .ZN(new_n4330_));
  AOI21_X1   g04074(.A1(\b[16] ), .A2(new_n1584_), .B(new_n4330_), .ZN(new_n4331_));
  OAI21_X1   g04075(.A1(new_n1563_), .A2(new_n1732_), .B(new_n4331_), .ZN(new_n4332_));
  XOR2_X1    g04076(.A1(new_n4332_), .A2(\a[17] ), .Z(new_n4333_));
  INV_X1     g04077(.I(new_n4333_), .ZN(new_n4334_));
  AOI21_X1   g04078(.A1(new_n4150_), .A2(new_n4140_), .B(new_n4334_), .ZN(new_n4335_));
  NOR3_X1    g04079(.A1(new_n4144_), .A2(new_n4146_), .A3(new_n4333_), .ZN(new_n4336_));
  NOR3_X1    g04080(.A1(new_n4335_), .A2(new_n4336_), .A3(new_n4329_), .ZN(new_n4337_));
  OAI21_X1   g04081(.A1(new_n4335_), .A2(new_n4336_), .B(new_n4329_), .ZN(new_n4338_));
  INV_X1     g04082(.I(new_n4338_), .ZN(new_n4339_));
  NOR2_X1    g04083(.A1(new_n4339_), .A2(new_n4337_), .ZN(new_n4340_));
  OAI22_X1   g04084(.A1(new_n993_), .A2(new_n2027_), .B1(new_n1860_), .B2(new_n997_), .ZN(new_n4341_));
  AOI21_X1   g04085(.A1(\b[19] ), .A2(new_n1486_), .B(new_n4341_), .ZN(new_n4342_));
  OAI21_X1   g04086(.A1(new_n3727_), .A2(new_n1323_), .B(new_n4342_), .ZN(new_n4343_));
  XOR2_X1    g04087(.A1(new_n4343_), .A2(\a[14] ), .Z(new_n4344_));
  OAI21_X1   g04088(.A1(new_n4161_), .A2(new_n4149_), .B(new_n4344_), .ZN(new_n4345_));
  INV_X1     g04089(.I(new_n4344_), .ZN(new_n4346_));
  NAND3_X1   g04090(.A1(new_n4154_), .A2(new_n4155_), .A3(new_n4346_), .ZN(new_n4347_));
  NAND3_X1   g04091(.A1(new_n4347_), .A2(new_n4345_), .A3(new_n4340_), .ZN(new_n4348_));
  AOI21_X1   g04092(.A1(new_n4347_), .A2(new_n4345_), .B(new_n4340_), .ZN(new_n4349_));
  INV_X1     g04093(.I(new_n4349_), .ZN(new_n4350_));
  NAND2_X1   g04094(.A1(new_n4350_), .A2(new_n4348_), .ZN(new_n4351_));
  OAI22_X1   g04095(.A1(new_n713_), .A2(new_n2495_), .B1(new_n2463_), .B2(new_n717_), .ZN(new_n4352_));
  AOI21_X1   g04096(.A1(\b[22] ), .A2(new_n1126_), .B(new_n4352_), .ZN(new_n4353_));
  OAI21_X1   g04097(.A1(new_n2506_), .A2(new_n986_), .B(new_n4353_), .ZN(new_n4354_));
  XOR2_X1    g04098(.A1(new_n4354_), .A2(\a[11] ), .Z(new_n4355_));
  INV_X1     g04099(.I(new_n4355_), .ZN(new_n4356_));
  OAI21_X1   g04100(.A1(new_n3987_), .A2(new_n4034_), .B(new_n4169_), .ZN(new_n4357_));
  AOI21_X1   g04101(.A1(new_n4357_), .A2(new_n4159_), .B(new_n4356_), .ZN(new_n4358_));
  AOI21_X1   g04102(.A1(new_n3978_), .A2(new_n4166_), .B(new_n4164_), .ZN(new_n4359_));
  NOR3_X1    g04103(.A1(new_n4359_), .A2(new_n4167_), .A3(new_n4355_), .ZN(new_n4360_));
  NOR3_X1    g04104(.A1(new_n4360_), .A2(new_n4358_), .A3(new_n4351_), .ZN(new_n4361_));
  INV_X1     g04105(.I(new_n4348_), .ZN(new_n4362_));
  NOR2_X1    g04106(.A1(new_n4362_), .A2(new_n4349_), .ZN(new_n4363_));
  OAI21_X1   g04107(.A1(new_n4359_), .A2(new_n4167_), .B(new_n4355_), .ZN(new_n4364_));
  NAND3_X1   g04108(.A1(new_n4357_), .A2(new_n4159_), .A3(new_n4356_), .ZN(new_n4365_));
  AOI21_X1   g04109(.A1(new_n4364_), .A2(new_n4365_), .B(new_n4363_), .ZN(new_n4366_));
  NOR2_X1    g04110(.A1(new_n4361_), .A2(new_n4366_), .ZN(new_n4367_));
  INV_X1     g04111(.I(new_n4179_), .ZN(new_n4368_));
  OAI22_X1   g04112(.A1(new_n610_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n612_), .ZN(new_n4369_));
  AOI21_X1   g04113(.A1(\b[25] ), .A2(new_n826_), .B(new_n4369_), .ZN(new_n4370_));
  OAI21_X1   g04114(.A1(new_n3165_), .A2(new_n624_), .B(new_n4370_), .ZN(new_n4371_));
  XOR2_X1    g04115(.A1(new_n4371_), .A2(\a[8] ), .Z(new_n4372_));
  OAI21_X1   g04116(.A1(new_n4181_), .A2(new_n4368_), .B(new_n4372_), .ZN(new_n4373_));
  INV_X1     g04117(.I(new_n4372_), .ZN(new_n4374_));
  OAI21_X1   g04118(.A1(new_n4003_), .A2(new_n3990_), .B(new_n3985_), .ZN(new_n4375_));
  AOI21_X1   g04119(.A1(new_n4375_), .A2(new_n4176_), .B(new_n4368_), .ZN(new_n4376_));
  NAND2_X1   g04120(.A1(new_n4376_), .A2(new_n4374_), .ZN(new_n4377_));
  NAND3_X1   g04121(.A1(new_n4377_), .A2(new_n4373_), .A3(new_n4367_), .ZN(new_n4378_));
  AOI21_X1   g04122(.A1(new_n4377_), .A2(new_n4373_), .B(new_n4367_), .ZN(new_n4379_));
  INV_X1     g04123(.I(new_n4379_), .ZN(new_n4380_));
  AOI21_X1   g04124(.A1(new_n4380_), .A2(new_n4378_), .B(new_n4234_), .ZN(new_n4381_));
  INV_X1     g04125(.I(new_n4234_), .ZN(new_n4382_));
  OR2_X2     g04126(.A1(new_n4361_), .A2(new_n4366_), .Z(new_n4383_));
  INV_X1     g04127(.I(new_n4373_), .ZN(new_n4384_));
  NOR3_X1    g04128(.A1(new_n4181_), .A2(new_n4368_), .A3(new_n4372_), .ZN(new_n4385_));
  NOR3_X1    g04129(.A1(new_n4384_), .A2(new_n4385_), .A3(new_n4383_), .ZN(new_n4386_));
  NOR3_X1    g04130(.A1(new_n4386_), .A2(new_n4379_), .A3(new_n4382_), .ZN(new_n4387_));
  OAI21_X1   g04131(.A1(new_n4381_), .A2(new_n4387_), .B(new_n4229_), .ZN(new_n4388_));
  OAI21_X1   g04132(.A1(new_n4200_), .A2(new_n4196_), .B(new_n4202_), .ZN(new_n4389_));
  OAI21_X1   g04133(.A1(new_n4386_), .A2(new_n4379_), .B(new_n4382_), .ZN(new_n4390_));
  NAND3_X1   g04134(.A1(new_n4380_), .A2(new_n4378_), .A3(new_n4234_), .ZN(new_n4391_));
  NAND3_X1   g04135(.A1(new_n4389_), .A2(new_n4390_), .A3(new_n4391_), .ZN(new_n4392_));
  NAND2_X1   g04136(.A1(new_n4392_), .A2(new_n4388_), .ZN(new_n4393_));
  NAND2_X1   g04137(.A1(new_n4393_), .A2(new_n4228_), .ZN(new_n4394_));
  INV_X1     g04138(.I(new_n4394_), .ZN(new_n4395_));
  NOR2_X1    g04139(.A1(new_n4393_), .A2(new_n4228_), .ZN(new_n4396_));
  NOR2_X1    g04140(.A1(new_n4395_), .A2(new_n4396_), .ZN(new_n4397_));
  XOR2_X1    g04141(.A1(new_n4397_), .A2(new_n4210_), .Z(\f[33] ));
  OAI21_X1   g04142(.A1(new_n4229_), .A2(new_n4387_), .B(new_n4390_), .ZN(new_n4399_));
  OAI21_X1   g04143(.A1(new_n3750_), .A2(new_n3739_), .B(new_n3752_), .ZN(new_n4400_));
  OAI21_X1   g04144(.A1(new_n4400_), .A2(new_n3983_), .B(new_n4166_), .ZN(new_n4401_));
  AOI21_X1   g04145(.A1(new_n4401_), .A2(new_n4169_), .B(new_n4167_), .ZN(new_n4402_));
  OAI21_X1   g04146(.A1(new_n4402_), .A2(new_n4356_), .B(new_n4351_), .ZN(new_n4403_));
  OAI22_X1   g04147(.A1(new_n713_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n717_), .ZN(new_n4404_));
  AOI21_X1   g04148(.A1(\b[23] ), .A2(new_n1126_), .B(new_n4404_), .ZN(new_n4405_));
  OAI21_X1   g04149(.A1(new_n2655_), .A2(new_n986_), .B(new_n4405_), .ZN(new_n4406_));
  XOR2_X1    g04150(.A1(new_n4406_), .A2(\a[11] ), .Z(new_n4407_));
  INV_X1     g04151(.I(new_n4337_), .ZN(new_n4408_));
  NAND2_X1   g04152(.A1(new_n4408_), .A2(new_n4338_), .ZN(new_n4409_));
  AOI21_X1   g04153(.A1(new_n3722_), .A2(new_n3533_), .B(new_n3723_), .ZN(new_n4410_));
  OAI21_X1   g04154(.A1(new_n3716_), .A2(new_n4410_), .B(new_n3724_), .ZN(new_n4411_));
  OAI21_X1   g04155(.A1(new_n4411_), .A2(new_n3962_), .B(new_n3957_), .ZN(new_n4412_));
  AOI21_X1   g04156(.A1(new_n4412_), .A2(new_n4153_), .B(new_n4149_), .ZN(new_n4413_));
  OAI21_X1   g04157(.A1(new_n4413_), .A2(new_n4346_), .B(new_n4409_), .ZN(new_n4414_));
  OAI22_X1   g04158(.A1(new_n993_), .A2(new_n2142_), .B1(new_n2027_), .B2(new_n997_), .ZN(new_n4415_));
  AOI21_X1   g04159(.A1(\b[20] ), .A2(new_n1486_), .B(new_n4415_), .ZN(new_n4416_));
  OAI21_X1   g04160(.A1(new_n2153_), .A2(new_n1323_), .B(new_n4416_), .ZN(new_n4417_));
  XOR2_X1    g04161(.A1(new_n4417_), .A2(\a[14] ), .Z(new_n4418_));
  INV_X1     g04162(.I(new_n4418_), .ZN(new_n4419_));
  INV_X1     g04163(.I(new_n4326_), .ZN(new_n4420_));
  NOR2_X1    g04164(.A1(new_n4420_), .A2(new_n4327_), .ZN(new_n4421_));
  AOI21_X1   g04165(.A1(new_n3707_), .A2(new_n3712_), .B(new_n3948_), .ZN(new_n4422_));
  AOI21_X1   g04166(.A1(new_n4422_), .A2(new_n3946_), .B(new_n4142_), .ZN(new_n4423_));
  OAI21_X1   g04167(.A1(new_n4423_), .A2(new_n4141_), .B(new_n4140_), .ZN(new_n4424_));
  AOI21_X1   g04168(.A1(new_n4424_), .A2(new_n4333_), .B(new_n4421_), .ZN(new_n4425_));
  OAI22_X1   g04169(.A1(new_n1592_), .A2(new_n1859_), .B1(new_n1553_), .B2(new_n1505_), .ZN(new_n4426_));
  AOI21_X1   g04170(.A1(\b[17] ), .A2(new_n1584_), .B(new_n4426_), .ZN(new_n4427_));
  NAND2_X1   g04171(.A1(new_n1695_), .A2(new_n1354_), .ZN(new_n4428_));
  NAND2_X1   g04172(.A1(new_n4428_), .A2(new_n4427_), .ZN(new_n4429_));
  NAND2_X1   g04173(.A1(new_n4429_), .A2(\a[17] ), .ZN(new_n4430_));
  NAND3_X1   g04174(.A1(new_n4428_), .A2(new_n1344_), .A3(new_n4427_), .ZN(new_n4431_));
  NAND2_X1   g04175(.A1(new_n4430_), .A2(new_n4431_), .ZN(new_n4432_));
  NAND2_X1   g04176(.A1(new_n4312_), .A2(new_n4292_), .ZN(new_n4433_));
  AOI21_X1   g04177(.A1(new_n4280_), .A2(new_n4275_), .B(new_n4285_), .ZN(new_n4434_));
  AOI21_X1   g04178(.A1(new_n4253_), .A2(new_n4256_), .B(new_n4258_), .ZN(new_n4435_));
  AOI21_X1   g04179(.A1(new_n4237_), .A2(new_n4262_), .B(new_n4435_), .ZN(new_n4436_));
  NOR2_X1    g04180(.A1(new_n4062_), .A2(new_n4248_), .ZN(new_n4437_));
  NAND2_X1   g04181(.A1(new_n4062_), .A2(new_n4248_), .ZN(new_n4438_));
  OAI21_X1   g04182(.A1(new_n4251_), .A2(new_n4437_), .B(new_n4438_), .ZN(new_n4439_));
  INV_X1     g04183(.I(new_n4439_), .ZN(new_n4440_));
  AOI22_X1   g04184(.A1(new_n3864_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n3869_), .ZN(new_n4441_));
  NAND2_X1   g04185(.A1(new_n4053_), .A2(\b[2] ), .ZN(new_n4442_));
  NAND2_X1   g04186(.A1(new_n1725_), .A2(new_n3872_), .ZN(new_n4443_));
  NAND3_X1   g04187(.A1(new_n4443_), .A2(new_n4441_), .A3(new_n4442_), .ZN(new_n4444_));
  XOR2_X1    g04188(.A1(new_n4444_), .A2(\a[32] ), .Z(new_n4445_));
  INV_X1     g04189(.I(\a[35] ), .ZN(new_n4446_));
  XOR2_X1    g04190(.A1(\a[32] ), .A2(\a[33] ), .Z(new_n4447_));
  XNOR2_X1   g04191(.A1(\a[34] ), .A2(\a[35] ), .ZN(new_n4448_));
  NAND2_X1   g04192(.A1(new_n4448_), .A2(new_n4447_), .ZN(new_n4449_));
  INV_X1     g04193(.I(\a[34] ), .ZN(new_n4450_));
  NOR3_X1    g04194(.A1(new_n4450_), .A2(\a[32] ), .A3(\a[33] ), .ZN(new_n4451_));
  NAND3_X1   g04195(.A1(new_n4450_), .A2(\a[32] ), .A3(\a[33] ), .ZN(new_n4452_));
  INV_X1     g04196(.I(new_n4452_), .ZN(new_n4453_));
  NOR2_X1    g04197(.A1(new_n4453_), .A2(new_n4451_), .ZN(new_n4454_));
  OAI22_X1   g04198(.A1(new_n275_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n258_), .ZN(new_n4455_));
  NOR2_X1    g04199(.A1(new_n4446_), .A2(\a[34] ), .ZN(new_n4456_));
  NOR2_X1    g04200(.A1(new_n4450_), .A2(\a[35] ), .ZN(new_n4457_));
  OAI21_X1   g04201(.A1(new_n4456_), .A2(new_n4457_), .B(new_n4447_), .ZN(new_n4458_));
  NOR2_X1    g04202(.A1(new_n4458_), .A2(new_n313_), .ZN(new_n4459_));
  NOR2_X1    g04203(.A1(new_n4455_), .A2(new_n4459_), .ZN(new_n4460_));
  NOR2_X1    g04204(.A1(new_n4460_), .A2(new_n4446_), .ZN(new_n4461_));
  NAND2_X1   g04205(.A1(new_n4460_), .A2(new_n4446_), .ZN(new_n4462_));
  INV_X1     g04206(.I(new_n4462_), .ZN(new_n4463_));
  NOR2_X1    g04207(.A1(new_n4248_), .A2(new_n4446_), .ZN(new_n4464_));
  NOR3_X1    g04208(.A1(new_n4463_), .A2(new_n4461_), .A3(new_n4464_), .ZN(new_n4465_));
  NAND2_X1   g04209(.A1(new_n4461_), .A2(new_n4249_), .ZN(new_n4466_));
  INV_X1     g04210(.I(new_n4466_), .ZN(new_n4467_));
  OAI21_X1   g04211(.A1(new_n4465_), .A2(new_n4467_), .B(new_n4445_), .ZN(new_n4468_));
  XOR2_X1    g04212(.A1(new_n4444_), .A2(new_n3876_), .Z(new_n4469_));
  INV_X1     g04213(.I(new_n4461_), .ZN(new_n4470_));
  INV_X1     g04214(.I(new_n4464_), .ZN(new_n4471_));
  NAND3_X1   g04215(.A1(new_n4470_), .A2(new_n4462_), .A3(new_n4471_), .ZN(new_n4472_));
  NAND3_X1   g04216(.A1(new_n4472_), .A2(new_n4469_), .A3(new_n4466_), .ZN(new_n4473_));
  AOI21_X1   g04217(.A1(new_n4468_), .A2(new_n4473_), .B(new_n4440_), .ZN(new_n4474_));
  AOI21_X1   g04218(.A1(new_n4472_), .A2(new_n4466_), .B(new_n4469_), .ZN(new_n4475_));
  NOR3_X1    g04219(.A1(new_n4465_), .A2(new_n4445_), .A3(new_n4467_), .ZN(new_n4476_));
  NOR3_X1    g04220(.A1(new_n4475_), .A2(new_n4476_), .A3(new_n4439_), .ZN(new_n4477_));
  NOR2_X1    g04221(.A1(new_n4474_), .A2(new_n4477_), .ZN(new_n4478_));
  OAI22_X1   g04222(.A1(new_n471_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n438_), .ZN(new_n4479_));
  AOI21_X1   g04223(.A1(\b[5] ), .A2(new_n3456_), .B(new_n4479_), .ZN(new_n4480_));
  OAI21_X1   g04224(.A1(new_n485_), .A2(new_n3261_), .B(new_n4480_), .ZN(new_n4481_));
  XOR2_X1    g04225(.A1(new_n4481_), .A2(\a[29] ), .Z(new_n4482_));
  INV_X1     g04226(.I(new_n4482_), .ZN(new_n4483_));
  NAND2_X1   g04227(.A1(new_n4478_), .A2(new_n4483_), .ZN(new_n4484_));
  OAI21_X1   g04228(.A1(new_n4475_), .A2(new_n4476_), .B(new_n4439_), .ZN(new_n4485_));
  NAND3_X1   g04229(.A1(new_n4440_), .A2(new_n4468_), .A3(new_n4473_), .ZN(new_n4486_));
  NAND2_X1   g04230(.A1(new_n4486_), .A2(new_n4485_), .ZN(new_n4487_));
  NAND2_X1   g04231(.A1(new_n4487_), .A2(new_n4482_), .ZN(new_n4488_));
  AOI21_X1   g04232(.A1(new_n4484_), .A2(new_n4488_), .B(new_n4436_), .ZN(new_n4489_));
  INV_X1     g04233(.I(new_n4435_), .ZN(new_n4490_));
  OAI21_X1   g04234(.A1(new_n4269_), .A2(new_n4266_), .B(new_n4490_), .ZN(new_n4491_));
  NAND2_X1   g04235(.A1(new_n4484_), .A2(new_n4488_), .ZN(new_n4492_));
  NOR2_X1    g04236(.A1(new_n4492_), .A2(new_n4491_), .ZN(new_n4493_));
  AOI22_X1   g04237(.A1(new_n2716_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n2719_), .ZN(new_n4494_));
  OAI21_X1   g04238(.A1(new_n577_), .A2(new_n2924_), .B(new_n4494_), .ZN(new_n4495_));
  AOI21_X1   g04239(.A1(new_n1059_), .A2(new_n2722_), .B(new_n4495_), .ZN(new_n4496_));
  XOR2_X1    g04240(.A1(new_n4496_), .A2(new_n2714_), .Z(new_n4497_));
  NOR3_X1    g04241(.A1(new_n4489_), .A2(new_n4493_), .A3(new_n4497_), .ZN(new_n4498_));
  NAND2_X1   g04242(.A1(new_n4492_), .A2(new_n4491_), .ZN(new_n4499_));
  NAND3_X1   g04243(.A1(new_n4436_), .A2(new_n4484_), .A3(new_n4488_), .ZN(new_n4500_));
  XOR2_X1    g04244(.A1(new_n4496_), .A2(\a[26] ), .Z(new_n4501_));
  AOI21_X1   g04245(.A1(new_n4499_), .A2(new_n4500_), .B(new_n4501_), .ZN(new_n4502_));
  NOR2_X1    g04246(.A1(new_n4498_), .A2(new_n4502_), .ZN(new_n4503_));
  NOR3_X1    g04247(.A1(new_n4503_), .A2(new_n4283_), .A3(new_n4434_), .ZN(new_n4504_));
  OAI21_X1   g04248(.A1(new_n4288_), .A2(new_n4286_), .B(new_n4271_), .ZN(new_n4505_));
  NAND3_X1   g04249(.A1(new_n4499_), .A2(new_n4500_), .A3(new_n4501_), .ZN(new_n4506_));
  OAI21_X1   g04250(.A1(new_n4489_), .A2(new_n4493_), .B(new_n4497_), .ZN(new_n4507_));
  NAND2_X1   g04251(.A1(new_n4507_), .A2(new_n4506_), .ZN(new_n4508_));
  AOI21_X1   g04252(.A1(new_n4505_), .A2(new_n4289_), .B(new_n4508_), .ZN(new_n4509_));
  AOI22_X1   g04253(.A1(new_n2202_), .A2(\b[13] ), .B1(\b[12] ), .B2(new_n2205_), .ZN(new_n4510_));
  OAI21_X1   g04254(.A1(new_n852_), .A2(new_n2370_), .B(new_n4510_), .ZN(new_n4511_));
  INV_X1     g04255(.I(new_n4511_), .ZN(new_n4512_));
  OAI21_X1   g04256(.A1(new_n1082_), .A2(new_n2197_), .B(new_n4512_), .ZN(new_n4513_));
  XOR2_X1    g04257(.A1(new_n4513_), .A2(\a[23] ), .Z(new_n4514_));
  NOR3_X1    g04258(.A1(new_n4514_), .A2(new_n4509_), .A3(new_n4504_), .ZN(new_n4515_));
  NAND3_X1   g04259(.A1(new_n4505_), .A2(new_n4508_), .A3(new_n4289_), .ZN(new_n4516_));
  OAI21_X1   g04260(.A1(new_n4283_), .A2(new_n4434_), .B(new_n4503_), .ZN(new_n4517_));
  XOR2_X1    g04261(.A1(new_n4513_), .A2(new_n2200_), .Z(new_n4518_));
  AOI21_X1   g04262(.A1(new_n4517_), .A2(new_n4516_), .B(new_n4518_), .ZN(new_n4519_));
  NOR2_X1    g04263(.A1(new_n4519_), .A2(new_n4515_), .ZN(new_n4520_));
  AOI21_X1   g04264(.A1(new_n4313_), .A2(new_n4433_), .B(new_n4520_), .ZN(new_n4521_));
  AOI21_X1   g04265(.A1(new_n4307_), .A2(new_n4296_), .B(new_n4291_), .ZN(new_n4522_));
  NAND3_X1   g04266(.A1(new_n4518_), .A2(new_n4517_), .A3(new_n4516_), .ZN(new_n4523_));
  OAI21_X1   g04267(.A1(new_n4504_), .A2(new_n4509_), .B(new_n4514_), .ZN(new_n4524_));
  NAND2_X1   g04268(.A1(new_n4524_), .A2(new_n4523_), .ZN(new_n4525_));
  NOR3_X1    g04269(.A1(new_n4525_), .A2(new_n4522_), .A3(new_n4308_), .ZN(new_n4526_));
  AOI22_X1   g04270(.A1(new_n1738_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n1743_), .ZN(new_n4527_));
  OAI21_X1   g04271(.A1(new_n1093_), .A2(new_n1931_), .B(new_n4527_), .ZN(new_n4528_));
  AOI21_X1   g04272(.A1(new_n1701_), .A2(new_n1746_), .B(new_n4528_), .ZN(new_n4529_));
  XOR2_X1    g04273(.A1(new_n4529_), .A2(new_n1736_), .Z(new_n4530_));
  INV_X1     g04274(.I(new_n4530_), .ZN(new_n4531_));
  OAI21_X1   g04275(.A1(new_n4521_), .A2(new_n4526_), .B(new_n4531_), .ZN(new_n4532_));
  OAI21_X1   g04276(.A1(new_n4522_), .A2(new_n4308_), .B(new_n4525_), .ZN(new_n4533_));
  NAND3_X1   g04277(.A1(new_n4433_), .A2(new_n4520_), .A3(new_n4313_), .ZN(new_n4534_));
  NAND3_X1   g04278(.A1(new_n4533_), .A2(new_n4534_), .A3(new_n4530_), .ZN(new_n4535_));
  NAND2_X1   g04279(.A1(new_n4532_), .A2(new_n4535_), .ZN(new_n4536_));
  AOI21_X1   g04280(.A1(new_n4133_), .A2(new_n4132_), .B(new_n4322_), .ZN(new_n4537_));
  OAI22_X1   g04281(.A1(new_n4537_), .A2(new_n4324_), .B1(new_n4309_), .B2(new_n4314_), .ZN(new_n4538_));
  AOI21_X1   g04282(.A1(new_n4538_), .A2(new_n4325_), .B(new_n4536_), .ZN(new_n4539_));
  OAI21_X1   g04283(.A1(new_n3942_), .A2(new_n3928_), .B(new_n3937_), .ZN(new_n4540_));
  OAI21_X1   g04284(.A1(new_n4540_), .A2(new_n4127_), .B(new_n4321_), .ZN(new_n4541_));
  NOR2_X1    g04285(.A1(new_n4541_), .A2(new_n4319_), .ZN(new_n4542_));
  AOI21_X1   g04286(.A1(new_n4533_), .A2(new_n4534_), .B(new_n4530_), .ZN(new_n4543_));
  NOR3_X1    g04287(.A1(new_n4521_), .A2(new_n4526_), .A3(new_n4531_), .ZN(new_n4544_));
  NOR2_X1    g04288(.A1(new_n4544_), .A2(new_n4543_), .ZN(new_n4545_));
  AOI21_X1   g04289(.A1(new_n4541_), .A2(new_n4319_), .B(new_n4315_), .ZN(new_n4546_));
  NOR3_X1    g04290(.A1(new_n4546_), .A2(new_n4545_), .A3(new_n4542_), .ZN(new_n4547_));
  NOR3_X1    g04291(.A1(new_n4547_), .A2(new_n4539_), .A3(new_n4432_), .ZN(new_n4548_));
  INV_X1     g04292(.I(new_n4432_), .ZN(new_n4549_));
  OAI21_X1   g04293(.A1(new_n4546_), .A2(new_n4542_), .B(new_n4545_), .ZN(new_n4550_));
  NAND3_X1   g04294(.A1(new_n4538_), .A2(new_n4536_), .A3(new_n4325_), .ZN(new_n4551_));
  AOI21_X1   g04295(.A1(new_n4550_), .A2(new_n4551_), .B(new_n4549_), .ZN(new_n4552_));
  NOR2_X1    g04296(.A1(new_n4552_), .A2(new_n4548_), .ZN(new_n4553_));
  NOR3_X1    g04297(.A1(new_n4425_), .A2(new_n4336_), .A3(new_n4553_), .ZN(new_n4554_));
  NAND3_X1   g04298(.A1(new_n4150_), .A2(new_n4140_), .A3(new_n4334_), .ZN(new_n4555_));
  NAND2_X1   g04299(.A1(new_n3843_), .A2(new_n3714_), .ZN(new_n4556_));
  OAI21_X1   g04300(.A1(new_n4556_), .A2(new_n3955_), .B(new_n4143_), .ZN(new_n4557_));
  AOI21_X1   g04301(.A1(new_n4557_), .A2(new_n4147_), .B(new_n4146_), .ZN(new_n4558_));
  OAI21_X1   g04302(.A1(new_n4558_), .A2(new_n4334_), .B(new_n4329_), .ZN(new_n4559_));
  NAND3_X1   g04303(.A1(new_n4550_), .A2(new_n4551_), .A3(new_n4549_), .ZN(new_n4560_));
  OAI21_X1   g04304(.A1(new_n4547_), .A2(new_n4539_), .B(new_n4432_), .ZN(new_n4561_));
  NAND2_X1   g04305(.A1(new_n4561_), .A2(new_n4560_), .ZN(new_n4562_));
  AOI21_X1   g04306(.A1(new_n4559_), .A2(new_n4555_), .B(new_n4562_), .ZN(new_n4563_));
  NOR3_X1    g04307(.A1(new_n4563_), .A2(new_n4554_), .A3(new_n4419_), .ZN(new_n4564_));
  NAND3_X1   g04308(.A1(new_n4559_), .A2(new_n4555_), .A3(new_n4562_), .ZN(new_n4565_));
  OAI21_X1   g04309(.A1(new_n4425_), .A2(new_n4336_), .B(new_n4553_), .ZN(new_n4566_));
  AOI21_X1   g04310(.A1(new_n4565_), .A2(new_n4566_), .B(new_n4418_), .ZN(new_n4567_));
  NOR2_X1    g04311(.A1(new_n4567_), .A2(new_n4564_), .ZN(new_n4568_));
  NAND3_X1   g04312(.A1(new_n4414_), .A2(new_n4347_), .A3(new_n4568_), .ZN(new_n4569_));
  AOI21_X1   g04313(.A1(new_n4154_), .A2(new_n4155_), .B(new_n4346_), .ZN(new_n4570_));
  OAI21_X1   g04314(.A1(new_n4340_), .A2(new_n4570_), .B(new_n4347_), .ZN(new_n4571_));
  NAND3_X1   g04315(.A1(new_n4565_), .A2(new_n4566_), .A3(new_n4418_), .ZN(new_n4572_));
  OAI21_X1   g04316(.A1(new_n4563_), .A2(new_n4554_), .B(new_n4419_), .ZN(new_n4573_));
  NAND2_X1   g04317(.A1(new_n4573_), .A2(new_n4572_), .ZN(new_n4574_));
  NAND2_X1   g04318(.A1(new_n4571_), .A2(new_n4574_), .ZN(new_n4575_));
  AOI21_X1   g04319(.A1(new_n4575_), .A2(new_n4569_), .B(new_n4407_), .ZN(new_n4576_));
  INV_X1     g04320(.I(new_n4407_), .ZN(new_n4577_));
  NOR3_X1    g04321(.A1(new_n4161_), .A2(new_n4149_), .A3(new_n4344_), .ZN(new_n4578_));
  AOI21_X1   g04322(.A1(new_n3747_), .A2(new_n3721_), .B(new_n3830_), .ZN(new_n4579_));
  AOI21_X1   g04323(.A1(new_n4579_), .A2(new_n3970_), .B(new_n3968_), .ZN(new_n4580_));
  OAI21_X1   g04324(.A1(new_n4580_), .A2(new_n4157_), .B(new_n4155_), .ZN(new_n4581_));
  AOI21_X1   g04325(.A1(new_n4581_), .A2(new_n4344_), .B(new_n4340_), .ZN(new_n4582_));
  NOR3_X1    g04326(.A1(new_n4582_), .A2(new_n4578_), .A3(new_n4574_), .ZN(new_n4583_));
  AOI21_X1   g04327(.A1(new_n4409_), .A2(new_n4345_), .B(new_n4578_), .ZN(new_n4584_));
  NOR2_X1    g04328(.A1(new_n4584_), .A2(new_n4568_), .ZN(new_n4585_));
  NOR3_X1    g04329(.A1(new_n4585_), .A2(new_n4577_), .A3(new_n4583_), .ZN(new_n4586_));
  NOR2_X1    g04330(.A1(new_n4576_), .A2(new_n4586_), .ZN(new_n4587_));
  NAND3_X1   g04331(.A1(new_n4587_), .A2(new_n4403_), .A3(new_n4365_), .ZN(new_n4588_));
  AOI21_X1   g04332(.A1(new_n3726_), .A2(new_n3751_), .B(new_n3743_), .ZN(new_n4589_));
  AOI21_X1   g04333(.A1(new_n4589_), .A2(new_n3977_), .B(new_n4034_), .ZN(new_n4590_));
  OAI21_X1   g04334(.A1(new_n4590_), .A2(new_n4164_), .B(new_n4159_), .ZN(new_n4591_));
  AOI21_X1   g04335(.A1(new_n4591_), .A2(new_n4355_), .B(new_n4363_), .ZN(new_n4592_));
  OAI22_X1   g04336(.A1(new_n4592_), .A2(new_n4360_), .B1(new_n4576_), .B2(new_n4586_), .ZN(new_n4593_));
  AOI22_X1   g04337(.A1(new_n518_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n636_), .ZN(new_n4594_));
  OAI21_X1   g04338(.A1(new_n3006_), .A2(new_n917_), .B(new_n4594_), .ZN(new_n4595_));
  AOI21_X1   g04339(.A1(new_n3807_), .A2(new_n618_), .B(new_n4595_), .ZN(new_n4596_));
  XOR2_X1    g04340(.A1(new_n4596_), .A2(new_n488_), .Z(new_n4597_));
  AOI21_X1   g04341(.A1(new_n4593_), .A2(new_n4588_), .B(new_n4597_), .ZN(new_n4598_));
  NAND3_X1   g04342(.A1(new_n4593_), .A2(new_n4588_), .A3(new_n4597_), .ZN(new_n4599_));
  INV_X1     g04343(.I(new_n4599_), .ZN(new_n4600_));
  NOR2_X1    g04344(.A1(new_n4600_), .A2(new_n4598_), .ZN(new_n4601_));
  OAI21_X1   g04345(.A1(new_n4184_), .A2(new_n4180_), .B(new_n4179_), .ZN(new_n4602_));
  AOI21_X1   g04346(.A1(new_n4602_), .A2(new_n4372_), .B(new_n4367_), .ZN(new_n4603_));
  OAI21_X1   g04347(.A1(new_n4385_), .A2(new_n4603_), .B(new_n4601_), .ZN(new_n4604_));
  INV_X1     g04348(.I(new_n4588_), .ZN(new_n4605_));
  AOI21_X1   g04349(.A1(new_n4351_), .A2(new_n4364_), .B(new_n4360_), .ZN(new_n4606_));
  NOR2_X1    g04350(.A1(new_n4606_), .A2(new_n4587_), .ZN(new_n4607_));
  INV_X1     g04351(.I(new_n4597_), .ZN(new_n4608_));
  OAI21_X1   g04352(.A1(new_n4605_), .A2(new_n4607_), .B(new_n4608_), .ZN(new_n4609_));
  NAND2_X1   g04353(.A1(new_n4609_), .A2(new_n4599_), .ZN(new_n4610_));
  OAI21_X1   g04354(.A1(new_n4376_), .A2(new_n4374_), .B(new_n4383_), .ZN(new_n4611_));
  NAND3_X1   g04355(.A1(new_n4610_), .A2(new_n4611_), .A3(new_n4377_), .ZN(new_n4612_));
  AOI22_X1   g04356(.A1(new_n800_), .A2(\b[30] ), .B1(\b[31] ), .B2(new_n333_), .ZN(new_n4613_));
  OAI21_X1   g04357(.A1(new_n3592_), .A2(new_n392_), .B(new_n4613_), .ZN(new_n4614_));
  INV_X1     g04358(.I(new_n4614_), .ZN(new_n4615_));
  NAND2_X1   g04359(.A1(new_n3795_), .A2(\b[31] ), .ZN(new_n4616_));
  NOR2_X1    g04360(.A1(new_n3792_), .A2(new_n3624_), .ZN(new_n4617_));
  AOI21_X1   g04361(.A1(new_n3624_), .A2(new_n3793_), .B(new_n4617_), .ZN(new_n4618_));
  NAND2_X1   g04362(.A1(new_n4618_), .A2(new_n4022_), .ZN(new_n4619_));
  NAND3_X1   g04363(.A1(new_n4619_), .A2(new_n4616_), .A3(new_n330_), .ZN(new_n4620_));
  AOI21_X1   g04364(.A1(new_n4620_), .A2(new_n4615_), .B(new_n312_), .ZN(new_n4621_));
  INV_X1     g04365(.I(new_n4621_), .ZN(new_n4622_));
  NAND3_X1   g04366(.A1(new_n4620_), .A2(new_n312_), .A3(new_n4615_), .ZN(new_n4623_));
  NAND2_X1   g04367(.A1(new_n4622_), .A2(new_n4623_), .ZN(new_n4624_));
  AOI21_X1   g04368(.A1(new_n4604_), .A2(new_n4612_), .B(new_n4624_), .ZN(new_n4625_));
  AOI21_X1   g04369(.A1(new_n4383_), .A2(new_n4373_), .B(new_n4385_), .ZN(new_n4626_));
  NOR2_X1    g04370(.A1(new_n4626_), .A2(new_n4610_), .ZN(new_n4627_));
  NOR3_X1    g04371(.A1(new_n4601_), .A2(new_n4603_), .A3(new_n4385_), .ZN(new_n4628_));
  INV_X1     g04372(.I(new_n4623_), .ZN(new_n4629_));
  NOR2_X1    g04373(.A1(new_n4629_), .A2(new_n4621_), .ZN(new_n4630_));
  NOR3_X1    g04374(.A1(new_n4627_), .A2(new_n4628_), .A3(new_n4630_), .ZN(new_n4631_));
  OAI21_X1   g04375(.A1(new_n4625_), .A2(new_n4631_), .B(new_n4399_), .ZN(new_n4632_));
  AOI21_X1   g04376(.A1(new_n4389_), .A2(new_n4391_), .B(new_n4381_), .ZN(new_n4633_));
  NOR2_X1    g04377(.A1(new_n4625_), .A2(new_n4631_), .ZN(new_n4634_));
  NAND2_X1   g04378(.A1(new_n4633_), .A2(new_n4634_), .ZN(new_n4635_));
  NAND2_X1   g04379(.A1(new_n4632_), .A2(new_n4635_), .ZN(new_n4636_));
  INV_X1     g04380(.I(new_n4636_), .ZN(new_n4637_));
  INV_X1     g04381(.I(\b[33] ), .ZN(new_n4638_));
  INV_X1     g04382(.I(\b[34] ), .ZN(new_n4639_));
  OAI22_X1   g04383(.A1(new_n277_), .A2(new_n4639_), .B1(new_n4638_), .B2(new_n262_), .ZN(new_n4640_));
  AOI21_X1   g04384(.A1(\b[32] ), .A2(new_n283_), .B(new_n4640_), .ZN(new_n4641_));
  OAI21_X1   g04385(.A1(new_n4217_), .A2(new_n4023_), .B(new_n4022_), .ZN(new_n4642_));
  NAND2_X1   g04386(.A1(new_n4219_), .A2(new_n4023_), .ZN(new_n4643_));
  NAND2_X1   g04387(.A1(new_n4642_), .A2(new_n4643_), .ZN(new_n4644_));
  XNOR2_X1   g04388(.A1(\b[33] ), .A2(\b[34] ), .ZN(new_n4645_));
  INV_X1     g04389(.I(new_n4645_), .ZN(new_n4646_));
  XOR2_X1    g04390(.A1(\b[33] ), .A2(\b[34] ), .Z(new_n4647_));
  NOR2_X1    g04391(.A1(new_n4644_), .A2(new_n4647_), .ZN(new_n4648_));
  AOI21_X1   g04392(.A1(new_n4644_), .A2(new_n4646_), .B(new_n4648_), .ZN(new_n4649_));
  OAI21_X1   g04393(.A1(new_n4649_), .A2(new_n279_), .B(new_n4641_), .ZN(new_n4650_));
  XOR2_X1    g04394(.A1(new_n4650_), .A2(\a[2] ), .Z(new_n4651_));
  INV_X1     g04395(.I(new_n4651_), .ZN(new_n4652_));
  INV_X1     g04396(.I(new_n4396_), .ZN(new_n4653_));
  AOI21_X1   g04397(.A1(new_n4210_), .A2(new_n4653_), .B(new_n4395_), .ZN(new_n4654_));
  NOR2_X1    g04398(.A1(new_n4654_), .A2(new_n4652_), .ZN(new_n4655_));
  NOR3_X1    g04399(.A1(new_n3785_), .A2(new_n3802_), .A3(new_n4016_), .ZN(new_n4656_));
  AOI21_X1   g04400(.A1(new_n3800_), .A2(new_n4017_), .B(new_n4656_), .ZN(new_n4657_));
  INV_X1     g04401(.I(new_n4207_), .ZN(new_n4658_));
  OAI21_X1   g04402(.A1(new_n4657_), .A2(new_n4658_), .B(new_n4206_), .ZN(new_n4659_));
  OAI21_X1   g04403(.A1(new_n4659_), .A2(new_n4396_), .B(new_n4394_), .ZN(new_n4660_));
  NOR2_X1    g04404(.A1(new_n4660_), .A2(new_n4651_), .ZN(new_n4661_));
  NOR2_X1    g04405(.A1(new_n4661_), .A2(new_n4655_), .ZN(new_n4662_));
  XOR2_X1    g04406(.A1(new_n4662_), .A2(new_n4637_), .Z(\f[34] ));
  AOI21_X1   g04407(.A1(new_n4660_), .A2(new_n4651_), .B(new_n4637_), .ZN(new_n4664_));
  NOR2_X1    g04408(.A1(new_n4664_), .A2(new_n4661_), .ZN(new_n4665_));
  INV_X1     g04409(.I(\b[35] ), .ZN(new_n4666_));
  OAI22_X1   g04410(.A1(new_n277_), .A2(new_n4666_), .B1(new_n4639_), .B2(new_n262_), .ZN(new_n4667_));
  AOI21_X1   g04411(.A1(\b[33] ), .A2(new_n283_), .B(new_n4667_), .ZN(new_n4668_));
  NAND2_X1   g04412(.A1(new_n4644_), .A2(new_n4638_), .ZN(new_n4669_));
  NOR2_X1    g04413(.A1(new_n4669_), .A2(new_n4639_), .ZN(new_n4670_));
  NAND3_X1   g04414(.A1(new_n4642_), .A2(new_n4643_), .A3(\b[33] ), .ZN(new_n4671_));
  NOR2_X1    g04415(.A1(new_n4671_), .A2(\b[34] ), .ZN(new_n4672_));
  OAI21_X1   g04416(.A1(new_n4670_), .A2(new_n4672_), .B(\b[35] ), .ZN(new_n4673_));
  NOR3_X1    g04417(.A1(new_n4670_), .A2(\b[35] ), .A3(new_n4672_), .ZN(new_n4674_));
  INV_X1     g04418(.I(new_n4674_), .ZN(new_n4675_));
  NAND2_X1   g04419(.A1(new_n4675_), .A2(new_n4673_), .ZN(new_n4676_));
  OAI21_X1   g04420(.A1(new_n4676_), .A2(new_n279_), .B(new_n4668_), .ZN(new_n4677_));
  XOR2_X1    g04421(.A1(new_n4677_), .A2(\a[2] ), .Z(new_n4678_));
  NOR3_X1    g04422(.A1(new_n4603_), .A2(new_n4385_), .A3(new_n4598_), .ZN(new_n4679_));
  AOI22_X1   g04423(.A1(new_n518_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n636_), .ZN(new_n4680_));
  OAI21_X1   g04424(.A1(new_n3158_), .A2(new_n917_), .B(new_n4680_), .ZN(new_n4681_));
  AOI21_X1   g04425(.A1(new_n4188_), .A2(new_n618_), .B(new_n4681_), .ZN(new_n4682_));
  XOR2_X1    g04426(.A1(new_n4682_), .A2(new_n488_), .Z(new_n4683_));
  AOI21_X1   g04427(.A1(new_n4403_), .A2(new_n4365_), .B(new_n4586_), .ZN(new_n4684_));
  OAI22_X1   g04428(.A1(new_n713_), .A2(new_n3006_), .B1(new_n2646_), .B2(new_n717_), .ZN(new_n4685_));
  AOI21_X1   g04429(.A1(\b[24] ), .A2(new_n1126_), .B(new_n4685_), .ZN(new_n4686_));
  OAI21_X1   g04430(.A1(new_n3016_), .A2(new_n986_), .B(new_n4686_), .ZN(new_n4687_));
  XOR2_X1    g04431(.A1(new_n4687_), .A2(\a[11] ), .Z(new_n4688_));
  INV_X1     g04432(.I(new_n4688_), .ZN(new_n4689_));
  AOI21_X1   g04433(.A1(new_n4550_), .A2(new_n4551_), .B(new_n4432_), .ZN(new_n4690_));
  NAND3_X1   g04434(.A1(new_n4538_), .A2(new_n4325_), .A3(new_n4532_), .ZN(new_n4691_));
  OAI22_X1   g04435(.A1(new_n1751_), .A2(new_n1432_), .B1(new_n1296_), .B2(new_n1754_), .ZN(new_n4692_));
  AOI21_X1   g04436(.A1(\b[15] ), .A2(new_n1939_), .B(new_n4692_), .ZN(new_n4693_));
  OAI21_X1   g04437(.A1(new_n1444_), .A2(new_n1757_), .B(new_n4693_), .ZN(new_n4694_));
  XOR2_X1    g04438(.A1(new_n4694_), .A2(\a[20] ), .Z(new_n4695_));
  INV_X1     g04439(.I(new_n4695_), .ZN(new_n4696_));
  NAND3_X1   g04440(.A1(new_n4433_), .A2(new_n4313_), .A3(new_n4523_), .ZN(new_n4697_));
  NOR2_X1    g04441(.A1(new_n4456_), .A2(new_n4457_), .ZN(new_n4698_));
  NOR2_X1    g04442(.A1(new_n4698_), .A2(new_n4247_), .ZN(new_n4699_));
  NAND2_X1   g04443(.A1(new_n4699_), .A2(new_n554_), .ZN(new_n4700_));
  NOR2_X1    g04444(.A1(new_n4449_), .A2(new_n276_), .ZN(new_n4701_));
  NOR2_X1    g04445(.A1(new_n4454_), .A2(new_n275_), .ZN(new_n4702_));
  NOR2_X1    g04446(.A1(new_n4701_), .A2(new_n4702_), .ZN(new_n4703_));
  NOR2_X1    g04447(.A1(new_n4456_), .A2(\a[32] ), .ZN(new_n4704_));
  NOR2_X1    g04448(.A1(new_n4457_), .A2(new_n3876_), .ZN(new_n4705_));
  NOR3_X1    g04449(.A1(new_n4704_), .A2(new_n4705_), .A3(new_n4447_), .ZN(new_n4706_));
  NAND2_X1   g04450(.A1(new_n4706_), .A2(\b[0] ), .ZN(new_n4707_));
  NAND3_X1   g04451(.A1(new_n4703_), .A2(new_n4700_), .A3(new_n4707_), .ZN(new_n4708_));
  XOR2_X1    g04452(.A1(new_n4708_), .A2(\a[35] ), .Z(new_n4709_));
  INV_X1     g04453(.I(new_n4460_), .ZN(new_n4710_));
  NOR3_X1    g04454(.A1(new_n4710_), .A2(new_n4446_), .A3(new_n4248_), .ZN(new_n4711_));
  NOR2_X1    g04455(.A1(new_n4709_), .A2(new_n4711_), .ZN(new_n4712_));
  INV_X1     g04456(.I(new_n4700_), .ZN(new_n4713_));
  INV_X1     g04457(.I(new_n4707_), .ZN(new_n4714_));
  NOR4_X1    g04458(.A1(new_n4714_), .A2(new_n4713_), .A3(new_n4701_), .A4(new_n4702_), .ZN(new_n4715_));
  NAND4_X1   g04459(.A1(new_n4715_), .A2(\a[35] ), .A3(new_n4249_), .A4(new_n4460_), .ZN(new_n4716_));
  INV_X1     g04460(.I(new_n4716_), .ZN(new_n4717_));
  NOR2_X1    g04461(.A1(new_n4712_), .A2(new_n4717_), .ZN(new_n4718_));
  OAI21_X1   g04462(.A1(new_n4440_), .A2(new_n4476_), .B(new_n4468_), .ZN(new_n4719_));
  NAND2_X1   g04463(.A1(new_n4719_), .A2(new_n4718_), .ZN(new_n4720_));
  XOR2_X1    g04464(.A1(new_n4708_), .A2(new_n4446_), .Z(new_n4721_));
  INV_X1     g04465(.I(new_n4711_), .ZN(new_n4722_));
  NAND2_X1   g04466(.A1(new_n4721_), .A2(new_n4722_), .ZN(new_n4723_));
  NAND2_X1   g04467(.A1(new_n4723_), .A2(new_n4716_), .ZN(new_n4724_));
  AOI21_X1   g04468(.A1(new_n4439_), .A2(new_n4473_), .B(new_n4475_), .ZN(new_n4725_));
  NAND2_X1   g04469(.A1(new_n4725_), .A2(new_n4724_), .ZN(new_n4726_));
  INV_X1     g04470(.I(new_n3872_), .ZN(new_n4727_));
  XNOR2_X1   g04471(.A1(\a[31] ), .A2(\a[32] ), .ZN(new_n4728_));
  NAND2_X1   g04472(.A1(new_n4728_), .A2(new_n4050_), .ZN(new_n4729_));
  INV_X1     g04473(.I(new_n3869_), .ZN(new_n4730_));
  OAI22_X1   g04474(.A1(new_n339_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n377_), .ZN(new_n4731_));
  AOI21_X1   g04475(.A1(\b[3] ), .A2(new_n4053_), .B(new_n4731_), .ZN(new_n4732_));
  OAI21_X1   g04476(.A1(new_n566_), .A2(new_n4727_), .B(new_n4732_), .ZN(new_n4733_));
  XOR2_X1    g04477(.A1(new_n4733_), .A2(new_n3876_), .Z(new_n4734_));
  AOI22_X1   g04478(.A1(new_n3267_), .A2(\b[8] ), .B1(\b[7] ), .B2(new_n3270_), .ZN(new_n4735_));
  OAI21_X1   g04479(.A1(new_n438_), .A2(new_n3475_), .B(new_n4735_), .ZN(new_n4736_));
  AOI21_X1   g04480(.A1(new_n799_), .A2(new_n3273_), .B(new_n4736_), .ZN(new_n4737_));
  XOR2_X1    g04481(.A1(new_n4737_), .A2(\a[29] ), .Z(new_n4738_));
  NAND2_X1   g04482(.A1(new_n4738_), .A2(new_n4734_), .ZN(new_n4739_));
  XOR2_X1    g04483(.A1(new_n4733_), .A2(\a[32] ), .Z(new_n4740_));
  OR2_X2     g04484(.A1(new_n4737_), .A2(new_n3264_), .Z(new_n4741_));
  NAND2_X1   g04485(.A1(new_n4737_), .A2(new_n3264_), .ZN(new_n4742_));
  NAND3_X1   g04486(.A1(new_n4741_), .A2(new_n4742_), .A3(new_n4740_), .ZN(new_n4743_));
  NAND4_X1   g04487(.A1(new_n4739_), .A2(new_n4720_), .A3(new_n4726_), .A4(new_n4743_), .ZN(new_n4744_));
  NOR2_X1    g04488(.A1(new_n4725_), .A2(new_n4724_), .ZN(new_n4745_));
  NOR2_X1    g04489(.A1(new_n4719_), .A2(new_n4718_), .ZN(new_n4746_));
  XOR2_X1    g04490(.A1(new_n4737_), .A2(new_n3264_), .Z(new_n4747_));
  NOR2_X1    g04491(.A1(new_n4747_), .A2(new_n4740_), .ZN(new_n4748_));
  NOR2_X1    g04492(.A1(new_n4738_), .A2(new_n4734_), .ZN(new_n4749_));
  OAI22_X1   g04493(.A1(new_n4748_), .A2(new_n4749_), .B1(new_n4745_), .B2(new_n4746_), .ZN(new_n4750_));
  NAND2_X1   g04494(.A1(new_n4750_), .A2(new_n4744_), .ZN(new_n4751_));
  NOR2_X1    g04495(.A1(new_n4487_), .A2(new_n4482_), .ZN(new_n4752_));
  OAI21_X1   g04496(.A1(new_n4436_), .A2(new_n4752_), .B(new_n4488_), .ZN(new_n4753_));
  NOR2_X1    g04497(.A1(new_n4751_), .A2(new_n4753_), .ZN(new_n4754_));
  NOR4_X1    g04498(.A1(new_n4748_), .A2(new_n4749_), .A3(new_n4745_), .A4(new_n4746_), .ZN(new_n4755_));
  AOI22_X1   g04499(.A1(new_n4739_), .A2(new_n4743_), .B1(new_n4720_), .B2(new_n4726_), .ZN(new_n4756_));
  NOR2_X1    g04500(.A1(new_n4755_), .A2(new_n4756_), .ZN(new_n4757_));
  NOR2_X1    g04501(.A1(new_n4478_), .A2(new_n4483_), .ZN(new_n4758_));
  AOI21_X1   g04502(.A1(new_n4491_), .A2(new_n4484_), .B(new_n4758_), .ZN(new_n4759_));
  NOR2_X1    g04503(.A1(new_n4757_), .A2(new_n4759_), .ZN(new_n4760_));
  OAI22_X1   g04504(.A1(new_n2703_), .A2(new_n852_), .B1(new_n776_), .B2(new_n2708_), .ZN(new_n4761_));
  AOI21_X1   g04505(.A1(\b[9] ), .A2(new_n2906_), .B(new_n4761_), .ZN(new_n4762_));
  OAI21_X1   g04506(.A1(new_n859_), .A2(new_n2711_), .B(new_n4762_), .ZN(new_n4763_));
  XOR2_X1    g04507(.A1(new_n4763_), .A2(\a[26] ), .Z(new_n4764_));
  NOR3_X1    g04508(.A1(new_n4760_), .A2(new_n4754_), .A3(new_n4764_), .ZN(new_n4765_));
  NAND2_X1   g04509(.A1(new_n4757_), .A2(new_n4759_), .ZN(new_n4766_));
  NAND2_X1   g04510(.A1(new_n4751_), .A2(new_n4753_), .ZN(new_n4767_));
  XOR2_X1    g04511(.A1(new_n4763_), .A2(new_n2714_), .Z(new_n4768_));
  AOI21_X1   g04512(.A1(new_n4766_), .A2(new_n4767_), .B(new_n4768_), .ZN(new_n4769_));
  NOR2_X1    g04513(.A1(new_n4769_), .A2(new_n4765_), .ZN(new_n4770_));
  OAI21_X1   g04514(.A1(new_n4434_), .A2(new_n4283_), .B(new_n4507_), .ZN(new_n4771_));
  NAND3_X1   g04515(.A1(new_n4770_), .A2(new_n4506_), .A3(new_n4771_), .ZN(new_n4772_));
  AOI21_X1   g04516(.A1(new_n4505_), .A2(new_n4289_), .B(new_n4502_), .ZN(new_n4773_));
  OAI22_X1   g04517(.A1(new_n4773_), .A2(new_n4498_), .B1(new_n4765_), .B2(new_n4769_), .ZN(new_n4774_));
  AOI22_X1   g04518(.A1(new_n2202_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n2205_), .ZN(new_n4775_));
  OAI21_X1   g04519(.A1(new_n941_), .A2(new_n2370_), .B(new_n4775_), .ZN(new_n4776_));
  AOI21_X1   g04520(.A1(new_n1449_), .A2(new_n2208_), .B(new_n4776_), .ZN(new_n4777_));
  XOR2_X1    g04521(.A1(new_n4777_), .A2(new_n2200_), .Z(new_n4778_));
  NAND3_X1   g04522(.A1(new_n4774_), .A2(new_n4772_), .A3(new_n4778_), .ZN(new_n4779_));
  NOR4_X1    g04523(.A1(new_n4773_), .A2(new_n4498_), .A3(new_n4765_), .A4(new_n4769_), .ZN(new_n4780_));
  AOI21_X1   g04524(.A1(new_n4506_), .A2(new_n4771_), .B(new_n4770_), .ZN(new_n4781_));
  XOR2_X1    g04525(.A1(new_n4777_), .A2(\a[23] ), .Z(new_n4782_));
  OAI21_X1   g04526(.A1(new_n4781_), .A2(new_n4780_), .B(new_n4782_), .ZN(new_n4783_));
  NAND2_X1   g04527(.A1(new_n4783_), .A2(new_n4779_), .ZN(new_n4784_));
  AOI21_X1   g04528(.A1(new_n4697_), .A2(new_n4524_), .B(new_n4784_), .ZN(new_n4785_));
  NOR3_X1    g04529(.A1(new_n4522_), .A2(new_n4308_), .A3(new_n4515_), .ZN(new_n4786_));
  NOR3_X1    g04530(.A1(new_n4781_), .A2(new_n4780_), .A3(new_n4782_), .ZN(new_n4787_));
  AOI21_X1   g04531(.A1(new_n4774_), .A2(new_n4772_), .B(new_n4778_), .ZN(new_n4788_));
  NOR2_X1    g04532(.A1(new_n4787_), .A2(new_n4788_), .ZN(new_n4789_));
  NOR3_X1    g04533(.A1(new_n4786_), .A2(new_n4789_), .A3(new_n4519_), .ZN(new_n4790_));
  NOR3_X1    g04534(.A1(new_n4696_), .A2(new_n4785_), .A3(new_n4790_), .ZN(new_n4791_));
  OAI21_X1   g04535(.A1(new_n4786_), .A2(new_n4519_), .B(new_n4789_), .ZN(new_n4792_));
  NAND3_X1   g04536(.A1(new_n4697_), .A2(new_n4784_), .A3(new_n4524_), .ZN(new_n4793_));
  AOI21_X1   g04537(.A1(new_n4793_), .A2(new_n4792_), .B(new_n4695_), .ZN(new_n4794_));
  NOR2_X1    g04538(.A1(new_n4791_), .A2(new_n4794_), .ZN(new_n4795_));
  AOI21_X1   g04539(.A1(new_n4691_), .A2(new_n4535_), .B(new_n4795_), .ZN(new_n4796_));
  NOR3_X1    g04540(.A1(new_n4546_), .A2(new_n4542_), .A3(new_n4543_), .ZN(new_n4797_));
  NAND3_X1   g04541(.A1(new_n4793_), .A2(new_n4792_), .A3(new_n4695_), .ZN(new_n4798_));
  OAI21_X1   g04542(.A1(new_n4785_), .A2(new_n4790_), .B(new_n4696_), .ZN(new_n4799_));
  NAND2_X1   g04543(.A1(new_n4799_), .A2(new_n4798_), .ZN(new_n4800_));
  NOR3_X1    g04544(.A1(new_n4797_), .A2(new_n4544_), .A3(new_n4800_), .ZN(new_n4801_));
  NOR2_X1    g04545(.A1(new_n4801_), .A2(new_n4796_), .ZN(new_n4802_));
  INV_X1     g04546(.I(new_n4802_), .ZN(new_n4803_));
  OAI21_X1   g04547(.A1(new_n4554_), .A2(new_n4690_), .B(new_n4803_), .ZN(new_n4804_));
  INV_X1     g04548(.I(new_n4690_), .ZN(new_n4805_));
  NAND3_X1   g04549(.A1(new_n4565_), .A2(new_n4805_), .A3(new_n4802_), .ZN(new_n4806_));
  AOI22_X1   g04550(.A1(new_n1006_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n1009_), .ZN(new_n4807_));
  OAI21_X1   g04551(.A1(new_n2027_), .A2(new_n1481_), .B(new_n4807_), .ZN(new_n4808_));
  INV_X1     g04552(.I(new_n4808_), .ZN(new_n4809_));
  OAI21_X1   g04553(.A1(new_n3552_), .A2(new_n1323_), .B(new_n4809_), .ZN(new_n4810_));
  NAND2_X1   g04554(.A1(new_n4810_), .A2(\a[14] ), .ZN(new_n4811_));
  AOI21_X1   g04555(.A1(new_n2470_), .A2(new_n1013_), .B(new_n4808_), .ZN(new_n4812_));
  NAND2_X1   g04556(.A1(new_n4812_), .A2(new_n1002_), .ZN(new_n4813_));
  OAI22_X1   g04557(.A1(new_n1592_), .A2(new_n1860_), .B1(new_n1859_), .B2(new_n1505_), .ZN(new_n4814_));
  AOI21_X1   g04558(.A1(\b[18] ), .A2(new_n1584_), .B(new_n4814_), .ZN(new_n4815_));
  OAI21_X1   g04559(.A1(new_n1871_), .A2(new_n1732_), .B(new_n4815_), .ZN(new_n4816_));
  XOR2_X1    g04560(.A1(new_n4816_), .A2(\a[17] ), .Z(new_n4817_));
  INV_X1     g04561(.I(new_n4817_), .ZN(new_n4818_));
  AOI21_X1   g04562(.A1(new_n4813_), .A2(new_n4811_), .B(new_n4818_), .ZN(new_n4819_));
  NOR2_X1    g04563(.A1(new_n4812_), .A2(new_n1002_), .ZN(new_n4820_));
  NOR2_X1    g04564(.A1(new_n4810_), .A2(\a[14] ), .ZN(new_n4821_));
  NOR3_X1    g04565(.A1(new_n4820_), .A2(new_n4821_), .A3(new_n4817_), .ZN(new_n4822_));
  NOR2_X1    g04566(.A1(new_n4819_), .A2(new_n4822_), .ZN(new_n4823_));
  AOI21_X1   g04567(.A1(new_n4804_), .A2(new_n4806_), .B(new_n4823_), .ZN(new_n4824_));
  AOI21_X1   g04568(.A1(new_n4565_), .A2(new_n4805_), .B(new_n4802_), .ZN(new_n4825_));
  NOR3_X1    g04569(.A1(new_n4554_), .A2(new_n4690_), .A3(new_n4803_), .ZN(new_n4826_));
  OR2_X2     g04570(.A1(new_n4819_), .A2(new_n4822_), .Z(new_n4827_));
  NOR3_X1    g04571(.A1(new_n4825_), .A2(new_n4827_), .A3(new_n4826_), .ZN(new_n4828_));
  NOR2_X1    g04572(.A1(new_n4828_), .A2(new_n4824_), .ZN(new_n4829_));
  AOI21_X1   g04573(.A1(new_n4569_), .A2(new_n4572_), .B(new_n4829_), .ZN(new_n4830_));
  OAI21_X1   g04574(.A1(new_n4826_), .A2(new_n4825_), .B(new_n4827_), .ZN(new_n4831_));
  NAND3_X1   g04575(.A1(new_n4804_), .A2(new_n4806_), .A3(new_n4823_), .ZN(new_n4832_));
  NAND2_X1   g04576(.A1(new_n4831_), .A2(new_n4832_), .ZN(new_n4833_));
  NOR3_X1    g04577(.A1(new_n4583_), .A2(new_n4564_), .A3(new_n4833_), .ZN(new_n4834_));
  NOR3_X1    g04578(.A1(new_n4830_), .A2(new_n4834_), .A3(new_n4689_), .ZN(new_n4835_));
  OAI21_X1   g04579(.A1(new_n4583_), .A2(new_n4564_), .B(new_n4833_), .ZN(new_n4836_));
  NAND3_X1   g04580(.A1(new_n4569_), .A2(new_n4572_), .A3(new_n4829_), .ZN(new_n4837_));
  AOI21_X1   g04581(.A1(new_n4837_), .A2(new_n4836_), .B(new_n4688_), .ZN(new_n4838_));
  NOR2_X1    g04582(.A1(new_n4838_), .A2(new_n4835_), .ZN(new_n4839_));
  OAI21_X1   g04583(.A1(new_n4684_), .A2(new_n4576_), .B(new_n4839_), .ZN(new_n4840_));
  INV_X1     g04584(.I(new_n4576_), .ZN(new_n4841_));
  INV_X1     g04585(.I(new_n4586_), .ZN(new_n4842_));
  OAI21_X1   g04586(.A1(new_n4592_), .A2(new_n4360_), .B(new_n4842_), .ZN(new_n4843_));
  NAND3_X1   g04587(.A1(new_n4837_), .A2(new_n4836_), .A3(new_n4688_), .ZN(new_n4844_));
  OAI21_X1   g04588(.A1(new_n4830_), .A2(new_n4834_), .B(new_n4689_), .ZN(new_n4845_));
  NAND2_X1   g04589(.A1(new_n4845_), .A2(new_n4844_), .ZN(new_n4846_));
  NAND3_X1   g04590(.A1(new_n4843_), .A2(new_n4841_), .A3(new_n4846_), .ZN(new_n4847_));
  NAND3_X1   g04591(.A1(new_n4847_), .A2(new_n4840_), .A3(new_n4683_), .ZN(new_n4848_));
  INV_X1     g04592(.I(new_n4683_), .ZN(new_n4849_));
  AOI21_X1   g04593(.A1(new_n4843_), .A2(new_n4841_), .B(new_n4846_), .ZN(new_n4850_));
  NOR3_X1    g04594(.A1(new_n4684_), .A2(new_n4839_), .A3(new_n4576_), .ZN(new_n4851_));
  OAI21_X1   g04595(.A1(new_n4850_), .A2(new_n4851_), .B(new_n4849_), .ZN(new_n4852_));
  NAND2_X1   g04596(.A1(new_n4852_), .A2(new_n4848_), .ZN(new_n4853_));
  OAI21_X1   g04597(.A1(new_n4679_), .A2(new_n4600_), .B(new_n4853_), .ZN(new_n4854_));
  AOI21_X1   g04598(.A1(new_n4626_), .A2(new_n4609_), .B(new_n4600_), .ZN(new_n4855_));
  NOR3_X1    g04599(.A1(new_n4850_), .A2(new_n4849_), .A3(new_n4851_), .ZN(new_n4856_));
  AOI21_X1   g04600(.A1(new_n4847_), .A2(new_n4840_), .B(new_n4683_), .ZN(new_n4857_));
  NOR2_X1    g04601(.A1(new_n4856_), .A2(new_n4857_), .ZN(new_n4858_));
  NAND2_X1   g04602(.A1(new_n4855_), .A2(new_n4858_), .ZN(new_n4859_));
  NAND2_X1   g04603(.A1(new_n4859_), .A2(new_n4854_), .ZN(new_n4860_));
  AOI22_X1   g04604(.A1(new_n800_), .A2(\b[31] ), .B1(\b[32] ), .B2(new_n333_), .ZN(new_n4861_));
  OAI21_X1   g04605(.A1(new_n3624_), .A2(new_n392_), .B(new_n4861_), .ZN(new_n4862_));
  AOI21_X1   g04606(.A1(new_n4030_), .A2(new_n330_), .B(new_n4862_), .ZN(new_n4863_));
  XOR2_X1    g04607(.A1(new_n4863_), .A2(new_n312_), .Z(new_n4864_));
  INV_X1     g04608(.I(new_n4864_), .ZN(new_n4865_));
  AOI21_X1   g04609(.A1(new_n4633_), .A2(new_n4634_), .B(new_n4625_), .ZN(new_n4866_));
  NOR2_X1    g04610(.A1(new_n4866_), .A2(new_n4865_), .ZN(new_n4867_));
  INV_X1     g04611(.I(new_n4625_), .ZN(new_n4868_));
  OAI21_X1   g04612(.A1(new_n4399_), .A2(new_n4631_), .B(new_n4868_), .ZN(new_n4869_));
  NOR2_X1    g04613(.A1(new_n4869_), .A2(new_n4864_), .ZN(new_n4870_));
  NOR3_X1    g04614(.A1(new_n4867_), .A2(new_n4870_), .A3(new_n4860_), .ZN(new_n4871_));
  INV_X1     g04615(.I(new_n4871_), .ZN(new_n4872_));
  OAI21_X1   g04616(.A1(new_n4867_), .A2(new_n4870_), .B(new_n4860_), .ZN(new_n4873_));
  AOI21_X1   g04617(.A1(new_n4872_), .A2(new_n4873_), .B(new_n4678_), .ZN(new_n4874_));
  INV_X1     g04618(.I(new_n4678_), .ZN(new_n4875_));
  INV_X1     g04619(.I(new_n4873_), .ZN(new_n4876_));
  NOR3_X1    g04620(.A1(new_n4876_), .A2(new_n4875_), .A3(new_n4871_), .ZN(new_n4877_));
  NOR2_X1    g04621(.A1(new_n4874_), .A2(new_n4877_), .ZN(new_n4878_));
  XOR2_X1    g04622(.A1(new_n4665_), .A2(new_n4878_), .Z(\f[35] ));
  INV_X1     g04623(.I(new_n4877_), .ZN(new_n4880_));
  NAND2_X1   g04624(.A1(new_n4654_), .A2(new_n4652_), .ZN(new_n4881_));
  OAI21_X1   g04625(.A1(new_n4654_), .A2(new_n4652_), .B(new_n4636_), .ZN(new_n4882_));
  OAI21_X1   g04626(.A1(new_n4876_), .A2(new_n4871_), .B(new_n4875_), .ZN(new_n4883_));
  NAND3_X1   g04627(.A1(new_n4882_), .A2(new_n4881_), .A3(new_n4883_), .ZN(new_n4884_));
  NAND2_X1   g04628(.A1(new_n4884_), .A2(new_n4880_), .ZN(new_n4885_));
  INV_X1     g04629(.I(\b[36] ), .ZN(new_n4886_));
  OAI22_X1   g04630(.A1(new_n277_), .A2(new_n4886_), .B1(new_n4666_), .B2(new_n262_), .ZN(new_n4887_));
  AOI21_X1   g04631(.A1(\b[34] ), .A2(new_n283_), .B(new_n4887_), .ZN(new_n4888_));
  XOR2_X1    g04632(.A1(\b[35] ), .A2(\b[36] ), .Z(new_n4889_));
  NAND2_X1   g04633(.A1(new_n4671_), .A2(new_n4639_), .ZN(new_n4890_));
  AOI22_X1   g04634(.A1(new_n4890_), .A2(\b[35] ), .B1(new_n4669_), .B2(\b[34] ), .ZN(new_n4891_));
  NOR2_X1    g04635(.A1(new_n4891_), .A2(new_n4889_), .ZN(new_n4892_));
  INV_X1     g04636(.I(new_n4889_), .ZN(new_n4893_));
  NAND2_X1   g04637(.A1(new_n4890_), .A2(\b[35] ), .ZN(new_n4894_));
  NAND2_X1   g04638(.A1(new_n4669_), .A2(\b[34] ), .ZN(new_n4895_));
  NAND2_X1   g04639(.A1(new_n4894_), .A2(new_n4895_), .ZN(new_n4896_));
  NOR2_X1    g04640(.A1(new_n4896_), .A2(new_n4893_), .ZN(new_n4897_));
  NOR2_X1    g04641(.A1(new_n4897_), .A2(new_n4892_), .ZN(new_n4898_));
  OAI21_X1   g04642(.A1(new_n4898_), .A2(new_n279_), .B(new_n4888_), .ZN(new_n4899_));
  XOR2_X1    g04643(.A1(new_n4899_), .A2(\a[2] ), .Z(new_n4900_));
  INV_X1     g04644(.I(new_n4860_), .ZN(new_n4901_));
  AOI21_X1   g04645(.A1(new_n4869_), .A2(new_n4864_), .B(new_n4901_), .ZN(new_n4902_));
  NOR2_X1    g04646(.A1(new_n4902_), .A2(new_n4870_), .ZN(new_n4903_));
  AOI22_X1   g04647(.A1(new_n800_), .A2(\b[32] ), .B1(\b[33] ), .B2(new_n333_), .ZN(new_n4904_));
  OAI21_X1   g04648(.A1(new_n4022_), .A2(new_n392_), .B(new_n4904_), .ZN(new_n4905_));
  AOI21_X1   g04649(.A1(new_n4223_), .A2(new_n330_), .B(new_n4905_), .ZN(new_n4906_));
  XOR2_X1    g04650(.A1(new_n4906_), .A2(new_n312_), .Z(new_n4907_));
  INV_X1     g04651(.I(new_n4907_), .ZN(new_n4908_));
  NAND2_X1   g04652(.A1(new_n4718_), .A2(new_n4740_), .ZN(new_n4909_));
  NOR2_X1    g04653(.A1(new_n4718_), .A2(new_n4740_), .ZN(new_n4910_));
  OAI21_X1   g04654(.A1(new_n4725_), .A2(new_n4910_), .B(new_n4909_), .ZN(new_n4911_));
  OAI22_X1   g04655(.A1(new_n377_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n438_), .ZN(new_n4912_));
  AOI21_X1   g04656(.A1(\b[4] ), .A2(new_n4053_), .B(new_n4912_), .ZN(new_n4913_));
  OAI21_X1   g04657(.A1(new_n450_), .A2(new_n4727_), .B(new_n4913_), .ZN(new_n4914_));
  XOR2_X1    g04658(.A1(new_n4914_), .A2(\a[32] ), .Z(new_n4915_));
  NAND2_X1   g04659(.A1(new_n4706_), .A2(\b[1] ), .ZN(new_n4916_));
  XOR2_X1    g04660(.A1(\a[34] ), .A2(\a[35] ), .Z(new_n4917_));
  NOR2_X1    g04661(.A1(new_n4247_), .A2(new_n4917_), .ZN(new_n4918_));
  INV_X1     g04662(.I(\a[33] ), .ZN(new_n4919_));
  NAND3_X1   g04663(.A1(new_n3876_), .A2(new_n4919_), .A3(\a[34] ), .ZN(new_n4920_));
  NAND2_X1   g04664(.A1(new_n4920_), .A2(new_n4452_), .ZN(new_n4921_));
  AOI22_X1   g04665(.A1(new_n4918_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n4921_), .ZN(new_n4922_));
  NAND2_X1   g04666(.A1(new_n299_), .A2(new_n4699_), .ZN(new_n4923_));
  NAND3_X1   g04667(.A1(new_n4923_), .A2(new_n4922_), .A3(new_n4916_), .ZN(new_n4924_));
  XOR2_X1    g04668(.A1(new_n4924_), .A2(\a[35] ), .Z(new_n4925_));
  XNOR2_X1   g04669(.A1(\a[35] ), .A2(\a[36] ), .ZN(new_n4926_));
  NOR2_X1    g04670(.A1(new_n4926_), .A2(new_n258_), .ZN(new_n4927_));
  INV_X1     g04671(.I(new_n4927_), .ZN(new_n4928_));
  NOR2_X1    g04672(.A1(new_n4925_), .A2(new_n4928_), .ZN(new_n4929_));
  XOR2_X1    g04673(.A1(new_n4924_), .A2(new_n4446_), .Z(new_n4930_));
  NOR2_X1    g04674(.A1(new_n4930_), .A2(new_n4927_), .ZN(new_n4931_));
  OAI21_X1   g04675(.A1(new_n4929_), .A2(new_n4931_), .B(new_n4716_), .ZN(new_n4932_));
  NAND2_X1   g04676(.A1(new_n4930_), .A2(new_n4927_), .ZN(new_n4933_));
  NAND2_X1   g04677(.A1(new_n4925_), .A2(new_n4928_), .ZN(new_n4934_));
  NAND3_X1   g04678(.A1(new_n4933_), .A2(new_n4934_), .A3(new_n4717_), .ZN(new_n4935_));
  NAND3_X1   g04679(.A1(new_n4932_), .A2(new_n4935_), .A3(new_n4915_), .ZN(new_n4936_));
  XOR2_X1    g04680(.A1(new_n4914_), .A2(new_n3876_), .Z(new_n4937_));
  AOI21_X1   g04681(.A1(new_n4933_), .A2(new_n4934_), .B(new_n4717_), .ZN(new_n4938_));
  NOR3_X1    g04682(.A1(new_n4929_), .A2(new_n4931_), .A3(new_n4716_), .ZN(new_n4939_));
  OAI21_X1   g04683(.A1(new_n4938_), .A2(new_n4939_), .B(new_n4937_), .ZN(new_n4940_));
  NAND2_X1   g04684(.A1(new_n4940_), .A2(new_n4936_), .ZN(new_n4941_));
  XOR2_X1    g04685(.A1(new_n4911_), .A2(new_n4941_), .Z(new_n4942_));
  INV_X1     g04686(.I(new_n4942_), .ZN(new_n4943_));
  AOI22_X1   g04687(.A1(new_n3267_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n3270_), .ZN(new_n4944_));
  OAI21_X1   g04688(.A1(new_n471_), .A2(new_n3475_), .B(new_n4944_), .ZN(new_n4945_));
  AOI21_X1   g04689(.A1(new_n676_), .A2(new_n3273_), .B(new_n4945_), .ZN(new_n4946_));
  XOR2_X1    g04690(.A1(new_n4946_), .A2(new_n3264_), .Z(new_n4947_));
  INV_X1     g04691(.I(new_n4947_), .ZN(new_n4948_));
  NAND2_X1   g04692(.A1(new_n4724_), .A2(new_n4734_), .ZN(new_n4949_));
  NAND2_X1   g04693(.A1(new_n4909_), .A2(new_n4949_), .ZN(new_n4950_));
  NOR2_X1    g04694(.A1(new_n4950_), .A2(new_n4725_), .ZN(new_n4951_));
  NOR2_X1    g04695(.A1(new_n4724_), .A2(new_n4734_), .ZN(new_n4952_));
  NOR2_X1    g04696(.A1(new_n4910_), .A2(new_n4952_), .ZN(new_n4953_));
  NOR2_X1    g04697(.A1(new_n4953_), .A2(new_n4719_), .ZN(new_n4954_));
  NOR3_X1    g04698(.A1(new_n4954_), .A2(new_n4951_), .A3(new_n4738_), .ZN(new_n4955_));
  AOI21_X1   g04699(.A1(new_n4757_), .A2(new_n4753_), .B(new_n4955_), .ZN(new_n4956_));
  NOR2_X1    g04700(.A1(new_n4956_), .A2(new_n4948_), .ZN(new_n4957_));
  NAND2_X1   g04701(.A1(new_n4953_), .A2(new_n4719_), .ZN(new_n4958_));
  NAND2_X1   g04702(.A1(new_n4950_), .A2(new_n4725_), .ZN(new_n4959_));
  NAND3_X1   g04703(.A1(new_n4958_), .A2(new_n4959_), .A3(new_n4747_), .ZN(new_n4960_));
  OAI21_X1   g04704(.A1(new_n4751_), .A2(new_n4759_), .B(new_n4960_), .ZN(new_n4961_));
  NOR2_X1    g04705(.A1(new_n4961_), .A2(new_n4947_), .ZN(new_n4962_));
  NOR3_X1    g04706(.A1(new_n4957_), .A2(new_n4962_), .A3(new_n4943_), .ZN(new_n4963_));
  NAND2_X1   g04707(.A1(new_n4961_), .A2(new_n4947_), .ZN(new_n4964_));
  NAND2_X1   g04708(.A1(new_n4956_), .A2(new_n4948_), .ZN(new_n4965_));
  AOI21_X1   g04709(.A1(new_n4965_), .A2(new_n4964_), .B(new_n4942_), .ZN(new_n4966_));
  NOR2_X1    g04710(.A1(new_n4966_), .A2(new_n4963_), .ZN(new_n4967_));
  INV_X1     g04711(.I(new_n4967_), .ZN(new_n4968_));
  INV_X1     g04712(.I(new_n4769_), .ZN(new_n4969_));
  AOI22_X1   g04713(.A1(new_n2716_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n2719_), .ZN(new_n4970_));
  OAI21_X1   g04714(.A1(new_n776_), .A2(new_n2924_), .B(new_n4970_), .ZN(new_n4971_));
  AOI21_X1   g04715(.A1(new_n1194_), .A2(new_n2722_), .B(new_n4971_), .ZN(new_n4972_));
  XOR2_X1    g04716(.A1(new_n4972_), .A2(new_n2714_), .Z(new_n4973_));
  INV_X1     g04717(.I(new_n4973_), .ZN(new_n4974_));
  AOI21_X1   g04718(.A1(new_n4772_), .A2(new_n4969_), .B(new_n4974_), .ZN(new_n4975_));
  NOR3_X1    g04719(.A1(new_n4780_), .A2(new_n4769_), .A3(new_n4973_), .ZN(new_n4976_));
  NOR3_X1    g04720(.A1(new_n4976_), .A2(new_n4975_), .A3(new_n4968_), .ZN(new_n4977_));
  OAI21_X1   g04721(.A1(new_n4780_), .A2(new_n4769_), .B(new_n4973_), .ZN(new_n4978_));
  NAND3_X1   g04722(.A1(new_n4772_), .A2(new_n4969_), .A3(new_n4974_), .ZN(new_n4979_));
  AOI21_X1   g04723(.A1(new_n4978_), .A2(new_n4979_), .B(new_n4967_), .ZN(new_n4980_));
  NOR2_X1    g04724(.A1(new_n4977_), .A2(new_n4980_), .ZN(new_n4981_));
  INV_X1     g04725(.I(new_n4981_), .ZN(new_n4982_));
  OAI22_X1   g04726(.A1(new_n2189_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n2194_), .ZN(new_n4983_));
  AOI21_X1   g04727(.A1(\b[13] ), .A2(new_n2361_), .B(new_n4983_), .ZN(new_n4984_));
  OAI21_X1   g04728(.A1(new_n1275_), .A2(new_n2197_), .B(new_n4984_), .ZN(new_n4985_));
  XOR2_X1    g04729(.A1(new_n4985_), .A2(\a[23] ), .Z(new_n4986_));
  INV_X1     g04730(.I(new_n4986_), .ZN(new_n4987_));
  AOI21_X1   g04731(.A1(new_n4792_), .A2(new_n4779_), .B(new_n4987_), .ZN(new_n4988_));
  NOR3_X1    g04732(.A1(new_n4785_), .A2(new_n4787_), .A3(new_n4986_), .ZN(new_n4989_));
  NOR3_X1    g04733(.A1(new_n4989_), .A2(new_n4988_), .A3(new_n4982_), .ZN(new_n4990_));
  OAI21_X1   g04734(.A1(new_n4785_), .A2(new_n4787_), .B(new_n4986_), .ZN(new_n4991_));
  NAND3_X1   g04735(.A1(new_n4792_), .A2(new_n4779_), .A3(new_n4987_), .ZN(new_n4992_));
  AOI21_X1   g04736(.A1(new_n4991_), .A2(new_n4992_), .B(new_n4981_), .ZN(new_n4993_));
  NOR2_X1    g04737(.A1(new_n4990_), .A2(new_n4993_), .ZN(new_n4994_));
  INV_X1     g04738(.I(new_n4994_), .ZN(new_n4995_));
  AOI22_X1   g04739(.A1(new_n1738_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n1743_), .ZN(new_n4996_));
  OAI21_X1   g04740(.A1(new_n1296_), .A2(new_n1931_), .B(new_n4996_), .ZN(new_n4997_));
  AOI21_X1   g04741(.A1(new_n2038_), .A2(new_n1746_), .B(new_n4997_), .ZN(new_n4998_));
  XOR2_X1    g04742(.A1(new_n4998_), .A2(new_n1736_), .Z(new_n4999_));
  INV_X1     g04743(.I(new_n4999_), .ZN(new_n5000_));
  OAI21_X1   g04744(.A1(new_n4797_), .A2(new_n4544_), .B(new_n4795_), .ZN(new_n5001_));
  AOI21_X1   g04745(.A1(new_n5001_), .A2(new_n4798_), .B(new_n5000_), .ZN(new_n5002_));
  AOI21_X1   g04746(.A1(new_n4691_), .A2(new_n4535_), .B(new_n4800_), .ZN(new_n5003_));
  NOR3_X1    g04747(.A1(new_n5003_), .A2(new_n4791_), .A3(new_n4999_), .ZN(new_n5004_));
  NOR3_X1    g04748(.A1(new_n5002_), .A2(new_n5004_), .A3(new_n4995_), .ZN(new_n5005_));
  OAI21_X1   g04749(.A1(new_n5003_), .A2(new_n4791_), .B(new_n4999_), .ZN(new_n5006_));
  NAND3_X1   g04750(.A1(new_n5001_), .A2(new_n4798_), .A3(new_n5000_), .ZN(new_n5007_));
  AOI21_X1   g04751(.A1(new_n5006_), .A2(new_n5007_), .B(new_n4994_), .ZN(new_n5008_));
  NOR2_X1    g04752(.A1(new_n5008_), .A2(new_n5005_), .ZN(new_n5009_));
  INV_X1     g04753(.I(new_n5009_), .ZN(new_n5010_));
  OAI22_X1   g04754(.A1(new_n1592_), .A2(new_n2027_), .B1(new_n1860_), .B2(new_n1505_), .ZN(new_n5011_));
  AOI21_X1   g04755(.A1(\b[19] ), .A2(new_n1584_), .B(new_n5011_), .ZN(new_n5012_));
  OAI21_X1   g04756(.A1(new_n3727_), .A2(new_n1732_), .B(new_n5012_), .ZN(new_n5013_));
  XOR2_X1    g04757(.A1(new_n5013_), .A2(\a[17] ), .Z(new_n5014_));
  NOR2_X1    g04758(.A1(new_n4802_), .A2(new_n4818_), .ZN(new_n5015_));
  OAI21_X1   g04759(.A1(new_n4797_), .A2(new_n4544_), .B(new_n4800_), .ZN(new_n5016_));
  NAND3_X1   g04760(.A1(new_n4691_), .A2(new_n4795_), .A3(new_n4535_), .ZN(new_n5017_));
  AOI21_X1   g04761(.A1(new_n5016_), .A2(new_n5017_), .B(new_n4817_), .ZN(new_n5018_));
  NOR3_X1    g04762(.A1(new_n4801_), .A2(new_n4796_), .A3(new_n4818_), .ZN(new_n5019_));
  NOR2_X1    g04763(.A1(new_n5019_), .A2(new_n5018_), .ZN(new_n5020_));
  AOI21_X1   g04764(.A1(new_n4565_), .A2(new_n4805_), .B(new_n5020_), .ZN(new_n5021_));
  OAI21_X1   g04765(.A1(new_n5021_), .A2(new_n5015_), .B(new_n5014_), .ZN(new_n5022_));
  INV_X1     g04766(.I(new_n5014_), .ZN(new_n5023_));
  INV_X1     g04767(.I(new_n5015_), .ZN(new_n5024_));
  OAI21_X1   g04768(.A1(new_n4801_), .A2(new_n4796_), .B(new_n4818_), .ZN(new_n5025_));
  NAND3_X1   g04769(.A1(new_n5016_), .A2(new_n5017_), .A3(new_n4817_), .ZN(new_n5026_));
  NAND2_X1   g04770(.A1(new_n5025_), .A2(new_n5026_), .ZN(new_n5027_));
  OAI21_X1   g04771(.A1(new_n4554_), .A2(new_n4690_), .B(new_n5027_), .ZN(new_n5028_));
  NAND3_X1   g04772(.A1(new_n5028_), .A2(new_n5023_), .A3(new_n5024_), .ZN(new_n5029_));
  NAND2_X1   g04773(.A1(new_n5022_), .A2(new_n5029_), .ZN(new_n5030_));
  NOR2_X1    g04774(.A1(new_n5030_), .A2(new_n5010_), .ZN(new_n5031_));
  AOI21_X1   g04775(.A1(new_n5028_), .A2(new_n5024_), .B(new_n5023_), .ZN(new_n5032_));
  NOR3_X1    g04776(.A1(new_n5021_), .A2(new_n5014_), .A3(new_n5015_), .ZN(new_n5033_));
  NOR2_X1    g04777(.A1(new_n5033_), .A2(new_n5032_), .ZN(new_n5034_));
  NOR2_X1    g04778(.A1(new_n5034_), .A2(new_n5009_), .ZN(new_n5035_));
  NOR2_X1    g04779(.A1(new_n5035_), .A2(new_n5031_), .ZN(new_n5036_));
  OAI22_X1   g04780(.A1(new_n993_), .A2(new_n2495_), .B1(new_n2463_), .B2(new_n997_), .ZN(new_n5037_));
  AOI21_X1   g04781(.A1(\b[22] ), .A2(new_n1486_), .B(new_n5037_), .ZN(new_n5038_));
  OAI21_X1   g04782(.A1(new_n2506_), .A2(new_n1323_), .B(new_n5038_), .ZN(new_n5039_));
  XOR2_X1    g04783(.A1(new_n5039_), .A2(\a[14] ), .Z(new_n5040_));
  NOR2_X1    g04784(.A1(new_n4820_), .A2(new_n4821_), .ZN(new_n5041_));
  NAND3_X1   g04785(.A1(new_n4565_), .A2(new_n4805_), .A3(new_n5020_), .ZN(new_n5042_));
  NAND3_X1   g04786(.A1(new_n5028_), .A2(new_n5042_), .A3(new_n5041_), .ZN(new_n5043_));
  INV_X1     g04787(.I(new_n5043_), .ZN(new_n5044_));
  OAI21_X1   g04788(.A1(new_n4830_), .A2(new_n5044_), .B(new_n5040_), .ZN(new_n5045_));
  INV_X1     g04789(.I(new_n5040_), .ZN(new_n5046_));
  NAND3_X1   g04790(.A1(new_n4836_), .A2(new_n5046_), .A3(new_n5043_), .ZN(new_n5047_));
  NAND3_X1   g04791(.A1(new_n5045_), .A2(new_n5047_), .A3(new_n5036_), .ZN(new_n5048_));
  NAND2_X1   g04792(.A1(new_n5034_), .A2(new_n5009_), .ZN(new_n5049_));
  NAND2_X1   g04793(.A1(new_n5030_), .A2(new_n5010_), .ZN(new_n5050_));
  NAND2_X1   g04794(.A1(new_n5049_), .A2(new_n5050_), .ZN(new_n5051_));
  NAND2_X1   g04795(.A1(new_n5045_), .A2(new_n5047_), .ZN(new_n5052_));
  NAND2_X1   g04796(.A1(new_n5052_), .A2(new_n5051_), .ZN(new_n5053_));
  NAND2_X1   g04797(.A1(new_n5053_), .A2(new_n5048_), .ZN(new_n5054_));
  OAI22_X1   g04798(.A1(new_n713_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n717_), .ZN(new_n5055_));
  AOI21_X1   g04799(.A1(\b[25] ), .A2(new_n1126_), .B(new_n5055_), .ZN(new_n5056_));
  OAI21_X1   g04800(.A1(new_n3165_), .A2(new_n986_), .B(new_n5056_), .ZN(new_n5057_));
  XOR2_X1    g04801(.A1(new_n5057_), .A2(\a[11] ), .Z(new_n5058_));
  INV_X1     g04802(.I(new_n5058_), .ZN(new_n5059_));
  NAND3_X1   g04803(.A1(new_n4843_), .A2(new_n4841_), .A3(new_n4839_), .ZN(new_n5060_));
  AOI21_X1   g04804(.A1(new_n5060_), .A2(new_n4844_), .B(new_n5059_), .ZN(new_n5061_));
  NOR3_X1    g04805(.A1(new_n4684_), .A2(new_n4576_), .A3(new_n4846_), .ZN(new_n5062_));
  NOR3_X1    g04806(.A1(new_n5062_), .A2(new_n4835_), .A3(new_n5058_), .ZN(new_n5063_));
  NOR3_X1    g04807(.A1(new_n5061_), .A2(new_n5063_), .A3(new_n5054_), .ZN(new_n5064_));
  XOR2_X1    g04808(.A1(new_n5052_), .A2(new_n5051_), .Z(new_n5065_));
  OAI21_X1   g04809(.A1(new_n5062_), .A2(new_n4835_), .B(new_n5058_), .ZN(new_n5066_));
  NAND3_X1   g04810(.A1(new_n5060_), .A2(new_n4844_), .A3(new_n5059_), .ZN(new_n5067_));
  AOI21_X1   g04811(.A1(new_n5067_), .A2(new_n5066_), .B(new_n5065_), .ZN(new_n5068_));
  NOR2_X1    g04812(.A1(new_n5068_), .A2(new_n5064_), .ZN(new_n5069_));
  INV_X1     g04813(.I(new_n5069_), .ZN(new_n5070_));
  AOI21_X1   g04814(.A1(new_n4847_), .A2(new_n4840_), .B(new_n4849_), .ZN(new_n5071_));
  INV_X1     g04815(.I(new_n5071_), .ZN(new_n5072_));
  AOI22_X1   g04816(.A1(new_n518_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n636_), .ZN(new_n5073_));
  OAI21_X1   g04817(.A1(new_n3185_), .A2(new_n917_), .B(new_n5073_), .ZN(new_n5074_));
  AOI21_X1   g04818(.A1(new_n4230_), .A2(new_n618_), .B(new_n5074_), .ZN(new_n5075_));
  XOR2_X1    g04819(.A1(new_n5075_), .A2(new_n488_), .Z(new_n5076_));
  INV_X1     g04820(.I(new_n5076_), .ZN(new_n5077_));
  AOI21_X1   g04821(.A1(new_n4854_), .A2(new_n5072_), .B(new_n5077_), .ZN(new_n5078_));
  NAND3_X1   g04822(.A1(new_n4611_), .A2(new_n4377_), .A3(new_n4609_), .ZN(new_n5079_));
  AOI21_X1   g04823(.A1(new_n5079_), .A2(new_n4599_), .B(new_n4858_), .ZN(new_n5080_));
  NOR3_X1    g04824(.A1(new_n5080_), .A2(new_n5071_), .A3(new_n5076_), .ZN(new_n5081_));
  NOR3_X1    g04825(.A1(new_n5078_), .A2(new_n5081_), .A3(new_n5070_), .ZN(new_n5082_));
  OAI21_X1   g04826(.A1(new_n5080_), .A2(new_n5071_), .B(new_n5076_), .ZN(new_n5083_));
  NAND3_X1   g04827(.A1(new_n4854_), .A2(new_n5072_), .A3(new_n5077_), .ZN(new_n5084_));
  AOI21_X1   g04828(.A1(new_n5084_), .A2(new_n5083_), .B(new_n5069_), .ZN(new_n5085_));
  OAI21_X1   g04829(.A1(new_n5085_), .A2(new_n5082_), .B(new_n4908_), .ZN(new_n5086_));
  NOR3_X1    g04830(.A1(new_n5085_), .A2(new_n5082_), .A3(new_n4908_), .ZN(new_n5087_));
  INV_X1     g04831(.I(new_n5087_), .ZN(new_n5088_));
  NAND2_X1   g04832(.A1(new_n5088_), .A2(new_n5086_), .ZN(new_n5089_));
  XOR2_X1    g04833(.A1(new_n4903_), .A2(new_n5089_), .Z(new_n5090_));
  NAND2_X1   g04834(.A1(new_n5090_), .A2(new_n4900_), .ZN(new_n5091_));
  INV_X1     g04835(.I(new_n4903_), .ZN(new_n5092_));
  NAND3_X1   g04836(.A1(new_n5092_), .A2(new_n5086_), .A3(new_n5088_), .ZN(new_n5093_));
  NAND2_X1   g04837(.A1(new_n5089_), .A2(new_n4903_), .ZN(new_n5094_));
  AOI21_X1   g04838(.A1(new_n5093_), .A2(new_n5094_), .B(new_n4900_), .ZN(new_n5095_));
  INV_X1     g04839(.I(new_n5095_), .ZN(new_n5096_));
  NAND2_X1   g04840(.A1(new_n5091_), .A2(new_n5096_), .ZN(new_n5097_));
  XOR2_X1    g04841(.A1(new_n4885_), .A2(new_n5097_), .Z(\f[36] ));
  NAND2_X1   g04842(.A1(new_n4866_), .A2(new_n4865_), .ZN(new_n5099_));
  OAI21_X1   g04843(.A1(new_n4866_), .A2(new_n4865_), .B(new_n4860_), .ZN(new_n5100_));
  NAND3_X1   g04844(.A1(new_n5100_), .A2(new_n5099_), .A3(new_n5086_), .ZN(new_n5101_));
  NAND2_X1   g04845(.A1(new_n5101_), .A2(new_n5088_), .ZN(new_n5102_));
  INV_X1     g04846(.I(new_n4649_), .ZN(new_n5103_));
  AOI22_X1   g04847(.A1(new_n800_), .A2(\b[33] ), .B1(\b[34] ), .B2(new_n333_), .ZN(new_n5104_));
  OAI21_X1   g04848(.A1(new_n4023_), .A2(new_n392_), .B(new_n5104_), .ZN(new_n5105_));
  AOI21_X1   g04849(.A1(new_n5103_), .A2(new_n330_), .B(new_n5105_), .ZN(new_n5106_));
  XOR2_X1    g04850(.A1(new_n5106_), .A2(\a[5] ), .Z(new_n5107_));
  AOI21_X1   g04851(.A1(new_n5070_), .A2(new_n5083_), .B(new_n5081_), .ZN(new_n5108_));
  AOI21_X1   g04852(.A1(new_n5054_), .A2(new_n5066_), .B(new_n5063_), .ZN(new_n5109_));
  NOR3_X1    g04853(.A1(new_n4830_), .A2(new_n5040_), .A3(new_n5044_), .ZN(new_n5110_));
  AOI21_X1   g04854(.A1(new_n5051_), .A2(new_n5045_), .B(new_n5110_), .ZN(new_n5111_));
  OAI22_X1   g04855(.A1(new_n993_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n997_), .ZN(new_n5112_));
  AOI21_X1   g04856(.A1(\b[23] ), .A2(new_n1486_), .B(new_n5112_), .ZN(new_n5113_));
  OAI21_X1   g04857(.A1(new_n2655_), .A2(new_n1323_), .B(new_n5113_), .ZN(new_n5114_));
  XOR2_X1    g04858(.A1(new_n5114_), .A2(\a[14] ), .Z(new_n5115_));
  INV_X1     g04859(.I(new_n5115_), .ZN(new_n5116_));
  NOR2_X1    g04860(.A1(new_n5032_), .A2(new_n5009_), .ZN(new_n5117_));
  OAI22_X1   g04861(.A1(new_n1592_), .A2(new_n2142_), .B1(new_n2027_), .B2(new_n1505_), .ZN(new_n5118_));
  AOI21_X1   g04862(.A1(\b[20] ), .A2(new_n1584_), .B(new_n5118_), .ZN(new_n5119_));
  OAI21_X1   g04863(.A1(new_n2153_), .A2(new_n1732_), .B(new_n5119_), .ZN(new_n5120_));
  XOR2_X1    g04864(.A1(new_n5120_), .A2(\a[17] ), .Z(new_n5121_));
  INV_X1     g04865(.I(new_n5121_), .ZN(new_n5122_));
  NAND2_X1   g04866(.A1(new_n5006_), .A2(new_n4995_), .ZN(new_n5123_));
  AOI22_X1   g04867(.A1(new_n1738_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n1743_), .ZN(new_n5124_));
  NAND2_X1   g04868(.A1(new_n1939_), .A2(\b[17] ), .ZN(new_n5125_));
  NAND2_X1   g04869(.A1(new_n1695_), .A2(new_n1746_), .ZN(new_n5126_));
  NAND3_X1   g04870(.A1(new_n5126_), .A2(new_n5124_), .A3(new_n5125_), .ZN(new_n5127_));
  XOR2_X1    g04871(.A1(new_n5127_), .A2(\a[20] ), .Z(new_n5128_));
  INV_X1     g04872(.I(new_n5128_), .ZN(new_n5129_));
  OAI21_X1   g04873(.A1(new_n4981_), .A2(new_n4988_), .B(new_n4992_), .ZN(new_n5130_));
  AOI22_X1   g04874(.A1(new_n2202_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n2205_), .ZN(new_n5131_));
  OAI21_X1   g04875(.A1(new_n1093_), .A2(new_n2370_), .B(new_n5131_), .ZN(new_n5132_));
  AOI21_X1   g04876(.A1(new_n1701_), .A2(new_n2208_), .B(new_n5132_), .ZN(new_n5133_));
  XOR2_X1    g04877(.A1(new_n5133_), .A2(new_n2200_), .Z(new_n5134_));
  INV_X1     g04878(.I(new_n5134_), .ZN(new_n5135_));
  NAND2_X1   g04879(.A1(new_n4978_), .A2(new_n4968_), .ZN(new_n5136_));
  OAI21_X1   g04880(.A1(new_n4956_), .A2(new_n4948_), .B(new_n4943_), .ZN(new_n5137_));
  AOI21_X1   g04881(.A1(new_n4719_), .A2(new_n4949_), .B(new_n4952_), .ZN(new_n5138_));
  NOR3_X1    g04882(.A1(new_n4938_), .A2(new_n4939_), .A3(new_n4937_), .ZN(new_n5139_));
  AOI21_X1   g04883(.A1(new_n4932_), .A2(new_n4935_), .B(new_n4915_), .ZN(new_n5140_));
  NOR2_X1    g04884(.A1(new_n5139_), .A2(new_n5140_), .ZN(new_n5141_));
  AOI21_X1   g04885(.A1(new_n4932_), .A2(new_n4935_), .B(new_n4937_), .ZN(new_n5142_));
  INV_X1     g04886(.I(new_n5142_), .ZN(new_n5143_));
  OAI21_X1   g04887(.A1(new_n5138_), .A2(new_n5141_), .B(new_n5143_), .ZN(new_n5144_));
  NAND2_X1   g04888(.A1(new_n4716_), .A2(new_n4928_), .ZN(new_n5145_));
  NOR2_X1    g04889(.A1(new_n4716_), .A2(new_n4928_), .ZN(new_n5146_));
  AOI21_X1   g04890(.A1(new_n4925_), .A2(new_n5145_), .B(new_n5146_), .ZN(new_n5147_));
  AOI22_X1   g04891(.A1(new_n4918_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n4921_), .ZN(new_n5148_));
  NAND2_X1   g04892(.A1(new_n4706_), .A2(\b[2] ), .ZN(new_n5149_));
  NAND2_X1   g04893(.A1(new_n1725_), .A2(new_n4699_), .ZN(new_n5150_));
  NAND3_X1   g04894(.A1(new_n5150_), .A2(new_n5148_), .A3(new_n5149_), .ZN(new_n5151_));
  XOR2_X1    g04895(.A1(new_n5151_), .A2(new_n4446_), .Z(new_n5152_));
  INV_X1     g04896(.I(new_n5152_), .ZN(new_n5153_));
  XOR2_X1    g04897(.A1(\a[37] ), .A2(\a[38] ), .Z(new_n5154_));
  NOR2_X1    g04898(.A1(new_n4926_), .A2(new_n5154_), .ZN(new_n5155_));
  INV_X1     g04899(.I(\a[36] ), .ZN(new_n5156_));
  NAND3_X1   g04900(.A1(new_n4446_), .A2(new_n5156_), .A3(\a[37] ), .ZN(new_n5157_));
  INV_X1     g04901(.I(\a[37] ), .ZN(new_n5158_));
  NAND3_X1   g04902(.A1(new_n5158_), .A2(\a[35] ), .A3(\a[36] ), .ZN(new_n5159_));
  NAND2_X1   g04903(.A1(new_n5157_), .A2(new_n5159_), .ZN(new_n5160_));
  AOI22_X1   g04904(.A1(new_n5155_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n5160_), .ZN(new_n5161_));
  INV_X1     g04905(.I(\a[38] ), .ZN(new_n5162_));
  NOR2_X1    g04906(.A1(new_n5162_), .A2(\a[37] ), .ZN(new_n5163_));
  NOR2_X1    g04907(.A1(new_n5158_), .A2(\a[38] ), .ZN(new_n5164_));
  NOR2_X1    g04908(.A1(new_n5163_), .A2(new_n5164_), .ZN(new_n5165_));
  NOR2_X1    g04909(.A1(new_n5165_), .A2(new_n4926_), .ZN(new_n5166_));
  NAND2_X1   g04910(.A1(new_n5166_), .A2(new_n263_), .ZN(new_n5167_));
  NAND2_X1   g04911(.A1(new_n5161_), .A2(new_n5167_), .ZN(new_n5168_));
  NAND2_X1   g04912(.A1(new_n5168_), .A2(\a[38] ), .ZN(new_n5169_));
  INV_X1     g04913(.I(new_n5168_), .ZN(new_n5170_));
  NAND2_X1   g04914(.A1(new_n5170_), .A2(new_n5162_), .ZN(new_n5171_));
  NOR2_X1    g04915(.A1(new_n4927_), .A2(new_n5162_), .ZN(new_n5172_));
  INV_X1     g04916(.I(new_n5172_), .ZN(new_n5173_));
  NAND3_X1   g04917(.A1(new_n5171_), .A2(new_n5169_), .A3(new_n5173_), .ZN(new_n5174_));
  NAND3_X1   g04918(.A1(new_n5168_), .A2(\a[38] ), .A3(new_n4928_), .ZN(new_n5175_));
  NAND2_X1   g04919(.A1(new_n5174_), .A2(new_n5175_), .ZN(new_n5176_));
  NAND2_X1   g04920(.A1(new_n5176_), .A2(new_n5153_), .ZN(new_n5177_));
  NAND3_X1   g04921(.A1(new_n5152_), .A2(new_n5174_), .A3(new_n5175_), .ZN(new_n5178_));
  AOI21_X1   g04922(.A1(new_n5177_), .A2(new_n5178_), .B(new_n5147_), .ZN(new_n5179_));
  NAND2_X1   g04923(.A1(new_n5145_), .A2(new_n4925_), .ZN(new_n5180_));
  INV_X1     g04924(.I(new_n5146_), .ZN(new_n5181_));
  NAND2_X1   g04925(.A1(new_n5180_), .A2(new_n5181_), .ZN(new_n5182_));
  AOI21_X1   g04926(.A1(new_n5174_), .A2(new_n5175_), .B(new_n5152_), .ZN(new_n5183_));
  INV_X1     g04927(.I(new_n5178_), .ZN(new_n5184_));
  NOR3_X1    g04928(.A1(new_n5182_), .A2(new_n5184_), .A3(new_n5183_), .ZN(new_n5185_));
  NOR2_X1    g04929(.A1(new_n5185_), .A2(new_n5179_), .ZN(new_n5186_));
  OAI22_X1   g04930(.A1(new_n438_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n471_), .ZN(new_n5187_));
  AOI21_X1   g04931(.A1(\b[5] ), .A2(new_n4053_), .B(new_n5187_), .ZN(new_n5188_));
  OAI21_X1   g04932(.A1(new_n485_), .A2(new_n4727_), .B(new_n5188_), .ZN(new_n5189_));
  XOR2_X1    g04933(.A1(new_n5189_), .A2(\a[32] ), .Z(new_n5190_));
  INV_X1     g04934(.I(new_n5190_), .ZN(new_n5191_));
  NAND2_X1   g04935(.A1(new_n5186_), .A2(new_n5191_), .ZN(new_n5192_));
  OAI21_X1   g04936(.A1(new_n5183_), .A2(new_n5184_), .B(new_n5182_), .ZN(new_n5193_));
  NAND3_X1   g04937(.A1(new_n5177_), .A2(new_n5147_), .A3(new_n5178_), .ZN(new_n5194_));
  NAND2_X1   g04938(.A1(new_n5193_), .A2(new_n5194_), .ZN(new_n5195_));
  NAND2_X1   g04939(.A1(new_n5195_), .A2(new_n5190_), .ZN(new_n5196_));
  NAND2_X1   g04940(.A1(new_n5196_), .A2(new_n5192_), .ZN(new_n5197_));
  NAND2_X1   g04941(.A1(new_n5197_), .A2(new_n5144_), .ZN(new_n5198_));
  AOI21_X1   g04942(.A1(new_n4911_), .A2(new_n4941_), .B(new_n5142_), .ZN(new_n5199_));
  NAND3_X1   g04943(.A1(new_n5199_), .A2(new_n5196_), .A3(new_n5192_), .ZN(new_n5200_));
  AOI22_X1   g04944(.A1(new_n3267_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n3270_), .ZN(new_n5201_));
  OAI21_X1   g04945(.A1(new_n577_), .A2(new_n3475_), .B(new_n5201_), .ZN(new_n5202_));
  AOI21_X1   g04946(.A1(new_n1059_), .A2(new_n3273_), .B(new_n5202_), .ZN(new_n5203_));
  XOR2_X1    g04947(.A1(new_n5203_), .A2(new_n3264_), .Z(new_n5204_));
  INV_X1     g04948(.I(new_n5204_), .ZN(new_n5205_));
  NAND3_X1   g04949(.A1(new_n5198_), .A2(new_n5200_), .A3(new_n5205_), .ZN(new_n5206_));
  AOI21_X1   g04950(.A1(new_n5192_), .A2(new_n5196_), .B(new_n5199_), .ZN(new_n5207_));
  INV_X1     g04951(.I(new_n5200_), .ZN(new_n5208_));
  OAI21_X1   g04952(.A1(new_n5208_), .A2(new_n5207_), .B(new_n5204_), .ZN(new_n5209_));
  NAND2_X1   g04953(.A1(new_n5209_), .A2(new_n5206_), .ZN(new_n5210_));
  NAND3_X1   g04954(.A1(new_n5210_), .A2(new_n5137_), .A3(new_n4965_), .ZN(new_n5211_));
  INV_X1     g04955(.I(new_n5211_), .ZN(new_n5212_));
  AOI21_X1   g04956(.A1(new_n4965_), .A2(new_n5137_), .B(new_n5210_), .ZN(new_n5213_));
  OAI22_X1   g04957(.A1(new_n2703_), .A2(new_n1070_), .B1(new_n941_), .B2(new_n2708_), .ZN(new_n5214_));
  AOI21_X1   g04958(.A1(\b[11] ), .A2(new_n2906_), .B(new_n5214_), .ZN(new_n5215_));
  OAI21_X1   g04959(.A1(new_n1082_), .A2(new_n2711_), .B(new_n5215_), .ZN(new_n5216_));
  XOR2_X1    g04960(.A1(new_n5216_), .A2(\a[26] ), .Z(new_n5217_));
  OAI21_X1   g04961(.A1(new_n5212_), .A2(new_n5213_), .B(new_n5217_), .ZN(new_n5218_));
  NAND2_X1   g04962(.A1(new_n5137_), .A2(new_n4965_), .ZN(new_n5219_));
  NAND3_X1   g04963(.A1(new_n5219_), .A2(new_n5206_), .A3(new_n5209_), .ZN(new_n5220_));
  XOR2_X1    g04964(.A1(new_n5216_), .A2(new_n2714_), .Z(new_n5221_));
  NAND3_X1   g04965(.A1(new_n5220_), .A2(new_n5221_), .A3(new_n5211_), .ZN(new_n5222_));
  NAND2_X1   g04966(.A1(new_n5218_), .A2(new_n5222_), .ZN(new_n5223_));
  AOI21_X1   g04967(.A1(new_n5136_), .A2(new_n4979_), .B(new_n5223_), .ZN(new_n5224_));
  OAI21_X1   g04968(.A1(new_n4967_), .A2(new_n4975_), .B(new_n4979_), .ZN(new_n5225_));
  AOI21_X1   g04969(.A1(new_n5220_), .A2(new_n5211_), .B(new_n5221_), .ZN(new_n5226_));
  NOR3_X1    g04970(.A1(new_n5212_), .A2(new_n5213_), .A3(new_n5217_), .ZN(new_n5227_));
  NOR2_X1    g04971(.A1(new_n5227_), .A2(new_n5226_), .ZN(new_n5228_));
  NOR2_X1    g04972(.A1(new_n5225_), .A2(new_n5228_), .ZN(new_n5229_));
  NOR3_X1    g04973(.A1(new_n5224_), .A2(new_n5229_), .A3(new_n5135_), .ZN(new_n5230_));
  NAND2_X1   g04974(.A1(new_n5225_), .A2(new_n5228_), .ZN(new_n5231_));
  NAND3_X1   g04975(.A1(new_n5136_), .A2(new_n5223_), .A3(new_n4979_), .ZN(new_n5232_));
  AOI21_X1   g04976(.A1(new_n5231_), .A2(new_n5232_), .B(new_n5134_), .ZN(new_n5233_));
  NOR2_X1    g04977(.A1(new_n5230_), .A2(new_n5233_), .ZN(new_n5234_));
  NOR2_X1    g04978(.A1(new_n5130_), .A2(new_n5234_), .ZN(new_n5235_));
  AOI21_X1   g04979(.A1(new_n4982_), .A2(new_n4991_), .B(new_n4989_), .ZN(new_n5236_));
  NAND3_X1   g04980(.A1(new_n5231_), .A2(new_n5232_), .A3(new_n5134_), .ZN(new_n5237_));
  OAI21_X1   g04981(.A1(new_n5224_), .A2(new_n5229_), .B(new_n5135_), .ZN(new_n5238_));
  NAND2_X1   g04982(.A1(new_n5238_), .A2(new_n5237_), .ZN(new_n5239_));
  NOR2_X1    g04983(.A1(new_n5236_), .A2(new_n5239_), .ZN(new_n5240_));
  NOR3_X1    g04984(.A1(new_n5240_), .A2(new_n5235_), .A3(new_n5129_), .ZN(new_n5241_));
  NAND2_X1   g04985(.A1(new_n4991_), .A2(new_n4982_), .ZN(new_n5242_));
  NAND3_X1   g04986(.A1(new_n5242_), .A2(new_n5239_), .A3(new_n4992_), .ZN(new_n5243_));
  NAND2_X1   g04987(.A1(new_n5130_), .A2(new_n5234_), .ZN(new_n5244_));
  AOI21_X1   g04988(.A1(new_n5244_), .A2(new_n5243_), .B(new_n5128_), .ZN(new_n5245_));
  NOR2_X1    g04989(.A1(new_n5241_), .A2(new_n5245_), .ZN(new_n5246_));
  NAND3_X1   g04990(.A1(new_n5123_), .A2(new_n5246_), .A3(new_n5007_), .ZN(new_n5247_));
  OAI21_X1   g04991(.A1(new_n4994_), .A2(new_n5002_), .B(new_n5007_), .ZN(new_n5248_));
  NAND3_X1   g04992(.A1(new_n5244_), .A2(new_n5243_), .A3(new_n5128_), .ZN(new_n5249_));
  OAI21_X1   g04993(.A1(new_n5240_), .A2(new_n5235_), .B(new_n5129_), .ZN(new_n5250_));
  NAND2_X1   g04994(.A1(new_n5250_), .A2(new_n5249_), .ZN(new_n5251_));
  NAND2_X1   g04995(.A1(new_n5248_), .A2(new_n5251_), .ZN(new_n5252_));
  AOI21_X1   g04996(.A1(new_n5252_), .A2(new_n5247_), .B(new_n5122_), .ZN(new_n5253_));
  NOR2_X1    g04997(.A1(new_n5248_), .A2(new_n5251_), .ZN(new_n5254_));
  AOI21_X1   g04998(.A1(new_n4995_), .A2(new_n5006_), .B(new_n5004_), .ZN(new_n5255_));
  NOR2_X1    g04999(.A1(new_n5255_), .A2(new_n5246_), .ZN(new_n5256_));
  NOR3_X1    g05000(.A1(new_n5256_), .A2(new_n5254_), .A3(new_n5121_), .ZN(new_n5257_));
  NOR2_X1    g05001(.A1(new_n5257_), .A2(new_n5253_), .ZN(new_n5258_));
  NOR3_X1    g05002(.A1(new_n5117_), .A2(new_n5258_), .A3(new_n5033_), .ZN(new_n5259_));
  AOI21_X1   g05003(.A1(new_n5010_), .A2(new_n5022_), .B(new_n5033_), .ZN(new_n5260_));
  OAI21_X1   g05004(.A1(new_n5256_), .A2(new_n5254_), .B(new_n5121_), .ZN(new_n5261_));
  NAND3_X1   g05005(.A1(new_n5252_), .A2(new_n5247_), .A3(new_n5122_), .ZN(new_n5262_));
  NAND2_X1   g05006(.A1(new_n5261_), .A2(new_n5262_), .ZN(new_n5263_));
  NOR2_X1    g05007(.A1(new_n5260_), .A2(new_n5263_), .ZN(new_n5264_));
  OAI21_X1   g05008(.A1(new_n5264_), .A2(new_n5259_), .B(new_n5116_), .ZN(new_n5265_));
  INV_X1     g05009(.I(new_n5265_), .ZN(new_n5266_));
  NOR3_X1    g05010(.A1(new_n5264_), .A2(new_n5259_), .A3(new_n5116_), .ZN(new_n5267_));
  NOR2_X1    g05011(.A1(new_n5266_), .A2(new_n5267_), .ZN(new_n5268_));
  NOR2_X1    g05012(.A1(new_n5111_), .A2(new_n5268_), .ZN(new_n5269_));
  AOI21_X1   g05013(.A1(new_n4836_), .A2(new_n5043_), .B(new_n5046_), .ZN(new_n5270_));
  OAI21_X1   g05014(.A1(new_n5036_), .A2(new_n5270_), .B(new_n5047_), .ZN(new_n5271_));
  INV_X1     g05015(.I(new_n5267_), .ZN(new_n5272_));
  NAND2_X1   g05016(.A1(new_n5272_), .A2(new_n5265_), .ZN(new_n5273_));
  NOR2_X1    g05017(.A1(new_n5273_), .A2(new_n5271_), .ZN(new_n5274_));
  OAI22_X1   g05018(.A1(new_n713_), .A2(new_n3185_), .B1(new_n3158_), .B2(new_n717_), .ZN(new_n5275_));
  AOI21_X1   g05019(.A1(\b[26] ), .A2(new_n1126_), .B(new_n5275_), .ZN(new_n5276_));
  OAI21_X1   g05020(.A1(new_n3196_), .A2(new_n986_), .B(new_n5276_), .ZN(new_n5277_));
  XOR2_X1    g05021(.A1(new_n5277_), .A2(\a[11] ), .Z(new_n5278_));
  INV_X1     g05022(.I(new_n5278_), .ZN(new_n5279_));
  OAI21_X1   g05023(.A1(new_n5269_), .A2(new_n5274_), .B(new_n5279_), .ZN(new_n5280_));
  OR3_X2     g05024(.A1(new_n5269_), .A2(new_n5274_), .A3(new_n5279_), .Z(new_n5281_));
  NAND2_X1   g05025(.A1(new_n5281_), .A2(new_n5280_), .ZN(new_n5282_));
  NOR2_X1    g05026(.A1(new_n5282_), .A2(new_n5109_), .ZN(new_n5283_));
  OAI21_X1   g05027(.A1(new_n5065_), .A2(new_n5061_), .B(new_n5067_), .ZN(new_n5284_));
  INV_X1     g05028(.I(new_n5280_), .ZN(new_n5285_));
  NOR3_X1    g05029(.A1(new_n5269_), .A2(new_n5274_), .A3(new_n5279_), .ZN(new_n5286_));
  NOR2_X1    g05030(.A1(new_n5285_), .A2(new_n5286_), .ZN(new_n5287_));
  NOR2_X1    g05031(.A1(new_n5287_), .A2(new_n5284_), .ZN(new_n5288_));
  AOI22_X1   g05032(.A1(new_n518_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n636_), .ZN(new_n5289_));
  OAI21_X1   g05033(.A1(new_n3592_), .A2(new_n917_), .B(new_n5289_), .ZN(new_n5290_));
  AOI21_X1   g05034(.A1(new_n3796_), .A2(new_n618_), .B(new_n5290_), .ZN(new_n5291_));
  XOR2_X1    g05035(.A1(new_n5291_), .A2(new_n488_), .Z(new_n5292_));
  OAI21_X1   g05036(.A1(new_n5288_), .A2(new_n5283_), .B(new_n5292_), .ZN(new_n5293_));
  NAND2_X1   g05037(.A1(new_n5287_), .A2(new_n5284_), .ZN(new_n5294_));
  NAND2_X1   g05038(.A1(new_n5282_), .A2(new_n5109_), .ZN(new_n5295_));
  XOR2_X1    g05039(.A1(new_n5291_), .A2(\a[8] ), .Z(new_n5296_));
  NAND3_X1   g05040(.A1(new_n5294_), .A2(new_n5296_), .A3(new_n5295_), .ZN(new_n5297_));
  NAND2_X1   g05041(.A1(new_n5293_), .A2(new_n5297_), .ZN(new_n5298_));
  NOR2_X1    g05042(.A1(new_n5108_), .A2(new_n5298_), .ZN(new_n5299_));
  OAI21_X1   g05043(.A1(new_n5069_), .A2(new_n5078_), .B(new_n5084_), .ZN(new_n5300_));
  AOI21_X1   g05044(.A1(new_n5294_), .A2(new_n5295_), .B(new_n5296_), .ZN(new_n5301_));
  NOR3_X1    g05045(.A1(new_n5288_), .A2(new_n5292_), .A3(new_n5283_), .ZN(new_n5302_));
  NOR2_X1    g05046(.A1(new_n5301_), .A2(new_n5302_), .ZN(new_n5303_));
  NOR2_X1    g05047(.A1(new_n5300_), .A2(new_n5303_), .ZN(new_n5304_));
  NOR3_X1    g05048(.A1(new_n5299_), .A2(new_n5304_), .A3(new_n5107_), .ZN(new_n5305_));
  XOR2_X1    g05049(.A1(new_n5106_), .A2(new_n312_), .Z(new_n5306_));
  NAND2_X1   g05050(.A1(new_n5300_), .A2(new_n5303_), .ZN(new_n5307_));
  NAND2_X1   g05051(.A1(new_n5108_), .A2(new_n5298_), .ZN(new_n5308_));
  AOI21_X1   g05052(.A1(new_n5308_), .A2(new_n5307_), .B(new_n5306_), .ZN(new_n5309_));
  NOR2_X1    g05053(.A1(new_n5309_), .A2(new_n5305_), .ZN(new_n5310_));
  XOR2_X1    g05054(.A1(new_n5102_), .A2(new_n5310_), .Z(new_n5311_));
  INV_X1     g05055(.I(\b[37] ), .ZN(new_n5312_));
  OAI22_X1   g05056(.A1(new_n277_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n262_), .ZN(new_n5313_));
  AOI21_X1   g05057(.A1(\b[35] ), .A2(new_n283_), .B(new_n5313_), .ZN(new_n5314_));
  AOI21_X1   g05058(.A1(new_n4896_), .A2(\b[36] ), .B(new_n4666_), .ZN(new_n5315_));
  NOR2_X1    g05059(.A1(new_n4896_), .A2(\b[36] ), .ZN(new_n5316_));
  NAND3_X1   g05060(.A1(new_n4894_), .A2(new_n4895_), .A3(new_n5312_), .ZN(new_n5317_));
  INV_X1     g05061(.I(new_n5317_), .ZN(new_n5318_));
  NOR2_X1    g05062(.A1(new_n4891_), .A2(new_n5312_), .ZN(new_n5319_));
  OAI22_X1   g05063(.A1(new_n5315_), .A2(new_n5316_), .B1(new_n5318_), .B2(new_n5319_), .ZN(new_n5320_));
  OR4_X2     g05064(.A1(new_n5315_), .A2(new_n5316_), .A3(new_n5318_), .A4(new_n5319_), .Z(new_n5321_));
  NAND2_X1   g05065(.A1(new_n5321_), .A2(new_n5320_), .ZN(new_n5322_));
  OAI21_X1   g05066(.A1(new_n5322_), .A2(new_n279_), .B(new_n5314_), .ZN(new_n5323_));
  XOR2_X1    g05067(.A1(new_n5323_), .A2(\a[2] ), .Z(new_n5324_));
  INV_X1     g05068(.I(new_n4900_), .ZN(new_n5325_));
  NOR2_X1    g05069(.A1(new_n5090_), .A2(new_n5325_), .ZN(new_n5326_));
  AOI22_X1   g05070(.A1(new_n4880_), .A2(new_n4884_), .B1(new_n5091_), .B2(new_n5096_), .ZN(new_n5327_));
  OAI21_X1   g05071(.A1(new_n5327_), .A2(new_n5326_), .B(new_n5324_), .ZN(new_n5328_));
  INV_X1     g05072(.I(new_n5324_), .ZN(new_n5329_));
  INV_X1     g05073(.I(new_n5326_), .ZN(new_n5330_));
  NOR3_X1    g05074(.A1(new_n4664_), .A2(new_n4661_), .A3(new_n4874_), .ZN(new_n5331_));
  NAND2_X1   g05075(.A1(new_n5093_), .A2(new_n5094_), .ZN(new_n5332_));
  NOR2_X1    g05076(.A1(new_n5332_), .A2(new_n5325_), .ZN(new_n5333_));
  OAI22_X1   g05077(.A1(new_n5331_), .A2(new_n4877_), .B1(new_n5333_), .B2(new_n5095_), .ZN(new_n5334_));
  NAND3_X1   g05078(.A1(new_n5334_), .A2(new_n5329_), .A3(new_n5330_), .ZN(new_n5335_));
  NAND2_X1   g05079(.A1(new_n5328_), .A2(new_n5335_), .ZN(new_n5336_));
  XOR2_X1    g05080(.A1(new_n5336_), .A2(new_n5311_), .Z(\f[37] ));
  INV_X1     g05081(.I(new_n5311_), .ZN(new_n5338_));
  AOI21_X1   g05082(.A1(new_n5334_), .A2(new_n5330_), .B(new_n5329_), .ZN(new_n5339_));
  OAI21_X1   g05083(.A1(new_n5338_), .A2(new_n5339_), .B(new_n5335_), .ZN(new_n5340_));
  INV_X1     g05084(.I(\b[38] ), .ZN(new_n5341_));
  OAI22_X1   g05085(.A1(new_n277_), .A2(new_n5341_), .B1(new_n5312_), .B2(new_n262_), .ZN(new_n5342_));
  AOI21_X1   g05086(.A1(\b[36] ), .A2(new_n283_), .B(new_n5342_), .ZN(new_n5343_));
  AOI21_X1   g05087(.A1(new_n5317_), .A2(\b[36] ), .B(\b[35] ), .ZN(new_n5344_));
  AOI21_X1   g05088(.A1(new_n4896_), .A2(\b[37] ), .B(\b[36] ), .ZN(new_n5345_));
  NOR2_X1    g05089(.A1(new_n5344_), .A2(new_n5345_), .ZN(new_n5346_));
  XNOR2_X1   g05090(.A1(\b[37] ), .A2(\b[38] ), .ZN(new_n5347_));
  XOR2_X1    g05091(.A1(\b[37] ), .A2(\b[38] ), .Z(new_n5348_));
  INV_X1     g05092(.I(new_n5348_), .ZN(new_n5349_));
  NAND2_X1   g05093(.A1(new_n5346_), .A2(new_n5349_), .ZN(new_n5350_));
  OAI21_X1   g05094(.A1(new_n5346_), .A2(new_n5347_), .B(new_n5350_), .ZN(new_n5351_));
  INV_X1     g05095(.I(new_n5351_), .ZN(new_n5352_));
  OAI21_X1   g05096(.A1(new_n5352_), .A2(new_n279_), .B(new_n5343_), .ZN(new_n5353_));
  XOR2_X1    g05097(.A1(new_n5353_), .A2(new_n270_), .Z(new_n5354_));
  INV_X1     g05098(.I(new_n5354_), .ZN(new_n5355_));
  OAI21_X1   g05099(.A1(new_n4855_), .A2(new_n4858_), .B(new_n5072_), .ZN(new_n5356_));
  AOI21_X1   g05100(.A1(new_n5356_), .A2(new_n5076_), .B(new_n5069_), .ZN(new_n5357_));
  OAI21_X1   g05101(.A1(new_n5357_), .A2(new_n5081_), .B(new_n5293_), .ZN(new_n5358_));
  AOI22_X1   g05102(.A1(new_n518_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n636_), .ZN(new_n5359_));
  OAI21_X1   g05103(.A1(new_n3624_), .A2(new_n917_), .B(new_n5359_), .ZN(new_n5360_));
  AOI21_X1   g05104(.A1(new_n4030_), .A2(new_n618_), .B(new_n5360_), .ZN(new_n5361_));
  XOR2_X1    g05105(.A1(new_n5361_), .A2(new_n488_), .Z(new_n5362_));
  INV_X1     g05106(.I(new_n5362_), .ZN(new_n5363_));
  OAI21_X1   g05107(.A1(new_n4363_), .A2(new_n4358_), .B(new_n4365_), .ZN(new_n5364_));
  AOI21_X1   g05108(.A1(new_n5364_), .A2(new_n4842_), .B(new_n4576_), .ZN(new_n5365_));
  AOI21_X1   g05109(.A1(new_n5365_), .A2(new_n4839_), .B(new_n4835_), .ZN(new_n5366_));
  OAI21_X1   g05110(.A1(new_n5366_), .A2(new_n5059_), .B(new_n5054_), .ZN(new_n5367_));
  AOI21_X1   g05111(.A1(new_n5367_), .A2(new_n5067_), .B(new_n5286_), .ZN(new_n5368_));
  INV_X1     g05112(.I(new_n4188_), .ZN(new_n5369_));
  OAI22_X1   g05113(.A1(new_n713_), .A2(new_n3592_), .B1(new_n3185_), .B2(new_n717_), .ZN(new_n5370_));
  AOI21_X1   g05114(.A1(\b[27] ), .A2(new_n1126_), .B(new_n5370_), .ZN(new_n5371_));
  OAI21_X1   g05115(.A1(new_n5369_), .A2(new_n986_), .B(new_n5371_), .ZN(new_n5372_));
  XOR2_X1    g05116(.A1(new_n5372_), .A2(\a[11] ), .Z(new_n5373_));
  AOI21_X1   g05117(.A1(new_n4584_), .A2(new_n4568_), .B(new_n4564_), .ZN(new_n5374_));
  OAI21_X1   g05118(.A1(new_n5374_), .A2(new_n4829_), .B(new_n5043_), .ZN(new_n5375_));
  AOI21_X1   g05119(.A1(new_n5375_), .A2(new_n5040_), .B(new_n5036_), .ZN(new_n5376_));
  OAI21_X1   g05120(.A1(new_n5376_), .A2(new_n5110_), .B(new_n5272_), .ZN(new_n5377_));
  OAI22_X1   g05121(.A1(new_n993_), .A2(new_n3006_), .B1(new_n2646_), .B2(new_n997_), .ZN(new_n5378_));
  AOI21_X1   g05122(.A1(\b[24] ), .A2(new_n1486_), .B(new_n5378_), .ZN(new_n5379_));
  OAI21_X1   g05123(.A1(new_n3016_), .A2(new_n1323_), .B(new_n5379_), .ZN(new_n5380_));
  XOR2_X1    g05124(.A1(new_n5380_), .A2(\a[14] ), .Z(new_n5381_));
  INV_X1     g05125(.I(new_n5381_), .ZN(new_n5382_));
  OAI21_X1   g05126(.A1(new_n4421_), .A2(new_n4335_), .B(new_n4555_), .ZN(new_n5383_));
  OAI21_X1   g05127(.A1(new_n5383_), .A2(new_n4553_), .B(new_n4805_), .ZN(new_n5384_));
  AOI21_X1   g05128(.A1(new_n5384_), .A2(new_n5027_), .B(new_n5015_), .ZN(new_n5385_));
  OAI21_X1   g05129(.A1(new_n5385_), .A2(new_n5023_), .B(new_n5010_), .ZN(new_n5386_));
  NAND3_X1   g05130(.A1(new_n5386_), .A2(new_n5263_), .A3(new_n5029_), .ZN(new_n5387_));
  NOR3_X1    g05131(.A1(new_n5256_), .A2(new_n5254_), .A3(new_n5122_), .ZN(new_n5388_));
  INV_X1     g05132(.I(new_n5388_), .ZN(new_n5389_));
  OAI22_X1   g05133(.A1(new_n1592_), .A2(new_n2463_), .B1(new_n2142_), .B2(new_n1505_), .ZN(new_n5390_));
  AOI21_X1   g05134(.A1(\b[21] ), .A2(new_n1584_), .B(new_n5390_), .ZN(new_n5391_));
  OAI21_X1   g05135(.A1(new_n3552_), .A2(new_n1732_), .B(new_n5391_), .ZN(new_n5392_));
  XOR2_X1    g05136(.A1(new_n5392_), .A2(\a[17] ), .Z(new_n5393_));
  AOI22_X1   g05137(.A1(new_n1738_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n1743_), .ZN(new_n5394_));
  OAI21_X1   g05138(.A1(new_n1553_), .A2(new_n1931_), .B(new_n5394_), .ZN(new_n5395_));
  AOI21_X1   g05139(.A1(new_n2452_), .A2(new_n1746_), .B(new_n5395_), .ZN(new_n5396_));
  XOR2_X1    g05140(.A1(new_n5396_), .A2(new_n1736_), .Z(new_n5397_));
  OAI22_X1   g05141(.A1(new_n2189_), .A2(new_n1432_), .B1(new_n1296_), .B2(new_n2194_), .ZN(new_n5398_));
  AOI21_X1   g05142(.A1(\b[15] ), .A2(new_n2361_), .B(new_n5398_), .ZN(new_n5399_));
  OAI21_X1   g05143(.A1(new_n1444_), .A2(new_n2197_), .B(new_n5399_), .ZN(new_n5400_));
  XOR2_X1    g05144(.A1(new_n5400_), .A2(\a[23] ), .Z(new_n5401_));
  NOR2_X1    g05145(.A1(new_n4975_), .A2(new_n4967_), .ZN(new_n5402_));
  OAI21_X1   g05146(.A1(new_n5402_), .A2(new_n4976_), .B(new_n5218_), .ZN(new_n5403_));
  OAI22_X1   g05147(.A1(new_n852_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n776_), .ZN(new_n5404_));
  AOI21_X1   g05148(.A1(\b[9] ), .A2(new_n3456_), .B(new_n5404_), .ZN(new_n5405_));
  OAI21_X1   g05149(.A1(new_n859_), .A2(new_n3261_), .B(new_n5405_), .ZN(new_n5406_));
  XOR2_X1    g05150(.A1(new_n5406_), .A2(\a[29] ), .Z(new_n5407_));
  NOR2_X1    g05151(.A1(new_n5195_), .A2(new_n5190_), .ZN(new_n5408_));
  AOI21_X1   g05152(.A1(new_n5199_), .A2(new_n5196_), .B(new_n5408_), .ZN(new_n5409_));
  INV_X1     g05153(.I(new_n4053_), .ZN(new_n5410_));
  AOI22_X1   g05154(.A1(new_n3864_), .A2(\b[8] ), .B1(\b[7] ), .B2(new_n3869_), .ZN(new_n5411_));
  OAI21_X1   g05155(.A1(new_n438_), .A2(new_n5410_), .B(new_n5411_), .ZN(new_n5412_));
  AOI21_X1   g05156(.A1(new_n799_), .A2(new_n3872_), .B(new_n5412_), .ZN(new_n5413_));
  XOR2_X1    g05157(.A1(new_n5413_), .A2(new_n3876_), .Z(new_n5414_));
  NAND2_X1   g05158(.A1(new_n5166_), .A2(new_n554_), .ZN(new_n5415_));
  AOI22_X1   g05159(.A1(new_n5155_), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n5160_), .ZN(new_n5416_));
  XOR2_X1    g05160(.A1(\a[35] ), .A2(\a[36] ), .Z(new_n5417_));
  NOR2_X1    g05161(.A1(new_n5163_), .A2(\a[35] ), .ZN(new_n5418_));
  AOI21_X1   g05162(.A1(\a[37] ), .A2(new_n5162_), .B(new_n4446_), .ZN(new_n5419_));
  NOR3_X1    g05163(.A1(new_n5418_), .A2(new_n5417_), .A3(new_n5419_), .ZN(new_n5420_));
  NAND2_X1   g05164(.A1(new_n5420_), .A2(\b[0] ), .ZN(new_n5421_));
  NAND3_X1   g05165(.A1(new_n5416_), .A2(new_n5421_), .A3(new_n5415_), .ZN(new_n5422_));
  XOR2_X1    g05166(.A1(new_n5422_), .A2(new_n5162_), .Z(new_n5423_));
  NOR3_X1    g05167(.A1(new_n5168_), .A2(new_n5162_), .A3(new_n4927_), .ZN(new_n5424_));
  INV_X1     g05168(.I(new_n5424_), .ZN(new_n5425_));
  NAND2_X1   g05169(.A1(new_n5423_), .A2(new_n5425_), .ZN(new_n5426_));
  OR4_X2     g05170(.A1(new_n5162_), .A2(new_n5422_), .A3(new_n4927_), .A4(new_n5168_), .Z(new_n5427_));
  OAI22_X1   g05171(.A1(new_n377_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n339_), .ZN(new_n5428_));
  AOI21_X1   g05172(.A1(\b[3] ), .A2(new_n4706_), .B(new_n5428_), .ZN(new_n5429_));
  OAI21_X1   g05173(.A1(new_n566_), .A2(new_n4458_), .B(new_n5429_), .ZN(new_n5430_));
  XOR2_X1    g05174(.A1(new_n5430_), .A2(\a[35] ), .Z(new_n5431_));
  AOI21_X1   g05175(.A1(new_n5426_), .A2(new_n5427_), .B(new_n5431_), .ZN(new_n5432_));
  NAND2_X1   g05176(.A1(new_n5426_), .A2(new_n5427_), .ZN(new_n5433_));
  XOR2_X1    g05177(.A1(new_n5430_), .A2(new_n4446_), .Z(new_n5434_));
  NOR2_X1    g05178(.A1(new_n5433_), .A2(new_n5434_), .ZN(new_n5435_));
  NOR2_X1    g05179(.A1(new_n5432_), .A2(new_n5435_), .ZN(new_n5436_));
  OAI21_X1   g05180(.A1(new_n5147_), .A2(new_n5184_), .B(new_n5177_), .ZN(new_n5437_));
  NAND2_X1   g05181(.A1(new_n5436_), .A2(new_n5437_), .ZN(new_n5438_));
  NAND2_X1   g05182(.A1(new_n5433_), .A2(new_n5434_), .ZN(new_n5439_));
  NAND3_X1   g05183(.A1(new_n5431_), .A2(new_n5426_), .A3(new_n5427_), .ZN(new_n5440_));
  NAND2_X1   g05184(.A1(new_n5439_), .A2(new_n5440_), .ZN(new_n5441_));
  AOI21_X1   g05185(.A1(new_n5182_), .A2(new_n5178_), .B(new_n5183_), .ZN(new_n5442_));
  NAND2_X1   g05186(.A1(new_n5441_), .A2(new_n5442_), .ZN(new_n5443_));
  NAND3_X1   g05187(.A1(new_n5438_), .A2(new_n5443_), .A3(new_n5414_), .ZN(new_n5444_));
  INV_X1     g05188(.I(new_n5414_), .ZN(new_n5445_));
  NOR2_X1    g05189(.A1(new_n5441_), .A2(new_n5442_), .ZN(new_n5446_));
  NOR2_X1    g05190(.A1(new_n5436_), .A2(new_n5437_), .ZN(new_n5447_));
  OAI21_X1   g05191(.A1(new_n5447_), .A2(new_n5446_), .B(new_n5445_), .ZN(new_n5448_));
  NAND3_X1   g05192(.A1(new_n5409_), .A2(new_n5444_), .A3(new_n5448_), .ZN(new_n5449_));
  NOR2_X1    g05193(.A1(new_n5186_), .A2(new_n5191_), .ZN(new_n5450_));
  OAI21_X1   g05194(.A1(new_n5144_), .A2(new_n5450_), .B(new_n5192_), .ZN(new_n5451_));
  NAND2_X1   g05195(.A1(new_n5448_), .A2(new_n5444_), .ZN(new_n5452_));
  NAND2_X1   g05196(.A1(new_n5452_), .A2(new_n5451_), .ZN(new_n5453_));
  AOI21_X1   g05197(.A1(new_n5449_), .A2(new_n5453_), .B(new_n5407_), .ZN(new_n5454_));
  XOR2_X1    g05198(.A1(new_n5406_), .A2(new_n3264_), .Z(new_n5455_));
  NOR2_X1    g05199(.A1(new_n5452_), .A2(new_n5451_), .ZN(new_n5456_));
  AOI21_X1   g05200(.A1(new_n5444_), .A2(new_n5448_), .B(new_n5409_), .ZN(new_n5457_));
  NOR3_X1    g05201(.A1(new_n5457_), .A2(new_n5456_), .A3(new_n5455_), .ZN(new_n5458_));
  NOR2_X1    g05202(.A1(new_n5458_), .A2(new_n5454_), .ZN(new_n5459_));
  AOI21_X1   g05203(.A1(new_n4961_), .A2(new_n4947_), .B(new_n4942_), .ZN(new_n5460_));
  OAI21_X1   g05204(.A1(new_n5460_), .A2(new_n4962_), .B(new_n5209_), .ZN(new_n5461_));
  NAND3_X1   g05205(.A1(new_n5459_), .A2(new_n5461_), .A3(new_n5206_), .ZN(new_n5462_));
  INV_X1     g05206(.I(new_n5206_), .ZN(new_n5463_));
  OAI21_X1   g05207(.A1(new_n5457_), .A2(new_n5456_), .B(new_n5455_), .ZN(new_n5464_));
  NAND3_X1   g05208(.A1(new_n5449_), .A2(new_n5453_), .A3(new_n5407_), .ZN(new_n5465_));
  NAND2_X1   g05209(.A1(new_n5464_), .A2(new_n5465_), .ZN(new_n5466_));
  AOI21_X1   g05210(.A1(new_n5198_), .A2(new_n5200_), .B(new_n5205_), .ZN(new_n5467_));
  AOI21_X1   g05211(.A1(new_n5137_), .A2(new_n4965_), .B(new_n5467_), .ZN(new_n5468_));
  OAI21_X1   g05212(.A1(new_n5468_), .A2(new_n5463_), .B(new_n5466_), .ZN(new_n5469_));
  AOI22_X1   g05213(.A1(new_n2716_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n2719_), .ZN(new_n5470_));
  OAI21_X1   g05214(.A1(new_n941_), .A2(new_n2924_), .B(new_n5470_), .ZN(new_n5471_));
  AOI21_X1   g05215(.A1(new_n1449_), .A2(new_n2722_), .B(new_n5471_), .ZN(new_n5472_));
  XOR2_X1    g05216(.A1(new_n5472_), .A2(new_n2714_), .Z(new_n5473_));
  NAND3_X1   g05217(.A1(new_n5469_), .A2(new_n5462_), .A3(new_n5473_), .ZN(new_n5474_));
  INV_X1     g05218(.I(new_n5474_), .ZN(new_n5475_));
  AOI21_X1   g05219(.A1(new_n5469_), .A2(new_n5462_), .B(new_n5473_), .ZN(new_n5476_));
  NOR2_X1    g05220(.A1(new_n5475_), .A2(new_n5476_), .ZN(new_n5477_));
  NAND3_X1   g05221(.A1(new_n5403_), .A2(new_n5477_), .A3(new_n5222_), .ZN(new_n5478_));
  AOI21_X1   g05222(.A1(new_n5136_), .A2(new_n4979_), .B(new_n5226_), .ZN(new_n5479_));
  INV_X1     g05223(.I(new_n5476_), .ZN(new_n5480_));
  NAND2_X1   g05224(.A1(new_n5480_), .A2(new_n5474_), .ZN(new_n5481_));
  OAI21_X1   g05225(.A1(new_n5479_), .A2(new_n5227_), .B(new_n5481_), .ZN(new_n5482_));
  AOI21_X1   g05226(.A1(new_n5482_), .A2(new_n5478_), .B(new_n5401_), .ZN(new_n5483_));
  INV_X1     g05227(.I(new_n5401_), .ZN(new_n5484_));
  NOR3_X1    g05228(.A1(new_n5479_), .A2(new_n5481_), .A3(new_n5227_), .ZN(new_n5485_));
  AOI21_X1   g05229(.A1(new_n5225_), .A2(new_n5218_), .B(new_n5227_), .ZN(new_n5486_));
  NOR2_X1    g05230(.A1(new_n5486_), .A2(new_n5477_), .ZN(new_n5487_));
  NOR3_X1    g05231(.A1(new_n5487_), .A2(new_n5485_), .A3(new_n5484_), .ZN(new_n5488_));
  NOR2_X1    g05232(.A1(new_n5488_), .A2(new_n5483_), .ZN(new_n5489_));
  AOI21_X1   g05233(.A1(new_n5231_), .A2(new_n5232_), .B(new_n5135_), .ZN(new_n5490_));
  INV_X1     g05234(.I(new_n5490_), .ZN(new_n5491_));
  OAI21_X1   g05235(.A1(new_n5130_), .A2(new_n5234_), .B(new_n5491_), .ZN(new_n5492_));
  NAND2_X1   g05236(.A1(new_n5492_), .A2(new_n5489_), .ZN(new_n5493_));
  OAI21_X1   g05237(.A1(new_n5487_), .A2(new_n5485_), .B(new_n5484_), .ZN(new_n5494_));
  NAND3_X1   g05238(.A1(new_n5482_), .A2(new_n5478_), .A3(new_n5401_), .ZN(new_n5495_));
  NAND2_X1   g05239(.A1(new_n5494_), .A2(new_n5495_), .ZN(new_n5496_));
  NAND3_X1   g05240(.A1(new_n5243_), .A2(new_n5496_), .A3(new_n5491_), .ZN(new_n5497_));
  AOI21_X1   g05241(.A1(new_n5493_), .A2(new_n5497_), .B(new_n5397_), .ZN(new_n5498_));
  INV_X1     g05242(.I(new_n5397_), .ZN(new_n5499_));
  AOI21_X1   g05243(.A1(new_n5243_), .A2(new_n5491_), .B(new_n5496_), .ZN(new_n5500_));
  NOR2_X1    g05244(.A1(new_n5492_), .A2(new_n5489_), .ZN(new_n5501_));
  NOR3_X1    g05245(.A1(new_n5501_), .A2(new_n5500_), .A3(new_n5499_), .ZN(new_n5502_));
  NOR2_X1    g05246(.A1(new_n5502_), .A2(new_n5498_), .ZN(new_n5503_));
  OAI21_X1   g05247(.A1(new_n5248_), .A2(new_n5251_), .B(new_n5249_), .ZN(new_n5504_));
  NAND2_X1   g05248(.A1(new_n5504_), .A2(new_n5503_), .ZN(new_n5505_));
  OAI21_X1   g05249(.A1(new_n5501_), .A2(new_n5500_), .B(new_n5499_), .ZN(new_n5506_));
  NAND3_X1   g05250(.A1(new_n5493_), .A2(new_n5497_), .A3(new_n5397_), .ZN(new_n5507_));
  NAND2_X1   g05251(.A1(new_n5506_), .A2(new_n5507_), .ZN(new_n5508_));
  NAND3_X1   g05252(.A1(new_n5247_), .A2(new_n5508_), .A3(new_n5249_), .ZN(new_n5509_));
  NAND3_X1   g05253(.A1(new_n5505_), .A2(new_n5509_), .A3(new_n5393_), .ZN(new_n5510_));
  INV_X1     g05254(.I(new_n5393_), .ZN(new_n5511_));
  AOI21_X1   g05255(.A1(new_n5247_), .A2(new_n5249_), .B(new_n5508_), .ZN(new_n5512_));
  NOR2_X1    g05256(.A1(new_n5504_), .A2(new_n5503_), .ZN(new_n5513_));
  OAI21_X1   g05257(.A1(new_n5513_), .A2(new_n5512_), .B(new_n5511_), .ZN(new_n5514_));
  NAND2_X1   g05258(.A1(new_n5514_), .A2(new_n5510_), .ZN(new_n5515_));
  AOI21_X1   g05259(.A1(new_n5387_), .A2(new_n5389_), .B(new_n5515_), .ZN(new_n5516_));
  OAI21_X1   g05260(.A1(new_n5009_), .A2(new_n5032_), .B(new_n5029_), .ZN(new_n5517_));
  OAI21_X1   g05261(.A1(new_n5517_), .A2(new_n5258_), .B(new_n5389_), .ZN(new_n5518_));
  NOR3_X1    g05262(.A1(new_n5513_), .A2(new_n5512_), .A3(new_n5511_), .ZN(new_n5519_));
  AOI21_X1   g05263(.A1(new_n5505_), .A2(new_n5509_), .B(new_n5393_), .ZN(new_n5520_));
  NOR2_X1    g05264(.A1(new_n5519_), .A2(new_n5520_), .ZN(new_n5521_));
  NOR2_X1    g05265(.A1(new_n5518_), .A2(new_n5521_), .ZN(new_n5522_));
  NOR3_X1    g05266(.A1(new_n5522_), .A2(new_n5516_), .A3(new_n5382_), .ZN(new_n5523_));
  OAI21_X1   g05267(.A1(new_n5259_), .A2(new_n5388_), .B(new_n5521_), .ZN(new_n5524_));
  NAND3_X1   g05268(.A1(new_n5387_), .A2(new_n5515_), .A3(new_n5389_), .ZN(new_n5525_));
  AOI21_X1   g05269(.A1(new_n5524_), .A2(new_n5525_), .B(new_n5381_), .ZN(new_n5526_));
  NOR2_X1    g05270(.A1(new_n5523_), .A2(new_n5526_), .ZN(new_n5527_));
  NAND3_X1   g05271(.A1(new_n5377_), .A2(new_n5527_), .A3(new_n5265_), .ZN(new_n5528_));
  OAI21_X1   g05272(.A1(new_n4571_), .A2(new_n4574_), .B(new_n4572_), .ZN(new_n5529_));
  AOI21_X1   g05273(.A1(new_n5529_), .A2(new_n4833_), .B(new_n5044_), .ZN(new_n5530_));
  OAI21_X1   g05274(.A1(new_n5530_), .A2(new_n5046_), .B(new_n5051_), .ZN(new_n5531_));
  AOI21_X1   g05275(.A1(new_n5531_), .A2(new_n5047_), .B(new_n5267_), .ZN(new_n5532_));
  NAND3_X1   g05276(.A1(new_n5524_), .A2(new_n5525_), .A3(new_n5381_), .ZN(new_n5533_));
  OAI21_X1   g05277(.A1(new_n5522_), .A2(new_n5516_), .B(new_n5382_), .ZN(new_n5534_));
  NAND2_X1   g05278(.A1(new_n5534_), .A2(new_n5533_), .ZN(new_n5535_));
  OAI21_X1   g05279(.A1(new_n5532_), .A2(new_n5266_), .B(new_n5535_), .ZN(new_n5536_));
  NAND3_X1   g05280(.A1(new_n5536_), .A2(new_n5528_), .A3(new_n5373_), .ZN(new_n5537_));
  XOR2_X1    g05281(.A1(new_n5372_), .A2(new_n722_), .Z(new_n5538_));
  NOR3_X1    g05282(.A1(new_n5532_), .A2(new_n5266_), .A3(new_n5535_), .ZN(new_n5539_));
  AOI21_X1   g05283(.A1(new_n5377_), .A2(new_n5265_), .B(new_n5527_), .ZN(new_n5540_));
  OAI21_X1   g05284(.A1(new_n5539_), .A2(new_n5540_), .B(new_n5538_), .ZN(new_n5541_));
  NAND2_X1   g05285(.A1(new_n5541_), .A2(new_n5537_), .ZN(new_n5542_));
  NOR3_X1    g05286(.A1(new_n5368_), .A2(new_n5285_), .A3(new_n5542_), .ZN(new_n5543_));
  AOI21_X1   g05287(.A1(new_n5284_), .A2(new_n5281_), .B(new_n5285_), .ZN(new_n5544_));
  NOR3_X1    g05288(.A1(new_n5539_), .A2(new_n5540_), .A3(new_n5538_), .ZN(new_n5545_));
  AOI21_X1   g05289(.A1(new_n5536_), .A2(new_n5528_), .B(new_n5373_), .ZN(new_n5546_));
  NOR2_X1    g05290(.A1(new_n5545_), .A2(new_n5546_), .ZN(new_n5547_));
  NOR2_X1    g05291(.A1(new_n5544_), .A2(new_n5547_), .ZN(new_n5548_));
  NOR3_X1    g05292(.A1(new_n5548_), .A2(new_n5543_), .A3(new_n5363_), .ZN(new_n5549_));
  OAI21_X1   g05293(.A1(new_n4606_), .A2(new_n4586_), .B(new_n4841_), .ZN(new_n5550_));
  OAI21_X1   g05294(.A1(new_n5550_), .A2(new_n4846_), .B(new_n4844_), .ZN(new_n5551_));
  AOI21_X1   g05295(.A1(new_n5551_), .A2(new_n5058_), .B(new_n5065_), .ZN(new_n5552_));
  OAI21_X1   g05296(.A1(new_n5552_), .A2(new_n5063_), .B(new_n5281_), .ZN(new_n5553_));
  NAND3_X1   g05297(.A1(new_n5553_), .A2(new_n5280_), .A3(new_n5547_), .ZN(new_n5554_));
  OAI21_X1   g05298(.A1(new_n5368_), .A2(new_n5285_), .B(new_n5542_), .ZN(new_n5555_));
  AOI21_X1   g05299(.A1(new_n5554_), .A2(new_n5555_), .B(new_n5362_), .ZN(new_n5556_));
  NOR2_X1    g05300(.A1(new_n5549_), .A2(new_n5556_), .ZN(new_n5557_));
  NAND3_X1   g05301(.A1(new_n5358_), .A2(new_n5557_), .A3(new_n5297_), .ZN(new_n5558_));
  OAI21_X1   g05302(.A1(new_n5108_), .A2(new_n5301_), .B(new_n5297_), .ZN(new_n5559_));
  NAND3_X1   g05303(.A1(new_n5554_), .A2(new_n5555_), .A3(new_n5362_), .ZN(new_n5560_));
  INV_X1     g05304(.I(new_n5556_), .ZN(new_n5561_));
  NAND2_X1   g05305(.A1(new_n5561_), .A2(new_n5560_), .ZN(new_n5562_));
  NAND2_X1   g05306(.A1(new_n5559_), .A2(new_n5562_), .ZN(new_n5563_));
  NAND2_X1   g05307(.A1(new_n5563_), .A2(new_n5558_), .ZN(new_n5564_));
  OAI22_X1   g05308(.A1(new_n321_), .A2(new_n4666_), .B1(new_n325_), .B2(new_n4639_), .ZN(new_n5565_));
  AOI21_X1   g05309(.A1(\b[33] ), .A2(new_n602_), .B(new_n5565_), .ZN(new_n5566_));
  OAI21_X1   g05310(.A1(new_n4676_), .A2(new_n318_), .B(new_n5566_), .ZN(new_n5567_));
  XOR2_X1    g05311(.A1(new_n5567_), .A2(\a[5] ), .Z(new_n5568_));
  INV_X1     g05312(.I(new_n5568_), .ZN(new_n5569_));
  NAND3_X1   g05313(.A1(new_n5084_), .A2(new_n5083_), .A3(new_n5069_), .ZN(new_n5570_));
  OAI21_X1   g05314(.A1(new_n5078_), .A2(new_n5081_), .B(new_n5070_), .ZN(new_n5571_));
  AOI21_X1   g05315(.A1(new_n5571_), .A2(new_n5570_), .B(new_n4907_), .ZN(new_n5572_));
  NOR3_X1    g05316(.A1(new_n4902_), .A2(new_n4870_), .A3(new_n5572_), .ZN(new_n5573_));
  OAI22_X1   g05317(.A1(new_n5573_), .A2(new_n5087_), .B1(new_n5309_), .B2(new_n5305_), .ZN(new_n5574_));
  AOI21_X1   g05318(.A1(new_n5308_), .A2(new_n5307_), .B(new_n5107_), .ZN(new_n5575_));
  INV_X1     g05319(.I(new_n5575_), .ZN(new_n5576_));
  AOI21_X1   g05320(.A1(new_n5574_), .A2(new_n5576_), .B(new_n5569_), .ZN(new_n5577_));
  NAND3_X1   g05321(.A1(new_n5308_), .A2(new_n5307_), .A3(new_n5306_), .ZN(new_n5578_));
  OAI21_X1   g05322(.A1(new_n5299_), .A2(new_n5304_), .B(new_n5107_), .ZN(new_n5579_));
  AOI22_X1   g05323(.A1(new_n5101_), .A2(new_n5088_), .B1(new_n5578_), .B2(new_n5579_), .ZN(new_n5580_));
  NOR3_X1    g05324(.A1(new_n5580_), .A2(new_n5568_), .A3(new_n5575_), .ZN(new_n5581_));
  NOR3_X1    g05325(.A1(new_n5581_), .A2(new_n5577_), .A3(new_n5564_), .ZN(new_n5582_));
  INV_X1     g05326(.I(new_n5564_), .ZN(new_n5583_));
  OAI21_X1   g05327(.A1(new_n5580_), .A2(new_n5575_), .B(new_n5568_), .ZN(new_n5584_));
  NAND3_X1   g05328(.A1(new_n5574_), .A2(new_n5569_), .A3(new_n5576_), .ZN(new_n5585_));
  AOI21_X1   g05329(.A1(new_n5584_), .A2(new_n5585_), .B(new_n5583_), .ZN(new_n5586_));
  NOR2_X1    g05330(.A1(new_n5582_), .A2(new_n5586_), .ZN(new_n5587_));
  NOR2_X1    g05331(.A1(new_n5587_), .A2(new_n5355_), .ZN(new_n5588_));
  INV_X1     g05332(.I(new_n5588_), .ZN(new_n5589_));
  NAND2_X1   g05333(.A1(new_n5587_), .A2(new_n5355_), .ZN(new_n5590_));
  NAND2_X1   g05334(.A1(new_n5589_), .A2(new_n5590_), .ZN(new_n5591_));
  XOR2_X1    g05335(.A1(new_n5340_), .A2(new_n5591_), .Z(\f[38] ));
  AOI21_X1   g05336(.A1(new_n5564_), .A2(new_n5584_), .B(new_n5581_), .ZN(new_n5593_));
  INV_X1     g05337(.I(new_n4898_), .ZN(new_n5594_));
  AOI22_X1   g05338(.A1(new_n800_), .A2(\b[35] ), .B1(\b[36] ), .B2(new_n333_), .ZN(new_n5595_));
  OAI21_X1   g05339(.A1(new_n4639_), .A2(new_n392_), .B(new_n5595_), .ZN(new_n5596_));
  AOI21_X1   g05340(.A1(new_n5594_), .A2(new_n330_), .B(new_n5596_), .ZN(new_n5597_));
  XOR2_X1    g05341(.A1(new_n5597_), .A2(new_n312_), .Z(new_n5598_));
  INV_X1     g05342(.I(new_n5427_), .ZN(new_n5599_));
  NAND2_X1   g05343(.A1(new_n5420_), .A2(\b[1] ), .ZN(new_n5600_));
  AOI22_X1   g05344(.A1(new_n5155_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n5160_), .ZN(new_n5601_));
  NAND2_X1   g05345(.A1(new_n299_), .A2(new_n5166_), .ZN(new_n5602_));
  NAND3_X1   g05346(.A1(new_n5602_), .A2(new_n5601_), .A3(new_n5600_), .ZN(new_n5603_));
  XOR2_X1    g05347(.A1(new_n5603_), .A2(new_n5162_), .Z(new_n5604_));
  XNOR2_X1   g05348(.A1(\a[38] ), .A2(\a[39] ), .ZN(new_n5605_));
  NOR2_X1    g05349(.A1(new_n5605_), .A2(new_n258_), .ZN(new_n5606_));
  INV_X1     g05350(.I(new_n5606_), .ZN(new_n5607_));
  NAND2_X1   g05351(.A1(new_n5604_), .A2(new_n5607_), .ZN(new_n5608_));
  XOR2_X1    g05352(.A1(new_n5603_), .A2(\a[38] ), .Z(new_n5609_));
  NAND2_X1   g05353(.A1(new_n5609_), .A2(new_n5606_), .ZN(new_n5610_));
  NAND2_X1   g05354(.A1(new_n5608_), .A2(new_n5610_), .ZN(new_n5611_));
  XOR2_X1    g05355(.A1(new_n5611_), .A2(new_n5599_), .Z(new_n5612_));
  OAI22_X1   g05356(.A1(new_n438_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n377_), .ZN(new_n5613_));
  AOI21_X1   g05357(.A1(\b[4] ), .A2(new_n4706_), .B(new_n5613_), .ZN(new_n5614_));
  OAI21_X1   g05358(.A1(new_n450_), .A2(new_n4458_), .B(new_n5614_), .ZN(new_n5615_));
  XOR2_X1    g05359(.A1(new_n5615_), .A2(\a[35] ), .Z(new_n5616_));
  OAI21_X1   g05360(.A1(new_n5442_), .A2(new_n5432_), .B(new_n5440_), .ZN(new_n5617_));
  NAND2_X1   g05361(.A1(new_n5617_), .A2(new_n5616_), .ZN(new_n5618_));
  INV_X1     g05362(.I(new_n5616_), .ZN(new_n5619_));
  AOI21_X1   g05363(.A1(new_n5437_), .A2(new_n5439_), .B(new_n5435_), .ZN(new_n5620_));
  NAND2_X1   g05364(.A1(new_n5620_), .A2(new_n5619_), .ZN(new_n5621_));
  NAND3_X1   g05365(.A1(new_n5618_), .A2(new_n5621_), .A3(new_n5612_), .ZN(new_n5622_));
  XOR2_X1    g05366(.A1(new_n5611_), .A2(new_n5427_), .Z(new_n5623_));
  NOR2_X1    g05367(.A1(new_n5620_), .A2(new_n5619_), .ZN(new_n5624_));
  NOR2_X1    g05368(.A1(new_n5617_), .A2(new_n5616_), .ZN(new_n5625_));
  OAI21_X1   g05369(.A1(new_n5625_), .A2(new_n5624_), .B(new_n5623_), .ZN(new_n5626_));
  NAND2_X1   g05370(.A1(new_n5626_), .A2(new_n5622_), .ZN(new_n5627_));
  AOI22_X1   g05371(.A1(new_n3864_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n3869_), .ZN(new_n5628_));
  OAI21_X1   g05372(.A1(new_n471_), .A2(new_n5410_), .B(new_n5628_), .ZN(new_n5629_));
  AOI21_X1   g05373(.A1(new_n676_), .A2(new_n3872_), .B(new_n5629_), .ZN(new_n5630_));
  XOR2_X1    g05374(.A1(new_n5630_), .A2(new_n3876_), .Z(new_n5631_));
  INV_X1     g05375(.I(new_n5631_), .ZN(new_n5632_));
  INV_X1     g05376(.I(new_n5444_), .ZN(new_n5633_));
  AOI21_X1   g05377(.A1(new_n5409_), .A2(new_n5448_), .B(new_n5633_), .ZN(new_n5634_));
  NOR2_X1    g05378(.A1(new_n5634_), .A2(new_n5632_), .ZN(new_n5635_));
  OAI21_X1   g05379(.A1(new_n5452_), .A2(new_n5451_), .B(new_n5444_), .ZN(new_n5636_));
  NOR2_X1    g05380(.A1(new_n5636_), .A2(new_n5631_), .ZN(new_n5637_));
  NOR3_X1    g05381(.A1(new_n5637_), .A2(new_n5635_), .A3(new_n5627_), .ZN(new_n5638_));
  NOR3_X1    g05382(.A1(new_n5625_), .A2(new_n5624_), .A3(new_n5623_), .ZN(new_n5639_));
  AOI21_X1   g05383(.A1(new_n5618_), .A2(new_n5621_), .B(new_n5612_), .ZN(new_n5640_));
  NOR2_X1    g05384(.A1(new_n5639_), .A2(new_n5640_), .ZN(new_n5641_));
  NAND2_X1   g05385(.A1(new_n5636_), .A2(new_n5631_), .ZN(new_n5642_));
  NAND2_X1   g05386(.A1(new_n5634_), .A2(new_n5632_), .ZN(new_n5643_));
  AOI21_X1   g05387(.A1(new_n5642_), .A2(new_n5643_), .B(new_n5641_), .ZN(new_n5644_));
  NOR2_X1    g05388(.A1(new_n5644_), .A2(new_n5638_), .ZN(new_n5645_));
  INV_X1     g05389(.I(new_n5645_), .ZN(new_n5646_));
  NOR3_X1    g05390(.A1(new_n5466_), .A2(new_n5468_), .A3(new_n5463_), .ZN(new_n5647_));
  AOI22_X1   g05391(.A1(new_n3267_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n3270_), .ZN(new_n5648_));
  OAI21_X1   g05392(.A1(new_n776_), .A2(new_n3475_), .B(new_n5648_), .ZN(new_n5649_));
  AOI21_X1   g05393(.A1(new_n1194_), .A2(new_n3273_), .B(new_n5649_), .ZN(new_n5650_));
  XOR2_X1    g05394(.A1(new_n5650_), .A2(new_n3264_), .Z(new_n5651_));
  OAI21_X1   g05395(.A1(new_n5647_), .A2(new_n5458_), .B(new_n5651_), .ZN(new_n5652_));
  INV_X1     g05396(.I(new_n5651_), .ZN(new_n5653_));
  NAND3_X1   g05397(.A1(new_n5462_), .A2(new_n5465_), .A3(new_n5653_), .ZN(new_n5654_));
  NAND2_X1   g05398(.A1(new_n5652_), .A2(new_n5654_), .ZN(new_n5655_));
  XOR2_X1    g05399(.A1(new_n5655_), .A2(new_n5646_), .Z(new_n5656_));
  OAI22_X1   g05400(.A1(new_n2703_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n2708_), .ZN(new_n5657_));
  AOI21_X1   g05401(.A1(\b[13] ), .A2(new_n2906_), .B(new_n5657_), .ZN(new_n5658_));
  OAI21_X1   g05402(.A1(new_n1275_), .A2(new_n2711_), .B(new_n5658_), .ZN(new_n5659_));
  XOR2_X1    g05403(.A1(new_n5659_), .A2(\a[26] ), .Z(new_n5660_));
  OAI21_X1   g05404(.A1(new_n5485_), .A2(new_n5475_), .B(new_n5660_), .ZN(new_n5661_));
  INV_X1     g05405(.I(new_n5660_), .ZN(new_n5662_));
  NAND3_X1   g05406(.A1(new_n5478_), .A2(new_n5474_), .A3(new_n5662_), .ZN(new_n5663_));
  NAND3_X1   g05407(.A1(new_n5661_), .A2(new_n5663_), .A3(new_n5656_), .ZN(new_n5664_));
  INV_X1     g05408(.I(new_n5664_), .ZN(new_n5665_));
  AOI21_X1   g05409(.A1(new_n5661_), .A2(new_n5663_), .B(new_n5656_), .ZN(new_n5666_));
  NOR2_X1    g05410(.A1(new_n5665_), .A2(new_n5666_), .ZN(new_n5667_));
  AOI22_X1   g05411(.A1(new_n2202_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n2205_), .ZN(new_n5668_));
  OAI21_X1   g05412(.A1(new_n1296_), .A2(new_n2370_), .B(new_n5668_), .ZN(new_n5669_));
  AOI21_X1   g05413(.A1(new_n2038_), .A2(new_n2208_), .B(new_n5669_), .ZN(new_n5670_));
  XOR2_X1    g05414(.A1(new_n5670_), .A2(new_n2200_), .Z(new_n5671_));
  OAI21_X1   g05415(.A1(new_n5500_), .A2(new_n5488_), .B(new_n5671_), .ZN(new_n5672_));
  INV_X1     g05416(.I(new_n5671_), .ZN(new_n5673_));
  AOI21_X1   g05417(.A1(new_n5492_), .A2(new_n5489_), .B(new_n5488_), .ZN(new_n5674_));
  NAND2_X1   g05418(.A1(new_n5674_), .A2(new_n5673_), .ZN(new_n5675_));
  NAND3_X1   g05419(.A1(new_n5675_), .A2(new_n5672_), .A3(new_n5667_), .ZN(new_n5676_));
  INV_X1     g05420(.I(new_n5676_), .ZN(new_n5677_));
  AOI21_X1   g05421(.A1(new_n5675_), .A2(new_n5672_), .B(new_n5667_), .ZN(new_n5678_));
  NOR2_X1    g05422(.A1(new_n5677_), .A2(new_n5678_), .ZN(new_n5679_));
  AOI22_X1   g05423(.A1(new_n1738_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n1743_), .ZN(new_n5680_));
  OAI21_X1   g05424(.A1(new_n1859_), .A2(new_n1931_), .B(new_n5680_), .ZN(new_n5681_));
  AOI21_X1   g05425(.A1(new_n2032_), .A2(new_n1746_), .B(new_n5681_), .ZN(new_n5682_));
  XOR2_X1    g05426(.A1(new_n5682_), .A2(new_n1736_), .Z(new_n5683_));
  AOI21_X1   g05427(.A1(new_n5255_), .A2(new_n5246_), .B(new_n5241_), .ZN(new_n5684_));
  OAI21_X1   g05428(.A1(new_n5684_), .A2(new_n5508_), .B(new_n5507_), .ZN(new_n5685_));
  NAND2_X1   g05429(.A1(new_n5685_), .A2(new_n5683_), .ZN(new_n5686_));
  INV_X1     g05430(.I(new_n5683_), .ZN(new_n5687_));
  AOI21_X1   g05431(.A1(new_n5504_), .A2(new_n5503_), .B(new_n5502_), .ZN(new_n5688_));
  NAND2_X1   g05432(.A1(new_n5688_), .A2(new_n5687_), .ZN(new_n5689_));
  NAND3_X1   g05433(.A1(new_n5686_), .A2(new_n5689_), .A3(new_n5679_), .ZN(new_n5690_));
  INV_X1     g05434(.I(new_n5678_), .ZN(new_n5691_));
  NAND2_X1   g05435(.A1(new_n5691_), .A2(new_n5676_), .ZN(new_n5692_));
  NOR2_X1    g05436(.A1(new_n5688_), .A2(new_n5687_), .ZN(new_n5693_));
  NOR2_X1    g05437(.A1(new_n5685_), .A2(new_n5683_), .ZN(new_n5694_));
  OAI21_X1   g05438(.A1(new_n5694_), .A2(new_n5693_), .B(new_n5692_), .ZN(new_n5695_));
  NAND2_X1   g05439(.A1(new_n5695_), .A2(new_n5690_), .ZN(new_n5696_));
  OAI22_X1   g05440(.A1(new_n1592_), .A2(new_n2495_), .B1(new_n2463_), .B2(new_n1505_), .ZN(new_n5697_));
  AOI21_X1   g05441(.A1(\b[22] ), .A2(new_n1584_), .B(new_n5697_), .ZN(new_n5698_));
  OAI21_X1   g05442(.A1(new_n2506_), .A2(new_n1732_), .B(new_n5698_), .ZN(new_n5699_));
  XOR2_X1    g05443(.A1(new_n5699_), .A2(\a[17] ), .Z(new_n5700_));
  INV_X1     g05444(.I(new_n5700_), .ZN(new_n5701_));
  AOI21_X1   g05445(.A1(new_n5524_), .A2(new_n5510_), .B(new_n5701_), .ZN(new_n5702_));
  NOR3_X1    g05446(.A1(new_n5516_), .A2(new_n5519_), .A3(new_n5700_), .ZN(new_n5703_));
  NOR3_X1    g05447(.A1(new_n5702_), .A2(new_n5703_), .A3(new_n5696_), .ZN(new_n5704_));
  INV_X1     g05448(.I(new_n5704_), .ZN(new_n5705_));
  OAI21_X1   g05449(.A1(new_n5702_), .A2(new_n5703_), .B(new_n5696_), .ZN(new_n5706_));
  NAND2_X1   g05450(.A1(new_n5705_), .A2(new_n5706_), .ZN(new_n5707_));
  OAI22_X1   g05451(.A1(new_n993_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n997_), .ZN(new_n5708_));
  AOI21_X1   g05452(.A1(\b[25] ), .A2(new_n1486_), .B(new_n5708_), .ZN(new_n5709_));
  OAI21_X1   g05453(.A1(new_n3165_), .A2(new_n1323_), .B(new_n5709_), .ZN(new_n5710_));
  XOR2_X1    g05454(.A1(new_n5710_), .A2(\a[14] ), .Z(new_n5711_));
  INV_X1     g05455(.I(new_n5711_), .ZN(new_n5712_));
  AOI21_X1   g05456(.A1(new_n5528_), .A2(new_n5533_), .B(new_n5712_), .ZN(new_n5713_));
  NOR3_X1    g05457(.A1(new_n5539_), .A2(new_n5523_), .A3(new_n5711_), .ZN(new_n5714_));
  NOR3_X1    g05458(.A1(new_n5714_), .A2(new_n5707_), .A3(new_n5713_), .ZN(new_n5715_));
  INV_X1     g05459(.I(new_n5706_), .ZN(new_n5716_));
  NOR2_X1    g05460(.A1(new_n5716_), .A2(new_n5704_), .ZN(new_n5717_));
  OAI21_X1   g05461(.A1(new_n5539_), .A2(new_n5523_), .B(new_n5711_), .ZN(new_n5718_));
  NAND3_X1   g05462(.A1(new_n5528_), .A2(new_n5533_), .A3(new_n5712_), .ZN(new_n5719_));
  AOI21_X1   g05463(.A1(new_n5718_), .A2(new_n5719_), .B(new_n5717_), .ZN(new_n5720_));
  OR2_X2     g05464(.A1(new_n5715_), .A2(new_n5720_), .Z(new_n5721_));
  OAI22_X1   g05465(.A1(new_n713_), .A2(new_n3624_), .B1(new_n3592_), .B2(new_n717_), .ZN(new_n5722_));
  AOI21_X1   g05466(.A1(\b[28] ), .A2(new_n1126_), .B(new_n5722_), .ZN(new_n5723_));
  OAI21_X1   g05467(.A1(new_n3634_), .A2(new_n986_), .B(new_n5723_), .ZN(new_n5724_));
  XOR2_X1    g05468(.A1(new_n5724_), .A2(\a[11] ), .Z(new_n5725_));
  INV_X1     g05469(.I(new_n5725_), .ZN(new_n5726_));
  AOI21_X1   g05470(.A1(new_n5554_), .A2(new_n5537_), .B(new_n5726_), .ZN(new_n5727_));
  NOR3_X1    g05471(.A1(new_n5543_), .A2(new_n5545_), .A3(new_n5725_), .ZN(new_n5728_));
  NOR3_X1    g05472(.A1(new_n5727_), .A2(new_n5728_), .A3(new_n5721_), .ZN(new_n5729_));
  NOR2_X1    g05473(.A1(new_n5715_), .A2(new_n5720_), .ZN(new_n5730_));
  OAI21_X1   g05474(.A1(new_n5543_), .A2(new_n5545_), .B(new_n5725_), .ZN(new_n5731_));
  NAND3_X1   g05475(.A1(new_n5554_), .A2(new_n5537_), .A3(new_n5726_), .ZN(new_n5732_));
  AOI21_X1   g05476(.A1(new_n5732_), .A2(new_n5731_), .B(new_n5730_), .ZN(new_n5733_));
  OR2_X2     g05477(.A1(new_n5729_), .A2(new_n5733_), .Z(new_n5734_));
  AOI22_X1   g05478(.A1(new_n518_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n636_), .ZN(new_n5735_));
  OAI21_X1   g05479(.A1(new_n4022_), .A2(new_n917_), .B(new_n5735_), .ZN(new_n5736_));
  AOI21_X1   g05480(.A1(new_n4223_), .A2(new_n618_), .B(new_n5736_), .ZN(new_n5737_));
  XOR2_X1    g05481(.A1(new_n5737_), .A2(new_n488_), .Z(new_n5738_));
  INV_X1     g05482(.I(new_n5738_), .ZN(new_n5739_));
  AOI21_X1   g05483(.A1(new_n5558_), .A2(new_n5560_), .B(new_n5739_), .ZN(new_n5740_));
  OAI21_X1   g05484(.A1(new_n5559_), .A2(new_n5562_), .B(new_n5560_), .ZN(new_n5741_));
  NOR2_X1    g05485(.A1(new_n5741_), .A2(new_n5738_), .ZN(new_n5742_));
  NOR3_X1    g05486(.A1(new_n5742_), .A2(new_n5734_), .A3(new_n5740_), .ZN(new_n5743_));
  INV_X1     g05487(.I(new_n5743_), .ZN(new_n5744_));
  OAI21_X1   g05488(.A1(new_n5742_), .A2(new_n5740_), .B(new_n5734_), .ZN(new_n5745_));
  AOI21_X1   g05489(.A1(new_n5744_), .A2(new_n5745_), .B(new_n5598_), .ZN(new_n5746_));
  INV_X1     g05490(.I(new_n5746_), .ZN(new_n5747_));
  INV_X1     g05491(.I(new_n5598_), .ZN(new_n5748_));
  NOR2_X1    g05492(.A1(new_n5729_), .A2(new_n5733_), .ZN(new_n5749_));
  INV_X1     g05493(.I(new_n5740_), .ZN(new_n5750_));
  NAND3_X1   g05494(.A1(new_n5558_), .A2(new_n5560_), .A3(new_n5739_), .ZN(new_n5751_));
  AOI21_X1   g05495(.A1(new_n5750_), .A2(new_n5751_), .B(new_n5749_), .ZN(new_n5752_));
  NOR3_X1    g05496(.A1(new_n5752_), .A2(new_n5748_), .A3(new_n5743_), .ZN(new_n5753_));
  INV_X1     g05497(.I(new_n5753_), .ZN(new_n5754_));
  NAND2_X1   g05498(.A1(new_n283_), .A2(\b[37] ), .ZN(new_n5755_));
  AOI22_X1   g05499(.A1(new_n267_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n261_), .ZN(new_n5756_));
  NOR3_X1    g05500(.A1(new_n5346_), .A2(\b[37] ), .A3(new_n5341_), .ZN(new_n5757_));
  NAND3_X1   g05501(.A1(new_n5346_), .A2(\b[37] ), .A3(new_n5341_), .ZN(new_n5758_));
  INV_X1     g05502(.I(new_n5758_), .ZN(new_n5759_));
  OAI21_X1   g05503(.A1(new_n5759_), .A2(new_n5757_), .B(\b[39] ), .ZN(new_n5760_));
  INV_X1     g05504(.I(\b[39] ), .ZN(new_n5761_));
  INV_X1     g05505(.I(new_n5757_), .ZN(new_n5762_));
  NAND3_X1   g05506(.A1(new_n5762_), .A2(new_n5761_), .A3(new_n5758_), .ZN(new_n5763_));
  NAND3_X1   g05507(.A1(new_n5763_), .A2(new_n5760_), .A3(new_n265_), .ZN(new_n5764_));
  NAND3_X1   g05508(.A1(new_n5764_), .A2(new_n5755_), .A3(new_n5756_), .ZN(new_n5765_));
  XOR2_X1    g05509(.A1(new_n5765_), .A2(\a[2] ), .Z(new_n5766_));
  AOI21_X1   g05510(.A1(new_n5747_), .A2(new_n5754_), .B(new_n5766_), .ZN(new_n5767_));
  XOR2_X1    g05511(.A1(new_n5765_), .A2(new_n270_), .Z(new_n5768_));
  NOR3_X1    g05512(.A1(new_n5768_), .A2(new_n5746_), .A3(new_n5753_), .ZN(new_n5769_));
  NOR3_X1    g05513(.A1(new_n5767_), .A2(new_n5769_), .A3(new_n5593_), .ZN(new_n5770_));
  OAI21_X1   g05514(.A1(new_n5583_), .A2(new_n5577_), .B(new_n5585_), .ZN(new_n5771_));
  OAI21_X1   g05515(.A1(new_n5746_), .A2(new_n5753_), .B(new_n5768_), .ZN(new_n5772_));
  NAND3_X1   g05516(.A1(new_n5766_), .A2(new_n5747_), .A3(new_n5754_), .ZN(new_n5773_));
  AOI21_X1   g05517(.A1(new_n5772_), .A2(new_n5773_), .B(new_n5771_), .ZN(new_n5774_));
  NOR2_X1    g05518(.A1(new_n5770_), .A2(new_n5774_), .ZN(new_n5775_));
  OAI21_X1   g05519(.A1(new_n5340_), .A2(new_n5588_), .B(new_n5590_), .ZN(new_n5776_));
  XOR2_X1    g05520(.A1(new_n5776_), .A2(new_n5775_), .Z(\f[39] ));
  OAI21_X1   g05521(.A1(new_n5746_), .A2(new_n5753_), .B(new_n5771_), .ZN(new_n5778_));
  NAND3_X1   g05522(.A1(new_n5747_), .A2(new_n5593_), .A3(new_n5754_), .ZN(new_n5779_));
  AOI21_X1   g05523(.A1(new_n5779_), .A2(new_n5778_), .B(new_n5768_), .ZN(new_n5780_));
  AOI21_X1   g05524(.A1(new_n5776_), .A2(new_n5775_), .B(new_n5780_), .ZN(new_n5781_));
  AOI22_X1   g05525(.A1(new_n267_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n261_), .ZN(new_n5782_));
  OAI21_X1   g05526(.A1(new_n5341_), .A2(new_n284_), .B(new_n5782_), .ZN(new_n5783_));
  XOR2_X1    g05527(.A1(\b[39] ), .A2(\b[40] ), .Z(new_n5784_));
  NAND2_X1   g05528(.A1(new_n5346_), .A2(\b[37] ), .ZN(new_n5785_));
  AOI21_X1   g05529(.A1(new_n5785_), .A2(new_n5341_), .B(new_n5761_), .ZN(new_n5786_));
  INV_X1     g05530(.I(new_n5346_), .ZN(new_n5787_));
  AOI21_X1   g05531(.A1(new_n5787_), .A2(new_n5312_), .B(new_n5341_), .ZN(new_n5788_));
  NOR2_X1    g05532(.A1(new_n5786_), .A2(new_n5788_), .ZN(new_n5789_));
  NOR2_X1    g05533(.A1(new_n5789_), .A2(new_n5784_), .ZN(new_n5790_));
  INV_X1     g05534(.I(new_n5790_), .ZN(new_n5791_));
  NAND2_X1   g05535(.A1(new_n5789_), .A2(new_n5784_), .ZN(new_n5792_));
  NAND2_X1   g05536(.A1(new_n5791_), .A2(new_n5792_), .ZN(new_n5793_));
  AOI21_X1   g05537(.A1(new_n5793_), .A2(new_n265_), .B(new_n5783_), .ZN(new_n5794_));
  XOR2_X1    g05538(.A1(new_n5794_), .A2(\a[2] ), .Z(new_n5795_));
  OAI21_X1   g05539(.A1(new_n5752_), .A2(new_n5743_), .B(new_n5598_), .ZN(new_n5796_));
  NOR3_X1    g05540(.A1(new_n5752_), .A2(new_n5598_), .A3(new_n5743_), .ZN(new_n5797_));
  OAI21_X1   g05541(.A1(new_n5771_), .A2(new_n5797_), .B(new_n5796_), .ZN(new_n5798_));
  AOI22_X1   g05542(.A1(new_n800_), .A2(\b[36] ), .B1(\b[37] ), .B2(new_n333_), .ZN(new_n5799_));
  OAI21_X1   g05543(.A1(new_n4666_), .A2(new_n392_), .B(new_n5799_), .ZN(new_n5800_));
  INV_X1     g05544(.I(new_n5800_), .ZN(new_n5801_));
  OAI21_X1   g05545(.A1(new_n5322_), .A2(new_n318_), .B(new_n5801_), .ZN(new_n5802_));
  XOR2_X1    g05546(.A1(new_n5802_), .A2(new_n312_), .Z(new_n5803_));
  AOI21_X1   g05547(.A1(new_n5300_), .A2(new_n5293_), .B(new_n5302_), .ZN(new_n5804_));
  AOI21_X1   g05548(.A1(new_n5804_), .A2(new_n5557_), .B(new_n5549_), .ZN(new_n5805_));
  OAI21_X1   g05549(.A1(new_n5805_), .A2(new_n5739_), .B(new_n5749_), .ZN(new_n5806_));
  OAI21_X1   g05550(.A1(new_n5721_), .A2(new_n5727_), .B(new_n5732_), .ZN(new_n5807_));
  OAI21_X1   g05551(.A1(new_n5707_), .A2(new_n5713_), .B(new_n5719_), .ZN(new_n5808_));
  OAI22_X1   g05552(.A1(new_n993_), .A2(new_n3185_), .B1(new_n3158_), .B2(new_n997_), .ZN(new_n5809_));
  AOI21_X1   g05553(.A1(\b[26] ), .A2(new_n1486_), .B(new_n5809_), .ZN(new_n5810_));
  OAI21_X1   g05554(.A1(new_n3196_), .A2(new_n1323_), .B(new_n5810_), .ZN(new_n5811_));
  XOR2_X1    g05555(.A1(new_n5811_), .A2(\a[14] ), .Z(new_n5812_));
  AOI21_X1   g05556(.A1(new_n5518_), .A2(new_n5521_), .B(new_n5519_), .ZN(new_n5813_));
  NAND2_X1   g05557(.A1(new_n5813_), .A2(new_n5701_), .ZN(new_n5814_));
  NOR3_X1    g05558(.A1(new_n5694_), .A2(new_n5693_), .A3(new_n5692_), .ZN(new_n5815_));
  AOI21_X1   g05559(.A1(new_n5686_), .A2(new_n5689_), .B(new_n5679_), .ZN(new_n5816_));
  NOR2_X1    g05560(.A1(new_n5816_), .A2(new_n5815_), .ZN(new_n5817_));
  OAI21_X1   g05561(.A1(new_n5813_), .A2(new_n5701_), .B(new_n5817_), .ZN(new_n5818_));
  OAI22_X1   g05562(.A1(new_n1592_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n1505_), .ZN(new_n5819_));
  AOI21_X1   g05563(.A1(\b[23] ), .A2(new_n1584_), .B(new_n5819_), .ZN(new_n5820_));
  OAI21_X1   g05564(.A1(new_n2655_), .A2(new_n1732_), .B(new_n5820_), .ZN(new_n5821_));
  XOR2_X1    g05565(.A1(new_n5821_), .A2(\a[17] ), .Z(new_n5822_));
  AOI21_X1   g05566(.A1(new_n5685_), .A2(new_n5683_), .B(new_n5692_), .ZN(new_n5823_));
  AOI22_X1   g05567(.A1(new_n1738_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n1743_), .ZN(new_n5824_));
  OAI21_X1   g05568(.A1(new_n1860_), .A2(new_n1931_), .B(new_n5824_), .ZN(new_n5825_));
  AOI21_X1   g05569(.A1(new_n2659_), .A2(new_n1746_), .B(new_n5825_), .ZN(new_n5826_));
  XOR2_X1    g05570(.A1(new_n5826_), .A2(new_n1736_), .Z(new_n5827_));
  OAI21_X1   g05571(.A1(new_n5674_), .A2(new_n5673_), .B(new_n5667_), .ZN(new_n5828_));
  AOI22_X1   g05572(.A1(new_n2202_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n2205_), .ZN(new_n5829_));
  OAI21_X1   g05573(.A1(new_n1432_), .A2(new_n2370_), .B(new_n5829_), .ZN(new_n5830_));
  AOI21_X1   g05574(.A1(new_n1695_), .A2(new_n2208_), .B(new_n5830_), .ZN(new_n5831_));
  XOR2_X1    g05575(.A1(new_n5831_), .A2(new_n2200_), .Z(new_n5832_));
  AOI21_X1   g05576(.A1(new_n4968_), .A2(new_n4978_), .B(new_n4976_), .ZN(new_n5833_));
  OAI21_X1   g05577(.A1(new_n5833_), .A2(new_n5226_), .B(new_n5222_), .ZN(new_n5834_));
  OAI21_X1   g05578(.A1(new_n5834_), .A2(new_n5481_), .B(new_n5474_), .ZN(new_n5835_));
  NOR2_X1    g05579(.A1(new_n5835_), .A2(new_n5660_), .ZN(new_n5836_));
  INV_X1     g05580(.I(new_n5654_), .ZN(new_n5837_));
  NAND2_X1   g05581(.A1(new_n5462_), .A2(new_n5465_), .ZN(new_n5838_));
  AOI21_X1   g05582(.A1(new_n5838_), .A2(new_n5651_), .B(new_n5646_), .ZN(new_n5839_));
  AOI21_X1   g05583(.A1(new_n5636_), .A2(new_n5631_), .B(new_n5627_), .ZN(new_n5840_));
  OAI21_X1   g05584(.A1(new_n5620_), .A2(new_n5619_), .B(new_n5612_), .ZN(new_n5841_));
  NAND2_X1   g05585(.A1(new_n5841_), .A2(new_n5621_), .ZN(new_n5842_));
  AOI22_X1   g05586(.A1(new_n5155_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n5160_), .ZN(new_n5843_));
  NAND2_X1   g05587(.A1(new_n5420_), .A2(\b[2] ), .ZN(new_n5844_));
  NAND2_X1   g05588(.A1(new_n1725_), .A2(new_n5166_), .ZN(new_n5845_));
  NAND3_X1   g05589(.A1(new_n5845_), .A2(new_n5843_), .A3(new_n5844_), .ZN(new_n5846_));
  XOR2_X1    g05590(.A1(new_n5846_), .A2(\a[38] ), .Z(new_n5847_));
  INV_X1     g05591(.I(new_n5847_), .ZN(new_n5848_));
  INV_X1     g05592(.I(\a[41] ), .ZN(new_n5849_));
  XOR2_X1    g05593(.A1(\a[38] ), .A2(\a[39] ), .Z(new_n5850_));
  XNOR2_X1   g05594(.A1(\a[40] ), .A2(\a[41] ), .ZN(new_n5851_));
  NAND2_X1   g05595(.A1(new_n5851_), .A2(new_n5850_), .ZN(new_n5852_));
  INV_X1     g05596(.I(\a[40] ), .ZN(new_n5853_));
  NOR3_X1    g05597(.A1(new_n5853_), .A2(\a[38] ), .A3(\a[39] ), .ZN(new_n5854_));
  INV_X1     g05598(.I(\a[39] ), .ZN(new_n5855_));
  NOR3_X1    g05599(.A1(new_n5162_), .A2(new_n5855_), .A3(\a[40] ), .ZN(new_n5856_));
  NOR2_X1    g05600(.A1(new_n5856_), .A2(new_n5854_), .ZN(new_n5857_));
  OAI22_X1   g05601(.A1(new_n5852_), .A2(new_n275_), .B1(new_n258_), .B2(new_n5857_), .ZN(new_n5858_));
  NOR2_X1    g05602(.A1(new_n5849_), .A2(\a[40] ), .ZN(new_n5859_));
  NOR2_X1    g05603(.A1(new_n5853_), .A2(\a[41] ), .ZN(new_n5860_));
  OAI21_X1   g05604(.A1(new_n5859_), .A2(new_n5860_), .B(new_n5850_), .ZN(new_n5861_));
  NOR2_X1    g05605(.A1(new_n5861_), .A2(new_n313_), .ZN(new_n5862_));
  NOR2_X1    g05606(.A1(new_n5858_), .A2(new_n5862_), .ZN(new_n5863_));
  NOR2_X1    g05607(.A1(new_n5863_), .A2(new_n5849_), .ZN(new_n5864_));
  INV_X1     g05608(.I(new_n5864_), .ZN(new_n5865_));
  NAND2_X1   g05609(.A1(new_n5863_), .A2(new_n5849_), .ZN(new_n5866_));
  NOR2_X1    g05610(.A1(new_n5606_), .A2(new_n5849_), .ZN(new_n5867_));
  INV_X1     g05611(.I(new_n5867_), .ZN(new_n5868_));
  NAND3_X1   g05612(.A1(new_n5865_), .A2(new_n5866_), .A3(new_n5868_), .ZN(new_n5869_));
  NAND2_X1   g05613(.A1(new_n5864_), .A2(new_n5607_), .ZN(new_n5870_));
  AOI21_X1   g05614(.A1(new_n5869_), .A2(new_n5870_), .B(new_n5848_), .ZN(new_n5871_));
  NAND2_X1   g05615(.A1(new_n5869_), .A2(new_n5870_), .ZN(new_n5872_));
  NOR2_X1    g05616(.A1(new_n5872_), .A2(new_n5847_), .ZN(new_n5873_));
  NOR2_X1    g05617(.A1(new_n5871_), .A2(new_n5873_), .ZN(new_n5874_));
  NOR2_X1    g05618(.A1(new_n5604_), .A2(new_n5607_), .ZN(new_n5875_));
  OAI21_X1   g05619(.A1(new_n5599_), .A2(new_n5875_), .B(new_n5608_), .ZN(new_n5876_));
  NOR2_X1    g05620(.A1(new_n5874_), .A2(new_n5876_), .ZN(new_n5877_));
  NAND2_X1   g05621(.A1(new_n5872_), .A2(new_n5847_), .ZN(new_n5878_));
  NAND3_X1   g05622(.A1(new_n5848_), .A2(new_n5869_), .A3(new_n5870_), .ZN(new_n5879_));
  NAND2_X1   g05623(.A1(new_n5878_), .A2(new_n5879_), .ZN(new_n5880_));
  NOR2_X1    g05624(.A1(new_n5609_), .A2(new_n5606_), .ZN(new_n5881_));
  AOI21_X1   g05625(.A1(new_n5427_), .A2(new_n5610_), .B(new_n5881_), .ZN(new_n5882_));
  NOR2_X1    g05626(.A1(new_n5880_), .A2(new_n5882_), .ZN(new_n5883_));
  OAI22_X1   g05627(.A1(new_n471_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n438_), .ZN(new_n5884_));
  AOI21_X1   g05628(.A1(\b[5] ), .A2(new_n4706_), .B(new_n5884_), .ZN(new_n5885_));
  OAI21_X1   g05629(.A1(new_n485_), .A2(new_n4458_), .B(new_n5885_), .ZN(new_n5886_));
  XOR2_X1    g05630(.A1(new_n5886_), .A2(\a[35] ), .Z(new_n5887_));
  NOR3_X1    g05631(.A1(new_n5877_), .A2(new_n5883_), .A3(new_n5887_), .ZN(new_n5888_));
  NAND2_X1   g05632(.A1(new_n5880_), .A2(new_n5882_), .ZN(new_n5889_));
  NAND2_X1   g05633(.A1(new_n5874_), .A2(new_n5876_), .ZN(new_n5890_));
  INV_X1     g05634(.I(new_n5887_), .ZN(new_n5891_));
  AOI21_X1   g05635(.A1(new_n5890_), .A2(new_n5889_), .B(new_n5891_), .ZN(new_n5892_));
  NOR2_X1    g05636(.A1(new_n5892_), .A2(new_n5888_), .ZN(new_n5893_));
  NAND2_X1   g05637(.A1(new_n5842_), .A2(new_n5893_), .ZN(new_n5894_));
  NAND3_X1   g05638(.A1(new_n5890_), .A2(new_n5889_), .A3(new_n5891_), .ZN(new_n5895_));
  OAI21_X1   g05639(.A1(new_n5877_), .A2(new_n5883_), .B(new_n5887_), .ZN(new_n5896_));
  NAND2_X1   g05640(.A1(new_n5895_), .A2(new_n5896_), .ZN(new_n5897_));
  NAND3_X1   g05641(.A1(new_n5897_), .A2(new_n5621_), .A3(new_n5841_), .ZN(new_n5898_));
  AOI22_X1   g05642(.A1(new_n3864_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n3869_), .ZN(new_n5899_));
  OAI21_X1   g05643(.A1(new_n577_), .A2(new_n5410_), .B(new_n5899_), .ZN(new_n5900_));
  AOI21_X1   g05644(.A1(new_n1059_), .A2(new_n3872_), .B(new_n5900_), .ZN(new_n5901_));
  XOR2_X1    g05645(.A1(new_n5901_), .A2(new_n3876_), .Z(new_n5902_));
  INV_X1     g05646(.I(new_n5902_), .ZN(new_n5903_));
  NAND3_X1   g05647(.A1(new_n5894_), .A2(new_n5898_), .A3(new_n5903_), .ZN(new_n5904_));
  INV_X1     g05648(.I(new_n5904_), .ZN(new_n5905_));
  AOI21_X1   g05649(.A1(new_n5894_), .A2(new_n5898_), .B(new_n5903_), .ZN(new_n5906_));
  OAI22_X1   g05650(.A1(new_n5905_), .A2(new_n5906_), .B1(new_n5840_), .B2(new_n5637_), .ZN(new_n5907_));
  OAI21_X1   g05651(.A1(new_n5634_), .A2(new_n5632_), .B(new_n5641_), .ZN(new_n5908_));
  INV_X1     g05652(.I(new_n5906_), .ZN(new_n5909_));
  NAND4_X1   g05653(.A1(new_n5909_), .A2(new_n5643_), .A3(new_n5908_), .A4(new_n5904_), .ZN(new_n5910_));
  OAI22_X1   g05654(.A1(new_n1070_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n941_), .ZN(new_n5911_));
  AOI21_X1   g05655(.A1(\b[11] ), .A2(new_n3456_), .B(new_n5911_), .ZN(new_n5912_));
  OAI21_X1   g05656(.A1(new_n1082_), .A2(new_n3261_), .B(new_n5912_), .ZN(new_n5913_));
  XOR2_X1    g05657(.A1(new_n5913_), .A2(\a[29] ), .Z(new_n5914_));
  AOI21_X1   g05658(.A1(new_n5907_), .A2(new_n5910_), .B(new_n5914_), .ZN(new_n5915_));
  AOI22_X1   g05659(.A1(new_n5909_), .A2(new_n5904_), .B1(new_n5908_), .B2(new_n5643_), .ZN(new_n5916_));
  NOR4_X1    g05660(.A1(new_n5905_), .A2(new_n5840_), .A3(new_n5637_), .A4(new_n5906_), .ZN(new_n5917_));
  XOR2_X1    g05661(.A1(new_n5913_), .A2(new_n3264_), .Z(new_n5918_));
  NOR3_X1    g05662(.A1(new_n5916_), .A2(new_n5917_), .A3(new_n5918_), .ZN(new_n5919_));
  NOR2_X1    g05663(.A1(new_n5919_), .A2(new_n5915_), .ZN(new_n5920_));
  OAI21_X1   g05664(.A1(new_n5839_), .A2(new_n5837_), .B(new_n5920_), .ZN(new_n5921_));
  NAND2_X1   g05665(.A1(new_n5652_), .A2(new_n5645_), .ZN(new_n5922_));
  OAI21_X1   g05666(.A1(new_n5916_), .A2(new_n5917_), .B(new_n5918_), .ZN(new_n5923_));
  NAND3_X1   g05667(.A1(new_n5907_), .A2(new_n5910_), .A3(new_n5914_), .ZN(new_n5924_));
  NAND2_X1   g05668(.A1(new_n5923_), .A2(new_n5924_), .ZN(new_n5925_));
  NAND3_X1   g05669(.A1(new_n5922_), .A2(new_n5654_), .A3(new_n5925_), .ZN(new_n5926_));
  AOI22_X1   g05670(.A1(new_n2716_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n2719_), .ZN(new_n5927_));
  OAI21_X1   g05671(.A1(new_n1093_), .A2(new_n2924_), .B(new_n5927_), .ZN(new_n5928_));
  AOI21_X1   g05672(.A1(new_n1701_), .A2(new_n2722_), .B(new_n5928_), .ZN(new_n5929_));
  XOR2_X1    g05673(.A1(new_n5929_), .A2(new_n2714_), .Z(new_n5930_));
  INV_X1     g05674(.I(new_n5930_), .ZN(new_n5931_));
  NAND3_X1   g05675(.A1(new_n5926_), .A2(new_n5921_), .A3(new_n5931_), .ZN(new_n5932_));
  AOI21_X1   g05676(.A1(new_n5922_), .A2(new_n5654_), .B(new_n5925_), .ZN(new_n5933_));
  NOR3_X1    g05677(.A1(new_n5839_), .A2(new_n5837_), .A3(new_n5920_), .ZN(new_n5934_));
  OAI21_X1   g05678(.A1(new_n5933_), .A2(new_n5934_), .B(new_n5930_), .ZN(new_n5935_));
  NAND2_X1   g05679(.A1(new_n5935_), .A2(new_n5932_), .ZN(new_n5936_));
  XOR2_X1    g05680(.A1(new_n5655_), .A2(new_n5645_), .Z(new_n5937_));
  AOI21_X1   g05681(.A1(new_n5835_), .A2(new_n5660_), .B(new_n5937_), .ZN(new_n5938_));
  NOR3_X1    g05682(.A1(new_n5938_), .A2(new_n5836_), .A3(new_n5936_), .ZN(new_n5939_));
  NOR3_X1    g05683(.A1(new_n5933_), .A2(new_n5934_), .A3(new_n5930_), .ZN(new_n5940_));
  AOI21_X1   g05684(.A1(new_n5926_), .A2(new_n5921_), .B(new_n5931_), .ZN(new_n5941_));
  NOR2_X1    g05685(.A1(new_n5941_), .A2(new_n5940_), .ZN(new_n5942_));
  AOI21_X1   g05686(.A1(new_n5486_), .A2(new_n5477_), .B(new_n5475_), .ZN(new_n5943_));
  OAI21_X1   g05687(.A1(new_n5943_), .A2(new_n5662_), .B(new_n5656_), .ZN(new_n5944_));
  AOI21_X1   g05688(.A1(new_n5944_), .A2(new_n5663_), .B(new_n5942_), .ZN(new_n5945_));
  OAI21_X1   g05689(.A1(new_n5939_), .A2(new_n5945_), .B(new_n5832_), .ZN(new_n5946_));
  INV_X1     g05690(.I(new_n5832_), .ZN(new_n5947_));
  NAND3_X1   g05691(.A1(new_n5944_), .A2(new_n5663_), .A3(new_n5942_), .ZN(new_n5948_));
  OAI21_X1   g05692(.A1(new_n5938_), .A2(new_n5836_), .B(new_n5936_), .ZN(new_n5949_));
  NAND3_X1   g05693(.A1(new_n5949_), .A2(new_n5948_), .A3(new_n5947_), .ZN(new_n5950_));
  NAND2_X1   g05694(.A1(new_n5946_), .A2(new_n5950_), .ZN(new_n5951_));
  NAND3_X1   g05695(.A1(new_n5828_), .A2(new_n5951_), .A3(new_n5675_), .ZN(new_n5952_));
  NOR3_X1    g05696(.A1(new_n5500_), .A2(new_n5488_), .A3(new_n5671_), .ZN(new_n5953_));
  INV_X1     g05697(.I(new_n5666_), .ZN(new_n5954_));
  NAND2_X1   g05698(.A1(new_n5954_), .A2(new_n5664_), .ZN(new_n5955_));
  AOI21_X1   g05699(.A1(new_n5236_), .A2(new_n5239_), .B(new_n5490_), .ZN(new_n5956_));
  OAI21_X1   g05700(.A1(new_n5956_), .A2(new_n5496_), .B(new_n5495_), .ZN(new_n5957_));
  AOI21_X1   g05701(.A1(new_n5957_), .A2(new_n5671_), .B(new_n5955_), .ZN(new_n5958_));
  AOI21_X1   g05702(.A1(new_n5949_), .A2(new_n5948_), .B(new_n5947_), .ZN(new_n5959_));
  NOR3_X1    g05703(.A1(new_n5939_), .A2(new_n5945_), .A3(new_n5832_), .ZN(new_n5960_));
  NOR2_X1    g05704(.A1(new_n5960_), .A2(new_n5959_), .ZN(new_n5961_));
  OAI21_X1   g05705(.A1(new_n5958_), .A2(new_n5953_), .B(new_n5961_), .ZN(new_n5962_));
  NAND3_X1   g05706(.A1(new_n5962_), .A2(new_n5952_), .A3(new_n5827_), .ZN(new_n5963_));
  INV_X1     g05707(.I(new_n5827_), .ZN(new_n5964_));
  NOR3_X1    g05708(.A1(new_n5958_), .A2(new_n5961_), .A3(new_n5953_), .ZN(new_n5965_));
  AOI21_X1   g05709(.A1(new_n5828_), .A2(new_n5675_), .B(new_n5951_), .ZN(new_n5966_));
  OAI21_X1   g05710(.A1(new_n5965_), .A2(new_n5966_), .B(new_n5964_), .ZN(new_n5967_));
  NAND2_X1   g05711(.A1(new_n5967_), .A2(new_n5963_), .ZN(new_n5968_));
  NOR3_X1    g05712(.A1(new_n5823_), .A2(new_n5694_), .A3(new_n5968_), .ZN(new_n5969_));
  OAI21_X1   g05713(.A1(new_n5688_), .A2(new_n5687_), .B(new_n5679_), .ZN(new_n5970_));
  NOR3_X1    g05714(.A1(new_n5965_), .A2(new_n5966_), .A3(new_n5964_), .ZN(new_n5971_));
  AOI21_X1   g05715(.A1(new_n5962_), .A2(new_n5952_), .B(new_n5827_), .ZN(new_n5972_));
  NOR2_X1    g05716(.A1(new_n5971_), .A2(new_n5972_), .ZN(new_n5973_));
  AOI21_X1   g05717(.A1(new_n5970_), .A2(new_n5689_), .B(new_n5973_), .ZN(new_n5974_));
  OAI21_X1   g05718(.A1(new_n5969_), .A2(new_n5974_), .B(new_n5822_), .ZN(new_n5975_));
  INV_X1     g05719(.I(new_n5822_), .ZN(new_n5976_));
  NAND3_X1   g05720(.A1(new_n5970_), .A2(new_n5973_), .A3(new_n5689_), .ZN(new_n5977_));
  OAI21_X1   g05721(.A1(new_n5823_), .A2(new_n5694_), .B(new_n5968_), .ZN(new_n5978_));
  NAND3_X1   g05722(.A1(new_n5978_), .A2(new_n5977_), .A3(new_n5976_), .ZN(new_n5979_));
  NAND2_X1   g05723(.A1(new_n5975_), .A2(new_n5979_), .ZN(new_n5980_));
  NAND3_X1   g05724(.A1(new_n5818_), .A2(new_n5814_), .A3(new_n5980_), .ZN(new_n5981_));
  AOI21_X1   g05725(.A1(new_n5260_), .A2(new_n5263_), .B(new_n5388_), .ZN(new_n5982_));
  OAI21_X1   g05726(.A1(new_n5982_), .A2(new_n5515_), .B(new_n5510_), .ZN(new_n5983_));
  AOI21_X1   g05727(.A1(new_n5983_), .A2(new_n5700_), .B(new_n5696_), .ZN(new_n5984_));
  AOI21_X1   g05728(.A1(new_n5978_), .A2(new_n5977_), .B(new_n5976_), .ZN(new_n5985_));
  NOR3_X1    g05729(.A1(new_n5969_), .A2(new_n5974_), .A3(new_n5822_), .ZN(new_n5986_));
  NOR2_X1    g05730(.A1(new_n5986_), .A2(new_n5985_), .ZN(new_n5987_));
  OAI21_X1   g05731(.A1(new_n5984_), .A2(new_n5703_), .B(new_n5987_), .ZN(new_n5988_));
  NAND3_X1   g05732(.A1(new_n5988_), .A2(new_n5981_), .A3(new_n5812_), .ZN(new_n5989_));
  INV_X1     g05733(.I(new_n5812_), .ZN(new_n5990_));
  NOR3_X1    g05734(.A1(new_n5984_), .A2(new_n5703_), .A3(new_n5987_), .ZN(new_n5991_));
  AOI21_X1   g05735(.A1(new_n5818_), .A2(new_n5814_), .B(new_n5980_), .ZN(new_n5992_));
  OAI21_X1   g05736(.A1(new_n5991_), .A2(new_n5992_), .B(new_n5990_), .ZN(new_n5993_));
  NAND2_X1   g05737(.A1(new_n5993_), .A2(new_n5989_), .ZN(new_n5994_));
  NAND2_X1   g05738(.A1(new_n5808_), .A2(new_n5994_), .ZN(new_n5995_));
  AOI21_X1   g05739(.A1(new_n5271_), .A2(new_n5272_), .B(new_n5266_), .ZN(new_n5996_));
  AOI21_X1   g05740(.A1(new_n5996_), .A2(new_n5527_), .B(new_n5523_), .ZN(new_n5997_));
  OAI21_X1   g05741(.A1(new_n5997_), .A2(new_n5712_), .B(new_n5717_), .ZN(new_n5998_));
  NOR3_X1    g05742(.A1(new_n5991_), .A2(new_n5992_), .A3(new_n5990_), .ZN(new_n5999_));
  AOI21_X1   g05743(.A1(new_n5988_), .A2(new_n5981_), .B(new_n5812_), .ZN(new_n6000_));
  NOR2_X1    g05744(.A1(new_n5999_), .A2(new_n6000_), .ZN(new_n6001_));
  NAND3_X1   g05745(.A1(new_n5998_), .A2(new_n5719_), .A3(new_n6001_), .ZN(new_n6002_));
  NAND2_X1   g05746(.A1(new_n4619_), .A2(new_n4616_), .ZN(new_n6003_));
  OAI22_X1   g05747(.A1(new_n713_), .A2(new_n4022_), .B1(new_n3624_), .B2(new_n717_), .ZN(new_n6004_));
  AOI21_X1   g05748(.A1(\b[29] ), .A2(new_n1126_), .B(new_n6004_), .ZN(new_n6005_));
  OAI21_X1   g05749(.A1(new_n6003_), .A2(new_n986_), .B(new_n6005_), .ZN(new_n6006_));
  XOR2_X1    g05750(.A1(new_n6006_), .A2(\a[11] ), .Z(new_n6007_));
  AOI21_X1   g05751(.A1(new_n5995_), .A2(new_n6002_), .B(new_n6007_), .ZN(new_n6008_));
  NAND3_X1   g05752(.A1(new_n5995_), .A2(new_n6002_), .A3(new_n6007_), .ZN(new_n6009_));
  INV_X1     g05753(.I(new_n6009_), .ZN(new_n6010_));
  NOR2_X1    g05754(.A1(new_n6010_), .A2(new_n6008_), .ZN(new_n6011_));
  NAND2_X1   g05755(.A1(new_n5807_), .A2(new_n6011_), .ZN(new_n6012_));
  AOI21_X1   g05756(.A1(new_n5730_), .A2(new_n5731_), .B(new_n5728_), .ZN(new_n6013_));
  INV_X1     g05757(.I(new_n6008_), .ZN(new_n6014_));
  NAND2_X1   g05758(.A1(new_n6014_), .A2(new_n6009_), .ZN(new_n6015_));
  NAND2_X1   g05759(.A1(new_n6013_), .A2(new_n6015_), .ZN(new_n6016_));
  AOI22_X1   g05760(.A1(new_n518_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n636_), .ZN(new_n6017_));
  OAI21_X1   g05761(.A1(new_n4023_), .A2(new_n917_), .B(new_n6017_), .ZN(new_n6018_));
  AOI21_X1   g05762(.A1(new_n5103_), .A2(new_n618_), .B(new_n6018_), .ZN(new_n6019_));
  XOR2_X1    g05763(.A1(new_n6019_), .A2(\a[8] ), .Z(new_n6020_));
  NAND3_X1   g05764(.A1(new_n6012_), .A2(new_n6016_), .A3(new_n6020_), .ZN(new_n6021_));
  NOR2_X1    g05765(.A1(new_n6013_), .A2(new_n6015_), .ZN(new_n6022_));
  NOR2_X1    g05766(.A1(new_n5807_), .A2(new_n6011_), .ZN(new_n6023_));
  XOR2_X1    g05767(.A1(new_n6019_), .A2(new_n488_), .Z(new_n6024_));
  OAI21_X1   g05768(.A1(new_n6023_), .A2(new_n6022_), .B(new_n6024_), .ZN(new_n6025_));
  NAND2_X1   g05769(.A1(new_n6025_), .A2(new_n6021_), .ZN(new_n6026_));
  AOI21_X1   g05770(.A1(new_n5751_), .A2(new_n5806_), .B(new_n6026_), .ZN(new_n6027_));
  OAI21_X1   g05771(.A1(new_n5734_), .A2(new_n5740_), .B(new_n5751_), .ZN(new_n6028_));
  NOR3_X1    g05772(.A1(new_n6023_), .A2(new_n6022_), .A3(new_n6024_), .ZN(new_n6029_));
  AOI21_X1   g05773(.A1(new_n6012_), .A2(new_n6016_), .B(new_n6020_), .ZN(new_n6030_));
  NOR2_X1    g05774(.A1(new_n6030_), .A2(new_n6029_), .ZN(new_n6031_));
  NOR2_X1    g05775(.A1(new_n6028_), .A2(new_n6031_), .ZN(new_n6032_));
  NOR3_X1    g05776(.A1(new_n6032_), .A2(new_n6027_), .A3(new_n5803_), .ZN(new_n6033_));
  XOR2_X1    g05777(.A1(new_n5802_), .A2(\a[5] ), .Z(new_n6034_));
  NAND2_X1   g05778(.A1(new_n6028_), .A2(new_n6031_), .ZN(new_n6035_));
  NAND3_X1   g05779(.A1(new_n6026_), .A2(new_n5806_), .A3(new_n5751_), .ZN(new_n6036_));
  AOI21_X1   g05780(.A1(new_n6035_), .A2(new_n6036_), .B(new_n6034_), .ZN(new_n6037_));
  NOR2_X1    g05781(.A1(new_n6033_), .A2(new_n6037_), .ZN(new_n6038_));
  XOR2_X1    g05782(.A1(new_n5798_), .A2(new_n6038_), .Z(new_n6039_));
  NOR2_X1    g05783(.A1(new_n6039_), .A2(new_n5795_), .ZN(new_n6040_));
  INV_X1     g05784(.I(new_n6040_), .ZN(new_n6041_));
  NAND2_X1   g05785(.A1(new_n6039_), .A2(new_n5795_), .ZN(new_n6042_));
  NAND2_X1   g05786(.A1(new_n6041_), .A2(new_n6042_), .ZN(new_n6043_));
  XOR2_X1    g05787(.A1(new_n5781_), .A2(new_n6043_), .Z(\f[40] ));
  OAI21_X1   g05788(.A1(new_n5781_), .A2(new_n6043_), .B(new_n6041_), .ZN(new_n6045_));
  NAND3_X1   g05789(.A1(new_n6035_), .A2(new_n6034_), .A3(new_n6036_), .ZN(new_n6046_));
  OAI21_X1   g05790(.A1(new_n6032_), .A2(new_n6027_), .B(new_n5803_), .ZN(new_n6047_));
  NAND2_X1   g05791(.A1(new_n6047_), .A2(new_n6046_), .ZN(new_n6048_));
  AOI21_X1   g05792(.A1(new_n6035_), .A2(new_n6036_), .B(new_n5803_), .ZN(new_n6049_));
  AOI21_X1   g05793(.A1(new_n5798_), .A2(new_n6048_), .B(new_n6049_), .ZN(new_n6050_));
  AOI22_X1   g05794(.A1(new_n800_), .A2(\b[37] ), .B1(\b[38] ), .B2(new_n333_), .ZN(new_n6051_));
  OAI21_X1   g05795(.A1(new_n4886_), .A2(new_n392_), .B(new_n6051_), .ZN(new_n6052_));
  AOI21_X1   g05796(.A1(new_n5351_), .A2(new_n330_), .B(new_n6052_), .ZN(new_n6053_));
  XOR2_X1    g05797(.A1(new_n6053_), .A2(new_n312_), .Z(new_n6054_));
  AOI22_X1   g05798(.A1(new_n518_), .A2(\b[35] ), .B1(\b[34] ), .B2(new_n636_), .ZN(new_n6055_));
  OAI21_X1   g05799(.A1(new_n4638_), .A2(new_n917_), .B(new_n6055_), .ZN(new_n6056_));
  INV_X1     g05800(.I(new_n6056_), .ZN(new_n6057_));
  NAND3_X1   g05801(.A1(new_n4675_), .A2(new_n618_), .A3(new_n4673_), .ZN(new_n6058_));
  AOI21_X1   g05802(.A1(new_n6058_), .A2(new_n6057_), .B(new_n488_), .ZN(new_n6059_));
  INV_X1     g05803(.I(new_n4673_), .ZN(new_n6060_));
  NOR3_X1    g05804(.A1(new_n6060_), .A2(new_n624_), .A3(new_n4674_), .ZN(new_n6061_));
  NOR3_X1    g05805(.A1(new_n6061_), .A2(\a[8] ), .A3(new_n6056_), .ZN(new_n6062_));
  NOR2_X1    g05806(.A1(new_n6062_), .A2(new_n6059_), .ZN(new_n6063_));
  OAI21_X1   g05807(.A1(new_n5109_), .A2(new_n5286_), .B(new_n5280_), .ZN(new_n6064_));
  OAI21_X1   g05808(.A1(new_n6064_), .A2(new_n5542_), .B(new_n5537_), .ZN(new_n6065_));
  AOI21_X1   g05809(.A1(new_n6065_), .A2(new_n5725_), .B(new_n5721_), .ZN(new_n6066_));
  OAI21_X1   g05810(.A1(new_n6066_), .A2(new_n5728_), .B(new_n6009_), .ZN(new_n6067_));
  OAI22_X1   g05811(.A1(new_n713_), .A2(new_n4023_), .B1(new_n4022_), .B2(new_n717_), .ZN(new_n6068_));
  AOI21_X1   g05812(.A1(\b[30] ), .A2(new_n1126_), .B(new_n6068_), .ZN(new_n6069_));
  OAI21_X1   g05813(.A1(new_n4031_), .A2(new_n986_), .B(new_n6069_), .ZN(new_n6070_));
  XOR2_X1    g05814(.A1(new_n6070_), .A2(new_n722_), .Z(new_n6071_));
  NOR3_X1    g05815(.A1(new_n5969_), .A2(new_n5974_), .A3(new_n5976_), .ZN(new_n6072_));
  OAI22_X1   g05816(.A1(new_n1592_), .A2(new_n3006_), .B1(new_n2646_), .B2(new_n1505_), .ZN(new_n6073_));
  AOI21_X1   g05817(.A1(\b[24] ), .A2(new_n1584_), .B(new_n6073_), .ZN(new_n6074_));
  OAI21_X1   g05818(.A1(new_n3016_), .A2(new_n1732_), .B(new_n6074_), .ZN(new_n6075_));
  XOR2_X1    g05819(.A1(new_n6075_), .A2(\a[17] ), .Z(new_n6076_));
  AOI22_X1   g05820(.A1(new_n1738_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n1743_), .ZN(new_n6077_));
  OAI21_X1   g05821(.A1(new_n2027_), .A2(new_n1931_), .B(new_n6077_), .ZN(new_n6078_));
  AOI21_X1   g05822(.A1(new_n2470_), .A2(new_n1746_), .B(new_n6078_), .ZN(new_n6079_));
  XOR2_X1    g05823(.A1(new_n6079_), .A2(new_n1736_), .Z(new_n6080_));
  INV_X1     g05824(.I(new_n6080_), .ZN(new_n6081_));
  AOI22_X1   g05825(.A1(new_n2202_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n2205_), .ZN(new_n6082_));
  OAI21_X1   g05826(.A1(new_n1553_), .A2(new_n2370_), .B(new_n6082_), .ZN(new_n6083_));
  AOI21_X1   g05827(.A1(new_n2452_), .A2(new_n2208_), .B(new_n6083_), .ZN(new_n6084_));
  XOR2_X1    g05828(.A1(new_n6084_), .A2(new_n2200_), .Z(new_n6085_));
  INV_X1     g05829(.I(new_n6085_), .ZN(new_n6086_));
  OAI22_X1   g05830(.A1(new_n2703_), .A2(new_n1432_), .B1(new_n1296_), .B2(new_n2708_), .ZN(new_n6087_));
  AOI21_X1   g05831(.A1(\b[15] ), .A2(new_n2906_), .B(new_n6087_), .ZN(new_n6088_));
  OAI21_X1   g05832(.A1(new_n1444_), .A2(new_n2711_), .B(new_n6088_), .ZN(new_n6089_));
  XOR2_X1    g05833(.A1(new_n6089_), .A2(\a[26] ), .Z(new_n6090_));
  OAI21_X1   g05834(.A1(new_n5839_), .A2(new_n5837_), .B(new_n5924_), .ZN(new_n6091_));
  AOI22_X1   g05835(.A1(new_n3267_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n3270_), .ZN(new_n6092_));
  OAI21_X1   g05836(.A1(new_n941_), .A2(new_n3475_), .B(new_n6092_), .ZN(new_n6093_));
  AOI21_X1   g05837(.A1(new_n1449_), .A2(new_n3273_), .B(new_n6093_), .ZN(new_n6094_));
  XOR2_X1    g05838(.A1(new_n6094_), .A2(new_n3264_), .Z(new_n6095_));
  INV_X1     g05839(.I(new_n6095_), .ZN(new_n6096_));
  NOR2_X1    g05840(.A1(new_n5840_), .A2(new_n5637_), .ZN(new_n6097_));
  AOI21_X1   g05841(.A1(new_n6097_), .A2(new_n5904_), .B(new_n5906_), .ZN(new_n6098_));
  INV_X1     g05842(.I(new_n4706_), .ZN(new_n6099_));
  AOI22_X1   g05843(.A1(new_n4918_), .A2(\b[8] ), .B1(\b[7] ), .B2(new_n4921_), .ZN(new_n6100_));
  OAI21_X1   g05844(.A1(new_n438_), .A2(new_n6099_), .B(new_n6100_), .ZN(new_n6101_));
  AOI21_X1   g05845(.A1(new_n799_), .A2(new_n4699_), .B(new_n6101_), .ZN(new_n6102_));
  XOR2_X1    g05846(.A1(new_n6102_), .A2(new_n4446_), .Z(new_n6103_));
  NOR2_X1    g05847(.A1(new_n5859_), .A2(new_n5860_), .ZN(new_n6104_));
  NOR2_X1    g05848(.A1(new_n6104_), .A2(new_n5605_), .ZN(new_n6105_));
  NAND2_X1   g05849(.A1(new_n6105_), .A2(new_n554_), .ZN(new_n6106_));
  XOR2_X1    g05850(.A1(\a[40] ), .A2(\a[41] ), .Z(new_n6107_));
  NOR2_X1    g05851(.A1(new_n5605_), .A2(new_n6107_), .ZN(new_n6108_));
  NAND3_X1   g05852(.A1(new_n5162_), .A2(new_n5855_), .A3(\a[40] ), .ZN(new_n6109_));
  NAND3_X1   g05853(.A1(new_n5853_), .A2(\a[38] ), .A3(\a[39] ), .ZN(new_n6110_));
  NAND2_X1   g05854(.A1(new_n6109_), .A2(new_n6110_), .ZN(new_n6111_));
  AOI22_X1   g05855(.A1(new_n6108_), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n6111_), .ZN(new_n6112_));
  NOR2_X1    g05856(.A1(new_n5859_), .A2(\a[38] ), .ZN(new_n6113_));
  AOI21_X1   g05857(.A1(\a[40] ), .A2(new_n5849_), .B(new_n5162_), .ZN(new_n6114_));
  NOR3_X1    g05858(.A1(new_n6113_), .A2(new_n5850_), .A3(new_n6114_), .ZN(new_n6115_));
  NAND2_X1   g05859(.A1(new_n6115_), .A2(\b[0] ), .ZN(new_n6116_));
  NAND3_X1   g05860(.A1(new_n6112_), .A2(new_n6116_), .A3(new_n6106_), .ZN(new_n6117_));
  XOR2_X1    g05861(.A1(new_n6117_), .A2(new_n5849_), .Z(new_n6118_));
  NAND3_X1   g05862(.A1(new_n5863_), .A2(\a[41] ), .A3(new_n5607_), .ZN(new_n6119_));
  NAND2_X1   g05863(.A1(new_n6118_), .A2(new_n6119_), .ZN(new_n6120_));
  INV_X1     g05864(.I(new_n5863_), .ZN(new_n6121_));
  OR4_X2     g05865(.A1(new_n5849_), .A2(new_n6121_), .A3(new_n5606_), .A4(new_n6117_), .Z(new_n6122_));
  NAND2_X1   g05866(.A1(new_n6120_), .A2(new_n6122_), .ZN(new_n6123_));
  INV_X1     g05867(.I(new_n5166_), .ZN(new_n6124_));
  XNOR2_X1   g05868(.A1(\a[37] ), .A2(\a[38] ), .ZN(new_n6125_));
  NAND2_X1   g05869(.A1(new_n6125_), .A2(new_n5417_), .ZN(new_n6126_));
  NOR3_X1    g05870(.A1(new_n5158_), .A2(\a[35] ), .A3(\a[36] ), .ZN(new_n6127_));
  INV_X1     g05871(.I(new_n5159_), .ZN(new_n6128_));
  NOR2_X1    g05872(.A1(new_n6128_), .A2(new_n6127_), .ZN(new_n6129_));
  OAI22_X1   g05873(.A1(new_n377_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n339_), .ZN(new_n6130_));
  AOI21_X1   g05874(.A1(\b[3] ), .A2(new_n5420_), .B(new_n6130_), .ZN(new_n6131_));
  OAI21_X1   g05875(.A1(new_n566_), .A2(new_n6124_), .B(new_n6131_), .ZN(new_n6132_));
  XOR2_X1    g05876(.A1(new_n6132_), .A2(new_n5162_), .Z(new_n6133_));
  XOR2_X1    g05877(.A1(new_n6123_), .A2(new_n6133_), .Z(new_n6134_));
  OAI21_X1   g05878(.A1(new_n5876_), .A2(new_n5873_), .B(new_n5878_), .ZN(new_n6135_));
  NAND2_X1   g05879(.A1(new_n6134_), .A2(new_n6135_), .ZN(new_n6136_));
  NAND2_X1   g05880(.A1(new_n6123_), .A2(new_n6133_), .ZN(new_n6137_));
  XOR2_X1    g05881(.A1(new_n6132_), .A2(\a[38] ), .Z(new_n6138_));
  NAND3_X1   g05882(.A1(new_n6138_), .A2(new_n6120_), .A3(new_n6122_), .ZN(new_n6139_));
  NAND2_X1   g05883(.A1(new_n6137_), .A2(new_n6139_), .ZN(new_n6140_));
  AOI21_X1   g05884(.A1(new_n5882_), .A2(new_n5879_), .B(new_n5871_), .ZN(new_n6141_));
  NAND2_X1   g05885(.A1(new_n6140_), .A2(new_n6141_), .ZN(new_n6142_));
  AOI21_X1   g05886(.A1(new_n6136_), .A2(new_n6142_), .B(new_n6103_), .ZN(new_n6143_));
  INV_X1     g05887(.I(new_n6103_), .ZN(new_n6144_));
  NOR2_X1    g05888(.A1(new_n6140_), .A2(new_n6141_), .ZN(new_n6145_));
  NOR2_X1    g05889(.A1(new_n6134_), .A2(new_n6135_), .ZN(new_n6146_));
  NOR3_X1    g05890(.A1(new_n6146_), .A2(new_n6145_), .A3(new_n6144_), .ZN(new_n6147_));
  NOR2_X1    g05891(.A1(new_n6147_), .A2(new_n6143_), .ZN(new_n6148_));
  AOI21_X1   g05892(.A1(new_n5617_), .A2(new_n5616_), .B(new_n5623_), .ZN(new_n6149_));
  OAI21_X1   g05893(.A1(new_n6149_), .A2(new_n5625_), .B(new_n5896_), .ZN(new_n6150_));
  NAND3_X1   g05894(.A1(new_n6148_), .A2(new_n5895_), .A3(new_n6150_), .ZN(new_n6151_));
  OAI21_X1   g05895(.A1(new_n6146_), .A2(new_n6145_), .B(new_n6144_), .ZN(new_n6152_));
  NAND3_X1   g05896(.A1(new_n6136_), .A2(new_n6142_), .A3(new_n6103_), .ZN(new_n6153_));
  NAND2_X1   g05897(.A1(new_n6152_), .A2(new_n6153_), .ZN(new_n6154_));
  NAND2_X1   g05898(.A1(new_n6150_), .A2(new_n5895_), .ZN(new_n6155_));
  NAND2_X1   g05899(.A1(new_n6155_), .A2(new_n6154_), .ZN(new_n6156_));
  OAI22_X1   g05900(.A1(new_n776_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n852_), .ZN(new_n6157_));
  AOI21_X1   g05901(.A1(\b[9] ), .A2(new_n4053_), .B(new_n6157_), .ZN(new_n6158_));
  OAI21_X1   g05902(.A1(new_n859_), .A2(new_n4727_), .B(new_n6158_), .ZN(new_n6159_));
  XOR2_X1    g05903(.A1(new_n6159_), .A2(\a[32] ), .Z(new_n6160_));
  NAND3_X1   g05904(.A1(new_n6156_), .A2(new_n6151_), .A3(new_n6160_), .ZN(new_n6161_));
  AOI21_X1   g05905(.A1(new_n5841_), .A2(new_n5621_), .B(new_n5892_), .ZN(new_n6162_));
  NOR3_X1    g05906(.A1(new_n6154_), .A2(new_n6162_), .A3(new_n5888_), .ZN(new_n6163_));
  AOI21_X1   g05907(.A1(new_n5895_), .A2(new_n6150_), .B(new_n6148_), .ZN(new_n6164_));
  INV_X1     g05908(.I(new_n6160_), .ZN(new_n6165_));
  OAI21_X1   g05909(.A1(new_n6164_), .A2(new_n6163_), .B(new_n6165_), .ZN(new_n6166_));
  NAND2_X1   g05910(.A1(new_n6166_), .A2(new_n6161_), .ZN(new_n6167_));
  NOR2_X1    g05911(.A1(new_n6098_), .A2(new_n6167_), .ZN(new_n6168_));
  NAND3_X1   g05912(.A1(new_n5908_), .A2(new_n5643_), .A3(new_n5904_), .ZN(new_n6169_));
  NAND2_X1   g05913(.A1(new_n6169_), .A2(new_n5909_), .ZN(new_n6170_));
  NOR3_X1    g05914(.A1(new_n6164_), .A2(new_n6163_), .A3(new_n6165_), .ZN(new_n6171_));
  AOI21_X1   g05915(.A1(new_n6156_), .A2(new_n6151_), .B(new_n6160_), .ZN(new_n6172_));
  NOR2_X1    g05916(.A1(new_n6171_), .A2(new_n6172_), .ZN(new_n6173_));
  NOR2_X1    g05917(.A1(new_n6170_), .A2(new_n6173_), .ZN(new_n6174_));
  NOR3_X1    g05918(.A1(new_n6168_), .A2(new_n6174_), .A3(new_n6096_), .ZN(new_n6175_));
  NAND2_X1   g05919(.A1(new_n6170_), .A2(new_n6173_), .ZN(new_n6176_));
  NAND2_X1   g05920(.A1(new_n6098_), .A2(new_n6167_), .ZN(new_n6177_));
  AOI21_X1   g05921(.A1(new_n6177_), .A2(new_n6176_), .B(new_n6095_), .ZN(new_n6178_));
  NOR2_X1    g05922(.A1(new_n6175_), .A2(new_n6178_), .ZN(new_n6179_));
  NAND3_X1   g05923(.A1(new_n6091_), .A2(new_n6179_), .A3(new_n5923_), .ZN(new_n6180_));
  AOI21_X1   g05924(.A1(new_n5922_), .A2(new_n5654_), .B(new_n5919_), .ZN(new_n6181_));
  NAND3_X1   g05925(.A1(new_n6177_), .A2(new_n6176_), .A3(new_n6095_), .ZN(new_n6182_));
  OAI21_X1   g05926(.A1(new_n6168_), .A2(new_n6174_), .B(new_n6096_), .ZN(new_n6183_));
  NAND2_X1   g05927(.A1(new_n6183_), .A2(new_n6182_), .ZN(new_n6184_));
  OAI21_X1   g05928(.A1(new_n6181_), .A2(new_n5915_), .B(new_n6184_), .ZN(new_n6185_));
  NAND3_X1   g05929(.A1(new_n6185_), .A2(new_n6180_), .A3(new_n6090_), .ZN(new_n6186_));
  INV_X1     g05930(.I(new_n6090_), .ZN(new_n6187_));
  NOR3_X1    g05931(.A1(new_n6181_), .A2(new_n6184_), .A3(new_n5915_), .ZN(new_n6188_));
  AOI21_X1   g05932(.A1(new_n6091_), .A2(new_n5923_), .B(new_n6179_), .ZN(new_n6189_));
  OAI21_X1   g05933(.A1(new_n6189_), .A2(new_n6188_), .B(new_n6187_), .ZN(new_n6190_));
  NAND2_X1   g05934(.A1(new_n6190_), .A2(new_n6186_), .ZN(new_n6191_));
  AOI21_X1   g05935(.A1(new_n5948_), .A2(new_n5935_), .B(new_n6191_), .ZN(new_n6192_));
  NOR3_X1    g05936(.A1(new_n6189_), .A2(new_n6188_), .A3(new_n6187_), .ZN(new_n6193_));
  AOI21_X1   g05937(.A1(new_n6185_), .A2(new_n6180_), .B(new_n6090_), .ZN(new_n6194_));
  NOR2_X1    g05938(.A1(new_n6193_), .A2(new_n6194_), .ZN(new_n6195_));
  NOR3_X1    g05939(.A1(new_n5939_), .A2(new_n5941_), .A3(new_n6195_), .ZN(new_n6196_));
  OAI21_X1   g05940(.A1(new_n6196_), .A2(new_n6192_), .B(new_n6086_), .ZN(new_n6197_));
  OAI21_X1   g05941(.A1(new_n5939_), .A2(new_n5941_), .B(new_n6195_), .ZN(new_n6198_));
  NAND3_X1   g05942(.A1(new_n5948_), .A2(new_n6191_), .A3(new_n5935_), .ZN(new_n6199_));
  NAND3_X1   g05943(.A1(new_n6198_), .A2(new_n6199_), .A3(new_n6085_), .ZN(new_n6200_));
  NAND2_X1   g05944(.A1(new_n6197_), .A2(new_n6200_), .ZN(new_n6201_));
  NOR3_X1    g05945(.A1(new_n5939_), .A2(new_n5945_), .A3(new_n5947_), .ZN(new_n6202_));
  INV_X1     g05946(.I(new_n6202_), .ZN(new_n6203_));
  AOI21_X1   g05947(.A1(new_n5952_), .A2(new_n6203_), .B(new_n6201_), .ZN(new_n6204_));
  AOI21_X1   g05948(.A1(new_n6198_), .A2(new_n6199_), .B(new_n6085_), .ZN(new_n6205_));
  NOR3_X1    g05949(.A1(new_n6196_), .A2(new_n6192_), .A3(new_n6086_), .ZN(new_n6206_));
  NOR2_X1    g05950(.A1(new_n6206_), .A2(new_n6205_), .ZN(new_n6207_));
  NOR3_X1    g05951(.A1(new_n5965_), .A2(new_n6207_), .A3(new_n6202_), .ZN(new_n6208_));
  NOR3_X1    g05952(.A1(new_n6208_), .A2(new_n6204_), .A3(new_n6081_), .ZN(new_n6209_));
  OAI21_X1   g05953(.A1(new_n5965_), .A2(new_n6202_), .B(new_n6207_), .ZN(new_n6210_));
  NAND3_X1   g05954(.A1(new_n5952_), .A2(new_n6201_), .A3(new_n6203_), .ZN(new_n6211_));
  AOI21_X1   g05955(.A1(new_n6210_), .A2(new_n6211_), .B(new_n6080_), .ZN(new_n6212_));
  NOR2_X1    g05956(.A1(new_n6209_), .A2(new_n6212_), .ZN(new_n6213_));
  OAI21_X1   g05957(.A1(new_n5969_), .A2(new_n5971_), .B(new_n6213_), .ZN(new_n6214_));
  NAND3_X1   g05958(.A1(new_n6210_), .A2(new_n6211_), .A3(new_n6080_), .ZN(new_n6215_));
  OAI21_X1   g05959(.A1(new_n6208_), .A2(new_n6204_), .B(new_n6081_), .ZN(new_n6216_));
  NAND2_X1   g05960(.A1(new_n6216_), .A2(new_n6215_), .ZN(new_n6217_));
  NAND3_X1   g05961(.A1(new_n5977_), .A2(new_n6217_), .A3(new_n5963_), .ZN(new_n6218_));
  NAND3_X1   g05962(.A1(new_n6214_), .A2(new_n6218_), .A3(new_n6076_), .ZN(new_n6219_));
  INV_X1     g05963(.I(new_n6076_), .ZN(new_n6220_));
  AOI21_X1   g05964(.A1(new_n5977_), .A2(new_n5963_), .B(new_n6217_), .ZN(new_n6221_));
  NOR3_X1    g05965(.A1(new_n5969_), .A2(new_n5971_), .A3(new_n6213_), .ZN(new_n6222_));
  OAI21_X1   g05966(.A1(new_n6222_), .A2(new_n6221_), .B(new_n6220_), .ZN(new_n6223_));
  NAND2_X1   g05967(.A1(new_n6223_), .A2(new_n6219_), .ZN(new_n6224_));
  OAI21_X1   g05968(.A1(new_n5991_), .A2(new_n6072_), .B(new_n6224_), .ZN(new_n6225_));
  INV_X1     g05969(.I(new_n6072_), .ZN(new_n6226_));
  NOR3_X1    g05970(.A1(new_n6222_), .A2(new_n6221_), .A3(new_n6220_), .ZN(new_n6227_));
  AOI21_X1   g05971(.A1(new_n6214_), .A2(new_n6218_), .B(new_n6076_), .ZN(new_n6228_));
  NOR2_X1    g05972(.A1(new_n6227_), .A2(new_n6228_), .ZN(new_n6229_));
  NAND3_X1   g05973(.A1(new_n5981_), .A2(new_n6229_), .A3(new_n6226_), .ZN(new_n6230_));
  OAI22_X1   g05974(.A1(new_n993_), .A2(new_n3592_), .B1(new_n3185_), .B2(new_n997_), .ZN(new_n6231_));
  AOI21_X1   g05975(.A1(\b[27] ), .A2(new_n1486_), .B(new_n6231_), .ZN(new_n6232_));
  OAI21_X1   g05976(.A1(new_n5369_), .A2(new_n1323_), .B(new_n6232_), .ZN(new_n6233_));
  XOR2_X1    g05977(.A1(new_n6233_), .A2(\a[14] ), .Z(new_n6234_));
  AOI21_X1   g05978(.A1(new_n6225_), .A2(new_n6230_), .B(new_n6234_), .ZN(new_n6235_));
  AOI21_X1   g05979(.A1(new_n5981_), .A2(new_n6226_), .B(new_n6229_), .ZN(new_n6236_));
  NOR3_X1    g05980(.A1(new_n5991_), .A2(new_n6072_), .A3(new_n6224_), .ZN(new_n6237_));
  XOR2_X1    g05981(.A1(new_n6233_), .A2(new_n1002_), .Z(new_n6238_));
  NOR3_X1    g05982(.A1(new_n6237_), .A2(new_n6236_), .A3(new_n6238_), .ZN(new_n6239_));
  NOR2_X1    g05983(.A1(new_n6239_), .A2(new_n6235_), .ZN(new_n6240_));
  AOI21_X1   g05984(.A1(new_n6002_), .A2(new_n5989_), .B(new_n6240_), .ZN(new_n6241_));
  OAI21_X1   g05985(.A1(new_n5111_), .A2(new_n5267_), .B(new_n5265_), .ZN(new_n6242_));
  OAI21_X1   g05986(.A1(new_n6242_), .A2(new_n5535_), .B(new_n5533_), .ZN(new_n6243_));
  AOI21_X1   g05987(.A1(new_n6243_), .A2(new_n5711_), .B(new_n5707_), .ZN(new_n6244_));
  NOR3_X1    g05988(.A1(new_n6244_), .A2(new_n5714_), .A3(new_n5994_), .ZN(new_n6245_));
  OAI21_X1   g05989(.A1(new_n6237_), .A2(new_n6236_), .B(new_n6238_), .ZN(new_n6246_));
  NAND3_X1   g05990(.A1(new_n6225_), .A2(new_n6230_), .A3(new_n6234_), .ZN(new_n6247_));
  NAND2_X1   g05991(.A1(new_n6246_), .A2(new_n6247_), .ZN(new_n6248_));
  NOR3_X1    g05992(.A1(new_n6245_), .A2(new_n5999_), .A3(new_n6248_), .ZN(new_n6249_));
  NOR3_X1    g05993(.A1(new_n6249_), .A2(new_n6241_), .A3(new_n6071_), .ZN(new_n6250_));
  XOR2_X1    g05994(.A1(new_n6070_), .A2(\a[11] ), .Z(new_n6251_));
  OAI21_X1   g05995(.A1(new_n6245_), .A2(new_n5999_), .B(new_n6248_), .ZN(new_n6252_));
  NAND3_X1   g05996(.A1(new_n6002_), .A2(new_n5989_), .A3(new_n6240_), .ZN(new_n6253_));
  AOI21_X1   g05997(.A1(new_n6252_), .A2(new_n6253_), .B(new_n6251_), .ZN(new_n6254_));
  NOR2_X1    g05998(.A1(new_n6250_), .A2(new_n6254_), .ZN(new_n6255_));
  NAND3_X1   g05999(.A1(new_n6067_), .A2(new_n6014_), .A3(new_n6255_), .ZN(new_n6256_));
  AOI21_X1   g06000(.A1(new_n5544_), .A2(new_n5547_), .B(new_n5545_), .ZN(new_n6257_));
  OAI21_X1   g06001(.A1(new_n6257_), .A2(new_n5726_), .B(new_n5730_), .ZN(new_n6258_));
  AOI21_X1   g06002(.A1(new_n6258_), .A2(new_n5732_), .B(new_n6010_), .ZN(new_n6259_));
  NAND3_X1   g06003(.A1(new_n6252_), .A2(new_n6253_), .A3(new_n6251_), .ZN(new_n6260_));
  OAI21_X1   g06004(.A1(new_n6249_), .A2(new_n6241_), .B(new_n6071_), .ZN(new_n6261_));
  NAND2_X1   g06005(.A1(new_n6261_), .A2(new_n6260_), .ZN(new_n6262_));
  OAI21_X1   g06006(.A1(new_n6259_), .A2(new_n6008_), .B(new_n6262_), .ZN(new_n6263_));
  AOI21_X1   g06007(.A1(new_n6263_), .A2(new_n6256_), .B(new_n6063_), .ZN(new_n6264_));
  OR2_X2     g06008(.A1(new_n6062_), .A2(new_n6059_), .Z(new_n6265_));
  NOR3_X1    g06009(.A1(new_n6259_), .A2(new_n6008_), .A3(new_n6262_), .ZN(new_n6266_));
  AOI21_X1   g06010(.A1(new_n6067_), .A2(new_n6014_), .B(new_n6255_), .ZN(new_n6267_));
  NOR3_X1    g06011(.A1(new_n6265_), .A2(new_n6266_), .A3(new_n6267_), .ZN(new_n6268_));
  NOR2_X1    g06012(.A1(new_n6268_), .A2(new_n6264_), .ZN(new_n6269_));
  AOI21_X1   g06013(.A1(new_n5741_), .A2(new_n5738_), .B(new_n5734_), .ZN(new_n6270_));
  NOR3_X1    g06014(.A1(new_n6270_), .A2(new_n5742_), .A3(new_n6029_), .ZN(new_n6271_));
  OAI21_X1   g06015(.A1(new_n6271_), .A2(new_n6030_), .B(new_n6269_), .ZN(new_n6272_));
  OAI21_X1   g06016(.A1(new_n6266_), .A2(new_n6267_), .B(new_n6265_), .ZN(new_n6273_));
  NAND3_X1   g06017(.A1(new_n6263_), .A2(new_n6256_), .A3(new_n6063_), .ZN(new_n6274_));
  NAND2_X1   g06018(.A1(new_n6273_), .A2(new_n6274_), .ZN(new_n6275_));
  NAND3_X1   g06019(.A1(new_n5806_), .A2(new_n5751_), .A3(new_n6021_), .ZN(new_n6276_));
  NAND3_X1   g06020(.A1(new_n6276_), .A2(new_n6025_), .A3(new_n6275_), .ZN(new_n6277_));
  NAND3_X1   g06021(.A1(new_n6272_), .A2(new_n6277_), .A3(new_n6054_), .ZN(new_n6278_));
  INV_X1     g06022(.I(new_n6278_), .ZN(new_n6279_));
  AOI21_X1   g06023(.A1(new_n6272_), .A2(new_n6277_), .B(new_n6054_), .ZN(new_n6280_));
  NOR2_X1    g06024(.A1(new_n6279_), .A2(new_n6280_), .ZN(new_n6281_));
  XOR2_X1    g06025(.A1(new_n6050_), .A2(new_n6281_), .Z(new_n6282_));
  INV_X1     g06026(.I(new_n6282_), .ZN(new_n6283_));
  INV_X1     g06027(.I(\b[40] ), .ZN(new_n6284_));
  INV_X1     g06028(.I(\b[41] ), .ZN(new_n6285_));
  OAI22_X1   g06029(.A1(new_n277_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n262_), .ZN(new_n6286_));
  AOI21_X1   g06030(.A1(\b[39] ), .A2(new_n283_), .B(new_n6286_), .ZN(new_n6287_));
  OAI21_X1   g06031(.A1(new_n5789_), .A2(new_n6284_), .B(\b[39] ), .ZN(new_n6288_));
  NAND2_X1   g06032(.A1(new_n5789_), .A2(new_n6284_), .ZN(new_n6289_));
  NAND2_X1   g06033(.A1(new_n6288_), .A2(new_n6289_), .ZN(new_n6290_));
  NAND2_X1   g06034(.A1(new_n5789_), .A2(new_n6285_), .ZN(new_n6291_));
  NOR2_X1    g06035(.A1(new_n5789_), .A2(new_n6285_), .ZN(new_n6292_));
  INV_X1     g06036(.I(new_n6292_), .ZN(new_n6293_));
  NAND2_X1   g06037(.A1(new_n6293_), .A2(new_n6291_), .ZN(new_n6294_));
  NAND2_X1   g06038(.A1(new_n6294_), .A2(new_n6290_), .ZN(new_n6295_));
  INV_X1     g06039(.I(new_n6291_), .ZN(new_n6296_));
  NOR2_X1    g06040(.A1(new_n6296_), .A2(new_n6292_), .ZN(new_n6297_));
  NAND3_X1   g06041(.A1(new_n6297_), .A2(new_n6288_), .A3(new_n6289_), .ZN(new_n6298_));
  NAND2_X1   g06042(.A1(new_n6298_), .A2(new_n6295_), .ZN(new_n6299_));
  OAI21_X1   g06043(.A1(new_n6299_), .A2(new_n279_), .B(new_n6287_), .ZN(new_n6300_));
  XOR2_X1    g06044(.A1(new_n6300_), .A2(\a[2] ), .Z(new_n6301_));
  NOR2_X1    g06045(.A1(new_n6283_), .A2(new_n6301_), .ZN(new_n6302_));
  NAND2_X1   g06046(.A1(new_n6283_), .A2(new_n6301_), .ZN(new_n6303_));
  INV_X1     g06047(.I(new_n6303_), .ZN(new_n6304_));
  NOR2_X1    g06048(.A1(new_n6304_), .A2(new_n6302_), .ZN(new_n6305_));
  XOR2_X1    g06049(.A1(new_n6305_), .A2(new_n6045_), .Z(\f[41] ));
  INV_X1     g06050(.I(new_n6302_), .ZN(new_n6307_));
  AOI21_X1   g06051(.A1(new_n6045_), .A2(new_n6307_), .B(new_n6304_), .ZN(new_n6308_));
  NAND2_X1   g06052(.A1(new_n5763_), .A2(new_n5760_), .ZN(new_n6309_));
  INV_X1     g06053(.I(new_n6309_), .ZN(new_n6310_));
  AOI22_X1   g06054(.A1(new_n800_), .A2(\b[38] ), .B1(\b[39] ), .B2(new_n333_), .ZN(new_n6311_));
  OAI21_X1   g06055(.A1(new_n5312_), .A2(new_n392_), .B(new_n6311_), .ZN(new_n6312_));
  AOI21_X1   g06056(.A1(new_n6310_), .A2(new_n330_), .B(new_n6312_), .ZN(new_n6313_));
  XOR2_X1    g06057(.A1(new_n6313_), .A2(new_n312_), .Z(new_n6314_));
  INV_X1     g06058(.I(new_n6122_), .ZN(new_n6315_));
  NAND2_X1   g06059(.A1(new_n6115_), .A2(\b[1] ), .ZN(new_n6316_));
  AOI22_X1   g06060(.A1(new_n6108_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n6111_), .ZN(new_n6317_));
  NAND2_X1   g06061(.A1(new_n299_), .A2(new_n6105_), .ZN(new_n6318_));
  NAND3_X1   g06062(.A1(new_n6318_), .A2(new_n6317_), .A3(new_n6316_), .ZN(new_n6319_));
  XOR2_X1    g06063(.A1(new_n6319_), .A2(new_n5849_), .Z(new_n6320_));
  XNOR2_X1   g06064(.A1(\a[41] ), .A2(\a[42] ), .ZN(new_n6321_));
  NOR2_X1    g06065(.A1(new_n6321_), .A2(new_n258_), .ZN(new_n6322_));
  INV_X1     g06066(.I(new_n6322_), .ZN(new_n6323_));
  NAND2_X1   g06067(.A1(new_n6320_), .A2(new_n6323_), .ZN(new_n6324_));
  XOR2_X1    g06068(.A1(new_n6319_), .A2(\a[41] ), .Z(new_n6325_));
  NAND2_X1   g06069(.A1(new_n6325_), .A2(new_n6322_), .ZN(new_n6326_));
  NAND2_X1   g06070(.A1(new_n6324_), .A2(new_n6326_), .ZN(new_n6327_));
  XOR2_X1    g06071(.A1(new_n6327_), .A2(new_n6315_), .Z(new_n6328_));
  INV_X1     g06072(.I(new_n6328_), .ZN(new_n6329_));
  OAI22_X1   g06073(.A1(new_n438_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n377_), .ZN(new_n6330_));
  AOI21_X1   g06074(.A1(\b[4] ), .A2(new_n5420_), .B(new_n6330_), .ZN(new_n6331_));
  OAI21_X1   g06075(.A1(new_n450_), .A2(new_n6124_), .B(new_n6331_), .ZN(new_n6332_));
  XOR2_X1    g06076(.A1(new_n6332_), .A2(\a[38] ), .Z(new_n6333_));
  INV_X1     g06077(.I(new_n6333_), .ZN(new_n6334_));
  NOR2_X1    g06078(.A1(new_n6123_), .A2(new_n6133_), .ZN(new_n6335_));
  AOI21_X1   g06079(.A1(new_n6135_), .A2(new_n6137_), .B(new_n6335_), .ZN(new_n6336_));
  NOR2_X1    g06080(.A1(new_n6336_), .A2(new_n6334_), .ZN(new_n6337_));
  NOR3_X1    g06081(.A1(new_n6145_), .A2(new_n6335_), .A3(new_n6333_), .ZN(new_n6338_));
  OR3_X2     g06082(.A1(new_n6338_), .A2(new_n6329_), .A3(new_n6337_), .Z(new_n6339_));
  OAI21_X1   g06083(.A1(new_n6338_), .A2(new_n6337_), .B(new_n6329_), .ZN(new_n6340_));
  NAND2_X1   g06084(.A1(new_n6339_), .A2(new_n6340_), .ZN(new_n6341_));
  AOI22_X1   g06085(.A1(new_n4918_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n4921_), .ZN(new_n6342_));
  OAI21_X1   g06086(.A1(new_n471_), .A2(new_n6099_), .B(new_n6342_), .ZN(new_n6343_));
  AOI21_X1   g06087(.A1(new_n676_), .A2(new_n4699_), .B(new_n6343_), .ZN(new_n6344_));
  XOR2_X1    g06088(.A1(new_n6344_), .A2(new_n4446_), .Z(new_n6345_));
  INV_X1     g06089(.I(new_n6345_), .ZN(new_n6346_));
  AOI21_X1   g06090(.A1(new_n6151_), .A2(new_n6153_), .B(new_n6346_), .ZN(new_n6347_));
  NOR3_X1    g06091(.A1(new_n6163_), .A2(new_n6147_), .A3(new_n6345_), .ZN(new_n6348_));
  NOR3_X1    g06092(.A1(new_n6347_), .A2(new_n6348_), .A3(new_n6341_), .ZN(new_n6349_));
  INV_X1     g06093(.I(new_n6341_), .ZN(new_n6350_));
  OAI21_X1   g06094(.A1(new_n6163_), .A2(new_n6147_), .B(new_n6345_), .ZN(new_n6351_));
  NAND3_X1   g06095(.A1(new_n6151_), .A2(new_n6153_), .A3(new_n6346_), .ZN(new_n6352_));
  AOI21_X1   g06096(.A1(new_n6351_), .A2(new_n6352_), .B(new_n6350_), .ZN(new_n6353_));
  NOR2_X1    g06097(.A1(new_n6349_), .A2(new_n6353_), .ZN(new_n6354_));
  AOI22_X1   g06098(.A1(new_n3864_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n3869_), .ZN(new_n6355_));
  OAI21_X1   g06099(.A1(new_n776_), .A2(new_n5410_), .B(new_n6355_), .ZN(new_n6356_));
  AOI21_X1   g06100(.A1(new_n1194_), .A2(new_n3872_), .B(new_n6356_), .ZN(new_n6357_));
  XOR2_X1    g06101(.A1(new_n6357_), .A2(\a[32] ), .Z(new_n6358_));
  INV_X1     g06102(.I(new_n6358_), .ZN(new_n6359_));
  OAI21_X1   g06103(.A1(new_n6098_), .A2(new_n6167_), .B(new_n6161_), .ZN(new_n6360_));
  NAND2_X1   g06104(.A1(new_n6360_), .A2(new_n6359_), .ZN(new_n6361_));
  AOI21_X1   g06105(.A1(new_n6170_), .A2(new_n6173_), .B(new_n6171_), .ZN(new_n6362_));
  NAND2_X1   g06106(.A1(new_n6362_), .A2(new_n6358_), .ZN(new_n6363_));
  NAND2_X1   g06107(.A1(new_n6361_), .A2(new_n6363_), .ZN(new_n6364_));
  XOR2_X1    g06108(.A1(new_n6364_), .A2(new_n6354_), .Z(new_n6365_));
  OAI22_X1   g06109(.A1(new_n1268_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n1093_), .ZN(new_n6366_));
  AOI21_X1   g06110(.A1(\b[13] ), .A2(new_n3456_), .B(new_n6366_), .ZN(new_n6367_));
  OAI21_X1   g06111(.A1(new_n1275_), .A2(new_n3261_), .B(new_n6367_), .ZN(new_n6368_));
  XOR2_X1    g06112(.A1(new_n6368_), .A2(\a[29] ), .Z(new_n6369_));
  INV_X1     g06113(.I(new_n6369_), .ZN(new_n6370_));
  AOI21_X1   g06114(.A1(new_n6180_), .A2(new_n6182_), .B(new_n6370_), .ZN(new_n6371_));
  NOR3_X1    g06115(.A1(new_n6188_), .A2(new_n6175_), .A3(new_n6369_), .ZN(new_n6372_));
  NOR3_X1    g06116(.A1(new_n6372_), .A2(new_n6371_), .A3(new_n6365_), .ZN(new_n6373_));
  INV_X1     g06117(.I(new_n6354_), .ZN(new_n6374_));
  XOR2_X1    g06118(.A1(new_n6364_), .A2(new_n6374_), .Z(new_n6375_));
  OAI21_X1   g06119(.A1(new_n6188_), .A2(new_n6175_), .B(new_n6369_), .ZN(new_n6376_));
  NAND3_X1   g06120(.A1(new_n6180_), .A2(new_n6182_), .A3(new_n6370_), .ZN(new_n6377_));
  AOI21_X1   g06121(.A1(new_n6376_), .A2(new_n6377_), .B(new_n6375_), .ZN(new_n6378_));
  NOR2_X1    g06122(.A1(new_n6373_), .A2(new_n6378_), .ZN(new_n6379_));
  INV_X1     g06123(.I(new_n6379_), .ZN(new_n6380_));
  AOI22_X1   g06124(.A1(new_n2716_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n2719_), .ZN(new_n6381_));
  OAI21_X1   g06125(.A1(new_n1296_), .A2(new_n2924_), .B(new_n6381_), .ZN(new_n6382_));
  AOI21_X1   g06126(.A1(new_n2038_), .A2(new_n2722_), .B(new_n6382_), .ZN(new_n6383_));
  XOR2_X1    g06127(.A1(new_n6383_), .A2(new_n2714_), .Z(new_n6384_));
  INV_X1     g06128(.I(new_n6384_), .ZN(new_n6385_));
  AOI21_X1   g06129(.A1(new_n6198_), .A2(new_n6186_), .B(new_n6385_), .ZN(new_n6386_));
  NOR3_X1    g06130(.A1(new_n6192_), .A2(new_n6193_), .A3(new_n6384_), .ZN(new_n6387_));
  NOR3_X1    g06131(.A1(new_n6386_), .A2(new_n6387_), .A3(new_n6380_), .ZN(new_n6388_));
  OAI21_X1   g06132(.A1(new_n6192_), .A2(new_n6193_), .B(new_n6384_), .ZN(new_n6389_));
  NAND3_X1   g06133(.A1(new_n6198_), .A2(new_n6186_), .A3(new_n6385_), .ZN(new_n6390_));
  AOI21_X1   g06134(.A1(new_n6390_), .A2(new_n6389_), .B(new_n6379_), .ZN(new_n6391_));
  NOR2_X1    g06135(.A1(new_n6391_), .A2(new_n6388_), .ZN(new_n6392_));
  INV_X1     g06136(.I(new_n6392_), .ZN(new_n6393_));
  AOI22_X1   g06137(.A1(new_n2202_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n2205_), .ZN(new_n6394_));
  OAI21_X1   g06138(.A1(new_n1859_), .A2(new_n2370_), .B(new_n6394_), .ZN(new_n6395_));
  AOI21_X1   g06139(.A1(new_n2032_), .A2(new_n2208_), .B(new_n6395_), .ZN(new_n6396_));
  XOR2_X1    g06140(.A1(new_n6396_), .A2(new_n2200_), .Z(new_n6397_));
  INV_X1     g06141(.I(new_n6397_), .ZN(new_n6398_));
  AOI21_X1   g06142(.A1(new_n6210_), .A2(new_n6200_), .B(new_n6398_), .ZN(new_n6399_));
  NOR3_X1    g06143(.A1(new_n6204_), .A2(new_n6206_), .A3(new_n6397_), .ZN(new_n6400_));
  NOR3_X1    g06144(.A1(new_n6399_), .A2(new_n6400_), .A3(new_n6393_), .ZN(new_n6401_));
  OAI21_X1   g06145(.A1(new_n6204_), .A2(new_n6206_), .B(new_n6397_), .ZN(new_n6402_));
  NAND3_X1   g06146(.A1(new_n6210_), .A2(new_n6200_), .A3(new_n6398_), .ZN(new_n6403_));
  AOI21_X1   g06147(.A1(new_n6403_), .A2(new_n6402_), .B(new_n6392_), .ZN(new_n6404_));
  NOR2_X1    g06148(.A1(new_n6404_), .A2(new_n6401_), .ZN(new_n6405_));
  INV_X1     g06149(.I(new_n6405_), .ZN(new_n6406_));
  AOI22_X1   g06150(.A1(new_n1738_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n1743_), .ZN(new_n6407_));
  OAI21_X1   g06151(.A1(new_n2142_), .A2(new_n1931_), .B(new_n6407_), .ZN(new_n6408_));
  AOI21_X1   g06152(.A1(new_n3033_), .A2(new_n1746_), .B(new_n6408_), .ZN(new_n6409_));
  XOR2_X1    g06153(.A1(new_n6409_), .A2(new_n1736_), .Z(new_n6410_));
  INV_X1     g06154(.I(new_n6410_), .ZN(new_n6411_));
  AOI21_X1   g06155(.A1(new_n6214_), .A2(new_n6215_), .B(new_n6411_), .ZN(new_n6412_));
  NOR3_X1    g06156(.A1(new_n6221_), .A2(new_n6209_), .A3(new_n6410_), .ZN(new_n6413_));
  NOR3_X1    g06157(.A1(new_n6412_), .A2(new_n6413_), .A3(new_n6406_), .ZN(new_n6414_));
  OAI21_X1   g06158(.A1(new_n6221_), .A2(new_n6209_), .B(new_n6410_), .ZN(new_n6415_));
  NAND3_X1   g06159(.A1(new_n6214_), .A2(new_n6215_), .A3(new_n6411_), .ZN(new_n6416_));
  AOI21_X1   g06160(.A1(new_n6416_), .A2(new_n6415_), .B(new_n6405_), .ZN(new_n6417_));
  NOR2_X1    g06161(.A1(new_n6417_), .A2(new_n6414_), .ZN(new_n6418_));
  INV_X1     g06162(.I(new_n6418_), .ZN(new_n6419_));
  OAI22_X1   g06163(.A1(new_n1592_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n1505_), .ZN(new_n6420_));
  AOI21_X1   g06164(.A1(\b[25] ), .A2(new_n1584_), .B(new_n6420_), .ZN(new_n6421_));
  OAI21_X1   g06165(.A1(new_n3165_), .A2(new_n1732_), .B(new_n6421_), .ZN(new_n6422_));
  XOR2_X1    g06166(.A1(new_n6422_), .A2(\a[17] ), .Z(new_n6423_));
  INV_X1     g06167(.I(new_n6423_), .ZN(new_n6424_));
  OAI21_X1   g06168(.A1(new_n5991_), .A2(new_n6072_), .B(new_n6229_), .ZN(new_n6425_));
  AOI21_X1   g06169(.A1(new_n6425_), .A2(new_n6219_), .B(new_n6424_), .ZN(new_n6426_));
  AOI21_X1   g06170(.A1(new_n5981_), .A2(new_n6226_), .B(new_n6224_), .ZN(new_n6427_));
  NOR3_X1    g06171(.A1(new_n6427_), .A2(new_n6227_), .A3(new_n6423_), .ZN(new_n6428_));
  NOR3_X1    g06172(.A1(new_n6426_), .A2(new_n6428_), .A3(new_n6419_), .ZN(new_n6429_));
  OAI21_X1   g06173(.A1(new_n6427_), .A2(new_n6227_), .B(new_n6423_), .ZN(new_n6430_));
  NAND3_X1   g06174(.A1(new_n6425_), .A2(new_n6219_), .A3(new_n6424_), .ZN(new_n6431_));
  AOI21_X1   g06175(.A1(new_n6431_), .A2(new_n6430_), .B(new_n6418_), .ZN(new_n6432_));
  NOR2_X1    g06176(.A1(new_n6432_), .A2(new_n6429_), .ZN(new_n6433_));
  OAI22_X1   g06177(.A1(new_n993_), .A2(new_n3624_), .B1(new_n3592_), .B2(new_n997_), .ZN(new_n6434_));
  AOI21_X1   g06178(.A1(\b[28] ), .A2(new_n1486_), .B(new_n6434_), .ZN(new_n6435_));
  OAI21_X1   g06179(.A1(new_n3634_), .A2(new_n1323_), .B(new_n6435_), .ZN(new_n6436_));
  XOR2_X1    g06180(.A1(new_n6436_), .A2(\a[14] ), .Z(new_n6437_));
  INV_X1     g06181(.I(new_n6437_), .ZN(new_n6438_));
  AOI21_X1   g06182(.A1(new_n6225_), .A2(new_n6230_), .B(new_n6238_), .ZN(new_n6439_));
  INV_X1     g06183(.I(new_n6439_), .ZN(new_n6440_));
  AOI21_X1   g06184(.A1(new_n6252_), .A2(new_n6440_), .B(new_n6438_), .ZN(new_n6441_));
  NOR3_X1    g06185(.A1(new_n6241_), .A2(new_n6437_), .A3(new_n6439_), .ZN(new_n6442_));
  NOR2_X1    g06186(.A1(new_n6441_), .A2(new_n6442_), .ZN(new_n6443_));
  NAND2_X1   g06187(.A1(new_n6443_), .A2(new_n6433_), .ZN(new_n6444_));
  INV_X1     g06188(.I(new_n6433_), .ZN(new_n6445_));
  OAI21_X1   g06189(.A1(new_n6241_), .A2(new_n6439_), .B(new_n6437_), .ZN(new_n6446_));
  NAND3_X1   g06190(.A1(new_n6252_), .A2(new_n6438_), .A3(new_n6440_), .ZN(new_n6447_));
  NAND2_X1   g06191(.A1(new_n6447_), .A2(new_n6446_), .ZN(new_n6448_));
  NAND2_X1   g06192(.A1(new_n6448_), .A2(new_n6445_), .ZN(new_n6449_));
  NAND2_X1   g06193(.A1(new_n6444_), .A2(new_n6449_), .ZN(new_n6450_));
  INV_X1     g06194(.I(new_n4223_), .ZN(new_n6451_));
  OAI22_X1   g06195(.A1(new_n713_), .A2(new_n4638_), .B1(new_n4023_), .B2(new_n717_), .ZN(new_n6452_));
  AOI21_X1   g06196(.A1(\b[31] ), .A2(new_n1126_), .B(new_n6452_), .ZN(new_n6453_));
  OAI21_X1   g06197(.A1(new_n6451_), .A2(new_n986_), .B(new_n6453_), .ZN(new_n6454_));
  XOR2_X1    g06198(.A1(new_n6454_), .A2(\a[11] ), .Z(new_n6455_));
  OAI21_X1   g06199(.A1(new_n6266_), .A2(new_n6250_), .B(new_n6455_), .ZN(new_n6456_));
  INV_X1     g06200(.I(new_n6455_), .ZN(new_n6457_));
  NAND3_X1   g06201(.A1(new_n6256_), .A2(new_n6260_), .A3(new_n6457_), .ZN(new_n6458_));
  NAND2_X1   g06202(.A1(new_n6456_), .A2(new_n6458_), .ZN(new_n6459_));
  NOR2_X1    g06203(.A1(new_n6459_), .A2(new_n6450_), .ZN(new_n6460_));
  NOR2_X1    g06204(.A1(new_n6448_), .A2(new_n6445_), .ZN(new_n6461_));
  NOR2_X1    g06205(.A1(new_n6443_), .A2(new_n6433_), .ZN(new_n6462_));
  NOR2_X1    g06206(.A1(new_n6462_), .A2(new_n6461_), .ZN(new_n6463_));
  AOI21_X1   g06207(.A1(new_n6456_), .A2(new_n6458_), .B(new_n6463_), .ZN(new_n6464_));
  NOR2_X1    g06208(.A1(new_n6460_), .A2(new_n6464_), .ZN(new_n6465_));
  AOI21_X1   g06209(.A1(new_n6276_), .A2(new_n6025_), .B(new_n6275_), .ZN(new_n6466_));
  AOI22_X1   g06210(.A1(new_n518_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n636_), .ZN(new_n6467_));
  OAI21_X1   g06211(.A1(new_n4639_), .A2(new_n917_), .B(new_n6467_), .ZN(new_n6468_));
  AOI21_X1   g06212(.A1(new_n5594_), .A2(new_n618_), .B(new_n6468_), .ZN(new_n6469_));
  XOR2_X1    g06213(.A1(new_n6469_), .A2(new_n488_), .Z(new_n6470_));
  OAI21_X1   g06214(.A1(new_n6466_), .A2(new_n6268_), .B(new_n6470_), .ZN(new_n6471_));
  INV_X1     g06215(.I(new_n6470_), .ZN(new_n6472_));
  NAND3_X1   g06216(.A1(new_n6272_), .A2(new_n6274_), .A3(new_n6472_), .ZN(new_n6473_));
  NAND3_X1   g06217(.A1(new_n6473_), .A2(new_n6471_), .A3(new_n6465_), .ZN(new_n6474_));
  XOR2_X1    g06218(.A1(new_n6459_), .A2(new_n6463_), .Z(new_n6475_));
  AOI21_X1   g06219(.A1(new_n6272_), .A2(new_n6274_), .B(new_n6472_), .ZN(new_n6476_));
  NOR3_X1    g06220(.A1(new_n6466_), .A2(new_n6268_), .A3(new_n6470_), .ZN(new_n6477_));
  OAI21_X1   g06221(.A1(new_n6476_), .A2(new_n6477_), .B(new_n6475_), .ZN(new_n6478_));
  AOI21_X1   g06222(.A1(new_n6478_), .A2(new_n6474_), .B(new_n6314_), .ZN(new_n6479_));
  XOR2_X1    g06223(.A1(new_n6313_), .A2(\a[5] ), .Z(new_n6480_));
  NOR3_X1    g06224(.A1(new_n6476_), .A2(new_n6477_), .A3(new_n6475_), .ZN(new_n6481_));
  AOI21_X1   g06225(.A1(new_n6473_), .A2(new_n6471_), .B(new_n6465_), .ZN(new_n6482_));
  NOR3_X1    g06226(.A1(new_n6482_), .A2(new_n6481_), .A3(new_n6480_), .ZN(new_n6483_));
  NOR2_X1    g06227(.A1(new_n6483_), .A2(new_n6479_), .ZN(new_n6484_));
  OAI21_X1   g06228(.A1(new_n6050_), .A2(new_n6280_), .B(new_n6278_), .ZN(new_n6485_));
  AOI22_X1   g06229(.A1(new_n267_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n261_), .ZN(new_n6486_));
  OAI21_X1   g06230(.A1(new_n6284_), .A2(new_n284_), .B(new_n6486_), .ZN(new_n6487_));
  AOI21_X1   g06231(.A1(new_n6291_), .A2(\b[40] ), .B(\b[39] ), .ZN(new_n6488_));
  NOR2_X1    g06232(.A1(new_n6292_), .A2(\b[40] ), .ZN(new_n6489_));
  INV_X1     g06233(.I(\b[42] ), .ZN(new_n6490_));
  NOR2_X1    g06234(.A1(new_n6490_), .A2(\b[41] ), .ZN(new_n6491_));
  NOR2_X1    g06235(.A1(new_n6285_), .A2(\b[42] ), .ZN(new_n6492_));
  OAI22_X1   g06236(.A1(new_n6488_), .A2(new_n6489_), .B1(new_n6491_), .B2(new_n6492_), .ZN(new_n6493_));
  NOR2_X1    g06237(.A1(new_n6488_), .A2(new_n6489_), .ZN(new_n6494_));
  NOR2_X1    g06238(.A1(new_n6285_), .A2(new_n6490_), .ZN(new_n6495_));
  NOR2_X1    g06239(.A1(\b[41] ), .A2(\b[42] ), .ZN(new_n6496_));
  OAI21_X1   g06240(.A1(new_n6495_), .A2(new_n6496_), .B(new_n6494_), .ZN(new_n6497_));
  AOI21_X1   g06241(.A1(new_n6497_), .A2(new_n6493_), .B(new_n279_), .ZN(new_n6498_));
  NOR2_X1    g06242(.A1(new_n6498_), .A2(new_n6487_), .ZN(new_n6499_));
  NOR2_X1    g06243(.A1(new_n6499_), .A2(new_n270_), .ZN(new_n6500_));
  NOR3_X1    g06244(.A1(new_n6498_), .A2(\a[2] ), .A3(new_n6487_), .ZN(new_n6501_));
  NOR2_X1    g06245(.A1(new_n6500_), .A2(new_n6501_), .ZN(new_n6502_));
  NOR2_X1    g06246(.A1(new_n6502_), .A2(new_n6485_), .ZN(new_n6503_));
  INV_X1     g06247(.I(new_n6503_), .ZN(new_n6504_));
  NAND2_X1   g06248(.A1(new_n6502_), .A2(new_n6485_), .ZN(new_n6505_));
  AOI21_X1   g06249(.A1(new_n6504_), .A2(new_n6505_), .B(new_n6484_), .ZN(new_n6506_));
  INV_X1     g06250(.I(new_n6484_), .ZN(new_n6507_));
  INV_X1     g06251(.I(new_n6505_), .ZN(new_n6508_));
  NOR3_X1    g06252(.A1(new_n6508_), .A2(new_n6507_), .A3(new_n6503_), .ZN(new_n6509_));
  NOR2_X1    g06253(.A1(new_n6506_), .A2(new_n6509_), .ZN(new_n6510_));
  XOR2_X1    g06254(.A1(new_n6308_), .A2(new_n6510_), .Z(\f[42] ));
  NAND3_X1   g06255(.A1(new_n6478_), .A2(new_n6474_), .A3(new_n6480_), .ZN(new_n6512_));
  AOI21_X1   g06256(.A1(new_n6478_), .A2(new_n6474_), .B(new_n6480_), .ZN(new_n6513_));
  OAI21_X1   g06257(.A1(new_n6485_), .A2(new_n6513_), .B(new_n6512_), .ZN(new_n6514_));
  NOR3_X1    g06258(.A1(new_n6266_), .A2(new_n6250_), .A3(new_n6455_), .ZN(new_n6515_));
  AOI21_X1   g06259(.A1(new_n6463_), .A2(new_n6456_), .B(new_n6515_), .ZN(new_n6516_));
  OAI22_X1   g06260(.A1(new_n713_), .A2(new_n4639_), .B1(new_n4638_), .B2(new_n717_), .ZN(new_n6517_));
  AOI21_X1   g06261(.A1(\b[32] ), .A2(new_n1126_), .B(new_n6517_), .ZN(new_n6518_));
  OAI21_X1   g06262(.A1(new_n4649_), .A2(new_n986_), .B(new_n6518_), .ZN(new_n6519_));
  XOR2_X1    g06263(.A1(new_n6519_), .A2(\a[11] ), .Z(new_n6520_));
  INV_X1     g06264(.I(new_n6520_), .ZN(new_n6521_));
  OAI21_X1   g06265(.A1(new_n5808_), .A2(new_n5994_), .B(new_n5989_), .ZN(new_n6522_));
  AOI21_X1   g06266(.A1(new_n6522_), .A2(new_n6248_), .B(new_n6439_), .ZN(new_n6523_));
  OAI21_X1   g06267(.A1(new_n6523_), .A2(new_n6438_), .B(new_n6433_), .ZN(new_n6524_));
  OAI21_X1   g06268(.A1(new_n6419_), .A2(new_n6426_), .B(new_n6431_), .ZN(new_n6525_));
  OAI22_X1   g06269(.A1(new_n1592_), .A2(new_n3185_), .B1(new_n3158_), .B2(new_n1505_), .ZN(new_n6526_));
  AOI21_X1   g06270(.A1(\b[26] ), .A2(new_n1584_), .B(new_n6526_), .ZN(new_n6527_));
  OAI21_X1   g06271(.A1(new_n3196_), .A2(new_n1732_), .B(new_n6527_), .ZN(new_n6528_));
  XOR2_X1    g06272(.A1(new_n6528_), .A2(\a[17] ), .Z(new_n6529_));
  INV_X1     g06273(.I(new_n6529_), .ZN(new_n6530_));
  NAND2_X1   g06274(.A1(new_n6415_), .A2(new_n6405_), .ZN(new_n6531_));
  OAI22_X1   g06275(.A1(new_n1751_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n1754_), .ZN(new_n6532_));
  AOI21_X1   g06276(.A1(\b[23] ), .A2(new_n1939_), .B(new_n6532_), .ZN(new_n6533_));
  OAI21_X1   g06277(.A1(new_n2655_), .A2(new_n1757_), .B(new_n6533_), .ZN(new_n6534_));
  XOR2_X1    g06278(.A1(new_n6534_), .A2(\a[20] ), .Z(new_n6535_));
  INV_X1     g06279(.I(new_n6535_), .ZN(new_n6536_));
  NOR2_X1    g06280(.A1(new_n6399_), .A2(new_n6393_), .ZN(new_n6537_));
  AOI22_X1   g06281(.A1(new_n2202_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n2205_), .ZN(new_n6538_));
  OAI21_X1   g06282(.A1(new_n1860_), .A2(new_n2370_), .B(new_n6538_), .ZN(new_n6539_));
  AOI21_X1   g06283(.A1(new_n2659_), .A2(new_n2208_), .B(new_n6539_), .ZN(new_n6540_));
  XOR2_X1    g06284(.A1(new_n6540_), .A2(new_n2200_), .Z(new_n6541_));
  INV_X1     g06285(.I(new_n6541_), .ZN(new_n6542_));
  NAND2_X1   g06286(.A1(new_n6389_), .A2(new_n6379_), .ZN(new_n6543_));
  AOI22_X1   g06287(.A1(new_n2716_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n2719_), .ZN(new_n6544_));
  OAI21_X1   g06288(.A1(new_n1432_), .A2(new_n2924_), .B(new_n6544_), .ZN(new_n6545_));
  AOI21_X1   g06289(.A1(new_n1695_), .A2(new_n2722_), .B(new_n6545_), .ZN(new_n6546_));
  XOR2_X1    g06290(.A1(new_n6546_), .A2(new_n2714_), .Z(new_n6547_));
  INV_X1     g06291(.I(new_n6547_), .ZN(new_n6548_));
  OAI21_X1   g06292(.A1(new_n6365_), .A2(new_n6371_), .B(new_n6377_), .ZN(new_n6549_));
  AOI22_X1   g06293(.A1(new_n3267_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n3270_), .ZN(new_n6550_));
  OAI21_X1   g06294(.A1(new_n1093_), .A2(new_n3475_), .B(new_n6550_), .ZN(new_n6551_));
  AOI21_X1   g06295(.A1(new_n1701_), .A2(new_n3273_), .B(new_n6551_), .ZN(new_n6552_));
  XOR2_X1    g06296(.A1(new_n6552_), .A2(new_n3264_), .Z(new_n6553_));
  OAI21_X1   g06297(.A1(new_n6362_), .A2(new_n6358_), .B(new_n6354_), .ZN(new_n6554_));
  NAND2_X1   g06298(.A1(new_n6554_), .A2(new_n6363_), .ZN(new_n6555_));
  OAI21_X1   g06299(.A1(new_n6155_), .A2(new_n6154_), .B(new_n6153_), .ZN(new_n6556_));
  AOI21_X1   g06300(.A1(new_n6556_), .A2(new_n6345_), .B(new_n6341_), .ZN(new_n6557_));
  NOR2_X1    g06301(.A1(new_n6557_), .A2(new_n6348_), .ZN(new_n6558_));
  OAI21_X1   g06302(.A1(new_n6336_), .A2(new_n6334_), .B(new_n6328_), .ZN(new_n6559_));
  INV_X1     g06303(.I(new_n6559_), .ZN(new_n6560_));
  NOR2_X1    g06304(.A1(new_n6560_), .A2(new_n6338_), .ZN(new_n6561_));
  AOI22_X1   g06305(.A1(new_n6108_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n6111_), .ZN(new_n6562_));
  NAND2_X1   g06306(.A1(new_n6115_), .A2(\b[2] ), .ZN(new_n6563_));
  NAND2_X1   g06307(.A1(new_n1725_), .A2(new_n6105_), .ZN(new_n6564_));
  NAND3_X1   g06308(.A1(new_n6564_), .A2(new_n6562_), .A3(new_n6563_), .ZN(new_n6565_));
  XOR2_X1    g06309(.A1(new_n6565_), .A2(new_n5849_), .Z(new_n6566_));
  INV_X1     g06310(.I(\a[44] ), .ZN(new_n6567_));
  XOR2_X1    g06311(.A1(\a[43] ), .A2(\a[44] ), .Z(new_n6568_));
  NOR2_X1    g06312(.A1(new_n6321_), .A2(new_n6568_), .ZN(new_n6569_));
  INV_X1     g06313(.I(\a[42] ), .ZN(new_n6570_));
  NAND3_X1   g06314(.A1(new_n5849_), .A2(new_n6570_), .A3(\a[43] ), .ZN(new_n6571_));
  INV_X1     g06315(.I(\a[43] ), .ZN(new_n6572_));
  NAND3_X1   g06316(.A1(new_n6572_), .A2(\a[41] ), .A3(\a[42] ), .ZN(new_n6573_));
  NAND2_X1   g06317(.A1(new_n6571_), .A2(new_n6573_), .ZN(new_n6574_));
  AOI22_X1   g06318(.A1(new_n6569_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n6574_), .ZN(new_n6575_));
  NOR2_X1    g06319(.A1(new_n6567_), .A2(\a[43] ), .ZN(new_n6576_));
  NOR2_X1    g06320(.A1(new_n6572_), .A2(\a[44] ), .ZN(new_n6577_));
  NOR2_X1    g06321(.A1(new_n6576_), .A2(new_n6577_), .ZN(new_n6578_));
  NOR2_X1    g06322(.A1(new_n6578_), .A2(new_n6321_), .ZN(new_n6579_));
  NAND2_X1   g06323(.A1(new_n6579_), .A2(new_n263_), .ZN(new_n6580_));
  NAND2_X1   g06324(.A1(new_n6575_), .A2(new_n6580_), .ZN(new_n6581_));
  INV_X1     g06325(.I(new_n6581_), .ZN(new_n6582_));
  NOR2_X1    g06326(.A1(new_n6582_), .A2(new_n6567_), .ZN(new_n6583_));
  NOR2_X1    g06327(.A1(new_n6581_), .A2(\a[44] ), .ZN(new_n6584_));
  NOR2_X1    g06328(.A1(new_n6583_), .A2(new_n6584_), .ZN(new_n6585_));
  NOR2_X1    g06329(.A1(new_n6322_), .A2(new_n6567_), .ZN(new_n6586_));
  INV_X1     g06330(.I(new_n6586_), .ZN(new_n6587_));
  NAND2_X1   g06331(.A1(new_n6585_), .A2(new_n6587_), .ZN(new_n6588_));
  NAND2_X1   g06332(.A1(new_n6583_), .A2(new_n6323_), .ZN(new_n6589_));
  AOI21_X1   g06333(.A1(new_n6588_), .A2(new_n6589_), .B(new_n6566_), .ZN(new_n6590_));
  INV_X1     g06334(.I(new_n6590_), .ZN(new_n6591_));
  NAND3_X1   g06335(.A1(new_n6588_), .A2(new_n6566_), .A3(new_n6589_), .ZN(new_n6592_));
  NAND2_X1   g06336(.A1(new_n6591_), .A2(new_n6592_), .ZN(new_n6593_));
  NOR2_X1    g06337(.A1(new_n6325_), .A2(new_n6322_), .ZN(new_n6594_));
  AOI21_X1   g06338(.A1(new_n6122_), .A2(new_n6326_), .B(new_n6594_), .ZN(new_n6595_));
  NAND2_X1   g06339(.A1(new_n6593_), .A2(new_n6595_), .ZN(new_n6596_));
  INV_X1     g06340(.I(new_n6592_), .ZN(new_n6597_));
  NOR2_X1    g06341(.A1(new_n6597_), .A2(new_n6590_), .ZN(new_n6598_));
  NAND2_X1   g06342(.A1(new_n6326_), .A2(new_n6122_), .ZN(new_n6599_));
  NAND2_X1   g06343(.A1(new_n6599_), .A2(new_n6324_), .ZN(new_n6600_));
  NAND2_X1   g06344(.A1(new_n6598_), .A2(new_n6600_), .ZN(new_n6601_));
  OAI22_X1   g06345(.A1(new_n471_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n438_), .ZN(new_n6602_));
  AOI21_X1   g06346(.A1(\b[5] ), .A2(new_n5420_), .B(new_n6602_), .ZN(new_n6603_));
  OAI21_X1   g06347(.A1(new_n485_), .A2(new_n6124_), .B(new_n6603_), .ZN(new_n6604_));
  XOR2_X1    g06348(.A1(new_n6604_), .A2(\a[38] ), .Z(new_n6605_));
  INV_X1     g06349(.I(new_n6605_), .ZN(new_n6606_));
  NAND3_X1   g06350(.A1(new_n6596_), .A2(new_n6601_), .A3(new_n6606_), .ZN(new_n6607_));
  NOR2_X1    g06351(.A1(new_n6598_), .A2(new_n6600_), .ZN(new_n6608_));
  NOR2_X1    g06352(.A1(new_n6593_), .A2(new_n6595_), .ZN(new_n6609_));
  OAI21_X1   g06353(.A1(new_n6609_), .A2(new_n6608_), .B(new_n6605_), .ZN(new_n6610_));
  NAND2_X1   g06354(.A1(new_n6610_), .A2(new_n6607_), .ZN(new_n6611_));
  NOR2_X1    g06355(.A1(new_n6561_), .A2(new_n6611_), .ZN(new_n6612_));
  NOR3_X1    g06356(.A1(new_n6609_), .A2(new_n6608_), .A3(new_n6605_), .ZN(new_n6613_));
  AOI21_X1   g06357(.A1(new_n6596_), .A2(new_n6601_), .B(new_n6606_), .ZN(new_n6614_));
  NOR2_X1    g06358(.A1(new_n6614_), .A2(new_n6613_), .ZN(new_n6615_));
  NOR3_X1    g06359(.A1(new_n6615_), .A2(new_n6338_), .A3(new_n6560_), .ZN(new_n6616_));
  AOI22_X1   g06360(.A1(new_n4918_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n4921_), .ZN(new_n6617_));
  OAI21_X1   g06361(.A1(new_n577_), .A2(new_n6099_), .B(new_n6617_), .ZN(new_n6618_));
  AOI21_X1   g06362(.A1(new_n1059_), .A2(new_n4699_), .B(new_n6618_), .ZN(new_n6619_));
  XOR2_X1    g06363(.A1(new_n6619_), .A2(new_n4446_), .Z(new_n6620_));
  NOR3_X1    g06364(.A1(new_n6612_), .A2(new_n6616_), .A3(new_n6620_), .ZN(new_n6621_));
  OAI21_X1   g06365(.A1(new_n6338_), .A2(new_n6560_), .B(new_n6615_), .ZN(new_n6622_));
  NAND2_X1   g06366(.A1(new_n6561_), .A2(new_n6611_), .ZN(new_n6623_));
  INV_X1     g06367(.I(new_n6620_), .ZN(new_n6624_));
  AOI21_X1   g06368(.A1(new_n6622_), .A2(new_n6623_), .B(new_n6624_), .ZN(new_n6625_));
  NOR2_X1    g06369(.A1(new_n6625_), .A2(new_n6621_), .ZN(new_n6626_));
  NOR2_X1    g06370(.A1(new_n6558_), .A2(new_n6626_), .ZN(new_n6627_));
  OAI21_X1   g06371(.A1(new_n6341_), .A2(new_n6347_), .B(new_n6352_), .ZN(new_n6628_));
  NAND3_X1   g06372(.A1(new_n6622_), .A2(new_n6623_), .A3(new_n6624_), .ZN(new_n6629_));
  OAI21_X1   g06373(.A1(new_n6612_), .A2(new_n6616_), .B(new_n6620_), .ZN(new_n6630_));
  NAND2_X1   g06374(.A1(new_n6629_), .A2(new_n6630_), .ZN(new_n6631_));
  NOR2_X1    g06375(.A1(new_n6628_), .A2(new_n6631_), .ZN(new_n6632_));
  OAI22_X1   g06376(.A1(new_n941_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n1070_), .ZN(new_n6633_));
  AOI21_X1   g06377(.A1(\b[11] ), .A2(new_n4053_), .B(new_n6633_), .ZN(new_n6634_));
  OAI21_X1   g06378(.A1(new_n1082_), .A2(new_n4727_), .B(new_n6634_), .ZN(new_n6635_));
  XOR2_X1    g06379(.A1(new_n6635_), .A2(\a[32] ), .Z(new_n6636_));
  INV_X1     g06380(.I(new_n6636_), .ZN(new_n6637_));
  NOR3_X1    g06381(.A1(new_n6627_), .A2(new_n6632_), .A3(new_n6637_), .ZN(new_n6638_));
  NAND2_X1   g06382(.A1(new_n6628_), .A2(new_n6631_), .ZN(new_n6639_));
  NAND2_X1   g06383(.A1(new_n6558_), .A2(new_n6626_), .ZN(new_n6640_));
  AOI21_X1   g06384(.A1(new_n6640_), .A2(new_n6639_), .B(new_n6636_), .ZN(new_n6641_));
  NOR2_X1    g06385(.A1(new_n6641_), .A2(new_n6638_), .ZN(new_n6642_));
  NAND2_X1   g06386(.A1(new_n6555_), .A2(new_n6642_), .ZN(new_n6643_));
  NAND3_X1   g06387(.A1(new_n6640_), .A2(new_n6639_), .A3(new_n6636_), .ZN(new_n6644_));
  OAI21_X1   g06388(.A1(new_n6627_), .A2(new_n6632_), .B(new_n6637_), .ZN(new_n6645_));
  NAND2_X1   g06389(.A1(new_n6645_), .A2(new_n6644_), .ZN(new_n6646_));
  NAND3_X1   g06390(.A1(new_n6646_), .A2(new_n6363_), .A3(new_n6554_), .ZN(new_n6647_));
  NAND3_X1   g06391(.A1(new_n6643_), .A2(new_n6647_), .A3(new_n6553_), .ZN(new_n6648_));
  INV_X1     g06392(.I(new_n6648_), .ZN(new_n6649_));
  AOI21_X1   g06393(.A1(new_n6643_), .A2(new_n6647_), .B(new_n6553_), .ZN(new_n6650_));
  NOR2_X1    g06394(.A1(new_n6649_), .A2(new_n6650_), .ZN(new_n6651_));
  NOR2_X1    g06395(.A1(new_n6549_), .A2(new_n6651_), .ZN(new_n6652_));
  NAND2_X1   g06396(.A1(new_n6376_), .A2(new_n6375_), .ZN(new_n6653_));
  INV_X1     g06397(.I(new_n6553_), .ZN(new_n6654_));
  AOI21_X1   g06398(.A1(new_n6363_), .A2(new_n6554_), .B(new_n6646_), .ZN(new_n6655_));
  NOR2_X1    g06399(.A1(new_n6555_), .A2(new_n6642_), .ZN(new_n6656_));
  OAI21_X1   g06400(.A1(new_n6655_), .A2(new_n6656_), .B(new_n6654_), .ZN(new_n6657_));
  NAND2_X1   g06401(.A1(new_n6657_), .A2(new_n6648_), .ZN(new_n6658_));
  AOI21_X1   g06402(.A1(new_n6653_), .A2(new_n6377_), .B(new_n6658_), .ZN(new_n6659_));
  NOR3_X1    g06403(.A1(new_n6652_), .A2(new_n6659_), .A3(new_n6548_), .ZN(new_n6660_));
  NAND3_X1   g06404(.A1(new_n6653_), .A2(new_n6658_), .A3(new_n6377_), .ZN(new_n6661_));
  NAND2_X1   g06405(.A1(new_n6549_), .A2(new_n6651_), .ZN(new_n6662_));
  AOI21_X1   g06406(.A1(new_n6662_), .A2(new_n6661_), .B(new_n6547_), .ZN(new_n6663_));
  NOR2_X1    g06407(.A1(new_n6660_), .A2(new_n6663_), .ZN(new_n6664_));
  NAND3_X1   g06408(.A1(new_n6543_), .A2(new_n6664_), .A3(new_n6390_), .ZN(new_n6665_));
  NOR2_X1    g06409(.A1(new_n6386_), .A2(new_n6380_), .ZN(new_n6666_));
  NAND3_X1   g06410(.A1(new_n6662_), .A2(new_n6661_), .A3(new_n6547_), .ZN(new_n6667_));
  OAI21_X1   g06411(.A1(new_n6652_), .A2(new_n6659_), .B(new_n6548_), .ZN(new_n6668_));
  NAND2_X1   g06412(.A1(new_n6668_), .A2(new_n6667_), .ZN(new_n6669_));
  OAI21_X1   g06413(.A1(new_n6666_), .A2(new_n6387_), .B(new_n6669_), .ZN(new_n6670_));
  AOI21_X1   g06414(.A1(new_n6670_), .A2(new_n6665_), .B(new_n6542_), .ZN(new_n6671_));
  NOR3_X1    g06415(.A1(new_n6666_), .A2(new_n6387_), .A3(new_n6669_), .ZN(new_n6672_));
  AOI21_X1   g06416(.A1(new_n6543_), .A2(new_n6390_), .B(new_n6664_), .ZN(new_n6673_));
  NOR3_X1    g06417(.A1(new_n6672_), .A2(new_n6673_), .A3(new_n6541_), .ZN(new_n6674_));
  NOR2_X1    g06418(.A1(new_n6674_), .A2(new_n6671_), .ZN(new_n6675_));
  NOR3_X1    g06419(.A1(new_n6537_), .A2(new_n6400_), .A3(new_n6675_), .ZN(new_n6676_));
  NAND2_X1   g06420(.A1(new_n6402_), .A2(new_n6392_), .ZN(new_n6677_));
  OAI21_X1   g06421(.A1(new_n6672_), .A2(new_n6673_), .B(new_n6541_), .ZN(new_n6678_));
  NAND3_X1   g06422(.A1(new_n6670_), .A2(new_n6665_), .A3(new_n6542_), .ZN(new_n6679_));
  NAND2_X1   g06423(.A1(new_n6678_), .A2(new_n6679_), .ZN(new_n6680_));
  AOI21_X1   g06424(.A1(new_n6677_), .A2(new_n6403_), .B(new_n6680_), .ZN(new_n6681_));
  NOR3_X1    g06425(.A1(new_n6676_), .A2(new_n6681_), .A3(new_n6536_), .ZN(new_n6682_));
  NAND3_X1   g06426(.A1(new_n6677_), .A2(new_n6680_), .A3(new_n6403_), .ZN(new_n6683_));
  OAI21_X1   g06427(.A1(new_n6393_), .A2(new_n6399_), .B(new_n6403_), .ZN(new_n6684_));
  NAND2_X1   g06428(.A1(new_n6684_), .A2(new_n6675_), .ZN(new_n6685_));
  AOI21_X1   g06429(.A1(new_n6685_), .A2(new_n6683_), .B(new_n6535_), .ZN(new_n6686_));
  NOR2_X1    g06430(.A1(new_n6686_), .A2(new_n6682_), .ZN(new_n6687_));
  NAND3_X1   g06431(.A1(new_n6531_), .A2(new_n6687_), .A3(new_n6416_), .ZN(new_n6688_));
  OAI21_X1   g06432(.A1(new_n6406_), .A2(new_n6412_), .B(new_n6416_), .ZN(new_n6689_));
  NAND3_X1   g06433(.A1(new_n6685_), .A2(new_n6683_), .A3(new_n6535_), .ZN(new_n6690_));
  OAI21_X1   g06434(.A1(new_n6676_), .A2(new_n6681_), .B(new_n6536_), .ZN(new_n6691_));
  NAND2_X1   g06435(.A1(new_n6690_), .A2(new_n6691_), .ZN(new_n6692_));
  NAND2_X1   g06436(.A1(new_n6689_), .A2(new_n6692_), .ZN(new_n6693_));
  AOI21_X1   g06437(.A1(new_n6693_), .A2(new_n6688_), .B(new_n6530_), .ZN(new_n6694_));
  NOR2_X1    g06438(.A1(new_n6412_), .A2(new_n6406_), .ZN(new_n6695_));
  NOR3_X1    g06439(.A1(new_n6695_), .A2(new_n6413_), .A3(new_n6692_), .ZN(new_n6696_));
  AOI21_X1   g06440(.A1(new_n6405_), .A2(new_n6415_), .B(new_n6413_), .ZN(new_n6697_));
  NOR2_X1    g06441(.A1(new_n6697_), .A2(new_n6687_), .ZN(new_n6698_));
  NOR3_X1    g06442(.A1(new_n6698_), .A2(new_n6696_), .A3(new_n6529_), .ZN(new_n6699_));
  NOR2_X1    g06443(.A1(new_n6699_), .A2(new_n6694_), .ZN(new_n6700_));
  NAND2_X1   g06444(.A1(new_n6525_), .A2(new_n6700_), .ZN(new_n6701_));
  NAND2_X1   g06445(.A1(new_n6430_), .A2(new_n6418_), .ZN(new_n6702_));
  OAI21_X1   g06446(.A1(new_n6698_), .A2(new_n6696_), .B(new_n6529_), .ZN(new_n6703_));
  NAND3_X1   g06447(.A1(new_n6693_), .A2(new_n6688_), .A3(new_n6530_), .ZN(new_n6704_));
  NAND2_X1   g06448(.A1(new_n6703_), .A2(new_n6704_), .ZN(new_n6705_));
  NAND3_X1   g06449(.A1(new_n6702_), .A2(new_n6705_), .A3(new_n6431_), .ZN(new_n6706_));
  OAI22_X1   g06450(.A1(new_n993_), .A2(new_n4022_), .B1(new_n3624_), .B2(new_n997_), .ZN(new_n6707_));
  AOI21_X1   g06451(.A1(\b[29] ), .A2(new_n1486_), .B(new_n6707_), .ZN(new_n6708_));
  OAI21_X1   g06452(.A1(new_n6003_), .A2(new_n1323_), .B(new_n6708_), .ZN(new_n6709_));
  XOR2_X1    g06453(.A1(new_n6709_), .A2(\a[14] ), .Z(new_n6710_));
  NAND3_X1   g06454(.A1(new_n6701_), .A2(new_n6706_), .A3(new_n6710_), .ZN(new_n6711_));
  AOI21_X1   g06455(.A1(new_n6418_), .A2(new_n6430_), .B(new_n6428_), .ZN(new_n6712_));
  NOR2_X1    g06456(.A1(new_n6712_), .A2(new_n6705_), .ZN(new_n6713_));
  NOR2_X1    g06457(.A1(new_n6426_), .A2(new_n6419_), .ZN(new_n6714_));
  NOR3_X1    g06458(.A1(new_n6714_), .A2(new_n6700_), .A3(new_n6428_), .ZN(new_n6715_));
  XOR2_X1    g06459(.A1(new_n6709_), .A2(new_n1002_), .Z(new_n6716_));
  OAI21_X1   g06460(.A1(new_n6713_), .A2(new_n6715_), .B(new_n6716_), .ZN(new_n6717_));
  NAND2_X1   g06461(.A1(new_n6717_), .A2(new_n6711_), .ZN(new_n6718_));
  AOI21_X1   g06462(.A1(new_n6524_), .A2(new_n6447_), .B(new_n6718_), .ZN(new_n6719_));
  AOI21_X1   g06463(.A1(new_n5717_), .A2(new_n5718_), .B(new_n5714_), .ZN(new_n6720_));
  AOI21_X1   g06464(.A1(new_n6720_), .A2(new_n6001_), .B(new_n5999_), .ZN(new_n6721_));
  OAI21_X1   g06465(.A1(new_n6721_), .A2(new_n6240_), .B(new_n6440_), .ZN(new_n6722_));
  AOI21_X1   g06466(.A1(new_n6722_), .A2(new_n6437_), .B(new_n6445_), .ZN(new_n6723_));
  NOR3_X1    g06467(.A1(new_n6713_), .A2(new_n6715_), .A3(new_n6716_), .ZN(new_n6724_));
  AOI21_X1   g06468(.A1(new_n6701_), .A2(new_n6706_), .B(new_n6710_), .ZN(new_n6725_));
  NOR2_X1    g06469(.A1(new_n6725_), .A2(new_n6724_), .ZN(new_n6726_));
  NOR3_X1    g06470(.A1(new_n6723_), .A2(new_n6442_), .A3(new_n6726_), .ZN(new_n6727_));
  NOR3_X1    g06471(.A1(new_n6727_), .A2(new_n6719_), .A3(new_n6521_), .ZN(new_n6728_));
  OAI21_X1   g06472(.A1(new_n6723_), .A2(new_n6442_), .B(new_n6726_), .ZN(new_n6729_));
  NAND3_X1   g06473(.A1(new_n6718_), .A2(new_n6524_), .A3(new_n6447_), .ZN(new_n6730_));
  AOI21_X1   g06474(.A1(new_n6729_), .A2(new_n6730_), .B(new_n6520_), .ZN(new_n6731_));
  NOR2_X1    g06475(.A1(new_n6728_), .A2(new_n6731_), .ZN(new_n6732_));
  NAND2_X1   g06476(.A1(new_n6516_), .A2(new_n6732_), .ZN(new_n6733_));
  AOI21_X1   g06477(.A1(new_n6256_), .A2(new_n6260_), .B(new_n6457_), .ZN(new_n6734_));
  OAI21_X1   g06478(.A1(new_n6450_), .A2(new_n6734_), .B(new_n6458_), .ZN(new_n6735_));
  NAND3_X1   g06479(.A1(new_n6729_), .A2(new_n6730_), .A3(new_n6520_), .ZN(new_n6736_));
  OAI21_X1   g06480(.A1(new_n6727_), .A2(new_n6719_), .B(new_n6521_), .ZN(new_n6737_));
  NAND2_X1   g06481(.A1(new_n6737_), .A2(new_n6736_), .ZN(new_n6738_));
  NAND2_X1   g06482(.A1(new_n6735_), .A2(new_n6738_), .ZN(new_n6739_));
  NAND2_X1   g06483(.A1(new_n6733_), .A2(new_n6739_), .ZN(new_n6740_));
  OAI22_X1   g06484(.A1(new_n610_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n612_), .ZN(new_n6741_));
  AOI21_X1   g06485(.A1(\b[35] ), .A2(new_n826_), .B(new_n6741_), .ZN(new_n6742_));
  OAI21_X1   g06486(.A1(new_n5322_), .A2(new_n624_), .B(new_n6742_), .ZN(new_n6743_));
  XOR2_X1    g06487(.A1(new_n6743_), .A2(\a[8] ), .Z(new_n6744_));
  XOR2_X1    g06488(.A1(new_n6740_), .A2(new_n6744_), .Z(new_n6745_));
  OAI21_X1   g06489(.A1(new_n6475_), .A2(new_n6476_), .B(new_n6473_), .ZN(new_n6746_));
  AOI22_X1   g06490(.A1(new_n800_), .A2(\b[39] ), .B1(\b[40] ), .B2(new_n333_), .ZN(new_n6747_));
  OAI21_X1   g06491(.A1(new_n5341_), .A2(new_n392_), .B(new_n6747_), .ZN(new_n6748_));
  INV_X1     g06492(.I(new_n6748_), .ZN(new_n6749_));
  INV_X1     g06493(.I(new_n5792_), .ZN(new_n6750_));
  OAI21_X1   g06494(.A1(new_n6750_), .A2(new_n5790_), .B(new_n330_), .ZN(new_n6751_));
  AOI21_X1   g06495(.A1(new_n6751_), .A2(new_n6749_), .B(new_n312_), .ZN(new_n6752_));
  AOI21_X1   g06496(.A1(new_n5791_), .A2(new_n5792_), .B(new_n318_), .ZN(new_n6753_));
  NOR3_X1    g06497(.A1(new_n6753_), .A2(\a[5] ), .A3(new_n6748_), .ZN(new_n6754_));
  NOR2_X1    g06498(.A1(new_n6754_), .A2(new_n6752_), .ZN(new_n6755_));
  NOR2_X1    g06499(.A1(new_n6746_), .A2(new_n6755_), .ZN(new_n6756_));
  OAI21_X1   g06500(.A1(new_n6028_), .A2(new_n6029_), .B(new_n6025_), .ZN(new_n6757_));
  AOI21_X1   g06501(.A1(new_n6757_), .A2(new_n6269_), .B(new_n6268_), .ZN(new_n6758_));
  OAI21_X1   g06502(.A1(new_n6758_), .A2(new_n6472_), .B(new_n6465_), .ZN(new_n6759_));
  OAI21_X1   g06503(.A1(new_n6753_), .A2(new_n6748_), .B(\a[5] ), .ZN(new_n6760_));
  NAND3_X1   g06504(.A1(new_n6751_), .A2(new_n312_), .A3(new_n6749_), .ZN(new_n6761_));
  NAND2_X1   g06505(.A1(new_n6760_), .A2(new_n6761_), .ZN(new_n6762_));
  AOI21_X1   g06506(.A1(new_n6759_), .A2(new_n6473_), .B(new_n6762_), .ZN(new_n6763_));
  OAI21_X1   g06507(.A1(new_n6756_), .A2(new_n6763_), .B(new_n6745_), .ZN(new_n6764_));
  INV_X1     g06508(.I(new_n6744_), .ZN(new_n6765_));
  XOR2_X1    g06509(.A1(new_n6740_), .A2(new_n6765_), .Z(new_n6766_));
  NAND3_X1   g06510(.A1(new_n6759_), .A2(new_n6762_), .A3(new_n6473_), .ZN(new_n6767_));
  NAND2_X1   g06511(.A1(new_n6272_), .A2(new_n6274_), .ZN(new_n6768_));
  AOI21_X1   g06512(.A1(new_n6768_), .A2(new_n6470_), .B(new_n6475_), .ZN(new_n6769_));
  OAI21_X1   g06513(.A1(new_n6769_), .A2(new_n6477_), .B(new_n6755_), .ZN(new_n6770_));
  NAND3_X1   g06514(.A1(new_n6770_), .A2(new_n6766_), .A3(new_n6767_), .ZN(new_n6771_));
  NAND2_X1   g06515(.A1(new_n6764_), .A2(new_n6771_), .ZN(new_n6772_));
  XOR2_X1    g06516(.A1(new_n6772_), .A2(new_n6514_), .Z(new_n6773_));
  INV_X1     g06517(.I(new_n6773_), .ZN(new_n6774_));
  INV_X1     g06518(.I(\b[43] ), .ZN(new_n6775_));
  OAI22_X1   g06519(.A1(new_n277_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n262_), .ZN(new_n6776_));
  AOI21_X1   g06520(.A1(\b[41] ), .A2(new_n283_), .B(new_n6776_), .ZN(new_n6777_));
  NOR3_X1    g06521(.A1(new_n6494_), .A2(\b[41] ), .A3(new_n6490_), .ZN(new_n6778_));
  NOR3_X1    g06522(.A1(new_n6488_), .A2(new_n6489_), .A3(new_n6285_), .ZN(new_n6779_));
  NAND2_X1   g06523(.A1(new_n6779_), .A2(new_n6490_), .ZN(new_n6780_));
  INV_X1     g06524(.I(new_n6780_), .ZN(new_n6781_));
  OAI21_X1   g06525(.A1(new_n6781_), .A2(new_n6778_), .B(\b[43] ), .ZN(new_n6782_));
  INV_X1     g06526(.I(new_n6778_), .ZN(new_n6783_));
  NAND3_X1   g06527(.A1(new_n6783_), .A2(new_n6775_), .A3(new_n6780_), .ZN(new_n6784_));
  NAND2_X1   g06528(.A1(new_n6784_), .A2(new_n6782_), .ZN(new_n6785_));
  OAI21_X1   g06529(.A1(new_n6785_), .A2(new_n279_), .B(new_n6777_), .ZN(new_n6786_));
  XOR2_X1    g06530(.A1(new_n6786_), .A2(\a[2] ), .Z(new_n6787_));
  INV_X1     g06531(.I(new_n6502_), .ZN(new_n6788_));
  XOR2_X1    g06532(.A1(new_n6484_), .A2(new_n6485_), .Z(new_n6789_));
  NOR2_X1    g06533(.A1(new_n6789_), .A2(new_n6788_), .ZN(new_n6790_));
  INV_X1     g06534(.I(new_n6790_), .ZN(new_n6791_));
  OAI21_X1   g06535(.A1(new_n6308_), .A2(new_n6510_), .B(new_n6791_), .ZN(new_n6792_));
  NAND2_X1   g06536(.A1(new_n6792_), .A2(new_n6787_), .ZN(new_n6793_));
  INV_X1     g06537(.I(new_n6787_), .ZN(new_n6794_));
  INV_X1     g06538(.I(new_n5775_), .ZN(new_n6795_));
  NOR3_X1    g06539(.A1(new_n5327_), .A2(new_n5324_), .A3(new_n5326_), .ZN(new_n6796_));
  AOI21_X1   g06540(.A1(new_n5311_), .A2(new_n5328_), .B(new_n6796_), .ZN(new_n6797_));
  INV_X1     g06541(.I(new_n5590_), .ZN(new_n6798_));
  AOI21_X1   g06542(.A1(new_n6797_), .A2(new_n5589_), .B(new_n6798_), .ZN(new_n6799_));
  INV_X1     g06543(.I(new_n5780_), .ZN(new_n6800_));
  OAI21_X1   g06544(.A1(new_n6799_), .A2(new_n6795_), .B(new_n6800_), .ZN(new_n6801_));
  AOI21_X1   g06545(.A1(new_n6801_), .A2(new_n6042_), .B(new_n6040_), .ZN(new_n6802_));
  OAI21_X1   g06546(.A1(new_n6802_), .A2(new_n6302_), .B(new_n6303_), .ZN(new_n6803_));
  OAI21_X1   g06547(.A1(new_n6508_), .A2(new_n6503_), .B(new_n6507_), .ZN(new_n6804_));
  NAND3_X1   g06548(.A1(new_n6504_), .A2(new_n6505_), .A3(new_n6484_), .ZN(new_n6805_));
  NAND2_X1   g06549(.A1(new_n6804_), .A2(new_n6805_), .ZN(new_n6806_));
  AOI21_X1   g06550(.A1(new_n6803_), .A2(new_n6806_), .B(new_n6790_), .ZN(new_n6807_));
  NAND2_X1   g06551(.A1(new_n6807_), .A2(new_n6794_), .ZN(new_n6808_));
  NAND2_X1   g06552(.A1(new_n6808_), .A2(new_n6793_), .ZN(new_n6809_));
  XOR2_X1    g06553(.A1(new_n6809_), .A2(new_n6774_), .Z(\f[43] ));
  NOR2_X1    g06554(.A1(new_n6792_), .A2(new_n6787_), .ZN(new_n6811_));
  AOI21_X1   g06555(.A1(new_n6792_), .A2(new_n6787_), .B(new_n6773_), .ZN(new_n6812_));
  NOR2_X1    g06556(.A1(new_n6812_), .A2(new_n6811_), .ZN(new_n6813_));
  NOR2_X1    g06557(.A1(new_n6745_), .A2(new_n6746_), .ZN(new_n6814_));
  AOI21_X1   g06558(.A1(new_n6465_), .A2(new_n6471_), .B(new_n6477_), .ZN(new_n6815_));
  NOR2_X1    g06559(.A1(new_n6766_), .A2(new_n6815_), .ZN(new_n6816_));
  OAI21_X1   g06560(.A1(new_n6816_), .A2(new_n6814_), .B(new_n6755_), .ZN(new_n6817_));
  OAI21_X1   g06561(.A1(new_n6772_), .A2(new_n6514_), .B(new_n6817_), .ZN(new_n6818_));
  AOI22_X1   g06562(.A1(new_n800_), .A2(\b[40] ), .B1(\b[41] ), .B2(new_n333_), .ZN(new_n6819_));
  OAI21_X1   g06563(.A1(new_n5761_), .A2(new_n392_), .B(new_n6819_), .ZN(new_n6820_));
  INV_X1     g06564(.I(new_n6820_), .ZN(new_n6821_));
  NAND3_X1   g06565(.A1(new_n6298_), .A2(new_n6295_), .A3(new_n330_), .ZN(new_n6822_));
  AOI21_X1   g06566(.A1(new_n6822_), .A2(new_n6821_), .B(new_n312_), .ZN(new_n6823_));
  NAND3_X1   g06567(.A1(new_n6822_), .A2(new_n312_), .A3(new_n6821_), .ZN(new_n6824_));
  INV_X1     g06568(.I(new_n6824_), .ZN(new_n6825_));
  NOR2_X1    g06569(.A1(new_n6825_), .A2(new_n6823_), .ZN(new_n6826_));
  AOI22_X1   g06570(.A1(new_n729_), .A2(\b[35] ), .B1(\b[34] ), .B2(new_n732_), .ZN(new_n6827_));
  OAI21_X1   g06571(.A1(new_n4638_), .A2(new_n1127_), .B(new_n6827_), .ZN(new_n6828_));
  INV_X1     g06572(.I(new_n6828_), .ZN(new_n6829_));
  NAND3_X1   g06573(.A1(new_n4675_), .A2(new_n724_), .A3(new_n4673_), .ZN(new_n6830_));
  AOI21_X1   g06574(.A1(new_n6830_), .A2(new_n6829_), .B(new_n722_), .ZN(new_n6831_));
  INV_X1     g06575(.I(new_n6831_), .ZN(new_n6832_));
  NAND3_X1   g06576(.A1(new_n6830_), .A2(new_n722_), .A3(new_n6829_), .ZN(new_n6833_));
  NAND2_X1   g06577(.A1(new_n6832_), .A2(new_n6833_), .ZN(new_n6834_));
  AOI21_X1   g06578(.A1(new_n6524_), .A2(new_n6447_), .B(new_n6724_), .ZN(new_n6835_));
  OAI22_X1   g06579(.A1(new_n993_), .A2(new_n4023_), .B1(new_n4022_), .B2(new_n997_), .ZN(new_n6836_));
  AOI21_X1   g06580(.A1(\b[30] ), .A2(new_n1486_), .B(new_n6836_), .ZN(new_n6837_));
  OAI21_X1   g06581(.A1(new_n4031_), .A2(new_n1323_), .B(new_n6837_), .ZN(new_n6838_));
  XOR2_X1    g06582(.A1(new_n6838_), .A2(\a[14] ), .Z(new_n6839_));
  NOR3_X1    g06583(.A1(new_n6698_), .A2(new_n6696_), .A3(new_n6530_), .ZN(new_n6840_));
  OAI22_X1   g06584(.A1(new_n1592_), .A2(new_n3592_), .B1(new_n3185_), .B2(new_n1505_), .ZN(new_n6841_));
  AOI21_X1   g06585(.A1(\b[27] ), .A2(new_n1584_), .B(new_n6841_), .ZN(new_n6842_));
  OAI21_X1   g06586(.A1(new_n5369_), .A2(new_n1732_), .B(new_n6842_), .ZN(new_n6843_));
  XOR2_X1    g06587(.A1(new_n6843_), .A2(\a[17] ), .Z(new_n6844_));
  INV_X1     g06588(.I(new_n6844_), .ZN(new_n6845_));
  AOI22_X1   g06589(.A1(new_n1738_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n1743_), .ZN(new_n6846_));
  OAI21_X1   g06590(.A1(new_n2495_), .A2(new_n1931_), .B(new_n6846_), .ZN(new_n6847_));
  AOI21_X1   g06591(.A1(new_n3407_), .A2(new_n1746_), .B(new_n6847_), .ZN(new_n6848_));
  XOR2_X1    g06592(.A1(new_n6848_), .A2(new_n1736_), .Z(new_n6849_));
  NOR3_X1    g06593(.A1(new_n6672_), .A2(new_n6673_), .A3(new_n6542_), .ZN(new_n6850_));
  AOI22_X1   g06594(.A1(new_n2202_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n2205_), .ZN(new_n6851_));
  OAI21_X1   g06595(.A1(new_n2027_), .A2(new_n2370_), .B(new_n6851_), .ZN(new_n6852_));
  AOI21_X1   g06596(.A1(new_n2470_), .A2(new_n2208_), .B(new_n6852_), .ZN(new_n6853_));
  XOR2_X1    g06597(.A1(new_n6853_), .A2(new_n2200_), .Z(new_n6854_));
  INV_X1     g06598(.I(new_n6854_), .ZN(new_n6855_));
  AOI22_X1   g06599(.A1(new_n2716_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n2719_), .ZN(new_n6856_));
  OAI21_X1   g06600(.A1(new_n1553_), .A2(new_n2924_), .B(new_n6856_), .ZN(new_n6857_));
  AOI21_X1   g06601(.A1(new_n2452_), .A2(new_n2722_), .B(new_n6857_), .ZN(new_n6858_));
  XOR2_X1    g06602(.A1(new_n6858_), .A2(new_n2714_), .Z(new_n6859_));
  INV_X1     g06603(.I(new_n6859_), .ZN(new_n6860_));
  AOI21_X1   g06604(.A1(new_n6643_), .A2(new_n6647_), .B(new_n6654_), .ZN(new_n6861_));
  INV_X1     g06605(.I(new_n6861_), .ZN(new_n6862_));
  OAI22_X1   g06606(.A1(new_n1432_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n1296_), .ZN(new_n6863_));
  AOI21_X1   g06607(.A1(\b[15] ), .A2(new_n3456_), .B(new_n6863_), .ZN(new_n6864_));
  OAI21_X1   g06608(.A1(new_n1444_), .A2(new_n3261_), .B(new_n6864_), .ZN(new_n6865_));
  XOR2_X1    g06609(.A1(new_n6865_), .A2(\a[29] ), .Z(new_n6866_));
  NOR2_X1    g06610(.A1(new_n6360_), .A2(new_n6359_), .ZN(new_n6867_));
  AOI21_X1   g06611(.A1(new_n6360_), .A2(new_n6359_), .B(new_n6374_), .ZN(new_n6868_));
  OAI21_X1   g06612(.A1(new_n6868_), .A2(new_n6867_), .B(new_n6644_), .ZN(new_n6869_));
  AOI22_X1   g06613(.A1(new_n3864_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n3869_), .ZN(new_n6870_));
  OAI21_X1   g06614(.A1(new_n941_), .A2(new_n5410_), .B(new_n6870_), .ZN(new_n6871_));
  AOI21_X1   g06615(.A1(new_n1449_), .A2(new_n3872_), .B(new_n6871_), .ZN(new_n6872_));
  XOR2_X1    g06616(.A1(new_n6872_), .A2(new_n3876_), .Z(new_n6873_));
  INV_X1     g06617(.I(new_n6873_), .ZN(new_n6874_));
  NAND2_X1   g06618(.A1(new_n6351_), .A2(new_n6350_), .ZN(new_n6875_));
  NAND3_X1   g06619(.A1(new_n6875_), .A2(new_n6352_), .A3(new_n6629_), .ZN(new_n6876_));
  INV_X1     g06620(.I(new_n5420_), .ZN(new_n6877_));
  AOI22_X1   g06621(.A1(new_n5155_), .A2(\b[8] ), .B1(\b[7] ), .B2(new_n5160_), .ZN(new_n6878_));
  OAI21_X1   g06622(.A1(new_n438_), .A2(new_n6877_), .B(new_n6878_), .ZN(new_n6879_));
  AOI21_X1   g06623(.A1(new_n799_), .A2(new_n5166_), .B(new_n6879_), .ZN(new_n6880_));
  XOR2_X1    g06624(.A1(new_n6880_), .A2(new_n5162_), .Z(new_n6881_));
  NAND2_X1   g06625(.A1(new_n6579_), .A2(new_n554_), .ZN(new_n6882_));
  AOI22_X1   g06626(.A1(new_n6569_), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n6574_), .ZN(new_n6883_));
  XOR2_X1    g06627(.A1(\a[41] ), .A2(\a[42] ), .Z(new_n6884_));
  NOR2_X1    g06628(.A1(new_n6576_), .A2(\a[41] ), .ZN(new_n6885_));
  NOR2_X1    g06629(.A1(new_n6577_), .A2(new_n5849_), .ZN(new_n6886_));
  NOR3_X1    g06630(.A1(new_n6885_), .A2(new_n6886_), .A3(new_n6884_), .ZN(new_n6887_));
  NAND2_X1   g06631(.A1(new_n6887_), .A2(\b[0] ), .ZN(new_n6888_));
  NAND3_X1   g06632(.A1(new_n6883_), .A2(new_n6888_), .A3(new_n6882_), .ZN(new_n6889_));
  XOR2_X1    g06633(.A1(new_n6889_), .A2(new_n6567_), .Z(new_n6890_));
  NOR3_X1    g06634(.A1(new_n6581_), .A2(new_n6567_), .A3(new_n6322_), .ZN(new_n6891_));
  INV_X1     g06635(.I(new_n6891_), .ZN(new_n6892_));
  NAND2_X1   g06636(.A1(new_n6890_), .A2(new_n6892_), .ZN(new_n6893_));
  OR4_X2     g06637(.A1(new_n6567_), .A2(new_n6889_), .A3(new_n6322_), .A4(new_n6581_), .Z(new_n6894_));
  OAI22_X1   g06638(.A1(new_n5852_), .A2(new_n377_), .B1(new_n339_), .B2(new_n5857_), .ZN(new_n6895_));
  AOI21_X1   g06639(.A1(\b[3] ), .A2(new_n6115_), .B(new_n6895_), .ZN(new_n6896_));
  OAI21_X1   g06640(.A1(new_n566_), .A2(new_n5861_), .B(new_n6896_), .ZN(new_n6897_));
  XOR2_X1    g06641(.A1(new_n6897_), .A2(\a[41] ), .Z(new_n6898_));
  AOI21_X1   g06642(.A1(new_n6893_), .A2(new_n6894_), .B(new_n6898_), .ZN(new_n6899_));
  NAND2_X1   g06643(.A1(new_n6893_), .A2(new_n6894_), .ZN(new_n6900_));
  XOR2_X1    g06644(.A1(new_n6897_), .A2(new_n5849_), .Z(new_n6901_));
  NOR2_X1    g06645(.A1(new_n6900_), .A2(new_n6901_), .ZN(new_n6902_));
  NOR2_X1    g06646(.A1(new_n6899_), .A2(new_n6902_), .ZN(new_n6903_));
  AOI21_X1   g06647(.A1(new_n6595_), .A2(new_n6592_), .B(new_n6590_), .ZN(new_n6904_));
  INV_X1     g06648(.I(new_n6904_), .ZN(new_n6905_));
  NAND2_X1   g06649(.A1(new_n6905_), .A2(new_n6903_), .ZN(new_n6906_));
  NAND2_X1   g06650(.A1(new_n6900_), .A2(new_n6901_), .ZN(new_n6907_));
  NAND3_X1   g06651(.A1(new_n6898_), .A2(new_n6893_), .A3(new_n6894_), .ZN(new_n6908_));
  NAND2_X1   g06652(.A1(new_n6907_), .A2(new_n6908_), .ZN(new_n6909_));
  NAND2_X1   g06653(.A1(new_n6909_), .A2(new_n6904_), .ZN(new_n6910_));
  AOI21_X1   g06654(.A1(new_n6906_), .A2(new_n6910_), .B(new_n6881_), .ZN(new_n6911_));
  INV_X1     g06655(.I(new_n6881_), .ZN(new_n6912_));
  NOR2_X1    g06656(.A1(new_n6909_), .A2(new_n6904_), .ZN(new_n6913_));
  NOR2_X1    g06657(.A1(new_n6905_), .A2(new_n6903_), .ZN(new_n6914_));
  NOR3_X1    g06658(.A1(new_n6914_), .A2(new_n6913_), .A3(new_n6912_), .ZN(new_n6915_));
  NOR2_X1    g06659(.A1(new_n6915_), .A2(new_n6911_), .ZN(new_n6916_));
  OAI21_X1   g06660(.A1(new_n6560_), .A2(new_n6338_), .B(new_n6610_), .ZN(new_n6917_));
  NAND3_X1   g06661(.A1(new_n6917_), .A2(new_n6916_), .A3(new_n6607_), .ZN(new_n6918_));
  OAI21_X1   g06662(.A1(new_n6914_), .A2(new_n6913_), .B(new_n6912_), .ZN(new_n6919_));
  NAND3_X1   g06663(.A1(new_n6906_), .A2(new_n6910_), .A3(new_n6881_), .ZN(new_n6920_));
  NAND2_X1   g06664(.A1(new_n6919_), .A2(new_n6920_), .ZN(new_n6921_));
  NAND2_X1   g06665(.A1(new_n6336_), .A2(new_n6334_), .ZN(new_n6922_));
  AOI21_X1   g06666(.A1(new_n6559_), .A2(new_n6922_), .B(new_n6614_), .ZN(new_n6923_));
  OAI21_X1   g06667(.A1(new_n6923_), .A2(new_n6613_), .B(new_n6921_), .ZN(new_n6924_));
  OAI22_X1   g06668(.A1(new_n852_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n776_), .ZN(new_n6925_));
  AOI21_X1   g06669(.A1(\b[9] ), .A2(new_n4706_), .B(new_n6925_), .ZN(new_n6926_));
  OAI21_X1   g06670(.A1(new_n859_), .A2(new_n4458_), .B(new_n6926_), .ZN(new_n6927_));
  XOR2_X1    g06671(.A1(new_n6927_), .A2(\a[35] ), .Z(new_n6928_));
  NAND3_X1   g06672(.A1(new_n6918_), .A2(new_n6924_), .A3(new_n6928_), .ZN(new_n6929_));
  NOR3_X1    g06673(.A1(new_n6921_), .A2(new_n6923_), .A3(new_n6613_), .ZN(new_n6930_));
  AOI21_X1   g06674(.A1(new_n6917_), .A2(new_n6607_), .B(new_n6916_), .ZN(new_n6931_));
  INV_X1     g06675(.I(new_n6928_), .ZN(new_n6932_));
  OAI21_X1   g06676(.A1(new_n6931_), .A2(new_n6930_), .B(new_n6932_), .ZN(new_n6933_));
  NAND2_X1   g06677(.A1(new_n6929_), .A2(new_n6933_), .ZN(new_n6934_));
  AOI21_X1   g06678(.A1(new_n6876_), .A2(new_n6630_), .B(new_n6934_), .ZN(new_n6935_));
  NOR3_X1    g06679(.A1(new_n6557_), .A2(new_n6348_), .A3(new_n6621_), .ZN(new_n6936_));
  NOR3_X1    g06680(.A1(new_n6931_), .A2(new_n6930_), .A3(new_n6932_), .ZN(new_n6937_));
  AOI21_X1   g06681(.A1(new_n6918_), .A2(new_n6924_), .B(new_n6928_), .ZN(new_n6938_));
  NOR2_X1    g06682(.A1(new_n6938_), .A2(new_n6937_), .ZN(new_n6939_));
  NOR3_X1    g06683(.A1(new_n6936_), .A2(new_n6939_), .A3(new_n6625_), .ZN(new_n6940_));
  NOR3_X1    g06684(.A1(new_n6935_), .A2(new_n6940_), .A3(new_n6874_), .ZN(new_n6941_));
  OAI21_X1   g06685(.A1(new_n6936_), .A2(new_n6625_), .B(new_n6939_), .ZN(new_n6942_));
  NAND3_X1   g06686(.A1(new_n6876_), .A2(new_n6630_), .A3(new_n6934_), .ZN(new_n6943_));
  AOI21_X1   g06687(.A1(new_n6943_), .A2(new_n6942_), .B(new_n6873_), .ZN(new_n6944_));
  NOR2_X1    g06688(.A1(new_n6941_), .A2(new_n6944_), .ZN(new_n6945_));
  NAND3_X1   g06689(.A1(new_n6869_), .A2(new_n6945_), .A3(new_n6645_), .ZN(new_n6946_));
  AOI21_X1   g06690(.A1(new_n6554_), .A2(new_n6363_), .B(new_n6638_), .ZN(new_n6947_));
  NAND3_X1   g06691(.A1(new_n6943_), .A2(new_n6942_), .A3(new_n6873_), .ZN(new_n6948_));
  OAI21_X1   g06692(.A1(new_n6935_), .A2(new_n6940_), .B(new_n6874_), .ZN(new_n6949_));
  NAND2_X1   g06693(.A1(new_n6949_), .A2(new_n6948_), .ZN(new_n6950_));
  OAI21_X1   g06694(.A1(new_n6947_), .A2(new_n6641_), .B(new_n6950_), .ZN(new_n6951_));
  NAND3_X1   g06695(.A1(new_n6946_), .A2(new_n6951_), .A3(new_n6866_), .ZN(new_n6952_));
  INV_X1     g06696(.I(new_n6866_), .ZN(new_n6953_));
  NOR3_X1    g06697(.A1(new_n6950_), .A2(new_n6947_), .A3(new_n6641_), .ZN(new_n6954_));
  AOI21_X1   g06698(.A1(new_n6869_), .A2(new_n6645_), .B(new_n6945_), .ZN(new_n6955_));
  OAI21_X1   g06699(.A1(new_n6955_), .A2(new_n6954_), .B(new_n6953_), .ZN(new_n6956_));
  NAND2_X1   g06700(.A1(new_n6952_), .A2(new_n6956_), .ZN(new_n6957_));
  AOI21_X1   g06701(.A1(new_n6661_), .A2(new_n6862_), .B(new_n6957_), .ZN(new_n6958_));
  OAI21_X1   g06702(.A1(new_n6549_), .A2(new_n6651_), .B(new_n6862_), .ZN(new_n6959_));
  INV_X1     g06703(.I(new_n6957_), .ZN(new_n6960_));
  NOR2_X1    g06704(.A1(new_n6959_), .A2(new_n6960_), .ZN(new_n6961_));
  OAI21_X1   g06705(.A1(new_n6961_), .A2(new_n6958_), .B(new_n6860_), .ZN(new_n6962_));
  NAND2_X1   g06706(.A1(new_n6959_), .A2(new_n6960_), .ZN(new_n6963_));
  NAND3_X1   g06707(.A1(new_n6661_), .A2(new_n6862_), .A3(new_n6957_), .ZN(new_n6964_));
  NAND3_X1   g06708(.A1(new_n6963_), .A2(new_n6964_), .A3(new_n6859_), .ZN(new_n6965_));
  NAND2_X1   g06709(.A1(new_n6962_), .A2(new_n6965_), .ZN(new_n6966_));
  AOI21_X1   g06710(.A1(new_n6665_), .A2(new_n6667_), .B(new_n6966_), .ZN(new_n6967_));
  AOI21_X1   g06711(.A1(new_n6963_), .A2(new_n6964_), .B(new_n6859_), .ZN(new_n6968_));
  NOR3_X1    g06712(.A1(new_n6961_), .A2(new_n6958_), .A3(new_n6860_), .ZN(new_n6969_));
  NOR2_X1    g06713(.A1(new_n6969_), .A2(new_n6968_), .ZN(new_n6970_));
  OAI21_X1   g06714(.A1(new_n6380_), .A2(new_n6386_), .B(new_n6390_), .ZN(new_n6971_));
  OAI21_X1   g06715(.A1(new_n6971_), .A2(new_n6669_), .B(new_n6667_), .ZN(new_n6972_));
  NOR2_X1    g06716(.A1(new_n6972_), .A2(new_n6970_), .ZN(new_n6973_));
  NOR3_X1    g06717(.A1(new_n6973_), .A2(new_n6967_), .A3(new_n6855_), .ZN(new_n6974_));
  NAND2_X1   g06718(.A1(new_n6972_), .A2(new_n6970_), .ZN(new_n6975_));
  NAND3_X1   g06719(.A1(new_n6665_), .A2(new_n6667_), .A3(new_n6966_), .ZN(new_n6976_));
  AOI21_X1   g06720(.A1(new_n6975_), .A2(new_n6976_), .B(new_n6854_), .ZN(new_n6977_));
  NOR2_X1    g06721(.A1(new_n6974_), .A2(new_n6977_), .ZN(new_n6978_));
  OAI21_X1   g06722(.A1(new_n6676_), .A2(new_n6850_), .B(new_n6978_), .ZN(new_n6979_));
  INV_X1     g06723(.I(new_n6850_), .ZN(new_n6980_));
  NAND3_X1   g06724(.A1(new_n6975_), .A2(new_n6976_), .A3(new_n6854_), .ZN(new_n6981_));
  OAI21_X1   g06725(.A1(new_n6973_), .A2(new_n6967_), .B(new_n6855_), .ZN(new_n6982_));
  NAND2_X1   g06726(.A1(new_n6982_), .A2(new_n6981_), .ZN(new_n6983_));
  NAND3_X1   g06727(.A1(new_n6683_), .A2(new_n6983_), .A3(new_n6980_), .ZN(new_n6984_));
  NAND3_X1   g06728(.A1(new_n6979_), .A2(new_n6984_), .A3(new_n6849_), .ZN(new_n6985_));
  INV_X1     g06729(.I(new_n6849_), .ZN(new_n6986_));
  AOI21_X1   g06730(.A1(new_n6683_), .A2(new_n6980_), .B(new_n6983_), .ZN(new_n6987_));
  OAI21_X1   g06731(.A1(new_n6684_), .A2(new_n6675_), .B(new_n6980_), .ZN(new_n6988_));
  NOR2_X1    g06732(.A1(new_n6988_), .A2(new_n6978_), .ZN(new_n6989_));
  OAI21_X1   g06733(.A1(new_n6989_), .A2(new_n6987_), .B(new_n6986_), .ZN(new_n6990_));
  NAND2_X1   g06734(.A1(new_n6990_), .A2(new_n6985_), .ZN(new_n6991_));
  AOI21_X1   g06735(.A1(new_n6688_), .A2(new_n6690_), .B(new_n6991_), .ZN(new_n6992_));
  OAI21_X1   g06736(.A1(new_n6689_), .A2(new_n6692_), .B(new_n6690_), .ZN(new_n6993_));
  NOR3_X1    g06737(.A1(new_n6989_), .A2(new_n6987_), .A3(new_n6986_), .ZN(new_n6994_));
  AOI21_X1   g06738(.A1(new_n6979_), .A2(new_n6984_), .B(new_n6849_), .ZN(new_n6995_));
  NOR2_X1    g06739(.A1(new_n6994_), .A2(new_n6995_), .ZN(new_n6996_));
  NOR2_X1    g06740(.A1(new_n6993_), .A2(new_n6996_), .ZN(new_n6997_));
  NOR3_X1    g06741(.A1(new_n6997_), .A2(new_n6845_), .A3(new_n6992_), .ZN(new_n6998_));
  OAI21_X1   g06742(.A1(new_n6696_), .A2(new_n6682_), .B(new_n6996_), .ZN(new_n6999_));
  NAND3_X1   g06743(.A1(new_n6688_), .A2(new_n6991_), .A3(new_n6690_), .ZN(new_n7000_));
  AOI21_X1   g06744(.A1(new_n6999_), .A2(new_n7000_), .B(new_n6844_), .ZN(new_n7001_));
  NOR2_X1    g06745(.A1(new_n6998_), .A2(new_n7001_), .ZN(new_n7002_));
  OAI21_X1   g06746(.A1(new_n6715_), .A2(new_n6840_), .B(new_n7002_), .ZN(new_n7003_));
  INV_X1     g06747(.I(new_n6840_), .ZN(new_n7004_));
  NAND3_X1   g06748(.A1(new_n6999_), .A2(new_n7000_), .A3(new_n6844_), .ZN(new_n7005_));
  OAI21_X1   g06749(.A1(new_n6997_), .A2(new_n6992_), .B(new_n6845_), .ZN(new_n7006_));
  NAND2_X1   g06750(.A1(new_n7006_), .A2(new_n7005_), .ZN(new_n7007_));
  NAND3_X1   g06751(.A1(new_n6706_), .A2(new_n7007_), .A3(new_n7004_), .ZN(new_n7008_));
  NAND3_X1   g06752(.A1(new_n7003_), .A2(new_n7008_), .A3(new_n6839_), .ZN(new_n7009_));
  XOR2_X1    g06753(.A1(new_n6838_), .A2(new_n1002_), .Z(new_n7010_));
  AOI21_X1   g06754(.A1(new_n6706_), .A2(new_n7004_), .B(new_n7007_), .ZN(new_n7011_));
  OAI21_X1   g06755(.A1(new_n6525_), .A2(new_n6700_), .B(new_n7004_), .ZN(new_n7012_));
  NOR2_X1    g06756(.A1(new_n7012_), .A2(new_n7002_), .ZN(new_n7013_));
  OAI21_X1   g06757(.A1(new_n7013_), .A2(new_n7011_), .B(new_n7010_), .ZN(new_n7014_));
  NAND2_X1   g06758(.A1(new_n7014_), .A2(new_n7009_), .ZN(new_n7015_));
  NOR3_X1    g06759(.A1(new_n6835_), .A2(new_n7015_), .A3(new_n6725_), .ZN(new_n7016_));
  OAI21_X1   g06760(.A1(new_n6723_), .A2(new_n6442_), .B(new_n6711_), .ZN(new_n7017_));
  NOR3_X1    g06761(.A1(new_n7013_), .A2(new_n7011_), .A3(new_n7010_), .ZN(new_n7018_));
  AOI21_X1   g06762(.A1(new_n7003_), .A2(new_n7008_), .B(new_n6839_), .ZN(new_n7019_));
  NOR2_X1    g06763(.A1(new_n7018_), .A2(new_n7019_), .ZN(new_n7020_));
  AOI21_X1   g06764(.A1(new_n7017_), .A2(new_n6717_), .B(new_n7020_), .ZN(new_n7021_));
  OAI21_X1   g06765(.A1(new_n7021_), .A2(new_n7016_), .B(new_n6834_), .ZN(new_n7022_));
  INV_X1     g06766(.I(new_n6833_), .ZN(new_n7023_));
  NOR2_X1    g06767(.A1(new_n7023_), .A2(new_n6831_), .ZN(new_n7024_));
  NAND3_X1   g06768(.A1(new_n7017_), .A2(new_n6717_), .A3(new_n7020_), .ZN(new_n7025_));
  OAI21_X1   g06769(.A1(new_n6835_), .A2(new_n6725_), .B(new_n7015_), .ZN(new_n7026_));
  NAND3_X1   g06770(.A1(new_n7025_), .A2(new_n7026_), .A3(new_n7024_), .ZN(new_n7027_));
  NAND2_X1   g06771(.A1(new_n7022_), .A2(new_n7027_), .ZN(new_n7028_));
  AOI21_X1   g06772(.A1(new_n6729_), .A2(new_n6730_), .B(new_n6521_), .ZN(new_n7029_));
  OAI21_X1   g06773(.A1(new_n6013_), .A2(new_n6010_), .B(new_n6014_), .ZN(new_n7030_));
  OAI21_X1   g06774(.A1(new_n7030_), .A2(new_n6262_), .B(new_n6260_), .ZN(new_n7031_));
  AOI21_X1   g06775(.A1(new_n7031_), .A2(new_n6455_), .B(new_n6450_), .ZN(new_n7032_));
  NOR3_X1    g06776(.A1(new_n7032_), .A2(new_n6732_), .A3(new_n6515_), .ZN(new_n7033_));
  OAI21_X1   g06777(.A1(new_n7033_), .A2(new_n7029_), .B(new_n7028_), .ZN(new_n7034_));
  AOI21_X1   g06778(.A1(new_n7025_), .A2(new_n7026_), .B(new_n7024_), .ZN(new_n7035_));
  NOR3_X1    g06779(.A1(new_n7021_), .A2(new_n6834_), .A3(new_n7016_), .ZN(new_n7036_));
  NOR2_X1    g06780(.A1(new_n7036_), .A2(new_n7035_), .ZN(new_n7037_));
  INV_X1     g06781(.I(new_n7029_), .ZN(new_n7038_));
  AOI21_X1   g06782(.A1(new_n5807_), .A2(new_n6009_), .B(new_n6008_), .ZN(new_n7039_));
  AOI21_X1   g06783(.A1(new_n7039_), .A2(new_n6255_), .B(new_n6250_), .ZN(new_n7040_));
  OAI21_X1   g06784(.A1(new_n7040_), .A2(new_n6457_), .B(new_n6463_), .ZN(new_n7041_));
  NAND3_X1   g06785(.A1(new_n7041_), .A2(new_n6458_), .A3(new_n6738_), .ZN(new_n7042_));
  NAND3_X1   g06786(.A1(new_n7042_), .A2(new_n7037_), .A3(new_n7038_), .ZN(new_n7043_));
  AOI22_X1   g06787(.A1(new_n518_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n636_), .ZN(new_n7044_));
  OAI21_X1   g06788(.A1(new_n4886_), .A2(new_n917_), .B(new_n7044_), .ZN(new_n7045_));
  AOI21_X1   g06789(.A1(new_n5351_), .A2(new_n618_), .B(new_n7045_), .ZN(new_n7046_));
  XOR2_X1    g06790(.A1(new_n7046_), .A2(\a[8] ), .Z(new_n7047_));
  NAND3_X1   g06791(.A1(new_n7043_), .A2(new_n7034_), .A3(new_n7047_), .ZN(new_n7048_));
  AOI21_X1   g06792(.A1(new_n7042_), .A2(new_n7038_), .B(new_n7037_), .ZN(new_n7049_));
  NOR3_X1    g06793(.A1(new_n7033_), .A2(new_n7028_), .A3(new_n7029_), .ZN(new_n7050_));
  INV_X1     g06794(.I(new_n7047_), .ZN(new_n7051_));
  OAI21_X1   g06795(.A1(new_n7049_), .A2(new_n7050_), .B(new_n7051_), .ZN(new_n7052_));
  NAND2_X1   g06796(.A1(new_n7052_), .A2(new_n7048_), .ZN(new_n7053_));
  AOI21_X1   g06797(.A1(new_n6733_), .A2(new_n6739_), .B(new_n6765_), .ZN(new_n7054_));
  INV_X1     g06798(.I(new_n7054_), .ZN(new_n7055_));
  NAND3_X1   g06799(.A1(new_n6765_), .A2(new_n6733_), .A3(new_n6739_), .ZN(new_n7056_));
  INV_X1     g06800(.I(new_n7056_), .ZN(new_n7057_));
  OAI21_X1   g06801(.A1(new_n6746_), .A2(new_n7057_), .B(new_n7055_), .ZN(new_n7058_));
  NAND2_X1   g06802(.A1(new_n7058_), .A2(new_n7053_), .ZN(new_n7059_));
  NOR3_X1    g06803(.A1(new_n7049_), .A2(new_n7050_), .A3(new_n7051_), .ZN(new_n7060_));
  AOI21_X1   g06804(.A1(new_n7043_), .A2(new_n7034_), .B(new_n7047_), .ZN(new_n7061_));
  NOR2_X1    g06805(.A1(new_n7060_), .A2(new_n7061_), .ZN(new_n7062_));
  NAND3_X1   g06806(.A1(new_n6759_), .A2(new_n6473_), .A3(new_n7056_), .ZN(new_n7063_));
  NAND3_X1   g06807(.A1(new_n7063_), .A2(new_n7062_), .A3(new_n7055_), .ZN(new_n7064_));
  NAND3_X1   g06808(.A1(new_n7059_), .A2(new_n6826_), .A3(new_n7064_), .ZN(new_n7065_));
  INV_X1     g06809(.I(new_n6823_), .ZN(new_n7066_));
  NAND2_X1   g06810(.A1(new_n7066_), .A2(new_n6824_), .ZN(new_n7067_));
  AOI21_X1   g06811(.A1(new_n6815_), .A2(new_n7056_), .B(new_n7054_), .ZN(new_n7068_));
  NOR2_X1    g06812(.A1(new_n7068_), .A2(new_n7062_), .ZN(new_n7069_));
  NOR2_X1    g06813(.A1(new_n7058_), .A2(new_n7053_), .ZN(new_n7070_));
  OAI21_X1   g06814(.A1(new_n7069_), .A2(new_n7070_), .B(new_n7067_), .ZN(new_n7071_));
  NAND2_X1   g06815(.A1(new_n7071_), .A2(new_n7065_), .ZN(new_n7072_));
  XOR2_X1    g06816(.A1(new_n7072_), .A2(new_n6818_), .Z(new_n7073_));
  INV_X1     g06817(.I(\b[44] ), .ZN(new_n7074_));
  OAI22_X1   g06818(.A1(new_n277_), .A2(new_n7074_), .B1(new_n6775_), .B2(new_n262_), .ZN(new_n7075_));
  AOI21_X1   g06819(.A1(\b[42] ), .A2(new_n283_), .B(new_n7075_), .ZN(new_n7076_));
  XOR2_X1    g06820(.A1(\b[43] ), .A2(\b[44] ), .Z(new_n7077_));
  OAI21_X1   g06821(.A1(new_n6779_), .A2(\b[42] ), .B(\b[43] ), .ZN(new_n7078_));
  OAI21_X1   g06822(.A1(new_n6494_), .A2(\b[41] ), .B(\b[42] ), .ZN(new_n7079_));
  NAND2_X1   g06823(.A1(new_n7078_), .A2(new_n7079_), .ZN(new_n7080_));
  XNOR2_X1   g06824(.A1(new_n7080_), .A2(new_n7077_), .ZN(new_n7081_));
  OAI21_X1   g06825(.A1(new_n7081_), .A2(new_n279_), .B(new_n7076_), .ZN(new_n7082_));
  XOR2_X1    g06826(.A1(new_n7082_), .A2(\a[2] ), .Z(new_n7083_));
  NOR2_X1    g06827(.A1(new_n7073_), .A2(new_n7083_), .ZN(new_n7084_));
  NAND2_X1   g06828(.A1(new_n7073_), .A2(new_n7083_), .ZN(new_n7085_));
  INV_X1     g06829(.I(new_n7085_), .ZN(new_n7086_));
  NOR2_X1    g06830(.A1(new_n7086_), .A2(new_n7084_), .ZN(new_n7087_));
  XOR2_X1    g06831(.A1(new_n6813_), .A2(new_n7087_), .Z(\f[44] ));
  INV_X1     g06832(.I(new_n7084_), .ZN(new_n7089_));
  OAI21_X1   g06833(.A1(new_n6812_), .A2(new_n6811_), .B(new_n7085_), .ZN(new_n7090_));
  NAND2_X1   g06834(.A1(new_n7090_), .A2(new_n7089_), .ZN(new_n7091_));
  NAND2_X1   g06835(.A1(new_n283_), .A2(\b[43] ), .ZN(new_n7092_));
  AOI22_X1   g06836(.A1(new_n267_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n261_), .ZN(new_n7093_));
  AOI21_X1   g06837(.A1(new_n7080_), .A2(\b[44] ), .B(new_n6775_), .ZN(new_n7094_));
  NOR2_X1    g06838(.A1(new_n7080_), .A2(\b[44] ), .ZN(new_n7095_));
  INV_X1     g06839(.I(\b[45] ), .ZN(new_n7096_));
  NAND3_X1   g06840(.A1(new_n7078_), .A2(new_n7079_), .A3(new_n7096_), .ZN(new_n7097_));
  INV_X1     g06841(.I(new_n7097_), .ZN(new_n7098_));
  AOI21_X1   g06842(.A1(new_n7078_), .A2(new_n7079_), .B(new_n7096_), .ZN(new_n7099_));
  OAI22_X1   g06843(.A1(new_n7094_), .A2(new_n7095_), .B1(new_n7098_), .B2(new_n7099_), .ZN(new_n7100_));
  OR4_X2     g06844(.A1(new_n7094_), .A2(new_n7095_), .A3(new_n7098_), .A4(new_n7099_), .Z(new_n7101_));
  NAND3_X1   g06845(.A1(new_n7101_), .A2(new_n265_), .A3(new_n7100_), .ZN(new_n7102_));
  NAND3_X1   g06846(.A1(new_n7102_), .A2(new_n7092_), .A3(new_n7093_), .ZN(new_n7103_));
  XOR2_X1    g06847(.A1(new_n7103_), .A2(new_n270_), .Z(new_n7104_));
  INV_X1     g06848(.I(new_n7104_), .ZN(new_n7105_));
  NAND2_X1   g06849(.A1(new_n6497_), .A2(new_n6493_), .ZN(new_n7106_));
  AOI22_X1   g06850(.A1(new_n800_), .A2(\b[41] ), .B1(\b[42] ), .B2(new_n333_), .ZN(new_n7107_));
  OAI21_X1   g06851(.A1(new_n6284_), .A2(new_n392_), .B(new_n7107_), .ZN(new_n7108_));
  AOI21_X1   g06852(.A1(new_n7106_), .A2(new_n330_), .B(new_n7108_), .ZN(new_n7109_));
  XOR2_X1    g06853(.A1(new_n7109_), .A2(new_n312_), .Z(new_n7110_));
  NAND2_X1   g06854(.A1(new_n6887_), .A2(\b[1] ), .ZN(new_n7111_));
  AOI22_X1   g06855(.A1(new_n6569_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n6574_), .ZN(new_n7112_));
  NAND2_X1   g06856(.A1(new_n299_), .A2(new_n6579_), .ZN(new_n7113_));
  NAND3_X1   g06857(.A1(new_n7113_), .A2(new_n7112_), .A3(new_n7111_), .ZN(new_n7114_));
  XOR2_X1    g06858(.A1(new_n7114_), .A2(new_n6567_), .Z(new_n7115_));
  XNOR2_X1   g06859(.A1(\a[44] ), .A2(\a[45] ), .ZN(new_n7116_));
  NOR2_X1    g06860(.A1(new_n7116_), .A2(new_n258_), .ZN(new_n7117_));
  INV_X1     g06861(.I(new_n7117_), .ZN(new_n7118_));
  NAND2_X1   g06862(.A1(new_n7115_), .A2(new_n7118_), .ZN(new_n7119_));
  XOR2_X1    g06863(.A1(new_n7114_), .A2(\a[44] ), .Z(new_n7120_));
  NAND2_X1   g06864(.A1(new_n7120_), .A2(new_n7117_), .ZN(new_n7121_));
  NAND2_X1   g06865(.A1(new_n7119_), .A2(new_n7121_), .ZN(new_n7122_));
  XOR2_X1    g06866(.A1(new_n7122_), .A2(new_n6894_), .Z(new_n7123_));
  OAI22_X1   g06867(.A1(new_n5852_), .A2(new_n438_), .B1(new_n377_), .B2(new_n5857_), .ZN(new_n7124_));
  AOI21_X1   g06868(.A1(\b[4] ), .A2(new_n6115_), .B(new_n7124_), .ZN(new_n7125_));
  OAI21_X1   g06869(.A1(new_n450_), .A2(new_n5861_), .B(new_n7125_), .ZN(new_n7126_));
  XOR2_X1    g06870(.A1(new_n7126_), .A2(\a[41] ), .Z(new_n7127_));
  OAI21_X1   g06871(.A1(new_n6904_), .A2(new_n6899_), .B(new_n6908_), .ZN(new_n7128_));
  NAND2_X1   g06872(.A1(new_n7128_), .A2(new_n7127_), .ZN(new_n7129_));
  NOR2_X1    g06873(.A1(new_n7128_), .A2(new_n7127_), .ZN(new_n7130_));
  INV_X1     g06874(.I(new_n7130_), .ZN(new_n7131_));
  NAND2_X1   g06875(.A1(new_n7131_), .A2(new_n7129_), .ZN(new_n7132_));
  XNOR2_X1   g06876(.A1(new_n7132_), .A2(new_n7123_), .ZN(new_n7133_));
  AOI22_X1   g06877(.A1(new_n5155_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n5160_), .ZN(new_n7134_));
  OAI21_X1   g06878(.A1(new_n471_), .A2(new_n6877_), .B(new_n7134_), .ZN(new_n7135_));
  AOI21_X1   g06879(.A1(new_n676_), .A2(new_n5166_), .B(new_n7135_), .ZN(new_n7136_));
  XOR2_X1    g06880(.A1(new_n7136_), .A2(new_n5162_), .Z(new_n7137_));
  INV_X1     g06881(.I(new_n7137_), .ZN(new_n7138_));
  AOI21_X1   g06882(.A1(new_n6918_), .A2(new_n6920_), .B(new_n7138_), .ZN(new_n7139_));
  NOR3_X1    g06883(.A1(new_n6930_), .A2(new_n6915_), .A3(new_n7137_), .ZN(new_n7140_));
  NOR3_X1    g06884(.A1(new_n7139_), .A2(new_n7133_), .A3(new_n7140_), .ZN(new_n7141_));
  XOR2_X1    g06885(.A1(new_n7132_), .A2(new_n7123_), .Z(new_n7142_));
  OAI21_X1   g06886(.A1(new_n6930_), .A2(new_n6915_), .B(new_n7137_), .ZN(new_n7143_));
  NAND3_X1   g06887(.A1(new_n6918_), .A2(new_n6920_), .A3(new_n7138_), .ZN(new_n7144_));
  AOI21_X1   g06888(.A1(new_n7144_), .A2(new_n7143_), .B(new_n7142_), .ZN(new_n7145_));
  NOR2_X1    g06889(.A1(new_n7141_), .A2(new_n7145_), .ZN(new_n7146_));
  AOI22_X1   g06890(.A1(new_n4918_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n4921_), .ZN(new_n7147_));
  OAI21_X1   g06891(.A1(new_n776_), .A2(new_n6099_), .B(new_n7147_), .ZN(new_n7148_));
  AOI21_X1   g06892(.A1(new_n1194_), .A2(new_n4699_), .B(new_n7148_), .ZN(new_n7149_));
  XOR2_X1    g06893(.A1(new_n7149_), .A2(new_n4446_), .Z(new_n7150_));
  OAI21_X1   g06894(.A1(new_n6935_), .A2(new_n6937_), .B(new_n7150_), .ZN(new_n7151_));
  INV_X1     g06895(.I(new_n7150_), .ZN(new_n7152_));
  NAND3_X1   g06896(.A1(new_n6942_), .A2(new_n6929_), .A3(new_n7152_), .ZN(new_n7153_));
  NAND2_X1   g06897(.A1(new_n7151_), .A2(new_n7153_), .ZN(new_n7154_));
  XOR2_X1    g06898(.A1(new_n7154_), .A2(new_n7146_), .Z(new_n7155_));
  OAI22_X1   g06899(.A1(new_n1093_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n1268_), .ZN(new_n7156_));
  AOI21_X1   g06900(.A1(\b[13] ), .A2(new_n4053_), .B(new_n7156_), .ZN(new_n7157_));
  OAI21_X1   g06901(.A1(new_n1275_), .A2(new_n4727_), .B(new_n7157_), .ZN(new_n7158_));
  XOR2_X1    g06902(.A1(new_n7158_), .A2(\a[32] ), .Z(new_n7159_));
  INV_X1     g06903(.I(new_n7159_), .ZN(new_n7160_));
  AOI21_X1   g06904(.A1(new_n6946_), .A2(new_n6948_), .B(new_n7160_), .ZN(new_n7161_));
  NOR3_X1    g06905(.A1(new_n6954_), .A2(new_n6941_), .A3(new_n7159_), .ZN(new_n7162_));
  NOR3_X1    g06906(.A1(new_n7161_), .A2(new_n7162_), .A3(new_n7155_), .ZN(new_n7163_));
  INV_X1     g06907(.I(new_n7146_), .ZN(new_n7164_));
  NOR2_X1    g06908(.A1(new_n7154_), .A2(new_n7164_), .ZN(new_n7165_));
  AOI21_X1   g06909(.A1(new_n7151_), .A2(new_n7153_), .B(new_n7146_), .ZN(new_n7166_));
  NOR2_X1    g06910(.A1(new_n7165_), .A2(new_n7166_), .ZN(new_n7167_));
  OAI21_X1   g06911(.A1(new_n6954_), .A2(new_n6941_), .B(new_n7159_), .ZN(new_n7168_));
  NAND3_X1   g06912(.A1(new_n6946_), .A2(new_n6948_), .A3(new_n7160_), .ZN(new_n7169_));
  AOI21_X1   g06913(.A1(new_n7169_), .A2(new_n7168_), .B(new_n7167_), .ZN(new_n7170_));
  NOR2_X1    g06914(.A1(new_n7163_), .A2(new_n7170_), .ZN(new_n7171_));
  INV_X1     g06915(.I(new_n6952_), .ZN(new_n7172_));
  AOI22_X1   g06916(.A1(new_n3267_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n3270_), .ZN(new_n7173_));
  OAI21_X1   g06917(.A1(new_n1296_), .A2(new_n3475_), .B(new_n7173_), .ZN(new_n7174_));
  AOI21_X1   g06918(.A1(new_n2038_), .A2(new_n3273_), .B(new_n7174_), .ZN(new_n7175_));
  XOR2_X1    g06919(.A1(new_n7175_), .A2(new_n3264_), .Z(new_n7176_));
  OAI21_X1   g06920(.A1(new_n6958_), .A2(new_n7172_), .B(new_n7176_), .ZN(new_n7177_));
  INV_X1     g06921(.I(new_n7176_), .ZN(new_n7178_));
  AOI21_X1   g06922(.A1(new_n6959_), .A2(new_n6956_), .B(new_n7172_), .ZN(new_n7179_));
  NAND2_X1   g06923(.A1(new_n7179_), .A2(new_n7178_), .ZN(new_n7180_));
  NAND3_X1   g06924(.A1(new_n7180_), .A2(new_n7177_), .A3(new_n7171_), .ZN(new_n7181_));
  INV_X1     g06925(.I(new_n7181_), .ZN(new_n7182_));
  AOI21_X1   g06926(.A1(new_n7180_), .A2(new_n7177_), .B(new_n7171_), .ZN(new_n7183_));
  NOR2_X1    g06927(.A1(new_n7182_), .A2(new_n7183_), .ZN(new_n7184_));
  AOI22_X1   g06928(.A1(new_n2716_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n2719_), .ZN(new_n7185_));
  OAI21_X1   g06929(.A1(new_n1859_), .A2(new_n2924_), .B(new_n7185_), .ZN(new_n7186_));
  AOI21_X1   g06930(.A1(new_n2032_), .A2(new_n2722_), .B(new_n7186_), .ZN(new_n7187_));
  XOR2_X1    g06931(.A1(new_n7187_), .A2(new_n2714_), .Z(new_n7188_));
  OAI21_X1   g06932(.A1(new_n6967_), .A2(new_n6969_), .B(new_n7188_), .ZN(new_n7189_));
  INV_X1     g06933(.I(new_n7188_), .ZN(new_n7190_));
  AOI21_X1   g06934(.A1(new_n6972_), .A2(new_n6970_), .B(new_n6969_), .ZN(new_n7191_));
  NAND2_X1   g06935(.A1(new_n7191_), .A2(new_n7190_), .ZN(new_n7192_));
  NAND3_X1   g06936(.A1(new_n7192_), .A2(new_n7189_), .A3(new_n7184_), .ZN(new_n7193_));
  INV_X1     g06937(.I(new_n7171_), .ZN(new_n7194_));
  NAND2_X1   g06938(.A1(new_n7180_), .A2(new_n7177_), .ZN(new_n7195_));
  NAND2_X1   g06939(.A1(new_n7195_), .A2(new_n7194_), .ZN(new_n7196_));
  NAND2_X1   g06940(.A1(new_n7196_), .A2(new_n7181_), .ZN(new_n7197_));
  INV_X1     g06941(.I(new_n7189_), .ZN(new_n7198_));
  NOR3_X1    g06942(.A1(new_n6967_), .A2(new_n6969_), .A3(new_n7188_), .ZN(new_n7199_));
  OAI21_X1   g06943(.A1(new_n7198_), .A2(new_n7199_), .B(new_n7197_), .ZN(new_n7200_));
  NAND2_X1   g06944(.A1(new_n7200_), .A2(new_n7193_), .ZN(new_n7201_));
  AOI22_X1   g06945(.A1(new_n2202_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n2205_), .ZN(new_n7202_));
  OAI21_X1   g06946(.A1(new_n2142_), .A2(new_n2370_), .B(new_n7202_), .ZN(new_n7203_));
  AOI21_X1   g06947(.A1(new_n3033_), .A2(new_n2208_), .B(new_n7203_), .ZN(new_n7204_));
  XOR2_X1    g06948(.A1(new_n7204_), .A2(new_n2200_), .Z(new_n7205_));
  INV_X1     g06949(.I(new_n7205_), .ZN(new_n7206_));
  AOI21_X1   g06950(.A1(new_n6988_), .A2(new_n6978_), .B(new_n6974_), .ZN(new_n7207_));
  NOR2_X1    g06951(.A1(new_n7207_), .A2(new_n7206_), .ZN(new_n7208_));
  NOR3_X1    g06952(.A1(new_n6987_), .A2(new_n6974_), .A3(new_n7205_), .ZN(new_n7209_));
  NOR3_X1    g06953(.A1(new_n7208_), .A2(new_n7209_), .A3(new_n7201_), .ZN(new_n7210_));
  NOR3_X1    g06954(.A1(new_n7198_), .A2(new_n7199_), .A3(new_n7197_), .ZN(new_n7211_));
  AOI21_X1   g06955(.A1(new_n7192_), .A2(new_n7189_), .B(new_n7184_), .ZN(new_n7212_));
  NOR2_X1    g06956(.A1(new_n7211_), .A2(new_n7212_), .ZN(new_n7213_));
  AOI21_X1   g06957(.A1(new_n6392_), .A2(new_n6402_), .B(new_n6400_), .ZN(new_n7214_));
  AOI21_X1   g06958(.A1(new_n7214_), .A2(new_n6680_), .B(new_n6850_), .ZN(new_n7215_));
  OAI21_X1   g06959(.A1(new_n7215_), .A2(new_n6983_), .B(new_n6981_), .ZN(new_n7216_));
  NAND2_X1   g06960(.A1(new_n7216_), .A2(new_n7205_), .ZN(new_n7217_));
  NAND3_X1   g06961(.A1(new_n6979_), .A2(new_n6981_), .A3(new_n7206_), .ZN(new_n7218_));
  AOI21_X1   g06962(.A1(new_n7217_), .A2(new_n7218_), .B(new_n7213_), .ZN(new_n7219_));
  NOR2_X1    g06963(.A1(new_n7210_), .A2(new_n7219_), .ZN(new_n7220_));
  OAI22_X1   g06964(.A1(new_n1751_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n1754_), .ZN(new_n7221_));
  AOI21_X1   g06965(.A1(\b[25] ), .A2(new_n1939_), .B(new_n7221_), .ZN(new_n7222_));
  OAI21_X1   g06966(.A1(new_n3165_), .A2(new_n1757_), .B(new_n7222_), .ZN(new_n7223_));
  XOR2_X1    g06967(.A1(new_n7223_), .A2(\a[20] ), .Z(new_n7224_));
  OAI21_X1   g06968(.A1(new_n6992_), .A2(new_n6994_), .B(new_n7224_), .ZN(new_n7225_));
  INV_X1     g06969(.I(new_n7224_), .ZN(new_n7226_));
  NAND3_X1   g06970(.A1(new_n6999_), .A2(new_n6985_), .A3(new_n7226_), .ZN(new_n7227_));
  NAND3_X1   g06971(.A1(new_n7227_), .A2(new_n7225_), .A3(new_n7220_), .ZN(new_n7228_));
  INV_X1     g06972(.I(new_n7228_), .ZN(new_n7229_));
  AOI21_X1   g06973(.A1(new_n7227_), .A2(new_n7225_), .B(new_n7220_), .ZN(new_n7230_));
  NOR2_X1    g06974(.A1(new_n7229_), .A2(new_n7230_), .ZN(new_n7231_));
  OAI22_X1   g06975(.A1(new_n1592_), .A2(new_n3624_), .B1(new_n3592_), .B2(new_n1505_), .ZN(new_n7232_));
  AOI21_X1   g06976(.A1(\b[28] ), .A2(new_n1584_), .B(new_n7232_), .ZN(new_n7233_));
  OAI21_X1   g06977(.A1(new_n3634_), .A2(new_n1732_), .B(new_n7233_), .ZN(new_n7234_));
  XOR2_X1    g06978(.A1(new_n7234_), .A2(\a[17] ), .Z(new_n7235_));
  OAI21_X1   g06979(.A1(new_n7011_), .A2(new_n6998_), .B(new_n7235_), .ZN(new_n7236_));
  INV_X1     g06980(.I(new_n7235_), .ZN(new_n7237_));
  NAND3_X1   g06981(.A1(new_n7003_), .A2(new_n7005_), .A3(new_n7237_), .ZN(new_n7238_));
  NAND3_X1   g06982(.A1(new_n7238_), .A2(new_n7236_), .A3(new_n7231_), .ZN(new_n7239_));
  AOI21_X1   g06983(.A1(new_n7238_), .A2(new_n7236_), .B(new_n7231_), .ZN(new_n7240_));
  INV_X1     g06984(.I(new_n7240_), .ZN(new_n7241_));
  NAND2_X1   g06985(.A1(new_n7241_), .A2(new_n7239_), .ZN(new_n7242_));
  OAI22_X1   g06986(.A1(new_n993_), .A2(new_n4638_), .B1(new_n4023_), .B2(new_n997_), .ZN(new_n7243_));
  AOI21_X1   g06987(.A1(\b[31] ), .A2(new_n1486_), .B(new_n7243_), .ZN(new_n7244_));
  OAI21_X1   g06988(.A1(new_n6451_), .A2(new_n1323_), .B(new_n7244_), .ZN(new_n7245_));
  XOR2_X1    g06989(.A1(new_n7245_), .A2(\a[14] ), .Z(new_n7246_));
  INV_X1     g06990(.I(new_n7246_), .ZN(new_n7247_));
  AOI21_X1   g06991(.A1(new_n7025_), .A2(new_n7009_), .B(new_n7247_), .ZN(new_n7248_));
  NOR3_X1    g06992(.A1(new_n7016_), .A2(new_n7018_), .A3(new_n7246_), .ZN(new_n7249_));
  NOR3_X1    g06993(.A1(new_n7248_), .A2(new_n7249_), .A3(new_n7242_), .ZN(new_n7250_));
  INV_X1     g06994(.I(new_n7239_), .ZN(new_n7251_));
  NOR2_X1    g06995(.A1(new_n7251_), .A2(new_n7240_), .ZN(new_n7252_));
  OAI21_X1   g06996(.A1(new_n7016_), .A2(new_n7018_), .B(new_n7246_), .ZN(new_n7253_));
  NAND3_X1   g06997(.A1(new_n7025_), .A2(new_n7009_), .A3(new_n7247_), .ZN(new_n7254_));
  AOI21_X1   g06998(.A1(new_n7254_), .A2(new_n7253_), .B(new_n7252_), .ZN(new_n7255_));
  NOR2_X1    g06999(.A1(new_n7250_), .A2(new_n7255_), .ZN(new_n7256_));
  INV_X1     g07000(.I(new_n7256_), .ZN(new_n7257_));
  OAI22_X1   g07001(.A1(new_n713_), .A2(new_n4886_), .B1(new_n4666_), .B2(new_n717_), .ZN(new_n7258_));
  AOI21_X1   g07002(.A1(\b[34] ), .A2(new_n1126_), .B(new_n7258_), .ZN(new_n7259_));
  OAI21_X1   g07003(.A1(new_n4898_), .A2(new_n986_), .B(new_n7259_), .ZN(new_n7260_));
  XOR2_X1    g07004(.A1(new_n7260_), .A2(\a[11] ), .Z(new_n7261_));
  INV_X1     g07005(.I(new_n7261_), .ZN(new_n7262_));
  OAI21_X1   g07006(.A1(new_n7033_), .A2(new_n7029_), .B(new_n7037_), .ZN(new_n7263_));
  AOI21_X1   g07007(.A1(new_n7263_), .A2(new_n7027_), .B(new_n7262_), .ZN(new_n7264_));
  AOI21_X1   g07008(.A1(new_n7042_), .A2(new_n7038_), .B(new_n7028_), .ZN(new_n7265_));
  NOR3_X1    g07009(.A1(new_n7265_), .A2(new_n7036_), .A3(new_n7261_), .ZN(new_n7266_));
  NOR3_X1    g07010(.A1(new_n7266_), .A2(new_n7264_), .A3(new_n7257_), .ZN(new_n7267_));
  OAI21_X1   g07011(.A1(new_n7265_), .A2(new_n7036_), .B(new_n7261_), .ZN(new_n7268_));
  NAND3_X1   g07012(.A1(new_n7263_), .A2(new_n7027_), .A3(new_n7262_), .ZN(new_n7269_));
  AOI21_X1   g07013(.A1(new_n7268_), .A2(new_n7269_), .B(new_n7256_), .ZN(new_n7270_));
  OR2_X2     g07014(.A1(new_n7267_), .A2(new_n7270_), .Z(new_n7271_));
  AOI22_X1   g07015(.A1(new_n518_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n636_), .ZN(new_n7272_));
  OAI21_X1   g07016(.A1(new_n5312_), .A2(new_n917_), .B(new_n7272_), .ZN(new_n7273_));
  AOI21_X1   g07017(.A1(new_n6310_), .A2(new_n618_), .B(new_n7273_), .ZN(new_n7274_));
  XOR2_X1    g07018(.A1(new_n7274_), .A2(new_n488_), .Z(new_n7275_));
  INV_X1     g07019(.I(new_n7275_), .ZN(new_n7276_));
  NOR3_X1    g07020(.A1(new_n6769_), .A2(new_n6477_), .A3(new_n7057_), .ZN(new_n7277_));
  OAI21_X1   g07021(.A1(new_n7277_), .A2(new_n7054_), .B(new_n7062_), .ZN(new_n7278_));
  AOI21_X1   g07022(.A1(new_n7278_), .A2(new_n7052_), .B(new_n7276_), .ZN(new_n7279_));
  AOI21_X1   g07023(.A1(new_n7063_), .A2(new_n7055_), .B(new_n7053_), .ZN(new_n7280_));
  NOR3_X1    g07024(.A1(new_n7280_), .A2(new_n7061_), .A3(new_n7275_), .ZN(new_n7281_));
  NOR3_X1    g07025(.A1(new_n7279_), .A2(new_n7281_), .A3(new_n7271_), .ZN(new_n7282_));
  NOR2_X1    g07026(.A1(new_n7267_), .A2(new_n7270_), .ZN(new_n7283_));
  OAI21_X1   g07027(.A1(new_n7280_), .A2(new_n7061_), .B(new_n7275_), .ZN(new_n7284_));
  NAND3_X1   g07028(.A1(new_n7278_), .A2(new_n7052_), .A3(new_n7276_), .ZN(new_n7285_));
  AOI21_X1   g07029(.A1(new_n7285_), .A2(new_n7284_), .B(new_n7283_), .ZN(new_n7286_));
  NOR3_X1    g07030(.A1(new_n7282_), .A2(new_n7286_), .A3(new_n7110_), .ZN(new_n7287_));
  INV_X1     g07031(.I(new_n7110_), .ZN(new_n7288_));
  NAND3_X1   g07032(.A1(new_n7285_), .A2(new_n7284_), .A3(new_n7283_), .ZN(new_n7289_));
  OAI21_X1   g07033(.A1(new_n7279_), .A2(new_n7281_), .B(new_n7271_), .ZN(new_n7290_));
  AOI21_X1   g07034(.A1(new_n7290_), .A2(new_n7289_), .B(new_n7288_), .ZN(new_n7291_));
  AOI21_X1   g07035(.A1(new_n5744_), .A2(new_n5745_), .B(new_n5748_), .ZN(new_n7292_));
  INV_X1     g07036(.I(new_n5797_), .ZN(new_n7293_));
  AOI21_X1   g07037(.A1(new_n5593_), .A2(new_n7293_), .B(new_n7292_), .ZN(new_n7294_));
  INV_X1     g07038(.I(new_n6049_), .ZN(new_n7295_));
  OAI21_X1   g07039(.A1(new_n7294_), .A2(new_n6038_), .B(new_n7295_), .ZN(new_n7296_));
  AOI21_X1   g07040(.A1(new_n7296_), .A2(new_n6281_), .B(new_n6279_), .ZN(new_n7297_));
  NOR3_X1    g07041(.A1(new_n6482_), .A2(new_n6481_), .A3(new_n6314_), .ZN(new_n7298_));
  OAI21_X1   g07042(.A1(new_n6482_), .A2(new_n6481_), .B(new_n6314_), .ZN(new_n7299_));
  AOI21_X1   g07043(.A1(new_n7297_), .A2(new_n7299_), .B(new_n7298_), .ZN(new_n7300_));
  AOI21_X1   g07044(.A1(new_n6770_), .A2(new_n6767_), .B(new_n6766_), .ZN(new_n7301_));
  NOR3_X1    g07045(.A1(new_n6756_), .A2(new_n6745_), .A3(new_n6763_), .ZN(new_n7302_));
  NOR2_X1    g07046(.A1(new_n7302_), .A2(new_n7301_), .ZN(new_n7303_));
  NAND2_X1   g07047(.A1(new_n6766_), .A2(new_n6815_), .ZN(new_n7304_));
  NAND2_X1   g07048(.A1(new_n6745_), .A2(new_n6746_), .ZN(new_n7305_));
  AOI21_X1   g07049(.A1(new_n7304_), .A2(new_n7305_), .B(new_n6762_), .ZN(new_n7306_));
  AOI21_X1   g07050(.A1(new_n7300_), .A2(new_n7303_), .B(new_n7306_), .ZN(new_n7307_));
  NOR3_X1    g07051(.A1(new_n7069_), .A2(new_n7070_), .A3(new_n7067_), .ZN(new_n7308_));
  AOI21_X1   g07052(.A1(new_n7059_), .A2(new_n7064_), .B(new_n6826_), .ZN(new_n7309_));
  NOR2_X1    g07053(.A1(new_n7308_), .A2(new_n7309_), .ZN(new_n7310_));
  AOI21_X1   g07054(.A1(new_n7059_), .A2(new_n7064_), .B(new_n7067_), .ZN(new_n7311_));
  INV_X1     g07055(.I(new_n7311_), .ZN(new_n7312_));
  OAI21_X1   g07056(.A1(new_n7310_), .A2(new_n7307_), .B(new_n7312_), .ZN(new_n7313_));
  NOR3_X1    g07057(.A1(new_n7313_), .A2(new_n7287_), .A3(new_n7291_), .ZN(new_n7314_));
  NAND3_X1   g07058(.A1(new_n7290_), .A2(new_n7289_), .A3(new_n7288_), .ZN(new_n7315_));
  OAI21_X1   g07059(.A1(new_n7282_), .A2(new_n7286_), .B(new_n7110_), .ZN(new_n7316_));
  AOI21_X1   g07060(.A1(new_n7072_), .A2(new_n6818_), .B(new_n7311_), .ZN(new_n7317_));
  AOI21_X1   g07061(.A1(new_n7315_), .A2(new_n7316_), .B(new_n7317_), .ZN(new_n7318_));
  OAI21_X1   g07062(.A1(new_n7314_), .A2(new_n7318_), .B(new_n7105_), .ZN(new_n7319_));
  NOR2_X1    g07063(.A1(new_n7318_), .A2(new_n7314_), .ZN(new_n7320_));
  NAND2_X1   g07064(.A1(new_n7320_), .A2(new_n7104_), .ZN(new_n7321_));
  NAND2_X1   g07065(.A1(new_n7319_), .A2(new_n7321_), .ZN(new_n7322_));
  XOR2_X1    g07066(.A1(new_n7091_), .A2(new_n7322_), .Z(\f[45] ));
  OAI21_X1   g07067(.A1(new_n7287_), .A2(new_n7317_), .B(new_n7316_), .ZN(new_n7324_));
  AOI22_X1   g07068(.A1(new_n800_), .A2(\b[42] ), .B1(\b[43] ), .B2(new_n333_), .ZN(new_n7325_));
  OAI21_X1   g07069(.A1(new_n6285_), .A2(new_n392_), .B(new_n7325_), .ZN(new_n7326_));
  INV_X1     g07070(.I(new_n7326_), .ZN(new_n7327_));
  NAND3_X1   g07071(.A1(new_n6784_), .A2(new_n6782_), .A3(new_n330_), .ZN(new_n7328_));
  AOI21_X1   g07072(.A1(new_n7328_), .A2(new_n7327_), .B(new_n312_), .ZN(new_n7329_));
  NAND3_X1   g07073(.A1(new_n7328_), .A2(new_n312_), .A3(new_n7327_), .ZN(new_n7330_));
  INV_X1     g07074(.I(new_n7330_), .ZN(new_n7331_));
  NOR2_X1    g07075(.A1(new_n7331_), .A2(new_n7329_), .ZN(new_n7332_));
  OAI21_X1   g07076(.A1(new_n7068_), .A2(new_n7053_), .B(new_n7052_), .ZN(new_n7333_));
  AOI21_X1   g07077(.A1(new_n7333_), .A2(new_n7275_), .B(new_n7271_), .ZN(new_n7334_));
  AOI22_X1   g07078(.A1(new_n518_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n636_), .ZN(new_n7335_));
  OAI21_X1   g07079(.A1(new_n5341_), .A2(new_n917_), .B(new_n7335_), .ZN(new_n7336_));
  AOI21_X1   g07080(.A1(new_n5793_), .A2(new_n618_), .B(new_n7336_), .ZN(new_n7337_));
  XOR2_X1    g07081(.A1(new_n7337_), .A2(\a[8] ), .Z(new_n7338_));
  AOI21_X1   g07082(.A1(new_n6516_), .A2(new_n6738_), .B(new_n7029_), .ZN(new_n7339_));
  OAI21_X1   g07083(.A1(new_n7339_), .A2(new_n7028_), .B(new_n7027_), .ZN(new_n7340_));
  AOI21_X1   g07084(.A1(new_n7340_), .A2(new_n7261_), .B(new_n7257_), .ZN(new_n7341_));
  AOI22_X1   g07085(.A1(new_n729_), .A2(\b[37] ), .B1(\b[36] ), .B2(new_n732_), .ZN(new_n7342_));
  OAI21_X1   g07086(.A1(new_n4666_), .A2(new_n1127_), .B(new_n7342_), .ZN(new_n7343_));
  INV_X1     g07087(.I(new_n7343_), .ZN(new_n7344_));
  OAI21_X1   g07088(.A1(new_n5322_), .A2(new_n986_), .B(new_n7344_), .ZN(new_n7345_));
  XOR2_X1    g07089(.A1(new_n7345_), .A2(\a[11] ), .Z(new_n7346_));
  OAI21_X1   g07090(.A1(new_n6445_), .A2(new_n6441_), .B(new_n6447_), .ZN(new_n7347_));
  AOI21_X1   g07091(.A1(new_n7347_), .A2(new_n6711_), .B(new_n6725_), .ZN(new_n7348_));
  AOI21_X1   g07092(.A1(new_n7348_), .A2(new_n7020_), .B(new_n7018_), .ZN(new_n7349_));
  OAI21_X1   g07093(.A1(new_n7349_), .A2(new_n7247_), .B(new_n7252_), .ZN(new_n7350_));
  OAI22_X1   g07094(.A1(new_n993_), .A2(new_n4639_), .B1(new_n4638_), .B2(new_n997_), .ZN(new_n7351_));
  AOI21_X1   g07095(.A1(\b[32] ), .A2(new_n1486_), .B(new_n7351_), .ZN(new_n7352_));
  OAI21_X1   g07096(.A1(new_n4649_), .A2(new_n1323_), .B(new_n7352_), .ZN(new_n7353_));
  XOR2_X1    g07097(.A1(new_n7353_), .A2(\a[14] ), .Z(new_n7354_));
  AOI21_X1   g07098(.A1(new_n6712_), .A2(new_n6705_), .B(new_n6840_), .ZN(new_n7355_));
  OAI21_X1   g07099(.A1(new_n7355_), .A2(new_n7007_), .B(new_n7005_), .ZN(new_n7356_));
  NOR2_X1    g07100(.A1(new_n7356_), .A2(new_n7235_), .ZN(new_n7357_));
  OR2_X2     g07101(.A1(new_n7210_), .A2(new_n7219_), .Z(new_n7358_));
  NAND2_X1   g07102(.A1(new_n7227_), .A2(new_n7225_), .ZN(new_n7359_));
  NAND2_X1   g07103(.A1(new_n7359_), .A2(new_n7358_), .ZN(new_n7360_));
  NAND2_X1   g07104(.A1(new_n7360_), .A2(new_n7228_), .ZN(new_n7361_));
  AOI21_X1   g07105(.A1(new_n7356_), .A2(new_n7235_), .B(new_n7361_), .ZN(new_n7362_));
  AOI21_X1   g07106(.A1(new_n6993_), .A2(new_n6996_), .B(new_n6994_), .ZN(new_n7363_));
  OAI21_X1   g07107(.A1(new_n7363_), .A2(new_n7226_), .B(new_n7220_), .ZN(new_n7364_));
  AOI22_X1   g07108(.A1(new_n1738_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n1743_), .ZN(new_n7365_));
  OAI21_X1   g07109(.A1(new_n3006_), .A2(new_n1931_), .B(new_n7365_), .ZN(new_n7366_));
  AOI21_X1   g07110(.A1(new_n3807_), .A2(new_n1746_), .B(new_n7366_), .ZN(new_n7367_));
  XOR2_X1    g07111(.A1(new_n7367_), .A2(new_n1736_), .Z(new_n7368_));
  AOI21_X1   g07112(.A1(new_n7216_), .A2(new_n7205_), .B(new_n7201_), .ZN(new_n7369_));
  OAI22_X1   g07113(.A1(new_n2189_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n2194_), .ZN(new_n7370_));
  AOI21_X1   g07114(.A1(\b[23] ), .A2(new_n2361_), .B(new_n7370_), .ZN(new_n7371_));
  OAI21_X1   g07115(.A1(new_n2655_), .A2(new_n2197_), .B(new_n7371_), .ZN(new_n7372_));
  XOR2_X1    g07116(.A1(new_n7372_), .A2(\a[23] ), .Z(new_n7373_));
  OAI21_X1   g07117(.A1(new_n7191_), .A2(new_n7190_), .B(new_n7184_), .ZN(new_n7374_));
  AOI22_X1   g07118(.A1(new_n2716_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n2719_), .ZN(new_n7375_));
  OAI21_X1   g07119(.A1(new_n1860_), .A2(new_n2924_), .B(new_n7375_), .ZN(new_n7376_));
  AOI21_X1   g07120(.A1(new_n2659_), .A2(new_n2722_), .B(new_n7376_), .ZN(new_n7377_));
  XOR2_X1    g07121(.A1(new_n7377_), .A2(new_n2714_), .Z(new_n7378_));
  NOR3_X1    g07122(.A1(new_n6958_), .A2(new_n7172_), .A3(new_n7176_), .ZN(new_n7379_));
  AOI21_X1   g07123(.A1(new_n6375_), .A2(new_n6376_), .B(new_n6372_), .ZN(new_n7380_));
  AOI21_X1   g07124(.A1(new_n7380_), .A2(new_n6658_), .B(new_n6861_), .ZN(new_n7381_));
  OAI21_X1   g07125(.A1(new_n7381_), .A2(new_n6957_), .B(new_n6952_), .ZN(new_n7382_));
  AOI21_X1   g07126(.A1(new_n7382_), .A2(new_n7176_), .B(new_n7194_), .ZN(new_n7383_));
  AOI22_X1   g07127(.A1(new_n3267_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n3270_), .ZN(new_n7384_));
  OAI21_X1   g07128(.A1(new_n1432_), .A2(new_n3475_), .B(new_n7384_), .ZN(new_n7385_));
  AOI21_X1   g07129(.A1(new_n1695_), .A2(new_n3273_), .B(new_n7385_), .ZN(new_n7386_));
  XOR2_X1    g07130(.A1(new_n7386_), .A2(new_n3264_), .Z(new_n7387_));
  NAND2_X1   g07131(.A1(new_n7168_), .A2(new_n7167_), .ZN(new_n7388_));
  AOI22_X1   g07132(.A1(new_n3864_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n3869_), .ZN(new_n7389_));
  OAI21_X1   g07133(.A1(new_n1093_), .A2(new_n5410_), .B(new_n7389_), .ZN(new_n7390_));
  AOI21_X1   g07134(.A1(new_n1701_), .A2(new_n3872_), .B(new_n7390_), .ZN(new_n7391_));
  XOR2_X1    g07135(.A1(new_n7391_), .A2(new_n3876_), .Z(new_n7392_));
  AOI21_X1   g07136(.A1(new_n6942_), .A2(new_n6929_), .B(new_n7152_), .ZN(new_n7393_));
  OAI21_X1   g07137(.A1(new_n7164_), .A2(new_n7393_), .B(new_n7153_), .ZN(new_n7394_));
  OAI21_X1   g07138(.A1(new_n7133_), .A2(new_n7139_), .B(new_n7144_), .ZN(new_n7395_));
  AOI21_X1   g07139(.A1(new_n7128_), .A2(new_n7127_), .B(new_n7123_), .ZN(new_n7396_));
  AOI22_X1   g07140(.A1(new_n6569_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n6574_), .ZN(new_n7397_));
  NAND2_X1   g07141(.A1(new_n6887_), .A2(\b[2] ), .ZN(new_n7398_));
  NAND2_X1   g07142(.A1(new_n1725_), .A2(new_n6579_), .ZN(new_n7399_));
  NAND3_X1   g07143(.A1(new_n7399_), .A2(new_n7397_), .A3(new_n7398_), .ZN(new_n7400_));
  XOR2_X1    g07144(.A1(new_n7400_), .A2(new_n6567_), .Z(new_n7401_));
  XOR2_X1    g07145(.A1(\a[46] ), .A2(\a[47] ), .Z(new_n7402_));
  NOR2_X1    g07146(.A1(new_n7116_), .A2(new_n7402_), .ZN(new_n7403_));
  INV_X1     g07147(.I(\a[45] ), .ZN(new_n7404_));
  NAND3_X1   g07148(.A1(new_n6567_), .A2(new_n7404_), .A3(\a[46] ), .ZN(new_n7405_));
  INV_X1     g07149(.I(\a[46] ), .ZN(new_n7406_));
  NAND3_X1   g07150(.A1(new_n7406_), .A2(\a[44] ), .A3(\a[45] ), .ZN(new_n7407_));
  NAND2_X1   g07151(.A1(new_n7405_), .A2(new_n7407_), .ZN(new_n7408_));
  AOI22_X1   g07152(.A1(new_n7403_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n7408_), .ZN(new_n7409_));
  INV_X1     g07153(.I(\a[47] ), .ZN(new_n7410_));
  NOR2_X1    g07154(.A1(new_n7410_), .A2(\a[46] ), .ZN(new_n7411_));
  NOR2_X1    g07155(.A1(new_n7406_), .A2(\a[47] ), .ZN(new_n7412_));
  NOR2_X1    g07156(.A1(new_n7411_), .A2(new_n7412_), .ZN(new_n7413_));
  NOR2_X1    g07157(.A1(new_n7413_), .A2(new_n7116_), .ZN(new_n7414_));
  NAND2_X1   g07158(.A1(new_n7414_), .A2(new_n263_), .ZN(new_n7415_));
  NAND2_X1   g07159(.A1(new_n7409_), .A2(new_n7415_), .ZN(new_n7416_));
  NAND2_X1   g07160(.A1(new_n7416_), .A2(\a[47] ), .ZN(new_n7417_));
  INV_X1     g07161(.I(new_n7416_), .ZN(new_n7418_));
  NAND2_X1   g07162(.A1(new_n7418_), .A2(new_n7410_), .ZN(new_n7419_));
  NOR2_X1    g07163(.A1(new_n7117_), .A2(new_n7410_), .ZN(new_n7420_));
  INV_X1     g07164(.I(new_n7420_), .ZN(new_n7421_));
  NAND3_X1   g07165(.A1(new_n7419_), .A2(new_n7417_), .A3(new_n7421_), .ZN(new_n7422_));
  NOR2_X1    g07166(.A1(new_n7417_), .A2(new_n7117_), .ZN(new_n7423_));
  INV_X1     g07167(.I(new_n7423_), .ZN(new_n7424_));
  AOI21_X1   g07168(.A1(new_n7422_), .A2(new_n7424_), .B(new_n7401_), .ZN(new_n7425_));
  NAND3_X1   g07169(.A1(new_n7401_), .A2(new_n7422_), .A3(new_n7424_), .ZN(new_n7426_));
  INV_X1     g07170(.I(new_n7426_), .ZN(new_n7427_));
  NOR2_X1    g07171(.A1(new_n7120_), .A2(new_n7117_), .ZN(new_n7428_));
  AOI21_X1   g07172(.A1(new_n6894_), .A2(new_n7121_), .B(new_n7428_), .ZN(new_n7429_));
  OAI21_X1   g07173(.A1(new_n7425_), .A2(new_n7427_), .B(new_n7429_), .ZN(new_n7430_));
  INV_X1     g07174(.I(new_n7430_), .ZN(new_n7431_));
  NOR3_X1    g07175(.A1(new_n7429_), .A2(new_n7425_), .A3(new_n7427_), .ZN(new_n7432_));
  OAI22_X1   g07176(.A1(new_n5852_), .A2(new_n471_), .B1(new_n438_), .B2(new_n5857_), .ZN(new_n7433_));
  AOI21_X1   g07177(.A1(\b[5] ), .A2(new_n6115_), .B(new_n7433_), .ZN(new_n7434_));
  OAI21_X1   g07178(.A1(new_n485_), .A2(new_n5861_), .B(new_n7434_), .ZN(new_n7435_));
  XOR2_X1    g07179(.A1(new_n7435_), .A2(\a[41] ), .Z(new_n7436_));
  NOR3_X1    g07180(.A1(new_n7431_), .A2(new_n7432_), .A3(new_n7436_), .ZN(new_n7437_));
  INV_X1     g07181(.I(new_n7432_), .ZN(new_n7438_));
  INV_X1     g07182(.I(new_n7436_), .ZN(new_n7439_));
  AOI21_X1   g07183(.A1(new_n7438_), .A2(new_n7430_), .B(new_n7439_), .ZN(new_n7440_));
  NOR2_X1    g07184(.A1(new_n7437_), .A2(new_n7440_), .ZN(new_n7441_));
  OAI21_X1   g07185(.A1(new_n7130_), .A2(new_n7396_), .B(new_n7441_), .ZN(new_n7442_));
  NOR3_X1    g07186(.A1(new_n7441_), .A2(new_n7130_), .A3(new_n7396_), .ZN(new_n7443_));
  INV_X1     g07187(.I(new_n7443_), .ZN(new_n7444_));
  AOI22_X1   g07188(.A1(new_n5155_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n5160_), .ZN(new_n7445_));
  OAI21_X1   g07189(.A1(new_n577_), .A2(new_n6877_), .B(new_n7445_), .ZN(new_n7446_));
  AOI21_X1   g07190(.A1(new_n1059_), .A2(new_n5166_), .B(new_n7446_), .ZN(new_n7447_));
  XOR2_X1    g07191(.A1(new_n7447_), .A2(new_n5162_), .Z(new_n7448_));
  INV_X1     g07192(.I(new_n7448_), .ZN(new_n7449_));
  NAND3_X1   g07193(.A1(new_n7444_), .A2(new_n7442_), .A3(new_n7449_), .ZN(new_n7450_));
  INV_X1     g07194(.I(new_n7442_), .ZN(new_n7451_));
  OAI21_X1   g07195(.A1(new_n7451_), .A2(new_n7443_), .B(new_n7448_), .ZN(new_n7452_));
  NAND2_X1   g07196(.A1(new_n7452_), .A2(new_n7450_), .ZN(new_n7453_));
  NAND2_X1   g07197(.A1(new_n7395_), .A2(new_n7453_), .ZN(new_n7454_));
  AOI21_X1   g07198(.A1(new_n7142_), .A2(new_n7143_), .B(new_n7140_), .ZN(new_n7455_));
  NOR3_X1    g07199(.A1(new_n7451_), .A2(new_n7443_), .A3(new_n7448_), .ZN(new_n7456_));
  AOI21_X1   g07200(.A1(new_n7444_), .A2(new_n7442_), .B(new_n7449_), .ZN(new_n7457_));
  NOR2_X1    g07201(.A1(new_n7456_), .A2(new_n7457_), .ZN(new_n7458_));
  NAND2_X1   g07202(.A1(new_n7455_), .A2(new_n7458_), .ZN(new_n7459_));
  OAI22_X1   g07203(.A1(new_n1070_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n941_), .ZN(new_n7460_));
  AOI21_X1   g07204(.A1(\b[11] ), .A2(new_n4706_), .B(new_n7460_), .ZN(new_n7461_));
  OAI21_X1   g07205(.A1(new_n1082_), .A2(new_n4458_), .B(new_n7461_), .ZN(new_n7462_));
  XOR2_X1    g07206(.A1(new_n7462_), .A2(\a[35] ), .Z(new_n7463_));
  AOI21_X1   g07207(.A1(new_n7454_), .A2(new_n7459_), .B(new_n7463_), .ZN(new_n7464_));
  NOR2_X1    g07208(.A1(new_n7455_), .A2(new_n7458_), .ZN(new_n7465_));
  NOR2_X1    g07209(.A1(new_n7139_), .A2(new_n7133_), .ZN(new_n7466_));
  NOR3_X1    g07210(.A1(new_n7466_), .A2(new_n7453_), .A3(new_n7140_), .ZN(new_n7467_));
  INV_X1     g07211(.I(new_n7463_), .ZN(new_n7468_));
  NOR3_X1    g07212(.A1(new_n7465_), .A2(new_n7467_), .A3(new_n7468_), .ZN(new_n7469_));
  NOR2_X1    g07213(.A1(new_n7464_), .A2(new_n7469_), .ZN(new_n7470_));
  NAND2_X1   g07214(.A1(new_n7394_), .A2(new_n7470_), .ZN(new_n7471_));
  OAI21_X1   g07215(.A1(new_n6628_), .A2(new_n6621_), .B(new_n6630_), .ZN(new_n7472_));
  AOI21_X1   g07216(.A1(new_n7472_), .A2(new_n6939_), .B(new_n6937_), .ZN(new_n7473_));
  OAI21_X1   g07217(.A1(new_n7473_), .A2(new_n7152_), .B(new_n7146_), .ZN(new_n7474_));
  OAI21_X1   g07218(.A1(new_n7465_), .A2(new_n7467_), .B(new_n7468_), .ZN(new_n7475_));
  NAND3_X1   g07219(.A1(new_n7454_), .A2(new_n7459_), .A3(new_n7463_), .ZN(new_n7476_));
  NAND2_X1   g07220(.A1(new_n7475_), .A2(new_n7476_), .ZN(new_n7477_));
  NAND3_X1   g07221(.A1(new_n7477_), .A2(new_n7474_), .A3(new_n7153_), .ZN(new_n7478_));
  NAND3_X1   g07222(.A1(new_n7471_), .A2(new_n7478_), .A3(new_n7392_), .ZN(new_n7479_));
  INV_X1     g07223(.I(new_n7392_), .ZN(new_n7480_));
  AOI21_X1   g07224(.A1(new_n7474_), .A2(new_n7153_), .B(new_n7477_), .ZN(new_n7481_));
  NOR3_X1    g07225(.A1(new_n6935_), .A2(new_n6937_), .A3(new_n7150_), .ZN(new_n7482_));
  NOR2_X1    g07226(.A1(new_n7393_), .A2(new_n7164_), .ZN(new_n7483_));
  NOR3_X1    g07227(.A1(new_n7483_), .A2(new_n7470_), .A3(new_n7482_), .ZN(new_n7484_));
  OAI21_X1   g07228(.A1(new_n7481_), .A2(new_n7484_), .B(new_n7480_), .ZN(new_n7485_));
  NAND2_X1   g07229(.A1(new_n7485_), .A2(new_n7479_), .ZN(new_n7486_));
  NAND3_X1   g07230(.A1(new_n7388_), .A2(new_n7486_), .A3(new_n7169_), .ZN(new_n7487_));
  NOR2_X1    g07231(.A1(new_n7161_), .A2(new_n7155_), .ZN(new_n7488_));
  NOR3_X1    g07232(.A1(new_n7481_), .A2(new_n7484_), .A3(new_n7480_), .ZN(new_n7489_));
  AOI21_X1   g07233(.A1(new_n7471_), .A2(new_n7478_), .B(new_n7392_), .ZN(new_n7490_));
  NOR2_X1    g07234(.A1(new_n7489_), .A2(new_n7490_), .ZN(new_n7491_));
  OAI21_X1   g07235(.A1(new_n7488_), .A2(new_n7162_), .B(new_n7491_), .ZN(new_n7492_));
  NAND3_X1   g07236(.A1(new_n7492_), .A2(new_n7487_), .A3(new_n7387_), .ZN(new_n7493_));
  INV_X1     g07237(.I(new_n7387_), .ZN(new_n7494_));
  NOR3_X1    g07238(.A1(new_n7488_), .A2(new_n7162_), .A3(new_n7491_), .ZN(new_n7495_));
  AOI21_X1   g07239(.A1(new_n7167_), .A2(new_n7168_), .B(new_n7162_), .ZN(new_n7496_));
  NOR2_X1    g07240(.A1(new_n7496_), .A2(new_n7486_), .ZN(new_n7497_));
  OAI21_X1   g07241(.A1(new_n7495_), .A2(new_n7497_), .B(new_n7494_), .ZN(new_n7498_));
  NAND2_X1   g07242(.A1(new_n7498_), .A2(new_n7493_), .ZN(new_n7499_));
  NOR3_X1    g07243(.A1(new_n7383_), .A2(new_n7499_), .A3(new_n7379_), .ZN(new_n7500_));
  OAI21_X1   g07244(.A1(new_n7179_), .A2(new_n7178_), .B(new_n7171_), .ZN(new_n7501_));
  NOR3_X1    g07245(.A1(new_n7495_), .A2(new_n7497_), .A3(new_n7494_), .ZN(new_n7502_));
  AOI21_X1   g07246(.A1(new_n7492_), .A2(new_n7487_), .B(new_n7387_), .ZN(new_n7503_));
  NOR2_X1    g07247(.A1(new_n7502_), .A2(new_n7503_), .ZN(new_n7504_));
  AOI21_X1   g07248(.A1(new_n7501_), .A2(new_n7180_), .B(new_n7504_), .ZN(new_n7505_));
  OAI21_X1   g07249(.A1(new_n7505_), .A2(new_n7500_), .B(new_n7378_), .ZN(new_n7506_));
  INV_X1     g07250(.I(new_n7378_), .ZN(new_n7507_));
  NAND3_X1   g07251(.A1(new_n7504_), .A2(new_n7501_), .A3(new_n7180_), .ZN(new_n7508_));
  OAI21_X1   g07252(.A1(new_n7383_), .A2(new_n7379_), .B(new_n7499_), .ZN(new_n7509_));
  NAND3_X1   g07253(.A1(new_n7509_), .A2(new_n7508_), .A3(new_n7507_), .ZN(new_n7510_));
  NAND2_X1   g07254(.A1(new_n7506_), .A2(new_n7510_), .ZN(new_n7511_));
  NAND3_X1   g07255(.A1(new_n7374_), .A2(new_n7192_), .A3(new_n7511_), .ZN(new_n7512_));
  AOI21_X1   g07256(.A1(new_n6379_), .A2(new_n6389_), .B(new_n6387_), .ZN(new_n7513_));
  AOI21_X1   g07257(.A1(new_n7513_), .A2(new_n6664_), .B(new_n6660_), .ZN(new_n7514_));
  OAI21_X1   g07258(.A1(new_n7514_), .A2(new_n6966_), .B(new_n6965_), .ZN(new_n7515_));
  AOI21_X1   g07259(.A1(new_n7515_), .A2(new_n7188_), .B(new_n7197_), .ZN(new_n7516_));
  AOI21_X1   g07260(.A1(new_n7509_), .A2(new_n7508_), .B(new_n7507_), .ZN(new_n7517_));
  NOR3_X1    g07261(.A1(new_n7505_), .A2(new_n7500_), .A3(new_n7378_), .ZN(new_n7518_));
  NOR2_X1    g07262(.A1(new_n7518_), .A2(new_n7517_), .ZN(new_n7519_));
  OAI21_X1   g07263(.A1(new_n7516_), .A2(new_n7199_), .B(new_n7519_), .ZN(new_n7520_));
  NAND3_X1   g07264(.A1(new_n7520_), .A2(new_n7512_), .A3(new_n7373_), .ZN(new_n7521_));
  INV_X1     g07265(.I(new_n7373_), .ZN(new_n7522_));
  NOR3_X1    g07266(.A1(new_n7516_), .A2(new_n7199_), .A3(new_n7519_), .ZN(new_n7523_));
  AOI21_X1   g07267(.A1(new_n7374_), .A2(new_n7192_), .B(new_n7511_), .ZN(new_n7524_));
  OAI21_X1   g07268(.A1(new_n7523_), .A2(new_n7524_), .B(new_n7522_), .ZN(new_n7525_));
  NAND2_X1   g07269(.A1(new_n7525_), .A2(new_n7521_), .ZN(new_n7526_));
  NOR3_X1    g07270(.A1(new_n7369_), .A2(new_n7526_), .A3(new_n7209_), .ZN(new_n7527_));
  OAI21_X1   g07271(.A1(new_n7207_), .A2(new_n7206_), .B(new_n7213_), .ZN(new_n7528_));
  NOR3_X1    g07272(.A1(new_n7523_), .A2(new_n7524_), .A3(new_n7522_), .ZN(new_n7529_));
  AOI21_X1   g07273(.A1(new_n7520_), .A2(new_n7512_), .B(new_n7373_), .ZN(new_n7530_));
  NOR2_X1    g07274(.A1(new_n7529_), .A2(new_n7530_), .ZN(new_n7531_));
  AOI21_X1   g07275(.A1(new_n7528_), .A2(new_n7218_), .B(new_n7531_), .ZN(new_n7532_));
  OAI21_X1   g07276(.A1(new_n7532_), .A2(new_n7527_), .B(new_n7368_), .ZN(new_n7533_));
  INV_X1     g07277(.I(new_n7368_), .ZN(new_n7534_));
  NAND3_X1   g07278(.A1(new_n7528_), .A2(new_n7531_), .A3(new_n7218_), .ZN(new_n7535_));
  OAI21_X1   g07279(.A1(new_n7369_), .A2(new_n7209_), .B(new_n7526_), .ZN(new_n7536_));
  NAND3_X1   g07280(.A1(new_n7536_), .A2(new_n7535_), .A3(new_n7534_), .ZN(new_n7537_));
  NAND2_X1   g07281(.A1(new_n7533_), .A2(new_n7537_), .ZN(new_n7538_));
  AOI21_X1   g07282(.A1(new_n7364_), .A2(new_n7227_), .B(new_n7538_), .ZN(new_n7539_));
  NOR3_X1    g07283(.A1(new_n6992_), .A2(new_n6994_), .A3(new_n7224_), .ZN(new_n7540_));
  AOI21_X1   g07284(.A1(new_n6697_), .A2(new_n6687_), .B(new_n6682_), .ZN(new_n7541_));
  OAI21_X1   g07285(.A1(new_n7541_), .A2(new_n6991_), .B(new_n6985_), .ZN(new_n7542_));
  AOI21_X1   g07286(.A1(new_n7224_), .A2(new_n7542_), .B(new_n7358_), .ZN(new_n7543_));
  AOI21_X1   g07287(.A1(new_n7536_), .A2(new_n7535_), .B(new_n7534_), .ZN(new_n7544_));
  NOR3_X1    g07288(.A1(new_n7532_), .A2(new_n7527_), .A3(new_n7368_), .ZN(new_n7545_));
  NOR2_X1    g07289(.A1(new_n7545_), .A2(new_n7544_), .ZN(new_n7546_));
  NOR3_X1    g07290(.A1(new_n7543_), .A2(new_n7540_), .A3(new_n7546_), .ZN(new_n7547_));
  OAI22_X1   g07291(.A1(new_n1592_), .A2(new_n4022_), .B1(new_n3624_), .B2(new_n1505_), .ZN(new_n7548_));
  AOI21_X1   g07292(.A1(\b[29] ), .A2(new_n1584_), .B(new_n7548_), .ZN(new_n7549_));
  OAI21_X1   g07293(.A1(new_n6003_), .A2(new_n1732_), .B(new_n7549_), .ZN(new_n7550_));
  XOR2_X1    g07294(.A1(new_n7550_), .A2(new_n1344_), .Z(new_n7551_));
  NOR3_X1    g07295(.A1(new_n7547_), .A2(new_n7539_), .A3(new_n7551_), .ZN(new_n7552_));
  OAI21_X1   g07296(.A1(new_n7543_), .A2(new_n7540_), .B(new_n7546_), .ZN(new_n7553_));
  NAND3_X1   g07297(.A1(new_n7364_), .A2(new_n7227_), .A3(new_n7538_), .ZN(new_n7554_));
  XOR2_X1    g07298(.A1(new_n7550_), .A2(\a[17] ), .Z(new_n7555_));
  AOI21_X1   g07299(.A1(new_n7553_), .A2(new_n7554_), .B(new_n7555_), .ZN(new_n7556_));
  NOR2_X1    g07300(.A1(new_n7552_), .A2(new_n7556_), .ZN(new_n7557_));
  OAI21_X1   g07301(.A1(new_n7362_), .A2(new_n7357_), .B(new_n7557_), .ZN(new_n7558_));
  AOI21_X1   g07302(.A1(new_n7012_), .A2(new_n7002_), .B(new_n6998_), .ZN(new_n7559_));
  OAI21_X1   g07303(.A1(new_n7559_), .A2(new_n7237_), .B(new_n7231_), .ZN(new_n7560_));
  NAND3_X1   g07304(.A1(new_n7553_), .A2(new_n7554_), .A3(new_n7555_), .ZN(new_n7561_));
  OAI21_X1   g07305(.A1(new_n7547_), .A2(new_n7539_), .B(new_n7551_), .ZN(new_n7562_));
  NAND2_X1   g07306(.A1(new_n7562_), .A2(new_n7561_), .ZN(new_n7563_));
  NAND3_X1   g07307(.A1(new_n7560_), .A2(new_n7563_), .A3(new_n7238_), .ZN(new_n7564_));
  NAND3_X1   g07308(.A1(new_n7558_), .A2(new_n7564_), .A3(new_n7354_), .ZN(new_n7565_));
  INV_X1     g07309(.I(new_n7354_), .ZN(new_n7566_));
  AOI21_X1   g07310(.A1(new_n7560_), .A2(new_n7238_), .B(new_n7563_), .ZN(new_n7567_));
  NOR3_X1    g07311(.A1(new_n7362_), .A2(new_n7557_), .A3(new_n7357_), .ZN(new_n7568_));
  OAI21_X1   g07312(.A1(new_n7568_), .A2(new_n7567_), .B(new_n7566_), .ZN(new_n7569_));
  NAND2_X1   g07313(.A1(new_n7569_), .A2(new_n7565_), .ZN(new_n7570_));
  NAND3_X1   g07314(.A1(new_n7350_), .A2(new_n7254_), .A3(new_n7570_), .ZN(new_n7571_));
  AOI21_X1   g07315(.A1(new_n6433_), .A2(new_n6446_), .B(new_n6442_), .ZN(new_n7572_));
  OAI21_X1   g07316(.A1(new_n7572_), .A2(new_n6724_), .B(new_n6717_), .ZN(new_n7573_));
  OAI21_X1   g07317(.A1(new_n7573_), .A2(new_n7015_), .B(new_n7009_), .ZN(new_n7574_));
  AOI21_X1   g07318(.A1(new_n7574_), .A2(new_n7246_), .B(new_n7242_), .ZN(new_n7575_));
  NOR3_X1    g07319(.A1(new_n7568_), .A2(new_n7567_), .A3(new_n7566_), .ZN(new_n7576_));
  AOI21_X1   g07320(.A1(new_n7558_), .A2(new_n7564_), .B(new_n7354_), .ZN(new_n7577_));
  NOR2_X1    g07321(.A1(new_n7576_), .A2(new_n7577_), .ZN(new_n7578_));
  OAI21_X1   g07322(.A1(new_n7575_), .A2(new_n7249_), .B(new_n7578_), .ZN(new_n7579_));
  NAND3_X1   g07323(.A1(new_n7571_), .A2(new_n7579_), .A3(new_n7346_), .ZN(new_n7580_));
  XOR2_X1    g07324(.A1(new_n7345_), .A2(new_n722_), .Z(new_n7581_));
  NOR3_X1    g07325(.A1(new_n7575_), .A2(new_n7249_), .A3(new_n7578_), .ZN(new_n7582_));
  AOI21_X1   g07326(.A1(new_n7350_), .A2(new_n7254_), .B(new_n7570_), .ZN(new_n7583_));
  OAI21_X1   g07327(.A1(new_n7583_), .A2(new_n7582_), .B(new_n7581_), .ZN(new_n7584_));
  NAND2_X1   g07328(.A1(new_n7584_), .A2(new_n7580_), .ZN(new_n7585_));
  NOR3_X1    g07329(.A1(new_n7341_), .A2(new_n7266_), .A3(new_n7585_), .ZN(new_n7586_));
  OAI21_X1   g07330(.A1(new_n6735_), .A2(new_n6732_), .B(new_n7038_), .ZN(new_n7587_));
  AOI21_X1   g07331(.A1(new_n7587_), .A2(new_n7037_), .B(new_n7036_), .ZN(new_n7588_));
  OAI21_X1   g07332(.A1(new_n7588_), .A2(new_n7262_), .B(new_n7256_), .ZN(new_n7589_));
  NOR3_X1    g07333(.A1(new_n7583_), .A2(new_n7582_), .A3(new_n7581_), .ZN(new_n7590_));
  AOI21_X1   g07334(.A1(new_n7571_), .A2(new_n7579_), .B(new_n7346_), .ZN(new_n7591_));
  NOR2_X1    g07335(.A1(new_n7591_), .A2(new_n7590_), .ZN(new_n7592_));
  AOI21_X1   g07336(.A1(new_n7589_), .A2(new_n7269_), .B(new_n7592_), .ZN(new_n7593_));
  NOR3_X1    g07337(.A1(new_n7586_), .A2(new_n7593_), .A3(new_n7338_), .ZN(new_n7594_));
  XOR2_X1    g07338(.A1(new_n7337_), .A2(new_n488_), .Z(new_n7595_));
  NAND3_X1   g07339(.A1(new_n7589_), .A2(new_n7592_), .A3(new_n7269_), .ZN(new_n7596_));
  OAI21_X1   g07340(.A1(new_n7341_), .A2(new_n7266_), .B(new_n7585_), .ZN(new_n7597_));
  AOI21_X1   g07341(.A1(new_n7597_), .A2(new_n7596_), .B(new_n7595_), .ZN(new_n7598_));
  NOR2_X1    g07342(.A1(new_n7594_), .A2(new_n7598_), .ZN(new_n7599_));
  OAI21_X1   g07343(.A1(new_n7334_), .A2(new_n7281_), .B(new_n7599_), .ZN(new_n7600_));
  AOI21_X1   g07344(.A1(new_n7058_), .A2(new_n7062_), .B(new_n7061_), .ZN(new_n7601_));
  OAI21_X1   g07345(.A1(new_n7601_), .A2(new_n7276_), .B(new_n7283_), .ZN(new_n7602_));
  NAND3_X1   g07346(.A1(new_n7597_), .A2(new_n7596_), .A3(new_n7595_), .ZN(new_n7603_));
  OAI21_X1   g07347(.A1(new_n7586_), .A2(new_n7593_), .B(new_n7338_), .ZN(new_n7604_));
  NAND2_X1   g07348(.A1(new_n7604_), .A2(new_n7603_), .ZN(new_n7605_));
  NAND3_X1   g07349(.A1(new_n7602_), .A2(new_n7285_), .A3(new_n7605_), .ZN(new_n7606_));
  NAND3_X1   g07350(.A1(new_n7600_), .A2(new_n7606_), .A3(new_n7332_), .ZN(new_n7607_));
  INV_X1     g07351(.I(new_n7329_), .ZN(new_n7608_));
  NAND2_X1   g07352(.A1(new_n7608_), .A2(new_n7330_), .ZN(new_n7609_));
  AOI21_X1   g07353(.A1(new_n7602_), .A2(new_n7285_), .B(new_n7605_), .ZN(new_n7610_));
  NOR3_X1    g07354(.A1(new_n7334_), .A2(new_n7281_), .A3(new_n7599_), .ZN(new_n7611_));
  OAI21_X1   g07355(.A1(new_n7611_), .A2(new_n7610_), .B(new_n7609_), .ZN(new_n7612_));
  NAND2_X1   g07356(.A1(new_n7612_), .A2(new_n7607_), .ZN(new_n7613_));
  XOR2_X1    g07357(.A1(new_n7613_), .A2(new_n7324_), .Z(new_n7614_));
  INV_X1     g07358(.I(new_n7614_), .ZN(new_n7615_));
  INV_X1     g07359(.I(new_n7319_), .ZN(new_n7616_));
  INV_X1     g07360(.I(\b[46] ), .ZN(new_n7617_));
  OAI22_X1   g07361(.A1(new_n277_), .A2(new_n7617_), .B1(new_n7096_), .B2(new_n262_), .ZN(new_n7618_));
  AOI21_X1   g07362(.A1(\b[44] ), .A2(new_n283_), .B(new_n7618_), .ZN(new_n7619_));
  AOI21_X1   g07363(.A1(new_n7097_), .A2(\b[44] ), .B(\b[43] ), .ZN(new_n7620_));
  NOR2_X1    g07364(.A1(new_n7099_), .A2(\b[44] ), .ZN(new_n7621_));
  NOR2_X1    g07365(.A1(new_n7620_), .A2(new_n7621_), .ZN(new_n7622_));
  XNOR2_X1   g07366(.A1(\b[45] ), .A2(\b[46] ), .ZN(new_n7623_));
  NOR2_X1    g07367(.A1(new_n7622_), .A2(new_n7623_), .ZN(new_n7624_));
  XOR2_X1    g07368(.A1(\b[45] ), .A2(\b[46] ), .Z(new_n7625_));
  NOR3_X1    g07369(.A1(new_n7620_), .A2(new_n7621_), .A3(new_n7625_), .ZN(new_n7626_));
  NOR2_X1    g07370(.A1(new_n7624_), .A2(new_n7626_), .ZN(new_n7627_));
  OAI21_X1   g07371(.A1(new_n7627_), .A2(new_n279_), .B(new_n7619_), .ZN(new_n7628_));
  XOR2_X1    g07372(.A1(new_n7628_), .A2(\a[2] ), .Z(new_n7629_));
  OAI21_X1   g07373(.A1(new_n6807_), .A2(new_n6794_), .B(new_n6774_), .ZN(new_n7630_));
  AOI21_X1   g07374(.A1(new_n7630_), .A2(new_n6808_), .B(new_n7086_), .ZN(new_n7631_));
  NOR3_X1    g07375(.A1(new_n7631_), .A2(new_n7322_), .A3(new_n7084_), .ZN(new_n7632_));
  OAI21_X1   g07376(.A1(new_n7632_), .A2(new_n7616_), .B(new_n7629_), .ZN(new_n7633_));
  INV_X1     g07377(.I(new_n7629_), .ZN(new_n7634_));
  NAND4_X1   g07378(.A1(new_n7090_), .A2(new_n7089_), .A3(new_n7319_), .A4(new_n7321_), .ZN(new_n7635_));
  NAND3_X1   g07379(.A1(new_n7635_), .A2(new_n7319_), .A3(new_n7634_), .ZN(new_n7636_));
  NAND2_X1   g07380(.A1(new_n7633_), .A2(new_n7636_), .ZN(new_n7637_));
  XOR2_X1    g07381(.A1(new_n7637_), .A2(new_n7615_), .Z(\f[46] ));
  AOI21_X1   g07382(.A1(new_n7635_), .A2(new_n7319_), .B(new_n7634_), .ZN(new_n7639_));
  OAI21_X1   g07383(.A1(new_n7614_), .A2(new_n7639_), .B(new_n7636_), .ZN(new_n7640_));
  AOI22_X1   g07384(.A1(new_n267_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n261_), .ZN(new_n7641_));
  OAI21_X1   g07385(.A1(new_n7096_), .A2(new_n284_), .B(new_n7641_), .ZN(new_n7642_));
  OAI21_X1   g07386(.A1(new_n7620_), .A2(new_n7621_), .B(new_n7096_), .ZN(new_n7643_));
  NOR2_X1    g07387(.A1(new_n7643_), .A2(new_n7617_), .ZN(new_n7644_));
  NOR4_X1    g07388(.A1(new_n7620_), .A2(new_n7621_), .A3(new_n7096_), .A4(\b[46] ), .ZN(new_n7645_));
  OAI21_X1   g07389(.A1(new_n7644_), .A2(new_n7645_), .B(\b[47] ), .ZN(new_n7646_));
  INV_X1     g07390(.I(new_n7646_), .ZN(new_n7647_));
  NOR3_X1    g07391(.A1(new_n7644_), .A2(\b[47] ), .A3(new_n7645_), .ZN(new_n7648_));
  NOR2_X1    g07392(.A1(new_n7647_), .A2(new_n7648_), .ZN(new_n7649_));
  AOI21_X1   g07393(.A1(new_n7649_), .A2(new_n265_), .B(new_n7642_), .ZN(new_n7650_));
  XOR2_X1    g07394(.A1(new_n7650_), .A2(new_n270_), .Z(new_n7651_));
  INV_X1     g07395(.I(new_n7651_), .ZN(new_n7652_));
  AOI21_X1   g07396(.A1(new_n7283_), .A2(new_n7284_), .B(new_n7281_), .ZN(new_n7653_));
  OAI21_X1   g07397(.A1(new_n7653_), .A2(new_n7594_), .B(new_n7604_), .ZN(new_n7654_));
  AOI22_X1   g07398(.A1(new_n518_), .A2(\b[41] ), .B1(\b[40] ), .B2(new_n636_), .ZN(new_n7655_));
  OAI21_X1   g07399(.A1(new_n5761_), .A2(new_n917_), .B(new_n7655_), .ZN(new_n7656_));
  INV_X1     g07400(.I(new_n7656_), .ZN(new_n7657_));
  NAND3_X1   g07401(.A1(new_n6298_), .A2(new_n6295_), .A3(new_n618_), .ZN(new_n7658_));
  AOI21_X1   g07402(.A1(new_n7658_), .A2(new_n7657_), .B(new_n488_), .ZN(new_n7659_));
  AOI21_X1   g07403(.A1(new_n6288_), .A2(new_n6289_), .B(new_n6297_), .ZN(new_n7660_));
  NOR2_X1    g07404(.A1(new_n6294_), .A2(new_n6290_), .ZN(new_n7661_));
  NOR3_X1    g07405(.A1(new_n7660_), .A2(new_n624_), .A3(new_n7661_), .ZN(new_n7662_));
  NOR3_X1    g07406(.A1(new_n7662_), .A2(\a[8] ), .A3(new_n7656_), .ZN(new_n7663_));
  NOR2_X1    g07407(.A1(new_n7663_), .A2(new_n7659_), .ZN(new_n7664_));
  OAI22_X1   g07408(.A1(new_n713_), .A2(new_n5341_), .B1(new_n5312_), .B2(new_n717_), .ZN(new_n7665_));
  AOI21_X1   g07409(.A1(\b[36] ), .A2(new_n1126_), .B(new_n7665_), .ZN(new_n7666_));
  OAI21_X1   g07410(.A1(new_n5352_), .A2(new_n986_), .B(new_n7666_), .ZN(new_n7667_));
  XOR2_X1    g07411(.A1(new_n7667_), .A2(\a[11] ), .Z(new_n7668_));
  AOI22_X1   g07412(.A1(new_n1006_), .A2(\b[35] ), .B1(\b[34] ), .B2(new_n1009_), .ZN(new_n7669_));
  OAI21_X1   g07413(.A1(new_n4638_), .A2(new_n1481_), .B(new_n7669_), .ZN(new_n7670_));
  INV_X1     g07414(.I(new_n7670_), .ZN(new_n7671_));
  OAI21_X1   g07415(.A1(new_n4676_), .A2(new_n1323_), .B(new_n7671_), .ZN(new_n7672_));
  XOR2_X1    g07416(.A1(new_n7672_), .A2(\a[14] ), .Z(new_n7673_));
  OAI21_X1   g07417(.A1(new_n7362_), .A2(new_n7357_), .B(new_n7561_), .ZN(new_n7674_));
  OAI22_X1   g07418(.A1(new_n1592_), .A2(new_n4023_), .B1(new_n4022_), .B2(new_n1505_), .ZN(new_n7675_));
  AOI21_X1   g07419(.A1(\b[30] ), .A2(new_n1584_), .B(new_n7675_), .ZN(new_n7676_));
  OAI21_X1   g07420(.A1(new_n4031_), .A2(new_n1732_), .B(new_n7676_), .ZN(new_n7677_));
  XOR2_X1    g07421(.A1(new_n7677_), .A2(\a[17] ), .Z(new_n7678_));
  INV_X1     g07422(.I(new_n7678_), .ZN(new_n7679_));
  NOR3_X1    g07423(.A1(new_n7532_), .A2(new_n7527_), .A3(new_n7534_), .ZN(new_n7680_));
  INV_X1     g07424(.I(new_n7680_), .ZN(new_n7681_));
  AOI22_X1   g07425(.A1(new_n1738_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n1743_), .ZN(new_n7682_));
  OAI21_X1   g07426(.A1(new_n3158_), .A2(new_n1931_), .B(new_n7682_), .ZN(new_n7683_));
  AOI21_X1   g07427(.A1(new_n4188_), .A2(new_n1746_), .B(new_n7683_), .ZN(new_n7684_));
  XOR2_X1    g07428(.A1(new_n7684_), .A2(new_n1736_), .Z(new_n7685_));
  AOI22_X1   g07429(.A1(new_n2202_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n2205_), .ZN(new_n7686_));
  OAI21_X1   g07430(.A1(new_n2495_), .A2(new_n2370_), .B(new_n7686_), .ZN(new_n7687_));
  AOI21_X1   g07431(.A1(new_n3407_), .A2(new_n2208_), .B(new_n7687_), .ZN(new_n7688_));
  XOR2_X1    g07432(.A1(new_n7688_), .A2(new_n2200_), .Z(new_n7689_));
  INV_X1     g07433(.I(new_n7689_), .ZN(new_n7690_));
  NOR3_X1    g07434(.A1(new_n7505_), .A2(new_n7500_), .A3(new_n7507_), .ZN(new_n7691_));
  INV_X1     g07435(.I(new_n7691_), .ZN(new_n7692_));
  AOI22_X1   g07436(.A1(new_n2716_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n2719_), .ZN(new_n7693_));
  OAI21_X1   g07437(.A1(new_n2027_), .A2(new_n2924_), .B(new_n7693_), .ZN(new_n7694_));
  AOI21_X1   g07438(.A1(new_n2470_), .A2(new_n2722_), .B(new_n7694_), .ZN(new_n7695_));
  XOR2_X1    g07439(.A1(new_n7695_), .A2(new_n2714_), .Z(new_n7696_));
  OAI22_X1   g07440(.A1(new_n1296_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n1432_), .ZN(new_n7697_));
  AOI21_X1   g07441(.A1(\b[15] ), .A2(new_n4053_), .B(new_n7697_), .ZN(new_n7698_));
  OAI21_X1   g07442(.A1(new_n1444_), .A2(new_n4727_), .B(new_n7698_), .ZN(new_n7699_));
  XOR2_X1    g07443(.A1(new_n7699_), .A2(\a[32] ), .Z(new_n7700_));
  OAI21_X1   g07444(.A1(new_n7394_), .A2(new_n7464_), .B(new_n7476_), .ZN(new_n7701_));
  AOI22_X1   g07445(.A1(new_n4918_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n4921_), .ZN(new_n7702_));
  OAI21_X1   g07446(.A1(new_n941_), .A2(new_n6099_), .B(new_n7702_), .ZN(new_n7703_));
  AOI21_X1   g07447(.A1(new_n1449_), .A2(new_n4699_), .B(new_n7703_), .ZN(new_n7704_));
  XOR2_X1    g07448(.A1(new_n7704_), .A2(new_n4446_), .Z(new_n7705_));
  INV_X1     g07449(.I(new_n7705_), .ZN(new_n7706_));
  AOI21_X1   g07450(.A1(new_n7455_), .A2(new_n7450_), .B(new_n7457_), .ZN(new_n7707_));
  INV_X1     g07451(.I(new_n6115_), .ZN(new_n7708_));
  AOI22_X1   g07452(.A1(new_n6108_), .A2(\b[8] ), .B1(\b[7] ), .B2(new_n6111_), .ZN(new_n7709_));
  OAI21_X1   g07453(.A1(new_n438_), .A2(new_n7708_), .B(new_n7709_), .ZN(new_n7710_));
  AOI21_X1   g07454(.A1(new_n799_), .A2(new_n6105_), .B(new_n7710_), .ZN(new_n7711_));
  XOR2_X1    g07455(.A1(new_n7711_), .A2(new_n5849_), .Z(new_n7712_));
  INV_X1     g07456(.I(new_n7712_), .ZN(new_n7713_));
  NAND2_X1   g07457(.A1(new_n7414_), .A2(new_n554_), .ZN(new_n7714_));
  AOI22_X1   g07458(.A1(new_n7403_), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n7408_), .ZN(new_n7715_));
  XOR2_X1    g07459(.A1(\a[44] ), .A2(\a[45] ), .Z(new_n7716_));
  NOR2_X1    g07460(.A1(new_n7411_), .A2(\a[44] ), .ZN(new_n7717_));
  NOR2_X1    g07461(.A1(new_n7412_), .A2(new_n6567_), .ZN(new_n7718_));
  NOR3_X1    g07462(.A1(new_n7717_), .A2(new_n7718_), .A3(new_n7716_), .ZN(new_n7719_));
  NAND2_X1   g07463(.A1(new_n7719_), .A2(\b[0] ), .ZN(new_n7720_));
  NAND3_X1   g07464(.A1(new_n7715_), .A2(new_n7720_), .A3(new_n7714_), .ZN(new_n7721_));
  XOR2_X1    g07465(.A1(new_n7721_), .A2(new_n7410_), .Z(new_n7722_));
  NOR3_X1    g07466(.A1(new_n7416_), .A2(new_n7410_), .A3(new_n7117_), .ZN(new_n7723_));
  INV_X1     g07467(.I(new_n7723_), .ZN(new_n7724_));
  NAND2_X1   g07468(.A1(new_n7722_), .A2(new_n7724_), .ZN(new_n7725_));
  OR4_X2     g07469(.A1(new_n7410_), .A2(new_n7721_), .A3(new_n7117_), .A4(new_n7416_), .Z(new_n7726_));
  NAND2_X1   g07470(.A1(new_n7725_), .A2(new_n7726_), .ZN(new_n7727_));
  INV_X1     g07471(.I(new_n6579_), .ZN(new_n7728_));
  INV_X1     g07472(.I(new_n6568_), .ZN(new_n7729_));
  NAND2_X1   g07473(.A1(new_n7729_), .A2(new_n6884_), .ZN(new_n7730_));
  INV_X1     g07474(.I(new_n6574_), .ZN(new_n7731_));
  OAI22_X1   g07475(.A1(new_n7730_), .A2(new_n377_), .B1(new_n339_), .B2(new_n7731_), .ZN(new_n7732_));
  AOI21_X1   g07476(.A1(\b[3] ), .A2(new_n6887_), .B(new_n7732_), .ZN(new_n7733_));
  OAI21_X1   g07477(.A1(new_n566_), .A2(new_n7728_), .B(new_n7733_), .ZN(new_n7734_));
  XOR2_X1    g07478(.A1(new_n7734_), .A2(new_n6567_), .Z(new_n7735_));
  NAND2_X1   g07479(.A1(new_n7735_), .A2(new_n7727_), .ZN(new_n7736_));
  INV_X1     g07480(.I(new_n7727_), .ZN(new_n7737_));
  XOR2_X1    g07481(.A1(new_n7734_), .A2(\a[44] ), .Z(new_n7738_));
  NAND2_X1   g07482(.A1(new_n7737_), .A2(new_n7738_), .ZN(new_n7739_));
  NAND2_X1   g07483(.A1(new_n7739_), .A2(new_n7736_), .ZN(new_n7740_));
  AOI21_X1   g07484(.A1(new_n7429_), .A2(new_n7426_), .B(new_n7425_), .ZN(new_n7741_));
  NOR2_X1    g07485(.A1(new_n7740_), .A2(new_n7741_), .ZN(new_n7742_));
  NOR2_X1    g07486(.A1(new_n7737_), .A2(new_n7738_), .ZN(new_n7743_));
  NOR2_X1    g07487(.A1(new_n7735_), .A2(new_n7727_), .ZN(new_n7744_));
  NOR2_X1    g07488(.A1(new_n7743_), .A2(new_n7744_), .ZN(new_n7745_));
  INV_X1     g07489(.I(new_n7741_), .ZN(new_n7746_));
  NOR2_X1    g07490(.A1(new_n7745_), .A2(new_n7746_), .ZN(new_n7747_));
  OAI21_X1   g07491(.A1(new_n7747_), .A2(new_n7742_), .B(new_n7713_), .ZN(new_n7748_));
  NAND2_X1   g07492(.A1(new_n7745_), .A2(new_n7746_), .ZN(new_n7749_));
  NAND2_X1   g07493(.A1(new_n7740_), .A2(new_n7741_), .ZN(new_n7750_));
  NAND3_X1   g07494(.A1(new_n7749_), .A2(new_n7750_), .A3(new_n7712_), .ZN(new_n7751_));
  NAND2_X1   g07495(.A1(new_n7748_), .A2(new_n7751_), .ZN(new_n7752_));
  INV_X1     g07496(.I(new_n7437_), .ZN(new_n7753_));
  OAI21_X1   g07497(.A1(new_n7431_), .A2(new_n7432_), .B(new_n7436_), .ZN(new_n7754_));
  OAI21_X1   g07498(.A1(new_n7396_), .A2(new_n7130_), .B(new_n7754_), .ZN(new_n7755_));
  NAND2_X1   g07499(.A1(new_n7755_), .A2(new_n7753_), .ZN(new_n7756_));
  NOR2_X1    g07500(.A1(new_n7756_), .A2(new_n7752_), .ZN(new_n7757_));
  AOI21_X1   g07501(.A1(new_n7749_), .A2(new_n7750_), .B(new_n7712_), .ZN(new_n7758_));
  NOR3_X1    g07502(.A1(new_n7747_), .A2(new_n7742_), .A3(new_n7713_), .ZN(new_n7759_));
  NOR2_X1    g07503(.A1(new_n7758_), .A2(new_n7759_), .ZN(new_n7760_));
  AOI21_X1   g07504(.A1(new_n7753_), .A2(new_n7755_), .B(new_n7760_), .ZN(new_n7761_));
  OAI22_X1   g07505(.A1(new_n852_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n776_), .ZN(new_n7762_));
  AOI21_X1   g07506(.A1(\b[9] ), .A2(new_n5420_), .B(new_n7762_), .ZN(new_n7763_));
  OAI21_X1   g07507(.A1(new_n859_), .A2(new_n6124_), .B(new_n7763_), .ZN(new_n7764_));
  XOR2_X1    g07508(.A1(new_n7764_), .A2(\a[38] ), .Z(new_n7765_));
  INV_X1     g07509(.I(new_n7765_), .ZN(new_n7766_));
  NOR3_X1    g07510(.A1(new_n7761_), .A2(new_n7757_), .A3(new_n7766_), .ZN(new_n7767_));
  NAND3_X1   g07511(.A1(new_n7760_), .A2(new_n7753_), .A3(new_n7755_), .ZN(new_n7768_));
  NAND2_X1   g07512(.A1(new_n7756_), .A2(new_n7752_), .ZN(new_n7769_));
  AOI21_X1   g07513(.A1(new_n7769_), .A2(new_n7768_), .B(new_n7765_), .ZN(new_n7770_));
  NOR2_X1    g07514(.A1(new_n7767_), .A2(new_n7770_), .ZN(new_n7771_));
  INV_X1     g07515(.I(new_n7771_), .ZN(new_n7772_));
  NOR2_X1    g07516(.A1(new_n7707_), .A2(new_n7772_), .ZN(new_n7773_));
  OAI21_X1   g07517(.A1(new_n7395_), .A2(new_n7456_), .B(new_n7452_), .ZN(new_n7774_));
  NOR2_X1    g07518(.A1(new_n7774_), .A2(new_n7771_), .ZN(new_n7775_));
  NOR3_X1    g07519(.A1(new_n7775_), .A2(new_n7773_), .A3(new_n7706_), .ZN(new_n7776_));
  NAND2_X1   g07520(.A1(new_n7774_), .A2(new_n7771_), .ZN(new_n7777_));
  NAND2_X1   g07521(.A1(new_n7707_), .A2(new_n7772_), .ZN(new_n7778_));
  AOI21_X1   g07522(.A1(new_n7777_), .A2(new_n7778_), .B(new_n7705_), .ZN(new_n7779_));
  NOR2_X1    g07523(.A1(new_n7779_), .A2(new_n7776_), .ZN(new_n7780_));
  NAND2_X1   g07524(.A1(new_n7701_), .A2(new_n7780_), .ZN(new_n7781_));
  NAND3_X1   g07525(.A1(new_n7474_), .A2(new_n7153_), .A3(new_n7475_), .ZN(new_n7782_));
  NAND3_X1   g07526(.A1(new_n7777_), .A2(new_n7778_), .A3(new_n7705_), .ZN(new_n7783_));
  OAI21_X1   g07527(.A1(new_n7775_), .A2(new_n7773_), .B(new_n7706_), .ZN(new_n7784_));
  NAND2_X1   g07528(.A1(new_n7784_), .A2(new_n7783_), .ZN(new_n7785_));
  NAND3_X1   g07529(.A1(new_n7785_), .A2(new_n7782_), .A3(new_n7476_), .ZN(new_n7786_));
  AOI21_X1   g07530(.A1(new_n7781_), .A2(new_n7786_), .B(new_n7700_), .ZN(new_n7787_));
  INV_X1     g07531(.I(new_n7700_), .ZN(new_n7788_));
  AOI21_X1   g07532(.A1(new_n7476_), .A2(new_n7782_), .B(new_n7785_), .ZN(new_n7789_));
  NOR2_X1    g07533(.A1(new_n7701_), .A2(new_n7780_), .ZN(new_n7790_));
  NOR3_X1    g07534(.A1(new_n7790_), .A2(new_n7789_), .A3(new_n7788_), .ZN(new_n7791_));
  NOR2_X1    g07535(.A1(new_n7791_), .A2(new_n7787_), .ZN(new_n7792_));
  AOI21_X1   g07536(.A1(new_n7471_), .A2(new_n7478_), .B(new_n7480_), .ZN(new_n7793_));
  OAI21_X1   g07537(.A1(new_n7495_), .A2(new_n7793_), .B(new_n7792_), .ZN(new_n7794_));
  OAI21_X1   g07538(.A1(new_n7790_), .A2(new_n7789_), .B(new_n7788_), .ZN(new_n7795_));
  NAND3_X1   g07539(.A1(new_n7781_), .A2(new_n7786_), .A3(new_n7700_), .ZN(new_n7796_));
  NAND2_X1   g07540(.A1(new_n7795_), .A2(new_n7796_), .ZN(new_n7797_));
  INV_X1     g07541(.I(new_n7793_), .ZN(new_n7798_));
  NAND3_X1   g07542(.A1(new_n7487_), .A2(new_n7797_), .A3(new_n7798_), .ZN(new_n7799_));
  AOI22_X1   g07543(.A1(new_n3267_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n3270_), .ZN(new_n7800_));
  OAI21_X1   g07544(.A1(new_n1553_), .A2(new_n3475_), .B(new_n7800_), .ZN(new_n7801_));
  AOI21_X1   g07545(.A1(new_n2452_), .A2(new_n3273_), .B(new_n7801_), .ZN(new_n7802_));
  XOR2_X1    g07546(.A1(new_n7802_), .A2(new_n3264_), .Z(new_n7803_));
  AOI21_X1   g07547(.A1(new_n7794_), .A2(new_n7799_), .B(new_n7803_), .ZN(new_n7804_));
  AOI21_X1   g07548(.A1(new_n7496_), .A2(new_n7486_), .B(new_n7793_), .ZN(new_n7805_));
  NOR2_X1    g07549(.A1(new_n7805_), .A2(new_n7797_), .ZN(new_n7806_));
  NOR3_X1    g07550(.A1(new_n7495_), .A2(new_n7792_), .A3(new_n7793_), .ZN(new_n7807_));
  INV_X1     g07551(.I(new_n7803_), .ZN(new_n7808_));
  NOR3_X1    g07552(.A1(new_n7807_), .A2(new_n7806_), .A3(new_n7808_), .ZN(new_n7809_));
  NOR2_X1    g07553(.A1(new_n7809_), .A2(new_n7804_), .ZN(new_n7810_));
  OAI21_X1   g07554(.A1(new_n7500_), .A2(new_n7502_), .B(new_n7810_), .ZN(new_n7811_));
  OAI21_X1   g07555(.A1(new_n7807_), .A2(new_n7806_), .B(new_n7808_), .ZN(new_n7812_));
  NAND3_X1   g07556(.A1(new_n7794_), .A2(new_n7799_), .A3(new_n7803_), .ZN(new_n7813_));
  NAND2_X1   g07557(.A1(new_n7812_), .A2(new_n7813_), .ZN(new_n7814_));
  NAND3_X1   g07558(.A1(new_n7508_), .A2(new_n7814_), .A3(new_n7493_), .ZN(new_n7815_));
  NAND3_X1   g07559(.A1(new_n7811_), .A2(new_n7815_), .A3(new_n7696_), .ZN(new_n7816_));
  INV_X1     g07560(.I(new_n7696_), .ZN(new_n7817_));
  AOI21_X1   g07561(.A1(new_n7508_), .A2(new_n7493_), .B(new_n7814_), .ZN(new_n7818_));
  NOR3_X1    g07562(.A1(new_n7500_), .A2(new_n7810_), .A3(new_n7502_), .ZN(new_n7819_));
  OAI21_X1   g07563(.A1(new_n7818_), .A2(new_n7819_), .B(new_n7817_), .ZN(new_n7820_));
  NAND2_X1   g07564(.A1(new_n7820_), .A2(new_n7816_), .ZN(new_n7821_));
  AOI21_X1   g07565(.A1(new_n7512_), .A2(new_n7692_), .B(new_n7821_), .ZN(new_n7822_));
  NOR3_X1    g07566(.A1(new_n7818_), .A2(new_n7819_), .A3(new_n7817_), .ZN(new_n7823_));
  AOI21_X1   g07567(.A1(new_n7811_), .A2(new_n7815_), .B(new_n7696_), .ZN(new_n7824_));
  NOR2_X1    g07568(.A1(new_n7823_), .A2(new_n7824_), .ZN(new_n7825_));
  NOR3_X1    g07569(.A1(new_n7523_), .A2(new_n7691_), .A3(new_n7825_), .ZN(new_n7826_));
  NOR3_X1    g07570(.A1(new_n7826_), .A2(new_n7822_), .A3(new_n7690_), .ZN(new_n7827_));
  OAI21_X1   g07571(.A1(new_n7523_), .A2(new_n7691_), .B(new_n7825_), .ZN(new_n7828_));
  NAND3_X1   g07572(.A1(new_n7512_), .A2(new_n7692_), .A3(new_n7821_), .ZN(new_n7829_));
  AOI21_X1   g07573(.A1(new_n7828_), .A2(new_n7829_), .B(new_n7689_), .ZN(new_n7830_));
  NOR2_X1    g07574(.A1(new_n7827_), .A2(new_n7830_), .ZN(new_n7831_));
  OAI21_X1   g07575(.A1(new_n7527_), .A2(new_n7529_), .B(new_n7831_), .ZN(new_n7832_));
  NAND3_X1   g07576(.A1(new_n7828_), .A2(new_n7829_), .A3(new_n7689_), .ZN(new_n7833_));
  OAI21_X1   g07577(.A1(new_n7826_), .A2(new_n7822_), .B(new_n7690_), .ZN(new_n7834_));
  NAND2_X1   g07578(.A1(new_n7834_), .A2(new_n7833_), .ZN(new_n7835_));
  NAND3_X1   g07579(.A1(new_n7535_), .A2(new_n7835_), .A3(new_n7521_), .ZN(new_n7836_));
  NAND3_X1   g07580(.A1(new_n7832_), .A2(new_n7836_), .A3(new_n7685_), .ZN(new_n7837_));
  INV_X1     g07581(.I(new_n7685_), .ZN(new_n7838_));
  AOI21_X1   g07582(.A1(new_n7535_), .A2(new_n7521_), .B(new_n7835_), .ZN(new_n7839_));
  NOR3_X1    g07583(.A1(new_n7527_), .A2(new_n7831_), .A3(new_n7529_), .ZN(new_n7840_));
  OAI21_X1   g07584(.A1(new_n7840_), .A2(new_n7839_), .B(new_n7838_), .ZN(new_n7841_));
  NAND2_X1   g07585(.A1(new_n7841_), .A2(new_n7837_), .ZN(new_n7842_));
  AOI21_X1   g07586(.A1(new_n7554_), .A2(new_n7681_), .B(new_n7842_), .ZN(new_n7843_));
  NOR3_X1    g07587(.A1(new_n7840_), .A2(new_n7839_), .A3(new_n7838_), .ZN(new_n7844_));
  AOI21_X1   g07588(.A1(new_n7832_), .A2(new_n7836_), .B(new_n7685_), .ZN(new_n7845_));
  NOR2_X1    g07589(.A1(new_n7844_), .A2(new_n7845_), .ZN(new_n7846_));
  NOR3_X1    g07590(.A1(new_n7547_), .A2(new_n7680_), .A3(new_n7846_), .ZN(new_n7847_));
  NOR3_X1    g07591(.A1(new_n7847_), .A2(new_n7679_), .A3(new_n7843_), .ZN(new_n7848_));
  OAI21_X1   g07592(.A1(new_n7547_), .A2(new_n7680_), .B(new_n7846_), .ZN(new_n7849_));
  NAND3_X1   g07593(.A1(new_n7554_), .A2(new_n7681_), .A3(new_n7842_), .ZN(new_n7850_));
  AOI21_X1   g07594(.A1(new_n7849_), .A2(new_n7850_), .B(new_n7678_), .ZN(new_n7851_));
  NOR2_X1    g07595(.A1(new_n7848_), .A2(new_n7851_), .ZN(new_n7852_));
  NAND3_X1   g07596(.A1(new_n7674_), .A2(new_n7852_), .A3(new_n7562_), .ZN(new_n7853_));
  AOI21_X1   g07597(.A1(new_n7560_), .A2(new_n7238_), .B(new_n7552_), .ZN(new_n7854_));
  NAND3_X1   g07598(.A1(new_n7849_), .A2(new_n7850_), .A3(new_n7678_), .ZN(new_n7855_));
  OAI21_X1   g07599(.A1(new_n7847_), .A2(new_n7843_), .B(new_n7679_), .ZN(new_n7856_));
  NAND2_X1   g07600(.A1(new_n7856_), .A2(new_n7855_), .ZN(new_n7857_));
  OAI21_X1   g07601(.A1(new_n7854_), .A2(new_n7556_), .B(new_n7857_), .ZN(new_n7858_));
  AOI21_X1   g07602(.A1(new_n7858_), .A2(new_n7853_), .B(new_n7673_), .ZN(new_n7859_));
  XOR2_X1    g07603(.A1(new_n7672_), .A2(new_n1002_), .Z(new_n7860_));
  NOR3_X1    g07604(.A1(new_n7854_), .A2(new_n7857_), .A3(new_n7556_), .ZN(new_n7861_));
  AOI21_X1   g07605(.A1(new_n7674_), .A2(new_n7562_), .B(new_n7852_), .ZN(new_n7862_));
  NOR3_X1    g07606(.A1(new_n7860_), .A2(new_n7862_), .A3(new_n7861_), .ZN(new_n7863_));
  NOR2_X1    g07607(.A1(new_n7859_), .A2(new_n7863_), .ZN(new_n7864_));
  AOI21_X1   g07608(.A1(new_n7558_), .A2(new_n7564_), .B(new_n7566_), .ZN(new_n7865_));
  OAI21_X1   g07609(.A1(new_n7582_), .A2(new_n7865_), .B(new_n7864_), .ZN(new_n7866_));
  OAI21_X1   g07610(.A1(new_n7861_), .A2(new_n7862_), .B(new_n7860_), .ZN(new_n7867_));
  NAND3_X1   g07611(.A1(new_n7673_), .A2(new_n7858_), .A3(new_n7853_), .ZN(new_n7868_));
  NAND2_X1   g07612(.A1(new_n7867_), .A2(new_n7868_), .ZN(new_n7869_));
  INV_X1     g07613(.I(new_n7865_), .ZN(new_n7870_));
  NAND3_X1   g07614(.A1(new_n7571_), .A2(new_n7869_), .A3(new_n7870_), .ZN(new_n7871_));
  AOI21_X1   g07615(.A1(new_n7866_), .A2(new_n7871_), .B(new_n7668_), .ZN(new_n7872_));
  XOR2_X1    g07616(.A1(new_n7667_), .A2(new_n722_), .Z(new_n7873_));
  AOI21_X1   g07617(.A1(new_n7571_), .A2(new_n7870_), .B(new_n7869_), .ZN(new_n7874_));
  NOR3_X1    g07618(.A1(new_n7582_), .A2(new_n7864_), .A3(new_n7865_), .ZN(new_n7875_));
  NOR3_X1    g07619(.A1(new_n7874_), .A2(new_n7875_), .A3(new_n7873_), .ZN(new_n7876_));
  NOR2_X1    g07620(.A1(new_n7872_), .A2(new_n7876_), .ZN(new_n7877_));
  OAI21_X1   g07621(.A1(new_n7586_), .A2(new_n7590_), .B(new_n7877_), .ZN(new_n7878_));
  OAI21_X1   g07622(.A1(new_n7874_), .A2(new_n7875_), .B(new_n7873_), .ZN(new_n7879_));
  NAND3_X1   g07623(.A1(new_n7866_), .A2(new_n7871_), .A3(new_n7668_), .ZN(new_n7880_));
  NAND2_X1   g07624(.A1(new_n7879_), .A2(new_n7880_), .ZN(new_n7881_));
  NAND3_X1   g07625(.A1(new_n7596_), .A2(new_n7881_), .A3(new_n7580_), .ZN(new_n7882_));
  NAND3_X1   g07626(.A1(new_n7878_), .A2(new_n7882_), .A3(new_n7664_), .ZN(new_n7883_));
  INV_X1     g07627(.I(new_n7659_), .ZN(new_n7884_));
  NAND3_X1   g07628(.A1(new_n7658_), .A2(new_n488_), .A3(new_n7657_), .ZN(new_n7885_));
  NAND2_X1   g07629(.A1(new_n7884_), .A2(new_n7885_), .ZN(new_n7886_));
  AOI21_X1   g07630(.A1(new_n7596_), .A2(new_n7580_), .B(new_n7881_), .ZN(new_n7887_));
  NOR3_X1    g07631(.A1(new_n7586_), .A2(new_n7590_), .A3(new_n7877_), .ZN(new_n7888_));
  OAI21_X1   g07632(.A1(new_n7888_), .A2(new_n7887_), .B(new_n7886_), .ZN(new_n7889_));
  NAND2_X1   g07633(.A1(new_n7889_), .A2(new_n7883_), .ZN(new_n7890_));
  NAND2_X1   g07634(.A1(new_n7654_), .A2(new_n7890_), .ZN(new_n7891_));
  OAI21_X1   g07635(.A1(new_n7334_), .A2(new_n7281_), .B(new_n7603_), .ZN(new_n7892_));
  NOR3_X1    g07636(.A1(new_n7888_), .A2(new_n7886_), .A3(new_n7887_), .ZN(new_n7893_));
  AOI21_X1   g07637(.A1(new_n7878_), .A2(new_n7882_), .B(new_n7664_), .ZN(new_n7894_));
  NOR2_X1    g07638(.A1(new_n7893_), .A2(new_n7894_), .ZN(new_n7895_));
  NAND3_X1   g07639(.A1(new_n7892_), .A2(new_n7604_), .A3(new_n7895_), .ZN(new_n7896_));
  NAND2_X1   g07640(.A1(new_n7891_), .A2(new_n7896_), .ZN(new_n7897_));
  INV_X1     g07641(.I(new_n7897_), .ZN(new_n7898_));
  AOI21_X1   g07642(.A1(new_n7313_), .A2(new_n7315_), .B(new_n7291_), .ZN(new_n7899_));
  NOR3_X1    g07643(.A1(new_n7611_), .A2(new_n7610_), .A3(new_n7609_), .ZN(new_n7900_));
  AOI21_X1   g07644(.A1(new_n7600_), .A2(new_n7606_), .B(new_n7332_), .ZN(new_n7901_));
  NOR2_X1    g07645(.A1(new_n7900_), .A2(new_n7901_), .ZN(new_n7902_));
  AOI21_X1   g07646(.A1(new_n7600_), .A2(new_n7606_), .B(new_n7609_), .ZN(new_n7903_));
  INV_X1     g07647(.I(new_n7903_), .ZN(new_n7904_));
  OAI21_X1   g07648(.A1(new_n7902_), .A2(new_n7899_), .B(new_n7904_), .ZN(new_n7905_));
  XOR2_X1    g07649(.A1(new_n7080_), .A2(new_n7077_), .Z(new_n7906_));
  AOI22_X1   g07650(.A1(new_n800_), .A2(\b[43] ), .B1(\b[44] ), .B2(new_n333_), .ZN(new_n7907_));
  OAI21_X1   g07651(.A1(new_n6490_), .A2(new_n392_), .B(new_n7907_), .ZN(new_n7908_));
  AOI21_X1   g07652(.A1(new_n7906_), .A2(new_n330_), .B(new_n7908_), .ZN(new_n7909_));
  XOR2_X1    g07653(.A1(new_n7909_), .A2(new_n312_), .Z(new_n7910_));
  NAND2_X1   g07654(.A1(new_n7905_), .A2(new_n7910_), .ZN(new_n7911_));
  AOI21_X1   g07655(.A1(new_n7613_), .A2(new_n7324_), .B(new_n7903_), .ZN(new_n7912_));
  INV_X1     g07656(.I(new_n7910_), .ZN(new_n7913_));
  NAND2_X1   g07657(.A1(new_n7912_), .A2(new_n7913_), .ZN(new_n7914_));
  NAND3_X1   g07658(.A1(new_n7911_), .A2(new_n7914_), .A3(new_n7898_), .ZN(new_n7915_));
  AOI21_X1   g07659(.A1(new_n7911_), .A2(new_n7914_), .B(new_n7898_), .ZN(new_n7916_));
  INV_X1     g07660(.I(new_n7916_), .ZN(new_n7917_));
  AOI21_X1   g07661(.A1(new_n7917_), .A2(new_n7915_), .B(new_n7652_), .ZN(new_n7918_));
  INV_X1     g07662(.I(new_n7915_), .ZN(new_n7919_));
  NOR3_X1    g07663(.A1(new_n7919_), .A2(new_n7651_), .A3(new_n7916_), .ZN(new_n7920_));
  NOR2_X1    g07664(.A1(new_n7918_), .A2(new_n7920_), .ZN(new_n7921_));
  XOR2_X1    g07665(.A1(new_n7640_), .A2(new_n7921_), .Z(\f[47] ));
  OAI21_X1   g07666(.A1(new_n7912_), .A2(new_n7913_), .B(new_n7897_), .ZN(new_n7923_));
  NAND2_X1   g07667(.A1(new_n7923_), .A2(new_n7914_), .ZN(new_n7924_));
  NAND2_X1   g07668(.A1(new_n7101_), .A2(new_n7100_), .ZN(new_n7925_));
  INV_X1     g07669(.I(new_n7925_), .ZN(new_n7926_));
  AOI22_X1   g07670(.A1(new_n800_), .A2(\b[44] ), .B1(\b[45] ), .B2(new_n333_), .ZN(new_n7927_));
  OAI21_X1   g07671(.A1(new_n6775_), .A2(new_n392_), .B(new_n7927_), .ZN(new_n7928_));
  AOI21_X1   g07672(.A1(new_n7926_), .A2(new_n330_), .B(new_n7928_), .ZN(new_n7929_));
  XOR2_X1    g07673(.A1(new_n7929_), .A2(\a[5] ), .Z(new_n7930_));
  NAND2_X1   g07674(.A1(new_n7719_), .A2(\b[1] ), .ZN(new_n7931_));
  AOI22_X1   g07675(.A1(new_n7403_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n7408_), .ZN(new_n7932_));
  NAND2_X1   g07676(.A1(new_n299_), .A2(new_n7414_), .ZN(new_n7933_));
  NAND3_X1   g07677(.A1(new_n7933_), .A2(new_n7932_), .A3(new_n7931_), .ZN(new_n7934_));
  XOR2_X1    g07678(.A1(new_n7934_), .A2(new_n7410_), .Z(new_n7935_));
  XNOR2_X1   g07679(.A1(\a[47] ), .A2(\a[48] ), .ZN(new_n7936_));
  NOR2_X1    g07680(.A1(new_n7936_), .A2(new_n258_), .ZN(new_n7937_));
  INV_X1     g07681(.I(new_n7937_), .ZN(new_n7938_));
  NAND2_X1   g07682(.A1(new_n7935_), .A2(new_n7938_), .ZN(new_n7939_));
  XOR2_X1    g07683(.A1(new_n7934_), .A2(\a[47] ), .Z(new_n7940_));
  NAND2_X1   g07684(.A1(new_n7940_), .A2(new_n7937_), .ZN(new_n7941_));
  NAND2_X1   g07685(.A1(new_n7939_), .A2(new_n7941_), .ZN(new_n7942_));
  XOR2_X1    g07686(.A1(new_n7942_), .A2(new_n7726_), .Z(new_n7943_));
  OAI22_X1   g07687(.A1(new_n7730_), .A2(new_n438_), .B1(new_n377_), .B2(new_n7731_), .ZN(new_n7944_));
  AOI21_X1   g07688(.A1(\b[4] ), .A2(new_n6887_), .B(new_n7944_), .ZN(new_n7945_));
  OAI21_X1   g07689(.A1(new_n450_), .A2(new_n7728_), .B(new_n7945_), .ZN(new_n7946_));
  XOR2_X1    g07690(.A1(new_n7946_), .A2(\a[44] ), .Z(new_n7947_));
  INV_X1     g07691(.I(new_n7947_), .ZN(new_n7948_));
  OAI21_X1   g07692(.A1(new_n7741_), .A2(new_n7743_), .B(new_n7739_), .ZN(new_n7949_));
  XOR2_X1    g07693(.A1(new_n7949_), .A2(new_n7948_), .Z(new_n7950_));
  XOR2_X1    g07694(.A1(new_n7950_), .A2(new_n7943_), .Z(new_n7951_));
  AOI22_X1   g07695(.A1(new_n6108_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n6111_), .ZN(new_n7952_));
  OAI21_X1   g07696(.A1(new_n471_), .A2(new_n7708_), .B(new_n7952_), .ZN(new_n7953_));
  AOI21_X1   g07697(.A1(new_n676_), .A2(new_n6105_), .B(new_n7953_), .ZN(new_n7954_));
  XOR2_X1    g07698(.A1(new_n7954_), .A2(new_n5849_), .Z(new_n7955_));
  NAND2_X1   g07699(.A1(new_n7768_), .A2(new_n7751_), .ZN(new_n7956_));
  NAND2_X1   g07700(.A1(new_n7956_), .A2(new_n7955_), .ZN(new_n7957_));
  INV_X1     g07701(.I(new_n7955_), .ZN(new_n7958_));
  NOR2_X1    g07702(.A1(new_n7757_), .A2(new_n7759_), .ZN(new_n7959_));
  NAND2_X1   g07703(.A1(new_n7959_), .A2(new_n7958_), .ZN(new_n7960_));
  NAND3_X1   g07704(.A1(new_n7960_), .A2(new_n7957_), .A3(new_n7951_), .ZN(new_n7961_));
  XNOR2_X1   g07705(.A1(new_n7950_), .A2(new_n7943_), .ZN(new_n7962_));
  NOR2_X1    g07706(.A1(new_n7959_), .A2(new_n7958_), .ZN(new_n7963_));
  NOR2_X1    g07707(.A1(new_n7956_), .A2(new_n7955_), .ZN(new_n7964_));
  OAI21_X1   g07708(.A1(new_n7963_), .A2(new_n7964_), .B(new_n7962_), .ZN(new_n7965_));
  NAND2_X1   g07709(.A1(new_n7965_), .A2(new_n7961_), .ZN(new_n7966_));
  AOI22_X1   g07710(.A1(new_n5155_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n5160_), .ZN(new_n7967_));
  OAI21_X1   g07711(.A1(new_n776_), .A2(new_n6877_), .B(new_n7967_), .ZN(new_n7968_));
  AOI21_X1   g07712(.A1(new_n1194_), .A2(new_n5166_), .B(new_n7968_), .ZN(new_n7969_));
  XOR2_X1    g07713(.A1(new_n7969_), .A2(new_n5162_), .Z(new_n7970_));
  INV_X1     g07714(.I(new_n7970_), .ZN(new_n7971_));
  AOI21_X1   g07715(.A1(new_n7774_), .A2(new_n7771_), .B(new_n7767_), .ZN(new_n7972_));
  NOR2_X1    g07716(.A1(new_n7972_), .A2(new_n7971_), .ZN(new_n7973_));
  INV_X1     g07717(.I(new_n7767_), .ZN(new_n7974_));
  OAI21_X1   g07718(.A1(new_n7707_), .A2(new_n7772_), .B(new_n7974_), .ZN(new_n7975_));
  NOR2_X1    g07719(.A1(new_n7975_), .A2(new_n7970_), .ZN(new_n7976_));
  NOR3_X1    g07720(.A1(new_n7973_), .A2(new_n7976_), .A3(new_n7966_), .ZN(new_n7977_));
  NOR3_X1    g07721(.A1(new_n7963_), .A2(new_n7964_), .A3(new_n7962_), .ZN(new_n7978_));
  AOI21_X1   g07722(.A1(new_n7960_), .A2(new_n7957_), .B(new_n7951_), .ZN(new_n7979_));
  NOR2_X1    g07723(.A1(new_n7978_), .A2(new_n7979_), .ZN(new_n7980_));
  NAND2_X1   g07724(.A1(new_n7975_), .A2(new_n7970_), .ZN(new_n7981_));
  NAND2_X1   g07725(.A1(new_n7972_), .A2(new_n7971_), .ZN(new_n7982_));
  AOI21_X1   g07726(.A1(new_n7982_), .A2(new_n7981_), .B(new_n7980_), .ZN(new_n7983_));
  NOR2_X1    g07727(.A1(new_n7983_), .A2(new_n7977_), .ZN(new_n7984_));
  OAI22_X1   g07728(.A1(new_n1268_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n1093_), .ZN(new_n7985_));
  AOI21_X1   g07729(.A1(\b[13] ), .A2(new_n4706_), .B(new_n7985_), .ZN(new_n7986_));
  OAI21_X1   g07730(.A1(new_n1275_), .A2(new_n4458_), .B(new_n7986_), .ZN(new_n7987_));
  XOR2_X1    g07731(.A1(new_n7987_), .A2(\a[35] ), .Z(new_n7988_));
  OAI21_X1   g07732(.A1(new_n7789_), .A2(new_n7776_), .B(new_n7988_), .ZN(new_n7989_));
  INV_X1     g07733(.I(new_n7988_), .ZN(new_n7990_));
  AOI21_X1   g07734(.A1(new_n7701_), .A2(new_n7780_), .B(new_n7776_), .ZN(new_n7991_));
  NAND2_X1   g07735(.A1(new_n7991_), .A2(new_n7990_), .ZN(new_n7992_));
  NAND3_X1   g07736(.A1(new_n7992_), .A2(new_n7989_), .A3(new_n7984_), .ZN(new_n7993_));
  OR2_X2     g07737(.A1(new_n7983_), .A2(new_n7977_), .Z(new_n7994_));
  NOR2_X1    g07738(.A1(new_n7991_), .A2(new_n7990_), .ZN(new_n7995_));
  NOR3_X1    g07739(.A1(new_n7789_), .A2(new_n7776_), .A3(new_n7988_), .ZN(new_n7996_));
  OAI21_X1   g07740(.A1(new_n7995_), .A2(new_n7996_), .B(new_n7994_), .ZN(new_n7997_));
  NAND2_X1   g07741(.A1(new_n7997_), .A2(new_n7993_), .ZN(new_n7998_));
  INV_X1     g07742(.I(new_n7998_), .ZN(new_n7999_));
  AOI22_X1   g07743(.A1(new_n3864_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n3869_), .ZN(new_n8000_));
  OAI21_X1   g07744(.A1(new_n1296_), .A2(new_n5410_), .B(new_n8000_), .ZN(new_n8001_));
  AOI21_X1   g07745(.A1(new_n2038_), .A2(new_n3872_), .B(new_n8001_), .ZN(new_n8002_));
  XOR2_X1    g07746(.A1(new_n8002_), .A2(new_n3876_), .Z(new_n8003_));
  OAI21_X1   g07747(.A1(new_n7805_), .A2(new_n7797_), .B(new_n7796_), .ZN(new_n8004_));
  NAND2_X1   g07748(.A1(new_n8004_), .A2(new_n8003_), .ZN(new_n8005_));
  INV_X1     g07749(.I(new_n8003_), .ZN(new_n8006_));
  NAND2_X1   g07750(.A1(new_n7487_), .A2(new_n7798_), .ZN(new_n8007_));
  AOI21_X1   g07751(.A1(new_n8007_), .A2(new_n7792_), .B(new_n7791_), .ZN(new_n8008_));
  NAND2_X1   g07752(.A1(new_n8008_), .A2(new_n8006_), .ZN(new_n8009_));
  NAND3_X1   g07753(.A1(new_n8009_), .A2(new_n7999_), .A3(new_n8005_), .ZN(new_n8010_));
  INV_X1     g07754(.I(new_n8005_), .ZN(new_n8011_));
  NOR2_X1    g07755(.A1(new_n8004_), .A2(new_n8003_), .ZN(new_n8012_));
  OAI21_X1   g07756(.A1(new_n8011_), .A2(new_n8012_), .B(new_n7998_), .ZN(new_n8013_));
  AND2_X2    g07757(.A1(new_n8013_), .A2(new_n8010_), .Z(new_n8014_));
  AOI22_X1   g07758(.A1(new_n3267_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n3270_), .ZN(new_n8015_));
  OAI21_X1   g07759(.A1(new_n1859_), .A2(new_n3475_), .B(new_n8015_), .ZN(new_n8016_));
  AOI21_X1   g07760(.A1(new_n2032_), .A2(new_n3273_), .B(new_n8016_), .ZN(new_n8017_));
  XOR2_X1    g07761(.A1(new_n8017_), .A2(new_n3264_), .Z(new_n8018_));
  OAI21_X1   g07762(.A1(new_n7818_), .A2(new_n7809_), .B(new_n8018_), .ZN(new_n8019_));
  NOR3_X1    g07763(.A1(new_n7818_), .A2(new_n7809_), .A3(new_n8018_), .ZN(new_n8020_));
  INV_X1     g07764(.I(new_n8020_), .ZN(new_n8021_));
  NAND3_X1   g07765(.A1(new_n8021_), .A2(new_n8014_), .A3(new_n8019_), .ZN(new_n8022_));
  NAND2_X1   g07766(.A1(new_n8013_), .A2(new_n8010_), .ZN(new_n8023_));
  INV_X1     g07767(.I(new_n8019_), .ZN(new_n8024_));
  OAI21_X1   g07768(.A1(new_n8024_), .A2(new_n8020_), .B(new_n8023_), .ZN(new_n8025_));
  NAND2_X1   g07769(.A1(new_n8025_), .A2(new_n8022_), .ZN(new_n8026_));
  AOI22_X1   g07770(.A1(new_n2716_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n2719_), .ZN(new_n8027_));
  OAI21_X1   g07771(.A1(new_n2142_), .A2(new_n2924_), .B(new_n8027_), .ZN(new_n8028_));
  AOI21_X1   g07772(.A1(new_n3033_), .A2(new_n2722_), .B(new_n8028_), .ZN(new_n8029_));
  XOR2_X1    g07773(.A1(new_n8029_), .A2(new_n2714_), .Z(new_n8030_));
  INV_X1     g07774(.I(new_n8030_), .ZN(new_n8031_));
  AOI21_X1   g07775(.A1(new_n7828_), .A2(new_n7816_), .B(new_n8031_), .ZN(new_n8032_));
  NOR3_X1    g07776(.A1(new_n7822_), .A2(new_n7823_), .A3(new_n8030_), .ZN(new_n8033_));
  NOR3_X1    g07777(.A1(new_n8032_), .A2(new_n8033_), .A3(new_n8026_), .ZN(new_n8034_));
  INV_X1     g07778(.I(new_n8026_), .ZN(new_n8035_));
  OAI21_X1   g07779(.A1(new_n7822_), .A2(new_n7823_), .B(new_n8030_), .ZN(new_n8036_));
  NAND3_X1   g07780(.A1(new_n7828_), .A2(new_n7816_), .A3(new_n8031_), .ZN(new_n8037_));
  AOI21_X1   g07781(.A1(new_n8036_), .A2(new_n8037_), .B(new_n8035_), .ZN(new_n8038_));
  NOR2_X1    g07782(.A1(new_n8038_), .A2(new_n8034_), .ZN(new_n8039_));
  INV_X1     g07783(.I(new_n8039_), .ZN(new_n8040_));
  OAI22_X1   g07784(.A1(new_n2189_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n2194_), .ZN(new_n8041_));
  AOI21_X1   g07785(.A1(\b[25] ), .A2(new_n2361_), .B(new_n8041_), .ZN(new_n8042_));
  OAI21_X1   g07786(.A1(new_n3165_), .A2(new_n2197_), .B(new_n8042_), .ZN(new_n8043_));
  XOR2_X1    g07787(.A1(new_n8043_), .A2(\a[23] ), .Z(new_n8044_));
  INV_X1     g07788(.I(new_n8044_), .ZN(new_n8045_));
  AOI21_X1   g07789(.A1(new_n7832_), .A2(new_n7833_), .B(new_n8045_), .ZN(new_n8046_));
  NOR3_X1    g07790(.A1(new_n7839_), .A2(new_n7827_), .A3(new_n8044_), .ZN(new_n8047_));
  NOR3_X1    g07791(.A1(new_n8046_), .A2(new_n8047_), .A3(new_n8040_), .ZN(new_n8048_));
  OAI21_X1   g07792(.A1(new_n7839_), .A2(new_n7827_), .B(new_n8044_), .ZN(new_n8049_));
  NAND3_X1   g07793(.A1(new_n7832_), .A2(new_n7833_), .A3(new_n8045_), .ZN(new_n8050_));
  AOI21_X1   g07794(.A1(new_n8050_), .A2(new_n8049_), .B(new_n8039_), .ZN(new_n8051_));
  NOR2_X1    g07795(.A1(new_n8051_), .A2(new_n8048_), .ZN(new_n8052_));
  INV_X1     g07796(.I(new_n8052_), .ZN(new_n8053_));
  AOI22_X1   g07797(.A1(new_n1738_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n1743_), .ZN(new_n8054_));
  OAI21_X1   g07798(.A1(new_n3185_), .A2(new_n1931_), .B(new_n8054_), .ZN(new_n8055_));
  AOI21_X1   g07799(.A1(new_n4230_), .A2(new_n1746_), .B(new_n8055_), .ZN(new_n8056_));
  XOR2_X1    g07800(.A1(new_n8056_), .A2(new_n1736_), .Z(new_n8057_));
  INV_X1     g07801(.I(new_n8057_), .ZN(new_n8058_));
  AOI21_X1   g07802(.A1(new_n7849_), .A2(new_n7837_), .B(new_n8058_), .ZN(new_n8059_));
  NOR3_X1    g07803(.A1(new_n7843_), .A2(new_n7844_), .A3(new_n8057_), .ZN(new_n8060_));
  NOR3_X1    g07804(.A1(new_n8059_), .A2(new_n8060_), .A3(new_n8053_), .ZN(new_n8061_));
  OAI21_X1   g07805(.A1(new_n7843_), .A2(new_n7844_), .B(new_n8057_), .ZN(new_n8062_));
  NAND3_X1   g07806(.A1(new_n7849_), .A2(new_n7837_), .A3(new_n8058_), .ZN(new_n8063_));
  AOI21_X1   g07807(.A1(new_n8063_), .A2(new_n8062_), .B(new_n8052_), .ZN(new_n8064_));
  NOR2_X1    g07808(.A1(new_n8061_), .A2(new_n8064_), .ZN(new_n8065_));
  OAI22_X1   g07809(.A1(new_n1592_), .A2(new_n4638_), .B1(new_n4023_), .B2(new_n1505_), .ZN(new_n8066_));
  AOI21_X1   g07810(.A1(\b[31] ), .A2(new_n1584_), .B(new_n8066_), .ZN(new_n8067_));
  OAI21_X1   g07811(.A1(new_n6451_), .A2(new_n1732_), .B(new_n8067_), .ZN(new_n8068_));
  XOR2_X1    g07812(.A1(new_n8068_), .A2(\a[17] ), .Z(new_n8069_));
  INV_X1     g07813(.I(new_n8069_), .ZN(new_n8070_));
  AOI21_X1   g07814(.A1(new_n7853_), .A2(new_n7855_), .B(new_n8070_), .ZN(new_n8071_));
  NOR3_X1    g07815(.A1(new_n7861_), .A2(new_n7848_), .A3(new_n8069_), .ZN(new_n8072_));
  NOR2_X1    g07816(.A1(new_n8072_), .A2(new_n8071_), .ZN(new_n8073_));
  NAND2_X1   g07817(.A1(new_n8073_), .A2(new_n8065_), .ZN(new_n8074_));
  INV_X1     g07818(.I(new_n8065_), .ZN(new_n8075_));
  OAI21_X1   g07819(.A1(new_n7861_), .A2(new_n7848_), .B(new_n8069_), .ZN(new_n8076_));
  NAND3_X1   g07820(.A1(new_n7853_), .A2(new_n7855_), .A3(new_n8070_), .ZN(new_n8077_));
  NAND2_X1   g07821(.A1(new_n8076_), .A2(new_n8077_), .ZN(new_n8078_));
  NAND2_X1   g07822(.A1(new_n8078_), .A2(new_n8075_), .ZN(new_n8079_));
  NAND2_X1   g07823(.A1(new_n8074_), .A2(new_n8079_), .ZN(new_n8080_));
  OAI22_X1   g07824(.A1(new_n993_), .A2(new_n4886_), .B1(new_n4666_), .B2(new_n997_), .ZN(new_n8081_));
  AOI21_X1   g07825(.A1(\b[34] ), .A2(new_n1486_), .B(new_n8081_), .ZN(new_n8082_));
  OAI21_X1   g07826(.A1(new_n4898_), .A2(new_n1323_), .B(new_n8082_), .ZN(new_n8083_));
  XOR2_X1    g07827(.A1(new_n8083_), .A2(\a[14] ), .Z(new_n8084_));
  INV_X1     g07828(.I(new_n8084_), .ZN(new_n8085_));
  AOI21_X1   g07829(.A1(new_n7866_), .A2(new_n7868_), .B(new_n8085_), .ZN(new_n8086_));
  NOR3_X1    g07830(.A1(new_n7874_), .A2(new_n7863_), .A3(new_n8084_), .ZN(new_n8087_));
  NOR3_X1    g07831(.A1(new_n8086_), .A2(new_n8087_), .A3(new_n8080_), .ZN(new_n8088_));
  NOR2_X1    g07832(.A1(new_n8078_), .A2(new_n8075_), .ZN(new_n8089_));
  NOR2_X1    g07833(.A1(new_n8073_), .A2(new_n8065_), .ZN(new_n8090_));
  NOR2_X1    g07834(.A1(new_n8090_), .A2(new_n8089_), .ZN(new_n8091_));
  OAI21_X1   g07835(.A1(new_n7874_), .A2(new_n7863_), .B(new_n8084_), .ZN(new_n8092_));
  NAND3_X1   g07836(.A1(new_n7866_), .A2(new_n7868_), .A3(new_n8085_), .ZN(new_n8093_));
  AOI21_X1   g07837(.A1(new_n8093_), .A2(new_n8092_), .B(new_n8091_), .ZN(new_n8094_));
  NOR2_X1    g07838(.A1(new_n8094_), .A2(new_n8088_), .ZN(new_n8095_));
  OAI22_X1   g07839(.A1(new_n713_), .A2(new_n5761_), .B1(new_n5341_), .B2(new_n717_), .ZN(new_n8096_));
  AOI21_X1   g07840(.A1(\b[37] ), .A2(new_n1126_), .B(new_n8096_), .ZN(new_n8097_));
  OAI21_X1   g07841(.A1(new_n6309_), .A2(new_n986_), .B(new_n8097_), .ZN(new_n8098_));
  XOR2_X1    g07842(.A1(new_n8098_), .A2(\a[11] ), .Z(new_n8099_));
  OAI21_X1   g07843(.A1(new_n7887_), .A2(new_n7876_), .B(new_n8099_), .ZN(new_n8100_));
  INV_X1     g07844(.I(new_n8099_), .ZN(new_n8101_));
  NAND3_X1   g07845(.A1(new_n7878_), .A2(new_n7880_), .A3(new_n8101_), .ZN(new_n8102_));
  NAND3_X1   g07846(.A1(new_n8102_), .A2(new_n8100_), .A3(new_n8095_), .ZN(new_n8103_));
  INV_X1     g07847(.I(new_n8095_), .ZN(new_n8104_));
  AOI21_X1   g07848(.A1(new_n7878_), .A2(new_n7880_), .B(new_n8101_), .ZN(new_n8105_));
  NOR3_X1    g07849(.A1(new_n7887_), .A2(new_n7876_), .A3(new_n8099_), .ZN(new_n8106_));
  OAI21_X1   g07850(.A1(new_n8105_), .A2(new_n8106_), .B(new_n8104_), .ZN(new_n8107_));
  NAND2_X1   g07851(.A1(new_n8107_), .A2(new_n8103_), .ZN(new_n8108_));
  INV_X1     g07852(.I(new_n8108_), .ZN(new_n8109_));
  AOI21_X1   g07853(.A1(new_n7602_), .A2(new_n7285_), .B(new_n7594_), .ZN(new_n8110_));
  NOR3_X1    g07854(.A1(new_n8110_), .A2(new_n7598_), .A3(new_n7890_), .ZN(new_n8111_));
  AOI22_X1   g07855(.A1(new_n518_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n636_), .ZN(new_n8112_));
  OAI21_X1   g07856(.A1(new_n6284_), .A2(new_n917_), .B(new_n8112_), .ZN(new_n8113_));
  AOI21_X1   g07857(.A1(new_n7106_), .A2(new_n618_), .B(new_n8113_), .ZN(new_n8114_));
  XOR2_X1    g07858(.A1(new_n8114_), .A2(new_n488_), .Z(new_n8115_));
  OAI21_X1   g07859(.A1(new_n8111_), .A2(new_n7893_), .B(new_n8115_), .ZN(new_n8116_));
  INV_X1     g07860(.I(new_n8115_), .ZN(new_n8117_));
  NAND3_X1   g07861(.A1(new_n7896_), .A2(new_n7883_), .A3(new_n8117_), .ZN(new_n8118_));
  NAND3_X1   g07862(.A1(new_n8116_), .A2(new_n8118_), .A3(new_n8109_), .ZN(new_n8119_));
  INV_X1     g07863(.I(new_n8119_), .ZN(new_n8120_));
  AOI21_X1   g07864(.A1(new_n8116_), .A2(new_n8118_), .B(new_n8109_), .ZN(new_n8121_));
  OAI21_X1   g07865(.A1(new_n8120_), .A2(new_n8121_), .B(new_n7930_), .ZN(new_n8122_));
  XOR2_X1    g07866(.A1(new_n7929_), .A2(new_n312_), .Z(new_n8123_));
  INV_X1     g07867(.I(new_n8121_), .ZN(new_n8124_));
  NAND3_X1   g07868(.A1(new_n8124_), .A2(new_n8119_), .A3(new_n8123_), .ZN(new_n8125_));
  INV_X1     g07869(.I(\b[47] ), .ZN(new_n8126_));
  INV_X1     g07870(.I(\b[48] ), .ZN(new_n8127_));
  OAI22_X1   g07871(.A1(new_n277_), .A2(new_n8127_), .B1(new_n8126_), .B2(new_n262_), .ZN(new_n8128_));
  AOI21_X1   g07872(.A1(\b[46] ), .A2(new_n283_), .B(new_n8128_), .ZN(new_n8129_));
  XOR2_X1    g07873(.A1(\b[47] ), .A2(\b[48] ), .Z(new_n8130_));
  NOR3_X1    g07874(.A1(new_n7620_), .A2(new_n7621_), .A3(new_n7096_), .ZN(new_n8131_));
  OAI21_X1   g07875(.A1(new_n8131_), .A2(\b[46] ), .B(\b[47] ), .ZN(new_n8132_));
  NAND2_X1   g07876(.A1(new_n7643_), .A2(\b[46] ), .ZN(new_n8133_));
  AOI21_X1   g07877(.A1(new_n8132_), .A2(new_n8133_), .B(new_n8130_), .ZN(new_n8134_));
  INV_X1     g07878(.I(new_n8130_), .ZN(new_n8135_));
  NAND2_X1   g07879(.A1(new_n8132_), .A2(new_n8133_), .ZN(new_n8136_));
  NOR2_X1    g07880(.A1(new_n8136_), .A2(new_n8135_), .ZN(new_n8137_));
  NOR2_X1    g07881(.A1(new_n8137_), .A2(new_n8134_), .ZN(new_n8138_));
  OAI21_X1   g07882(.A1(new_n8138_), .A2(new_n279_), .B(new_n8129_), .ZN(new_n8139_));
  XOR2_X1    g07883(.A1(new_n8139_), .A2(\a[2] ), .Z(new_n8140_));
  INV_X1     g07884(.I(new_n8140_), .ZN(new_n8141_));
  NAND3_X1   g07885(.A1(new_n8141_), .A2(new_n8125_), .A3(new_n8122_), .ZN(new_n8142_));
  INV_X1     g07886(.I(new_n8122_), .ZN(new_n8143_));
  NOR3_X1    g07887(.A1(new_n8120_), .A2(new_n8121_), .A3(new_n7930_), .ZN(new_n8144_));
  OAI21_X1   g07888(.A1(new_n8143_), .A2(new_n8144_), .B(new_n8140_), .ZN(new_n8145_));
  AOI21_X1   g07889(.A1(new_n8145_), .A2(new_n8142_), .B(new_n7924_), .ZN(new_n8146_));
  NOR2_X1    g07890(.A1(new_n7905_), .A2(new_n7910_), .ZN(new_n8147_));
  AOI21_X1   g07891(.A1(new_n7905_), .A2(new_n7910_), .B(new_n7898_), .ZN(new_n8148_));
  NOR2_X1    g07892(.A1(new_n8148_), .A2(new_n8147_), .ZN(new_n8149_));
  NOR3_X1    g07893(.A1(new_n8143_), .A2(new_n8144_), .A3(new_n8140_), .ZN(new_n8150_));
  AOI21_X1   g07894(.A1(new_n8122_), .A2(new_n8125_), .B(new_n8141_), .ZN(new_n8151_));
  NOR3_X1    g07895(.A1(new_n8150_), .A2(new_n8151_), .A3(new_n8149_), .ZN(new_n8152_));
  NOR2_X1    g07896(.A1(new_n8152_), .A2(new_n8146_), .ZN(new_n8153_));
  INV_X1     g07897(.I(new_n8153_), .ZN(new_n8154_));
  NOR3_X1    g07898(.A1(new_n7919_), .A2(new_n7652_), .A3(new_n7916_), .ZN(new_n8155_));
  INV_X1     g07899(.I(new_n8155_), .ZN(new_n8156_));
  OAI21_X1   g07900(.A1(new_n7640_), .A2(new_n7921_), .B(new_n8156_), .ZN(new_n8157_));
  XOR2_X1    g07901(.A1(new_n8157_), .A2(new_n8154_), .Z(\f[48] ));
  OAI21_X1   g07902(.A1(new_n8143_), .A2(new_n8144_), .B(new_n7924_), .ZN(new_n8159_));
  NAND3_X1   g07903(.A1(new_n8149_), .A2(new_n8122_), .A3(new_n8125_), .ZN(new_n8160_));
  AOI21_X1   g07904(.A1(new_n8159_), .A2(new_n8160_), .B(new_n8141_), .ZN(new_n8161_));
  AOI21_X1   g07905(.A1(new_n8157_), .A2(new_n8154_), .B(new_n8161_), .ZN(new_n8162_));
  AOI22_X1   g07906(.A1(new_n267_), .A2(\b[49] ), .B1(\b[48] ), .B2(new_n261_), .ZN(new_n8163_));
  OAI21_X1   g07907(.A1(new_n8126_), .A2(new_n284_), .B(new_n8163_), .ZN(new_n8164_));
  INV_X1     g07908(.I(new_n8164_), .ZN(new_n8165_));
  AOI21_X1   g07909(.A1(new_n8136_), .A2(\b[48] ), .B(new_n8126_), .ZN(new_n8166_));
  NOR2_X1    g07910(.A1(new_n8136_), .A2(\b[48] ), .ZN(new_n8167_));
  INV_X1     g07911(.I(\b[49] ), .ZN(new_n8168_));
  NAND3_X1   g07912(.A1(new_n8132_), .A2(new_n8133_), .A3(new_n8168_), .ZN(new_n8169_));
  NAND2_X1   g07913(.A1(new_n8136_), .A2(\b[49] ), .ZN(new_n8170_));
  NAND2_X1   g07914(.A1(new_n8170_), .A2(new_n8169_), .ZN(new_n8171_));
  OAI21_X1   g07915(.A1(new_n8166_), .A2(new_n8167_), .B(new_n8171_), .ZN(new_n8172_));
  OR3_X2     g07916(.A1(new_n8171_), .A2(new_n8166_), .A3(new_n8167_), .Z(new_n8173_));
  NAND3_X1   g07917(.A1(new_n8173_), .A2(new_n265_), .A3(new_n8172_), .ZN(new_n8174_));
  AOI21_X1   g07918(.A1(new_n8174_), .A2(new_n8165_), .B(new_n270_), .ZN(new_n8175_));
  AND3_X2    g07919(.A1(new_n8174_), .A2(new_n270_), .A3(new_n8165_), .Z(new_n8176_));
  NOR2_X1    g07920(.A1(new_n8176_), .A2(new_n8175_), .ZN(new_n8177_));
  OAI21_X1   g07921(.A1(new_n8120_), .A2(new_n8121_), .B(new_n8123_), .ZN(new_n8178_));
  NOR3_X1    g07922(.A1(new_n8120_), .A2(new_n8121_), .A3(new_n8123_), .ZN(new_n8179_));
  OAI21_X1   g07923(.A1(new_n7924_), .A2(new_n8179_), .B(new_n8178_), .ZN(new_n8180_));
  NAND2_X1   g07924(.A1(new_n8177_), .A2(new_n8180_), .ZN(new_n8181_));
  INV_X1     g07925(.I(new_n8181_), .ZN(new_n8182_));
  NOR2_X1    g07926(.A1(new_n8177_), .A2(new_n8180_), .ZN(new_n8183_));
  AOI22_X1   g07927(.A1(new_n800_), .A2(\b[45] ), .B1(\b[46] ), .B2(new_n333_), .ZN(new_n8184_));
  OAI21_X1   g07928(.A1(new_n7074_), .A2(new_n392_), .B(new_n8184_), .ZN(new_n8185_));
  INV_X1     g07929(.I(new_n8185_), .ZN(new_n8186_));
  OAI21_X1   g07930(.A1(new_n7627_), .A2(new_n318_), .B(new_n8186_), .ZN(new_n8187_));
  XOR2_X1    g07931(.A1(new_n8187_), .A2(\a[5] ), .Z(new_n8188_));
  AOI22_X1   g07932(.A1(new_n518_), .A2(\b[43] ), .B1(\b[42] ), .B2(new_n636_), .ZN(new_n8189_));
  OAI21_X1   g07933(.A1(new_n6285_), .A2(new_n917_), .B(new_n8189_), .ZN(new_n8190_));
  INV_X1     g07934(.I(new_n8190_), .ZN(new_n8191_));
  NAND3_X1   g07935(.A1(new_n6782_), .A2(new_n6784_), .A3(new_n618_), .ZN(new_n8192_));
  NAND2_X1   g07936(.A1(new_n8192_), .A2(new_n8191_), .ZN(new_n8193_));
  XOR2_X1    g07937(.A1(new_n8193_), .A2(\a[8] ), .Z(new_n8194_));
  NOR2_X1    g07938(.A1(new_n6750_), .A2(new_n5790_), .ZN(new_n8195_));
  OAI22_X1   g07939(.A1(new_n713_), .A2(new_n6284_), .B1(new_n5761_), .B2(new_n717_), .ZN(new_n8196_));
  AOI21_X1   g07940(.A1(\b[38] ), .A2(new_n1126_), .B(new_n8196_), .ZN(new_n8197_));
  OAI21_X1   g07941(.A1(new_n8195_), .A2(new_n986_), .B(new_n8197_), .ZN(new_n8198_));
  XOR2_X1    g07942(.A1(new_n8198_), .A2(\a[11] ), .Z(new_n8199_));
  OAI22_X1   g07943(.A1(new_n993_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n997_), .ZN(new_n8200_));
  AOI21_X1   g07944(.A1(\b[35] ), .A2(new_n1486_), .B(new_n8200_), .ZN(new_n8201_));
  OAI21_X1   g07945(.A1(new_n5322_), .A2(new_n1323_), .B(new_n8201_), .ZN(new_n8202_));
  XOR2_X1    g07946(.A1(new_n8202_), .A2(\a[14] ), .Z(new_n8203_));
  OAI22_X1   g07947(.A1(new_n1592_), .A2(new_n4639_), .B1(new_n4638_), .B2(new_n1505_), .ZN(new_n8204_));
  AOI21_X1   g07948(.A1(\b[32] ), .A2(new_n1584_), .B(new_n8204_), .ZN(new_n8205_));
  OAI21_X1   g07949(.A1(new_n4649_), .A2(new_n1732_), .B(new_n8205_), .ZN(new_n8206_));
  XOR2_X1    g07950(.A1(new_n8206_), .A2(\a[17] ), .Z(new_n8207_));
  NOR2_X1    g07951(.A1(new_n8046_), .A2(new_n8040_), .ZN(new_n8208_));
  AOI22_X1   g07952(.A1(new_n2202_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n2205_), .ZN(new_n8209_));
  OAI21_X1   g07953(.A1(new_n3006_), .A2(new_n2370_), .B(new_n8209_), .ZN(new_n8210_));
  AOI21_X1   g07954(.A1(new_n3807_), .A2(new_n2208_), .B(new_n8210_), .ZN(new_n8211_));
  XOR2_X1    g07955(.A1(new_n8211_), .A2(new_n2200_), .Z(new_n8212_));
  INV_X1     g07956(.I(new_n8212_), .ZN(new_n8213_));
  OAI22_X1   g07957(.A1(new_n2703_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n2708_), .ZN(new_n8214_));
  AOI21_X1   g07958(.A1(\b[23] ), .A2(new_n2906_), .B(new_n8214_), .ZN(new_n8215_));
  OAI21_X1   g07959(.A1(new_n2655_), .A2(new_n2711_), .B(new_n8215_), .ZN(new_n8216_));
  XOR2_X1    g07960(.A1(new_n8216_), .A2(\a[26] ), .Z(new_n8217_));
  INV_X1     g07961(.I(new_n8217_), .ZN(new_n8218_));
  AOI22_X1   g07962(.A1(new_n3267_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n3270_), .ZN(new_n8219_));
  OAI21_X1   g07963(.A1(new_n1860_), .A2(new_n3475_), .B(new_n8219_), .ZN(new_n8220_));
  AOI21_X1   g07964(.A1(new_n2659_), .A2(new_n3273_), .B(new_n8220_), .ZN(new_n8221_));
  XOR2_X1    g07965(.A1(new_n8221_), .A2(new_n3264_), .Z(new_n8222_));
  INV_X1     g07966(.I(new_n8222_), .ZN(new_n8223_));
  AOI22_X1   g07967(.A1(new_n3864_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n3869_), .ZN(new_n8224_));
  OAI21_X1   g07968(.A1(new_n1432_), .A2(new_n5410_), .B(new_n8224_), .ZN(new_n8225_));
  AOI21_X1   g07969(.A1(new_n1695_), .A2(new_n3872_), .B(new_n8225_), .ZN(new_n8226_));
  XOR2_X1    g07970(.A1(new_n8226_), .A2(new_n3876_), .Z(new_n8227_));
  INV_X1     g07971(.I(new_n8227_), .ZN(new_n8228_));
  AOI21_X1   g07972(.A1(new_n7975_), .A2(new_n7970_), .B(new_n7966_), .ZN(new_n8229_));
  AOI21_X1   g07973(.A1(new_n7956_), .A2(new_n7955_), .B(new_n7962_), .ZN(new_n8230_));
  NOR2_X1    g07974(.A1(new_n7949_), .A2(new_n7947_), .ZN(new_n8231_));
  AOI21_X1   g07975(.A1(new_n7949_), .A2(new_n7947_), .B(new_n7943_), .ZN(new_n8232_));
  NOR2_X1    g07976(.A1(new_n8232_), .A2(new_n8231_), .ZN(new_n8233_));
  INV_X1     g07977(.I(new_n8233_), .ZN(new_n8234_));
  AOI22_X1   g07978(.A1(new_n7403_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n7408_), .ZN(new_n8235_));
  NAND2_X1   g07979(.A1(new_n7719_), .A2(\b[2] ), .ZN(new_n8236_));
  NAND2_X1   g07980(.A1(new_n1725_), .A2(new_n7414_), .ZN(new_n8237_));
  NAND3_X1   g07981(.A1(new_n8237_), .A2(new_n8235_), .A3(new_n8236_), .ZN(new_n8238_));
  XOR2_X1    g07982(.A1(new_n8238_), .A2(new_n7410_), .Z(new_n8239_));
  XOR2_X1    g07983(.A1(\a[49] ), .A2(\a[50] ), .Z(new_n8240_));
  NOR2_X1    g07984(.A1(new_n7936_), .A2(new_n8240_), .ZN(new_n8241_));
  INV_X1     g07985(.I(\a[48] ), .ZN(new_n8242_));
  NAND3_X1   g07986(.A1(new_n7410_), .A2(new_n8242_), .A3(\a[49] ), .ZN(new_n8243_));
  INV_X1     g07987(.I(\a[49] ), .ZN(new_n8244_));
  NAND3_X1   g07988(.A1(new_n8244_), .A2(\a[47] ), .A3(\a[48] ), .ZN(new_n8245_));
  NAND2_X1   g07989(.A1(new_n8243_), .A2(new_n8245_), .ZN(new_n8246_));
  AOI22_X1   g07990(.A1(new_n8241_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n8246_), .ZN(new_n8247_));
  INV_X1     g07991(.I(\a[50] ), .ZN(new_n8248_));
  NOR2_X1    g07992(.A1(new_n8248_), .A2(\a[49] ), .ZN(new_n8249_));
  NOR2_X1    g07993(.A1(new_n8244_), .A2(\a[50] ), .ZN(new_n8250_));
  NOR2_X1    g07994(.A1(new_n8249_), .A2(new_n8250_), .ZN(new_n8251_));
  NOR2_X1    g07995(.A1(new_n8251_), .A2(new_n7936_), .ZN(new_n8252_));
  NAND2_X1   g07996(.A1(new_n8252_), .A2(new_n263_), .ZN(new_n8253_));
  NAND2_X1   g07997(.A1(new_n8247_), .A2(new_n8253_), .ZN(new_n8254_));
  NAND2_X1   g07998(.A1(new_n8254_), .A2(\a[50] ), .ZN(new_n8255_));
  INV_X1     g07999(.I(new_n8254_), .ZN(new_n8256_));
  NAND2_X1   g08000(.A1(new_n8256_), .A2(new_n8248_), .ZN(new_n8257_));
  NOR2_X1    g08001(.A1(new_n7937_), .A2(new_n8248_), .ZN(new_n8258_));
  INV_X1     g08002(.I(new_n8258_), .ZN(new_n8259_));
  NAND3_X1   g08003(.A1(new_n8257_), .A2(new_n8255_), .A3(new_n8259_), .ZN(new_n8260_));
  NOR2_X1    g08004(.A1(new_n8255_), .A2(new_n7937_), .ZN(new_n8261_));
  INV_X1     g08005(.I(new_n8261_), .ZN(new_n8262_));
  AOI21_X1   g08006(.A1(new_n8260_), .A2(new_n8262_), .B(new_n8239_), .ZN(new_n8263_));
  NAND3_X1   g08007(.A1(new_n8239_), .A2(new_n8260_), .A3(new_n8262_), .ZN(new_n8264_));
  INV_X1     g08008(.I(new_n8264_), .ZN(new_n8265_));
  NOR2_X1    g08009(.A1(new_n8265_), .A2(new_n8263_), .ZN(new_n8266_));
  NOR2_X1    g08010(.A1(new_n7940_), .A2(new_n7937_), .ZN(new_n8267_));
  AOI21_X1   g08011(.A1(new_n7726_), .A2(new_n7941_), .B(new_n8267_), .ZN(new_n8268_));
  INV_X1     g08012(.I(new_n8268_), .ZN(new_n8269_));
  NOR2_X1    g08013(.A1(new_n8269_), .A2(new_n8266_), .ZN(new_n8270_));
  NOR3_X1    g08014(.A1(new_n8268_), .A2(new_n8263_), .A3(new_n8265_), .ZN(new_n8271_));
  NOR2_X1    g08015(.A1(new_n8270_), .A2(new_n8271_), .ZN(new_n8272_));
  OAI22_X1   g08016(.A1(new_n7730_), .A2(new_n471_), .B1(new_n438_), .B2(new_n7731_), .ZN(new_n8273_));
  AOI21_X1   g08017(.A1(\b[5] ), .A2(new_n6887_), .B(new_n8273_), .ZN(new_n8274_));
  OAI21_X1   g08018(.A1(new_n485_), .A2(new_n7728_), .B(new_n8274_), .ZN(new_n8275_));
  XOR2_X1    g08019(.A1(new_n8275_), .A2(\a[44] ), .Z(new_n8276_));
  INV_X1     g08020(.I(new_n8276_), .ZN(new_n8277_));
  XOR2_X1    g08021(.A1(new_n8272_), .A2(new_n8277_), .Z(new_n8278_));
  NAND2_X1   g08022(.A1(new_n8234_), .A2(new_n8278_), .ZN(new_n8279_));
  XOR2_X1    g08023(.A1(new_n8272_), .A2(new_n8276_), .Z(new_n8280_));
  NAND2_X1   g08024(.A1(new_n8280_), .A2(new_n8233_), .ZN(new_n8281_));
  AOI22_X1   g08025(.A1(new_n6108_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n6111_), .ZN(new_n8282_));
  OAI21_X1   g08026(.A1(new_n577_), .A2(new_n7708_), .B(new_n8282_), .ZN(new_n8283_));
  AOI21_X1   g08027(.A1(new_n1059_), .A2(new_n6105_), .B(new_n8283_), .ZN(new_n8284_));
  XOR2_X1    g08028(.A1(new_n8284_), .A2(new_n5849_), .Z(new_n8285_));
  INV_X1     g08029(.I(new_n8285_), .ZN(new_n8286_));
  NAND3_X1   g08030(.A1(new_n8279_), .A2(new_n8281_), .A3(new_n8286_), .ZN(new_n8287_));
  NOR2_X1    g08031(.A1(new_n8280_), .A2(new_n8233_), .ZN(new_n8288_));
  NOR2_X1    g08032(.A1(new_n8234_), .A2(new_n8278_), .ZN(new_n8289_));
  OAI21_X1   g08033(.A1(new_n8289_), .A2(new_n8288_), .B(new_n8285_), .ZN(new_n8290_));
  NAND2_X1   g08034(.A1(new_n8290_), .A2(new_n8287_), .ZN(new_n8291_));
  OAI21_X1   g08035(.A1(new_n8230_), .A2(new_n7964_), .B(new_n8291_), .ZN(new_n8292_));
  OAI21_X1   g08036(.A1(new_n7959_), .A2(new_n7958_), .B(new_n7951_), .ZN(new_n8293_));
  NOR3_X1    g08037(.A1(new_n8289_), .A2(new_n8288_), .A3(new_n8285_), .ZN(new_n8294_));
  AOI21_X1   g08038(.A1(new_n8279_), .A2(new_n8281_), .B(new_n8286_), .ZN(new_n8295_));
  NOR2_X1    g08039(.A1(new_n8294_), .A2(new_n8295_), .ZN(new_n8296_));
  NAND3_X1   g08040(.A1(new_n8293_), .A2(new_n8296_), .A3(new_n7960_), .ZN(new_n8297_));
  OAI22_X1   g08041(.A1(new_n1070_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n941_), .ZN(new_n8298_));
  AOI21_X1   g08042(.A1(\b[11] ), .A2(new_n5420_), .B(new_n8298_), .ZN(new_n8299_));
  OAI21_X1   g08043(.A1(new_n1082_), .A2(new_n6124_), .B(new_n8299_), .ZN(new_n8300_));
  XOR2_X1    g08044(.A1(new_n8300_), .A2(\a[38] ), .Z(new_n8301_));
  AOI21_X1   g08045(.A1(new_n8292_), .A2(new_n8297_), .B(new_n8301_), .ZN(new_n8302_));
  AOI21_X1   g08046(.A1(new_n8293_), .A2(new_n7960_), .B(new_n8296_), .ZN(new_n8303_));
  NOR3_X1    g08047(.A1(new_n8230_), .A2(new_n7964_), .A3(new_n8291_), .ZN(new_n8304_));
  INV_X1     g08048(.I(new_n8301_), .ZN(new_n8305_));
  NOR3_X1    g08049(.A1(new_n8303_), .A2(new_n8304_), .A3(new_n8305_), .ZN(new_n8306_));
  NOR2_X1    g08050(.A1(new_n8306_), .A2(new_n8302_), .ZN(new_n8307_));
  OAI21_X1   g08051(.A1(new_n8229_), .A2(new_n7976_), .B(new_n8307_), .ZN(new_n8308_));
  OAI21_X1   g08052(.A1(new_n7972_), .A2(new_n7971_), .B(new_n7980_), .ZN(new_n8309_));
  OAI21_X1   g08053(.A1(new_n8303_), .A2(new_n8304_), .B(new_n8305_), .ZN(new_n8310_));
  NAND3_X1   g08054(.A1(new_n8292_), .A2(new_n8297_), .A3(new_n8301_), .ZN(new_n8311_));
  NAND2_X1   g08055(.A1(new_n8310_), .A2(new_n8311_), .ZN(new_n8312_));
  NAND3_X1   g08056(.A1(new_n8309_), .A2(new_n8312_), .A3(new_n7982_), .ZN(new_n8313_));
  AOI22_X1   g08057(.A1(new_n4918_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n4921_), .ZN(new_n8314_));
  OAI21_X1   g08058(.A1(new_n1093_), .A2(new_n6099_), .B(new_n8314_), .ZN(new_n8315_));
  AOI21_X1   g08059(.A1(new_n1701_), .A2(new_n4699_), .B(new_n8315_), .ZN(new_n8316_));
  XOR2_X1    g08060(.A1(new_n8316_), .A2(new_n4446_), .Z(new_n8317_));
  INV_X1     g08061(.I(new_n8317_), .ZN(new_n8318_));
  NAND3_X1   g08062(.A1(new_n8308_), .A2(new_n8313_), .A3(new_n8318_), .ZN(new_n8319_));
  AOI21_X1   g08063(.A1(new_n8309_), .A2(new_n7982_), .B(new_n8312_), .ZN(new_n8320_));
  NOR3_X1    g08064(.A1(new_n8307_), .A2(new_n8229_), .A3(new_n7976_), .ZN(new_n8321_));
  OAI21_X1   g08065(.A1(new_n8320_), .A2(new_n8321_), .B(new_n8317_), .ZN(new_n8322_));
  NAND2_X1   g08066(.A1(new_n8322_), .A2(new_n8319_), .ZN(new_n8323_));
  NOR2_X1    g08067(.A1(new_n7483_), .A2(new_n7482_), .ZN(new_n8324_));
  AOI21_X1   g08068(.A1(new_n8324_), .A2(new_n7475_), .B(new_n7469_), .ZN(new_n8325_));
  OAI21_X1   g08069(.A1(new_n8325_), .A2(new_n7785_), .B(new_n7783_), .ZN(new_n8326_));
  AOI21_X1   g08070(.A1(new_n8326_), .A2(new_n7988_), .B(new_n7994_), .ZN(new_n8327_));
  NOR3_X1    g08071(.A1(new_n8327_), .A2(new_n7996_), .A3(new_n8323_), .ZN(new_n8328_));
  NOR3_X1    g08072(.A1(new_n8320_), .A2(new_n8321_), .A3(new_n8317_), .ZN(new_n8329_));
  AOI21_X1   g08073(.A1(new_n8308_), .A2(new_n8313_), .B(new_n8318_), .ZN(new_n8330_));
  NOR2_X1    g08074(.A1(new_n8329_), .A2(new_n8330_), .ZN(new_n8331_));
  OAI21_X1   g08075(.A1(new_n7991_), .A2(new_n7990_), .B(new_n7984_), .ZN(new_n8332_));
  AOI21_X1   g08076(.A1(new_n8332_), .A2(new_n7992_), .B(new_n8331_), .ZN(new_n8333_));
  OAI21_X1   g08077(.A1(new_n8328_), .A2(new_n8333_), .B(new_n8228_), .ZN(new_n8334_));
  NAND3_X1   g08078(.A1(new_n8332_), .A2(new_n8331_), .A3(new_n7992_), .ZN(new_n8335_));
  OAI21_X1   g08079(.A1(new_n8327_), .A2(new_n7996_), .B(new_n8323_), .ZN(new_n8336_));
  NAND3_X1   g08080(.A1(new_n8336_), .A2(new_n8335_), .A3(new_n8227_), .ZN(new_n8337_));
  NAND2_X1   g08081(.A1(new_n8334_), .A2(new_n8337_), .ZN(new_n8338_));
  AOI21_X1   g08082(.A1(new_n8004_), .A2(new_n8003_), .B(new_n7998_), .ZN(new_n8339_));
  NOR3_X1    g08083(.A1(new_n8338_), .A2(new_n8339_), .A3(new_n8012_), .ZN(new_n8340_));
  AOI21_X1   g08084(.A1(new_n8336_), .A2(new_n8335_), .B(new_n8227_), .ZN(new_n8341_));
  NOR3_X1    g08085(.A1(new_n8328_), .A2(new_n8333_), .A3(new_n8228_), .ZN(new_n8342_));
  NOR2_X1    g08086(.A1(new_n8342_), .A2(new_n8341_), .ZN(new_n8343_));
  OAI21_X1   g08087(.A1(new_n8008_), .A2(new_n8006_), .B(new_n7999_), .ZN(new_n8344_));
  AOI21_X1   g08088(.A1(new_n8344_), .A2(new_n8009_), .B(new_n8343_), .ZN(new_n8345_));
  OAI21_X1   g08089(.A1(new_n8345_), .A2(new_n8340_), .B(new_n8223_), .ZN(new_n8346_));
  NAND3_X1   g08090(.A1(new_n8344_), .A2(new_n8343_), .A3(new_n8009_), .ZN(new_n8347_));
  OAI21_X1   g08091(.A1(new_n8339_), .A2(new_n8012_), .B(new_n8338_), .ZN(new_n8348_));
  NAND3_X1   g08092(.A1(new_n8347_), .A2(new_n8348_), .A3(new_n8222_), .ZN(new_n8349_));
  NAND2_X1   g08093(.A1(new_n8349_), .A2(new_n8346_), .ZN(new_n8350_));
  NOR2_X1    g08094(.A1(new_n7500_), .A2(new_n7502_), .ZN(new_n8351_));
  OAI21_X1   g08095(.A1(new_n8351_), .A2(new_n7814_), .B(new_n7813_), .ZN(new_n8352_));
  AOI21_X1   g08096(.A1(new_n8352_), .A2(new_n8018_), .B(new_n8023_), .ZN(new_n8353_));
  NOR3_X1    g08097(.A1(new_n8353_), .A2(new_n8020_), .A3(new_n8350_), .ZN(new_n8354_));
  AOI21_X1   g08098(.A1(new_n8347_), .A2(new_n8348_), .B(new_n8222_), .ZN(new_n8355_));
  NOR3_X1    g08099(.A1(new_n8345_), .A2(new_n8340_), .A3(new_n8223_), .ZN(new_n8356_));
  NOR2_X1    g08100(.A1(new_n8355_), .A2(new_n8356_), .ZN(new_n8357_));
  NAND2_X1   g08101(.A1(new_n8019_), .A2(new_n8014_), .ZN(new_n8358_));
  AOI21_X1   g08102(.A1(new_n8358_), .A2(new_n8021_), .B(new_n8357_), .ZN(new_n8359_));
  OAI21_X1   g08103(.A1(new_n8359_), .A2(new_n8354_), .B(new_n8218_), .ZN(new_n8360_));
  NAND3_X1   g08104(.A1(new_n8358_), .A2(new_n8021_), .A3(new_n8357_), .ZN(new_n8361_));
  OAI21_X1   g08105(.A1(new_n8353_), .A2(new_n8020_), .B(new_n8350_), .ZN(new_n8362_));
  NAND3_X1   g08106(.A1(new_n8361_), .A2(new_n8362_), .A3(new_n8217_), .ZN(new_n8363_));
  NAND2_X1   g08107(.A1(new_n8360_), .A2(new_n8363_), .ZN(new_n8364_));
  AOI21_X1   g08108(.A1(new_n7184_), .A2(new_n7189_), .B(new_n7199_), .ZN(new_n8365_));
  AOI21_X1   g08109(.A1(new_n8365_), .A2(new_n7511_), .B(new_n7691_), .ZN(new_n8366_));
  OAI21_X1   g08110(.A1(new_n8366_), .A2(new_n7821_), .B(new_n7816_), .ZN(new_n8367_));
  AOI21_X1   g08111(.A1(new_n8367_), .A2(new_n8030_), .B(new_n8026_), .ZN(new_n8368_));
  NOR3_X1    g08112(.A1(new_n8368_), .A2(new_n8364_), .A3(new_n8033_), .ZN(new_n8369_));
  AOI21_X1   g08113(.A1(new_n8361_), .A2(new_n8362_), .B(new_n8217_), .ZN(new_n8370_));
  NOR3_X1    g08114(.A1(new_n8359_), .A2(new_n8354_), .A3(new_n8218_), .ZN(new_n8371_));
  NOR2_X1    g08115(.A1(new_n8370_), .A2(new_n8371_), .ZN(new_n8372_));
  AOI21_X1   g08116(.A1(new_n8035_), .A2(new_n8036_), .B(new_n8033_), .ZN(new_n8373_));
  NOR2_X1    g08117(.A1(new_n8373_), .A2(new_n8372_), .ZN(new_n8374_));
  OAI21_X1   g08118(.A1(new_n8374_), .A2(new_n8369_), .B(new_n8213_), .ZN(new_n8375_));
  NAND2_X1   g08119(.A1(new_n8035_), .A2(new_n8036_), .ZN(new_n8376_));
  NAND3_X1   g08120(.A1(new_n8376_), .A2(new_n8037_), .A3(new_n8372_), .ZN(new_n8377_));
  OAI21_X1   g08121(.A1(new_n8368_), .A2(new_n8033_), .B(new_n8364_), .ZN(new_n8378_));
  NAND3_X1   g08122(.A1(new_n8377_), .A2(new_n8378_), .A3(new_n8212_), .ZN(new_n8379_));
  NAND2_X1   g08123(.A1(new_n8375_), .A2(new_n8379_), .ZN(new_n8380_));
  OAI21_X1   g08124(.A1(new_n8208_), .A2(new_n8047_), .B(new_n8380_), .ZN(new_n8381_));
  NAND2_X1   g08125(.A1(new_n8049_), .A2(new_n8039_), .ZN(new_n8382_));
  AOI21_X1   g08126(.A1(new_n8377_), .A2(new_n8378_), .B(new_n8212_), .ZN(new_n8383_));
  NOR3_X1    g08127(.A1(new_n8374_), .A2(new_n8369_), .A3(new_n8213_), .ZN(new_n8384_));
  NOR2_X1    g08128(.A1(new_n8384_), .A2(new_n8383_), .ZN(new_n8385_));
  NAND3_X1   g08129(.A1(new_n8382_), .A2(new_n8385_), .A3(new_n8050_), .ZN(new_n8386_));
  AOI22_X1   g08130(.A1(new_n1738_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n1743_), .ZN(new_n8387_));
  OAI21_X1   g08131(.A1(new_n3592_), .A2(new_n1931_), .B(new_n8387_), .ZN(new_n8388_));
  AOI21_X1   g08132(.A1(new_n3796_), .A2(new_n1746_), .B(new_n8388_), .ZN(new_n8389_));
  XOR2_X1    g08133(.A1(new_n8389_), .A2(new_n1736_), .Z(new_n8390_));
  AOI21_X1   g08134(.A1(new_n8381_), .A2(new_n8386_), .B(new_n8390_), .ZN(new_n8391_));
  AOI21_X1   g08135(.A1(new_n8039_), .A2(new_n8049_), .B(new_n8047_), .ZN(new_n8392_));
  NOR2_X1    g08136(.A1(new_n8392_), .A2(new_n8385_), .ZN(new_n8393_));
  NOR3_X1    g08137(.A1(new_n8208_), .A2(new_n8047_), .A3(new_n8380_), .ZN(new_n8394_));
  INV_X1     g08138(.I(new_n8390_), .ZN(new_n8395_));
  NOR3_X1    g08139(.A1(new_n8393_), .A2(new_n8395_), .A3(new_n8394_), .ZN(new_n8396_));
  NOR2_X1    g08140(.A1(new_n8396_), .A2(new_n8391_), .ZN(new_n8397_));
  NAND2_X1   g08141(.A1(new_n8062_), .A2(new_n8052_), .ZN(new_n8398_));
  NAND3_X1   g08142(.A1(new_n8398_), .A2(new_n8397_), .A3(new_n8063_), .ZN(new_n8399_));
  OAI21_X1   g08143(.A1(new_n8393_), .A2(new_n8394_), .B(new_n8395_), .ZN(new_n8400_));
  NAND3_X1   g08144(.A1(new_n8381_), .A2(new_n8386_), .A3(new_n8390_), .ZN(new_n8401_));
  NAND2_X1   g08145(.A1(new_n8400_), .A2(new_n8401_), .ZN(new_n8402_));
  AOI21_X1   g08146(.A1(new_n7220_), .A2(new_n7225_), .B(new_n7540_), .ZN(new_n8403_));
  AOI21_X1   g08147(.A1(new_n8403_), .A2(new_n7538_), .B(new_n7680_), .ZN(new_n8404_));
  OAI21_X1   g08148(.A1(new_n8404_), .A2(new_n7842_), .B(new_n7837_), .ZN(new_n8405_));
  AOI21_X1   g08149(.A1(new_n8405_), .A2(new_n8057_), .B(new_n8053_), .ZN(new_n8406_));
  OAI21_X1   g08150(.A1(new_n8406_), .A2(new_n8060_), .B(new_n8402_), .ZN(new_n8407_));
  AOI21_X1   g08151(.A1(new_n8407_), .A2(new_n8399_), .B(new_n8207_), .ZN(new_n8408_));
  INV_X1     g08152(.I(new_n8207_), .ZN(new_n8409_));
  NOR3_X1    g08153(.A1(new_n8406_), .A2(new_n8402_), .A3(new_n8060_), .ZN(new_n8410_));
  AOI21_X1   g08154(.A1(new_n8052_), .A2(new_n8062_), .B(new_n8060_), .ZN(new_n8411_));
  NOR2_X1    g08155(.A1(new_n8411_), .A2(new_n8397_), .ZN(new_n8412_));
  NOR3_X1    g08156(.A1(new_n8412_), .A2(new_n8410_), .A3(new_n8409_), .ZN(new_n8413_));
  NOR2_X1    g08157(.A1(new_n8413_), .A2(new_n8408_), .ZN(new_n8414_));
  NAND2_X1   g08158(.A1(new_n8076_), .A2(new_n8065_), .ZN(new_n8415_));
  NAND3_X1   g08159(.A1(new_n8415_), .A2(new_n8077_), .A3(new_n8414_), .ZN(new_n8416_));
  OAI21_X1   g08160(.A1(new_n8412_), .A2(new_n8410_), .B(new_n8409_), .ZN(new_n8417_));
  NAND3_X1   g08161(.A1(new_n8407_), .A2(new_n8399_), .A3(new_n8207_), .ZN(new_n8418_));
  NAND2_X1   g08162(.A1(new_n8417_), .A2(new_n8418_), .ZN(new_n8419_));
  NOR2_X1    g08163(.A1(new_n8071_), .A2(new_n8075_), .ZN(new_n8420_));
  OAI21_X1   g08164(.A1(new_n8420_), .A2(new_n8072_), .B(new_n8419_), .ZN(new_n8421_));
  AOI21_X1   g08165(.A1(new_n8416_), .A2(new_n8421_), .B(new_n8203_), .ZN(new_n8422_));
  XOR2_X1    g08166(.A1(new_n8202_), .A2(new_n1002_), .Z(new_n8423_));
  NOR3_X1    g08167(.A1(new_n8420_), .A2(new_n8072_), .A3(new_n8419_), .ZN(new_n8424_));
  AOI21_X1   g08168(.A1(new_n8415_), .A2(new_n8077_), .B(new_n8414_), .ZN(new_n8425_));
  NOR3_X1    g08169(.A1(new_n8425_), .A2(new_n8424_), .A3(new_n8423_), .ZN(new_n8426_));
  NOR2_X1    g08170(.A1(new_n8422_), .A2(new_n8426_), .ZN(new_n8427_));
  OAI21_X1   g08171(.A1(new_n7242_), .A2(new_n7248_), .B(new_n7254_), .ZN(new_n8428_));
  OAI21_X1   g08172(.A1(new_n8428_), .A2(new_n7578_), .B(new_n7870_), .ZN(new_n8429_));
  AOI21_X1   g08173(.A1(new_n8429_), .A2(new_n7864_), .B(new_n7863_), .ZN(new_n8430_));
  OAI21_X1   g08174(.A1(new_n8430_), .A2(new_n8085_), .B(new_n8091_), .ZN(new_n8431_));
  NAND3_X1   g08175(.A1(new_n8431_), .A2(new_n8093_), .A3(new_n8427_), .ZN(new_n8432_));
  OAI21_X1   g08176(.A1(new_n8425_), .A2(new_n8424_), .B(new_n8423_), .ZN(new_n8433_));
  NAND3_X1   g08177(.A1(new_n8416_), .A2(new_n8421_), .A3(new_n8203_), .ZN(new_n8434_));
  NAND2_X1   g08178(.A1(new_n8433_), .A2(new_n8434_), .ZN(new_n8435_));
  AOI21_X1   g08179(.A1(new_n7252_), .A2(new_n7253_), .B(new_n7249_), .ZN(new_n8436_));
  AOI21_X1   g08180(.A1(new_n8436_), .A2(new_n7570_), .B(new_n7865_), .ZN(new_n8437_));
  OAI21_X1   g08181(.A1(new_n8437_), .A2(new_n7869_), .B(new_n7868_), .ZN(new_n8438_));
  AOI21_X1   g08182(.A1(new_n8438_), .A2(new_n8084_), .B(new_n8080_), .ZN(new_n8439_));
  OAI21_X1   g08183(.A1(new_n8439_), .A2(new_n8087_), .B(new_n8435_), .ZN(new_n8440_));
  AOI21_X1   g08184(.A1(new_n8432_), .A2(new_n8440_), .B(new_n8199_), .ZN(new_n8441_));
  XOR2_X1    g08185(.A1(new_n8198_), .A2(new_n722_), .Z(new_n8442_));
  NOR3_X1    g08186(.A1(new_n8439_), .A2(new_n8435_), .A3(new_n8087_), .ZN(new_n8443_));
  AOI21_X1   g08187(.A1(new_n8431_), .A2(new_n8093_), .B(new_n8427_), .ZN(new_n8444_));
  NOR3_X1    g08188(.A1(new_n8444_), .A2(new_n8443_), .A3(new_n8442_), .ZN(new_n8445_));
  NOR2_X1    g08189(.A1(new_n8441_), .A2(new_n8445_), .ZN(new_n8446_));
  OAI21_X1   g08190(.A1(new_n7257_), .A2(new_n7264_), .B(new_n7269_), .ZN(new_n8447_));
  OAI21_X1   g08191(.A1(new_n8447_), .A2(new_n7585_), .B(new_n7580_), .ZN(new_n8448_));
  AOI21_X1   g08192(.A1(new_n8448_), .A2(new_n7877_), .B(new_n7876_), .ZN(new_n8449_));
  OAI21_X1   g08193(.A1(new_n8449_), .A2(new_n8101_), .B(new_n8095_), .ZN(new_n8450_));
  NAND3_X1   g08194(.A1(new_n8450_), .A2(new_n8102_), .A3(new_n8446_), .ZN(new_n8451_));
  OAI21_X1   g08195(.A1(new_n8444_), .A2(new_n8443_), .B(new_n8442_), .ZN(new_n8452_));
  NAND3_X1   g08196(.A1(new_n8432_), .A2(new_n8440_), .A3(new_n8199_), .ZN(new_n8453_));
  NAND2_X1   g08197(.A1(new_n8452_), .A2(new_n8453_), .ZN(new_n8454_));
  AOI21_X1   g08198(.A1(new_n7256_), .A2(new_n7268_), .B(new_n7266_), .ZN(new_n8455_));
  AOI21_X1   g08199(.A1(new_n8455_), .A2(new_n7592_), .B(new_n7590_), .ZN(new_n8456_));
  OAI21_X1   g08200(.A1(new_n8456_), .A2(new_n7881_), .B(new_n7880_), .ZN(new_n8457_));
  AOI21_X1   g08201(.A1(new_n8457_), .A2(new_n8099_), .B(new_n8104_), .ZN(new_n8458_));
  OAI21_X1   g08202(.A1(new_n8458_), .A2(new_n8106_), .B(new_n8454_), .ZN(new_n8459_));
  AOI21_X1   g08203(.A1(new_n8459_), .A2(new_n8451_), .B(new_n8194_), .ZN(new_n8460_));
  XOR2_X1    g08204(.A1(new_n8193_), .A2(new_n488_), .Z(new_n8461_));
  NOR3_X1    g08205(.A1(new_n8458_), .A2(new_n8106_), .A3(new_n8454_), .ZN(new_n8462_));
  AOI21_X1   g08206(.A1(new_n8450_), .A2(new_n8102_), .B(new_n8446_), .ZN(new_n8463_));
  NOR3_X1    g08207(.A1(new_n8462_), .A2(new_n8463_), .A3(new_n8461_), .ZN(new_n8464_));
  NOR2_X1    g08208(.A1(new_n8464_), .A2(new_n8460_), .ZN(new_n8465_));
  NAND2_X1   g08209(.A1(new_n8116_), .A2(new_n8109_), .ZN(new_n8466_));
  NAND3_X1   g08210(.A1(new_n8466_), .A2(new_n8118_), .A3(new_n8465_), .ZN(new_n8467_));
  NOR3_X1    g08211(.A1(new_n8111_), .A2(new_n7893_), .A3(new_n8115_), .ZN(new_n8468_));
  OAI21_X1   g08212(.A1(new_n8462_), .A2(new_n8463_), .B(new_n8461_), .ZN(new_n8469_));
  NAND3_X1   g08213(.A1(new_n8459_), .A2(new_n8451_), .A3(new_n8194_), .ZN(new_n8470_));
  NAND2_X1   g08214(.A1(new_n8469_), .A2(new_n8470_), .ZN(new_n8471_));
  OAI21_X1   g08215(.A1(new_n7654_), .A2(new_n7890_), .B(new_n7883_), .ZN(new_n8472_));
  AOI21_X1   g08216(.A1(new_n8472_), .A2(new_n8115_), .B(new_n8108_), .ZN(new_n8473_));
  OAI21_X1   g08217(.A1(new_n8473_), .A2(new_n8468_), .B(new_n8471_), .ZN(new_n8474_));
  NAND3_X1   g08218(.A1(new_n8467_), .A2(new_n8474_), .A3(new_n8188_), .ZN(new_n8475_));
  INV_X1     g08219(.I(new_n8188_), .ZN(new_n8476_));
  NOR3_X1    g08220(.A1(new_n8473_), .A2(new_n8471_), .A3(new_n8468_), .ZN(new_n8477_));
  AOI21_X1   g08221(.A1(new_n8466_), .A2(new_n8118_), .B(new_n8465_), .ZN(new_n8478_));
  OAI21_X1   g08222(.A1(new_n8478_), .A2(new_n8477_), .B(new_n8476_), .ZN(new_n8479_));
  NAND2_X1   g08223(.A1(new_n8479_), .A2(new_n8475_), .ZN(new_n8480_));
  OAI21_X1   g08224(.A1(new_n8182_), .A2(new_n8183_), .B(new_n8480_), .ZN(new_n8481_));
  INV_X1     g08225(.I(new_n8183_), .ZN(new_n8482_));
  NOR3_X1    g08226(.A1(new_n8478_), .A2(new_n8477_), .A3(new_n8476_), .ZN(new_n8483_));
  AOI21_X1   g08227(.A1(new_n8467_), .A2(new_n8474_), .B(new_n8188_), .ZN(new_n8484_));
  NOR2_X1    g08228(.A1(new_n8483_), .A2(new_n8484_), .ZN(new_n8485_));
  NAND3_X1   g08229(.A1(new_n8482_), .A2(new_n8181_), .A3(new_n8485_), .ZN(new_n8486_));
  NAND2_X1   g08230(.A1(new_n8481_), .A2(new_n8486_), .ZN(new_n8487_));
  XOR2_X1    g08231(.A1(new_n8162_), .A2(new_n8487_), .Z(\f[49] ));
  NOR3_X1    g08232(.A1(new_n7632_), .A2(new_n7616_), .A3(new_n7629_), .ZN(new_n8489_));
  AOI21_X1   g08233(.A1(new_n7615_), .A2(new_n7633_), .B(new_n8489_), .ZN(new_n8490_));
  INV_X1     g08234(.I(new_n7921_), .ZN(new_n8491_));
  AOI21_X1   g08235(.A1(new_n8490_), .A2(new_n8491_), .B(new_n8155_), .ZN(new_n8492_));
  INV_X1     g08236(.I(new_n8161_), .ZN(new_n8493_));
  OAI21_X1   g08237(.A1(new_n8492_), .A2(new_n8153_), .B(new_n8493_), .ZN(new_n8494_));
  INV_X1     g08238(.I(new_n8487_), .ZN(new_n8495_));
  INV_X1     g08239(.I(new_n8177_), .ZN(new_n8496_));
  XOR2_X1    g08240(.A1(new_n8180_), .A2(new_n8480_), .Z(new_n8497_));
  NOR2_X1    g08241(.A1(new_n8497_), .A2(new_n8496_), .ZN(new_n8498_));
  AOI21_X1   g08242(.A1(new_n8494_), .A2(new_n8495_), .B(new_n8498_), .ZN(new_n8499_));
  INV_X1     g08243(.I(\b[50] ), .ZN(new_n8500_));
  OAI22_X1   g08244(.A1(new_n277_), .A2(new_n8500_), .B1(new_n8168_), .B2(new_n262_), .ZN(new_n8501_));
  AOI21_X1   g08245(.A1(\b[48] ), .A2(new_n283_), .B(new_n8501_), .ZN(new_n8502_));
  AOI21_X1   g08246(.A1(new_n8169_), .A2(\b[48] ), .B(\b[47] ), .ZN(new_n8503_));
  AOI21_X1   g08247(.A1(new_n8136_), .A2(\b[49] ), .B(\b[48] ), .ZN(new_n8504_));
  NOR2_X1    g08248(.A1(new_n8503_), .A2(new_n8504_), .ZN(new_n8505_));
  XNOR2_X1   g08249(.A1(\b[49] ), .A2(\b[50] ), .ZN(new_n8506_));
  NOR2_X1    g08250(.A1(new_n8505_), .A2(new_n8506_), .ZN(new_n8507_));
  XOR2_X1    g08251(.A1(\b[49] ), .A2(\b[50] ), .Z(new_n8508_));
  INV_X1     g08252(.I(new_n8508_), .ZN(new_n8509_));
  AOI21_X1   g08253(.A1(new_n8505_), .A2(new_n8509_), .B(new_n8507_), .ZN(new_n8510_));
  OAI21_X1   g08254(.A1(new_n8510_), .A2(new_n279_), .B(new_n8502_), .ZN(new_n8511_));
  XOR2_X1    g08255(.A1(new_n8511_), .A2(\a[2] ), .Z(new_n8512_));
  INV_X1     g08256(.I(new_n8512_), .ZN(new_n8513_));
  AOI21_X1   g08257(.A1(new_n8109_), .A2(new_n8116_), .B(new_n8468_), .ZN(new_n8514_));
  AOI21_X1   g08258(.A1(new_n8514_), .A2(new_n8465_), .B(new_n8464_), .ZN(new_n8515_));
  AOI22_X1   g08259(.A1(new_n518_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n636_), .ZN(new_n8516_));
  OAI21_X1   g08260(.A1(new_n6490_), .A2(new_n917_), .B(new_n8516_), .ZN(new_n8517_));
  AOI21_X1   g08261(.A1(new_n7906_), .A2(new_n618_), .B(new_n8517_), .ZN(new_n8518_));
  XOR2_X1    g08262(.A1(new_n8518_), .A2(new_n488_), .Z(new_n8519_));
  OAI22_X1   g08263(.A1(new_n713_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n717_), .ZN(new_n8520_));
  AOI21_X1   g08264(.A1(\b[39] ), .A2(new_n1126_), .B(new_n8520_), .ZN(new_n8521_));
  NAND3_X1   g08265(.A1(new_n6298_), .A2(new_n6295_), .A3(new_n724_), .ZN(new_n8522_));
  AOI21_X1   g08266(.A1(new_n8522_), .A2(new_n8521_), .B(new_n722_), .ZN(new_n8523_));
  NAND3_X1   g08267(.A1(new_n8522_), .A2(new_n722_), .A3(new_n8521_), .ZN(new_n8524_));
  INV_X1     g08268(.I(new_n8524_), .ZN(new_n8525_));
  NOR2_X1    g08269(.A1(new_n8525_), .A2(new_n8523_), .ZN(new_n8526_));
  OAI22_X1   g08270(.A1(new_n993_), .A2(new_n5341_), .B1(new_n5312_), .B2(new_n997_), .ZN(new_n8527_));
  AOI21_X1   g08271(.A1(\b[36] ), .A2(new_n1486_), .B(new_n8527_), .ZN(new_n8528_));
  OAI21_X1   g08272(.A1(new_n5352_), .A2(new_n1323_), .B(new_n8528_), .ZN(new_n8529_));
  XOR2_X1    g08273(.A1(new_n8529_), .A2(\a[14] ), .Z(new_n8530_));
  AOI22_X1   g08274(.A1(new_n1586_), .A2(\b[35] ), .B1(\b[34] ), .B2(new_n1495_), .ZN(new_n8531_));
  OAI21_X1   g08275(.A1(new_n4638_), .A2(new_n1917_), .B(new_n8531_), .ZN(new_n8532_));
  INV_X1     g08276(.I(new_n8532_), .ZN(new_n8533_));
  OAI21_X1   g08277(.A1(new_n4676_), .A2(new_n1732_), .B(new_n8533_), .ZN(new_n8534_));
  XOR2_X1    g08278(.A1(new_n8534_), .A2(\a[17] ), .Z(new_n8535_));
  AOI22_X1   g08279(.A1(new_n1738_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n1743_), .ZN(new_n8536_));
  OAI21_X1   g08280(.A1(new_n3624_), .A2(new_n1931_), .B(new_n8536_), .ZN(new_n8537_));
  AOI21_X1   g08281(.A1(new_n4030_), .A2(new_n1746_), .B(new_n8537_), .ZN(new_n8538_));
  XOR2_X1    g08282(.A1(new_n8538_), .A2(new_n1736_), .Z(new_n8539_));
  INV_X1     g08283(.I(new_n8539_), .ZN(new_n8540_));
  AOI22_X1   g08284(.A1(new_n2202_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n2205_), .ZN(new_n8541_));
  OAI21_X1   g08285(.A1(new_n3158_), .A2(new_n2370_), .B(new_n8541_), .ZN(new_n8542_));
  AOI21_X1   g08286(.A1(new_n4188_), .A2(new_n2208_), .B(new_n8542_), .ZN(new_n8543_));
  XOR2_X1    g08287(.A1(new_n8543_), .A2(new_n2200_), .Z(new_n8544_));
  AOI22_X1   g08288(.A1(new_n2716_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n2719_), .ZN(new_n8545_));
  OAI21_X1   g08289(.A1(new_n2495_), .A2(new_n2924_), .B(new_n8545_), .ZN(new_n8546_));
  AOI21_X1   g08290(.A1(new_n3407_), .A2(new_n2722_), .B(new_n8546_), .ZN(new_n8547_));
  XOR2_X1    g08291(.A1(new_n8547_), .A2(new_n2714_), .Z(new_n8548_));
  INV_X1     g08292(.I(new_n8548_), .ZN(new_n8549_));
  AOI22_X1   g08293(.A1(new_n3267_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n3270_), .ZN(new_n8550_));
  OAI21_X1   g08294(.A1(new_n2027_), .A2(new_n3475_), .B(new_n8550_), .ZN(new_n8551_));
  AOI21_X1   g08295(.A1(new_n2470_), .A2(new_n3273_), .B(new_n8551_), .ZN(new_n8552_));
  XOR2_X1    g08296(.A1(new_n8552_), .A2(new_n3264_), .Z(new_n8553_));
  OAI22_X1   g08297(.A1(new_n1432_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n1296_), .ZN(new_n8554_));
  AOI21_X1   g08298(.A1(\b[15] ), .A2(new_n4706_), .B(new_n8554_), .ZN(new_n8555_));
  OAI21_X1   g08299(.A1(new_n1444_), .A2(new_n4458_), .B(new_n8555_), .ZN(new_n8556_));
  XOR2_X1    g08300(.A1(new_n8556_), .A2(\a[35] ), .Z(new_n8557_));
  NAND3_X1   g08301(.A1(new_n8309_), .A2(new_n7982_), .A3(new_n8310_), .ZN(new_n8558_));
  AOI22_X1   g08302(.A1(new_n5155_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n5160_), .ZN(new_n8559_));
  OAI21_X1   g08303(.A1(new_n941_), .A2(new_n6877_), .B(new_n8559_), .ZN(new_n8560_));
  AOI21_X1   g08304(.A1(new_n1449_), .A2(new_n5166_), .B(new_n8560_), .ZN(new_n8561_));
  XOR2_X1    g08305(.A1(new_n8561_), .A2(new_n5162_), .Z(new_n8562_));
  AOI21_X1   g08306(.A1(new_n8293_), .A2(new_n7960_), .B(new_n8295_), .ZN(new_n8563_));
  NAND2_X1   g08307(.A1(new_n8272_), .A2(new_n8277_), .ZN(new_n8564_));
  INV_X1     g08308(.I(new_n6887_), .ZN(new_n8565_));
  AOI22_X1   g08309(.A1(new_n6569_), .A2(\b[8] ), .B1(\b[7] ), .B2(new_n6574_), .ZN(new_n8566_));
  OAI21_X1   g08310(.A1(new_n438_), .A2(new_n8565_), .B(new_n8566_), .ZN(new_n8567_));
  AOI21_X1   g08311(.A1(new_n799_), .A2(new_n6579_), .B(new_n8567_), .ZN(new_n8568_));
  XOR2_X1    g08312(.A1(new_n8568_), .A2(new_n6567_), .Z(new_n8569_));
  INV_X1     g08313(.I(new_n8569_), .ZN(new_n8570_));
  AOI22_X1   g08314(.A1(new_n8241_), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n8246_), .ZN(new_n8571_));
  XOR2_X1    g08315(.A1(\a[47] ), .A2(\a[48] ), .Z(new_n8572_));
  NOR2_X1    g08316(.A1(new_n8249_), .A2(\a[47] ), .ZN(new_n8573_));
  NOR2_X1    g08317(.A1(new_n8250_), .A2(new_n7410_), .ZN(new_n8574_));
  NOR3_X1    g08318(.A1(new_n8573_), .A2(new_n8574_), .A3(new_n8572_), .ZN(new_n8575_));
  NAND2_X1   g08319(.A1(new_n8575_), .A2(\b[0] ), .ZN(new_n8576_));
  NAND2_X1   g08320(.A1(new_n8252_), .A2(new_n554_), .ZN(new_n8577_));
  NAND3_X1   g08321(.A1(new_n8571_), .A2(new_n8576_), .A3(new_n8577_), .ZN(new_n8578_));
  XOR2_X1    g08322(.A1(new_n8578_), .A2(new_n8248_), .Z(new_n8579_));
  NOR3_X1    g08323(.A1(new_n8254_), .A2(new_n8248_), .A3(new_n7937_), .ZN(new_n8580_));
  INV_X1     g08324(.I(new_n8580_), .ZN(new_n8581_));
  NAND2_X1   g08325(.A1(new_n8579_), .A2(new_n8581_), .ZN(new_n8582_));
  OR4_X2     g08326(.A1(new_n8248_), .A2(new_n8578_), .A3(new_n7937_), .A4(new_n8254_), .Z(new_n8583_));
  NAND2_X1   g08327(.A1(new_n8582_), .A2(new_n8583_), .ZN(new_n8584_));
  INV_X1     g08328(.I(new_n7414_), .ZN(new_n8585_));
  XNOR2_X1   g08329(.A1(\a[46] ), .A2(\a[47] ), .ZN(new_n8586_));
  NAND2_X1   g08330(.A1(new_n8586_), .A2(new_n7716_), .ZN(new_n8587_));
  INV_X1     g08331(.I(new_n7408_), .ZN(new_n8588_));
  OAI22_X1   g08332(.A1(new_n339_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n377_), .ZN(new_n8589_));
  AOI21_X1   g08333(.A1(\b[3] ), .A2(new_n7719_), .B(new_n8589_), .ZN(new_n8590_));
  OAI21_X1   g08334(.A1(new_n566_), .A2(new_n8585_), .B(new_n8590_), .ZN(new_n8591_));
  XOR2_X1    g08335(.A1(new_n8591_), .A2(new_n7410_), .Z(new_n8592_));
  NAND2_X1   g08336(.A1(new_n8592_), .A2(new_n8584_), .ZN(new_n8593_));
  XOR2_X1    g08337(.A1(new_n8591_), .A2(\a[47] ), .Z(new_n8594_));
  NAND3_X1   g08338(.A1(new_n8594_), .A2(new_n8582_), .A3(new_n8583_), .ZN(new_n8595_));
  NAND2_X1   g08339(.A1(new_n8595_), .A2(new_n8593_), .ZN(new_n8596_));
  AOI21_X1   g08340(.A1(new_n8268_), .A2(new_n8264_), .B(new_n8263_), .ZN(new_n8597_));
  NOR2_X1    g08341(.A1(new_n8596_), .A2(new_n8597_), .ZN(new_n8598_));
  NAND2_X1   g08342(.A1(new_n8596_), .A2(new_n8597_), .ZN(new_n8599_));
  INV_X1     g08343(.I(new_n8599_), .ZN(new_n8600_));
  OAI21_X1   g08344(.A1(new_n8600_), .A2(new_n8598_), .B(new_n8570_), .ZN(new_n8601_));
  INV_X1     g08345(.I(new_n8598_), .ZN(new_n8602_));
  NAND3_X1   g08346(.A1(new_n8602_), .A2(new_n8599_), .A3(new_n8569_), .ZN(new_n8603_));
  OAI22_X1   g08347(.A1(new_n8232_), .A2(new_n8231_), .B1(new_n8272_), .B2(new_n8277_), .ZN(new_n8604_));
  NAND4_X1   g08348(.A1(new_n8604_), .A2(new_n8564_), .A3(new_n8601_), .A4(new_n8603_), .ZN(new_n8605_));
  AOI22_X1   g08349(.A1(new_n8604_), .A2(new_n8564_), .B1(new_n8601_), .B2(new_n8603_), .ZN(new_n8606_));
  INV_X1     g08350(.I(new_n8606_), .ZN(new_n8607_));
  OAI22_X1   g08351(.A1(new_n5852_), .A2(new_n852_), .B1(new_n776_), .B2(new_n5857_), .ZN(new_n8608_));
  AOI21_X1   g08352(.A1(\b[9] ), .A2(new_n6115_), .B(new_n8608_), .ZN(new_n8609_));
  OAI21_X1   g08353(.A1(new_n859_), .A2(new_n5861_), .B(new_n8609_), .ZN(new_n8610_));
  XOR2_X1    g08354(.A1(new_n8610_), .A2(\a[41] ), .Z(new_n8611_));
  NAND3_X1   g08355(.A1(new_n8607_), .A2(new_n8605_), .A3(new_n8611_), .ZN(new_n8612_));
  INV_X1     g08356(.I(new_n8605_), .ZN(new_n8613_));
  INV_X1     g08357(.I(new_n8611_), .ZN(new_n8614_));
  OAI21_X1   g08358(.A1(new_n8613_), .A2(new_n8606_), .B(new_n8614_), .ZN(new_n8615_));
  NAND2_X1   g08359(.A1(new_n8612_), .A2(new_n8615_), .ZN(new_n8616_));
  NOR3_X1    g08360(.A1(new_n8563_), .A2(new_n8294_), .A3(new_n8616_), .ZN(new_n8617_));
  OAI21_X1   g08361(.A1(new_n8230_), .A2(new_n7964_), .B(new_n8290_), .ZN(new_n8618_));
  AND2_X2    g08362(.A1(new_n8612_), .A2(new_n8615_), .Z(new_n8619_));
  AOI21_X1   g08363(.A1(new_n8618_), .A2(new_n8287_), .B(new_n8619_), .ZN(new_n8620_));
  OAI21_X1   g08364(.A1(new_n8620_), .A2(new_n8617_), .B(new_n8562_), .ZN(new_n8621_));
  INV_X1     g08365(.I(new_n8562_), .ZN(new_n8622_));
  NAND3_X1   g08366(.A1(new_n8618_), .A2(new_n8619_), .A3(new_n8287_), .ZN(new_n8623_));
  OAI21_X1   g08367(.A1(new_n8563_), .A2(new_n8294_), .B(new_n8616_), .ZN(new_n8624_));
  NAND3_X1   g08368(.A1(new_n8623_), .A2(new_n8624_), .A3(new_n8622_), .ZN(new_n8625_));
  NAND2_X1   g08369(.A1(new_n8621_), .A2(new_n8625_), .ZN(new_n8626_));
  AOI21_X1   g08370(.A1(new_n8558_), .A2(new_n8311_), .B(new_n8626_), .ZN(new_n8627_));
  NOR3_X1    g08371(.A1(new_n8229_), .A2(new_n7976_), .A3(new_n8302_), .ZN(new_n8628_));
  AOI21_X1   g08372(.A1(new_n8623_), .A2(new_n8624_), .B(new_n8622_), .ZN(new_n8629_));
  NOR3_X1    g08373(.A1(new_n8620_), .A2(new_n8617_), .A3(new_n8562_), .ZN(new_n8630_));
  NOR2_X1    g08374(.A1(new_n8630_), .A2(new_n8629_), .ZN(new_n8631_));
  NOR3_X1    g08375(.A1(new_n8628_), .A2(new_n8631_), .A3(new_n8306_), .ZN(new_n8632_));
  NOR3_X1    g08376(.A1(new_n8627_), .A2(new_n8632_), .A3(new_n8557_), .ZN(new_n8633_));
  INV_X1     g08377(.I(new_n8557_), .ZN(new_n8634_));
  OAI21_X1   g08378(.A1(new_n8306_), .A2(new_n8628_), .B(new_n8631_), .ZN(new_n8635_));
  NAND3_X1   g08379(.A1(new_n8558_), .A2(new_n8626_), .A3(new_n8311_), .ZN(new_n8636_));
  AOI21_X1   g08380(.A1(new_n8635_), .A2(new_n8636_), .B(new_n8634_), .ZN(new_n8637_));
  NOR2_X1    g08381(.A1(new_n8633_), .A2(new_n8637_), .ZN(new_n8638_));
  OAI21_X1   g08382(.A1(new_n8328_), .A2(new_n8330_), .B(new_n8638_), .ZN(new_n8639_));
  NAND3_X1   g08383(.A1(new_n8635_), .A2(new_n8636_), .A3(new_n8634_), .ZN(new_n8640_));
  OAI21_X1   g08384(.A1(new_n8627_), .A2(new_n8632_), .B(new_n8557_), .ZN(new_n8641_));
  NAND2_X1   g08385(.A1(new_n8641_), .A2(new_n8640_), .ZN(new_n8642_));
  NAND3_X1   g08386(.A1(new_n8335_), .A2(new_n8642_), .A3(new_n8322_), .ZN(new_n8643_));
  AOI22_X1   g08387(.A1(new_n3864_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n3869_), .ZN(new_n8644_));
  OAI21_X1   g08388(.A1(new_n1553_), .A2(new_n5410_), .B(new_n8644_), .ZN(new_n8645_));
  AOI21_X1   g08389(.A1(new_n2452_), .A2(new_n3872_), .B(new_n8645_), .ZN(new_n8646_));
  XOR2_X1    g08390(.A1(new_n8646_), .A2(new_n3876_), .Z(new_n8647_));
  AOI21_X1   g08391(.A1(new_n8639_), .A2(new_n8643_), .B(new_n8647_), .ZN(new_n8648_));
  AOI21_X1   g08392(.A1(new_n8335_), .A2(new_n8322_), .B(new_n8642_), .ZN(new_n8649_));
  NOR3_X1    g08393(.A1(new_n8328_), .A2(new_n8330_), .A3(new_n8638_), .ZN(new_n8650_));
  INV_X1     g08394(.I(new_n8647_), .ZN(new_n8651_));
  NOR3_X1    g08395(.A1(new_n8650_), .A2(new_n8649_), .A3(new_n8651_), .ZN(new_n8652_));
  NOR2_X1    g08396(.A1(new_n8652_), .A2(new_n8648_), .ZN(new_n8653_));
  OAI21_X1   g08397(.A1(new_n8340_), .A2(new_n8342_), .B(new_n8653_), .ZN(new_n8654_));
  OAI21_X1   g08398(.A1(new_n8650_), .A2(new_n8649_), .B(new_n8651_), .ZN(new_n8655_));
  NAND3_X1   g08399(.A1(new_n8639_), .A2(new_n8643_), .A3(new_n8647_), .ZN(new_n8656_));
  NAND2_X1   g08400(.A1(new_n8655_), .A2(new_n8656_), .ZN(new_n8657_));
  NAND3_X1   g08401(.A1(new_n8347_), .A2(new_n8337_), .A3(new_n8657_), .ZN(new_n8658_));
  NAND3_X1   g08402(.A1(new_n8654_), .A2(new_n8658_), .A3(new_n8553_), .ZN(new_n8659_));
  INV_X1     g08403(.I(new_n8553_), .ZN(new_n8660_));
  AOI21_X1   g08404(.A1(new_n8347_), .A2(new_n8337_), .B(new_n8657_), .ZN(new_n8661_));
  NOR3_X1    g08405(.A1(new_n8653_), .A2(new_n8340_), .A3(new_n8342_), .ZN(new_n8662_));
  OAI21_X1   g08406(.A1(new_n8661_), .A2(new_n8662_), .B(new_n8660_), .ZN(new_n8663_));
  NAND2_X1   g08407(.A1(new_n8659_), .A2(new_n8663_), .ZN(new_n8664_));
  AOI21_X1   g08408(.A1(new_n8361_), .A2(new_n8349_), .B(new_n8664_), .ZN(new_n8665_));
  NOR3_X1    g08409(.A1(new_n8661_), .A2(new_n8662_), .A3(new_n8660_), .ZN(new_n8666_));
  AOI21_X1   g08410(.A1(new_n8654_), .A2(new_n8658_), .B(new_n8553_), .ZN(new_n8667_));
  NOR2_X1    g08411(.A1(new_n8667_), .A2(new_n8666_), .ZN(new_n8668_));
  NOR3_X1    g08412(.A1(new_n8354_), .A2(new_n8356_), .A3(new_n8668_), .ZN(new_n8669_));
  NOR3_X1    g08413(.A1(new_n8665_), .A2(new_n8669_), .A3(new_n8549_), .ZN(new_n8670_));
  OAI21_X1   g08414(.A1(new_n8354_), .A2(new_n8356_), .B(new_n8668_), .ZN(new_n8671_));
  NAND3_X1   g08415(.A1(new_n8361_), .A2(new_n8349_), .A3(new_n8664_), .ZN(new_n8672_));
  AOI21_X1   g08416(.A1(new_n8671_), .A2(new_n8672_), .B(new_n8548_), .ZN(new_n8673_));
  NOR2_X1    g08417(.A1(new_n8670_), .A2(new_n8673_), .ZN(new_n8674_));
  OAI21_X1   g08418(.A1(new_n8369_), .A2(new_n8371_), .B(new_n8674_), .ZN(new_n8675_));
  NAND3_X1   g08419(.A1(new_n8671_), .A2(new_n8672_), .A3(new_n8548_), .ZN(new_n8676_));
  OAI21_X1   g08420(.A1(new_n8665_), .A2(new_n8669_), .B(new_n8549_), .ZN(new_n8677_));
  NAND2_X1   g08421(.A1(new_n8677_), .A2(new_n8676_), .ZN(new_n8678_));
  NAND3_X1   g08422(.A1(new_n8377_), .A2(new_n8363_), .A3(new_n8678_), .ZN(new_n8679_));
  NAND3_X1   g08423(.A1(new_n8679_), .A2(new_n8675_), .A3(new_n8544_), .ZN(new_n8680_));
  INV_X1     g08424(.I(new_n8544_), .ZN(new_n8681_));
  AOI21_X1   g08425(.A1(new_n8377_), .A2(new_n8363_), .B(new_n8678_), .ZN(new_n8682_));
  OAI21_X1   g08426(.A1(new_n8026_), .A2(new_n8032_), .B(new_n8037_), .ZN(new_n8683_));
  OAI21_X1   g08427(.A1(new_n8683_), .A2(new_n8364_), .B(new_n8363_), .ZN(new_n8684_));
  NOR2_X1    g08428(.A1(new_n8684_), .A2(new_n8674_), .ZN(new_n8685_));
  OAI21_X1   g08429(.A1(new_n8685_), .A2(new_n8682_), .B(new_n8681_), .ZN(new_n8686_));
  NAND2_X1   g08430(.A1(new_n8686_), .A2(new_n8680_), .ZN(new_n8687_));
  AOI21_X1   g08431(.A1(new_n8386_), .A2(new_n8379_), .B(new_n8687_), .ZN(new_n8688_));
  NOR3_X1    g08432(.A1(new_n8685_), .A2(new_n8682_), .A3(new_n8681_), .ZN(new_n8689_));
  AOI21_X1   g08433(.A1(new_n8679_), .A2(new_n8675_), .B(new_n8544_), .ZN(new_n8690_));
  NOR2_X1    g08434(.A1(new_n8689_), .A2(new_n8690_), .ZN(new_n8691_));
  NOR3_X1    g08435(.A1(new_n8394_), .A2(new_n8691_), .A3(new_n8384_), .ZN(new_n8692_));
  NOR3_X1    g08436(.A1(new_n8688_), .A2(new_n8692_), .A3(new_n8540_), .ZN(new_n8693_));
  OAI21_X1   g08437(.A1(new_n8394_), .A2(new_n8384_), .B(new_n8691_), .ZN(new_n8694_));
  NAND3_X1   g08438(.A1(new_n8386_), .A2(new_n8687_), .A3(new_n8379_), .ZN(new_n8695_));
  AOI21_X1   g08439(.A1(new_n8694_), .A2(new_n8695_), .B(new_n8539_), .ZN(new_n8696_));
  NOR2_X1    g08440(.A1(new_n8693_), .A2(new_n8696_), .ZN(new_n8697_));
  OAI21_X1   g08441(.A1(new_n8410_), .A2(new_n8396_), .B(new_n8697_), .ZN(new_n8698_));
  NAND3_X1   g08442(.A1(new_n8694_), .A2(new_n8695_), .A3(new_n8539_), .ZN(new_n8699_));
  OAI21_X1   g08443(.A1(new_n8688_), .A2(new_n8692_), .B(new_n8540_), .ZN(new_n8700_));
  NAND2_X1   g08444(.A1(new_n8700_), .A2(new_n8699_), .ZN(new_n8701_));
  NAND3_X1   g08445(.A1(new_n8399_), .A2(new_n8701_), .A3(new_n8401_), .ZN(new_n8702_));
  AOI21_X1   g08446(.A1(new_n8698_), .A2(new_n8702_), .B(new_n8535_), .ZN(new_n8703_));
  XOR2_X1    g08447(.A1(new_n8534_), .A2(new_n1344_), .Z(new_n8704_));
  AOI21_X1   g08448(.A1(new_n8399_), .A2(new_n8401_), .B(new_n8701_), .ZN(new_n8705_));
  NOR3_X1    g08449(.A1(new_n8410_), .A2(new_n8697_), .A3(new_n8396_), .ZN(new_n8706_));
  NOR3_X1    g08450(.A1(new_n8706_), .A2(new_n8705_), .A3(new_n8704_), .ZN(new_n8707_));
  NOR2_X1    g08451(.A1(new_n8707_), .A2(new_n8703_), .ZN(new_n8708_));
  OAI21_X1   g08452(.A1(new_n8424_), .A2(new_n8413_), .B(new_n8708_), .ZN(new_n8709_));
  OAI21_X1   g08453(.A1(new_n8706_), .A2(new_n8705_), .B(new_n8704_), .ZN(new_n8710_));
  NAND3_X1   g08454(.A1(new_n8698_), .A2(new_n8702_), .A3(new_n8535_), .ZN(new_n8711_));
  NAND2_X1   g08455(.A1(new_n8710_), .A2(new_n8711_), .ZN(new_n8712_));
  NAND3_X1   g08456(.A1(new_n8416_), .A2(new_n8418_), .A3(new_n8712_), .ZN(new_n8713_));
  AOI21_X1   g08457(.A1(new_n8709_), .A2(new_n8713_), .B(new_n8530_), .ZN(new_n8714_));
  XOR2_X1    g08458(.A1(new_n8529_), .A2(new_n1002_), .Z(new_n8715_));
  AOI21_X1   g08459(.A1(new_n8416_), .A2(new_n8418_), .B(new_n8712_), .ZN(new_n8716_));
  OAI21_X1   g08460(.A1(new_n8075_), .A2(new_n8071_), .B(new_n8077_), .ZN(new_n8717_));
  OAI21_X1   g08461(.A1(new_n8717_), .A2(new_n8419_), .B(new_n8418_), .ZN(new_n8718_));
  NOR2_X1    g08462(.A1(new_n8718_), .A2(new_n8708_), .ZN(new_n8719_));
  NOR3_X1    g08463(.A1(new_n8719_), .A2(new_n8716_), .A3(new_n8715_), .ZN(new_n8720_));
  NOR2_X1    g08464(.A1(new_n8720_), .A2(new_n8714_), .ZN(new_n8721_));
  OAI21_X1   g08465(.A1(new_n8443_), .A2(new_n8426_), .B(new_n8721_), .ZN(new_n8722_));
  OAI21_X1   g08466(.A1(new_n8719_), .A2(new_n8716_), .B(new_n8715_), .ZN(new_n8723_));
  NAND3_X1   g08467(.A1(new_n8709_), .A2(new_n8713_), .A3(new_n8530_), .ZN(new_n8724_));
  NAND2_X1   g08468(.A1(new_n8723_), .A2(new_n8724_), .ZN(new_n8725_));
  NAND3_X1   g08469(.A1(new_n8432_), .A2(new_n8434_), .A3(new_n8725_), .ZN(new_n8726_));
  AOI21_X1   g08470(.A1(new_n8722_), .A2(new_n8726_), .B(new_n8526_), .ZN(new_n8727_));
  INV_X1     g08471(.I(new_n8523_), .ZN(new_n8728_));
  NAND2_X1   g08472(.A1(new_n8728_), .A2(new_n8524_), .ZN(new_n8729_));
  AOI21_X1   g08473(.A1(new_n8432_), .A2(new_n8434_), .B(new_n8725_), .ZN(new_n8730_));
  NOR3_X1    g08474(.A1(new_n8443_), .A2(new_n8721_), .A3(new_n8426_), .ZN(new_n8731_));
  NOR3_X1    g08475(.A1(new_n8730_), .A2(new_n8731_), .A3(new_n8729_), .ZN(new_n8732_));
  NOR2_X1    g08476(.A1(new_n8727_), .A2(new_n8732_), .ZN(new_n8733_));
  OAI21_X1   g08477(.A1(new_n8462_), .A2(new_n8445_), .B(new_n8733_), .ZN(new_n8734_));
  OAI21_X1   g08478(.A1(new_n8730_), .A2(new_n8731_), .B(new_n8729_), .ZN(new_n8735_));
  NAND3_X1   g08479(.A1(new_n8722_), .A2(new_n8726_), .A3(new_n8526_), .ZN(new_n8736_));
  NAND2_X1   g08480(.A1(new_n8736_), .A2(new_n8735_), .ZN(new_n8737_));
  NAND3_X1   g08481(.A1(new_n8451_), .A2(new_n8737_), .A3(new_n8453_), .ZN(new_n8738_));
  NAND3_X1   g08482(.A1(new_n8734_), .A2(new_n8738_), .A3(new_n8519_), .ZN(new_n8739_));
  INV_X1     g08483(.I(new_n8519_), .ZN(new_n8740_));
  AOI21_X1   g08484(.A1(new_n8451_), .A2(new_n8453_), .B(new_n8737_), .ZN(new_n8741_));
  NOR3_X1    g08485(.A1(new_n8462_), .A2(new_n8445_), .A3(new_n8733_), .ZN(new_n8742_));
  OAI21_X1   g08486(.A1(new_n8742_), .A2(new_n8741_), .B(new_n8740_), .ZN(new_n8743_));
  NAND2_X1   g08487(.A1(new_n8743_), .A2(new_n8739_), .ZN(new_n8744_));
  NAND2_X1   g08488(.A1(new_n8515_), .A2(new_n8744_), .ZN(new_n8745_));
  NOR3_X1    g08489(.A1(new_n8742_), .A2(new_n8740_), .A3(new_n8741_), .ZN(new_n8746_));
  AOI21_X1   g08490(.A1(new_n8734_), .A2(new_n8738_), .B(new_n8519_), .ZN(new_n8747_));
  NOR2_X1    g08491(.A1(new_n8746_), .A2(new_n8747_), .ZN(new_n8748_));
  OAI21_X1   g08492(.A1(new_n8477_), .A2(new_n8464_), .B(new_n8748_), .ZN(new_n8749_));
  NAND2_X1   g08493(.A1(new_n8745_), .A2(new_n8749_), .ZN(new_n8750_));
  AOI22_X1   g08494(.A1(new_n800_), .A2(\b[46] ), .B1(\b[47] ), .B2(new_n333_), .ZN(new_n8751_));
  OAI21_X1   g08495(.A1(new_n7096_), .A2(new_n392_), .B(new_n8751_), .ZN(new_n8752_));
  AOI21_X1   g08496(.A1(new_n7649_), .A2(new_n330_), .B(new_n8752_), .ZN(new_n8753_));
  XOR2_X1    g08497(.A1(new_n8753_), .A2(new_n312_), .Z(new_n8754_));
  INV_X1     g08498(.I(new_n8754_), .ZN(new_n8755_));
  AOI21_X1   g08499(.A1(new_n8180_), .A2(new_n8479_), .B(new_n8483_), .ZN(new_n8756_));
  NOR2_X1    g08500(.A1(new_n8756_), .A2(new_n8755_), .ZN(new_n8757_));
  AOI21_X1   g08501(.A1(new_n8124_), .A2(new_n8119_), .B(new_n7930_), .ZN(new_n8758_));
  NAND3_X1   g08502(.A1(new_n8124_), .A2(new_n8119_), .A3(new_n7930_), .ZN(new_n8759_));
  AOI21_X1   g08503(.A1(new_n8149_), .A2(new_n8759_), .B(new_n8758_), .ZN(new_n8760_));
  OAI21_X1   g08504(.A1(new_n8760_), .A2(new_n8480_), .B(new_n8475_), .ZN(new_n8761_));
  NOR2_X1    g08505(.A1(new_n8761_), .A2(new_n8754_), .ZN(new_n8762_));
  NOR3_X1    g08506(.A1(new_n8762_), .A2(new_n8757_), .A3(new_n8750_), .ZN(new_n8763_));
  OAI21_X1   g08507(.A1(new_n8762_), .A2(new_n8757_), .B(new_n8750_), .ZN(new_n8764_));
  INV_X1     g08508(.I(new_n8764_), .ZN(new_n8765_));
  OAI21_X1   g08509(.A1(new_n8765_), .A2(new_n8763_), .B(new_n8513_), .ZN(new_n8766_));
  NOR3_X1    g08510(.A1(new_n8765_), .A2(new_n8513_), .A3(new_n8763_), .ZN(new_n8767_));
  INV_X1     g08511(.I(new_n8767_), .ZN(new_n8768_));
  NAND2_X1   g08512(.A1(new_n8768_), .A2(new_n8766_), .ZN(new_n8769_));
  XOR2_X1    g08513(.A1(new_n8769_), .A2(new_n8499_), .Z(\f[50] ));
  INV_X1     g08514(.I(new_n8498_), .ZN(new_n8771_));
  OAI21_X1   g08515(.A1(new_n8162_), .A2(new_n8487_), .B(new_n8771_), .ZN(new_n8772_));
  OAI21_X1   g08516(.A1(new_n8772_), .A2(new_n8767_), .B(new_n8766_), .ZN(new_n8773_));
  NAND2_X1   g08517(.A1(new_n283_), .A2(\b[49] ), .ZN(new_n8774_));
  AOI22_X1   g08518(.A1(new_n267_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n261_), .ZN(new_n8775_));
  INV_X1     g08519(.I(\b[51] ), .ZN(new_n8776_));
  OAI21_X1   g08520(.A1(new_n8503_), .A2(new_n8504_), .B(new_n8168_), .ZN(new_n8777_));
  NOR2_X1    g08521(.A1(new_n8777_), .A2(new_n8500_), .ZN(new_n8778_));
  NOR3_X1    g08522(.A1(new_n8503_), .A2(new_n8504_), .A3(new_n8168_), .ZN(new_n8779_));
  AOI21_X1   g08523(.A1(new_n8500_), .A2(new_n8779_), .B(new_n8778_), .ZN(new_n8780_));
  NOR2_X1    g08524(.A1(new_n8780_), .A2(new_n8776_), .ZN(new_n8781_));
  AND2_X2    g08525(.A1(new_n8780_), .A2(new_n8776_), .Z(new_n8782_));
  NOR2_X1    g08526(.A1(new_n8782_), .A2(new_n8781_), .ZN(new_n8783_));
  NAND2_X1   g08527(.A1(new_n8783_), .A2(new_n265_), .ZN(new_n8784_));
  NAND3_X1   g08528(.A1(new_n8784_), .A2(new_n8774_), .A3(new_n8775_), .ZN(new_n8785_));
  XOR2_X1    g08529(.A1(new_n8785_), .A2(\a[2] ), .Z(new_n8786_));
  NAND2_X1   g08530(.A1(new_n8180_), .A2(new_n8485_), .ZN(new_n8787_));
  NAND3_X1   g08531(.A1(new_n8787_), .A2(new_n8475_), .A3(new_n8755_), .ZN(new_n8788_));
  OAI21_X1   g08532(.A1(new_n8756_), .A2(new_n8755_), .B(new_n8750_), .ZN(new_n8789_));
  NAND2_X1   g08533(.A1(new_n8789_), .A2(new_n8788_), .ZN(new_n8790_));
  INV_X1     g08534(.I(new_n8790_), .ZN(new_n8791_));
  INV_X1     g08535(.I(new_n8138_), .ZN(new_n8792_));
  AOI22_X1   g08536(.A1(new_n800_), .A2(\b[47] ), .B1(\b[48] ), .B2(new_n333_), .ZN(new_n8793_));
  OAI21_X1   g08537(.A1(new_n7617_), .A2(new_n392_), .B(new_n8793_), .ZN(new_n8794_));
  AOI21_X1   g08538(.A1(new_n8792_), .A2(new_n330_), .B(new_n8794_), .ZN(new_n8795_));
  XOR2_X1    g08539(.A1(new_n8795_), .A2(new_n312_), .Z(new_n8796_));
  INV_X1     g08540(.I(new_n8796_), .ZN(new_n8797_));
  NAND2_X1   g08541(.A1(new_n8575_), .A2(\b[1] ), .ZN(new_n8798_));
  AOI22_X1   g08542(.A1(new_n8241_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n8246_), .ZN(new_n8799_));
  NAND2_X1   g08543(.A1(new_n299_), .A2(new_n8252_), .ZN(new_n8800_));
  NAND3_X1   g08544(.A1(new_n8800_), .A2(new_n8799_), .A3(new_n8798_), .ZN(new_n8801_));
  XOR2_X1    g08545(.A1(new_n8801_), .A2(\a[50] ), .Z(new_n8802_));
  XNOR2_X1   g08546(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n8803_));
  NOR2_X1    g08547(.A1(new_n8803_), .A2(new_n258_), .ZN(new_n8804_));
  NOR2_X1    g08548(.A1(new_n8802_), .A2(new_n8804_), .ZN(new_n8805_));
  INV_X1     g08549(.I(new_n8805_), .ZN(new_n8806_));
  NAND2_X1   g08550(.A1(new_n8802_), .A2(new_n8804_), .ZN(new_n8807_));
  NAND2_X1   g08551(.A1(new_n8806_), .A2(new_n8807_), .ZN(new_n8808_));
  XNOR2_X1   g08552(.A1(new_n8808_), .A2(new_n8583_), .ZN(new_n8809_));
  OAI22_X1   g08553(.A1(new_n377_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n438_), .ZN(new_n8810_));
  AOI21_X1   g08554(.A1(\b[4] ), .A2(new_n7719_), .B(new_n8810_), .ZN(new_n8811_));
  OAI21_X1   g08555(.A1(new_n450_), .A2(new_n8585_), .B(new_n8811_), .ZN(new_n8812_));
  XOR2_X1    g08556(.A1(new_n8812_), .A2(\a[47] ), .Z(new_n8813_));
  INV_X1     g08557(.I(new_n8595_), .ZN(new_n8814_));
  NOR2_X1    g08558(.A1(new_n8598_), .A2(new_n8814_), .ZN(new_n8815_));
  INV_X1     g08559(.I(new_n8815_), .ZN(new_n8816_));
  NAND2_X1   g08560(.A1(new_n8816_), .A2(new_n8813_), .ZN(new_n8817_));
  INV_X1     g08561(.I(new_n8813_), .ZN(new_n8818_));
  NAND2_X1   g08562(.A1(new_n8815_), .A2(new_n8818_), .ZN(new_n8819_));
  NAND3_X1   g08563(.A1(new_n8817_), .A2(new_n8819_), .A3(new_n8809_), .ZN(new_n8820_));
  INV_X1     g08564(.I(new_n8809_), .ZN(new_n8821_));
  NAND2_X1   g08565(.A1(new_n8817_), .A2(new_n8819_), .ZN(new_n8822_));
  NAND2_X1   g08566(.A1(new_n8822_), .A2(new_n8821_), .ZN(new_n8823_));
  NAND2_X1   g08567(.A1(new_n8823_), .A2(new_n8820_), .ZN(new_n8824_));
  AOI22_X1   g08568(.A1(new_n6569_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n6574_), .ZN(new_n8825_));
  OAI21_X1   g08569(.A1(new_n471_), .A2(new_n8565_), .B(new_n8825_), .ZN(new_n8826_));
  AOI21_X1   g08570(.A1(new_n676_), .A2(new_n6579_), .B(new_n8826_), .ZN(new_n8827_));
  XOR2_X1    g08571(.A1(new_n8827_), .A2(new_n6567_), .Z(new_n8828_));
  NAND2_X1   g08572(.A1(new_n8605_), .A2(new_n8603_), .ZN(new_n8829_));
  NAND2_X1   g08573(.A1(new_n8829_), .A2(new_n8828_), .ZN(new_n8830_));
  INV_X1     g08574(.I(new_n8830_), .ZN(new_n8831_));
  NOR2_X1    g08575(.A1(new_n8829_), .A2(new_n8828_), .ZN(new_n8832_));
  NOR3_X1    g08576(.A1(new_n8831_), .A2(new_n8824_), .A3(new_n8832_), .ZN(new_n8833_));
  INV_X1     g08577(.I(new_n8820_), .ZN(new_n8834_));
  AOI21_X1   g08578(.A1(new_n8817_), .A2(new_n8819_), .B(new_n8809_), .ZN(new_n8835_));
  NOR2_X1    g08579(.A1(new_n8834_), .A2(new_n8835_), .ZN(new_n8836_));
  INV_X1     g08580(.I(new_n8832_), .ZN(new_n8837_));
  AOI21_X1   g08581(.A1(new_n8837_), .A2(new_n8830_), .B(new_n8836_), .ZN(new_n8838_));
  NOR2_X1    g08582(.A1(new_n8838_), .A2(new_n8833_), .ZN(new_n8839_));
  AOI22_X1   g08583(.A1(new_n6108_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n6111_), .ZN(new_n8840_));
  OAI21_X1   g08584(.A1(new_n776_), .A2(new_n7708_), .B(new_n8840_), .ZN(new_n8841_));
  AOI21_X1   g08585(.A1(new_n1194_), .A2(new_n6105_), .B(new_n8841_), .ZN(new_n8842_));
  XOR2_X1    g08586(.A1(new_n8842_), .A2(new_n5849_), .Z(new_n8843_));
  NAND2_X1   g08587(.A1(new_n8623_), .A2(new_n8612_), .ZN(new_n8844_));
  NAND2_X1   g08588(.A1(new_n8844_), .A2(new_n8843_), .ZN(new_n8845_));
  INV_X1     g08589(.I(new_n8843_), .ZN(new_n8846_));
  INV_X1     g08590(.I(new_n8612_), .ZN(new_n8847_));
  NOR2_X1    g08591(.A1(new_n8617_), .A2(new_n8847_), .ZN(new_n8848_));
  NAND2_X1   g08592(.A1(new_n8848_), .A2(new_n8846_), .ZN(new_n8849_));
  NAND3_X1   g08593(.A1(new_n8845_), .A2(new_n8849_), .A3(new_n8839_), .ZN(new_n8850_));
  INV_X1     g08594(.I(new_n8839_), .ZN(new_n8851_));
  NOR2_X1    g08595(.A1(new_n8848_), .A2(new_n8846_), .ZN(new_n8852_));
  NOR2_X1    g08596(.A1(new_n8844_), .A2(new_n8843_), .ZN(new_n8853_));
  OAI21_X1   g08597(.A1(new_n8853_), .A2(new_n8852_), .B(new_n8851_), .ZN(new_n8854_));
  NAND2_X1   g08598(.A1(new_n8854_), .A2(new_n8850_), .ZN(new_n8855_));
  OAI22_X1   g08599(.A1(new_n1268_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n1093_), .ZN(new_n8856_));
  AOI21_X1   g08600(.A1(\b[13] ), .A2(new_n5420_), .B(new_n8856_), .ZN(new_n8857_));
  OAI21_X1   g08601(.A1(new_n1275_), .A2(new_n6124_), .B(new_n8857_), .ZN(new_n8858_));
  XOR2_X1    g08602(.A1(new_n8858_), .A2(\a[38] ), .Z(new_n8859_));
  INV_X1     g08603(.I(new_n8859_), .ZN(new_n8860_));
  NAND2_X1   g08604(.A1(new_n8558_), .A2(new_n8311_), .ZN(new_n8861_));
  NOR3_X1    g08605(.A1(new_n8620_), .A2(new_n8617_), .A3(new_n8622_), .ZN(new_n8862_));
  AOI21_X1   g08606(.A1(new_n8861_), .A2(new_n8626_), .B(new_n8862_), .ZN(new_n8863_));
  NOR2_X1    g08607(.A1(new_n8863_), .A2(new_n8860_), .ZN(new_n8864_));
  NOR2_X1    g08608(.A1(new_n8628_), .A2(new_n8306_), .ZN(new_n8865_));
  INV_X1     g08609(.I(new_n8862_), .ZN(new_n8866_));
  OAI21_X1   g08610(.A1(new_n8865_), .A2(new_n8631_), .B(new_n8866_), .ZN(new_n8867_));
  NOR2_X1    g08611(.A1(new_n8867_), .A2(new_n8859_), .ZN(new_n8868_));
  NOR3_X1    g08612(.A1(new_n8864_), .A2(new_n8868_), .A3(new_n8855_), .ZN(new_n8869_));
  NOR3_X1    g08613(.A1(new_n8853_), .A2(new_n8852_), .A3(new_n8851_), .ZN(new_n8870_));
  AOI21_X1   g08614(.A1(new_n8845_), .A2(new_n8849_), .B(new_n8839_), .ZN(new_n8871_));
  NOR2_X1    g08615(.A1(new_n8871_), .A2(new_n8870_), .ZN(new_n8872_));
  NAND2_X1   g08616(.A1(new_n8867_), .A2(new_n8859_), .ZN(new_n8873_));
  NAND2_X1   g08617(.A1(new_n8863_), .A2(new_n8860_), .ZN(new_n8874_));
  AOI21_X1   g08618(.A1(new_n8874_), .A2(new_n8873_), .B(new_n8872_), .ZN(new_n8875_));
  NOR2_X1    g08619(.A1(new_n8875_), .A2(new_n8869_), .ZN(new_n8876_));
  AOI22_X1   g08620(.A1(new_n4918_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n4921_), .ZN(new_n8877_));
  OAI21_X1   g08621(.A1(new_n1296_), .A2(new_n6099_), .B(new_n8877_), .ZN(new_n8878_));
  AOI21_X1   g08622(.A1(new_n2038_), .A2(new_n4699_), .B(new_n8878_), .ZN(new_n8879_));
  XOR2_X1    g08623(.A1(new_n8879_), .A2(new_n4446_), .Z(new_n8880_));
  AOI21_X1   g08624(.A1(new_n7984_), .A2(new_n7989_), .B(new_n7996_), .ZN(new_n8881_));
  AOI21_X1   g08625(.A1(new_n8881_), .A2(new_n8331_), .B(new_n8330_), .ZN(new_n8882_));
  OAI21_X1   g08626(.A1(new_n8882_), .A2(new_n8642_), .B(new_n8641_), .ZN(new_n8883_));
  NAND2_X1   g08627(.A1(new_n8883_), .A2(new_n8880_), .ZN(new_n8884_));
  INV_X1     g08628(.I(new_n8880_), .ZN(new_n8885_));
  NOR2_X1    g08629(.A1(new_n8649_), .A2(new_n8637_), .ZN(new_n8886_));
  NAND2_X1   g08630(.A1(new_n8886_), .A2(new_n8885_), .ZN(new_n8887_));
  NAND3_X1   g08631(.A1(new_n8884_), .A2(new_n8887_), .A3(new_n8876_), .ZN(new_n8888_));
  OR2_X2     g08632(.A1(new_n8875_), .A2(new_n8869_), .Z(new_n8889_));
  NOR2_X1    g08633(.A1(new_n8886_), .A2(new_n8885_), .ZN(new_n8890_));
  NOR2_X1    g08634(.A1(new_n8883_), .A2(new_n8880_), .ZN(new_n8891_));
  OAI21_X1   g08635(.A1(new_n8891_), .A2(new_n8890_), .B(new_n8889_), .ZN(new_n8892_));
  NAND2_X1   g08636(.A1(new_n8892_), .A2(new_n8888_), .ZN(new_n8893_));
  AOI22_X1   g08637(.A1(new_n3864_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n3869_), .ZN(new_n8894_));
  OAI21_X1   g08638(.A1(new_n1859_), .A2(new_n5410_), .B(new_n8894_), .ZN(new_n8895_));
  AOI21_X1   g08639(.A1(new_n2032_), .A2(new_n3872_), .B(new_n8895_), .ZN(new_n8896_));
  XOR2_X1    g08640(.A1(new_n8896_), .A2(new_n3876_), .Z(new_n8897_));
  INV_X1     g08641(.I(new_n8897_), .ZN(new_n8898_));
  AOI21_X1   g08642(.A1(new_n8654_), .A2(new_n8656_), .B(new_n8898_), .ZN(new_n8899_));
  NOR3_X1    g08643(.A1(new_n8661_), .A2(new_n8652_), .A3(new_n8897_), .ZN(new_n8900_));
  NOR3_X1    g08644(.A1(new_n8899_), .A2(new_n8900_), .A3(new_n8893_), .ZN(new_n8901_));
  INV_X1     g08645(.I(new_n8893_), .ZN(new_n8902_));
  OAI21_X1   g08646(.A1(new_n8661_), .A2(new_n8652_), .B(new_n8897_), .ZN(new_n8903_));
  NAND3_X1   g08647(.A1(new_n8654_), .A2(new_n8656_), .A3(new_n8898_), .ZN(new_n8904_));
  AOI21_X1   g08648(.A1(new_n8903_), .A2(new_n8904_), .B(new_n8902_), .ZN(new_n8905_));
  OR2_X2     g08649(.A1(new_n8901_), .A2(new_n8905_), .Z(new_n8906_));
  AOI22_X1   g08650(.A1(new_n3267_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n3270_), .ZN(new_n8907_));
  OAI21_X1   g08651(.A1(new_n2142_), .A2(new_n3475_), .B(new_n8907_), .ZN(new_n8908_));
  AOI21_X1   g08652(.A1(new_n3033_), .A2(new_n3273_), .B(new_n8908_), .ZN(new_n8909_));
  XOR2_X1    g08653(.A1(new_n8909_), .A2(new_n3264_), .Z(new_n8910_));
  INV_X1     g08654(.I(new_n8910_), .ZN(new_n8911_));
  AOI21_X1   g08655(.A1(new_n8671_), .A2(new_n8659_), .B(new_n8911_), .ZN(new_n8912_));
  NOR3_X1    g08656(.A1(new_n8665_), .A2(new_n8666_), .A3(new_n8910_), .ZN(new_n8913_));
  NOR3_X1    g08657(.A1(new_n8913_), .A2(new_n8912_), .A3(new_n8906_), .ZN(new_n8914_));
  NOR2_X1    g08658(.A1(new_n8901_), .A2(new_n8905_), .ZN(new_n8915_));
  OAI21_X1   g08659(.A1(new_n8665_), .A2(new_n8666_), .B(new_n8910_), .ZN(new_n8916_));
  NAND3_X1   g08660(.A1(new_n8671_), .A2(new_n8659_), .A3(new_n8911_), .ZN(new_n8917_));
  AOI21_X1   g08661(.A1(new_n8916_), .A2(new_n8917_), .B(new_n8915_), .ZN(new_n8918_));
  OR2_X2     g08662(.A1(new_n8914_), .A2(new_n8918_), .Z(new_n8919_));
  OAI22_X1   g08663(.A1(new_n2703_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n2708_), .ZN(new_n8920_));
  AOI21_X1   g08664(.A1(\b[25] ), .A2(new_n2906_), .B(new_n8920_), .ZN(new_n8921_));
  OAI21_X1   g08665(.A1(new_n3165_), .A2(new_n2711_), .B(new_n8921_), .ZN(new_n8922_));
  XOR2_X1    g08666(.A1(new_n8922_), .A2(\a[26] ), .Z(new_n8923_));
  AOI21_X1   g08667(.A1(new_n8373_), .A2(new_n8372_), .B(new_n8371_), .ZN(new_n8924_));
  OAI21_X1   g08668(.A1(new_n8924_), .A2(new_n8678_), .B(new_n8676_), .ZN(new_n8925_));
  NAND2_X1   g08669(.A1(new_n8925_), .A2(new_n8923_), .ZN(new_n8926_));
  INV_X1     g08670(.I(new_n8923_), .ZN(new_n8927_));
  NAND3_X1   g08671(.A1(new_n8675_), .A2(new_n8676_), .A3(new_n8927_), .ZN(new_n8928_));
  NAND2_X1   g08672(.A1(new_n8926_), .A2(new_n8928_), .ZN(new_n8929_));
  XOR2_X1    g08673(.A1(new_n8929_), .A2(new_n8919_), .Z(new_n8930_));
  AOI22_X1   g08674(.A1(new_n2202_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n2205_), .ZN(new_n8931_));
  OAI21_X1   g08675(.A1(new_n3185_), .A2(new_n2370_), .B(new_n8931_), .ZN(new_n8932_));
  AOI21_X1   g08676(.A1(new_n4230_), .A2(new_n2208_), .B(new_n8932_), .ZN(new_n8933_));
  XOR2_X1    g08677(.A1(new_n8933_), .A2(new_n2200_), .Z(new_n8934_));
  OAI21_X1   g08678(.A1(new_n8688_), .A2(new_n8689_), .B(new_n8934_), .ZN(new_n8935_));
  INV_X1     g08679(.I(new_n8934_), .ZN(new_n8936_));
  NAND3_X1   g08680(.A1(new_n8694_), .A2(new_n8680_), .A3(new_n8936_), .ZN(new_n8937_));
  NAND3_X1   g08681(.A1(new_n8937_), .A2(new_n8935_), .A3(new_n8930_), .ZN(new_n8938_));
  NOR2_X1    g08682(.A1(new_n8914_), .A2(new_n8918_), .ZN(new_n8939_));
  NAND3_X1   g08683(.A1(new_n8926_), .A2(new_n8928_), .A3(new_n8939_), .ZN(new_n8940_));
  NAND2_X1   g08684(.A1(new_n8929_), .A2(new_n8919_), .ZN(new_n8941_));
  NAND2_X1   g08685(.A1(new_n8941_), .A2(new_n8940_), .ZN(new_n8942_));
  AOI21_X1   g08686(.A1(new_n8694_), .A2(new_n8680_), .B(new_n8936_), .ZN(new_n8943_));
  AOI21_X1   g08687(.A1(new_n8392_), .A2(new_n8385_), .B(new_n8384_), .ZN(new_n8944_));
  OAI21_X1   g08688(.A1(new_n8944_), .A2(new_n8687_), .B(new_n8680_), .ZN(new_n8945_));
  NOR2_X1    g08689(.A1(new_n8945_), .A2(new_n8934_), .ZN(new_n8946_));
  OAI21_X1   g08690(.A1(new_n8946_), .A2(new_n8943_), .B(new_n8942_), .ZN(new_n8947_));
  NAND2_X1   g08691(.A1(new_n8947_), .A2(new_n8938_), .ZN(new_n8948_));
  INV_X1     g08692(.I(new_n8948_), .ZN(new_n8949_));
  AOI22_X1   g08693(.A1(new_n1738_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n1743_), .ZN(new_n8950_));
  OAI21_X1   g08694(.A1(new_n4022_), .A2(new_n1931_), .B(new_n8950_), .ZN(new_n8951_));
  AOI21_X1   g08695(.A1(new_n4223_), .A2(new_n1746_), .B(new_n8951_), .ZN(new_n8952_));
  XOR2_X1    g08696(.A1(new_n8952_), .A2(new_n1736_), .Z(new_n8953_));
  AOI21_X1   g08697(.A1(new_n8411_), .A2(new_n8397_), .B(new_n8396_), .ZN(new_n8954_));
  OAI21_X1   g08698(.A1(new_n8954_), .A2(new_n8701_), .B(new_n8699_), .ZN(new_n8955_));
  NAND2_X1   g08699(.A1(new_n8955_), .A2(new_n8953_), .ZN(new_n8956_));
  INV_X1     g08700(.I(new_n8953_), .ZN(new_n8957_));
  NAND3_X1   g08701(.A1(new_n8698_), .A2(new_n8699_), .A3(new_n8957_), .ZN(new_n8958_));
  NAND3_X1   g08702(.A1(new_n8956_), .A2(new_n8958_), .A3(new_n8949_), .ZN(new_n8959_));
  AOI21_X1   g08703(.A1(new_n8956_), .A2(new_n8958_), .B(new_n8949_), .ZN(new_n8960_));
  INV_X1     g08704(.I(new_n8960_), .ZN(new_n8961_));
  NAND2_X1   g08705(.A1(new_n8961_), .A2(new_n8959_), .ZN(new_n8962_));
  OAI22_X1   g08706(.A1(new_n1592_), .A2(new_n4886_), .B1(new_n4666_), .B2(new_n1505_), .ZN(new_n8963_));
  AOI21_X1   g08707(.A1(\b[34] ), .A2(new_n1584_), .B(new_n8963_), .ZN(new_n8964_));
  OAI21_X1   g08708(.A1(new_n4898_), .A2(new_n1732_), .B(new_n8964_), .ZN(new_n8965_));
  XOR2_X1    g08709(.A1(new_n8965_), .A2(\a[17] ), .Z(new_n8966_));
  INV_X1     g08710(.I(new_n8966_), .ZN(new_n8967_));
  AOI21_X1   g08711(.A1(new_n8709_), .A2(new_n8711_), .B(new_n8967_), .ZN(new_n8968_));
  NOR3_X1    g08712(.A1(new_n8716_), .A2(new_n8707_), .A3(new_n8966_), .ZN(new_n8969_));
  NOR3_X1    g08713(.A1(new_n8969_), .A2(new_n8968_), .A3(new_n8962_), .ZN(new_n8970_));
  OAI21_X1   g08714(.A1(new_n8969_), .A2(new_n8968_), .B(new_n8962_), .ZN(new_n8971_));
  INV_X1     g08715(.I(new_n8971_), .ZN(new_n8972_));
  NOR2_X1    g08716(.A1(new_n8972_), .A2(new_n8970_), .ZN(new_n8973_));
  OAI22_X1   g08717(.A1(new_n993_), .A2(new_n5761_), .B1(new_n5341_), .B2(new_n997_), .ZN(new_n8974_));
  AOI21_X1   g08718(.A1(\b[37] ), .A2(new_n1486_), .B(new_n8974_), .ZN(new_n8975_));
  OAI21_X1   g08719(.A1(new_n6309_), .A2(new_n1323_), .B(new_n8975_), .ZN(new_n8976_));
  XOR2_X1    g08720(.A1(new_n8976_), .A2(\a[14] ), .Z(new_n8977_));
  OAI21_X1   g08721(.A1(new_n8730_), .A2(new_n8720_), .B(new_n8977_), .ZN(new_n8978_));
  INV_X1     g08722(.I(new_n8977_), .ZN(new_n8979_));
  NAND3_X1   g08723(.A1(new_n8722_), .A2(new_n8724_), .A3(new_n8979_), .ZN(new_n8980_));
  NAND3_X1   g08724(.A1(new_n8978_), .A2(new_n8980_), .A3(new_n8973_), .ZN(new_n8981_));
  INV_X1     g08725(.I(new_n8970_), .ZN(new_n8982_));
  NAND2_X1   g08726(.A1(new_n8982_), .A2(new_n8971_), .ZN(new_n8983_));
  AOI21_X1   g08727(.A1(new_n8722_), .A2(new_n8724_), .B(new_n8979_), .ZN(new_n8984_));
  NOR3_X1    g08728(.A1(new_n8730_), .A2(new_n8720_), .A3(new_n8977_), .ZN(new_n8985_));
  OAI21_X1   g08729(.A1(new_n8985_), .A2(new_n8984_), .B(new_n8983_), .ZN(new_n8986_));
  NAND2_X1   g08730(.A1(new_n8986_), .A2(new_n8981_), .ZN(new_n8987_));
  INV_X1     g08731(.I(new_n7106_), .ZN(new_n8988_));
  OAI22_X1   g08732(.A1(new_n713_), .A2(new_n6490_), .B1(new_n6285_), .B2(new_n717_), .ZN(new_n8989_));
  AOI21_X1   g08733(.A1(\b[40] ), .A2(new_n1126_), .B(new_n8989_), .ZN(new_n8990_));
  OAI21_X1   g08734(.A1(new_n8988_), .A2(new_n986_), .B(new_n8990_), .ZN(new_n8991_));
  XOR2_X1    g08735(.A1(new_n8991_), .A2(\a[11] ), .Z(new_n8992_));
  INV_X1     g08736(.I(new_n8992_), .ZN(new_n8993_));
  AOI21_X1   g08737(.A1(new_n8734_), .A2(new_n8736_), .B(new_n8993_), .ZN(new_n8994_));
  NOR3_X1    g08738(.A1(new_n8741_), .A2(new_n8732_), .A3(new_n8992_), .ZN(new_n8995_));
  NOR3_X1    g08739(.A1(new_n8994_), .A2(new_n8995_), .A3(new_n8987_), .ZN(new_n8996_));
  INV_X1     g08740(.I(new_n8987_), .ZN(new_n8997_));
  OAI21_X1   g08741(.A1(new_n8741_), .A2(new_n8732_), .B(new_n8992_), .ZN(new_n8998_));
  NAND3_X1   g08742(.A1(new_n8734_), .A2(new_n8736_), .A3(new_n8993_), .ZN(new_n8999_));
  AOI21_X1   g08743(.A1(new_n8999_), .A2(new_n8998_), .B(new_n8997_), .ZN(new_n9000_));
  NOR2_X1    g08744(.A1(new_n8996_), .A2(new_n9000_), .ZN(new_n9001_));
  AOI21_X1   g08745(.A1(new_n8467_), .A2(new_n8470_), .B(new_n8744_), .ZN(new_n9002_));
  AOI22_X1   g08746(.A1(new_n518_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n636_), .ZN(new_n9003_));
  OAI21_X1   g08747(.A1(new_n6775_), .A2(new_n917_), .B(new_n9003_), .ZN(new_n9004_));
  AOI21_X1   g08748(.A1(new_n7926_), .A2(new_n618_), .B(new_n9004_), .ZN(new_n9005_));
  XOR2_X1    g08749(.A1(new_n9005_), .A2(new_n488_), .Z(new_n9006_));
  OAI21_X1   g08750(.A1(new_n9002_), .A2(new_n8746_), .B(new_n9006_), .ZN(new_n9007_));
  INV_X1     g08751(.I(new_n9006_), .ZN(new_n9008_));
  NAND3_X1   g08752(.A1(new_n8749_), .A2(new_n8739_), .A3(new_n9008_), .ZN(new_n9009_));
  NAND3_X1   g08753(.A1(new_n9007_), .A2(new_n9009_), .A3(new_n9001_), .ZN(new_n9010_));
  OR2_X2     g08754(.A1(new_n8996_), .A2(new_n9000_), .Z(new_n9011_));
  AOI21_X1   g08755(.A1(new_n8749_), .A2(new_n8739_), .B(new_n9008_), .ZN(new_n9012_));
  NOR3_X1    g08756(.A1(new_n9002_), .A2(new_n8746_), .A3(new_n9006_), .ZN(new_n9013_));
  OAI21_X1   g08757(.A1(new_n9013_), .A2(new_n9012_), .B(new_n9011_), .ZN(new_n9014_));
  AOI21_X1   g08758(.A1(new_n9014_), .A2(new_n9010_), .B(new_n8797_), .ZN(new_n9015_));
  NOR3_X1    g08759(.A1(new_n9013_), .A2(new_n9012_), .A3(new_n9011_), .ZN(new_n9016_));
  AOI21_X1   g08760(.A1(new_n9007_), .A2(new_n9009_), .B(new_n9001_), .ZN(new_n9017_));
  NOR3_X1    g08761(.A1(new_n9016_), .A2(new_n9017_), .A3(new_n8796_), .ZN(new_n9018_));
  NOR3_X1    g08762(.A1(new_n8791_), .A2(new_n9015_), .A3(new_n9018_), .ZN(new_n9019_));
  INV_X1     g08763(.I(new_n9015_), .ZN(new_n9020_));
  NAND3_X1   g08764(.A1(new_n9014_), .A2(new_n9010_), .A3(new_n8797_), .ZN(new_n9021_));
  AOI21_X1   g08765(.A1(new_n9020_), .A2(new_n9021_), .B(new_n8790_), .ZN(new_n9022_));
  OAI21_X1   g08766(.A1(new_n9019_), .A2(new_n9022_), .B(new_n8786_), .ZN(new_n9023_));
  NOR3_X1    g08767(.A1(new_n9019_), .A2(new_n8786_), .A3(new_n9022_), .ZN(new_n9024_));
  INV_X1     g08768(.I(new_n9024_), .ZN(new_n9025_));
  NAND2_X1   g08769(.A1(new_n9025_), .A2(new_n9023_), .ZN(new_n9026_));
  XOR2_X1    g08770(.A1(new_n9026_), .A2(new_n8773_), .Z(\f[51] ));
  INV_X1     g08771(.I(new_n8766_), .ZN(new_n9028_));
  AOI21_X1   g08772(.A1(new_n8499_), .A2(new_n8768_), .B(new_n9028_), .ZN(new_n9029_));
  INV_X1     g08773(.I(new_n9023_), .ZN(new_n9030_));
  AOI21_X1   g08774(.A1(new_n9029_), .A2(new_n9025_), .B(new_n9030_), .ZN(new_n9031_));
  INV_X1     g08775(.I(\b[52] ), .ZN(new_n9032_));
  OAI22_X1   g08776(.A1(new_n277_), .A2(new_n9032_), .B1(new_n8776_), .B2(new_n262_), .ZN(new_n9033_));
  AOI21_X1   g08777(.A1(\b[50] ), .A2(new_n283_), .B(new_n9033_), .ZN(new_n9034_));
  XOR2_X1    g08778(.A1(\b[51] ), .A2(\b[52] ), .Z(new_n9035_));
  INV_X1     g08779(.I(new_n9035_), .ZN(new_n9036_));
  OAI21_X1   g08780(.A1(new_n8779_), .A2(\b[50] ), .B(\b[51] ), .ZN(new_n9037_));
  NAND2_X1   g08781(.A1(new_n8777_), .A2(\b[50] ), .ZN(new_n9038_));
  NAND2_X1   g08782(.A1(new_n9037_), .A2(new_n9038_), .ZN(new_n9039_));
  NAND2_X1   g08783(.A1(new_n9039_), .A2(new_n9036_), .ZN(new_n9040_));
  INV_X1     g08784(.I(new_n9040_), .ZN(new_n9041_));
  NOR2_X1    g08785(.A1(new_n9039_), .A2(new_n9036_), .ZN(new_n9042_));
  NOR2_X1    g08786(.A1(new_n9041_), .A2(new_n9042_), .ZN(new_n9043_));
  OAI21_X1   g08787(.A1(new_n9043_), .A2(new_n279_), .B(new_n9034_), .ZN(new_n9044_));
  XOR2_X1    g08788(.A1(new_n9044_), .A2(\a[2] ), .Z(new_n9045_));
  INV_X1     g08789(.I(new_n9045_), .ZN(new_n9046_));
  INV_X1     g08790(.I(new_n8750_), .ZN(new_n9047_));
  AOI21_X1   g08791(.A1(new_n8761_), .A2(new_n8754_), .B(new_n9047_), .ZN(new_n9048_));
  NOR3_X1    g08792(.A1(new_n9048_), .A2(new_n9018_), .A3(new_n8762_), .ZN(new_n9049_));
  NAND2_X1   g08793(.A1(new_n8173_), .A2(new_n8172_), .ZN(new_n9050_));
  OAI22_X1   g08794(.A1(new_n321_), .A2(new_n8168_), .B1(new_n325_), .B2(new_n8127_), .ZN(new_n9051_));
  AOI21_X1   g08795(.A1(\b[47] ), .A2(new_n602_), .B(new_n9051_), .ZN(new_n9052_));
  OAI21_X1   g08796(.A1(new_n9050_), .A2(new_n318_), .B(new_n9052_), .ZN(new_n9053_));
  XOR2_X1    g08797(.A1(new_n9053_), .A2(\a[5] ), .Z(new_n9054_));
  INV_X1     g08798(.I(new_n9054_), .ZN(new_n9055_));
  AOI21_X1   g08799(.A1(new_n8095_), .A2(new_n8100_), .B(new_n8106_), .ZN(new_n9056_));
  AOI21_X1   g08800(.A1(new_n9056_), .A2(new_n8446_), .B(new_n8445_), .ZN(new_n9057_));
  OAI21_X1   g08801(.A1(new_n9057_), .A2(new_n8737_), .B(new_n8736_), .ZN(new_n9058_));
  AOI21_X1   g08802(.A1(new_n9058_), .A2(new_n8992_), .B(new_n8987_), .ZN(new_n9059_));
  OAI22_X1   g08803(.A1(new_n713_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n717_), .ZN(new_n9060_));
  AOI21_X1   g08804(.A1(\b[41] ), .A2(new_n1126_), .B(new_n9060_), .ZN(new_n9061_));
  OAI21_X1   g08805(.A1(new_n6785_), .A2(new_n986_), .B(new_n9061_), .ZN(new_n9062_));
  XOR2_X1    g08806(.A1(new_n9062_), .A2(new_n722_), .Z(new_n9063_));
  AOI21_X1   g08807(.A1(new_n8091_), .A2(new_n8092_), .B(new_n8087_), .ZN(new_n9064_));
  AOI21_X1   g08808(.A1(new_n9064_), .A2(new_n8427_), .B(new_n8426_), .ZN(new_n9065_));
  OAI21_X1   g08809(.A1(new_n9065_), .A2(new_n8725_), .B(new_n8724_), .ZN(new_n9066_));
  AOI21_X1   g08810(.A1(new_n9066_), .A2(new_n8977_), .B(new_n8983_), .ZN(new_n9067_));
  OAI22_X1   g08811(.A1(new_n993_), .A2(new_n6284_), .B1(new_n5761_), .B2(new_n997_), .ZN(new_n9068_));
  AOI21_X1   g08812(.A1(\b[38] ), .A2(new_n1486_), .B(new_n9068_), .ZN(new_n9069_));
  OAI21_X1   g08813(.A1(new_n8195_), .A2(new_n1323_), .B(new_n9069_), .ZN(new_n9070_));
  XOR2_X1    g08814(.A1(new_n9070_), .A2(\a[14] ), .Z(new_n9071_));
  NAND3_X1   g08815(.A1(new_n8709_), .A2(new_n8711_), .A3(new_n8967_), .ZN(new_n9072_));
  INV_X1     g08816(.I(new_n8959_), .ZN(new_n9073_));
  NOR2_X1    g08817(.A1(new_n9073_), .A2(new_n8960_), .ZN(new_n9074_));
  AOI21_X1   g08818(.A1(new_n8718_), .A2(new_n8708_), .B(new_n8707_), .ZN(new_n9075_));
  OAI21_X1   g08819(.A1(new_n9075_), .A2(new_n8967_), .B(new_n9074_), .ZN(new_n9076_));
  OAI22_X1   g08820(.A1(new_n1592_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n1505_), .ZN(new_n9077_));
  AOI21_X1   g08821(.A1(\b[35] ), .A2(new_n1584_), .B(new_n9077_), .ZN(new_n9078_));
  OAI21_X1   g08822(.A1(new_n5322_), .A2(new_n1732_), .B(new_n9078_), .ZN(new_n9079_));
  XOR2_X1    g08823(.A1(new_n9079_), .A2(\a[17] ), .Z(new_n9080_));
  NOR2_X1    g08824(.A1(new_n8955_), .A2(new_n8953_), .ZN(new_n9081_));
  AOI21_X1   g08825(.A1(new_n8955_), .A2(new_n8953_), .B(new_n8948_), .ZN(new_n9082_));
  AOI22_X1   g08826(.A1(new_n1738_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n1743_), .ZN(new_n9083_));
  OAI21_X1   g08827(.A1(new_n4023_), .A2(new_n1931_), .B(new_n9083_), .ZN(new_n9084_));
  AOI21_X1   g08828(.A1(new_n5103_), .A2(new_n1746_), .B(new_n9084_), .ZN(new_n9085_));
  XOR2_X1    g08829(.A1(new_n9085_), .A2(new_n1736_), .Z(new_n9086_));
  NAND2_X1   g08830(.A1(new_n8935_), .A2(new_n8930_), .ZN(new_n9087_));
  AOI22_X1   g08831(.A1(new_n2202_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n2205_), .ZN(new_n9088_));
  OAI21_X1   g08832(.A1(new_n3592_), .A2(new_n2370_), .B(new_n9088_), .ZN(new_n9089_));
  AOI21_X1   g08833(.A1(new_n3796_), .A2(new_n2208_), .B(new_n9089_), .ZN(new_n9090_));
  XOR2_X1    g08834(.A1(new_n9090_), .A2(new_n2200_), .Z(new_n9091_));
  NOR2_X1    g08835(.A1(new_n8925_), .A2(new_n8923_), .ZN(new_n9092_));
  AOI21_X1   g08836(.A1(new_n8925_), .A2(new_n8923_), .B(new_n8919_), .ZN(new_n9093_));
  NAND2_X1   g08837(.A1(new_n8916_), .A2(new_n8915_), .ZN(new_n9094_));
  OAI22_X1   g08838(.A1(new_n2646_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n2495_), .ZN(new_n9095_));
  AOI21_X1   g08839(.A1(\b[23] ), .A2(new_n3456_), .B(new_n9095_), .ZN(new_n9096_));
  OAI21_X1   g08840(.A1(new_n2655_), .A2(new_n3261_), .B(new_n9096_), .ZN(new_n9097_));
  XOR2_X1    g08841(.A1(new_n9097_), .A2(\a[29] ), .Z(new_n9098_));
  AOI22_X1   g08842(.A1(new_n3864_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n3869_), .ZN(new_n9099_));
  OAI21_X1   g08843(.A1(new_n1860_), .A2(new_n5410_), .B(new_n9099_), .ZN(new_n9100_));
  AOI21_X1   g08844(.A1(new_n2659_), .A2(new_n3872_), .B(new_n9100_), .ZN(new_n9101_));
  XOR2_X1    g08845(.A1(new_n9101_), .A2(new_n3876_), .Z(new_n9102_));
  OAI21_X1   g08846(.A1(new_n8886_), .A2(new_n8885_), .B(new_n8876_), .ZN(new_n9103_));
  AOI21_X1   g08847(.A1(new_n8867_), .A2(new_n8859_), .B(new_n8855_), .ZN(new_n9104_));
  NOR2_X1    g08848(.A1(new_n9104_), .A2(new_n8868_), .ZN(new_n9105_));
  AOI22_X1   g08849(.A1(new_n5155_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n5160_), .ZN(new_n9106_));
  OAI21_X1   g08850(.A1(new_n1093_), .A2(new_n6877_), .B(new_n9106_), .ZN(new_n9107_));
  AOI21_X1   g08851(.A1(new_n1701_), .A2(new_n5166_), .B(new_n9107_), .ZN(new_n9108_));
  XOR2_X1    g08852(.A1(new_n9108_), .A2(new_n5162_), .Z(new_n9109_));
  INV_X1     g08853(.I(new_n9109_), .ZN(new_n9110_));
  OAI21_X1   g08854(.A1(new_n8848_), .A2(new_n8846_), .B(new_n8839_), .ZN(new_n9111_));
  NAND2_X1   g08855(.A1(new_n8830_), .A2(new_n8836_), .ZN(new_n9112_));
  OAI21_X1   g08856(.A1(new_n8815_), .A2(new_n8818_), .B(new_n8809_), .ZN(new_n9113_));
  INV_X1     g08857(.I(new_n8575_), .ZN(new_n9114_));
  AOI22_X1   g08858(.A1(new_n8241_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n8246_), .ZN(new_n9115_));
  OAI21_X1   g08859(.A1(new_n276_), .A2(new_n9114_), .B(new_n9115_), .ZN(new_n9116_));
  AOI21_X1   g08860(.A1(new_n1725_), .A2(new_n8252_), .B(new_n9116_), .ZN(new_n9117_));
  XOR2_X1    g08861(.A1(new_n9117_), .A2(\a[50] ), .Z(new_n9118_));
  INV_X1     g08862(.I(\a[51] ), .ZN(new_n9119_));
  NAND3_X1   g08863(.A1(new_n8248_), .A2(new_n9119_), .A3(\a[52] ), .ZN(new_n9120_));
  INV_X1     g08864(.I(\a[52] ), .ZN(new_n9121_));
  NAND3_X1   g08865(.A1(new_n9121_), .A2(\a[50] ), .A3(\a[51] ), .ZN(new_n9122_));
  NAND2_X1   g08866(.A1(new_n9120_), .A2(new_n9122_), .ZN(new_n9123_));
  XOR2_X1    g08867(.A1(\a[52] ), .A2(\a[53] ), .Z(new_n9124_));
  NOR2_X1    g08868(.A1(new_n8803_), .A2(new_n9124_), .ZN(new_n9125_));
  AOI22_X1   g08869(.A1(new_n9125_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n9123_), .ZN(new_n9126_));
  XOR2_X1    g08870(.A1(\a[52] ), .A2(\a[53] ), .Z(new_n9127_));
  INV_X1     g08871(.I(new_n9127_), .ZN(new_n9128_));
  NOR2_X1    g08872(.A1(new_n9128_), .A2(new_n8803_), .ZN(new_n9129_));
  NAND2_X1   g08873(.A1(new_n9129_), .A2(new_n263_), .ZN(new_n9130_));
  NAND2_X1   g08874(.A1(new_n9130_), .A2(new_n9126_), .ZN(new_n9131_));
  NAND2_X1   g08875(.A1(new_n9131_), .A2(\a[53] ), .ZN(new_n9132_));
  INV_X1     g08876(.I(\a[53] ), .ZN(new_n9133_));
  XOR2_X1    g08877(.A1(new_n9131_), .A2(new_n9133_), .Z(new_n9134_));
  NOR2_X1    g08878(.A1(new_n8804_), .A2(new_n9133_), .ZN(new_n9135_));
  OAI22_X1   g08879(.A1(new_n9134_), .A2(new_n9135_), .B1(new_n8804_), .B2(new_n9132_), .ZN(new_n9136_));
  AOI21_X1   g08880(.A1(new_n8583_), .A2(new_n8807_), .B(new_n8805_), .ZN(new_n9137_));
  XOR2_X1    g08881(.A1(new_n9137_), .A2(new_n9136_), .Z(new_n9138_));
  NAND2_X1   g08882(.A1(new_n9138_), .A2(new_n9118_), .ZN(new_n9139_));
  INV_X1     g08883(.I(new_n9118_), .ZN(new_n9140_));
  NAND2_X1   g08884(.A1(new_n9137_), .A2(new_n9136_), .ZN(new_n9141_));
  OR2_X2     g08885(.A1(new_n9137_), .A2(new_n9136_), .Z(new_n9142_));
  NAND2_X1   g08886(.A1(new_n9142_), .A2(new_n9141_), .ZN(new_n9143_));
  NAND2_X1   g08887(.A1(new_n9143_), .A2(new_n9140_), .ZN(new_n9144_));
  OAI22_X1   g08888(.A1(new_n438_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n471_), .ZN(new_n9145_));
  AOI21_X1   g08889(.A1(\b[5] ), .A2(new_n7719_), .B(new_n9145_), .ZN(new_n9146_));
  OAI21_X1   g08890(.A1(new_n485_), .A2(new_n8585_), .B(new_n9146_), .ZN(new_n9147_));
  XOR2_X1    g08891(.A1(new_n9147_), .A2(\a[47] ), .Z(new_n9148_));
  INV_X1     g08892(.I(new_n9148_), .ZN(new_n9149_));
  NAND3_X1   g08893(.A1(new_n9144_), .A2(new_n9139_), .A3(new_n9149_), .ZN(new_n9150_));
  NOR2_X1    g08894(.A1(new_n9143_), .A2(new_n9140_), .ZN(new_n9151_));
  NOR2_X1    g08895(.A1(new_n9138_), .A2(new_n9118_), .ZN(new_n9152_));
  OAI21_X1   g08896(.A1(new_n9151_), .A2(new_n9152_), .B(new_n9148_), .ZN(new_n9153_));
  NAND2_X1   g08897(.A1(new_n9153_), .A2(new_n9150_), .ZN(new_n9154_));
  AOI21_X1   g08898(.A1(new_n8819_), .A2(new_n9113_), .B(new_n9154_), .ZN(new_n9155_));
  NAND2_X1   g08899(.A1(new_n9113_), .A2(new_n8819_), .ZN(new_n9156_));
  NOR3_X1    g08900(.A1(new_n9151_), .A2(new_n9152_), .A3(new_n9148_), .ZN(new_n9157_));
  AOI21_X1   g08901(.A1(new_n9144_), .A2(new_n9139_), .B(new_n9149_), .ZN(new_n9158_));
  NOR2_X1    g08902(.A1(new_n9157_), .A2(new_n9158_), .ZN(new_n9159_));
  NOR2_X1    g08903(.A1(new_n9159_), .A2(new_n9156_), .ZN(new_n9160_));
  AOI22_X1   g08904(.A1(new_n6569_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n6574_), .ZN(new_n9161_));
  OAI21_X1   g08905(.A1(new_n577_), .A2(new_n8565_), .B(new_n9161_), .ZN(new_n9162_));
  AOI21_X1   g08906(.A1(new_n1059_), .A2(new_n6579_), .B(new_n9162_), .ZN(new_n9163_));
  XOR2_X1    g08907(.A1(new_n9163_), .A2(new_n6567_), .Z(new_n9164_));
  NOR3_X1    g08908(.A1(new_n9155_), .A2(new_n9160_), .A3(new_n9164_), .ZN(new_n9165_));
  NAND2_X1   g08909(.A1(new_n9159_), .A2(new_n9156_), .ZN(new_n9166_));
  NAND3_X1   g08910(.A1(new_n9154_), .A2(new_n8819_), .A3(new_n9113_), .ZN(new_n9167_));
  INV_X1     g08911(.I(new_n9164_), .ZN(new_n9168_));
  AOI21_X1   g08912(.A1(new_n9167_), .A2(new_n9166_), .B(new_n9168_), .ZN(new_n9169_));
  NOR2_X1    g08913(.A1(new_n9165_), .A2(new_n9169_), .ZN(new_n9170_));
  AOI21_X1   g08914(.A1(new_n8837_), .A2(new_n9112_), .B(new_n9170_), .ZN(new_n9171_));
  AOI21_X1   g08915(.A1(new_n8829_), .A2(new_n8828_), .B(new_n8824_), .ZN(new_n9172_));
  NAND3_X1   g08916(.A1(new_n9167_), .A2(new_n9166_), .A3(new_n9168_), .ZN(new_n9173_));
  OAI21_X1   g08917(.A1(new_n9155_), .A2(new_n9160_), .B(new_n9164_), .ZN(new_n9174_));
  NAND2_X1   g08918(.A1(new_n9174_), .A2(new_n9173_), .ZN(new_n9175_));
  NOR3_X1    g08919(.A1(new_n9172_), .A2(new_n9175_), .A3(new_n8832_), .ZN(new_n9176_));
  OAI22_X1   g08920(.A1(new_n5852_), .A2(new_n1070_), .B1(new_n941_), .B2(new_n5857_), .ZN(new_n9177_));
  AOI21_X1   g08921(.A1(\b[11] ), .A2(new_n6115_), .B(new_n9177_), .ZN(new_n9178_));
  OAI21_X1   g08922(.A1(new_n1082_), .A2(new_n5861_), .B(new_n9178_), .ZN(new_n9179_));
  XOR2_X1    g08923(.A1(new_n9179_), .A2(\a[41] ), .Z(new_n9180_));
  INV_X1     g08924(.I(new_n9180_), .ZN(new_n9181_));
  OAI21_X1   g08925(.A1(new_n9171_), .A2(new_n9176_), .B(new_n9181_), .ZN(new_n9182_));
  OAI21_X1   g08926(.A1(new_n9172_), .A2(new_n8832_), .B(new_n9175_), .ZN(new_n9183_));
  NAND3_X1   g08927(.A1(new_n9170_), .A2(new_n9112_), .A3(new_n8837_), .ZN(new_n9184_));
  NAND3_X1   g08928(.A1(new_n9183_), .A2(new_n9184_), .A3(new_n9180_), .ZN(new_n9185_));
  NAND2_X1   g08929(.A1(new_n9182_), .A2(new_n9185_), .ZN(new_n9186_));
  AOI21_X1   g08930(.A1(new_n9111_), .A2(new_n8849_), .B(new_n9186_), .ZN(new_n9187_));
  AOI21_X1   g08931(.A1(new_n8844_), .A2(new_n8843_), .B(new_n8851_), .ZN(new_n9188_));
  AOI21_X1   g08932(.A1(new_n9183_), .A2(new_n9184_), .B(new_n9180_), .ZN(new_n9189_));
  NOR3_X1    g08933(.A1(new_n9171_), .A2(new_n9176_), .A3(new_n9181_), .ZN(new_n9190_));
  NOR2_X1    g08934(.A1(new_n9190_), .A2(new_n9189_), .ZN(new_n9191_));
  NOR3_X1    g08935(.A1(new_n9188_), .A2(new_n8853_), .A3(new_n9191_), .ZN(new_n9192_));
  NOR3_X1    g08936(.A1(new_n9192_), .A2(new_n9187_), .A3(new_n9110_), .ZN(new_n9193_));
  OAI21_X1   g08937(.A1(new_n9188_), .A2(new_n8853_), .B(new_n9191_), .ZN(new_n9194_));
  NAND3_X1   g08938(.A1(new_n9111_), .A2(new_n8849_), .A3(new_n9186_), .ZN(new_n9195_));
  AOI21_X1   g08939(.A1(new_n9194_), .A2(new_n9195_), .B(new_n9109_), .ZN(new_n9196_));
  NOR2_X1    g08940(.A1(new_n9193_), .A2(new_n9196_), .ZN(new_n9197_));
  NOR2_X1    g08941(.A1(new_n9105_), .A2(new_n9197_), .ZN(new_n9198_));
  NAND3_X1   g08942(.A1(new_n9194_), .A2(new_n9195_), .A3(new_n9109_), .ZN(new_n9199_));
  OAI21_X1   g08943(.A1(new_n9192_), .A2(new_n9187_), .B(new_n9110_), .ZN(new_n9200_));
  NAND2_X1   g08944(.A1(new_n9200_), .A2(new_n9199_), .ZN(new_n9201_));
  NOR3_X1    g08945(.A1(new_n9104_), .A2(new_n9201_), .A3(new_n8868_), .ZN(new_n9202_));
  AOI22_X1   g08946(.A1(new_n4918_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n4921_), .ZN(new_n9203_));
  OAI21_X1   g08947(.A1(new_n1432_), .A2(new_n6099_), .B(new_n9203_), .ZN(new_n9204_));
  AOI21_X1   g08948(.A1(new_n1695_), .A2(new_n4699_), .B(new_n9204_), .ZN(new_n9205_));
  XOR2_X1    g08949(.A1(new_n9205_), .A2(new_n4446_), .Z(new_n9206_));
  NOR3_X1    g08950(.A1(new_n9198_), .A2(new_n9202_), .A3(new_n9206_), .ZN(new_n9207_));
  OAI21_X1   g08951(.A1(new_n9104_), .A2(new_n8868_), .B(new_n9201_), .ZN(new_n9208_));
  INV_X1     g08952(.I(new_n9202_), .ZN(new_n9209_));
  INV_X1     g08953(.I(new_n9206_), .ZN(new_n9210_));
  AOI21_X1   g08954(.A1(new_n9209_), .A2(new_n9208_), .B(new_n9210_), .ZN(new_n9211_));
  NOR2_X1    g08955(.A1(new_n9211_), .A2(new_n9207_), .ZN(new_n9212_));
  NAND3_X1   g08956(.A1(new_n9212_), .A2(new_n9103_), .A3(new_n8887_), .ZN(new_n9213_));
  AOI21_X1   g08957(.A1(new_n8883_), .A2(new_n8880_), .B(new_n8889_), .ZN(new_n9214_));
  NAND3_X1   g08958(.A1(new_n9209_), .A2(new_n9208_), .A3(new_n9210_), .ZN(new_n9215_));
  OAI21_X1   g08959(.A1(new_n9198_), .A2(new_n9202_), .B(new_n9206_), .ZN(new_n9216_));
  NAND2_X1   g08960(.A1(new_n9215_), .A2(new_n9216_), .ZN(new_n9217_));
  OAI21_X1   g08961(.A1(new_n9214_), .A2(new_n8891_), .B(new_n9217_), .ZN(new_n9218_));
  AOI21_X1   g08962(.A1(new_n9218_), .A2(new_n9213_), .B(new_n9102_), .ZN(new_n9219_));
  INV_X1     g08963(.I(new_n9102_), .ZN(new_n9220_));
  NOR3_X1    g08964(.A1(new_n9214_), .A2(new_n9217_), .A3(new_n8891_), .ZN(new_n9221_));
  AOI21_X1   g08965(.A1(new_n9103_), .A2(new_n8887_), .B(new_n9212_), .ZN(new_n9222_));
  NOR3_X1    g08966(.A1(new_n9222_), .A2(new_n9221_), .A3(new_n9220_), .ZN(new_n9223_));
  NOR2_X1    g08967(.A1(new_n9223_), .A2(new_n9219_), .ZN(new_n9224_));
  OAI21_X1   g08968(.A1(new_n8893_), .A2(new_n8899_), .B(new_n8904_), .ZN(new_n9225_));
  NAND2_X1   g08969(.A1(new_n9225_), .A2(new_n9224_), .ZN(new_n9226_));
  OAI21_X1   g08970(.A1(new_n9222_), .A2(new_n9221_), .B(new_n9220_), .ZN(new_n9227_));
  NAND3_X1   g08971(.A1(new_n9218_), .A2(new_n9213_), .A3(new_n9102_), .ZN(new_n9228_));
  NAND2_X1   g08972(.A1(new_n9227_), .A2(new_n9228_), .ZN(new_n9229_));
  AOI21_X1   g08973(.A1(new_n8902_), .A2(new_n8903_), .B(new_n8900_), .ZN(new_n9230_));
  NAND2_X1   g08974(.A1(new_n9230_), .A2(new_n9229_), .ZN(new_n9231_));
  NAND3_X1   g08975(.A1(new_n9231_), .A2(new_n9226_), .A3(new_n9098_), .ZN(new_n9232_));
  INV_X1     g08976(.I(new_n9098_), .ZN(new_n9233_));
  NAND2_X1   g08977(.A1(new_n8903_), .A2(new_n8902_), .ZN(new_n9234_));
  AOI21_X1   g08978(.A1(new_n9234_), .A2(new_n8904_), .B(new_n9229_), .ZN(new_n9235_));
  NOR2_X1    g08979(.A1(new_n8899_), .A2(new_n8893_), .ZN(new_n9236_));
  NOR3_X1    g08980(.A1(new_n9236_), .A2(new_n9224_), .A3(new_n8900_), .ZN(new_n9237_));
  OAI21_X1   g08981(.A1(new_n9237_), .A2(new_n9235_), .B(new_n9233_), .ZN(new_n9238_));
  NAND2_X1   g08982(.A1(new_n9232_), .A2(new_n9238_), .ZN(new_n9239_));
  AOI21_X1   g08983(.A1(new_n9094_), .A2(new_n8917_), .B(new_n9239_), .ZN(new_n9240_));
  AOI21_X1   g08984(.A1(new_n8014_), .A2(new_n8019_), .B(new_n8020_), .ZN(new_n9241_));
  AOI21_X1   g08985(.A1(new_n9241_), .A2(new_n8357_), .B(new_n8356_), .ZN(new_n9242_));
  OAI21_X1   g08986(.A1(new_n9242_), .A2(new_n8664_), .B(new_n8659_), .ZN(new_n9243_));
  AOI21_X1   g08987(.A1(new_n9243_), .A2(new_n8910_), .B(new_n8906_), .ZN(new_n9244_));
  NOR3_X1    g08988(.A1(new_n9237_), .A2(new_n9235_), .A3(new_n9233_), .ZN(new_n9245_));
  AOI21_X1   g08989(.A1(new_n9231_), .A2(new_n9226_), .B(new_n9098_), .ZN(new_n9246_));
  NOR2_X1    g08990(.A1(new_n9246_), .A2(new_n9245_), .ZN(new_n9247_));
  NOR3_X1    g08991(.A1(new_n9247_), .A2(new_n9244_), .A3(new_n8913_), .ZN(new_n9248_));
  AOI22_X1   g08992(.A1(new_n2716_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n2719_), .ZN(new_n9249_));
  OAI21_X1   g08993(.A1(new_n3006_), .A2(new_n2924_), .B(new_n9249_), .ZN(new_n9250_));
  AOI21_X1   g08994(.A1(new_n3807_), .A2(new_n2722_), .B(new_n9250_), .ZN(new_n9251_));
  XOR2_X1    g08995(.A1(new_n9251_), .A2(new_n2714_), .Z(new_n9252_));
  INV_X1     g08996(.I(new_n9252_), .ZN(new_n9253_));
  NOR3_X1    g08997(.A1(new_n9240_), .A2(new_n9248_), .A3(new_n9253_), .ZN(new_n9254_));
  OAI21_X1   g08998(.A1(new_n9244_), .A2(new_n8913_), .B(new_n9247_), .ZN(new_n9255_));
  NAND3_X1   g08999(.A1(new_n9094_), .A2(new_n8917_), .A3(new_n9239_), .ZN(new_n9256_));
  AOI21_X1   g09000(.A1(new_n9256_), .A2(new_n9255_), .B(new_n9252_), .ZN(new_n9257_));
  NOR2_X1    g09001(.A1(new_n9257_), .A2(new_n9254_), .ZN(new_n9258_));
  OAI21_X1   g09002(.A1(new_n9093_), .A2(new_n9092_), .B(new_n9258_), .ZN(new_n9259_));
  AOI21_X1   g09003(.A1(new_n8684_), .A2(new_n8674_), .B(new_n8670_), .ZN(new_n9260_));
  OAI21_X1   g09004(.A1(new_n9260_), .A2(new_n8927_), .B(new_n8939_), .ZN(new_n9261_));
  NAND3_X1   g09005(.A1(new_n9256_), .A2(new_n9255_), .A3(new_n9252_), .ZN(new_n9262_));
  OAI21_X1   g09006(.A1(new_n9240_), .A2(new_n9248_), .B(new_n9253_), .ZN(new_n9263_));
  NAND2_X1   g09007(.A1(new_n9262_), .A2(new_n9263_), .ZN(new_n9264_));
  NAND3_X1   g09008(.A1(new_n9264_), .A2(new_n9261_), .A3(new_n8928_), .ZN(new_n9265_));
  NAND3_X1   g09009(.A1(new_n9259_), .A2(new_n9265_), .A3(new_n9091_), .ZN(new_n9266_));
  INV_X1     g09010(.I(new_n9091_), .ZN(new_n9267_));
  AOI21_X1   g09011(.A1(new_n8928_), .A2(new_n9261_), .B(new_n9264_), .ZN(new_n9268_));
  NOR3_X1    g09012(.A1(new_n9093_), .A2(new_n9258_), .A3(new_n9092_), .ZN(new_n9269_));
  OAI21_X1   g09013(.A1(new_n9268_), .A2(new_n9269_), .B(new_n9267_), .ZN(new_n9270_));
  NAND2_X1   g09014(.A1(new_n9270_), .A2(new_n9266_), .ZN(new_n9271_));
  NAND3_X1   g09015(.A1(new_n9087_), .A2(new_n8937_), .A3(new_n9271_), .ZN(new_n9272_));
  AOI21_X1   g09016(.A1(new_n8945_), .A2(new_n8934_), .B(new_n8942_), .ZN(new_n9273_));
  NOR3_X1    g09017(.A1(new_n9268_), .A2(new_n9269_), .A3(new_n9267_), .ZN(new_n9274_));
  AOI21_X1   g09018(.A1(new_n9259_), .A2(new_n9265_), .B(new_n9091_), .ZN(new_n9275_));
  NOR2_X1    g09019(.A1(new_n9274_), .A2(new_n9275_), .ZN(new_n9276_));
  OAI21_X1   g09020(.A1(new_n9273_), .A2(new_n8946_), .B(new_n9276_), .ZN(new_n9277_));
  NAND3_X1   g09021(.A1(new_n9272_), .A2(new_n9277_), .A3(new_n9086_), .ZN(new_n9278_));
  INV_X1     g09022(.I(new_n9086_), .ZN(new_n9279_));
  NOR3_X1    g09023(.A1(new_n9273_), .A2(new_n9276_), .A3(new_n8946_), .ZN(new_n9280_));
  AOI21_X1   g09024(.A1(new_n9087_), .A2(new_n8937_), .B(new_n9271_), .ZN(new_n9281_));
  OAI21_X1   g09025(.A1(new_n9281_), .A2(new_n9280_), .B(new_n9279_), .ZN(new_n9282_));
  NAND2_X1   g09026(.A1(new_n9282_), .A2(new_n9278_), .ZN(new_n9283_));
  NOR3_X1    g09027(.A1(new_n9082_), .A2(new_n9283_), .A3(new_n9081_), .ZN(new_n9284_));
  OAI21_X1   g09028(.A1(new_n8053_), .A2(new_n8059_), .B(new_n8063_), .ZN(new_n9285_));
  OAI21_X1   g09029(.A1(new_n9285_), .A2(new_n8402_), .B(new_n8401_), .ZN(new_n9286_));
  AOI21_X1   g09030(.A1(new_n9286_), .A2(new_n8697_), .B(new_n8693_), .ZN(new_n9287_));
  OAI21_X1   g09031(.A1(new_n9287_), .A2(new_n8957_), .B(new_n8949_), .ZN(new_n9288_));
  NOR3_X1    g09032(.A1(new_n9281_), .A2(new_n9279_), .A3(new_n9280_), .ZN(new_n9289_));
  AOI21_X1   g09033(.A1(new_n9272_), .A2(new_n9277_), .B(new_n9086_), .ZN(new_n9290_));
  NOR2_X1    g09034(.A1(new_n9289_), .A2(new_n9290_), .ZN(new_n9291_));
  AOI21_X1   g09035(.A1(new_n9288_), .A2(new_n8958_), .B(new_n9291_), .ZN(new_n9292_));
  OAI21_X1   g09036(.A1(new_n9292_), .A2(new_n9284_), .B(new_n9080_), .ZN(new_n9293_));
  INV_X1     g09037(.I(new_n9080_), .ZN(new_n9294_));
  NAND3_X1   g09038(.A1(new_n9288_), .A2(new_n9291_), .A3(new_n8958_), .ZN(new_n9295_));
  OAI21_X1   g09039(.A1(new_n9082_), .A2(new_n9081_), .B(new_n9283_), .ZN(new_n9296_));
  NAND3_X1   g09040(.A1(new_n9296_), .A2(new_n9295_), .A3(new_n9294_), .ZN(new_n9297_));
  NAND2_X1   g09041(.A1(new_n9293_), .A2(new_n9297_), .ZN(new_n9298_));
  NAND3_X1   g09042(.A1(new_n9076_), .A2(new_n9072_), .A3(new_n9298_), .ZN(new_n9299_));
  AOI21_X1   g09043(.A1(new_n8065_), .A2(new_n8076_), .B(new_n8072_), .ZN(new_n9300_));
  AOI21_X1   g09044(.A1(new_n9300_), .A2(new_n8414_), .B(new_n8413_), .ZN(new_n9301_));
  OAI21_X1   g09045(.A1(new_n9301_), .A2(new_n8712_), .B(new_n8711_), .ZN(new_n9302_));
  AOI21_X1   g09046(.A1(new_n9302_), .A2(new_n8966_), .B(new_n8962_), .ZN(new_n9303_));
  AOI21_X1   g09047(.A1(new_n9296_), .A2(new_n9295_), .B(new_n9294_), .ZN(new_n9304_));
  NOR3_X1    g09048(.A1(new_n9292_), .A2(new_n9284_), .A3(new_n9080_), .ZN(new_n9305_));
  NOR2_X1    g09049(.A1(new_n9304_), .A2(new_n9305_), .ZN(new_n9306_));
  OAI21_X1   g09050(.A1(new_n9303_), .A2(new_n8969_), .B(new_n9306_), .ZN(new_n9307_));
  NAND3_X1   g09051(.A1(new_n9307_), .A2(new_n9299_), .A3(new_n9071_), .ZN(new_n9308_));
  INV_X1     g09052(.I(new_n9071_), .ZN(new_n9309_));
  NOR3_X1    g09053(.A1(new_n9303_), .A2(new_n8969_), .A3(new_n9306_), .ZN(new_n9310_));
  AOI21_X1   g09054(.A1(new_n9076_), .A2(new_n9072_), .B(new_n9298_), .ZN(new_n9311_));
  OAI21_X1   g09055(.A1(new_n9310_), .A2(new_n9311_), .B(new_n9309_), .ZN(new_n9312_));
  NAND2_X1   g09056(.A1(new_n9312_), .A2(new_n9308_), .ZN(new_n9313_));
  NOR3_X1    g09057(.A1(new_n9067_), .A2(new_n8985_), .A3(new_n9313_), .ZN(new_n9314_));
  AOI21_X1   g09058(.A1(new_n8973_), .A2(new_n8978_), .B(new_n8985_), .ZN(new_n9315_));
  NOR3_X1    g09059(.A1(new_n9310_), .A2(new_n9311_), .A3(new_n9309_), .ZN(new_n9316_));
  AOI21_X1   g09060(.A1(new_n9307_), .A2(new_n9299_), .B(new_n9071_), .ZN(new_n9317_));
  NOR2_X1    g09061(.A1(new_n9316_), .A2(new_n9317_), .ZN(new_n9318_));
  NOR2_X1    g09062(.A1(new_n9315_), .A2(new_n9318_), .ZN(new_n9319_));
  OAI21_X1   g09063(.A1(new_n9319_), .A2(new_n9314_), .B(new_n9063_), .ZN(new_n9320_));
  INV_X1     g09064(.I(new_n9063_), .ZN(new_n9321_));
  OAI21_X1   g09065(.A1(new_n8080_), .A2(new_n8086_), .B(new_n8093_), .ZN(new_n9322_));
  OAI21_X1   g09066(.A1(new_n9322_), .A2(new_n8435_), .B(new_n8434_), .ZN(new_n9323_));
  AOI21_X1   g09067(.A1(new_n9323_), .A2(new_n8721_), .B(new_n8720_), .ZN(new_n9324_));
  OAI21_X1   g09068(.A1(new_n9324_), .A2(new_n8979_), .B(new_n8973_), .ZN(new_n9325_));
  NAND3_X1   g09069(.A1(new_n9325_), .A2(new_n9318_), .A3(new_n8980_), .ZN(new_n9326_));
  OAI21_X1   g09070(.A1(new_n8983_), .A2(new_n8984_), .B(new_n8980_), .ZN(new_n9327_));
  NAND2_X1   g09071(.A1(new_n9327_), .A2(new_n9313_), .ZN(new_n9328_));
  NAND3_X1   g09072(.A1(new_n9328_), .A2(new_n9321_), .A3(new_n9326_), .ZN(new_n9329_));
  NAND2_X1   g09073(.A1(new_n9320_), .A2(new_n9329_), .ZN(new_n9330_));
  NOR3_X1    g09074(.A1(new_n9330_), .A2(new_n9059_), .A3(new_n8995_), .ZN(new_n9331_));
  AOI21_X1   g09075(.A1(new_n8997_), .A2(new_n8998_), .B(new_n8995_), .ZN(new_n9332_));
  AOI21_X1   g09076(.A1(new_n9328_), .A2(new_n9326_), .B(new_n9321_), .ZN(new_n9333_));
  NOR3_X1    g09077(.A1(new_n9319_), .A2(new_n9314_), .A3(new_n9063_), .ZN(new_n9334_));
  NOR2_X1    g09078(.A1(new_n9333_), .A2(new_n9334_), .ZN(new_n9335_));
  NOR2_X1    g09079(.A1(new_n9332_), .A2(new_n9335_), .ZN(new_n9336_));
  INV_X1     g09080(.I(new_n7627_), .ZN(new_n9337_));
  AOI22_X1   g09081(.A1(new_n518_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n636_), .ZN(new_n9338_));
  OAI21_X1   g09082(.A1(new_n7074_), .A2(new_n917_), .B(new_n9338_), .ZN(new_n9339_));
  AOI21_X1   g09083(.A1(new_n9337_), .A2(new_n618_), .B(new_n9339_), .ZN(new_n9340_));
  XOR2_X1    g09084(.A1(new_n9340_), .A2(new_n488_), .Z(new_n9341_));
  INV_X1     g09085(.I(new_n9341_), .ZN(new_n9342_));
  OAI21_X1   g09086(.A1(new_n9336_), .A2(new_n9331_), .B(new_n9342_), .ZN(new_n9343_));
  NAND2_X1   g09087(.A1(new_n9332_), .A2(new_n9335_), .ZN(new_n9344_));
  OAI21_X1   g09088(.A1(new_n8995_), .A2(new_n9059_), .B(new_n9330_), .ZN(new_n9345_));
  NAND3_X1   g09089(.A1(new_n9344_), .A2(new_n9345_), .A3(new_n9341_), .ZN(new_n9346_));
  NAND2_X1   g09090(.A1(new_n9343_), .A2(new_n9346_), .ZN(new_n9347_));
  AOI21_X1   g09091(.A1(new_n7896_), .A2(new_n7883_), .B(new_n8117_), .ZN(new_n9348_));
  OAI21_X1   g09092(.A1(new_n8108_), .A2(new_n9348_), .B(new_n8118_), .ZN(new_n9349_));
  OAI21_X1   g09093(.A1(new_n9349_), .A2(new_n8471_), .B(new_n8470_), .ZN(new_n9350_));
  AOI21_X1   g09094(.A1(new_n9350_), .A2(new_n8748_), .B(new_n8746_), .ZN(new_n9351_));
  OAI21_X1   g09095(.A1(new_n9351_), .A2(new_n9008_), .B(new_n9001_), .ZN(new_n9352_));
  AOI21_X1   g09096(.A1(new_n9009_), .A2(new_n9352_), .B(new_n9347_), .ZN(new_n9353_));
  AOI21_X1   g09097(.A1(new_n9344_), .A2(new_n9345_), .B(new_n9341_), .ZN(new_n9354_));
  NOR3_X1    g09098(.A1(new_n9336_), .A2(new_n9331_), .A3(new_n9342_), .ZN(new_n9355_));
  NOR2_X1    g09099(.A1(new_n9354_), .A2(new_n9355_), .ZN(new_n9356_));
  OAI21_X1   g09100(.A1(new_n8515_), .A2(new_n8744_), .B(new_n8739_), .ZN(new_n9357_));
  AOI21_X1   g09101(.A1(new_n9357_), .A2(new_n9006_), .B(new_n9011_), .ZN(new_n9358_));
  NOR3_X1    g09102(.A1(new_n9356_), .A2(new_n9358_), .A3(new_n9013_), .ZN(new_n9359_));
  NOR3_X1    g09103(.A1(new_n9353_), .A2(new_n9359_), .A3(new_n9055_), .ZN(new_n9360_));
  OAI21_X1   g09104(.A1(new_n9013_), .A2(new_n9358_), .B(new_n9356_), .ZN(new_n9361_));
  NAND3_X1   g09105(.A1(new_n9347_), .A2(new_n9352_), .A3(new_n9009_), .ZN(new_n9362_));
  AOI21_X1   g09106(.A1(new_n9361_), .A2(new_n9362_), .B(new_n9054_), .ZN(new_n9363_));
  OAI22_X1   g09107(.A1(new_n9049_), .A2(new_n9015_), .B1(new_n9360_), .B2(new_n9363_), .ZN(new_n9364_));
  NOR2_X1    g09108(.A1(new_n9049_), .A2(new_n9015_), .ZN(new_n9365_));
  NOR2_X1    g09109(.A1(new_n9360_), .A2(new_n9363_), .ZN(new_n9366_));
  NAND2_X1   g09110(.A1(new_n9365_), .A2(new_n9366_), .ZN(new_n9367_));
  NAND2_X1   g09111(.A1(new_n9367_), .A2(new_n9364_), .ZN(new_n9368_));
  NOR2_X1    g09112(.A1(new_n9368_), .A2(new_n9046_), .ZN(new_n9369_));
  INV_X1     g09113(.I(new_n9369_), .ZN(new_n9370_));
  NAND2_X1   g09114(.A1(new_n9368_), .A2(new_n9046_), .ZN(new_n9371_));
  NAND2_X1   g09115(.A1(new_n9370_), .A2(new_n9371_), .ZN(new_n9372_));
  XOR2_X1    g09116(.A1(new_n9372_), .A2(new_n9031_), .Z(\f[52] ));
  OAI21_X1   g09117(.A1(new_n8773_), .A2(new_n9024_), .B(new_n9023_), .ZN(new_n9374_));
  AOI21_X1   g09118(.A1(new_n9374_), .A2(new_n9371_), .B(new_n9369_), .ZN(new_n9375_));
  INV_X1     g09119(.I(\b[53] ), .ZN(new_n9376_));
  OAI22_X1   g09120(.A1(new_n277_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n262_), .ZN(new_n9377_));
  AOI21_X1   g09121(.A1(\b[51] ), .A2(new_n283_), .B(new_n9377_), .ZN(new_n9378_));
  AOI21_X1   g09122(.A1(new_n9039_), .A2(\b[52] ), .B(new_n8776_), .ZN(new_n9379_));
  NOR2_X1    g09123(.A1(new_n9039_), .A2(\b[52] ), .ZN(new_n9380_));
  NOR2_X1    g09124(.A1(new_n9379_), .A2(new_n9380_), .ZN(new_n9381_));
  NAND3_X1   g09125(.A1(new_n9037_), .A2(new_n9038_), .A3(new_n9376_), .ZN(new_n9382_));
  NAND2_X1   g09126(.A1(new_n9039_), .A2(\b[53] ), .ZN(new_n9383_));
  NAND2_X1   g09127(.A1(new_n9383_), .A2(new_n9382_), .ZN(new_n9384_));
  XOR2_X1    g09128(.A1(new_n9381_), .A2(new_n9384_), .Z(new_n9385_));
  OAI21_X1   g09129(.A1(new_n9385_), .A2(new_n279_), .B(new_n9378_), .ZN(new_n9386_));
  XOR2_X1    g09130(.A1(new_n9386_), .A2(\a[2] ), .Z(new_n9387_));
  INV_X1     g09131(.I(new_n9387_), .ZN(new_n9388_));
  NOR3_X1    g09132(.A1(new_n9358_), .A2(new_n9013_), .A3(new_n9354_), .ZN(new_n9389_));
  AOI22_X1   g09133(.A1(new_n518_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n636_), .ZN(new_n9390_));
  OAI21_X1   g09134(.A1(new_n7096_), .A2(new_n917_), .B(new_n9390_), .ZN(new_n9391_));
  INV_X1     g09135(.I(new_n9391_), .ZN(new_n9392_));
  NAND2_X1   g09136(.A1(new_n7649_), .A2(new_n618_), .ZN(new_n9393_));
  AOI21_X1   g09137(.A1(new_n9393_), .A2(new_n9392_), .B(new_n488_), .ZN(new_n9394_));
  NAND3_X1   g09138(.A1(new_n9393_), .A2(new_n488_), .A3(new_n9392_), .ZN(new_n9395_));
  INV_X1     g09139(.I(new_n9395_), .ZN(new_n9396_));
  NOR2_X1    g09140(.A1(new_n9396_), .A2(new_n9394_), .ZN(new_n9397_));
  OAI21_X1   g09141(.A1(new_n8104_), .A2(new_n8105_), .B(new_n8102_), .ZN(new_n9398_));
  OAI21_X1   g09142(.A1(new_n9398_), .A2(new_n8454_), .B(new_n8453_), .ZN(new_n9399_));
  AOI21_X1   g09143(.A1(new_n9399_), .A2(new_n8733_), .B(new_n8732_), .ZN(new_n9400_));
  OAI21_X1   g09144(.A1(new_n9400_), .A2(new_n8993_), .B(new_n8997_), .ZN(new_n9401_));
  AOI21_X1   g09145(.A1(new_n9401_), .A2(new_n8999_), .B(new_n9334_), .ZN(new_n9402_));
  OAI22_X1   g09146(.A1(new_n713_), .A2(new_n7074_), .B1(new_n6775_), .B2(new_n717_), .ZN(new_n9403_));
  AOI21_X1   g09147(.A1(\b[42] ), .A2(new_n1126_), .B(new_n9403_), .ZN(new_n9404_));
  OAI21_X1   g09148(.A1(new_n7081_), .A2(new_n986_), .B(new_n9404_), .ZN(new_n9405_));
  XOR2_X1    g09149(.A1(new_n9405_), .A2(new_n722_), .Z(new_n9406_));
  AOI22_X1   g09150(.A1(new_n1006_), .A2(\b[41] ), .B1(\b[40] ), .B2(new_n1009_), .ZN(new_n9407_));
  OAI21_X1   g09151(.A1(new_n5761_), .A2(new_n1481_), .B(new_n9407_), .ZN(new_n9408_));
  INV_X1     g09152(.I(new_n9408_), .ZN(new_n9409_));
  NAND3_X1   g09153(.A1(new_n6298_), .A2(new_n6295_), .A3(new_n1013_), .ZN(new_n9410_));
  NAND2_X1   g09154(.A1(new_n9410_), .A2(new_n9409_), .ZN(new_n9411_));
  XOR2_X1    g09155(.A1(new_n9411_), .A2(new_n1002_), .Z(new_n9412_));
  OAI22_X1   g09156(.A1(new_n1592_), .A2(new_n5341_), .B1(new_n5312_), .B2(new_n1505_), .ZN(new_n9413_));
  AOI21_X1   g09157(.A1(\b[36] ), .A2(new_n1584_), .B(new_n9413_), .ZN(new_n9414_));
  OAI21_X1   g09158(.A1(new_n5352_), .A2(new_n1732_), .B(new_n9414_), .ZN(new_n9415_));
  XOR2_X1    g09159(.A1(new_n9415_), .A2(\a[17] ), .Z(new_n9416_));
  INV_X1     g09160(.I(new_n9416_), .ZN(new_n9417_));
  OAI22_X1   g09161(.A1(new_n1751_), .A2(new_n4666_), .B1(new_n4639_), .B2(new_n1754_), .ZN(new_n9418_));
  AOI21_X1   g09162(.A1(\b[33] ), .A2(new_n1939_), .B(new_n9418_), .ZN(new_n9419_));
  OAI21_X1   g09163(.A1(new_n4676_), .A2(new_n1757_), .B(new_n9419_), .ZN(new_n9420_));
  XOR2_X1    g09164(.A1(new_n9420_), .A2(\a[20] ), .Z(new_n9421_));
  INV_X1     g09165(.I(new_n9421_), .ZN(new_n9422_));
  AOI21_X1   g09166(.A1(new_n9259_), .A2(new_n9265_), .B(new_n9267_), .ZN(new_n9423_));
  INV_X1     g09167(.I(new_n9423_), .ZN(new_n9424_));
  AOI22_X1   g09168(.A1(new_n2202_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n2205_), .ZN(new_n9425_));
  OAI21_X1   g09169(.A1(new_n3624_), .A2(new_n2370_), .B(new_n9425_), .ZN(new_n9426_));
  AOI21_X1   g09170(.A1(new_n4030_), .A2(new_n2208_), .B(new_n9426_), .ZN(new_n9427_));
  XOR2_X1    g09171(.A1(new_n9427_), .A2(new_n2200_), .Z(new_n9428_));
  AOI21_X1   g09172(.A1(new_n9261_), .A2(new_n8928_), .B(new_n9254_), .ZN(new_n9429_));
  NOR2_X1    g09173(.A1(new_n9429_), .A2(new_n9257_), .ZN(new_n9430_));
  AOI22_X1   g09174(.A1(new_n2716_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n2719_), .ZN(new_n9431_));
  OAI21_X1   g09175(.A1(new_n3158_), .A2(new_n2924_), .B(new_n9431_), .ZN(new_n9432_));
  AOI21_X1   g09176(.A1(new_n4188_), .A2(new_n2722_), .B(new_n9432_), .ZN(new_n9433_));
  XOR2_X1    g09177(.A1(new_n9433_), .A2(new_n2714_), .Z(new_n9434_));
  INV_X1     g09178(.I(new_n9434_), .ZN(new_n9435_));
  AOI21_X1   g09179(.A1(new_n9231_), .A2(new_n9226_), .B(new_n9233_), .ZN(new_n9436_));
  INV_X1     g09180(.I(new_n9436_), .ZN(new_n9437_));
  OAI21_X1   g09181(.A1(new_n9236_), .A2(new_n8900_), .B(new_n9228_), .ZN(new_n9438_));
  AOI22_X1   g09182(.A1(new_n3864_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n3869_), .ZN(new_n9439_));
  OAI21_X1   g09183(.A1(new_n2027_), .A2(new_n5410_), .B(new_n9439_), .ZN(new_n9440_));
  AOI21_X1   g09184(.A1(new_n2470_), .A2(new_n3872_), .B(new_n9440_), .ZN(new_n9441_));
  XOR2_X1    g09185(.A1(new_n9441_), .A2(new_n3876_), .Z(new_n9442_));
  AOI21_X1   g09186(.A1(new_n9103_), .A2(new_n8887_), .B(new_n9211_), .ZN(new_n9443_));
  AOI21_X1   g09187(.A1(new_n9194_), .A2(new_n9195_), .B(new_n9110_), .ZN(new_n9444_));
  NOR3_X1    g09188(.A1(new_n9197_), .A2(new_n9104_), .A3(new_n8868_), .ZN(new_n9445_));
  OAI22_X1   g09189(.A1(new_n1432_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n1296_), .ZN(new_n9446_));
  AOI21_X1   g09190(.A1(\b[15] ), .A2(new_n5420_), .B(new_n9446_), .ZN(new_n9447_));
  OAI21_X1   g09191(.A1(new_n1444_), .A2(new_n6124_), .B(new_n9447_), .ZN(new_n9448_));
  XOR2_X1    g09192(.A1(new_n9448_), .A2(\a[38] ), .Z(new_n9449_));
  NAND3_X1   g09193(.A1(new_n9111_), .A2(new_n8849_), .A3(new_n9182_), .ZN(new_n9450_));
  AOI22_X1   g09194(.A1(new_n6108_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n6111_), .ZN(new_n9451_));
  OAI21_X1   g09195(.A1(new_n941_), .A2(new_n7708_), .B(new_n9451_), .ZN(new_n9452_));
  AOI21_X1   g09196(.A1(new_n1449_), .A2(new_n6105_), .B(new_n9452_), .ZN(new_n9453_));
  XOR2_X1    g09197(.A1(new_n9453_), .A2(\a[41] ), .Z(new_n9454_));
  INV_X1     g09198(.I(new_n9454_), .ZN(new_n9455_));
  AOI21_X1   g09199(.A1(new_n9112_), .A2(new_n8837_), .B(new_n9169_), .ZN(new_n9456_));
  AOI21_X1   g09200(.A1(new_n9113_), .A2(new_n8819_), .B(new_n9158_), .ZN(new_n9457_));
  NOR2_X1    g09201(.A1(new_n9457_), .A2(new_n9157_), .ZN(new_n9458_));
  NAND2_X1   g09202(.A1(new_n9141_), .A2(new_n9118_), .ZN(new_n9459_));
  INV_X1     g09203(.I(new_n8252_), .ZN(new_n9460_));
  INV_X1     g09204(.I(new_n8241_), .ZN(new_n9461_));
  INV_X1     g09205(.I(new_n8246_), .ZN(new_n9462_));
  OAI22_X1   g09206(.A1(new_n9461_), .A2(new_n377_), .B1(new_n339_), .B2(new_n9462_), .ZN(new_n9463_));
  AOI21_X1   g09207(.A1(\b[3] ), .A2(new_n8575_), .B(new_n9463_), .ZN(new_n9464_));
  OAI21_X1   g09208(.A1(new_n566_), .A2(new_n9460_), .B(new_n9464_), .ZN(new_n9465_));
  XOR2_X1    g09209(.A1(new_n9465_), .A2(\a[50] ), .Z(new_n9466_));
  AOI22_X1   g09210(.A1(new_n9125_), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n9123_), .ZN(new_n9467_));
  NOR4_X1    g09211(.A1(new_n8248_), .A2(new_n9119_), .A3(new_n9121_), .A4(\a[53] ), .ZN(new_n9468_));
  NOR4_X1    g09212(.A1(new_n9133_), .A2(\a[50] ), .A3(\a[51] ), .A4(\a[52] ), .ZN(new_n9469_));
  NOR2_X1    g09213(.A1(new_n9468_), .A2(new_n9469_), .ZN(new_n9470_));
  INV_X1     g09214(.I(new_n9470_), .ZN(new_n9471_));
  NAND2_X1   g09215(.A1(new_n9471_), .A2(\b[0] ), .ZN(new_n9472_));
  NAND2_X1   g09216(.A1(new_n9129_), .A2(new_n554_), .ZN(new_n9473_));
  NAND3_X1   g09217(.A1(new_n9473_), .A2(new_n9467_), .A3(new_n9472_), .ZN(new_n9474_));
  NAND2_X1   g09218(.A1(new_n9474_), .A2(\a[53] ), .ZN(new_n9475_));
  NAND4_X1   g09219(.A1(new_n9473_), .A2(new_n9467_), .A3(new_n9472_), .A4(new_n9133_), .ZN(new_n9476_));
  NOR3_X1    g09220(.A1(new_n9131_), .A2(new_n9133_), .A3(new_n8804_), .ZN(new_n9477_));
  NAND3_X1   g09221(.A1(new_n9475_), .A2(new_n9477_), .A3(new_n9476_), .ZN(new_n9478_));
  INV_X1     g09222(.I(new_n9478_), .ZN(new_n9479_));
  AOI21_X1   g09223(.A1(new_n9476_), .A2(new_n9475_), .B(new_n9477_), .ZN(new_n9480_));
  NOR2_X1    g09224(.A1(new_n9479_), .A2(new_n9480_), .ZN(new_n9481_));
  NOR2_X1    g09225(.A1(new_n9466_), .A2(new_n9481_), .ZN(new_n9482_));
  AND2_X2    g09226(.A1(new_n9466_), .A2(new_n9481_), .Z(new_n9483_));
  NOR2_X1    g09227(.A1(new_n9483_), .A2(new_n9482_), .ZN(new_n9484_));
  NAND3_X1   g09228(.A1(new_n9484_), .A2(new_n9142_), .A3(new_n9459_), .ZN(new_n9485_));
  INV_X1     g09229(.I(new_n9485_), .ZN(new_n9486_));
  AOI21_X1   g09230(.A1(new_n9142_), .A2(new_n9459_), .B(new_n9484_), .ZN(new_n9487_));
  INV_X1     g09231(.I(new_n7719_), .ZN(new_n9488_));
  AOI22_X1   g09232(.A1(new_n7403_), .A2(\b[8] ), .B1(\b[7] ), .B2(new_n7408_), .ZN(new_n9489_));
  OAI21_X1   g09233(.A1(new_n438_), .A2(new_n9488_), .B(new_n9489_), .ZN(new_n9490_));
  AOI21_X1   g09234(.A1(new_n799_), .A2(new_n7414_), .B(new_n9490_), .ZN(new_n9491_));
  XOR2_X1    g09235(.A1(new_n9491_), .A2(new_n7410_), .Z(new_n9492_));
  INV_X1     g09236(.I(new_n9492_), .ZN(new_n9493_));
  OAI21_X1   g09237(.A1(new_n9486_), .A2(new_n9487_), .B(new_n9493_), .ZN(new_n9494_));
  INV_X1     g09238(.I(new_n9487_), .ZN(new_n9495_));
  NAND3_X1   g09239(.A1(new_n9495_), .A2(new_n9485_), .A3(new_n9492_), .ZN(new_n9496_));
  NAND2_X1   g09240(.A1(new_n9496_), .A2(new_n9494_), .ZN(new_n9497_));
  NOR2_X1    g09241(.A1(new_n9458_), .A2(new_n9497_), .ZN(new_n9498_));
  AOI21_X1   g09242(.A1(new_n9495_), .A2(new_n9485_), .B(new_n9492_), .ZN(new_n9499_));
  NOR3_X1    g09243(.A1(new_n9486_), .A2(new_n9487_), .A3(new_n9493_), .ZN(new_n9500_));
  NOR2_X1    g09244(.A1(new_n9499_), .A2(new_n9500_), .ZN(new_n9501_));
  NOR3_X1    g09245(.A1(new_n9501_), .A2(new_n9457_), .A3(new_n9157_), .ZN(new_n9502_));
  OAI22_X1   g09246(.A1(new_n7730_), .A2(new_n852_), .B1(new_n776_), .B2(new_n7731_), .ZN(new_n9503_));
  AOI21_X1   g09247(.A1(\b[9] ), .A2(new_n6887_), .B(new_n9503_), .ZN(new_n9504_));
  OAI21_X1   g09248(.A1(new_n859_), .A2(new_n7728_), .B(new_n9504_), .ZN(new_n9505_));
  XOR2_X1    g09249(.A1(new_n9505_), .A2(\a[44] ), .Z(new_n9506_));
  OAI21_X1   g09250(.A1(new_n9498_), .A2(new_n9502_), .B(new_n9506_), .ZN(new_n9507_));
  NAND2_X1   g09251(.A1(new_n9156_), .A2(new_n9153_), .ZN(new_n9508_));
  NAND2_X1   g09252(.A1(new_n9508_), .A2(new_n9150_), .ZN(new_n9509_));
  NAND2_X1   g09253(.A1(new_n9509_), .A2(new_n9501_), .ZN(new_n9510_));
  NAND2_X1   g09254(.A1(new_n9458_), .A2(new_n9497_), .ZN(new_n9511_));
  INV_X1     g09255(.I(new_n9506_), .ZN(new_n9512_));
  NAND3_X1   g09256(.A1(new_n9510_), .A2(new_n9511_), .A3(new_n9512_), .ZN(new_n9513_));
  NAND2_X1   g09257(.A1(new_n9513_), .A2(new_n9507_), .ZN(new_n9514_));
  NOR3_X1    g09258(.A1(new_n9514_), .A2(new_n9456_), .A3(new_n9165_), .ZN(new_n9515_));
  OAI21_X1   g09259(.A1(new_n9172_), .A2(new_n8832_), .B(new_n9174_), .ZN(new_n9516_));
  AOI21_X1   g09260(.A1(new_n9510_), .A2(new_n9511_), .B(new_n9512_), .ZN(new_n9517_));
  NOR3_X1    g09261(.A1(new_n9498_), .A2(new_n9502_), .A3(new_n9506_), .ZN(new_n9518_));
  NOR2_X1    g09262(.A1(new_n9517_), .A2(new_n9518_), .ZN(new_n9519_));
  AOI21_X1   g09263(.A1(new_n9516_), .A2(new_n9173_), .B(new_n9519_), .ZN(new_n9520_));
  OAI21_X1   g09264(.A1(new_n9520_), .A2(new_n9515_), .B(new_n9455_), .ZN(new_n9521_));
  NAND3_X1   g09265(.A1(new_n9516_), .A2(new_n9519_), .A3(new_n9173_), .ZN(new_n9522_));
  OAI21_X1   g09266(.A1(new_n9456_), .A2(new_n9165_), .B(new_n9514_), .ZN(new_n9523_));
  NAND3_X1   g09267(.A1(new_n9523_), .A2(new_n9522_), .A3(new_n9454_), .ZN(new_n9524_));
  NAND2_X1   g09268(.A1(new_n9521_), .A2(new_n9524_), .ZN(new_n9525_));
  AOI21_X1   g09269(.A1(new_n9450_), .A2(new_n9185_), .B(new_n9525_), .ZN(new_n9526_));
  NOR3_X1    g09270(.A1(new_n9188_), .A2(new_n8853_), .A3(new_n9189_), .ZN(new_n9527_));
  AOI21_X1   g09271(.A1(new_n9523_), .A2(new_n9522_), .B(new_n9454_), .ZN(new_n9528_));
  NOR3_X1    g09272(.A1(new_n9520_), .A2(new_n9455_), .A3(new_n9515_), .ZN(new_n9529_));
  NOR2_X1    g09273(.A1(new_n9529_), .A2(new_n9528_), .ZN(new_n9530_));
  NOR3_X1    g09274(.A1(new_n9527_), .A2(new_n9530_), .A3(new_n9190_), .ZN(new_n9531_));
  NOR3_X1    g09275(.A1(new_n9531_), .A2(new_n9526_), .A3(new_n9449_), .ZN(new_n9532_));
  INV_X1     g09276(.I(new_n9449_), .ZN(new_n9533_));
  OAI21_X1   g09277(.A1(new_n9527_), .A2(new_n9190_), .B(new_n9530_), .ZN(new_n9534_));
  NAND3_X1   g09278(.A1(new_n9450_), .A2(new_n9525_), .A3(new_n9185_), .ZN(new_n9535_));
  AOI21_X1   g09279(.A1(new_n9534_), .A2(new_n9535_), .B(new_n9533_), .ZN(new_n9536_));
  NOR2_X1    g09280(.A1(new_n9532_), .A2(new_n9536_), .ZN(new_n9537_));
  NOR3_X1    g09281(.A1(new_n9445_), .A2(new_n9537_), .A3(new_n9444_), .ZN(new_n9538_));
  INV_X1     g09282(.I(new_n9444_), .ZN(new_n9539_));
  OAI21_X1   g09283(.A1(new_n8863_), .A2(new_n8860_), .B(new_n8872_), .ZN(new_n9540_));
  NAND3_X1   g09284(.A1(new_n9540_), .A2(new_n9201_), .A3(new_n8874_), .ZN(new_n9541_));
  NAND3_X1   g09285(.A1(new_n9534_), .A2(new_n9535_), .A3(new_n9533_), .ZN(new_n9542_));
  OAI21_X1   g09286(.A1(new_n9531_), .A2(new_n9526_), .B(new_n9449_), .ZN(new_n9543_));
  NAND2_X1   g09287(.A1(new_n9543_), .A2(new_n9542_), .ZN(new_n9544_));
  AOI21_X1   g09288(.A1(new_n9541_), .A2(new_n9539_), .B(new_n9544_), .ZN(new_n9545_));
  AOI22_X1   g09289(.A1(new_n4918_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n4921_), .ZN(new_n9546_));
  OAI21_X1   g09290(.A1(new_n1553_), .A2(new_n6099_), .B(new_n9546_), .ZN(new_n9547_));
  AOI21_X1   g09291(.A1(new_n2452_), .A2(new_n4699_), .B(new_n9547_), .ZN(new_n9548_));
  XOR2_X1    g09292(.A1(new_n9548_), .A2(new_n4446_), .Z(new_n9549_));
  INV_X1     g09293(.I(new_n9549_), .ZN(new_n9550_));
  OAI21_X1   g09294(.A1(new_n9545_), .A2(new_n9538_), .B(new_n9550_), .ZN(new_n9551_));
  NAND3_X1   g09295(.A1(new_n9541_), .A2(new_n9544_), .A3(new_n9539_), .ZN(new_n9552_));
  OAI21_X1   g09296(.A1(new_n9445_), .A2(new_n9444_), .B(new_n9537_), .ZN(new_n9553_));
  NAND3_X1   g09297(.A1(new_n9553_), .A2(new_n9552_), .A3(new_n9549_), .ZN(new_n9554_));
  NAND2_X1   g09298(.A1(new_n9551_), .A2(new_n9554_), .ZN(new_n9555_));
  NOR3_X1    g09299(.A1(new_n9443_), .A2(new_n9555_), .A3(new_n9207_), .ZN(new_n9556_));
  OAI21_X1   g09300(.A1(new_n9214_), .A2(new_n8891_), .B(new_n9216_), .ZN(new_n9557_));
  AOI21_X1   g09301(.A1(new_n9553_), .A2(new_n9552_), .B(new_n9549_), .ZN(new_n9558_));
  NOR3_X1    g09302(.A1(new_n9545_), .A2(new_n9538_), .A3(new_n9550_), .ZN(new_n9559_));
  NOR2_X1    g09303(.A1(new_n9559_), .A2(new_n9558_), .ZN(new_n9560_));
  AOI21_X1   g09304(.A1(new_n9557_), .A2(new_n9215_), .B(new_n9560_), .ZN(new_n9561_));
  OAI21_X1   g09305(.A1(new_n9561_), .A2(new_n9556_), .B(new_n9442_), .ZN(new_n9562_));
  INV_X1     g09306(.I(new_n9442_), .ZN(new_n9563_));
  NAND3_X1   g09307(.A1(new_n9557_), .A2(new_n9560_), .A3(new_n9215_), .ZN(new_n9564_));
  OAI21_X1   g09308(.A1(new_n9443_), .A2(new_n9207_), .B(new_n9555_), .ZN(new_n9565_));
  NAND3_X1   g09309(.A1(new_n9564_), .A2(new_n9565_), .A3(new_n9563_), .ZN(new_n9566_));
  NAND2_X1   g09310(.A1(new_n9562_), .A2(new_n9566_), .ZN(new_n9567_));
  NAND3_X1   g09311(.A1(new_n9438_), .A2(new_n9227_), .A3(new_n9567_), .ZN(new_n9568_));
  OAI21_X1   g09312(.A1(new_n9230_), .A2(new_n9223_), .B(new_n9227_), .ZN(new_n9569_));
  AOI21_X1   g09313(.A1(new_n9564_), .A2(new_n9565_), .B(new_n9563_), .ZN(new_n9570_));
  NOR3_X1    g09314(.A1(new_n9561_), .A2(new_n9556_), .A3(new_n9442_), .ZN(new_n9571_));
  NOR2_X1    g09315(.A1(new_n9571_), .A2(new_n9570_), .ZN(new_n9572_));
  NAND2_X1   g09316(.A1(new_n9569_), .A2(new_n9572_), .ZN(new_n9573_));
  AOI22_X1   g09317(.A1(new_n3267_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n3270_), .ZN(new_n9574_));
  OAI21_X1   g09318(.A1(new_n2495_), .A2(new_n3475_), .B(new_n9574_), .ZN(new_n9575_));
  AOI21_X1   g09319(.A1(new_n3407_), .A2(new_n3273_), .B(new_n9575_), .ZN(new_n9576_));
  XOR2_X1    g09320(.A1(new_n9576_), .A2(\a[29] ), .Z(new_n9577_));
  INV_X1     g09321(.I(new_n9577_), .ZN(new_n9578_));
  NAND3_X1   g09322(.A1(new_n9573_), .A2(new_n9568_), .A3(new_n9578_), .ZN(new_n9579_));
  AOI21_X1   g09323(.A1(new_n9234_), .A2(new_n8904_), .B(new_n9223_), .ZN(new_n9580_));
  NOR3_X1    g09324(.A1(new_n9580_), .A2(new_n9219_), .A3(new_n9572_), .ZN(new_n9581_));
  AOI21_X1   g09325(.A1(new_n9225_), .A2(new_n9228_), .B(new_n9219_), .ZN(new_n9582_));
  NOR2_X1    g09326(.A1(new_n9582_), .A2(new_n9567_), .ZN(new_n9583_));
  OAI21_X1   g09327(.A1(new_n9583_), .A2(new_n9581_), .B(new_n9577_), .ZN(new_n9584_));
  NAND2_X1   g09328(.A1(new_n9584_), .A2(new_n9579_), .ZN(new_n9585_));
  AOI21_X1   g09329(.A1(new_n9256_), .A2(new_n9437_), .B(new_n9585_), .ZN(new_n9586_));
  NOR3_X1    g09330(.A1(new_n9583_), .A2(new_n9581_), .A3(new_n9577_), .ZN(new_n9587_));
  AOI21_X1   g09331(.A1(new_n9573_), .A2(new_n9568_), .B(new_n9578_), .ZN(new_n9588_));
  NOR2_X1    g09332(.A1(new_n9588_), .A2(new_n9587_), .ZN(new_n9589_));
  NOR3_X1    g09333(.A1(new_n9589_), .A2(new_n9248_), .A3(new_n9436_), .ZN(new_n9590_));
  NOR3_X1    g09334(.A1(new_n9586_), .A2(new_n9590_), .A3(new_n9435_), .ZN(new_n9591_));
  OAI21_X1   g09335(.A1(new_n8906_), .A2(new_n8912_), .B(new_n8917_), .ZN(new_n9592_));
  OAI21_X1   g09336(.A1(new_n9592_), .A2(new_n9247_), .B(new_n9437_), .ZN(new_n9593_));
  NAND2_X1   g09337(.A1(new_n9593_), .A2(new_n9589_), .ZN(new_n9594_));
  NOR2_X1    g09338(.A1(new_n9244_), .A2(new_n8913_), .ZN(new_n9595_));
  AOI21_X1   g09339(.A1(new_n9595_), .A2(new_n9239_), .B(new_n9436_), .ZN(new_n9596_));
  NAND2_X1   g09340(.A1(new_n9596_), .A2(new_n9585_), .ZN(new_n9597_));
  AOI21_X1   g09341(.A1(new_n9597_), .A2(new_n9594_), .B(new_n9434_), .ZN(new_n9598_));
  NOR2_X1    g09342(.A1(new_n9598_), .A2(new_n9591_), .ZN(new_n9599_));
  NAND2_X1   g09343(.A1(new_n9430_), .A2(new_n9599_), .ZN(new_n9600_));
  NAND3_X1   g09344(.A1(new_n9597_), .A2(new_n9594_), .A3(new_n9434_), .ZN(new_n9601_));
  OAI21_X1   g09345(.A1(new_n9586_), .A2(new_n9590_), .B(new_n9435_), .ZN(new_n9602_));
  NAND2_X1   g09346(.A1(new_n9601_), .A2(new_n9602_), .ZN(new_n9603_));
  OAI21_X1   g09347(.A1(new_n9429_), .A2(new_n9257_), .B(new_n9603_), .ZN(new_n9604_));
  NAND3_X1   g09348(.A1(new_n9600_), .A2(new_n9428_), .A3(new_n9604_), .ZN(new_n9605_));
  INV_X1     g09349(.I(new_n9428_), .ZN(new_n9606_));
  NOR3_X1    g09350(.A1(new_n9603_), .A2(new_n9429_), .A3(new_n9257_), .ZN(new_n9607_));
  NOR2_X1    g09351(.A1(new_n9430_), .A2(new_n9599_), .ZN(new_n9608_));
  OAI21_X1   g09352(.A1(new_n9608_), .A2(new_n9607_), .B(new_n9606_), .ZN(new_n9609_));
  NAND2_X1   g09353(.A1(new_n9609_), .A2(new_n9605_), .ZN(new_n9610_));
  AOI21_X1   g09354(.A1(new_n9272_), .A2(new_n9424_), .B(new_n9610_), .ZN(new_n9611_));
  NOR3_X1    g09355(.A1(new_n9608_), .A2(new_n9607_), .A3(new_n9606_), .ZN(new_n9612_));
  AOI21_X1   g09356(.A1(new_n9600_), .A2(new_n9604_), .B(new_n9428_), .ZN(new_n9613_));
  NOR2_X1    g09357(.A1(new_n9612_), .A2(new_n9613_), .ZN(new_n9614_));
  NOR3_X1    g09358(.A1(new_n9614_), .A2(new_n9280_), .A3(new_n9423_), .ZN(new_n9615_));
  OAI21_X1   g09359(.A1(new_n9611_), .A2(new_n9615_), .B(new_n9422_), .ZN(new_n9616_));
  OAI21_X1   g09360(.A1(new_n8942_), .A2(new_n8943_), .B(new_n8937_), .ZN(new_n9617_));
  OAI21_X1   g09361(.A1(new_n9617_), .A2(new_n9276_), .B(new_n9424_), .ZN(new_n9618_));
  NAND2_X1   g09362(.A1(new_n9618_), .A2(new_n9614_), .ZN(new_n9619_));
  NAND3_X1   g09363(.A1(new_n9272_), .A2(new_n9610_), .A3(new_n9424_), .ZN(new_n9620_));
  NAND3_X1   g09364(.A1(new_n9619_), .A2(new_n9620_), .A3(new_n9421_), .ZN(new_n9621_));
  NAND2_X1   g09365(.A1(new_n9621_), .A2(new_n9616_), .ZN(new_n9622_));
  AOI21_X1   g09366(.A1(new_n9295_), .A2(new_n9278_), .B(new_n9622_), .ZN(new_n9623_));
  AOI21_X1   g09367(.A1(new_n9619_), .A2(new_n9620_), .B(new_n9421_), .ZN(new_n9624_));
  NOR3_X1    g09368(.A1(new_n9611_), .A2(new_n9615_), .A3(new_n9422_), .ZN(new_n9625_));
  NOR2_X1    g09369(.A1(new_n9624_), .A2(new_n9625_), .ZN(new_n9626_));
  NOR3_X1    g09370(.A1(new_n9626_), .A2(new_n9284_), .A3(new_n9289_), .ZN(new_n9627_));
  OAI21_X1   g09371(.A1(new_n9623_), .A2(new_n9627_), .B(new_n9417_), .ZN(new_n9628_));
  OAI21_X1   g09372(.A1(new_n9289_), .A2(new_n9284_), .B(new_n9626_), .ZN(new_n9629_));
  NAND3_X1   g09373(.A1(new_n9295_), .A2(new_n9622_), .A3(new_n9278_), .ZN(new_n9630_));
  NAND3_X1   g09374(.A1(new_n9629_), .A2(new_n9630_), .A3(new_n9416_), .ZN(new_n9631_));
  NAND2_X1   g09375(.A1(new_n9628_), .A2(new_n9631_), .ZN(new_n9632_));
  NOR3_X1    g09376(.A1(new_n9292_), .A2(new_n9284_), .A3(new_n9294_), .ZN(new_n9633_));
  INV_X1     g09377(.I(new_n9633_), .ZN(new_n9634_));
  AOI21_X1   g09378(.A1(new_n9299_), .A2(new_n9634_), .B(new_n9632_), .ZN(new_n9635_));
  AOI21_X1   g09379(.A1(new_n9629_), .A2(new_n9630_), .B(new_n9416_), .ZN(new_n9636_));
  NOR3_X1    g09380(.A1(new_n9623_), .A2(new_n9627_), .A3(new_n9417_), .ZN(new_n9637_));
  NOR2_X1    g09381(.A1(new_n9636_), .A2(new_n9637_), .ZN(new_n9638_));
  NOR3_X1    g09382(.A1(new_n9310_), .A2(new_n9638_), .A3(new_n9633_), .ZN(new_n9639_));
  OAI21_X1   g09383(.A1(new_n9635_), .A2(new_n9639_), .B(new_n9412_), .ZN(new_n9640_));
  AOI21_X1   g09384(.A1(new_n9410_), .A2(new_n9409_), .B(new_n1002_), .ZN(new_n9641_));
  NOR2_X1    g09385(.A1(new_n9411_), .A2(\a[14] ), .ZN(new_n9642_));
  NOR2_X1    g09386(.A1(new_n9642_), .A2(new_n9641_), .ZN(new_n9643_));
  OAI21_X1   g09387(.A1(new_n9310_), .A2(new_n9633_), .B(new_n9638_), .ZN(new_n9644_));
  NAND3_X1   g09388(.A1(new_n9299_), .A2(new_n9632_), .A3(new_n9634_), .ZN(new_n9645_));
  NAND3_X1   g09389(.A1(new_n9644_), .A2(new_n9645_), .A3(new_n9643_), .ZN(new_n9646_));
  NAND2_X1   g09390(.A1(new_n9640_), .A2(new_n9646_), .ZN(new_n9647_));
  AOI21_X1   g09391(.A1(new_n9326_), .A2(new_n9308_), .B(new_n9647_), .ZN(new_n9648_));
  AOI21_X1   g09392(.A1(new_n9644_), .A2(new_n9645_), .B(new_n9643_), .ZN(new_n9649_));
  NOR3_X1    g09393(.A1(new_n9635_), .A2(new_n9639_), .A3(new_n9412_), .ZN(new_n9650_));
  NOR2_X1    g09394(.A1(new_n9650_), .A2(new_n9649_), .ZN(new_n9651_));
  NOR3_X1    g09395(.A1(new_n9314_), .A2(new_n9316_), .A3(new_n9651_), .ZN(new_n9652_));
  NOR3_X1    g09396(.A1(new_n9652_), .A2(new_n9648_), .A3(new_n9406_), .ZN(new_n9653_));
  XOR2_X1    g09397(.A1(new_n9405_), .A2(\a[11] ), .Z(new_n9654_));
  OAI21_X1   g09398(.A1(new_n9314_), .A2(new_n9316_), .B(new_n9651_), .ZN(new_n9655_));
  NAND3_X1   g09399(.A1(new_n9326_), .A2(new_n9647_), .A3(new_n9308_), .ZN(new_n9656_));
  AOI21_X1   g09400(.A1(new_n9655_), .A2(new_n9656_), .B(new_n9654_), .ZN(new_n9657_));
  NOR2_X1    g09401(.A1(new_n9653_), .A2(new_n9657_), .ZN(new_n9658_));
  OAI21_X1   g09402(.A1(new_n9402_), .A2(new_n9333_), .B(new_n9658_), .ZN(new_n9659_));
  OAI21_X1   g09403(.A1(new_n9059_), .A2(new_n8995_), .B(new_n9329_), .ZN(new_n9660_));
  NAND3_X1   g09404(.A1(new_n9655_), .A2(new_n9656_), .A3(new_n9654_), .ZN(new_n9661_));
  OAI21_X1   g09405(.A1(new_n9652_), .A2(new_n9648_), .B(new_n9406_), .ZN(new_n9662_));
  NAND2_X1   g09406(.A1(new_n9662_), .A2(new_n9661_), .ZN(new_n9663_));
  NAND3_X1   g09407(.A1(new_n9660_), .A2(new_n9320_), .A3(new_n9663_), .ZN(new_n9664_));
  NAND3_X1   g09408(.A1(new_n9659_), .A2(new_n9664_), .A3(new_n9397_), .ZN(new_n9665_));
  INV_X1     g09409(.I(new_n9394_), .ZN(new_n9666_));
  NAND2_X1   g09410(.A1(new_n9666_), .A2(new_n9395_), .ZN(new_n9667_));
  AOI21_X1   g09411(.A1(new_n9660_), .A2(new_n9320_), .B(new_n9663_), .ZN(new_n9668_));
  NOR3_X1    g09412(.A1(new_n9402_), .A2(new_n9333_), .A3(new_n9658_), .ZN(new_n9669_));
  OAI21_X1   g09413(.A1(new_n9669_), .A2(new_n9668_), .B(new_n9667_), .ZN(new_n9670_));
  NAND2_X1   g09414(.A1(new_n9670_), .A2(new_n9665_), .ZN(new_n9671_));
  OAI21_X1   g09415(.A1(new_n9389_), .A2(new_n9355_), .B(new_n9671_), .ZN(new_n9672_));
  NAND3_X1   g09416(.A1(new_n9352_), .A2(new_n9009_), .A3(new_n9343_), .ZN(new_n9673_));
  NOR3_X1    g09417(.A1(new_n9669_), .A2(new_n9668_), .A3(new_n9667_), .ZN(new_n9674_));
  AOI21_X1   g09418(.A1(new_n9659_), .A2(new_n9664_), .B(new_n9397_), .ZN(new_n9675_));
  NOR2_X1    g09419(.A1(new_n9674_), .A2(new_n9675_), .ZN(new_n9676_));
  NAND3_X1   g09420(.A1(new_n9673_), .A2(new_n9676_), .A3(new_n9346_), .ZN(new_n9677_));
  NAND2_X1   g09421(.A1(new_n9672_), .A2(new_n9677_), .ZN(new_n9678_));
  INV_X1     g09422(.I(new_n9678_), .ZN(new_n9679_));
  NAND3_X1   g09423(.A1(new_n8789_), .A2(new_n9021_), .A3(new_n8788_), .ZN(new_n9680_));
  NAND3_X1   g09424(.A1(new_n9361_), .A2(new_n9054_), .A3(new_n9362_), .ZN(new_n9681_));
  OAI21_X1   g09425(.A1(new_n9353_), .A2(new_n9359_), .B(new_n9055_), .ZN(new_n9682_));
  AOI22_X1   g09426(.A1(new_n9680_), .A2(new_n9020_), .B1(new_n9681_), .B2(new_n9682_), .ZN(new_n9683_));
  INV_X1     g09427(.I(new_n8510_), .ZN(new_n9684_));
  AOI22_X1   g09428(.A1(new_n800_), .A2(\b[49] ), .B1(\b[50] ), .B2(new_n333_), .ZN(new_n9685_));
  OAI21_X1   g09429(.A1(new_n8127_), .A2(new_n392_), .B(new_n9685_), .ZN(new_n9686_));
  AOI21_X1   g09430(.A1(new_n9684_), .A2(new_n330_), .B(new_n9686_), .ZN(new_n9687_));
  XOR2_X1    g09431(.A1(new_n9687_), .A2(new_n312_), .Z(new_n9688_));
  AOI21_X1   g09432(.A1(new_n9361_), .A2(new_n9362_), .B(new_n9055_), .ZN(new_n9689_));
  OAI21_X1   g09433(.A1(new_n9683_), .A2(new_n9689_), .B(new_n9688_), .ZN(new_n9690_));
  INV_X1     g09434(.I(new_n9688_), .ZN(new_n9691_));
  INV_X1     g09435(.I(new_n9689_), .ZN(new_n9692_));
  NAND3_X1   g09436(.A1(new_n9364_), .A2(new_n9691_), .A3(new_n9692_), .ZN(new_n9693_));
  NAND3_X1   g09437(.A1(new_n9693_), .A2(new_n9690_), .A3(new_n9679_), .ZN(new_n9694_));
  INV_X1     g09438(.I(new_n9694_), .ZN(new_n9695_));
  AOI21_X1   g09439(.A1(new_n9693_), .A2(new_n9690_), .B(new_n9679_), .ZN(new_n9696_));
  OAI21_X1   g09440(.A1(new_n9695_), .A2(new_n9696_), .B(new_n9388_), .ZN(new_n9697_));
  INV_X1     g09441(.I(new_n9696_), .ZN(new_n9698_));
  NAND3_X1   g09442(.A1(new_n9698_), .A2(new_n9694_), .A3(new_n9387_), .ZN(new_n9699_));
  NAND2_X1   g09443(.A1(new_n9699_), .A2(new_n9697_), .ZN(new_n9700_));
  XOR2_X1    g09444(.A1(new_n9700_), .A2(new_n9375_), .Z(\f[53] ));
  AOI21_X1   g09445(.A1(new_n9698_), .A2(new_n9694_), .B(new_n9387_), .ZN(new_n9702_));
  AOI21_X1   g09446(.A1(new_n9375_), .A2(new_n9699_), .B(new_n9702_), .ZN(new_n9703_));
  AOI22_X1   g09447(.A1(new_n800_), .A2(\b[50] ), .B1(\b[51] ), .B2(new_n333_), .ZN(new_n9704_));
  OAI21_X1   g09448(.A1(new_n8168_), .A2(new_n392_), .B(new_n9704_), .ZN(new_n9705_));
  AOI21_X1   g09449(.A1(new_n8783_), .A2(new_n330_), .B(new_n9705_), .ZN(new_n9706_));
  XOR2_X1    g09450(.A1(new_n9706_), .A2(new_n312_), .Z(new_n9707_));
  INV_X1     g09451(.I(new_n9707_), .ZN(new_n9708_));
  NOR2_X1    g09452(.A1(new_n9445_), .A2(new_n9444_), .ZN(new_n9709_));
  AOI21_X1   g09453(.A1(new_n9709_), .A2(new_n9543_), .B(new_n9532_), .ZN(new_n9710_));
  INV_X1     g09454(.I(new_n9710_), .ZN(new_n9711_));
  AOI22_X1   g09455(.A1(new_n5155_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n5160_), .ZN(new_n9712_));
  OAI21_X1   g09456(.A1(new_n1296_), .A2(new_n6877_), .B(new_n9712_), .ZN(new_n9713_));
  AOI21_X1   g09457(.A1(new_n2038_), .A2(new_n5166_), .B(new_n9713_), .ZN(new_n9714_));
  XOR2_X1    g09458(.A1(new_n9714_), .A2(new_n5162_), .Z(new_n9715_));
  INV_X1     g09459(.I(new_n9715_), .ZN(new_n9716_));
  AOI21_X1   g09460(.A1(new_n9509_), .A2(new_n9496_), .B(new_n9499_), .ZN(new_n9717_));
  AOI21_X1   g09461(.A1(new_n9459_), .A2(new_n9142_), .B(new_n9483_), .ZN(new_n9718_));
  NOR2_X1    g09462(.A1(new_n9718_), .A2(new_n9482_), .ZN(new_n9719_));
  OAI22_X1   g09463(.A1(new_n9461_), .A2(new_n438_), .B1(new_n377_), .B2(new_n9462_), .ZN(new_n9720_));
  AOI21_X1   g09464(.A1(\b[4] ), .A2(new_n8575_), .B(new_n9720_), .ZN(new_n9721_));
  OAI21_X1   g09465(.A1(new_n450_), .A2(new_n9460_), .B(new_n9721_), .ZN(new_n9722_));
  XOR2_X1    g09466(.A1(new_n9722_), .A2(\a[50] ), .Z(new_n9723_));
  INV_X1     g09467(.I(new_n9723_), .ZN(new_n9724_));
  AOI22_X1   g09468(.A1(new_n9125_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n9123_), .ZN(new_n9725_));
  OAI21_X1   g09469(.A1(new_n275_), .A2(new_n9470_), .B(new_n9725_), .ZN(new_n9726_));
  AOI21_X1   g09470(.A1(new_n299_), .A2(new_n9129_), .B(new_n9726_), .ZN(new_n9727_));
  XOR2_X1    g09471(.A1(new_n9727_), .A2(new_n9133_), .Z(new_n9728_));
  XNOR2_X1   g09472(.A1(\a[53] ), .A2(\a[54] ), .ZN(new_n9729_));
  NOR2_X1    g09473(.A1(new_n9729_), .A2(new_n258_), .ZN(new_n9730_));
  NAND2_X1   g09474(.A1(new_n9728_), .A2(new_n9730_), .ZN(new_n9731_));
  XOR2_X1    g09475(.A1(new_n9727_), .A2(\a[53] ), .Z(new_n9732_));
  INV_X1     g09476(.I(new_n9730_), .ZN(new_n9733_));
  NAND2_X1   g09477(.A1(new_n9732_), .A2(new_n9733_), .ZN(new_n9734_));
  NAND2_X1   g09478(.A1(new_n9731_), .A2(new_n9734_), .ZN(new_n9735_));
  XOR2_X1    g09479(.A1(new_n9735_), .A2(new_n9479_), .Z(new_n9736_));
  AND2_X2    g09480(.A1(new_n9736_), .A2(new_n9724_), .Z(new_n9737_));
  NOR2_X1    g09481(.A1(new_n9736_), .A2(new_n9724_), .ZN(new_n9738_));
  NOR2_X1    g09482(.A1(new_n9737_), .A2(new_n9738_), .ZN(new_n9739_));
  XOR2_X1    g09483(.A1(new_n9739_), .A2(new_n9719_), .Z(new_n9740_));
  AOI22_X1   g09484(.A1(new_n7403_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n7408_), .ZN(new_n9741_));
  OAI21_X1   g09485(.A1(new_n471_), .A2(new_n9488_), .B(new_n9741_), .ZN(new_n9742_));
  AOI21_X1   g09486(.A1(new_n676_), .A2(new_n7414_), .B(new_n9742_), .ZN(new_n9743_));
  XOR2_X1    g09487(.A1(new_n9743_), .A2(new_n7410_), .Z(new_n9744_));
  INV_X1     g09488(.I(new_n9744_), .ZN(new_n9745_));
  XOR2_X1    g09489(.A1(new_n9740_), .A2(new_n9745_), .Z(new_n9746_));
  XOR2_X1    g09490(.A1(new_n9746_), .A2(new_n9717_), .Z(new_n9747_));
  INV_X1     g09491(.I(new_n9747_), .ZN(new_n9748_));
  AOI22_X1   g09492(.A1(new_n6569_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n6574_), .ZN(new_n9749_));
  OAI21_X1   g09493(.A1(new_n776_), .A2(new_n8565_), .B(new_n9749_), .ZN(new_n9750_));
  AOI21_X1   g09494(.A1(new_n1194_), .A2(new_n6579_), .B(new_n9750_), .ZN(new_n9751_));
  XOR2_X1    g09495(.A1(new_n9751_), .A2(new_n6567_), .Z(new_n9752_));
  NAND2_X1   g09496(.A1(new_n9522_), .A2(new_n9507_), .ZN(new_n9753_));
  NAND2_X1   g09497(.A1(new_n9753_), .A2(new_n9752_), .ZN(new_n9754_));
  INV_X1     g09498(.I(new_n9754_), .ZN(new_n9755_));
  NOR2_X1    g09499(.A1(new_n9753_), .A2(new_n9752_), .ZN(new_n9756_));
  NOR3_X1    g09500(.A1(new_n9755_), .A2(new_n9748_), .A3(new_n9756_), .ZN(new_n9757_));
  INV_X1     g09501(.I(new_n9756_), .ZN(new_n9758_));
  AOI21_X1   g09502(.A1(new_n9758_), .A2(new_n9754_), .B(new_n9747_), .ZN(new_n9759_));
  NOR2_X1    g09503(.A1(new_n9759_), .A2(new_n9757_), .ZN(new_n9760_));
  OAI22_X1   g09504(.A1(new_n5852_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n5857_), .ZN(new_n9761_));
  AOI21_X1   g09505(.A1(\b[13] ), .A2(new_n6115_), .B(new_n9761_), .ZN(new_n9762_));
  OAI21_X1   g09506(.A1(new_n1275_), .A2(new_n5861_), .B(new_n9762_), .ZN(new_n9763_));
  XOR2_X1    g09507(.A1(new_n9763_), .A2(\a[41] ), .Z(new_n9764_));
  AOI21_X1   g09508(.A1(new_n9185_), .A2(new_n9450_), .B(new_n9530_), .ZN(new_n9765_));
  NOR3_X1    g09509(.A1(new_n9520_), .A2(new_n9454_), .A3(new_n9515_), .ZN(new_n9766_));
  OAI21_X1   g09510(.A1(new_n9765_), .A2(new_n9766_), .B(new_n9764_), .ZN(new_n9767_));
  NOR3_X1    g09511(.A1(new_n9765_), .A2(new_n9764_), .A3(new_n9766_), .ZN(new_n9768_));
  INV_X1     g09512(.I(new_n9768_), .ZN(new_n9769_));
  NAND3_X1   g09513(.A1(new_n9769_), .A2(new_n9760_), .A3(new_n9767_), .ZN(new_n9770_));
  AOI21_X1   g09514(.A1(new_n9769_), .A2(new_n9767_), .B(new_n9760_), .ZN(new_n9771_));
  INV_X1     g09515(.I(new_n9771_), .ZN(new_n9772_));
  NAND3_X1   g09516(.A1(new_n9772_), .A2(new_n9770_), .A3(new_n9716_), .ZN(new_n9773_));
  INV_X1     g09517(.I(new_n9770_), .ZN(new_n9774_));
  OAI21_X1   g09518(.A1(new_n9774_), .A2(new_n9771_), .B(new_n9715_), .ZN(new_n9775_));
  NAND2_X1   g09519(.A1(new_n9773_), .A2(new_n9775_), .ZN(new_n9776_));
  XOR2_X1    g09520(.A1(new_n9776_), .A2(new_n9711_), .Z(new_n9777_));
  AOI22_X1   g09521(.A1(new_n4918_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n4921_), .ZN(new_n9778_));
  OAI21_X1   g09522(.A1(new_n1859_), .A2(new_n6099_), .B(new_n9778_), .ZN(new_n9779_));
  AOI21_X1   g09523(.A1(new_n2032_), .A2(new_n4699_), .B(new_n9779_), .ZN(new_n9780_));
  XOR2_X1    g09524(.A1(new_n9780_), .A2(new_n4446_), .Z(new_n9781_));
  INV_X1     g09525(.I(new_n9781_), .ZN(new_n9782_));
  AOI21_X1   g09526(.A1(new_n9564_), .A2(new_n9554_), .B(new_n9782_), .ZN(new_n9783_));
  NOR3_X1    g09527(.A1(new_n9556_), .A2(new_n9559_), .A3(new_n9781_), .ZN(new_n9784_));
  NOR3_X1    g09528(.A1(new_n9783_), .A2(new_n9784_), .A3(new_n9777_), .ZN(new_n9785_));
  XOR2_X1    g09529(.A1(new_n9776_), .A2(new_n9710_), .Z(new_n9786_));
  OAI21_X1   g09530(.A1(new_n9556_), .A2(new_n9559_), .B(new_n9781_), .ZN(new_n9787_));
  NAND3_X1   g09531(.A1(new_n9564_), .A2(new_n9554_), .A3(new_n9782_), .ZN(new_n9788_));
  AOI21_X1   g09532(.A1(new_n9788_), .A2(new_n9787_), .B(new_n9786_), .ZN(new_n9789_));
  NOR2_X1    g09533(.A1(new_n9785_), .A2(new_n9789_), .ZN(new_n9790_));
  AOI22_X1   g09534(.A1(new_n3864_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n3869_), .ZN(new_n9791_));
  OAI21_X1   g09535(.A1(new_n2142_), .A2(new_n5410_), .B(new_n9791_), .ZN(new_n9792_));
  AOI21_X1   g09536(.A1(new_n3033_), .A2(new_n3872_), .B(new_n9792_), .ZN(new_n9793_));
  XOR2_X1    g09537(.A1(new_n9793_), .A2(new_n3876_), .Z(new_n9794_));
  NOR3_X1    g09538(.A1(new_n9561_), .A2(new_n9556_), .A3(new_n9563_), .ZN(new_n9795_));
  OAI21_X1   g09539(.A1(new_n9581_), .A2(new_n9795_), .B(new_n9794_), .ZN(new_n9796_));
  INV_X1     g09540(.I(new_n9794_), .ZN(new_n9797_));
  INV_X1     g09541(.I(new_n9795_), .ZN(new_n9798_));
  NAND3_X1   g09542(.A1(new_n9568_), .A2(new_n9797_), .A3(new_n9798_), .ZN(new_n9799_));
  NAND3_X1   g09543(.A1(new_n9796_), .A2(new_n9799_), .A3(new_n9790_), .ZN(new_n9800_));
  INV_X1     g09544(.I(new_n9800_), .ZN(new_n9801_));
  AOI21_X1   g09545(.A1(new_n9796_), .A2(new_n9799_), .B(new_n9790_), .ZN(new_n9802_));
  NOR2_X1    g09546(.A1(new_n9801_), .A2(new_n9802_), .ZN(new_n9803_));
  OAI22_X1   g09547(.A1(new_n3158_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n3006_), .ZN(new_n9804_));
  AOI21_X1   g09548(.A1(\b[25] ), .A2(new_n3456_), .B(new_n9804_), .ZN(new_n9805_));
  OAI21_X1   g09549(.A1(new_n3165_), .A2(new_n3261_), .B(new_n9805_), .ZN(new_n9806_));
  XOR2_X1    g09550(.A1(new_n9806_), .A2(\a[29] ), .Z(new_n9807_));
  OAI21_X1   g09551(.A1(new_n9586_), .A2(new_n9587_), .B(new_n9807_), .ZN(new_n9808_));
  INV_X1     g09552(.I(new_n9807_), .ZN(new_n9809_));
  NAND3_X1   g09553(.A1(new_n9594_), .A2(new_n9579_), .A3(new_n9809_), .ZN(new_n9810_));
  AND3_X2    g09554(.A1(new_n9810_), .A2(new_n9803_), .A3(new_n9808_), .Z(new_n9811_));
  AOI21_X1   g09555(.A1(new_n9810_), .A2(new_n9808_), .B(new_n9803_), .ZN(new_n9812_));
  NOR2_X1    g09556(.A1(new_n9811_), .A2(new_n9812_), .ZN(new_n9813_));
  AOI22_X1   g09557(.A1(new_n2716_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n2719_), .ZN(new_n9814_));
  OAI21_X1   g09558(.A1(new_n3185_), .A2(new_n2924_), .B(new_n9814_), .ZN(new_n9815_));
  AOI21_X1   g09559(.A1(new_n4230_), .A2(new_n2722_), .B(new_n9815_), .ZN(new_n9816_));
  XOR2_X1    g09560(.A1(new_n9816_), .A2(new_n2714_), .Z(new_n9817_));
  NOR2_X1    g09561(.A1(new_n9093_), .A2(new_n9092_), .ZN(new_n9818_));
  OAI21_X1   g09562(.A1(new_n9818_), .A2(new_n9254_), .B(new_n9263_), .ZN(new_n9819_));
  OAI21_X1   g09563(.A1(new_n9819_), .A2(new_n9603_), .B(new_n9601_), .ZN(new_n9820_));
  NAND2_X1   g09564(.A1(new_n9820_), .A2(new_n9817_), .ZN(new_n9821_));
  INV_X1     g09565(.I(new_n9817_), .ZN(new_n9822_));
  AOI21_X1   g09566(.A1(new_n9430_), .A2(new_n9599_), .B(new_n9591_), .ZN(new_n9823_));
  NAND2_X1   g09567(.A1(new_n9823_), .A2(new_n9822_), .ZN(new_n9824_));
  NAND3_X1   g09568(.A1(new_n9821_), .A2(new_n9824_), .A3(new_n9813_), .ZN(new_n9825_));
  NAND3_X1   g09569(.A1(new_n9810_), .A2(new_n9808_), .A3(new_n9803_), .ZN(new_n9826_));
  INV_X1     g09570(.I(new_n9812_), .ZN(new_n9827_));
  NAND2_X1   g09571(.A1(new_n9827_), .A2(new_n9826_), .ZN(new_n9828_));
  NOR2_X1    g09572(.A1(new_n9823_), .A2(new_n9822_), .ZN(new_n9829_));
  NOR2_X1    g09573(.A1(new_n9820_), .A2(new_n9817_), .ZN(new_n9830_));
  OAI21_X1   g09574(.A1(new_n9830_), .A2(new_n9829_), .B(new_n9828_), .ZN(new_n9831_));
  NAND2_X1   g09575(.A1(new_n9831_), .A2(new_n9825_), .ZN(new_n9832_));
  AOI22_X1   g09576(.A1(new_n2202_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n2205_), .ZN(new_n9833_));
  OAI21_X1   g09577(.A1(new_n4022_), .A2(new_n2370_), .B(new_n9833_), .ZN(new_n9834_));
  AOI21_X1   g09578(.A1(new_n4223_), .A2(new_n2208_), .B(new_n9834_), .ZN(new_n9835_));
  XOR2_X1    g09579(.A1(new_n9835_), .A2(new_n2200_), .Z(new_n9836_));
  INV_X1     g09580(.I(new_n9836_), .ZN(new_n9837_));
  AOI21_X1   g09581(.A1(new_n9618_), .A2(new_n9614_), .B(new_n9612_), .ZN(new_n9838_));
  NOR2_X1    g09582(.A1(new_n9838_), .A2(new_n9837_), .ZN(new_n9839_));
  NOR2_X1    g09583(.A1(new_n9280_), .A2(new_n9423_), .ZN(new_n9840_));
  OAI21_X1   g09584(.A1(new_n9840_), .A2(new_n9610_), .B(new_n9605_), .ZN(new_n9841_));
  NOR2_X1    g09585(.A1(new_n9841_), .A2(new_n9836_), .ZN(new_n9842_));
  NOR3_X1    g09586(.A1(new_n9842_), .A2(new_n9839_), .A3(new_n9832_), .ZN(new_n9843_));
  NOR3_X1    g09587(.A1(new_n9830_), .A2(new_n9829_), .A3(new_n9828_), .ZN(new_n9844_));
  AOI21_X1   g09588(.A1(new_n9821_), .A2(new_n9824_), .B(new_n9813_), .ZN(new_n9845_));
  NOR2_X1    g09589(.A1(new_n9844_), .A2(new_n9845_), .ZN(new_n9846_));
  NAND2_X1   g09590(.A1(new_n9841_), .A2(new_n9836_), .ZN(new_n9847_));
  NAND2_X1   g09591(.A1(new_n9838_), .A2(new_n9837_), .ZN(new_n9848_));
  AOI21_X1   g09592(.A1(new_n9847_), .A2(new_n9848_), .B(new_n9846_), .ZN(new_n9849_));
  NOR2_X1    g09593(.A1(new_n9843_), .A2(new_n9849_), .ZN(new_n9850_));
  AOI22_X1   g09594(.A1(new_n1738_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n1743_), .ZN(new_n9851_));
  OAI21_X1   g09595(.A1(new_n4639_), .A2(new_n1931_), .B(new_n9851_), .ZN(new_n9852_));
  AOI21_X1   g09596(.A1(new_n5594_), .A2(new_n1746_), .B(new_n9852_), .ZN(new_n9853_));
  XOR2_X1    g09597(.A1(new_n9853_), .A2(new_n1736_), .Z(new_n9854_));
  NOR2_X1    g09598(.A1(new_n9284_), .A2(new_n9289_), .ZN(new_n9855_));
  OAI21_X1   g09599(.A1(new_n9855_), .A2(new_n9622_), .B(new_n9621_), .ZN(new_n9856_));
  NAND2_X1   g09600(.A1(new_n9856_), .A2(new_n9854_), .ZN(new_n9857_));
  INV_X1     g09601(.I(new_n9854_), .ZN(new_n9858_));
  NAND2_X1   g09602(.A1(new_n9295_), .A2(new_n9278_), .ZN(new_n9859_));
  AOI21_X1   g09603(.A1(new_n9859_), .A2(new_n9626_), .B(new_n9625_), .ZN(new_n9860_));
  NAND2_X1   g09604(.A1(new_n9860_), .A2(new_n9858_), .ZN(new_n9861_));
  NAND3_X1   g09605(.A1(new_n9861_), .A2(new_n9857_), .A3(new_n9850_), .ZN(new_n9862_));
  NAND3_X1   g09606(.A1(new_n9847_), .A2(new_n9848_), .A3(new_n9846_), .ZN(new_n9863_));
  OAI21_X1   g09607(.A1(new_n9842_), .A2(new_n9839_), .B(new_n9832_), .ZN(new_n9864_));
  NAND2_X1   g09608(.A1(new_n9864_), .A2(new_n9863_), .ZN(new_n9865_));
  NOR2_X1    g09609(.A1(new_n9860_), .A2(new_n9858_), .ZN(new_n9866_));
  NOR2_X1    g09610(.A1(new_n9856_), .A2(new_n9854_), .ZN(new_n9867_));
  OAI21_X1   g09611(.A1(new_n9866_), .A2(new_n9867_), .B(new_n9865_), .ZN(new_n9868_));
  NAND2_X1   g09612(.A1(new_n9868_), .A2(new_n9862_), .ZN(new_n9869_));
  OAI22_X1   g09613(.A1(new_n1592_), .A2(new_n5761_), .B1(new_n5341_), .B2(new_n1505_), .ZN(new_n9870_));
  AOI21_X1   g09614(.A1(\b[37] ), .A2(new_n1584_), .B(new_n9870_), .ZN(new_n9871_));
  OAI21_X1   g09615(.A1(new_n6309_), .A2(new_n1732_), .B(new_n9871_), .ZN(new_n9872_));
  XOR2_X1    g09616(.A1(new_n9872_), .A2(\a[17] ), .Z(new_n9873_));
  OAI21_X1   g09617(.A1(new_n9635_), .A2(new_n9637_), .B(new_n9873_), .ZN(new_n9874_));
  INV_X1     g09618(.I(new_n9874_), .ZN(new_n9875_));
  NOR2_X1    g09619(.A1(new_n9310_), .A2(new_n9633_), .ZN(new_n9876_));
  OAI21_X1   g09620(.A1(new_n9876_), .A2(new_n9632_), .B(new_n9631_), .ZN(new_n9877_));
  NOR2_X1    g09621(.A1(new_n9877_), .A2(new_n9873_), .ZN(new_n9878_));
  NOR3_X1    g09622(.A1(new_n9875_), .A2(new_n9878_), .A3(new_n9869_), .ZN(new_n9879_));
  NOR3_X1    g09623(.A1(new_n9866_), .A2(new_n9867_), .A3(new_n9865_), .ZN(new_n9880_));
  AOI21_X1   g09624(.A1(new_n9861_), .A2(new_n9857_), .B(new_n9850_), .ZN(new_n9881_));
  NOR2_X1    g09625(.A1(new_n9881_), .A2(new_n9880_), .ZN(new_n9882_));
  INV_X1     g09626(.I(new_n9873_), .ZN(new_n9883_));
  OAI21_X1   g09627(.A1(new_n8962_), .A2(new_n8968_), .B(new_n9072_), .ZN(new_n9884_));
  OAI21_X1   g09628(.A1(new_n9884_), .A2(new_n9306_), .B(new_n9634_), .ZN(new_n9885_));
  AOI21_X1   g09629(.A1(new_n9885_), .A2(new_n9638_), .B(new_n9637_), .ZN(new_n9886_));
  NAND2_X1   g09630(.A1(new_n9886_), .A2(new_n9883_), .ZN(new_n9887_));
  AOI21_X1   g09631(.A1(new_n9887_), .A2(new_n9874_), .B(new_n9882_), .ZN(new_n9888_));
  NOR2_X1    g09632(.A1(new_n9879_), .A2(new_n9888_), .ZN(new_n9889_));
  OAI22_X1   g09633(.A1(new_n993_), .A2(new_n6490_), .B1(new_n6285_), .B2(new_n997_), .ZN(new_n9890_));
  AOI21_X1   g09634(.A1(\b[40] ), .A2(new_n1486_), .B(new_n9890_), .ZN(new_n9891_));
  OAI21_X1   g09635(.A1(new_n8988_), .A2(new_n1323_), .B(new_n9891_), .ZN(new_n9892_));
  XOR2_X1    g09636(.A1(new_n9892_), .A2(\a[14] ), .Z(new_n9893_));
  OAI21_X1   g09637(.A1(new_n9648_), .A2(new_n9650_), .B(new_n9893_), .ZN(new_n9894_));
  INV_X1     g09638(.I(new_n9893_), .ZN(new_n9895_));
  NAND3_X1   g09639(.A1(new_n9655_), .A2(new_n9646_), .A3(new_n9895_), .ZN(new_n9896_));
  NAND3_X1   g09640(.A1(new_n9896_), .A2(new_n9894_), .A3(new_n9889_), .ZN(new_n9897_));
  AOI21_X1   g09641(.A1(new_n9896_), .A2(new_n9894_), .B(new_n9889_), .ZN(new_n9898_));
  INV_X1     g09642(.I(new_n9898_), .ZN(new_n9899_));
  NAND2_X1   g09643(.A1(new_n9899_), .A2(new_n9897_), .ZN(new_n9900_));
  OAI22_X1   g09644(.A1(new_n713_), .A2(new_n7096_), .B1(new_n7074_), .B2(new_n717_), .ZN(new_n9901_));
  AOI21_X1   g09645(.A1(\b[43] ), .A2(new_n1126_), .B(new_n9901_), .ZN(new_n9902_));
  OAI21_X1   g09646(.A1(new_n7925_), .A2(new_n986_), .B(new_n9902_), .ZN(new_n9903_));
  XOR2_X1    g09647(.A1(new_n9903_), .A2(\a[11] ), .Z(new_n9904_));
  INV_X1     g09648(.I(new_n9904_), .ZN(new_n9905_));
  OAI21_X1   g09649(.A1(new_n8987_), .A2(new_n8994_), .B(new_n8999_), .ZN(new_n9906_));
  AOI21_X1   g09650(.A1(new_n9906_), .A2(new_n9329_), .B(new_n9333_), .ZN(new_n9907_));
  AOI21_X1   g09651(.A1(new_n9907_), .A2(new_n9658_), .B(new_n9653_), .ZN(new_n9908_));
  NOR2_X1    g09652(.A1(new_n9908_), .A2(new_n9905_), .ZN(new_n9909_));
  OAI21_X1   g09653(.A1(new_n9332_), .A2(new_n9334_), .B(new_n9320_), .ZN(new_n9910_));
  OAI21_X1   g09654(.A1(new_n9910_), .A2(new_n9663_), .B(new_n9661_), .ZN(new_n9911_));
  NOR2_X1    g09655(.A1(new_n9911_), .A2(new_n9904_), .ZN(new_n9912_));
  NOR3_X1    g09656(.A1(new_n9909_), .A2(new_n9912_), .A3(new_n9900_), .ZN(new_n9913_));
  INV_X1     g09657(.I(new_n9897_), .ZN(new_n9914_));
  NOR2_X1    g09658(.A1(new_n9914_), .A2(new_n9898_), .ZN(new_n9915_));
  NAND2_X1   g09659(.A1(new_n9911_), .A2(new_n9904_), .ZN(new_n9916_));
  NAND2_X1   g09660(.A1(new_n9908_), .A2(new_n9905_), .ZN(new_n9917_));
  AOI21_X1   g09661(.A1(new_n9917_), .A2(new_n9916_), .B(new_n9915_), .ZN(new_n9918_));
  NOR2_X1    g09662(.A1(new_n9918_), .A2(new_n9913_), .ZN(new_n9919_));
  AOI21_X1   g09663(.A1(new_n9673_), .A2(new_n9346_), .B(new_n9676_), .ZN(new_n9920_));
  AOI22_X1   g09664(.A1(new_n518_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n636_), .ZN(new_n9921_));
  OAI21_X1   g09665(.A1(new_n7617_), .A2(new_n917_), .B(new_n9921_), .ZN(new_n9922_));
  AOI21_X1   g09666(.A1(new_n8792_), .A2(new_n618_), .B(new_n9922_), .ZN(new_n9923_));
  XOR2_X1    g09667(.A1(new_n9923_), .A2(new_n488_), .Z(new_n9924_));
  AOI21_X1   g09668(.A1(new_n9659_), .A2(new_n9664_), .B(new_n9667_), .ZN(new_n9925_));
  OAI21_X1   g09669(.A1(new_n9920_), .A2(new_n9925_), .B(new_n9924_), .ZN(new_n9926_));
  INV_X1     g09670(.I(new_n9924_), .ZN(new_n9927_));
  INV_X1     g09671(.I(new_n9925_), .ZN(new_n9928_));
  NAND3_X1   g09672(.A1(new_n9672_), .A2(new_n9927_), .A3(new_n9928_), .ZN(new_n9929_));
  NAND3_X1   g09673(.A1(new_n9929_), .A2(new_n9926_), .A3(new_n9919_), .ZN(new_n9930_));
  INV_X1     g09674(.I(new_n9919_), .ZN(new_n9931_));
  AOI21_X1   g09675(.A1(new_n9672_), .A2(new_n9928_), .B(new_n9927_), .ZN(new_n9932_));
  NOR3_X1    g09676(.A1(new_n9920_), .A2(new_n9924_), .A3(new_n9925_), .ZN(new_n9933_));
  OAI21_X1   g09677(.A1(new_n9932_), .A2(new_n9933_), .B(new_n9931_), .ZN(new_n9934_));
  NAND3_X1   g09678(.A1(new_n9934_), .A2(new_n9930_), .A3(new_n9708_), .ZN(new_n9935_));
  NOR3_X1    g09679(.A1(new_n9932_), .A2(new_n9933_), .A3(new_n9931_), .ZN(new_n9936_));
  AOI21_X1   g09680(.A1(new_n9929_), .A2(new_n9926_), .B(new_n9919_), .ZN(new_n9937_));
  OAI21_X1   g09681(.A1(new_n9936_), .A2(new_n9937_), .B(new_n9707_), .ZN(new_n9938_));
  NAND2_X1   g09682(.A1(new_n9938_), .A2(new_n9935_), .ZN(new_n9939_));
  NOR3_X1    g09683(.A1(new_n9683_), .A2(new_n9688_), .A3(new_n9689_), .ZN(new_n9940_));
  AOI21_X1   g09684(.A1(new_n9678_), .A2(new_n9690_), .B(new_n9940_), .ZN(new_n9941_));
  INV_X1     g09685(.I(\b[54] ), .ZN(new_n9942_));
  OAI22_X1   g09686(.A1(new_n277_), .A2(new_n9942_), .B1(new_n9376_), .B2(new_n262_), .ZN(new_n9943_));
  AOI21_X1   g09687(.A1(\b[52] ), .A2(new_n283_), .B(new_n9943_), .ZN(new_n9944_));
  AOI21_X1   g09688(.A1(new_n9382_), .A2(\b[52] ), .B(\b[51] ), .ZN(new_n9945_));
  AOI21_X1   g09689(.A1(new_n9039_), .A2(\b[53] ), .B(\b[52] ), .ZN(new_n9946_));
  NOR2_X1    g09690(.A1(new_n9945_), .A2(new_n9946_), .ZN(new_n9947_));
  XNOR2_X1   g09691(.A1(\b[53] ), .A2(\b[54] ), .ZN(new_n9948_));
  NOR2_X1    g09692(.A1(new_n9947_), .A2(new_n9948_), .ZN(new_n9949_));
  XOR2_X1    g09693(.A1(\b[53] ), .A2(\b[54] ), .Z(new_n9950_));
  NOR3_X1    g09694(.A1(new_n9945_), .A2(new_n9946_), .A3(new_n9950_), .ZN(new_n9951_));
  NOR2_X1    g09695(.A1(new_n9949_), .A2(new_n9951_), .ZN(new_n9952_));
  OAI21_X1   g09696(.A1(new_n9952_), .A2(new_n279_), .B(new_n9944_), .ZN(new_n9953_));
  XOR2_X1    g09697(.A1(new_n9953_), .A2(\a[2] ), .Z(new_n9954_));
  INV_X1     g09698(.I(new_n9954_), .ZN(new_n9955_));
  NAND2_X1   g09699(.A1(new_n9941_), .A2(new_n9955_), .ZN(new_n9956_));
  AOI21_X1   g09700(.A1(new_n9364_), .A2(new_n9692_), .B(new_n9691_), .ZN(new_n9957_));
  OAI21_X1   g09701(.A1(new_n9679_), .A2(new_n9957_), .B(new_n9693_), .ZN(new_n9958_));
  NAND2_X1   g09702(.A1(new_n9958_), .A2(new_n9954_), .ZN(new_n9959_));
  AOI21_X1   g09703(.A1(new_n9959_), .A2(new_n9956_), .B(new_n9939_), .ZN(new_n9960_));
  NOR3_X1    g09704(.A1(new_n9936_), .A2(new_n9937_), .A3(new_n9707_), .ZN(new_n9961_));
  AOI21_X1   g09705(.A1(new_n9934_), .A2(new_n9930_), .B(new_n9708_), .ZN(new_n9962_));
  NOR2_X1    g09706(.A1(new_n9961_), .A2(new_n9962_), .ZN(new_n9963_));
  NOR2_X1    g09707(.A1(new_n9958_), .A2(new_n9954_), .ZN(new_n9964_));
  NOR2_X1    g09708(.A1(new_n9941_), .A2(new_n9955_), .ZN(new_n9965_));
  NOR3_X1    g09709(.A1(new_n9964_), .A2(new_n9965_), .A3(new_n9963_), .ZN(new_n9966_));
  NOR2_X1    g09710(.A1(new_n9960_), .A2(new_n9966_), .ZN(new_n9967_));
  XOR2_X1    g09711(.A1(new_n9967_), .A2(new_n9703_), .Z(\f[54] ));
  NAND2_X1   g09712(.A1(new_n283_), .A2(\b[53] ), .ZN(new_n9969_));
  AOI22_X1   g09713(.A1(new_n267_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n261_), .ZN(new_n9970_));
  INV_X1     g09714(.I(new_n9970_), .ZN(new_n9971_));
  INV_X1     g09715(.I(\b[55] ), .ZN(new_n9972_));
  OAI21_X1   g09716(.A1(new_n9945_), .A2(new_n9946_), .B(new_n9376_), .ZN(new_n9973_));
  NOR2_X1    g09717(.A1(new_n9973_), .A2(new_n9942_), .ZN(new_n9974_));
  NOR3_X1    g09718(.A1(new_n9945_), .A2(new_n9946_), .A3(new_n9376_), .ZN(new_n9975_));
  AOI21_X1   g09719(.A1(new_n9942_), .A2(new_n9975_), .B(new_n9974_), .ZN(new_n9976_));
  NOR2_X1    g09720(.A1(new_n9976_), .A2(new_n9972_), .ZN(new_n9977_));
  AND2_X2    g09721(.A1(new_n9976_), .A2(new_n9972_), .Z(new_n9978_));
  NOR2_X1    g09722(.A1(new_n9978_), .A2(new_n9977_), .ZN(new_n9979_));
  AOI21_X1   g09723(.A1(new_n9979_), .A2(new_n265_), .B(new_n9971_), .ZN(new_n9980_));
  AND3_X2    g09724(.A1(new_n9980_), .A2(\a[2] ), .A3(new_n9969_), .Z(new_n9981_));
  AOI21_X1   g09725(.A1(new_n9980_), .A2(new_n9969_), .B(\a[2] ), .ZN(new_n9982_));
  NOR2_X1    g09726(.A1(new_n9981_), .A2(new_n9982_), .ZN(new_n9983_));
  OAI21_X1   g09727(.A1(new_n9365_), .A2(new_n9366_), .B(new_n9692_), .ZN(new_n9984_));
  AOI21_X1   g09728(.A1(new_n9984_), .A2(new_n9688_), .B(new_n9679_), .ZN(new_n9985_));
  NOR3_X1    g09729(.A1(new_n9985_), .A2(new_n9940_), .A3(new_n9961_), .ZN(new_n9986_));
  INV_X1     g09730(.I(new_n9043_), .ZN(new_n9987_));
  AOI22_X1   g09731(.A1(new_n800_), .A2(\b[51] ), .B1(\b[52] ), .B2(new_n333_), .ZN(new_n9988_));
  OAI21_X1   g09732(.A1(new_n8500_), .A2(new_n392_), .B(new_n9988_), .ZN(new_n9989_));
  AOI21_X1   g09733(.A1(new_n9987_), .A2(new_n330_), .B(new_n9989_), .ZN(new_n9990_));
  XOR2_X1    g09734(.A1(new_n9990_), .A2(new_n312_), .Z(new_n9991_));
  INV_X1     g09735(.I(new_n9991_), .ZN(new_n9992_));
  AOI21_X1   g09736(.A1(new_n9919_), .A2(new_n9926_), .B(new_n9933_), .ZN(new_n9993_));
  OAI21_X1   g09737(.A1(new_n9908_), .A2(new_n9905_), .B(new_n9915_), .ZN(new_n9994_));
  OAI21_X1   g09738(.A1(new_n9327_), .A2(new_n9313_), .B(new_n9308_), .ZN(new_n9995_));
  AOI21_X1   g09739(.A1(new_n9995_), .A2(new_n9651_), .B(new_n9650_), .ZN(new_n9996_));
  OAI21_X1   g09740(.A1(new_n9996_), .A2(new_n9895_), .B(new_n9889_), .ZN(new_n9997_));
  NAND2_X1   g09741(.A1(new_n9997_), .A2(new_n9896_), .ZN(new_n9998_));
  OAI22_X1   g09742(.A1(new_n993_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n997_), .ZN(new_n9999_));
  AOI21_X1   g09743(.A1(\b[41] ), .A2(new_n1486_), .B(new_n9999_), .ZN(new_n10000_));
  OAI21_X1   g09744(.A1(new_n6785_), .A2(new_n1323_), .B(new_n10000_), .ZN(new_n10001_));
  XOR2_X1    g09745(.A1(new_n10001_), .A2(\a[14] ), .Z(new_n10002_));
  INV_X1     g09746(.I(new_n10002_), .ZN(new_n10003_));
  AOI21_X1   g09747(.A1(new_n9877_), .A2(new_n9873_), .B(new_n9869_), .ZN(new_n10004_));
  OAI22_X1   g09748(.A1(new_n1592_), .A2(new_n6284_), .B1(new_n5761_), .B2(new_n1505_), .ZN(new_n10005_));
  AOI21_X1   g09749(.A1(\b[38] ), .A2(new_n1584_), .B(new_n10005_), .ZN(new_n10006_));
  OAI21_X1   g09750(.A1(new_n8195_), .A2(new_n1732_), .B(new_n10006_), .ZN(new_n10007_));
  XOR2_X1    g09751(.A1(new_n10007_), .A2(\a[17] ), .Z(new_n10008_));
  OAI21_X1   g09752(.A1(new_n9860_), .A2(new_n9858_), .B(new_n9850_), .ZN(new_n10009_));
  OAI22_X1   g09753(.A1(new_n1751_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n1754_), .ZN(new_n10010_));
  AOI21_X1   g09754(.A1(\b[35] ), .A2(new_n1939_), .B(new_n10010_), .ZN(new_n10011_));
  OAI21_X1   g09755(.A1(new_n5322_), .A2(new_n1757_), .B(new_n10011_), .ZN(new_n10012_));
  XOR2_X1    g09756(.A1(new_n10012_), .A2(\a[20] ), .Z(new_n10013_));
  AOI21_X1   g09757(.A1(new_n9841_), .A2(new_n9836_), .B(new_n9832_), .ZN(new_n10014_));
  AOI22_X1   g09758(.A1(new_n2202_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n2205_), .ZN(new_n10015_));
  OAI21_X1   g09759(.A1(new_n4023_), .A2(new_n2370_), .B(new_n10015_), .ZN(new_n10016_));
  AOI21_X1   g09760(.A1(new_n5103_), .A2(new_n2208_), .B(new_n10016_), .ZN(new_n10017_));
  XOR2_X1    g09761(.A1(new_n10017_), .A2(new_n2200_), .Z(new_n10018_));
  OAI21_X1   g09762(.A1(new_n9823_), .A2(new_n9822_), .B(new_n9813_), .ZN(new_n10019_));
  AOI22_X1   g09763(.A1(new_n2716_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n2719_), .ZN(new_n10020_));
  OAI21_X1   g09764(.A1(new_n3592_), .A2(new_n2924_), .B(new_n10020_), .ZN(new_n10021_));
  AOI21_X1   g09765(.A1(new_n3796_), .A2(new_n2722_), .B(new_n10021_), .ZN(new_n10022_));
  XOR2_X1    g09766(.A1(new_n10022_), .A2(new_n2714_), .Z(new_n10023_));
  NOR3_X1    g09767(.A1(new_n9586_), .A2(new_n9587_), .A3(new_n9807_), .ZN(new_n10024_));
  OAI21_X1   g09768(.A1(new_n9569_), .A2(new_n9572_), .B(new_n9798_), .ZN(new_n10025_));
  NOR2_X1    g09769(.A1(new_n10025_), .A2(new_n9794_), .ZN(new_n10026_));
  OR2_X2     g09770(.A1(new_n9785_), .A2(new_n9789_), .Z(new_n10027_));
  AOI21_X1   g09771(.A1(new_n10025_), .A2(new_n9794_), .B(new_n10027_), .ZN(new_n10028_));
  AOI22_X1   g09772(.A1(new_n4918_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n4921_), .ZN(new_n10029_));
  OAI21_X1   g09773(.A1(new_n1860_), .A2(new_n6099_), .B(new_n10029_), .ZN(new_n10030_));
  AOI21_X1   g09774(.A1(new_n2659_), .A2(new_n4699_), .B(new_n10030_), .ZN(new_n10031_));
  XOR2_X1    g09775(.A1(new_n10031_), .A2(new_n4446_), .Z(new_n10032_));
  NOR3_X1    g09776(.A1(new_n9774_), .A2(new_n9771_), .A3(new_n9715_), .ZN(new_n10033_));
  AOI21_X1   g09777(.A1(new_n9711_), .A2(new_n9775_), .B(new_n10033_), .ZN(new_n10034_));
  AOI21_X1   g09778(.A1(new_n9760_), .A2(new_n9767_), .B(new_n9768_), .ZN(new_n10035_));
  NAND2_X1   g09779(.A1(new_n9754_), .A2(new_n9747_), .ZN(new_n10036_));
  NAND2_X1   g09780(.A1(new_n10036_), .A2(new_n9758_), .ZN(new_n10037_));
  NAND2_X1   g09781(.A1(new_n10035_), .A2(new_n10037_), .ZN(new_n10038_));
  NOR2_X1    g09782(.A1(new_n10035_), .A2(new_n10037_), .ZN(new_n10039_));
  INV_X1     g09783(.I(new_n10039_), .ZN(new_n10040_));
  AOI22_X1   g09784(.A1(new_n6108_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n6111_), .ZN(new_n10041_));
  OAI21_X1   g09785(.A1(new_n1093_), .A2(new_n7708_), .B(new_n10041_), .ZN(new_n10042_));
  AOI21_X1   g09786(.A1(new_n1701_), .A2(new_n6105_), .B(new_n10042_), .ZN(new_n10043_));
  XOR2_X1    g09787(.A1(new_n10043_), .A2(new_n5849_), .Z(new_n10044_));
  NOR2_X1    g09788(.A1(new_n9740_), .A2(new_n9744_), .ZN(new_n10045_));
  AOI21_X1   g09789(.A1(new_n9740_), .A2(new_n9744_), .B(new_n9717_), .ZN(new_n10046_));
  NOR2_X1    g09790(.A1(new_n10046_), .A2(new_n10045_), .ZN(new_n10047_));
  INV_X1     g09791(.I(new_n10047_), .ZN(new_n10048_));
  NOR2_X1    g09792(.A1(new_n9738_), .A2(new_n9719_), .ZN(new_n10049_));
  NOR2_X1    g09793(.A1(new_n10049_), .A2(new_n9737_), .ZN(new_n10050_));
  NAND2_X1   g09794(.A1(new_n9734_), .A2(new_n9479_), .ZN(new_n10051_));
  NAND2_X1   g09795(.A1(new_n10051_), .A2(new_n9731_), .ZN(new_n10052_));
  AOI22_X1   g09796(.A1(new_n9125_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n9123_), .ZN(new_n10053_));
  OAI21_X1   g09797(.A1(new_n276_), .A2(new_n9470_), .B(new_n10053_), .ZN(new_n10054_));
  AOI21_X1   g09798(.A1(new_n1725_), .A2(new_n9129_), .B(new_n10054_), .ZN(new_n10055_));
  XOR2_X1    g09799(.A1(new_n10055_), .A2(\a[53] ), .Z(new_n10056_));
  INV_X1     g09800(.I(\a[56] ), .ZN(new_n10057_));
  INV_X1     g09801(.I(\a[54] ), .ZN(new_n10058_));
  NAND3_X1   g09802(.A1(new_n9133_), .A2(new_n10058_), .A3(\a[55] ), .ZN(new_n10059_));
  INV_X1     g09803(.I(\a[55] ), .ZN(new_n10060_));
  NAND3_X1   g09804(.A1(new_n10060_), .A2(\a[53] ), .A3(\a[54] ), .ZN(new_n10061_));
  NAND2_X1   g09805(.A1(new_n10059_), .A2(new_n10061_), .ZN(new_n10062_));
  XOR2_X1    g09806(.A1(\a[55] ), .A2(\a[56] ), .Z(new_n10063_));
  NOR2_X1    g09807(.A1(new_n9729_), .A2(new_n10063_), .ZN(new_n10064_));
  AOI22_X1   g09808(.A1(new_n10064_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n10062_), .ZN(new_n10065_));
  XOR2_X1    g09809(.A1(\a[55] ), .A2(\a[56] ), .Z(new_n10066_));
  INV_X1     g09810(.I(new_n10066_), .ZN(new_n10067_));
  NOR2_X1    g09811(.A1(new_n10067_), .A2(new_n9729_), .ZN(new_n10068_));
  INV_X1     g09812(.I(new_n10068_), .ZN(new_n10069_));
  OAI21_X1   g09813(.A1(new_n313_), .A2(new_n10069_), .B(new_n10065_), .ZN(new_n10070_));
  OR3_X2     g09814(.A1(new_n10070_), .A2(new_n10057_), .A3(new_n9730_), .Z(new_n10071_));
  XOR2_X1    g09815(.A1(new_n10070_), .A2(new_n10057_), .Z(new_n10072_));
  NAND2_X1   g09816(.A1(new_n9733_), .A2(\a[56] ), .ZN(new_n10073_));
  NAND2_X1   g09817(.A1(new_n10072_), .A2(new_n10073_), .ZN(new_n10074_));
  NAND2_X1   g09818(.A1(new_n10074_), .A2(new_n10071_), .ZN(new_n10075_));
  OR2_X2     g09819(.A1(new_n10075_), .A2(new_n10056_), .Z(new_n10076_));
  NAND2_X1   g09820(.A1(new_n10075_), .A2(new_n10056_), .ZN(new_n10077_));
  NAND2_X1   g09821(.A1(new_n10076_), .A2(new_n10077_), .ZN(new_n10078_));
  XOR2_X1    g09822(.A1(new_n10078_), .A2(new_n10052_), .Z(new_n10079_));
  OAI22_X1   g09823(.A1(new_n9461_), .A2(new_n471_), .B1(new_n438_), .B2(new_n9462_), .ZN(new_n10080_));
  AOI21_X1   g09824(.A1(\b[5] ), .A2(new_n8575_), .B(new_n10080_), .ZN(new_n10081_));
  OAI21_X1   g09825(.A1(new_n485_), .A2(new_n9460_), .B(new_n10081_), .ZN(new_n10082_));
  XOR2_X1    g09826(.A1(new_n10082_), .A2(\a[50] ), .Z(new_n10083_));
  INV_X1     g09827(.I(new_n10083_), .ZN(new_n10084_));
  NAND2_X1   g09828(.A1(new_n10079_), .A2(new_n10084_), .ZN(new_n10085_));
  INV_X1     g09829(.I(new_n10079_), .ZN(new_n10086_));
  NAND2_X1   g09830(.A1(new_n10086_), .A2(new_n10083_), .ZN(new_n10087_));
  NAND2_X1   g09831(.A1(new_n10087_), .A2(new_n10085_), .ZN(new_n10088_));
  XOR2_X1    g09832(.A1(new_n10088_), .A2(new_n10050_), .Z(new_n10089_));
  AOI22_X1   g09833(.A1(new_n7403_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n7408_), .ZN(new_n10090_));
  OAI21_X1   g09834(.A1(new_n577_), .A2(new_n9488_), .B(new_n10090_), .ZN(new_n10091_));
  AOI21_X1   g09835(.A1(new_n1059_), .A2(new_n7414_), .B(new_n10091_), .ZN(new_n10092_));
  XOR2_X1    g09836(.A1(new_n10092_), .A2(new_n7410_), .Z(new_n10093_));
  INV_X1     g09837(.I(new_n10093_), .ZN(new_n10094_));
  NAND2_X1   g09838(.A1(new_n10089_), .A2(new_n10094_), .ZN(new_n10095_));
  XNOR2_X1   g09839(.A1(new_n10088_), .A2(new_n10050_), .ZN(new_n10096_));
  NAND2_X1   g09840(.A1(new_n10096_), .A2(new_n10093_), .ZN(new_n10097_));
  NAND3_X1   g09841(.A1(new_n10048_), .A2(new_n10095_), .A3(new_n10097_), .ZN(new_n10098_));
  NOR2_X1    g09842(.A1(new_n10096_), .A2(new_n10093_), .ZN(new_n10099_));
  NOR2_X1    g09843(.A1(new_n10089_), .A2(new_n10094_), .ZN(new_n10100_));
  OAI21_X1   g09844(.A1(new_n10099_), .A2(new_n10100_), .B(new_n10047_), .ZN(new_n10101_));
  OAI22_X1   g09845(.A1(new_n7730_), .A2(new_n1070_), .B1(new_n941_), .B2(new_n7731_), .ZN(new_n10102_));
  AOI21_X1   g09846(.A1(\b[11] ), .A2(new_n6887_), .B(new_n10102_), .ZN(new_n10103_));
  OAI21_X1   g09847(.A1(new_n1082_), .A2(new_n7728_), .B(new_n10103_), .ZN(new_n10104_));
  XOR2_X1    g09848(.A1(new_n10104_), .A2(\a[44] ), .Z(new_n10105_));
  INV_X1     g09849(.I(new_n10105_), .ZN(new_n10106_));
  NAND3_X1   g09850(.A1(new_n10098_), .A2(new_n10101_), .A3(new_n10106_), .ZN(new_n10107_));
  NAND2_X1   g09851(.A1(new_n10098_), .A2(new_n10101_), .ZN(new_n10108_));
  NAND2_X1   g09852(.A1(new_n10108_), .A2(new_n10105_), .ZN(new_n10109_));
  NAND2_X1   g09853(.A1(new_n10109_), .A2(new_n10107_), .ZN(new_n10110_));
  XNOR2_X1   g09854(.A1(new_n10110_), .A2(new_n10044_), .ZN(new_n10111_));
  NAND3_X1   g09855(.A1(new_n10040_), .A2(new_n10038_), .A3(new_n10111_), .ZN(new_n10112_));
  INV_X1     g09856(.I(new_n10038_), .ZN(new_n10113_));
  INV_X1     g09857(.I(new_n10111_), .ZN(new_n10114_));
  OAI21_X1   g09858(.A1(new_n10113_), .A2(new_n10039_), .B(new_n10114_), .ZN(new_n10115_));
  AOI22_X1   g09859(.A1(new_n5155_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n5160_), .ZN(new_n10116_));
  OAI21_X1   g09860(.A1(new_n1432_), .A2(new_n6877_), .B(new_n10116_), .ZN(new_n10117_));
  AOI21_X1   g09861(.A1(new_n1695_), .A2(new_n5166_), .B(new_n10117_), .ZN(new_n10118_));
  XOR2_X1    g09862(.A1(new_n10118_), .A2(new_n5162_), .Z(new_n10119_));
  INV_X1     g09863(.I(new_n10119_), .ZN(new_n10120_));
  NAND3_X1   g09864(.A1(new_n10115_), .A2(new_n10112_), .A3(new_n10120_), .ZN(new_n10121_));
  NOR3_X1    g09865(.A1(new_n10113_), .A2(new_n10039_), .A3(new_n10114_), .ZN(new_n10122_));
  AOI21_X1   g09866(.A1(new_n10040_), .A2(new_n10038_), .B(new_n10111_), .ZN(new_n10123_));
  OAI21_X1   g09867(.A1(new_n10123_), .A2(new_n10122_), .B(new_n10119_), .ZN(new_n10124_));
  NAND3_X1   g09868(.A1(new_n10124_), .A2(new_n10121_), .A3(new_n10034_), .ZN(new_n10125_));
  AOI21_X1   g09869(.A1(new_n10124_), .A2(new_n10121_), .B(new_n10034_), .ZN(new_n10126_));
  INV_X1     g09870(.I(new_n10126_), .ZN(new_n10127_));
  AOI21_X1   g09871(.A1(new_n10127_), .A2(new_n10125_), .B(new_n10032_), .ZN(new_n10128_));
  INV_X1     g09872(.I(new_n10032_), .ZN(new_n10129_));
  AOI21_X1   g09873(.A1(new_n9772_), .A2(new_n9770_), .B(new_n9716_), .ZN(new_n10130_));
  OAI21_X1   g09874(.A1(new_n9710_), .A2(new_n10130_), .B(new_n9773_), .ZN(new_n10131_));
  INV_X1     g09875(.I(new_n10121_), .ZN(new_n10132_));
  AOI21_X1   g09876(.A1(new_n10115_), .A2(new_n10112_), .B(new_n10120_), .ZN(new_n10133_));
  NOR3_X1    g09877(.A1(new_n10132_), .A2(new_n10133_), .A3(new_n10131_), .ZN(new_n10134_));
  NOR3_X1    g09878(.A1(new_n10134_), .A2(new_n10126_), .A3(new_n10129_), .ZN(new_n10135_));
  NOR2_X1    g09879(.A1(new_n10128_), .A2(new_n10135_), .ZN(new_n10136_));
  NOR3_X1    g09880(.A1(new_n10028_), .A2(new_n10026_), .A3(new_n10136_), .ZN(new_n10137_));
  AOI21_X1   g09881(.A1(new_n9582_), .A2(new_n9567_), .B(new_n9795_), .ZN(new_n10138_));
  OAI21_X1   g09882(.A1(new_n10138_), .A2(new_n9797_), .B(new_n9790_), .ZN(new_n10139_));
  INV_X1     g09883(.I(new_n10136_), .ZN(new_n10140_));
  AOI21_X1   g09884(.A1(new_n10139_), .A2(new_n9799_), .B(new_n10140_), .ZN(new_n10141_));
  AOI21_X1   g09885(.A1(new_n9786_), .A2(new_n9787_), .B(new_n9784_), .ZN(new_n10142_));
  OAI22_X1   g09886(.A1(new_n2495_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n2646_), .ZN(new_n10143_));
  AOI21_X1   g09887(.A1(\b[23] ), .A2(new_n4053_), .B(new_n10143_), .ZN(new_n10144_));
  OAI21_X1   g09888(.A1(new_n2655_), .A2(new_n4727_), .B(new_n10144_), .ZN(new_n10145_));
  XOR2_X1    g09889(.A1(new_n10145_), .A2(\a[32] ), .Z(new_n10146_));
  XOR2_X1    g09890(.A1(new_n10142_), .A2(new_n10146_), .Z(new_n10147_));
  INV_X1     g09891(.I(new_n10147_), .ZN(new_n10148_));
  NOR3_X1    g09892(.A1(new_n10137_), .A2(new_n10141_), .A3(new_n10148_), .ZN(new_n10149_));
  NAND3_X1   g09893(.A1(new_n10139_), .A2(new_n9799_), .A3(new_n10140_), .ZN(new_n10150_));
  OAI21_X1   g09894(.A1(new_n10028_), .A2(new_n10026_), .B(new_n10136_), .ZN(new_n10151_));
  AOI21_X1   g09895(.A1(new_n10151_), .A2(new_n10150_), .B(new_n10147_), .ZN(new_n10152_));
  AOI22_X1   g09896(.A1(new_n3267_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n3270_), .ZN(new_n10153_));
  OAI21_X1   g09897(.A1(new_n3006_), .A2(new_n3475_), .B(new_n10153_), .ZN(new_n10154_));
  AOI21_X1   g09898(.A1(new_n3807_), .A2(new_n3273_), .B(new_n10154_), .ZN(new_n10155_));
  XOR2_X1    g09899(.A1(new_n10155_), .A2(new_n3264_), .Z(new_n10156_));
  NOR3_X1    g09900(.A1(new_n10149_), .A2(new_n10152_), .A3(new_n10156_), .ZN(new_n10157_));
  NAND3_X1   g09901(.A1(new_n10151_), .A2(new_n10150_), .A3(new_n10147_), .ZN(new_n10158_));
  OAI21_X1   g09902(.A1(new_n10137_), .A2(new_n10141_), .B(new_n10148_), .ZN(new_n10159_));
  INV_X1     g09903(.I(new_n10156_), .ZN(new_n10160_));
  AOI21_X1   g09904(.A1(new_n10159_), .A2(new_n10158_), .B(new_n10160_), .ZN(new_n10161_));
  INV_X1     g09905(.I(new_n9802_), .ZN(new_n10162_));
  NAND2_X1   g09906(.A1(new_n10162_), .A2(new_n9800_), .ZN(new_n10163_));
  OAI21_X1   g09907(.A1(new_n9596_), .A2(new_n9585_), .B(new_n9579_), .ZN(new_n10164_));
  AOI21_X1   g09908(.A1(new_n10164_), .A2(new_n9807_), .B(new_n10163_), .ZN(new_n10165_));
  NOR4_X1    g09909(.A1(new_n10165_), .A2(new_n10157_), .A3(new_n10161_), .A4(new_n10024_), .ZN(new_n10166_));
  NAND3_X1   g09910(.A1(new_n10159_), .A2(new_n10158_), .A3(new_n10160_), .ZN(new_n10167_));
  OAI21_X1   g09911(.A1(new_n10149_), .A2(new_n10152_), .B(new_n10156_), .ZN(new_n10168_));
  AOI21_X1   g09912(.A1(new_n9593_), .A2(new_n9589_), .B(new_n9587_), .ZN(new_n10169_));
  OAI21_X1   g09913(.A1(new_n10169_), .A2(new_n9809_), .B(new_n9803_), .ZN(new_n10170_));
  AOI22_X1   g09914(.A1(new_n10170_), .A2(new_n9810_), .B1(new_n10168_), .B2(new_n10167_), .ZN(new_n10171_));
  OAI21_X1   g09915(.A1(new_n10166_), .A2(new_n10171_), .B(new_n10023_), .ZN(new_n10172_));
  INV_X1     g09916(.I(new_n10023_), .ZN(new_n10173_));
  NAND4_X1   g09917(.A1(new_n10170_), .A2(new_n10168_), .A3(new_n9810_), .A4(new_n10167_), .ZN(new_n10174_));
  OAI22_X1   g09918(.A1(new_n10165_), .A2(new_n10024_), .B1(new_n10157_), .B2(new_n10161_), .ZN(new_n10175_));
  NAND3_X1   g09919(.A1(new_n10175_), .A2(new_n10174_), .A3(new_n10173_), .ZN(new_n10176_));
  NAND2_X1   g09920(.A1(new_n10172_), .A2(new_n10176_), .ZN(new_n10177_));
  NAND3_X1   g09921(.A1(new_n10019_), .A2(new_n10177_), .A3(new_n9824_), .ZN(new_n10178_));
  AOI21_X1   g09922(.A1(new_n9820_), .A2(new_n9817_), .B(new_n9828_), .ZN(new_n10179_));
  AOI21_X1   g09923(.A1(new_n10175_), .A2(new_n10174_), .B(new_n10173_), .ZN(new_n10180_));
  NOR3_X1    g09924(.A1(new_n10166_), .A2(new_n10171_), .A3(new_n10023_), .ZN(new_n10181_));
  NOR2_X1    g09925(.A1(new_n10181_), .A2(new_n10180_), .ZN(new_n10182_));
  OAI21_X1   g09926(.A1(new_n10179_), .A2(new_n9830_), .B(new_n10182_), .ZN(new_n10183_));
  NAND3_X1   g09927(.A1(new_n10183_), .A2(new_n10178_), .A3(new_n10018_), .ZN(new_n10184_));
  INV_X1     g09928(.I(new_n10018_), .ZN(new_n10185_));
  NOR3_X1    g09929(.A1(new_n10179_), .A2(new_n9830_), .A3(new_n10182_), .ZN(new_n10186_));
  AOI21_X1   g09930(.A1(new_n10019_), .A2(new_n9824_), .B(new_n10177_), .ZN(new_n10187_));
  OAI21_X1   g09931(.A1(new_n10186_), .A2(new_n10187_), .B(new_n10185_), .ZN(new_n10188_));
  NAND2_X1   g09932(.A1(new_n10188_), .A2(new_n10184_), .ZN(new_n10189_));
  NOR3_X1    g09933(.A1(new_n10014_), .A2(new_n9842_), .A3(new_n10189_), .ZN(new_n10190_));
  OAI21_X1   g09934(.A1(new_n9838_), .A2(new_n9837_), .B(new_n9846_), .ZN(new_n10191_));
  NOR3_X1    g09935(.A1(new_n10186_), .A2(new_n10187_), .A3(new_n10185_), .ZN(new_n10192_));
  AOI21_X1   g09936(.A1(new_n10183_), .A2(new_n10178_), .B(new_n10018_), .ZN(new_n10193_));
  NOR2_X1    g09937(.A1(new_n10192_), .A2(new_n10193_), .ZN(new_n10194_));
  AOI21_X1   g09938(.A1(new_n10191_), .A2(new_n9848_), .B(new_n10194_), .ZN(new_n10195_));
  OAI21_X1   g09939(.A1(new_n10190_), .A2(new_n10195_), .B(new_n10013_), .ZN(new_n10196_));
  INV_X1     g09940(.I(new_n10013_), .ZN(new_n10197_));
  NAND3_X1   g09941(.A1(new_n10191_), .A2(new_n10194_), .A3(new_n9848_), .ZN(new_n10198_));
  OAI21_X1   g09942(.A1(new_n10014_), .A2(new_n9842_), .B(new_n10189_), .ZN(new_n10199_));
  NAND3_X1   g09943(.A1(new_n10199_), .A2(new_n10198_), .A3(new_n10197_), .ZN(new_n10200_));
  NAND2_X1   g09944(.A1(new_n10196_), .A2(new_n10200_), .ZN(new_n10201_));
  NAND3_X1   g09945(.A1(new_n10009_), .A2(new_n9861_), .A3(new_n10201_), .ZN(new_n10202_));
  AOI21_X1   g09946(.A1(new_n9856_), .A2(new_n9854_), .B(new_n9865_), .ZN(new_n10203_));
  AOI21_X1   g09947(.A1(new_n10199_), .A2(new_n10198_), .B(new_n10197_), .ZN(new_n10204_));
  NOR3_X1    g09948(.A1(new_n10190_), .A2(new_n10195_), .A3(new_n10013_), .ZN(new_n10205_));
  NOR2_X1    g09949(.A1(new_n10205_), .A2(new_n10204_), .ZN(new_n10206_));
  OAI21_X1   g09950(.A1(new_n10203_), .A2(new_n9867_), .B(new_n10206_), .ZN(new_n10207_));
  NAND3_X1   g09951(.A1(new_n10202_), .A2(new_n10207_), .A3(new_n10008_), .ZN(new_n10208_));
  INV_X1     g09952(.I(new_n10008_), .ZN(new_n10209_));
  NOR3_X1    g09953(.A1(new_n10203_), .A2(new_n9867_), .A3(new_n10206_), .ZN(new_n10210_));
  AOI21_X1   g09954(.A1(new_n10009_), .A2(new_n9861_), .B(new_n10201_), .ZN(new_n10211_));
  OAI21_X1   g09955(.A1(new_n10211_), .A2(new_n10210_), .B(new_n10209_), .ZN(new_n10212_));
  NAND2_X1   g09956(.A1(new_n10212_), .A2(new_n10208_), .ZN(new_n10213_));
  NOR3_X1    g09957(.A1(new_n10004_), .A2(new_n9878_), .A3(new_n10213_), .ZN(new_n10214_));
  OAI21_X1   g09958(.A1(new_n9886_), .A2(new_n9883_), .B(new_n9882_), .ZN(new_n10215_));
  NOR3_X1    g09959(.A1(new_n10211_), .A2(new_n10210_), .A3(new_n10209_), .ZN(new_n10216_));
  AOI21_X1   g09960(.A1(new_n10202_), .A2(new_n10207_), .B(new_n10008_), .ZN(new_n10217_));
  NOR2_X1    g09961(.A1(new_n10217_), .A2(new_n10216_), .ZN(new_n10218_));
  AOI21_X1   g09962(.A1(new_n10215_), .A2(new_n9887_), .B(new_n10218_), .ZN(new_n10219_));
  OAI21_X1   g09963(.A1(new_n10214_), .A2(new_n10219_), .B(new_n10003_), .ZN(new_n10220_));
  NOR3_X1    g09964(.A1(new_n10214_), .A2(new_n10219_), .A3(new_n10003_), .ZN(new_n10221_));
  INV_X1     g09965(.I(new_n10221_), .ZN(new_n10222_));
  NAND2_X1   g09966(.A1(new_n10222_), .A2(new_n10220_), .ZN(new_n10223_));
  NOR2_X1    g09967(.A1(new_n9998_), .A2(new_n10223_), .ZN(new_n10224_));
  NOR3_X1    g09968(.A1(new_n9648_), .A2(new_n9650_), .A3(new_n9893_), .ZN(new_n10225_));
  AOI21_X1   g09969(.A1(new_n9889_), .A2(new_n9894_), .B(new_n10225_), .ZN(new_n10226_));
  NAND3_X1   g09970(.A1(new_n10215_), .A2(new_n10218_), .A3(new_n9887_), .ZN(new_n10227_));
  INV_X1     g09971(.I(new_n10219_), .ZN(new_n10228_));
  AOI21_X1   g09972(.A1(new_n10228_), .A2(new_n10227_), .B(new_n10002_), .ZN(new_n10229_));
  NOR2_X1    g09973(.A1(new_n10229_), .A2(new_n10221_), .ZN(new_n10230_));
  NOR2_X1    g09974(.A1(new_n10226_), .A2(new_n10230_), .ZN(new_n10231_));
  OAI22_X1   g09975(.A1(new_n713_), .A2(new_n7617_), .B1(new_n7096_), .B2(new_n717_), .ZN(new_n10232_));
  AOI21_X1   g09976(.A1(\b[44] ), .A2(new_n1126_), .B(new_n10232_), .ZN(new_n10233_));
  OAI21_X1   g09977(.A1(new_n7627_), .A2(new_n986_), .B(new_n10233_), .ZN(new_n10234_));
  XOR2_X1    g09978(.A1(new_n10234_), .A2(\a[11] ), .Z(new_n10235_));
  INV_X1     g09979(.I(new_n10235_), .ZN(new_n10236_));
  OAI21_X1   g09980(.A1(new_n10224_), .A2(new_n10231_), .B(new_n10236_), .ZN(new_n10237_));
  NAND2_X1   g09981(.A1(new_n10226_), .A2(new_n10230_), .ZN(new_n10238_));
  NAND2_X1   g09982(.A1(new_n9998_), .A2(new_n10223_), .ZN(new_n10239_));
  NAND3_X1   g09983(.A1(new_n10239_), .A2(new_n10238_), .A3(new_n10235_), .ZN(new_n10240_));
  NAND2_X1   g09984(.A1(new_n10237_), .A2(new_n10240_), .ZN(new_n10241_));
  AOI21_X1   g09985(.A1(new_n9994_), .A2(new_n9917_), .B(new_n10241_), .ZN(new_n10242_));
  AOI21_X1   g09986(.A1(new_n9911_), .A2(new_n9904_), .B(new_n9900_), .ZN(new_n10243_));
  AOI21_X1   g09987(.A1(new_n10239_), .A2(new_n10238_), .B(new_n10235_), .ZN(new_n10244_));
  NOR3_X1    g09988(.A1(new_n10224_), .A2(new_n10231_), .A3(new_n10236_), .ZN(new_n10245_));
  NOR2_X1    g09989(.A1(new_n10245_), .A2(new_n10244_), .ZN(new_n10246_));
  NOR3_X1    g09990(.A1(new_n10246_), .A2(new_n10243_), .A3(new_n9912_), .ZN(new_n10247_));
  OAI22_X1   g09991(.A1(new_n610_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n612_), .ZN(new_n10248_));
  AOI21_X1   g09992(.A1(\b[47] ), .A2(new_n826_), .B(new_n10248_), .ZN(new_n10249_));
  OAI21_X1   g09993(.A1(new_n9050_), .A2(new_n624_), .B(new_n10249_), .ZN(new_n10250_));
  XOR2_X1    g09994(.A1(new_n10250_), .A2(\a[8] ), .Z(new_n10251_));
  OAI21_X1   g09995(.A1(new_n10242_), .A2(new_n10247_), .B(new_n10251_), .ZN(new_n10252_));
  OAI21_X1   g09996(.A1(new_n9912_), .A2(new_n10243_), .B(new_n10246_), .ZN(new_n10253_));
  NAND3_X1   g09997(.A1(new_n10241_), .A2(new_n9994_), .A3(new_n9917_), .ZN(new_n10254_));
  INV_X1     g09998(.I(new_n10251_), .ZN(new_n10255_));
  NAND3_X1   g09999(.A1(new_n10253_), .A2(new_n10254_), .A3(new_n10255_), .ZN(new_n10256_));
  NAND2_X1   g10000(.A1(new_n10252_), .A2(new_n10256_), .ZN(new_n10257_));
  NOR2_X1    g10001(.A1(new_n9993_), .A2(new_n10257_), .ZN(new_n10258_));
  OAI21_X1   g10002(.A1(new_n9931_), .A2(new_n9932_), .B(new_n9929_), .ZN(new_n10259_));
  AOI21_X1   g10003(.A1(new_n10253_), .A2(new_n10254_), .B(new_n10255_), .ZN(new_n10260_));
  NOR3_X1    g10004(.A1(new_n10242_), .A2(new_n10247_), .A3(new_n10251_), .ZN(new_n10261_));
  NOR2_X1    g10005(.A1(new_n10260_), .A2(new_n10261_), .ZN(new_n10262_));
  NOR2_X1    g10006(.A1(new_n10259_), .A2(new_n10262_), .ZN(new_n10263_));
  NOR3_X1    g10007(.A1(new_n10263_), .A2(new_n10258_), .A3(new_n9992_), .ZN(new_n10264_));
  NOR2_X1    g10008(.A1(new_n9932_), .A2(new_n9931_), .ZN(new_n10265_));
  OAI21_X1   g10009(.A1(new_n10265_), .A2(new_n9933_), .B(new_n10262_), .ZN(new_n10266_));
  NAND2_X1   g10010(.A1(new_n9926_), .A2(new_n9919_), .ZN(new_n10267_));
  NAND3_X1   g10011(.A1(new_n10267_), .A2(new_n10257_), .A3(new_n9929_), .ZN(new_n10268_));
  AOI21_X1   g10012(.A1(new_n10266_), .A2(new_n10268_), .B(new_n9991_), .ZN(new_n10269_));
  OAI22_X1   g10013(.A1(new_n9986_), .A2(new_n9962_), .B1(new_n10264_), .B2(new_n10269_), .ZN(new_n10270_));
  AOI21_X1   g10014(.A1(new_n9941_), .A2(new_n9935_), .B(new_n9962_), .ZN(new_n10271_));
  NOR2_X1    g10015(.A1(new_n10264_), .A2(new_n10269_), .ZN(new_n10272_));
  NAND2_X1   g10016(.A1(new_n10271_), .A2(new_n10272_), .ZN(new_n10273_));
  AOI21_X1   g10017(.A1(new_n10273_), .A2(new_n10270_), .B(new_n9983_), .ZN(new_n10274_));
  INV_X1     g10018(.I(new_n9983_), .ZN(new_n10275_));
  NAND2_X1   g10019(.A1(new_n9680_), .A2(new_n9020_), .ZN(new_n10276_));
  NAND2_X1   g10020(.A1(new_n9682_), .A2(new_n9681_), .ZN(new_n10277_));
  AOI21_X1   g10021(.A1(new_n10276_), .A2(new_n10277_), .B(new_n9689_), .ZN(new_n10278_));
  OAI21_X1   g10022(.A1(new_n10278_), .A2(new_n9691_), .B(new_n9678_), .ZN(new_n10279_));
  NAND3_X1   g10023(.A1(new_n10279_), .A2(new_n9693_), .A3(new_n9935_), .ZN(new_n10280_));
  NAND3_X1   g10024(.A1(new_n10266_), .A2(new_n10268_), .A3(new_n9991_), .ZN(new_n10281_));
  OAI21_X1   g10025(.A1(new_n10263_), .A2(new_n10258_), .B(new_n9992_), .ZN(new_n10282_));
  AOI22_X1   g10026(.A1(new_n10280_), .A2(new_n9938_), .B1(new_n10281_), .B2(new_n10282_), .ZN(new_n10283_));
  OAI21_X1   g10027(.A1(new_n9958_), .A2(new_n9961_), .B(new_n9938_), .ZN(new_n10284_));
  NAND2_X1   g10028(.A1(new_n10282_), .A2(new_n10281_), .ZN(new_n10285_));
  NOR2_X1    g10029(.A1(new_n10284_), .A2(new_n10285_), .ZN(new_n10286_));
  NOR3_X1    g10030(.A1(new_n10286_), .A2(new_n10275_), .A3(new_n10283_), .ZN(new_n10287_));
  NOR2_X1    g10031(.A1(new_n10287_), .A2(new_n10274_), .ZN(new_n10288_));
  NAND2_X1   g10032(.A1(new_n9941_), .A2(new_n9939_), .ZN(new_n10289_));
  NAND2_X1   g10033(.A1(new_n9958_), .A2(new_n9963_), .ZN(new_n10290_));
  AOI21_X1   g10034(.A1(new_n10290_), .A2(new_n10289_), .B(new_n9955_), .ZN(new_n10291_));
  AOI21_X1   g10035(.A1(new_n9967_), .A2(new_n9703_), .B(new_n10291_), .ZN(new_n10292_));
  XOR2_X1    g10036(.A1(new_n10292_), .A2(new_n10288_), .Z(\f[55] ));
  OAI21_X1   g10037(.A1(new_n10286_), .A2(new_n10283_), .B(new_n10275_), .ZN(new_n10294_));
  NAND3_X1   g10038(.A1(new_n10273_), .A2(new_n10270_), .A3(new_n9983_), .ZN(new_n10295_));
  NAND2_X1   g10039(.A1(new_n10294_), .A2(new_n10295_), .ZN(new_n10296_));
  INV_X1     g10040(.I(new_n9371_), .ZN(new_n10297_));
  OAI21_X1   g10041(.A1(new_n9031_), .A2(new_n10297_), .B(new_n9370_), .ZN(new_n10298_));
  NOR3_X1    g10042(.A1(new_n9695_), .A2(new_n9388_), .A3(new_n9696_), .ZN(new_n10299_));
  OAI21_X1   g10043(.A1(new_n10298_), .A2(new_n10299_), .B(new_n9697_), .ZN(new_n10300_));
  OAI21_X1   g10044(.A1(new_n9964_), .A2(new_n9965_), .B(new_n9963_), .ZN(new_n10301_));
  NAND3_X1   g10045(.A1(new_n9959_), .A2(new_n9956_), .A3(new_n9939_), .ZN(new_n10302_));
  NAND2_X1   g10046(.A1(new_n10301_), .A2(new_n10302_), .ZN(new_n10303_));
  INV_X1     g10047(.I(new_n10291_), .ZN(new_n10304_));
  OAI21_X1   g10048(.A1(new_n10300_), .A2(new_n10303_), .B(new_n10304_), .ZN(new_n10305_));
  NOR3_X1    g10049(.A1(new_n10286_), .A2(new_n9983_), .A3(new_n10283_), .ZN(new_n10306_));
  AOI21_X1   g10050(.A1(new_n10305_), .A2(new_n10296_), .B(new_n10306_), .ZN(new_n10307_));
  INV_X1     g10051(.I(\b[56] ), .ZN(new_n10308_));
  OAI22_X1   g10052(.A1(new_n277_), .A2(new_n10308_), .B1(new_n9972_), .B2(new_n262_), .ZN(new_n10309_));
  AOI21_X1   g10053(.A1(\b[54] ), .A2(new_n283_), .B(new_n10309_), .ZN(new_n10310_));
  XOR2_X1    g10054(.A1(\b[55] ), .A2(\b[56] ), .Z(new_n10311_));
  INV_X1     g10055(.I(new_n10311_), .ZN(new_n10312_));
  OAI21_X1   g10056(.A1(new_n9975_), .A2(\b[54] ), .B(\b[55] ), .ZN(new_n10313_));
  NAND2_X1   g10057(.A1(new_n9973_), .A2(\b[54] ), .ZN(new_n10314_));
  NAND2_X1   g10058(.A1(new_n10313_), .A2(new_n10314_), .ZN(new_n10315_));
  NAND2_X1   g10059(.A1(new_n10315_), .A2(new_n10312_), .ZN(new_n10316_));
  NAND3_X1   g10060(.A1(new_n10313_), .A2(new_n10314_), .A3(new_n10311_), .ZN(new_n10317_));
  NAND2_X1   g10061(.A1(new_n10316_), .A2(new_n10317_), .ZN(new_n10318_));
  INV_X1     g10062(.I(new_n10318_), .ZN(new_n10319_));
  OAI21_X1   g10063(.A1(new_n10319_), .A2(new_n279_), .B(new_n10310_), .ZN(new_n10320_));
  XOR2_X1    g10064(.A1(new_n10320_), .A2(\a[2] ), .Z(new_n10321_));
  INV_X1     g10065(.I(new_n10321_), .ZN(new_n10322_));
  AOI22_X1   g10066(.A1(new_n518_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n636_), .ZN(new_n10323_));
  OAI21_X1   g10067(.A1(new_n8127_), .A2(new_n917_), .B(new_n10323_), .ZN(new_n10324_));
  AOI21_X1   g10068(.A1(new_n9684_), .A2(new_n618_), .B(new_n10324_), .ZN(new_n10325_));
  XOR2_X1    g10069(.A1(new_n10325_), .A2(new_n488_), .Z(new_n10326_));
  NAND3_X1   g10070(.A1(new_n9994_), .A2(new_n9917_), .A3(new_n10237_), .ZN(new_n10327_));
  OAI22_X1   g10071(.A1(new_n713_), .A2(new_n8126_), .B1(new_n7617_), .B2(new_n717_), .ZN(new_n10328_));
  AOI21_X1   g10072(.A1(\b[45] ), .A2(new_n1126_), .B(new_n10328_), .ZN(new_n10329_));
  NAND2_X1   g10073(.A1(new_n7649_), .A2(new_n724_), .ZN(new_n10330_));
  AOI21_X1   g10074(.A1(new_n10330_), .A2(new_n10329_), .B(new_n722_), .ZN(new_n10331_));
  NAND3_X1   g10075(.A1(new_n10330_), .A2(new_n722_), .A3(new_n10329_), .ZN(new_n10332_));
  INV_X1     g10076(.I(new_n10332_), .ZN(new_n10333_));
  NOR2_X1    g10077(.A1(new_n10333_), .A2(new_n10331_), .ZN(new_n10334_));
  AOI21_X1   g10078(.A1(new_n9997_), .A2(new_n9896_), .B(new_n10221_), .ZN(new_n10335_));
  OAI22_X1   g10079(.A1(new_n993_), .A2(new_n7074_), .B1(new_n6775_), .B2(new_n997_), .ZN(new_n10336_));
  AOI21_X1   g10080(.A1(\b[42] ), .A2(new_n1486_), .B(new_n10336_), .ZN(new_n10337_));
  OAI21_X1   g10081(.A1(new_n7081_), .A2(new_n1323_), .B(new_n10337_), .ZN(new_n10338_));
  XOR2_X1    g10082(.A1(new_n10338_), .A2(\a[14] ), .Z(new_n10339_));
  INV_X1     g10083(.I(new_n10339_), .ZN(new_n10340_));
  OAI22_X1   g10084(.A1(new_n1592_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n1505_), .ZN(new_n10341_));
  AOI21_X1   g10085(.A1(\b[39] ), .A2(new_n1584_), .B(new_n10341_), .ZN(new_n10342_));
  OAI21_X1   g10086(.A1(new_n6299_), .A2(new_n1732_), .B(new_n10342_), .ZN(new_n10343_));
  XOR2_X1    g10087(.A1(new_n10343_), .A2(new_n1344_), .Z(new_n10344_));
  AOI22_X1   g10088(.A1(new_n1738_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n1743_), .ZN(new_n10345_));
  OAI21_X1   g10089(.A1(new_n4886_), .A2(new_n1931_), .B(new_n10345_), .ZN(new_n10346_));
  AOI21_X1   g10090(.A1(new_n5351_), .A2(new_n1746_), .B(new_n10346_), .ZN(new_n10347_));
  XOR2_X1    g10091(.A1(new_n10347_), .A2(new_n1736_), .Z(new_n10348_));
  INV_X1     g10092(.I(new_n10348_), .ZN(new_n10349_));
  OAI22_X1   g10093(.A1(new_n2189_), .A2(new_n4666_), .B1(new_n4639_), .B2(new_n2194_), .ZN(new_n10350_));
  AOI21_X1   g10094(.A1(\b[33] ), .A2(new_n2361_), .B(new_n10350_), .ZN(new_n10351_));
  OAI21_X1   g10095(.A1(new_n4676_), .A2(new_n2197_), .B(new_n10351_), .ZN(new_n10352_));
  XOR2_X1    g10096(.A1(new_n10352_), .A2(\a[23] ), .Z(new_n10353_));
  INV_X1     g10097(.I(new_n10353_), .ZN(new_n10354_));
  NOR3_X1    g10098(.A1(new_n10166_), .A2(new_n10171_), .A3(new_n10173_), .ZN(new_n10355_));
  INV_X1     g10099(.I(new_n10355_), .ZN(new_n10356_));
  AOI22_X1   g10100(.A1(new_n2716_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n2719_), .ZN(new_n10357_));
  OAI21_X1   g10101(.A1(new_n3624_), .A2(new_n2924_), .B(new_n10357_), .ZN(new_n10358_));
  AOI21_X1   g10102(.A1(new_n4030_), .A2(new_n2722_), .B(new_n10358_), .ZN(new_n10359_));
  XOR2_X1    g10103(.A1(new_n10359_), .A2(new_n2714_), .Z(new_n10360_));
  NAND2_X1   g10104(.A1(new_n10139_), .A2(new_n9799_), .ZN(new_n10361_));
  INV_X1     g10105(.I(new_n10146_), .ZN(new_n10362_));
  NAND2_X1   g10106(.A1(new_n10361_), .A2(new_n10362_), .ZN(new_n10363_));
  XNOR2_X1   g10107(.A1(new_n10136_), .A2(new_n10142_), .ZN(new_n10364_));
  OAI21_X1   g10108(.A1(new_n10361_), .A2(new_n10362_), .B(new_n10364_), .ZN(new_n10365_));
  NOR2_X1    g10109(.A1(new_n10142_), .A2(new_n10135_), .ZN(new_n10366_));
  NAND2_X1   g10110(.A1(new_n10124_), .A2(new_n10131_), .ZN(new_n10367_));
  NOR2_X1    g10111(.A1(new_n10035_), .A2(new_n10044_), .ZN(new_n10368_));
  XOR2_X1    g10112(.A1(new_n10110_), .A2(new_n10037_), .Z(new_n10369_));
  AOI21_X1   g10113(.A1(new_n10035_), .A2(new_n10044_), .B(new_n10369_), .ZN(new_n10370_));
  NOR2_X1    g10114(.A1(new_n10370_), .A2(new_n10368_), .ZN(new_n10371_));
  OAI22_X1   g10115(.A1(new_n5852_), .A2(new_n1432_), .B1(new_n1296_), .B2(new_n5857_), .ZN(new_n10372_));
  AOI21_X1   g10116(.A1(\b[15] ), .A2(new_n6115_), .B(new_n10372_), .ZN(new_n10373_));
  OAI21_X1   g10117(.A1(new_n1444_), .A2(new_n5861_), .B(new_n10373_), .ZN(new_n10374_));
  XOR2_X1    g10118(.A1(new_n10374_), .A2(\a[41] ), .Z(new_n10375_));
  AOI22_X1   g10119(.A1(new_n6569_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n6574_), .ZN(new_n10376_));
  OAI21_X1   g10120(.A1(new_n941_), .A2(new_n8565_), .B(new_n10376_), .ZN(new_n10377_));
  AOI21_X1   g10121(.A1(new_n1449_), .A2(new_n6579_), .B(new_n10377_), .ZN(new_n10378_));
  XOR2_X1    g10122(.A1(new_n10378_), .A2(new_n6567_), .Z(new_n10379_));
  NOR2_X1    g10123(.A1(new_n10047_), .A2(new_n10100_), .ZN(new_n10380_));
  OAI22_X1   g10124(.A1(new_n776_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n852_), .ZN(new_n10381_));
  AOI21_X1   g10125(.A1(\b[9] ), .A2(new_n7719_), .B(new_n10381_), .ZN(new_n10382_));
  OAI21_X1   g10126(.A1(new_n859_), .A2(new_n8585_), .B(new_n10382_), .ZN(new_n10383_));
  XOR2_X1    g10127(.A1(new_n10383_), .A2(\a[47] ), .Z(new_n10384_));
  OAI21_X1   g10128(.A1(new_n10049_), .A2(new_n9737_), .B(new_n10087_), .ZN(new_n10385_));
  NAND3_X1   g10129(.A1(new_n10076_), .A2(new_n10051_), .A3(new_n9731_), .ZN(new_n10386_));
  NAND2_X1   g10130(.A1(new_n10386_), .A2(new_n10077_), .ZN(new_n10387_));
  INV_X1     g10131(.I(new_n9129_), .ZN(new_n10388_));
  INV_X1     g10132(.I(new_n9123_), .ZN(new_n10389_));
  INV_X1     g10133(.I(new_n9125_), .ZN(new_n10390_));
  OAI22_X1   g10134(.A1(new_n10390_), .A2(new_n377_), .B1(new_n339_), .B2(new_n10389_), .ZN(new_n10391_));
  AOI21_X1   g10135(.A1(\b[3] ), .A2(new_n9471_), .B(new_n10391_), .ZN(new_n10392_));
  OAI21_X1   g10136(.A1(new_n566_), .A2(new_n10388_), .B(new_n10392_), .ZN(new_n10393_));
  XOR2_X1    g10137(.A1(new_n10393_), .A2(\a[53] ), .Z(new_n10394_));
  INV_X1     g10138(.I(new_n10070_), .ZN(new_n10395_));
  AOI22_X1   g10139(.A1(new_n10064_), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n10062_), .ZN(new_n10396_));
  NOR4_X1    g10140(.A1(new_n9133_), .A2(new_n10058_), .A3(new_n10060_), .A4(\a[56] ), .ZN(new_n10397_));
  NOR4_X1    g10141(.A1(new_n10057_), .A2(\a[53] ), .A3(\a[54] ), .A4(\a[55] ), .ZN(new_n10398_));
  NOR2_X1    g10142(.A1(new_n10397_), .A2(new_n10398_), .ZN(new_n10399_));
  OAI21_X1   g10143(.A1(new_n258_), .A2(new_n10399_), .B(new_n10396_), .ZN(new_n10400_));
  AOI21_X1   g10144(.A1(new_n554_), .A2(new_n10068_), .B(new_n10400_), .ZN(new_n10401_));
  AND4_X2    g10145(.A1(\a[56] ), .A2(new_n10401_), .A3(new_n9733_), .A4(new_n10395_), .Z(new_n10402_));
  INV_X1     g10146(.I(new_n10071_), .ZN(new_n10403_));
  XOR2_X1    g10147(.A1(new_n10401_), .A2(new_n10057_), .Z(new_n10404_));
  NOR2_X1    g10148(.A1(new_n10404_), .A2(new_n10403_), .ZN(new_n10405_));
  NOR2_X1    g10149(.A1(new_n10405_), .A2(new_n10402_), .ZN(new_n10406_));
  NOR2_X1    g10150(.A1(new_n10406_), .A2(new_n10394_), .ZN(new_n10407_));
  INV_X1     g10151(.I(new_n10407_), .ZN(new_n10408_));
  NAND2_X1   g10152(.A1(new_n10406_), .A2(new_n10394_), .ZN(new_n10409_));
  NAND2_X1   g10153(.A1(new_n10408_), .A2(new_n10409_), .ZN(new_n10410_));
  NOR2_X1    g10154(.A1(new_n10410_), .A2(new_n10387_), .ZN(new_n10411_));
  NAND2_X1   g10155(.A1(new_n10410_), .A2(new_n10387_), .ZN(new_n10412_));
  INV_X1     g10156(.I(new_n10412_), .ZN(new_n10413_));
  AOI22_X1   g10157(.A1(new_n8241_), .A2(\b[8] ), .B1(\b[7] ), .B2(new_n8246_), .ZN(new_n10414_));
  OAI21_X1   g10158(.A1(new_n438_), .A2(new_n9114_), .B(new_n10414_), .ZN(new_n10415_));
  AOI21_X1   g10159(.A1(new_n799_), .A2(new_n8252_), .B(new_n10415_), .ZN(new_n10416_));
  XOR2_X1    g10160(.A1(new_n10416_), .A2(new_n8248_), .Z(new_n10417_));
  INV_X1     g10161(.I(new_n10417_), .ZN(new_n10418_));
  NOR3_X1    g10162(.A1(new_n10413_), .A2(new_n10411_), .A3(new_n10418_), .ZN(new_n10419_));
  INV_X1     g10163(.I(new_n10411_), .ZN(new_n10420_));
  AOI21_X1   g10164(.A1(new_n10420_), .A2(new_n10412_), .B(new_n10417_), .ZN(new_n10421_));
  NOR2_X1    g10165(.A1(new_n10421_), .A2(new_n10419_), .ZN(new_n10422_));
  NAND3_X1   g10166(.A1(new_n10422_), .A2(new_n10385_), .A3(new_n10085_), .ZN(new_n10423_));
  INV_X1     g10167(.I(new_n10085_), .ZN(new_n10424_));
  AOI21_X1   g10168(.A1(new_n10086_), .A2(new_n10083_), .B(new_n10050_), .ZN(new_n10425_));
  OR2_X2     g10169(.A1(new_n10421_), .A2(new_n10419_), .Z(new_n10426_));
  OAI21_X1   g10170(.A1(new_n10424_), .A2(new_n10425_), .B(new_n10426_), .ZN(new_n10427_));
  NAND3_X1   g10171(.A1(new_n10427_), .A2(new_n10384_), .A3(new_n10423_), .ZN(new_n10428_));
  INV_X1     g10172(.I(new_n10384_), .ZN(new_n10429_));
  NOR3_X1    g10173(.A1(new_n10426_), .A2(new_n10425_), .A3(new_n10424_), .ZN(new_n10430_));
  AOI21_X1   g10174(.A1(new_n10085_), .A2(new_n10385_), .B(new_n10422_), .ZN(new_n10431_));
  OAI21_X1   g10175(.A1(new_n10430_), .A2(new_n10431_), .B(new_n10429_), .ZN(new_n10432_));
  NAND2_X1   g10176(.A1(new_n10428_), .A2(new_n10432_), .ZN(new_n10433_));
  NOR3_X1    g10177(.A1(new_n10380_), .A2(new_n10433_), .A3(new_n10099_), .ZN(new_n10434_));
  INV_X1     g10178(.I(new_n10434_), .ZN(new_n10435_));
  OAI21_X1   g10179(.A1(new_n10380_), .A2(new_n10099_), .B(new_n10433_), .ZN(new_n10436_));
  AOI21_X1   g10180(.A1(new_n10435_), .A2(new_n10436_), .B(new_n10379_), .ZN(new_n10437_));
  INV_X1     g10181(.I(new_n10379_), .ZN(new_n10438_));
  INV_X1     g10182(.I(new_n10436_), .ZN(new_n10439_));
  NOR3_X1    g10183(.A1(new_n10439_), .A2(new_n10434_), .A3(new_n10438_), .ZN(new_n10440_));
  NOR2_X1    g10184(.A1(new_n10440_), .A2(new_n10437_), .ZN(new_n10441_));
  NAND3_X1   g10185(.A1(new_n10036_), .A2(new_n9758_), .A3(new_n10107_), .ZN(new_n10442_));
  NAND2_X1   g10186(.A1(new_n10442_), .A2(new_n10109_), .ZN(new_n10443_));
  NAND2_X1   g10187(.A1(new_n10443_), .A2(new_n10441_), .ZN(new_n10444_));
  OAI21_X1   g10188(.A1(new_n10439_), .A2(new_n10434_), .B(new_n10438_), .ZN(new_n10445_));
  NAND3_X1   g10189(.A1(new_n10435_), .A2(new_n10436_), .A3(new_n10379_), .ZN(new_n10446_));
  NAND2_X1   g10190(.A1(new_n10445_), .A2(new_n10446_), .ZN(new_n10447_));
  NAND3_X1   g10191(.A1(new_n10447_), .A2(new_n10109_), .A3(new_n10442_), .ZN(new_n10448_));
  AOI21_X1   g10192(.A1(new_n10444_), .A2(new_n10448_), .B(new_n10375_), .ZN(new_n10449_));
  INV_X1     g10193(.I(new_n10375_), .ZN(new_n10450_));
  AOI21_X1   g10194(.A1(new_n10109_), .A2(new_n10442_), .B(new_n10447_), .ZN(new_n10451_));
  NOR2_X1    g10195(.A1(new_n10443_), .A2(new_n10441_), .ZN(new_n10452_));
  NOR3_X1    g10196(.A1(new_n10452_), .A2(new_n10451_), .A3(new_n10450_), .ZN(new_n10453_));
  NOR2_X1    g10197(.A1(new_n10453_), .A2(new_n10449_), .ZN(new_n10454_));
  NOR2_X1    g10198(.A1(new_n10371_), .A2(new_n10454_), .ZN(new_n10455_));
  OAI21_X1   g10199(.A1(new_n10452_), .A2(new_n10451_), .B(new_n10450_), .ZN(new_n10456_));
  NAND3_X1   g10200(.A1(new_n10444_), .A2(new_n10375_), .A3(new_n10448_), .ZN(new_n10457_));
  NAND2_X1   g10201(.A1(new_n10456_), .A2(new_n10457_), .ZN(new_n10458_));
  NOR3_X1    g10202(.A1(new_n10458_), .A2(new_n10368_), .A3(new_n10370_), .ZN(new_n10459_));
  AOI22_X1   g10203(.A1(new_n5155_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n5160_), .ZN(new_n10460_));
  OAI21_X1   g10204(.A1(new_n1553_), .A2(new_n6877_), .B(new_n10460_), .ZN(new_n10461_));
  AOI21_X1   g10205(.A1(new_n2452_), .A2(new_n5166_), .B(new_n10461_), .ZN(new_n10462_));
  XOR2_X1    g10206(.A1(new_n10462_), .A2(new_n5162_), .Z(new_n10463_));
  INV_X1     g10207(.I(new_n10463_), .ZN(new_n10464_));
  OAI21_X1   g10208(.A1(new_n10455_), .A2(new_n10459_), .B(new_n10464_), .ZN(new_n10465_));
  OAI21_X1   g10209(.A1(new_n10370_), .A2(new_n10368_), .B(new_n10458_), .ZN(new_n10466_));
  NAND2_X1   g10210(.A1(new_n10371_), .A2(new_n10454_), .ZN(new_n10467_));
  NAND3_X1   g10211(.A1(new_n10467_), .A2(new_n10466_), .A3(new_n10463_), .ZN(new_n10468_));
  NAND4_X1   g10212(.A1(new_n10367_), .A2(new_n10121_), .A3(new_n10465_), .A4(new_n10468_), .ZN(new_n10469_));
  OAI21_X1   g10213(.A1(new_n10034_), .A2(new_n10133_), .B(new_n10121_), .ZN(new_n10470_));
  NAND2_X1   g10214(.A1(new_n10465_), .A2(new_n10468_), .ZN(new_n10471_));
  NAND2_X1   g10215(.A1(new_n10470_), .A2(new_n10471_), .ZN(new_n10472_));
  AOI22_X1   g10216(.A1(new_n4918_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n4921_), .ZN(new_n10473_));
  OAI21_X1   g10217(.A1(new_n2027_), .A2(new_n6099_), .B(new_n10473_), .ZN(new_n10474_));
  AOI21_X1   g10218(.A1(new_n2470_), .A2(new_n4699_), .B(new_n10474_), .ZN(new_n10475_));
  XOR2_X1    g10219(.A1(new_n10475_), .A2(new_n4446_), .Z(new_n10476_));
  NAND3_X1   g10220(.A1(new_n10472_), .A2(new_n10469_), .A3(new_n10476_), .ZN(new_n10477_));
  NOR2_X1    g10221(.A1(new_n10470_), .A2(new_n10471_), .ZN(new_n10478_));
  AOI22_X1   g10222(.A1(new_n10367_), .A2(new_n10121_), .B1(new_n10465_), .B2(new_n10468_), .ZN(new_n10479_));
  INV_X1     g10223(.I(new_n10476_), .ZN(new_n10480_));
  OAI21_X1   g10224(.A1(new_n10478_), .A2(new_n10479_), .B(new_n10480_), .ZN(new_n10481_));
  NAND2_X1   g10225(.A1(new_n10481_), .A2(new_n10477_), .ZN(new_n10482_));
  NOR3_X1    g10226(.A1(new_n10482_), .A2(new_n10128_), .A3(new_n10366_), .ZN(new_n10483_));
  NOR2_X1    g10227(.A1(new_n10366_), .A2(new_n10128_), .ZN(new_n10484_));
  NOR3_X1    g10228(.A1(new_n10478_), .A2(new_n10479_), .A3(new_n10480_), .ZN(new_n10485_));
  AOI21_X1   g10229(.A1(new_n10472_), .A2(new_n10469_), .B(new_n10476_), .ZN(new_n10486_));
  NOR2_X1    g10230(.A1(new_n10485_), .A2(new_n10486_), .ZN(new_n10487_));
  NOR2_X1    g10231(.A1(new_n10484_), .A2(new_n10487_), .ZN(new_n10488_));
  NOR2_X1    g10232(.A1(new_n10488_), .A2(new_n10483_), .ZN(new_n10489_));
  NAND3_X1   g10233(.A1(new_n10365_), .A2(new_n10363_), .A3(new_n10489_), .ZN(new_n10490_));
  NOR2_X1    g10234(.A1(new_n10028_), .A2(new_n10026_), .ZN(new_n10491_));
  NOR2_X1    g10235(.A1(new_n10491_), .A2(new_n10146_), .ZN(new_n10492_));
  XOR2_X1    g10236(.A1(new_n10136_), .A2(new_n10142_), .Z(new_n10493_));
  AOI21_X1   g10237(.A1(new_n10491_), .A2(new_n10146_), .B(new_n10493_), .ZN(new_n10494_));
  INV_X1     g10238(.I(new_n10489_), .ZN(new_n10495_));
  OAI21_X1   g10239(.A1(new_n10494_), .A2(new_n10492_), .B(new_n10495_), .ZN(new_n10496_));
  AOI22_X1   g10240(.A1(new_n3267_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n3270_), .ZN(new_n10497_));
  OAI21_X1   g10241(.A1(new_n3158_), .A2(new_n3475_), .B(new_n10497_), .ZN(new_n10498_));
  AOI21_X1   g10242(.A1(new_n4188_), .A2(new_n3273_), .B(new_n10498_), .ZN(new_n10499_));
  XOR2_X1    g10243(.A1(new_n10499_), .A2(\a[29] ), .Z(new_n10500_));
  AOI22_X1   g10244(.A1(new_n3864_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n3869_), .ZN(new_n10501_));
  OAI21_X1   g10245(.A1(new_n2495_), .A2(new_n5410_), .B(new_n10501_), .ZN(new_n10502_));
  AOI21_X1   g10246(.A1(new_n3407_), .A2(new_n3872_), .B(new_n10502_), .ZN(new_n10503_));
  XOR2_X1    g10247(.A1(new_n10503_), .A2(new_n3876_), .Z(new_n10504_));
  XOR2_X1    g10248(.A1(new_n10500_), .A2(new_n10504_), .Z(new_n10505_));
  AOI21_X1   g10249(.A1(new_n10496_), .A2(new_n10490_), .B(new_n10505_), .ZN(new_n10506_));
  NOR3_X1    g10250(.A1(new_n10494_), .A2(new_n10492_), .A3(new_n10495_), .ZN(new_n10507_));
  AOI21_X1   g10251(.A1(new_n10365_), .A2(new_n10363_), .B(new_n10489_), .ZN(new_n10508_));
  INV_X1     g10252(.I(new_n10505_), .ZN(new_n10509_));
  NOR3_X1    g10253(.A1(new_n10507_), .A2(new_n10508_), .A3(new_n10509_), .ZN(new_n10510_));
  OAI22_X1   g10254(.A1(new_n10166_), .A2(new_n10161_), .B1(new_n10506_), .B2(new_n10510_), .ZN(new_n10511_));
  OAI21_X1   g10255(.A1(new_n10507_), .A2(new_n10508_), .B(new_n10509_), .ZN(new_n10512_));
  NAND3_X1   g10256(.A1(new_n10496_), .A2(new_n10490_), .A3(new_n10505_), .ZN(new_n10513_));
  NAND4_X1   g10257(.A1(new_n10174_), .A2(new_n10168_), .A3(new_n10512_), .A4(new_n10513_), .ZN(new_n10514_));
  NAND3_X1   g10258(.A1(new_n10511_), .A2(new_n10514_), .A3(new_n10360_), .ZN(new_n10515_));
  INV_X1     g10259(.I(new_n10360_), .ZN(new_n10516_));
  AOI22_X1   g10260(.A1(new_n10174_), .A2(new_n10168_), .B1(new_n10512_), .B2(new_n10513_), .ZN(new_n10517_));
  NOR4_X1    g10261(.A1(new_n10166_), .A2(new_n10161_), .A3(new_n10506_), .A4(new_n10510_), .ZN(new_n10518_));
  OAI21_X1   g10262(.A1(new_n10518_), .A2(new_n10517_), .B(new_n10516_), .ZN(new_n10519_));
  NAND2_X1   g10263(.A1(new_n10519_), .A2(new_n10515_), .ZN(new_n10520_));
  AOI21_X1   g10264(.A1(new_n10178_), .A2(new_n10356_), .B(new_n10520_), .ZN(new_n10521_));
  NOR3_X1    g10265(.A1(new_n10518_), .A2(new_n10517_), .A3(new_n10516_), .ZN(new_n10522_));
  AOI21_X1   g10266(.A1(new_n10511_), .A2(new_n10514_), .B(new_n10360_), .ZN(new_n10523_));
  NOR2_X1    g10267(.A1(new_n10522_), .A2(new_n10523_), .ZN(new_n10524_));
  NOR3_X1    g10268(.A1(new_n10186_), .A2(new_n10524_), .A3(new_n10355_), .ZN(new_n10525_));
  OAI21_X1   g10269(.A1(new_n10521_), .A2(new_n10525_), .B(new_n10354_), .ZN(new_n10526_));
  OAI21_X1   g10270(.A1(new_n10186_), .A2(new_n10355_), .B(new_n10524_), .ZN(new_n10527_));
  NAND3_X1   g10271(.A1(new_n10178_), .A2(new_n10520_), .A3(new_n10356_), .ZN(new_n10528_));
  NAND3_X1   g10272(.A1(new_n10527_), .A2(new_n10528_), .A3(new_n10353_), .ZN(new_n10529_));
  NAND2_X1   g10273(.A1(new_n10526_), .A2(new_n10529_), .ZN(new_n10530_));
  AOI21_X1   g10274(.A1(new_n10198_), .A2(new_n10184_), .B(new_n10530_), .ZN(new_n10531_));
  AOI21_X1   g10275(.A1(new_n10527_), .A2(new_n10528_), .B(new_n10353_), .ZN(new_n10532_));
  NOR3_X1    g10276(.A1(new_n10521_), .A2(new_n10525_), .A3(new_n10354_), .ZN(new_n10533_));
  NOR2_X1    g10277(.A1(new_n10533_), .A2(new_n10532_), .ZN(new_n10534_));
  NOR3_X1    g10278(.A1(new_n10190_), .A2(new_n10534_), .A3(new_n10192_), .ZN(new_n10535_));
  OAI21_X1   g10279(.A1(new_n10535_), .A2(new_n10531_), .B(new_n10349_), .ZN(new_n10536_));
  OAI21_X1   g10280(.A1(new_n10190_), .A2(new_n10192_), .B(new_n10534_), .ZN(new_n10537_));
  NAND3_X1   g10281(.A1(new_n10198_), .A2(new_n10530_), .A3(new_n10184_), .ZN(new_n10538_));
  NAND3_X1   g10282(.A1(new_n10537_), .A2(new_n10538_), .A3(new_n10348_), .ZN(new_n10539_));
  NAND2_X1   g10283(.A1(new_n10536_), .A2(new_n10539_), .ZN(new_n10540_));
  NOR3_X1    g10284(.A1(new_n10190_), .A2(new_n10195_), .A3(new_n10197_), .ZN(new_n10541_));
  INV_X1     g10285(.I(new_n10541_), .ZN(new_n10542_));
  AOI21_X1   g10286(.A1(new_n10202_), .A2(new_n10542_), .B(new_n10540_), .ZN(new_n10543_));
  AOI21_X1   g10287(.A1(new_n10537_), .A2(new_n10538_), .B(new_n10348_), .ZN(new_n10544_));
  NOR3_X1    g10288(.A1(new_n10535_), .A2(new_n10531_), .A3(new_n10349_), .ZN(new_n10545_));
  NOR2_X1    g10289(.A1(new_n10545_), .A2(new_n10544_), .ZN(new_n10546_));
  NOR3_X1    g10290(.A1(new_n10210_), .A2(new_n10541_), .A3(new_n10546_), .ZN(new_n10547_));
  OAI21_X1   g10291(.A1(new_n10547_), .A2(new_n10543_), .B(new_n10344_), .ZN(new_n10548_));
  XOR2_X1    g10292(.A1(new_n10343_), .A2(\a[17] ), .Z(new_n10549_));
  OAI21_X1   g10293(.A1(new_n10210_), .A2(new_n10541_), .B(new_n10546_), .ZN(new_n10550_));
  NAND3_X1   g10294(.A1(new_n10202_), .A2(new_n10540_), .A3(new_n10542_), .ZN(new_n10551_));
  NAND3_X1   g10295(.A1(new_n10550_), .A2(new_n10551_), .A3(new_n10549_), .ZN(new_n10552_));
  NAND2_X1   g10296(.A1(new_n10548_), .A2(new_n10552_), .ZN(new_n10553_));
  AOI21_X1   g10297(.A1(new_n10227_), .A2(new_n10208_), .B(new_n10553_), .ZN(new_n10554_));
  AOI21_X1   g10298(.A1(new_n10550_), .A2(new_n10551_), .B(new_n10549_), .ZN(new_n10555_));
  NOR3_X1    g10299(.A1(new_n10547_), .A2(new_n10543_), .A3(new_n10344_), .ZN(new_n10556_));
  NOR2_X1    g10300(.A1(new_n10556_), .A2(new_n10555_), .ZN(new_n10557_));
  NOR3_X1    g10301(.A1(new_n10214_), .A2(new_n10557_), .A3(new_n10216_), .ZN(new_n10558_));
  NOR3_X1    g10302(.A1(new_n10558_), .A2(new_n10554_), .A3(new_n10340_), .ZN(new_n10559_));
  OAI21_X1   g10303(.A1(new_n10214_), .A2(new_n10216_), .B(new_n10557_), .ZN(new_n10560_));
  NAND3_X1   g10304(.A1(new_n10227_), .A2(new_n10553_), .A3(new_n10208_), .ZN(new_n10561_));
  AOI21_X1   g10305(.A1(new_n10560_), .A2(new_n10561_), .B(new_n10339_), .ZN(new_n10562_));
  NOR2_X1    g10306(.A1(new_n10559_), .A2(new_n10562_), .ZN(new_n10563_));
  OAI21_X1   g10307(.A1(new_n10335_), .A2(new_n10229_), .B(new_n10563_), .ZN(new_n10564_));
  NAND3_X1   g10308(.A1(new_n9887_), .A2(new_n9882_), .A3(new_n9874_), .ZN(new_n10565_));
  OAI21_X1   g10309(.A1(new_n9875_), .A2(new_n9878_), .B(new_n9869_), .ZN(new_n10566_));
  NAND2_X1   g10310(.A1(new_n10566_), .A2(new_n10565_), .ZN(new_n10567_));
  AOI21_X1   g10311(.A1(new_n9315_), .A2(new_n9318_), .B(new_n9316_), .ZN(new_n10568_));
  OAI21_X1   g10312(.A1(new_n10568_), .A2(new_n9647_), .B(new_n9646_), .ZN(new_n10569_));
  AOI21_X1   g10313(.A1(new_n10569_), .A2(new_n9893_), .B(new_n10567_), .ZN(new_n10570_));
  OAI21_X1   g10314(.A1(new_n10570_), .A2(new_n10225_), .B(new_n10222_), .ZN(new_n10571_));
  NAND3_X1   g10315(.A1(new_n10560_), .A2(new_n10561_), .A3(new_n10339_), .ZN(new_n10572_));
  OAI21_X1   g10316(.A1(new_n10558_), .A2(new_n10554_), .B(new_n10340_), .ZN(new_n10573_));
  NAND2_X1   g10317(.A1(new_n10573_), .A2(new_n10572_), .ZN(new_n10574_));
  NAND3_X1   g10318(.A1(new_n10571_), .A2(new_n10574_), .A3(new_n10220_), .ZN(new_n10575_));
  NAND3_X1   g10319(.A1(new_n10564_), .A2(new_n10575_), .A3(new_n10334_), .ZN(new_n10576_));
  INV_X1     g10320(.I(new_n10334_), .ZN(new_n10577_));
  AOI21_X1   g10321(.A1(new_n10571_), .A2(new_n10220_), .B(new_n10574_), .ZN(new_n10578_));
  NOR3_X1    g10322(.A1(new_n10335_), .A2(new_n10563_), .A3(new_n10229_), .ZN(new_n10579_));
  OAI21_X1   g10323(.A1(new_n10578_), .A2(new_n10579_), .B(new_n10577_), .ZN(new_n10580_));
  NAND2_X1   g10324(.A1(new_n10580_), .A2(new_n10576_), .ZN(new_n10581_));
  AOI21_X1   g10325(.A1(new_n10327_), .A2(new_n10240_), .B(new_n10581_), .ZN(new_n10582_));
  NOR3_X1    g10326(.A1(new_n10243_), .A2(new_n9912_), .A3(new_n10244_), .ZN(new_n10583_));
  NOR3_X1    g10327(.A1(new_n10578_), .A2(new_n10579_), .A3(new_n10577_), .ZN(new_n10584_));
  AOI21_X1   g10328(.A1(new_n10564_), .A2(new_n10575_), .B(new_n10334_), .ZN(new_n10585_));
  NOR2_X1    g10329(.A1(new_n10585_), .A2(new_n10584_), .ZN(new_n10586_));
  NOR3_X1    g10330(.A1(new_n10583_), .A2(new_n10586_), .A3(new_n10245_), .ZN(new_n10587_));
  NOR3_X1    g10331(.A1(new_n10582_), .A2(new_n10587_), .A3(new_n10326_), .ZN(new_n10588_));
  INV_X1     g10332(.I(new_n10326_), .ZN(new_n10589_));
  OAI21_X1   g10333(.A1(new_n10583_), .A2(new_n10245_), .B(new_n10586_), .ZN(new_n10590_));
  NAND3_X1   g10334(.A1(new_n10327_), .A2(new_n10240_), .A3(new_n10581_), .ZN(new_n10591_));
  AOI21_X1   g10335(.A1(new_n10591_), .A2(new_n10590_), .B(new_n10589_), .ZN(new_n10592_));
  OR2_X2     g10336(.A1(new_n10592_), .A2(new_n10588_), .Z(new_n10593_));
  OAI21_X1   g10337(.A1(new_n9993_), .A2(new_n10260_), .B(new_n10256_), .ZN(new_n10594_));
  XOR2_X1    g10338(.A1(new_n10594_), .A2(new_n10593_), .Z(new_n10595_));
  INV_X1     g10339(.I(new_n10595_), .ZN(new_n10596_));
  OAI22_X1   g10340(.A1(new_n321_), .A2(new_n9376_), .B1(new_n325_), .B2(new_n9032_), .ZN(new_n10597_));
  AOI21_X1   g10341(.A1(\b[51] ), .A2(new_n602_), .B(new_n10597_), .ZN(new_n10598_));
  OAI21_X1   g10342(.A1(new_n9385_), .A2(new_n318_), .B(new_n10598_), .ZN(new_n10599_));
  XOR2_X1    g10343(.A1(new_n10599_), .A2(\a[5] ), .Z(new_n10600_));
  INV_X1     g10344(.I(new_n10600_), .ZN(new_n10601_));
  AOI21_X1   g10345(.A1(new_n10266_), .A2(new_n10268_), .B(new_n9992_), .ZN(new_n10602_));
  INV_X1     g10346(.I(new_n10602_), .ZN(new_n10603_));
  AOI21_X1   g10347(.A1(new_n10270_), .A2(new_n10603_), .B(new_n10601_), .ZN(new_n10604_));
  NOR3_X1    g10348(.A1(new_n10283_), .A2(new_n10600_), .A3(new_n10602_), .ZN(new_n10605_));
  NOR3_X1    g10349(.A1(new_n10604_), .A2(new_n10605_), .A3(new_n10596_), .ZN(new_n10606_));
  OAI21_X1   g10350(.A1(new_n10283_), .A2(new_n10602_), .B(new_n10600_), .ZN(new_n10607_));
  NAND3_X1   g10351(.A1(new_n10270_), .A2(new_n10601_), .A3(new_n10603_), .ZN(new_n10608_));
  AOI21_X1   g10352(.A1(new_n10608_), .A2(new_n10607_), .B(new_n10595_), .ZN(new_n10609_));
  OAI21_X1   g10353(.A1(new_n10606_), .A2(new_n10609_), .B(new_n10322_), .ZN(new_n10610_));
  NAND3_X1   g10354(.A1(new_n10608_), .A2(new_n10607_), .A3(new_n10595_), .ZN(new_n10611_));
  OAI21_X1   g10355(.A1(new_n10604_), .A2(new_n10605_), .B(new_n10596_), .ZN(new_n10612_));
  NAND3_X1   g10356(.A1(new_n10612_), .A2(new_n10611_), .A3(new_n10321_), .ZN(new_n10613_));
  NAND2_X1   g10357(.A1(new_n10610_), .A2(new_n10613_), .ZN(new_n10614_));
  XOR2_X1    g10358(.A1(new_n10614_), .A2(new_n10307_), .Z(\f[56] ));
  INV_X1     g10359(.I(new_n10306_), .ZN(new_n10616_));
  OAI21_X1   g10360(.A1(new_n10292_), .A2(new_n10288_), .B(new_n10616_), .ZN(new_n10617_));
  NOR3_X1    g10361(.A1(new_n10606_), .A2(new_n10609_), .A3(new_n10322_), .ZN(new_n10618_));
  AOI21_X1   g10362(.A1(new_n10617_), .A2(new_n10610_), .B(new_n10618_), .ZN(new_n10619_));
  NAND2_X1   g10363(.A1(new_n283_), .A2(\b[55] ), .ZN(new_n10620_));
  AOI22_X1   g10364(.A1(new_n267_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n261_), .ZN(new_n10621_));
  AOI21_X1   g10365(.A1(new_n10315_), .A2(\b[56] ), .B(new_n9972_), .ZN(new_n10622_));
  NOR2_X1    g10366(.A1(new_n10315_), .A2(\b[56] ), .ZN(new_n10623_));
  NOR2_X1    g10367(.A1(new_n10622_), .A2(new_n10623_), .ZN(new_n10624_));
  INV_X1     g10368(.I(\b[57] ), .ZN(new_n10625_));
  NAND3_X1   g10369(.A1(new_n10313_), .A2(new_n10314_), .A3(new_n10625_), .ZN(new_n10626_));
  NAND2_X1   g10370(.A1(new_n10315_), .A2(\b[57] ), .ZN(new_n10627_));
  AND2_X2    g10371(.A1(new_n10627_), .A2(new_n10626_), .Z(new_n10628_));
  NOR2_X1    g10372(.A1(new_n10628_), .A2(new_n10624_), .ZN(new_n10629_));
  AND2_X2    g10373(.A1(new_n10628_), .A2(new_n10624_), .Z(new_n10630_));
  NOR2_X1    g10374(.A1(new_n10630_), .A2(new_n10629_), .ZN(new_n10631_));
  NAND2_X1   g10375(.A1(new_n10631_), .A2(new_n265_), .ZN(new_n10632_));
  NAND3_X1   g10376(.A1(new_n10632_), .A2(new_n10620_), .A3(new_n10621_), .ZN(new_n10633_));
  XOR2_X1    g10377(.A1(new_n10633_), .A2(new_n270_), .Z(new_n10634_));
  OAI21_X1   g10378(.A1(new_n10271_), .A2(new_n10272_), .B(new_n10603_), .ZN(new_n10635_));
  AOI21_X1   g10379(.A1(new_n10635_), .A2(new_n10600_), .B(new_n10595_), .ZN(new_n10636_));
  NOR2_X1    g10380(.A1(new_n10592_), .A2(new_n10588_), .ZN(new_n10637_));
  AOI21_X1   g10381(.A1(new_n10259_), .A2(new_n10252_), .B(new_n10261_), .ZN(new_n10638_));
  AOI21_X1   g10382(.A1(new_n10638_), .A2(new_n10637_), .B(new_n10592_), .ZN(new_n10639_));
  AOI22_X1   g10383(.A1(new_n518_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n636_), .ZN(new_n10640_));
  OAI21_X1   g10384(.A1(new_n8168_), .A2(new_n917_), .B(new_n10640_), .ZN(new_n10641_));
  AOI21_X1   g10385(.A1(new_n8783_), .A2(new_n618_), .B(new_n10641_), .ZN(new_n10642_));
  XOR2_X1    g10386(.A1(new_n10642_), .A2(new_n488_), .Z(new_n10643_));
  INV_X1     g10387(.I(new_n10643_), .ZN(new_n10644_));
  NAND2_X1   g10388(.A1(new_n10470_), .A2(new_n10468_), .ZN(new_n10645_));
  NAND2_X1   g10389(.A1(new_n10645_), .A2(new_n10465_), .ZN(new_n10646_));
  AOI22_X1   g10390(.A1(new_n5155_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n5160_), .ZN(new_n10647_));
  OAI21_X1   g10391(.A1(new_n1859_), .A2(new_n6877_), .B(new_n10647_), .ZN(new_n10648_));
  AOI21_X1   g10392(.A1(new_n2032_), .A2(new_n5166_), .B(new_n10648_), .ZN(new_n10649_));
  XOR2_X1    g10393(.A1(new_n10649_), .A2(new_n5162_), .Z(new_n10650_));
  INV_X1     g10394(.I(new_n10650_), .ZN(new_n10651_));
  AOI22_X1   g10395(.A1(new_n6108_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n6111_), .ZN(new_n10652_));
  OAI21_X1   g10396(.A1(new_n1296_), .A2(new_n7708_), .B(new_n10652_), .ZN(new_n10653_));
  AOI21_X1   g10397(.A1(new_n2038_), .A2(new_n6105_), .B(new_n10653_), .ZN(new_n10654_));
  XOR2_X1    g10398(.A1(new_n10654_), .A2(new_n5849_), .Z(new_n10655_));
  INV_X1     g10399(.I(new_n10655_), .ZN(new_n10656_));
  AOI21_X1   g10400(.A1(new_n10387_), .A2(new_n10409_), .B(new_n10407_), .ZN(new_n10657_));
  AOI22_X1   g10401(.A1(new_n9125_), .A2(\b[6] ), .B1(\b[5] ), .B2(new_n9123_), .ZN(new_n10658_));
  OAI21_X1   g10402(.A1(new_n339_), .A2(new_n9470_), .B(new_n10658_), .ZN(new_n10659_));
  AOI21_X1   g10403(.A1(new_n916_), .A2(new_n9129_), .B(new_n10659_), .ZN(new_n10660_));
  XOR2_X1    g10404(.A1(new_n10660_), .A2(new_n9133_), .Z(new_n10661_));
  INV_X1     g10405(.I(new_n10661_), .ZN(new_n10662_));
  AOI22_X1   g10406(.A1(new_n10064_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n10062_), .ZN(new_n10663_));
  OAI21_X1   g10407(.A1(new_n275_), .A2(new_n10399_), .B(new_n10663_), .ZN(new_n10664_));
  AOI21_X1   g10408(.A1(new_n299_), .A2(new_n10068_), .B(new_n10664_), .ZN(new_n10665_));
  XOR2_X1    g10409(.A1(new_n10665_), .A2(\a[56] ), .Z(new_n10666_));
  NAND2_X1   g10410(.A1(\a[56] ), .A2(\a[57] ), .ZN(new_n10667_));
  NOR2_X1    g10411(.A1(\a[56] ), .A2(\a[57] ), .ZN(new_n10668_));
  INV_X1     g10412(.I(new_n10668_), .ZN(new_n10669_));
  NAND2_X1   g10413(.A1(new_n10669_), .A2(new_n10667_), .ZN(new_n10670_));
  NOR2_X1    g10414(.A1(new_n10670_), .A2(new_n258_), .ZN(new_n10671_));
  INV_X1     g10415(.I(new_n10671_), .ZN(new_n10672_));
  OR2_X2     g10416(.A1(new_n10666_), .A2(new_n10672_), .Z(new_n10673_));
  NAND2_X1   g10417(.A1(new_n10666_), .A2(new_n10672_), .ZN(new_n10674_));
  NAND2_X1   g10418(.A1(new_n10673_), .A2(new_n10674_), .ZN(new_n10675_));
  XOR2_X1    g10419(.A1(new_n10675_), .A2(new_n10402_), .Z(new_n10676_));
  NAND2_X1   g10420(.A1(new_n10676_), .A2(new_n10662_), .ZN(new_n10677_));
  NOR2_X1    g10421(.A1(new_n10676_), .A2(new_n10662_), .ZN(new_n10678_));
  INV_X1     g10422(.I(new_n10678_), .ZN(new_n10679_));
  NAND2_X1   g10423(.A1(new_n10679_), .A2(new_n10677_), .ZN(new_n10680_));
  XNOR2_X1   g10424(.A1(new_n10680_), .A2(new_n10657_), .ZN(new_n10681_));
  AOI22_X1   g10425(.A1(new_n8241_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n8246_), .ZN(new_n10682_));
  OAI21_X1   g10426(.A1(new_n471_), .A2(new_n9114_), .B(new_n10682_), .ZN(new_n10683_));
  AOI21_X1   g10427(.A1(new_n676_), .A2(new_n8252_), .B(new_n10683_), .ZN(new_n10684_));
  XOR2_X1    g10428(.A1(new_n10684_), .A2(new_n8248_), .Z(new_n10685_));
  INV_X1     g10429(.I(new_n10685_), .ZN(new_n10686_));
  NOR2_X1    g10430(.A1(new_n10430_), .A2(new_n10419_), .ZN(new_n10687_));
  NOR2_X1    g10431(.A1(new_n10687_), .A2(new_n10686_), .ZN(new_n10688_));
  NOR3_X1    g10432(.A1(new_n10430_), .A2(new_n10419_), .A3(new_n10685_), .ZN(new_n10689_));
  NOR2_X1    g10433(.A1(new_n10688_), .A2(new_n10689_), .ZN(new_n10690_));
  XOR2_X1    g10434(.A1(new_n10690_), .A2(new_n10681_), .Z(new_n10691_));
  INV_X1     g10435(.I(new_n10691_), .ZN(new_n10692_));
  AOI22_X1   g10436(.A1(new_n7403_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n7408_), .ZN(new_n10693_));
  OAI21_X1   g10437(.A1(new_n776_), .A2(new_n9488_), .B(new_n10693_), .ZN(new_n10694_));
  AOI21_X1   g10438(.A1(new_n1194_), .A2(new_n7414_), .B(new_n10694_), .ZN(new_n10695_));
  XOR2_X1    g10439(.A1(new_n10695_), .A2(new_n7410_), .Z(new_n10696_));
  NOR3_X1    g10440(.A1(new_n10430_), .A2(new_n10429_), .A3(new_n10431_), .ZN(new_n10697_));
  NOR2_X1    g10441(.A1(new_n10434_), .A2(new_n10697_), .ZN(new_n10698_));
  INV_X1     g10442(.I(new_n10698_), .ZN(new_n10699_));
  NAND2_X1   g10443(.A1(new_n10699_), .A2(new_n10696_), .ZN(new_n10700_));
  INV_X1     g10444(.I(new_n10696_), .ZN(new_n10701_));
  NAND2_X1   g10445(.A1(new_n10698_), .A2(new_n10701_), .ZN(new_n10702_));
  NAND2_X1   g10446(.A1(new_n10700_), .A2(new_n10702_), .ZN(new_n10703_));
  NOR2_X1    g10447(.A1(new_n10703_), .A2(new_n10692_), .ZN(new_n10704_));
  AOI21_X1   g10448(.A1(new_n10700_), .A2(new_n10702_), .B(new_n10691_), .ZN(new_n10705_));
  NOR2_X1    g10449(.A1(new_n10704_), .A2(new_n10705_), .ZN(new_n10706_));
  OAI22_X1   g10450(.A1(new_n7730_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n7731_), .ZN(new_n10707_));
  AOI21_X1   g10451(.A1(\b[13] ), .A2(new_n6887_), .B(new_n10707_), .ZN(new_n10708_));
  OAI21_X1   g10452(.A1(new_n1275_), .A2(new_n7728_), .B(new_n10708_), .ZN(new_n10709_));
  XOR2_X1    g10453(.A1(new_n10709_), .A2(\a[44] ), .Z(new_n10710_));
  OAI21_X1   g10454(.A1(new_n10451_), .A2(new_n10440_), .B(new_n10710_), .ZN(new_n10711_));
  INV_X1     g10455(.I(new_n10710_), .ZN(new_n10712_));
  NAND3_X1   g10456(.A1(new_n10444_), .A2(new_n10446_), .A3(new_n10712_), .ZN(new_n10713_));
  AND3_X2    g10457(.A1(new_n10713_), .A2(new_n10711_), .A3(new_n10706_), .Z(new_n10714_));
  AOI21_X1   g10458(.A1(new_n10711_), .A2(new_n10713_), .B(new_n10706_), .ZN(new_n10715_));
  OAI21_X1   g10459(.A1(new_n10714_), .A2(new_n10715_), .B(new_n10656_), .ZN(new_n10716_));
  NAND3_X1   g10460(.A1(new_n10711_), .A2(new_n10713_), .A3(new_n10706_), .ZN(new_n10717_));
  XOR2_X1    g10461(.A1(new_n10703_), .A2(new_n10691_), .Z(new_n10718_));
  NAND2_X1   g10462(.A1(new_n10713_), .A2(new_n10711_), .ZN(new_n10719_));
  NAND2_X1   g10463(.A1(new_n10719_), .A2(new_n10718_), .ZN(new_n10720_));
  NAND3_X1   g10464(.A1(new_n10720_), .A2(new_n10655_), .A3(new_n10717_), .ZN(new_n10721_));
  NAND2_X1   g10465(.A1(new_n10721_), .A2(new_n10716_), .ZN(new_n10722_));
  NOR2_X1    g10466(.A1(new_n10371_), .A2(new_n10453_), .ZN(new_n10723_));
  NOR3_X1    g10467(.A1(new_n10722_), .A2(new_n10449_), .A3(new_n10723_), .ZN(new_n10724_));
  AOI21_X1   g10468(.A1(new_n10720_), .A2(new_n10717_), .B(new_n10655_), .ZN(new_n10725_));
  NOR3_X1    g10469(.A1(new_n10714_), .A2(new_n10715_), .A3(new_n10656_), .ZN(new_n10726_));
  NOR2_X1    g10470(.A1(new_n10725_), .A2(new_n10726_), .ZN(new_n10727_));
  INV_X1     g10471(.I(new_n10723_), .ZN(new_n10728_));
  AOI21_X1   g10472(.A1(new_n10456_), .A2(new_n10728_), .B(new_n10727_), .ZN(new_n10729_));
  OAI21_X1   g10473(.A1(new_n10729_), .A2(new_n10724_), .B(new_n10651_), .ZN(new_n10730_));
  NAND3_X1   g10474(.A1(new_n10727_), .A2(new_n10728_), .A3(new_n10456_), .ZN(new_n10731_));
  OAI21_X1   g10475(.A1(new_n10723_), .A2(new_n10449_), .B(new_n10722_), .ZN(new_n10732_));
  NAND3_X1   g10476(.A1(new_n10732_), .A2(new_n10731_), .A3(new_n10650_), .ZN(new_n10733_));
  NAND2_X1   g10477(.A1(new_n10730_), .A2(new_n10733_), .ZN(new_n10734_));
  XNOR2_X1   g10478(.A1(new_n10734_), .A2(new_n10646_), .ZN(new_n10735_));
  AOI22_X1   g10479(.A1(new_n4918_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n4921_), .ZN(new_n10736_));
  OAI21_X1   g10480(.A1(new_n2142_), .A2(new_n6099_), .B(new_n10736_), .ZN(new_n10737_));
  AOI21_X1   g10481(.A1(new_n3033_), .A2(new_n4699_), .B(new_n10737_), .ZN(new_n10738_));
  XOR2_X1    g10482(.A1(new_n10738_), .A2(new_n4446_), .Z(new_n10739_));
  NAND2_X1   g10483(.A1(new_n10484_), .A2(new_n10487_), .ZN(new_n10740_));
  NAND2_X1   g10484(.A1(new_n10740_), .A2(new_n10477_), .ZN(new_n10741_));
  NAND2_X1   g10485(.A1(new_n10741_), .A2(new_n10739_), .ZN(new_n10742_));
  INV_X1     g10486(.I(new_n10739_), .ZN(new_n10743_));
  NOR2_X1    g10487(.A1(new_n10483_), .A2(new_n10485_), .ZN(new_n10744_));
  NAND2_X1   g10488(.A1(new_n10744_), .A2(new_n10743_), .ZN(new_n10745_));
  NAND3_X1   g10489(.A1(new_n10742_), .A2(new_n10745_), .A3(new_n10735_), .ZN(new_n10746_));
  XOR2_X1    g10490(.A1(new_n10734_), .A2(new_n10646_), .Z(new_n10747_));
  NOR2_X1    g10491(.A1(new_n10744_), .A2(new_n10743_), .ZN(new_n10748_));
  NOR2_X1    g10492(.A1(new_n10741_), .A2(new_n10739_), .ZN(new_n10749_));
  OAI21_X1   g10493(.A1(new_n10749_), .A2(new_n10748_), .B(new_n10747_), .ZN(new_n10750_));
  NAND2_X1   g10494(.A1(new_n10750_), .A2(new_n10746_), .ZN(new_n10751_));
  OAI22_X1   g10495(.A1(new_n3006_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n3158_), .ZN(new_n10752_));
  AOI21_X1   g10496(.A1(\b[25] ), .A2(new_n4053_), .B(new_n10752_), .ZN(new_n10753_));
  OAI21_X1   g10497(.A1(new_n3165_), .A2(new_n4727_), .B(new_n10753_), .ZN(new_n10754_));
  XOR2_X1    g10498(.A1(new_n10754_), .A2(\a[32] ), .Z(new_n10755_));
  INV_X1     g10499(.I(new_n10755_), .ZN(new_n10756_));
  OAI21_X1   g10500(.A1(new_n10128_), .A2(new_n10366_), .B(new_n10482_), .ZN(new_n10757_));
  NAND3_X1   g10501(.A1(new_n10740_), .A2(new_n10757_), .A3(new_n10504_), .ZN(new_n10758_));
  INV_X1     g10502(.I(new_n10504_), .ZN(new_n10759_));
  NOR3_X1    g10503(.A1(new_n10488_), .A2(new_n10483_), .A3(new_n10759_), .ZN(new_n10760_));
  AOI21_X1   g10504(.A1(new_n10740_), .A2(new_n10757_), .B(new_n10504_), .ZN(new_n10761_));
  NOR2_X1    g10505(.A1(new_n10761_), .A2(new_n10760_), .ZN(new_n10762_));
  NAND3_X1   g10506(.A1(new_n10365_), .A2(new_n10762_), .A3(new_n10363_), .ZN(new_n10763_));
  AOI21_X1   g10507(.A1(new_n10763_), .A2(new_n10758_), .B(new_n10756_), .ZN(new_n10764_));
  OAI21_X1   g10508(.A1(new_n10488_), .A2(new_n10483_), .B(new_n10759_), .ZN(new_n10765_));
  NAND2_X1   g10509(.A1(new_n10758_), .A2(new_n10765_), .ZN(new_n10766_));
  NOR3_X1    g10510(.A1(new_n10494_), .A2(new_n10766_), .A3(new_n10492_), .ZN(new_n10767_));
  NOR3_X1    g10511(.A1(new_n10767_), .A2(new_n10755_), .A3(new_n10760_), .ZN(new_n10768_));
  NOR3_X1    g10512(.A1(new_n10768_), .A2(new_n10764_), .A3(new_n10751_), .ZN(new_n10769_));
  AND2_X2    g10513(.A1(new_n10750_), .A2(new_n10746_), .Z(new_n10770_));
  OAI21_X1   g10514(.A1(new_n10767_), .A2(new_n10760_), .B(new_n10755_), .ZN(new_n10771_));
  NAND3_X1   g10515(.A1(new_n10763_), .A2(new_n10756_), .A3(new_n10758_), .ZN(new_n10772_));
  AOI21_X1   g10516(.A1(new_n10771_), .A2(new_n10772_), .B(new_n10770_), .ZN(new_n10773_));
  OR2_X2     g10517(.A1(new_n10773_), .A2(new_n10769_), .Z(new_n10774_));
  AOI22_X1   g10518(.A1(new_n3267_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n3270_), .ZN(new_n10775_));
  OAI21_X1   g10519(.A1(new_n3185_), .A2(new_n3475_), .B(new_n10775_), .ZN(new_n10776_));
  AOI21_X1   g10520(.A1(new_n4230_), .A2(new_n3273_), .B(new_n10776_), .ZN(new_n10777_));
  XOR2_X1    g10521(.A1(new_n10777_), .A2(new_n3264_), .Z(new_n10778_));
  AOI21_X1   g10522(.A1(new_n10363_), .A2(new_n10365_), .B(new_n10762_), .ZN(new_n10779_));
  NOR3_X1    g10523(.A1(new_n10779_), .A2(new_n10767_), .A3(new_n10500_), .ZN(new_n10780_));
  INV_X1     g10524(.I(new_n10780_), .ZN(new_n10781_));
  NAND2_X1   g10525(.A1(new_n10511_), .A2(new_n10781_), .ZN(new_n10782_));
  NAND2_X1   g10526(.A1(new_n10782_), .A2(new_n10778_), .ZN(new_n10783_));
  INV_X1     g10527(.I(new_n10778_), .ZN(new_n10784_));
  NOR2_X1    g10528(.A1(new_n10517_), .A2(new_n10780_), .ZN(new_n10785_));
  NAND2_X1   g10529(.A1(new_n10785_), .A2(new_n10784_), .ZN(new_n10786_));
  NAND2_X1   g10530(.A1(new_n10783_), .A2(new_n10786_), .ZN(new_n10787_));
  XOR2_X1    g10531(.A1(new_n10787_), .A2(new_n10774_), .Z(new_n10788_));
  AOI22_X1   g10532(.A1(new_n2716_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n2719_), .ZN(new_n10789_));
  OAI21_X1   g10533(.A1(new_n4022_), .A2(new_n2924_), .B(new_n10789_), .ZN(new_n10790_));
  AOI21_X1   g10534(.A1(new_n4223_), .A2(new_n2722_), .B(new_n10790_), .ZN(new_n10791_));
  XOR2_X1    g10535(.A1(new_n10791_), .A2(new_n2714_), .Z(new_n10792_));
  INV_X1     g10536(.I(new_n10792_), .ZN(new_n10793_));
  AOI21_X1   g10537(.A1(new_n10527_), .A2(new_n10515_), .B(new_n10793_), .ZN(new_n10794_));
  INV_X1     g10538(.I(new_n10794_), .ZN(new_n10795_));
  NAND3_X1   g10539(.A1(new_n10527_), .A2(new_n10515_), .A3(new_n10793_), .ZN(new_n10796_));
  AND3_X2    g10540(.A1(new_n10795_), .A2(new_n10788_), .A3(new_n10796_), .Z(new_n10797_));
  AOI21_X1   g10541(.A1(new_n10795_), .A2(new_n10796_), .B(new_n10788_), .ZN(new_n10798_));
  NOR2_X1    g10542(.A1(new_n10797_), .A2(new_n10798_), .ZN(new_n10799_));
  INV_X1     g10543(.I(new_n10799_), .ZN(new_n10800_));
  AOI22_X1   g10544(.A1(new_n2202_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n2205_), .ZN(new_n10801_));
  OAI21_X1   g10545(.A1(new_n4639_), .A2(new_n2370_), .B(new_n10801_), .ZN(new_n10802_));
  AOI21_X1   g10546(.A1(new_n5594_), .A2(new_n2208_), .B(new_n10802_), .ZN(new_n10803_));
  XOR2_X1    g10547(.A1(new_n10803_), .A2(new_n2200_), .Z(new_n10804_));
  INV_X1     g10548(.I(new_n10804_), .ZN(new_n10805_));
  NOR2_X1    g10549(.A1(new_n10531_), .A2(new_n10533_), .ZN(new_n10806_));
  NOR2_X1    g10550(.A1(new_n10806_), .A2(new_n10805_), .ZN(new_n10807_));
  NAND2_X1   g10551(.A1(new_n10537_), .A2(new_n10529_), .ZN(new_n10808_));
  NOR2_X1    g10552(.A1(new_n10808_), .A2(new_n10804_), .ZN(new_n10809_));
  NOR3_X1    g10553(.A1(new_n10809_), .A2(new_n10807_), .A3(new_n10800_), .ZN(new_n10810_));
  NAND2_X1   g10554(.A1(new_n10808_), .A2(new_n10804_), .ZN(new_n10811_));
  NAND2_X1   g10555(.A1(new_n10806_), .A2(new_n10805_), .ZN(new_n10812_));
  AOI21_X1   g10556(.A1(new_n10811_), .A2(new_n10812_), .B(new_n10799_), .ZN(new_n10813_));
  NOR2_X1    g10557(.A1(new_n10810_), .A2(new_n10813_), .ZN(new_n10814_));
  INV_X1     g10558(.I(new_n10814_), .ZN(new_n10815_));
  AOI22_X1   g10559(.A1(new_n1738_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n1743_), .ZN(new_n10816_));
  OAI21_X1   g10560(.A1(new_n5312_), .A2(new_n1931_), .B(new_n10816_), .ZN(new_n10817_));
  AOI21_X1   g10561(.A1(new_n6310_), .A2(new_n1746_), .B(new_n10817_), .ZN(new_n10818_));
  XOR2_X1    g10562(.A1(new_n10818_), .A2(new_n1736_), .Z(new_n10819_));
  INV_X1     g10563(.I(new_n10819_), .ZN(new_n10820_));
  AOI21_X1   g10564(.A1(new_n10550_), .A2(new_n10539_), .B(new_n10820_), .ZN(new_n10821_));
  NOR3_X1    g10565(.A1(new_n10543_), .A2(new_n10545_), .A3(new_n10819_), .ZN(new_n10822_));
  NOR3_X1    g10566(.A1(new_n10815_), .A2(new_n10822_), .A3(new_n10821_), .ZN(new_n10823_));
  OAI21_X1   g10567(.A1(new_n10543_), .A2(new_n10545_), .B(new_n10819_), .ZN(new_n10824_));
  NAND3_X1   g10568(.A1(new_n10550_), .A2(new_n10539_), .A3(new_n10820_), .ZN(new_n10825_));
  AOI21_X1   g10569(.A1(new_n10824_), .A2(new_n10825_), .B(new_n10814_), .ZN(new_n10826_));
  NOR2_X1    g10570(.A1(new_n10823_), .A2(new_n10826_), .ZN(new_n10827_));
  INV_X1     g10571(.I(new_n10827_), .ZN(new_n10828_));
  OAI22_X1   g10572(.A1(new_n1592_), .A2(new_n6490_), .B1(new_n6285_), .B2(new_n1505_), .ZN(new_n10829_));
  AOI21_X1   g10573(.A1(\b[40] ), .A2(new_n1584_), .B(new_n10829_), .ZN(new_n10830_));
  OAI21_X1   g10574(.A1(new_n8988_), .A2(new_n1732_), .B(new_n10830_), .ZN(new_n10831_));
  XOR2_X1    g10575(.A1(new_n10831_), .A2(\a[17] ), .Z(new_n10832_));
  OAI21_X1   g10576(.A1(new_n10554_), .A2(new_n10556_), .B(new_n10832_), .ZN(new_n10833_));
  INV_X1     g10577(.I(new_n10833_), .ZN(new_n10834_));
  NOR3_X1    g10578(.A1(new_n10554_), .A2(new_n10556_), .A3(new_n10832_), .ZN(new_n10835_));
  NOR3_X1    g10579(.A1(new_n10834_), .A2(new_n10828_), .A3(new_n10835_), .ZN(new_n10836_));
  INV_X1     g10580(.I(new_n10835_), .ZN(new_n10837_));
  AOI21_X1   g10581(.A1(new_n10837_), .A2(new_n10833_), .B(new_n10827_), .ZN(new_n10838_));
  NOR2_X1    g10582(.A1(new_n10838_), .A2(new_n10836_), .ZN(new_n10839_));
  OAI22_X1   g10583(.A1(new_n993_), .A2(new_n7096_), .B1(new_n7074_), .B2(new_n997_), .ZN(new_n10840_));
  AOI21_X1   g10584(.A1(\b[43] ), .A2(new_n1486_), .B(new_n10840_), .ZN(new_n10841_));
  OAI21_X1   g10585(.A1(new_n7925_), .A2(new_n1323_), .B(new_n10841_), .ZN(new_n10842_));
  XOR2_X1    g10586(.A1(new_n10842_), .A2(\a[14] ), .Z(new_n10843_));
  OAI21_X1   g10587(.A1(new_n10226_), .A2(new_n10221_), .B(new_n10220_), .ZN(new_n10844_));
  OAI21_X1   g10588(.A1(new_n10844_), .A2(new_n10574_), .B(new_n10572_), .ZN(new_n10845_));
  NAND2_X1   g10589(.A1(new_n10845_), .A2(new_n10843_), .ZN(new_n10846_));
  NOR2_X1    g10590(.A1(new_n10845_), .A2(new_n10843_), .ZN(new_n10847_));
  INV_X1     g10591(.I(new_n10847_), .ZN(new_n10848_));
  NAND3_X1   g10592(.A1(new_n10848_), .A2(new_n10839_), .A3(new_n10846_), .ZN(new_n10849_));
  OR2_X2     g10593(.A1(new_n10838_), .A2(new_n10836_), .Z(new_n10850_));
  INV_X1     g10594(.I(new_n10846_), .ZN(new_n10851_));
  OAI21_X1   g10595(.A1(new_n10851_), .A2(new_n10847_), .B(new_n10850_), .ZN(new_n10852_));
  NAND2_X1   g10596(.A1(new_n10852_), .A2(new_n10849_), .ZN(new_n10853_));
  OAI22_X1   g10597(.A1(new_n713_), .A2(new_n8127_), .B1(new_n8126_), .B2(new_n717_), .ZN(new_n10854_));
  AOI21_X1   g10598(.A1(\b[46] ), .A2(new_n1126_), .B(new_n10854_), .ZN(new_n10855_));
  OAI21_X1   g10599(.A1(new_n8138_), .A2(new_n986_), .B(new_n10855_), .ZN(new_n10856_));
  XOR2_X1    g10600(.A1(new_n10856_), .A2(\a[11] ), .Z(new_n10857_));
  INV_X1     g10601(.I(new_n10857_), .ZN(new_n10858_));
  OAI21_X1   g10602(.A1(new_n10583_), .A2(new_n10245_), .B(new_n10581_), .ZN(new_n10859_));
  AOI21_X1   g10603(.A1(new_n10564_), .A2(new_n10575_), .B(new_n10577_), .ZN(new_n10860_));
  INV_X1     g10604(.I(new_n10860_), .ZN(new_n10861_));
  AOI21_X1   g10605(.A1(new_n10859_), .A2(new_n10861_), .B(new_n10858_), .ZN(new_n10862_));
  AOI21_X1   g10606(.A1(new_n10327_), .A2(new_n10240_), .B(new_n10586_), .ZN(new_n10863_));
  NOR3_X1    g10607(.A1(new_n10863_), .A2(new_n10857_), .A3(new_n10860_), .ZN(new_n10864_));
  NOR3_X1    g10608(.A1(new_n10864_), .A2(new_n10862_), .A3(new_n10853_), .ZN(new_n10865_));
  NOR3_X1    g10609(.A1(new_n10851_), .A2(new_n10850_), .A3(new_n10847_), .ZN(new_n10866_));
  AOI21_X1   g10610(.A1(new_n10848_), .A2(new_n10846_), .B(new_n10839_), .ZN(new_n10867_));
  NOR2_X1    g10611(.A1(new_n10867_), .A2(new_n10866_), .ZN(new_n10868_));
  OAI21_X1   g10612(.A1(new_n10863_), .A2(new_n10860_), .B(new_n10857_), .ZN(new_n10869_));
  NAND3_X1   g10613(.A1(new_n10859_), .A2(new_n10858_), .A3(new_n10861_), .ZN(new_n10870_));
  AOI21_X1   g10614(.A1(new_n10869_), .A2(new_n10870_), .B(new_n10868_), .ZN(new_n10871_));
  OAI21_X1   g10615(.A1(new_n10865_), .A2(new_n10871_), .B(new_n10644_), .ZN(new_n10872_));
  NAND3_X1   g10616(.A1(new_n10869_), .A2(new_n10870_), .A3(new_n10868_), .ZN(new_n10873_));
  OAI21_X1   g10617(.A1(new_n10864_), .A2(new_n10862_), .B(new_n10853_), .ZN(new_n10874_));
  NAND3_X1   g10618(.A1(new_n10874_), .A2(new_n10873_), .A3(new_n10643_), .ZN(new_n10875_));
  NAND2_X1   g10619(.A1(new_n10872_), .A2(new_n10875_), .ZN(new_n10876_));
  NOR2_X1    g10620(.A1(new_n10876_), .A2(new_n10639_), .ZN(new_n10877_));
  INV_X1     g10621(.I(new_n10592_), .ZN(new_n10878_));
  OAI21_X1   g10622(.A1(new_n10594_), .A2(new_n10593_), .B(new_n10878_), .ZN(new_n10879_));
  AOI21_X1   g10623(.A1(new_n10874_), .A2(new_n10873_), .B(new_n10643_), .ZN(new_n10880_));
  NOR3_X1    g10624(.A1(new_n10865_), .A2(new_n10871_), .A3(new_n10644_), .ZN(new_n10881_));
  NOR2_X1    g10625(.A1(new_n10881_), .A2(new_n10880_), .ZN(new_n10882_));
  NOR2_X1    g10626(.A1(new_n10882_), .A2(new_n10879_), .ZN(new_n10883_));
  INV_X1     g10627(.I(new_n9952_), .ZN(new_n10884_));
  AOI22_X1   g10628(.A1(new_n800_), .A2(\b[53] ), .B1(\b[54] ), .B2(new_n333_), .ZN(new_n10885_));
  OAI21_X1   g10629(.A1(new_n9032_), .A2(new_n392_), .B(new_n10885_), .ZN(new_n10886_));
  AOI21_X1   g10630(.A1(new_n10884_), .A2(new_n330_), .B(new_n10886_), .ZN(new_n10887_));
  XOR2_X1    g10631(.A1(new_n10887_), .A2(new_n312_), .Z(new_n10888_));
  NOR3_X1    g10632(.A1(new_n10883_), .A2(new_n10877_), .A3(new_n10888_), .ZN(new_n10889_));
  NAND3_X1   g10633(.A1(new_n10879_), .A2(new_n10872_), .A3(new_n10875_), .ZN(new_n10890_));
  NAND2_X1   g10634(.A1(new_n10876_), .A2(new_n10639_), .ZN(new_n10891_));
  INV_X1     g10635(.I(new_n10888_), .ZN(new_n10892_));
  AOI21_X1   g10636(.A1(new_n10891_), .A2(new_n10890_), .B(new_n10892_), .ZN(new_n10893_));
  NOR2_X1    g10637(.A1(new_n10889_), .A2(new_n10893_), .ZN(new_n10894_));
  NOR3_X1    g10638(.A1(new_n10894_), .A2(new_n10636_), .A3(new_n10605_), .ZN(new_n10895_));
  AOI21_X1   g10639(.A1(new_n10284_), .A2(new_n10285_), .B(new_n10602_), .ZN(new_n10896_));
  OAI21_X1   g10640(.A1(new_n10896_), .A2(new_n10601_), .B(new_n10596_), .ZN(new_n10897_));
  NAND3_X1   g10641(.A1(new_n10891_), .A2(new_n10890_), .A3(new_n10892_), .ZN(new_n10898_));
  OAI21_X1   g10642(.A1(new_n10883_), .A2(new_n10877_), .B(new_n10888_), .ZN(new_n10899_));
  NAND2_X1   g10643(.A1(new_n10899_), .A2(new_n10898_), .ZN(new_n10900_));
  AOI21_X1   g10644(.A1(new_n10608_), .A2(new_n10897_), .B(new_n10900_), .ZN(new_n10901_));
  NOR3_X1    g10645(.A1(new_n10901_), .A2(new_n10895_), .A3(new_n10634_), .ZN(new_n10902_));
  XOR2_X1    g10646(.A1(new_n10633_), .A2(\a[2] ), .Z(new_n10903_));
  NAND3_X1   g10647(.A1(new_n10897_), .A2(new_n10900_), .A3(new_n10608_), .ZN(new_n10904_));
  OAI21_X1   g10648(.A1(new_n10605_), .A2(new_n10636_), .B(new_n10894_), .ZN(new_n10905_));
  AOI21_X1   g10649(.A1(new_n10905_), .A2(new_n10904_), .B(new_n10903_), .ZN(new_n10906_));
  NOR2_X1    g10650(.A1(new_n10906_), .A2(new_n10902_), .ZN(new_n10907_));
  XOR2_X1    g10651(.A1(new_n10907_), .A2(new_n10619_), .Z(\f[57] ));
  OAI21_X1   g10652(.A1(new_n10636_), .A2(new_n10605_), .B(new_n10899_), .ZN(new_n10909_));
  NAND2_X1   g10653(.A1(new_n10909_), .A2(new_n10898_), .ZN(new_n10910_));
  AOI22_X1   g10654(.A1(new_n800_), .A2(\b[54] ), .B1(\b[55] ), .B2(new_n333_), .ZN(new_n10911_));
  OAI21_X1   g10655(.A1(new_n9376_), .A2(new_n392_), .B(new_n10911_), .ZN(new_n10912_));
  AOI21_X1   g10656(.A1(new_n9979_), .A2(new_n330_), .B(new_n10912_), .ZN(new_n10913_));
  XOR2_X1    g10657(.A1(new_n10913_), .A2(new_n312_), .Z(new_n10914_));
  NOR2_X1    g10658(.A1(new_n10865_), .A2(new_n10871_), .ZN(new_n10915_));
  OAI21_X1   g10659(.A1(new_n10639_), .A2(new_n10644_), .B(new_n10915_), .ZN(new_n10916_));
  NAND2_X1   g10660(.A1(new_n10639_), .A2(new_n10644_), .ZN(new_n10917_));
  AOI22_X1   g10661(.A1(new_n518_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n636_), .ZN(new_n10918_));
  OAI21_X1   g10662(.A1(new_n8500_), .A2(new_n917_), .B(new_n10918_), .ZN(new_n10919_));
  AOI21_X1   g10663(.A1(new_n9987_), .A2(new_n618_), .B(new_n10919_), .ZN(new_n10920_));
  XOR2_X1    g10664(.A1(new_n10920_), .A2(new_n488_), .Z(new_n10921_));
  NAND2_X1   g10665(.A1(new_n10869_), .A2(new_n10868_), .ZN(new_n10922_));
  NAND2_X1   g10666(.A1(new_n10846_), .A2(new_n10839_), .ZN(new_n10923_));
  NAND2_X1   g10667(.A1(new_n10923_), .A2(new_n10848_), .ZN(new_n10924_));
  OAI22_X1   g10668(.A1(new_n993_), .A2(new_n7617_), .B1(new_n7096_), .B2(new_n997_), .ZN(new_n10925_));
  AOI21_X1   g10669(.A1(\b[44] ), .A2(new_n1486_), .B(new_n10925_), .ZN(new_n10926_));
  OAI21_X1   g10670(.A1(new_n7627_), .A2(new_n1323_), .B(new_n10926_), .ZN(new_n10927_));
  XOR2_X1    g10671(.A1(new_n10927_), .A2(\a[14] ), .Z(new_n10928_));
  INV_X1     g10672(.I(new_n10928_), .ZN(new_n10929_));
  NAND2_X1   g10673(.A1(new_n10560_), .A2(new_n10552_), .ZN(new_n10930_));
  AOI21_X1   g10674(.A1(new_n10930_), .A2(new_n10832_), .B(new_n10828_), .ZN(new_n10931_));
  OAI21_X1   g10675(.A1(new_n10815_), .A2(new_n10821_), .B(new_n10825_), .ZN(new_n10932_));
  NAND2_X1   g10676(.A1(new_n10811_), .A2(new_n10799_), .ZN(new_n10933_));
  NAND2_X1   g10677(.A1(new_n10933_), .A2(new_n10812_), .ZN(new_n10934_));
  INV_X1     g10678(.I(new_n10934_), .ZN(new_n10935_));
  NOR2_X1    g10679(.A1(new_n10932_), .A2(new_n10935_), .ZN(new_n10936_));
  AOI21_X1   g10680(.A1(new_n10814_), .A2(new_n10824_), .B(new_n10822_), .ZN(new_n10937_));
  NOR2_X1    g10681(.A1(new_n10937_), .A2(new_n10934_), .ZN(new_n10938_));
  AOI22_X1   g10682(.A1(new_n1738_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n1743_), .ZN(new_n10939_));
  OAI21_X1   g10683(.A1(new_n5341_), .A2(new_n1931_), .B(new_n10939_), .ZN(new_n10940_));
  AOI21_X1   g10684(.A1(new_n5793_), .A2(new_n1746_), .B(new_n10940_), .ZN(new_n10941_));
  XOR2_X1    g10685(.A1(new_n10941_), .A2(new_n1736_), .Z(new_n10942_));
  INV_X1     g10686(.I(new_n10942_), .ZN(new_n10943_));
  OAI22_X1   g10687(.A1(new_n2189_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n2194_), .ZN(new_n10944_));
  AOI21_X1   g10688(.A1(\b[35] ), .A2(new_n2361_), .B(new_n10944_), .ZN(new_n10945_));
  OAI21_X1   g10689(.A1(new_n5322_), .A2(new_n2197_), .B(new_n10945_), .ZN(new_n10946_));
  XOR2_X1    g10690(.A1(new_n10946_), .A2(\a[23] ), .Z(new_n10947_));
  NAND2_X1   g10691(.A1(new_n10795_), .A2(new_n10788_), .ZN(new_n10948_));
  AOI22_X1   g10692(.A1(new_n2716_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n2719_), .ZN(new_n10949_));
  OAI21_X1   g10693(.A1(new_n4023_), .A2(new_n2924_), .B(new_n10949_), .ZN(new_n10950_));
  AOI21_X1   g10694(.A1(new_n5103_), .A2(new_n2722_), .B(new_n10950_), .ZN(new_n10951_));
  XOR2_X1    g10695(.A1(new_n10951_), .A2(new_n2714_), .Z(new_n10952_));
  NOR2_X1    g10696(.A1(new_n10773_), .A2(new_n10769_), .ZN(new_n10953_));
  OAI21_X1   g10697(.A1(new_n10785_), .A2(new_n10784_), .B(new_n10953_), .ZN(new_n10954_));
  NAND2_X1   g10698(.A1(new_n10954_), .A2(new_n10786_), .ZN(new_n10955_));
  OAI21_X1   g10699(.A1(new_n10751_), .A2(new_n10764_), .B(new_n10772_), .ZN(new_n10956_));
  AOI22_X1   g10700(.A1(new_n5155_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n5160_), .ZN(new_n10957_));
  OAI21_X1   g10701(.A1(new_n1860_), .A2(new_n6877_), .B(new_n10957_), .ZN(new_n10958_));
  AOI21_X1   g10702(.A1(new_n2659_), .A2(new_n5166_), .B(new_n10958_), .ZN(new_n10959_));
  XOR2_X1    g10703(.A1(new_n10959_), .A2(new_n5162_), .Z(new_n10960_));
  NAND2_X1   g10704(.A1(new_n10718_), .A2(new_n10711_), .ZN(new_n10961_));
  NAND2_X1   g10705(.A1(new_n10961_), .A2(new_n10713_), .ZN(new_n10962_));
  INV_X1     g10706(.I(new_n10702_), .ZN(new_n10963_));
  AOI21_X1   g10707(.A1(new_n10696_), .A2(new_n10699_), .B(new_n10691_), .ZN(new_n10964_));
  NOR2_X1    g10708(.A1(new_n10964_), .A2(new_n10963_), .ZN(new_n10965_));
  NOR2_X1    g10709(.A1(new_n10688_), .A2(new_n10681_), .ZN(new_n10966_));
  NOR2_X1    g10710(.A1(new_n10966_), .A2(new_n10689_), .ZN(new_n10967_));
  INV_X1     g10711(.I(new_n10967_), .ZN(new_n10968_));
  OAI21_X1   g10712(.A1(new_n10657_), .A2(new_n10678_), .B(new_n10677_), .ZN(new_n10969_));
  NAND2_X1   g10713(.A1(new_n10674_), .A2(new_n10402_), .ZN(new_n10970_));
  NAND2_X1   g10714(.A1(new_n10970_), .A2(new_n10673_), .ZN(new_n10971_));
  AOI22_X1   g10715(.A1(new_n10064_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n10062_), .ZN(new_n10972_));
  OAI21_X1   g10716(.A1(new_n276_), .A2(new_n10399_), .B(new_n10972_), .ZN(new_n10973_));
  AOI21_X1   g10717(.A1(new_n1725_), .A2(new_n10068_), .B(new_n10973_), .ZN(new_n10974_));
  XOR2_X1    g10718(.A1(new_n10974_), .A2(new_n10057_), .Z(new_n10975_));
  INV_X1     g10719(.I(\a[58] ), .ZN(new_n10976_));
  OR3_X2     g10720(.A1(new_n10976_), .A2(\a[56] ), .A3(\a[57] ), .Z(new_n10977_));
  NAND3_X1   g10721(.A1(new_n10976_), .A2(\a[56] ), .A3(\a[57] ), .ZN(new_n10978_));
  NAND2_X1   g10722(.A1(new_n10977_), .A2(new_n10978_), .ZN(new_n10979_));
  XOR2_X1    g10723(.A1(\a[58] ), .A2(\a[59] ), .Z(new_n10980_));
  NOR2_X1    g10724(.A1(new_n10670_), .A2(new_n10980_), .ZN(new_n10981_));
  AOI22_X1   g10725(.A1(new_n10981_), .A2(\b[1] ), .B1(new_n10979_), .B2(\b[0] ), .ZN(new_n10982_));
  XNOR2_X1   g10726(.A1(\a[58] ), .A2(\a[59] ), .ZN(new_n10983_));
  NOR2_X1    g10727(.A1(new_n10670_), .A2(new_n10983_), .ZN(new_n10984_));
  INV_X1     g10728(.I(new_n10984_), .ZN(new_n10985_));
  OAI21_X1   g10729(.A1(new_n313_), .A2(new_n10985_), .B(new_n10982_), .ZN(new_n10986_));
  XOR2_X1    g10730(.A1(new_n10986_), .A2(\a[59] ), .Z(new_n10987_));
  NAND3_X1   g10731(.A1(new_n10987_), .A2(\a[59] ), .A3(new_n10672_), .ZN(new_n10988_));
  INV_X1     g10732(.I(\a[59] ), .ZN(new_n10989_));
  INV_X1     g10733(.I(new_n10987_), .ZN(new_n10990_));
  OAI21_X1   g10734(.A1(new_n10989_), .A2(new_n10671_), .B(new_n10990_), .ZN(new_n10991_));
  NAND3_X1   g10735(.A1(new_n10991_), .A2(new_n10975_), .A3(new_n10988_), .ZN(new_n10992_));
  INV_X1     g10736(.I(new_n10975_), .ZN(new_n10993_));
  NAND2_X1   g10737(.A1(new_n10991_), .A2(new_n10988_), .ZN(new_n10994_));
  NAND2_X1   g10738(.A1(new_n10994_), .A2(new_n10993_), .ZN(new_n10995_));
  NAND2_X1   g10739(.A1(new_n10995_), .A2(new_n10992_), .ZN(new_n10996_));
  XNOR2_X1   g10740(.A1(new_n10996_), .A2(new_n10971_), .ZN(new_n10997_));
  OAI22_X1   g10741(.A1(new_n10390_), .A2(new_n471_), .B1(new_n438_), .B2(new_n10389_), .ZN(new_n10998_));
  AOI21_X1   g10742(.A1(\b[5] ), .A2(new_n9471_), .B(new_n10998_), .ZN(new_n10999_));
  OAI21_X1   g10743(.A1(new_n485_), .A2(new_n10388_), .B(new_n10999_), .ZN(new_n11000_));
  XOR2_X1    g10744(.A1(new_n11000_), .A2(\a[53] ), .Z(new_n11001_));
  OR2_X2     g10745(.A1(new_n10997_), .A2(new_n11001_), .Z(new_n11002_));
  NAND2_X1   g10746(.A1(new_n10997_), .A2(new_n11001_), .ZN(new_n11003_));
  NAND2_X1   g10747(.A1(new_n11002_), .A2(new_n11003_), .ZN(new_n11004_));
  XNOR2_X1   g10748(.A1(new_n11004_), .A2(new_n10969_), .ZN(new_n11005_));
  INV_X1     g10749(.I(new_n11005_), .ZN(new_n11006_));
  AOI22_X1   g10750(.A1(new_n8241_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n8246_), .ZN(new_n11007_));
  OAI21_X1   g10751(.A1(new_n577_), .A2(new_n9114_), .B(new_n11007_), .ZN(new_n11008_));
  AOI21_X1   g10752(.A1(new_n1059_), .A2(new_n8252_), .B(new_n11008_), .ZN(new_n11009_));
  XOR2_X1    g10753(.A1(new_n11009_), .A2(new_n8248_), .Z(new_n11010_));
  NOR2_X1    g10754(.A1(new_n11006_), .A2(new_n11010_), .ZN(new_n11011_));
  NAND2_X1   g10755(.A1(new_n11006_), .A2(new_n11010_), .ZN(new_n11012_));
  INV_X1     g10756(.I(new_n11012_), .ZN(new_n11013_));
  NOR2_X1    g10757(.A1(new_n11013_), .A2(new_n11011_), .ZN(new_n11014_));
  NAND2_X1   g10758(.A1(new_n10968_), .A2(new_n11014_), .ZN(new_n11015_));
  INV_X1     g10759(.I(new_n11011_), .ZN(new_n11016_));
  NAND2_X1   g10760(.A1(new_n11016_), .A2(new_n11012_), .ZN(new_n11017_));
  NAND2_X1   g10761(.A1(new_n11017_), .A2(new_n10967_), .ZN(new_n11018_));
  OAI22_X1   g10762(.A1(new_n941_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n1070_), .ZN(new_n11019_));
  AOI21_X1   g10763(.A1(\b[11] ), .A2(new_n7719_), .B(new_n11019_), .ZN(new_n11020_));
  OAI21_X1   g10764(.A1(new_n1082_), .A2(new_n8585_), .B(new_n11020_), .ZN(new_n11021_));
  XOR2_X1    g10765(.A1(new_n11021_), .A2(\a[47] ), .Z(new_n11022_));
  INV_X1     g10766(.I(new_n11022_), .ZN(new_n11023_));
  NAND3_X1   g10767(.A1(new_n11015_), .A2(new_n11018_), .A3(new_n11023_), .ZN(new_n11024_));
  NOR2_X1    g10768(.A1(new_n11017_), .A2(new_n10967_), .ZN(new_n11025_));
  INV_X1     g10769(.I(new_n11018_), .ZN(new_n11026_));
  OAI21_X1   g10770(.A1(new_n11026_), .A2(new_n11025_), .B(new_n11022_), .ZN(new_n11027_));
  AOI21_X1   g10771(.A1(new_n11024_), .A2(new_n11027_), .B(new_n10965_), .ZN(new_n11028_));
  INV_X1     g10772(.I(new_n11024_), .ZN(new_n11029_));
  AOI21_X1   g10773(.A1(new_n11015_), .A2(new_n11018_), .B(new_n11023_), .ZN(new_n11030_));
  NOR4_X1    g10774(.A1(new_n10964_), .A2(new_n10963_), .A3(new_n11029_), .A4(new_n11030_), .ZN(new_n11031_));
  AOI22_X1   g10775(.A1(new_n6569_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n6574_), .ZN(new_n11032_));
  OAI21_X1   g10776(.A1(new_n1093_), .A2(new_n8565_), .B(new_n11032_), .ZN(new_n11033_));
  AOI21_X1   g10777(.A1(new_n1701_), .A2(new_n6579_), .B(new_n11033_), .ZN(new_n11034_));
  XOR2_X1    g10778(.A1(new_n11034_), .A2(new_n6567_), .Z(new_n11035_));
  INV_X1     g10779(.I(new_n11035_), .ZN(new_n11036_));
  OAI21_X1   g10780(.A1(new_n11028_), .A2(new_n11031_), .B(new_n11036_), .ZN(new_n11037_));
  INV_X1     g10781(.I(new_n11037_), .ZN(new_n11038_));
  NOR3_X1    g10782(.A1(new_n11028_), .A2(new_n11031_), .A3(new_n11036_), .ZN(new_n11039_));
  NOR2_X1    g10783(.A1(new_n11038_), .A2(new_n11039_), .ZN(new_n11040_));
  XOR2_X1    g10784(.A1(new_n11040_), .A2(new_n10962_), .Z(new_n11041_));
  INV_X1     g10785(.I(new_n11041_), .ZN(new_n11042_));
  AOI22_X1   g10786(.A1(new_n6108_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n6111_), .ZN(new_n11043_));
  OAI21_X1   g10787(.A1(new_n1432_), .A2(new_n7708_), .B(new_n11043_), .ZN(new_n11044_));
  AOI21_X1   g10788(.A1(new_n1695_), .A2(new_n6105_), .B(new_n11044_), .ZN(new_n11045_));
  XOR2_X1    g10789(.A1(new_n11045_), .A2(new_n5849_), .Z(new_n11046_));
  INV_X1     g10790(.I(new_n11046_), .ZN(new_n11047_));
  AOI21_X1   g10791(.A1(new_n10731_), .A2(new_n10721_), .B(new_n11047_), .ZN(new_n11048_));
  NOR3_X1    g10792(.A1(new_n10724_), .A2(new_n10726_), .A3(new_n11046_), .ZN(new_n11049_));
  NOR3_X1    g10793(.A1(new_n11049_), .A2(new_n11048_), .A3(new_n11042_), .ZN(new_n11050_));
  OAI21_X1   g10794(.A1(new_n10724_), .A2(new_n10726_), .B(new_n11046_), .ZN(new_n11051_));
  NAND3_X1   g10795(.A1(new_n10731_), .A2(new_n10721_), .A3(new_n11047_), .ZN(new_n11052_));
  AOI21_X1   g10796(.A1(new_n11051_), .A2(new_n11052_), .B(new_n11041_), .ZN(new_n11053_));
  NOR3_X1    g10797(.A1(new_n11050_), .A2(new_n11053_), .A3(new_n10960_), .ZN(new_n11054_));
  INV_X1     g10798(.I(new_n10960_), .ZN(new_n11055_));
  NAND3_X1   g10799(.A1(new_n11051_), .A2(new_n11052_), .A3(new_n11041_), .ZN(new_n11056_));
  OAI21_X1   g10800(.A1(new_n11049_), .A2(new_n11048_), .B(new_n11042_), .ZN(new_n11057_));
  AOI21_X1   g10801(.A1(new_n11057_), .A2(new_n11056_), .B(new_n11055_), .ZN(new_n11058_));
  NOR2_X1    g10802(.A1(new_n11054_), .A2(new_n11058_), .ZN(new_n11059_));
  NAND2_X1   g10803(.A1(new_n10646_), .A2(new_n10733_), .ZN(new_n11060_));
  NAND2_X1   g10804(.A1(new_n11060_), .A2(new_n10730_), .ZN(new_n11061_));
  OAI22_X1   g10805(.A1(new_n2646_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n2495_), .ZN(new_n11062_));
  AOI21_X1   g10806(.A1(\b[23] ), .A2(new_n4706_), .B(new_n11062_), .ZN(new_n11063_));
  OAI21_X1   g10807(.A1(new_n2655_), .A2(new_n4458_), .B(new_n11063_), .ZN(new_n11064_));
  XOR2_X1    g10808(.A1(new_n11064_), .A2(\a[35] ), .Z(new_n11065_));
  NOR2_X1    g10809(.A1(new_n11061_), .A2(new_n11065_), .ZN(new_n11066_));
  NAND2_X1   g10810(.A1(new_n11061_), .A2(new_n11065_), .ZN(new_n11067_));
  INV_X1     g10811(.I(new_n11067_), .ZN(new_n11068_));
  OAI21_X1   g10812(.A1(new_n11068_), .A2(new_n11066_), .B(new_n11059_), .ZN(new_n11069_));
  INV_X1     g10813(.I(new_n11069_), .ZN(new_n11070_));
  NOR3_X1    g10814(.A1(new_n11068_), .A2(new_n11059_), .A3(new_n11066_), .ZN(new_n11071_));
  NOR2_X1    g10815(.A1(new_n11070_), .A2(new_n11071_), .ZN(new_n11072_));
  OAI21_X1   g10816(.A1(new_n10744_), .A2(new_n10743_), .B(new_n10735_), .ZN(new_n11073_));
  AOI22_X1   g10817(.A1(new_n3864_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n3869_), .ZN(new_n11074_));
  OAI21_X1   g10818(.A1(new_n3006_), .A2(new_n5410_), .B(new_n11074_), .ZN(new_n11075_));
  AOI21_X1   g10819(.A1(new_n3807_), .A2(new_n3872_), .B(new_n11075_), .ZN(new_n11076_));
  XOR2_X1    g10820(.A1(new_n11076_), .A2(new_n3876_), .Z(new_n11077_));
  INV_X1     g10821(.I(new_n11077_), .ZN(new_n11078_));
  NAND3_X1   g10822(.A1(new_n11073_), .A2(new_n10745_), .A3(new_n11078_), .ZN(new_n11079_));
  INV_X1     g10823(.I(new_n11079_), .ZN(new_n11080_));
  AOI21_X1   g10824(.A1(new_n11073_), .A2(new_n10745_), .B(new_n11078_), .ZN(new_n11081_));
  OAI21_X1   g10825(.A1(new_n11080_), .A2(new_n11081_), .B(new_n11072_), .ZN(new_n11082_));
  OR3_X2     g10826(.A1(new_n11068_), .A2(new_n11059_), .A3(new_n11066_), .Z(new_n11083_));
  NAND2_X1   g10827(.A1(new_n11083_), .A2(new_n11069_), .ZN(new_n11084_));
  AOI21_X1   g10828(.A1(new_n10741_), .A2(new_n10739_), .B(new_n10747_), .ZN(new_n11085_));
  OAI21_X1   g10829(.A1(new_n11085_), .A2(new_n10749_), .B(new_n11077_), .ZN(new_n11086_));
  NAND3_X1   g10830(.A1(new_n11084_), .A2(new_n11079_), .A3(new_n11086_), .ZN(new_n11087_));
  NAND2_X1   g10831(.A1(new_n11082_), .A2(new_n11087_), .ZN(new_n11088_));
  NAND2_X1   g10832(.A1(new_n10956_), .A2(new_n11088_), .ZN(new_n11089_));
  AOI21_X1   g10833(.A1(new_n10770_), .A2(new_n10771_), .B(new_n10768_), .ZN(new_n11090_));
  AOI21_X1   g10834(.A1(new_n11086_), .A2(new_n11079_), .B(new_n11084_), .ZN(new_n11091_));
  NOR3_X1    g10835(.A1(new_n11080_), .A2(new_n11072_), .A3(new_n11081_), .ZN(new_n11092_));
  NOR2_X1    g10836(.A1(new_n11092_), .A2(new_n11091_), .ZN(new_n11093_));
  NAND2_X1   g10837(.A1(new_n11090_), .A2(new_n11093_), .ZN(new_n11094_));
  AOI22_X1   g10838(.A1(new_n3267_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n3270_), .ZN(new_n11095_));
  OAI21_X1   g10839(.A1(new_n3592_), .A2(new_n3475_), .B(new_n11095_), .ZN(new_n11096_));
  AOI21_X1   g10840(.A1(new_n3796_), .A2(new_n3273_), .B(new_n11096_), .ZN(new_n11097_));
  XOR2_X1    g10841(.A1(new_n11097_), .A2(new_n3264_), .Z(new_n11098_));
  AOI21_X1   g10842(.A1(new_n11094_), .A2(new_n11089_), .B(new_n11098_), .ZN(new_n11099_));
  NOR2_X1    g10843(.A1(new_n11090_), .A2(new_n11093_), .ZN(new_n11100_));
  NOR2_X1    g10844(.A1(new_n10956_), .A2(new_n11088_), .ZN(new_n11101_));
  INV_X1     g10845(.I(new_n11098_), .ZN(new_n11102_));
  NOR3_X1    g10846(.A1(new_n11100_), .A2(new_n11101_), .A3(new_n11102_), .ZN(new_n11103_));
  NOR2_X1    g10847(.A1(new_n11099_), .A2(new_n11103_), .ZN(new_n11104_));
  NAND2_X1   g10848(.A1(new_n10955_), .A2(new_n11104_), .ZN(new_n11105_));
  OAI21_X1   g10849(.A1(new_n11100_), .A2(new_n11101_), .B(new_n11102_), .ZN(new_n11106_));
  NAND3_X1   g10850(.A1(new_n11094_), .A2(new_n11089_), .A3(new_n11098_), .ZN(new_n11107_));
  NAND2_X1   g10851(.A1(new_n11106_), .A2(new_n11107_), .ZN(new_n11108_));
  NAND3_X1   g10852(.A1(new_n11108_), .A2(new_n10954_), .A3(new_n10786_), .ZN(new_n11109_));
  NAND3_X1   g10853(.A1(new_n11105_), .A2(new_n10952_), .A3(new_n11109_), .ZN(new_n11110_));
  INV_X1     g10854(.I(new_n10952_), .ZN(new_n11111_));
  AOI21_X1   g10855(.A1(new_n10786_), .A2(new_n10954_), .B(new_n11108_), .ZN(new_n11112_));
  NOR2_X1    g10856(.A1(new_n10782_), .A2(new_n10778_), .ZN(new_n11113_));
  AOI21_X1   g10857(.A1(new_n10782_), .A2(new_n10778_), .B(new_n10774_), .ZN(new_n11114_));
  NOR3_X1    g10858(.A1(new_n11104_), .A2(new_n11114_), .A3(new_n11113_), .ZN(new_n11115_));
  OAI21_X1   g10859(.A1(new_n11112_), .A2(new_n11115_), .B(new_n11111_), .ZN(new_n11116_));
  NAND2_X1   g10860(.A1(new_n11110_), .A2(new_n11116_), .ZN(new_n11117_));
  NAND3_X1   g10861(.A1(new_n10948_), .A2(new_n10796_), .A3(new_n11117_), .ZN(new_n11118_));
  XOR2_X1    g10862(.A1(new_n10787_), .A2(new_n10953_), .Z(new_n11119_));
  OAI21_X1   g10863(.A1(new_n11119_), .A2(new_n10794_), .B(new_n10796_), .ZN(new_n11120_));
  NOR3_X1    g10864(.A1(new_n11112_), .A2(new_n11115_), .A3(new_n11111_), .ZN(new_n11121_));
  AOI21_X1   g10865(.A1(new_n11105_), .A2(new_n11109_), .B(new_n10952_), .ZN(new_n11122_));
  NOR2_X1    g10866(.A1(new_n11122_), .A2(new_n11121_), .ZN(new_n11123_));
  NAND2_X1   g10867(.A1(new_n11120_), .A2(new_n11123_), .ZN(new_n11124_));
  NAND3_X1   g10868(.A1(new_n11118_), .A2(new_n11124_), .A3(new_n10947_), .ZN(new_n11125_));
  INV_X1     g10869(.I(new_n10947_), .ZN(new_n11126_));
  NOR2_X1    g10870(.A1(new_n11120_), .A2(new_n11123_), .ZN(new_n11127_));
  AOI21_X1   g10871(.A1(new_n10948_), .A2(new_n10796_), .B(new_n11117_), .ZN(new_n11128_));
  OAI21_X1   g10872(.A1(new_n11128_), .A2(new_n11127_), .B(new_n11126_), .ZN(new_n11129_));
  NAND2_X1   g10873(.A1(new_n11129_), .A2(new_n11125_), .ZN(new_n11130_));
  XOR2_X1    g10874(.A1(new_n11130_), .A2(new_n10943_), .Z(new_n11131_));
  INV_X1     g10875(.I(new_n11131_), .ZN(new_n11132_));
  NOR3_X1    g10876(.A1(new_n10938_), .A2(new_n10936_), .A3(new_n11132_), .ZN(new_n11133_));
  NAND2_X1   g10877(.A1(new_n10824_), .A2(new_n10814_), .ZN(new_n11134_));
  NAND3_X1   g10878(.A1(new_n11134_), .A2(new_n10825_), .A3(new_n10934_), .ZN(new_n11135_));
  NAND2_X1   g10879(.A1(new_n10932_), .A2(new_n10935_), .ZN(new_n11136_));
  AOI21_X1   g10880(.A1(new_n11136_), .A2(new_n11135_), .B(new_n11131_), .ZN(new_n11137_));
  OAI22_X1   g10881(.A1(new_n1592_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n1505_), .ZN(new_n11138_));
  AOI21_X1   g10882(.A1(\b[41] ), .A2(new_n1584_), .B(new_n11138_), .ZN(new_n11139_));
  OAI21_X1   g10883(.A1(new_n6785_), .A2(new_n1732_), .B(new_n11139_), .ZN(new_n11140_));
  XOR2_X1    g10884(.A1(new_n11140_), .A2(\a[17] ), .Z(new_n11141_));
  NOR3_X1    g10885(.A1(new_n11133_), .A2(new_n11137_), .A3(new_n11141_), .ZN(new_n11142_));
  NAND3_X1   g10886(.A1(new_n11136_), .A2(new_n11135_), .A3(new_n11131_), .ZN(new_n11143_));
  INV_X1     g10887(.I(new_n11137_), .ZN(new_n11144_));
  INV_X1     g10888(.I(new_n11141_), .ZN(new_n11145_));
  AOI21_X1   g10889(.A1(new_n11144_), .A2(new_n11143_), .B(new_n11145_), .ZN(new_n11146_));
  NOR4_X1    g10890(.A1(new_n11146_), .A2(new_n10835_), .A3(new_n10931_), .A4(new_n11142_), .ZN(new_n11147_));
  AOI21_X1   g10891(.A1(new_n10827_), .A2(new_n10833_), .B(new_n10835_), .ZN(new_n11148_));
  NAND3_X1   g10892(.A1(new_n11144_), .A2(new_n11143_), .A3(new_n11145_), .ZN(new_n11149_));
  OAI21_X1   g10893(.A1(new_n11133_), .A2(new_n11137_), .B(new_n11141_), .ZN(new_n11150_));
  AOI21_X1   g10894(.A1(new_n11149_), .A2(new_n11150_), .B(new_n11148_), .ZN(new_n11151_));
  OAI21_X1   g10895(.A1(new_n11147_), .A2(new_n11151_), .B(new_n10929_), .ZN(new_n11152_));
  NAND3_X1   g10896(.A1(new_n11149_), .A2(new_n11148_), .A3(new_n11150_), .ZN(new_n11153_));
  OAI22_X1   g10897(.A1(new_n11146_), .A2(new_n11142_), .B1(new_n10835_), .B2(new_n10931_), .ZN(new_n11154_));
  NAND3_X1   g10898(.A1(new_n11154_), .A2(new_n11153_), .A3(new_n10928_), .ZN(new_n11155_));
  NAND2_X1   g10899(.A1(new_n11152_), .A2(new_n11155_), .ZN(new_n11156_));
  INV_X1     g10900(.I(new_n11156_), .ZN(new_n11157_));
  NAND2_X1   g10901(.A1(new_n10924_), .A2(new_n11157_), .ZN(new_n11158_));
  NAND3_X1   g10902(.A1(new_n11156_), .A2(new_n10923_), .A3(new_n10848_), .ZN(new_n11159_));
  OAI22_X1   g10903(.A1(new_n713_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n717_), .ZN(new_n11160_));
  AOI21_X1   g10904(.A1(\b[47] ), .A2(new_n1126_), .B(new_n11160_), .ZN(new_n11161_));
  OAI21_X1   g10905(.A1(new_n9050_), .A2(new_n986_), .B(new_n11161_), .ZN(new_n11162_));
  XOR2_X1    g10906(.A1(new_n11162_), .A2(\a[11] ), .Z(new_n11163_));
  INV_X1     g10907(.I(new_n11163_), .ZN(new_n11164_));
  NAND3_X1   g10908(.A1(new_n11158_), .A2(new_n11159_), .A3(new_n11164_), .ZN(new_n11165_));
  AOI21_X1   g10909(.A1(new_n10923_), .A2(new_n10848_), .B(new_n11156_), .ZN(new_n11166_));
  INV_X1     g10910(.I(new_n11159_), .ZN(new_n11167_));
  OAI21_X1   g10911(.A1(new_n11167_), .A2(new_n11166_), .B(new_n11163_), .ZN(new_n11168_));
  NAND2_X1   g10912(.A1(new_n11168_), .A2(new_n11165_), .ZN(new_n11169_));
  AOI21_X1   g10913(.A1(new_n10870_), .A2(new_n10922_), .B(new_n11169_), .ZN(new_n11170_));
  NAND2_X1   g10914(.A1(new_n10922_), .A2(new_n10870_), .ZN(new_n11171_));
  NOR3_X1    g10915(.A1(new_n11167_), .A2(new_n11166_), .A3(new_n11163_), .ZN(new_n11172_));
  AOI21_X1   g10916(.A1(new_n11158_), .A2(new_n11159_), .B(new_n11164_), .ZN(new_n11173_));
  NOR2_X1    g10917(.A1(new_n11172_), .A2(new_n11173_), .ZN(new_n11174_));
  NOR2_X1    g10918(.A1(new_n11171_), .A2(new_n11174_), .ZN(new_n11175_));
  OAI21_X1   g10919(.A1(new_n11170_), .A2(new_n11175_), .B(new_n10921_), .ZN(new_n11176_));
  INV_X1     g10920(.I(new_n10921_), .ZN(new_n11177_));
  NAND2_X1   g10921(.A1(new_n11171_), .A2(new_n11174_), .ZN(new_n11178_));
  NAND3_X1   g10922(.A1(new_n11169_), .A2(new_n10922_), .A3(new_n10870_), .ZN(new_n11179_));
  NAND3_X1   g10923(.A1(new_n11178_), .A2(new_n11179_), .A3(new_n11177_), .ZN(new_n11180_));
  NAND2_X1   g10924(.A1(new_n11176_), .A2(new_n11180_), .ZN(new_n11181_));
  AOI21_X1   g10925(.A1(new_n10916_), .A2(new_n10917_), .B(new_n11181_), .ZN(new_n11182_));
  NAND2_X1   g10926(.A1(new_n10916_), .A2(new_n10917_), .ZN(new_n11183_));
  AOI21_X1   g10927(.A1(new_n11178_), .A2(new_n11179_), .B(new_n11177_), .ZN(new_n11184_));
  NOR3_X1    g10928(.A1(new_n11170_), .A2(new_n11175_), .A3(new_n10921_), .ZN(new_n11185_));
  NOR2_X1    g10929(.A1(new_n11185_), .A2(new_n11184_), .ZN(new_n11186_));
  NOR2_X1    g10930(.A1(new_n11183_), .A2(new_n11186_), .ZN(new_n11187_));
  OAI21_X1   g10931(.A1(new_n11182_), .A2(new_n11187_), .B(new_n10914_), .ZN(new_n11188_));
  INV_X1     g10932(.I(new_n10914_), .ZN(new_n11189_));
  NAND2_X1   g10933(.A1(new_n11183_), .A2(new_n11186_), .ZN(new_n11190_));
  NAND3_X1   g10934(.A1(new_n11181_), .A2(new_n10916_), .A3(new_n10917_), .ZN(new_n11191_));
  NAND3_X1   g10935(.A1(new_n11190_), .A2(new_n11191_), .A3(new_n11189_), .ZN(new_n11192_));
  NAND2_X1   g10936(.A1(new_n11188_), .A2(new_n11192_), .ZN(new_n11193_));
  XOR2_X1    g10937(.A1(new_n10910_), .A2(new_n11193_), .Z(new_n11194_));
  INV_X1     g10938(.I(\b[58] ), .ZN(new_n11195_));
  OAI22_X1   g10939(.A1(new_n277_), .A2(new_n11195_), .B1(new_n10625_), .B2(new_n262_), .ZN(new_n11196_));
  AOI21_X1   g10940(.A1(\b[56] ), .A2(new_n283_), .B(new_n11196_), .ZN(new_n11197_));
  AOI21_X1   g10941(.A1(new_n10626_), .A2(\b[56] ), .B(\b[55] ), .ZN(new_n11198_));
  AOI21_X1   g10942(.A1(new_n10315_), .A2(\b[57] ), .B(\b[56] ), .ZN(new_n11199_));
  NOR2_X1    g10943(.A1(new_n11198_), .A2(new_n11199_), .ZN(new_n11200_));
  XNOR2_X1   g10944(.A1(\b[57] ), .A2(\b[58] ), .ZN(new_n11201_));
  NOR2_X1    g10945(.A1(new_n11200_), .A2(new_n11201_), .ZN(new_n11202_));
  INV_X1     g10946(.I(new_n11200_), .ZN(new_n11203_));
  XOR2_X1    g10947(.A1(\b[57] ), .A2(\b[58] ), .Z(new_n11204_));
  NOR2_X1    g10948(.A1(new_n11203_), .A2(new_n11204_), .ZN(new_n11205_));
  NOR2_X1    g10949(.A1(new_n11205_), .A2(new_n11202_), .ZN(new_n11206_));
  OAI21_X1   g10950(.A1(new_n11206_), .A2(new_n279_), .B(new_n11197_), .ZN(new_n11207_));
  XOR2_X1    g10951(.A1(new_n11207_), .A2(\a[2] ), .Z(new_n11208_));
  INV_X1     g10952(.I(new_n11208_), .ZN(new_n11209_));
  AOI21_X1   g10953(.A1(new_n10612_), .A2(new_n10611_), .B(new_n10321_), .ZN(new_n11210_));
  OAI21_X1   g10954(.A1(new_n10307_), .A2(new_n11210_), .B(new_n10613_), .ZN(new_n11211_));
  NAND3_X1   g10955(.A1(new_n10905_), .A2(new_n10904_), .A3(new_n10903_), .ZN(new_n11212_));
  OAI21_X1   g10956(.A1(new_n10901_), .A2(new_n10895_), .B(new_n10634_), .ZN(new_n11213_));
  NAND2_X1   g10957(.A1(new_n11212_), .A2(new_n11213_), .ZN(new_n11214_));
  AOI21_X1   g10958(.A1(new_n10905_), .A2(new_n10904_), .B(new_n10634_), .ZN(new_n11215_));
  AOI21_X1   g10959(.A1(new_n11214_), .A2(new_n11211_), .B(new_n11215_), .ZN(new_n11216_));
  NOR2_X1    g10960(.A1(new_n11216_), .A2(new_n11209_), .ZN(new_n11217_));
  INV_X1     g10961(.I(new_n11215_), .ZN(new_n11218_));
  OAI21_X1   g10962(.A1(new_n10907_), .A2(new_n10619_), .B(new_n11218_), .ZN(new_n11219_));
  NOR2_X1    g10963(.A1(new_n11219_), .A2(new_n11208_), .ZN(new_n11220_));
  NOR2_X1    g10964(.A1(new_n11217_), .A2(new_n11220_), .ZN(new_n11221_));
  XOR2_X1    g10965(.A1(new_n11221_), .A2(new_n11194_), .Z(\f[58] ));
  NAND2_X1   g10966(.A1(new_n11216_), .A2(new_n11209_), .ZN(new_n11223_));
  XNOR2_X1   g10967(.A1(new_n10910_), .A2(new_n11193_), .ZN(new_n11224_));
  OAI21_X1   g10968(.A1(new_n11216_), .A2(new_n11209_), .B(new_n11224_), .ZN(new_n11225_));
  NAND2_X1   g10969(.A1(new_n11225_), .A2(new_n11223_), .ZN(new_n11226_));
  NOR2_X1    g10970(.A1(new_n10862_), .A2(new_n10853_), .ZN(new_n11227_));
  OAI21_X1   g10971(.A1(new_n11227_), .A2(new_n10864_), .B(new_n11168_), .ZN(new_n11228_));
  OAI22_X1   g10972(.A1(new_n713_), .A2(new_n8500_), .B1(new_n8168_), .B2(new_n717_), .ZN(new_n11229_));
  AOI21_X1   g10973(.A1(\b[48] ), .A2(new_n1126_), .B(new_n11229_), .ZN(new_n11230_));
  OAI21_X1   g10974(.A1(new_n8510_), .A2(new_n986_), .B(new_n11230_), .ZN(new_n11231_));
  XOR2_X1    g10975(.A1(new_n11231_), .A2(\a[11] ), .Z(new_n11232_));
  INV_X1     g10976(.I(new_n11232_), .ZN(new_n11233_));
  AOI21_X1   g10977(.A1(new_n11154_), .A2(new_n11153_), .B(new_n10928_), .ZN(new_n11234_));
  INV_X1     g10978(.I(new_n11155_), .ZN(new_n11235_));
  AOI21_X1   g10979(.A1(new_n10923_), .A2(new_n10848_), .B(new_n11235_), .ZN(new_n11236_));
  INV_X1     g10980(.I(new_n7649_), .ZN(new_n11237_));
  OAI22_X1   g10981(.A1(new_n993_), .A2(new_n8126_), .B1(new_n7617_), .B2(new_n997_), .ZN(new_n11238_));
  AOI21_X1   g10982(.A1(\b[45] ), .A2(new_n1486_), .B(new_n11238_), .ZN(new_n11239_));
  OAI21_X1   g10983(.A1(new_n11237_), .A2(new_n1323_), .B(new_n11239_), .ZN(new_n11240_));
  XOR2_X1    g10984(.A1(new_n11240_), .A2(\a[14] ), .Z(new_n11241_));
  OAI21_X1   g10985(.A1(new_n11148_), .A2(new_n11146_), .B(new_n11149_), .ZN(new_n11242_));
  NOR2_X1    g10986(.A1(new_n10937_), .A2(new_n10942_), .ZN(new_n11243_));
  NAND2_X1   g10987(.A1(new_n10934_), .A2(new_n11130_), .ZN(new_n11244_));
  NOR3_X1    g10988(.A1(new_n11128_), .A2(new_n11127_), .A3(new_n11126_), .ZN(new_n11245_));
  AOI21_X1   g10989(.A1(new_n11118_), .A2(new_n11124_), .B(new_n10947_), .ZN(new_n11246_));
  NOR2_X1    g10990(.A1(new_n11245_), .A2(new_n11246_), .ZN(new_n11247_));
  NAND3_X1   g10991(.A1(new_n10933_), .A2(new_n11247_), .A3(new_n10812_), .ZN(new_n11248_));
  AOI22_X1   g10992(.A1(new_n10937_), .A2(new_n10942_), .B1(new_n11244_), .B2(new_n11248_), .ZN(new_n11249_));
  OAI22_X1   g10993(.A1(new_n1751_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n1754_), .ZN(new_n11250_));
  AOI21_X1   g10994(.A1(\b[39] ), .A2(new_n1939_), .B(new_n11250_), .ZN(new_n11251_));
  OAI21_X1   g10995(.A1(new_n6299_), .A2(new_n1757_), .B(new_n11251_), .ZN(new_n11252_));
  XOR2_X1    g10996(.A1(new_n11252_), .A2(\a[20] ), .Z(new_n11253_));
  NOR2_X1    g10997(.A1(new_n10807_), .A2(new_n10800_), .ZN(new_n11254_));
  NOR3_X1    g10998(.A1(new_n11254_), .A2(new_n10809_), .A3(new_n11130_), .ZN(new_n11255_));
  AOI22_X1   g10999(.A1(new_n2202_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n2205_), .ZN(new_n11256_));
  OAI21_X1   g11000(.A1(new_n4886_), .A2(new_n2370_), .B(new_n11256_), .ZN(new_n11257_));
  AOI21_X1   g11001(.A1(new_n5351_), .A2(new_n2208_), .B(new_n11257_), .ZN(new_n11258_));
  XOR2_X1    g11002(.A1(new_n11258_), .A2(new_n2200_), .Z(new_n11259_));
  OAI22_X1   g11003(.A1(new_n2703_), .A2(new_n4666_), .B1(new_n4639_), .B2(new_n2708_), .ZN(new_n11260_));
  AOI21_X1   g11004(.A1(\b[33] ), .A2(new_n2906_), .B(new_n11260_), .ZN(new_n11261_));
  OAI21_X1   g11005(.A1(new_n4676_), .A2(new_n2711_), .B(new_n11261_), .ZN(new_n11262_));
  XOR2_X1    g11006(.A1(new_n11262_), .A2(\a[26] ), .Z(new_n11263_));
  AOI21_X1   g11007(.A1(new_n10955_), .A2(new_n11107_), .B(new_n11099_), .ZN(new_n11264_));
  NOR2_X1    g11008(.A1(new_n11090_), .A2(new_n11077_), .ZN(new_n11265_));
  NAND2_X1   g11009(.A1(new_n11073_), .A2(new_n10745_), .ZN(new_n11266_));
  XOR2_X1    g11010(.A1(new_n11084_), .A2(new_n11266_), .Z(new_n11267_));
  AOI21_X1   g11011(.A1(new_n11090_), .A2(new_n11077_), .B(new_n11267_), .ZN(new_n11268_));
  AOI22_X1   g11012(.A1(new_n4918_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n4921_), .ZN(new_n11269_));
  OAI21_X1   g11013(.A1(new_n2495_), .A2(new_n6099_), .B(new_n11269_), .ZN(new_n11270_));
  AOI21_X1   g11014(.A1(new_n3407_), .A2(new_n4699_), .B(new_n11270_), .ZN(new_n11271_));
  XOR2_X1    g11015(.A1(new_n11271_), .A2(new_n4446_), .Z(new_n11272_));
  NOR2_X1    g11016(.A1(new_n11054_), .A2(new_n11061_), .ZN(new_n11273_));
  NOR3_X1    g11017(.A1(new_n11273_), .A2(new_n11058_), .A3(new_n11272_), .ZN(new_n11274_));
  INV_X1     g11018(.I(new_n11274_), .ZN(new_n11275_));
  OAI21_X1   g11019(.A1(new_n11273_), .A2(new_n11058_), .B(new_n11272_), .ZN(new_n11276_));
  NAND2_X1   g11020(.A1(new_n11051_), .A2(new_n11041_), .ZN(new_n11277_));
  AOI21_X1   g11021(.A1(new_n10961_), .A2(new_n10713_), .B(new_n11039_), .ZN(new_n11278_));
  NOR2_X1    g11022(.A1(new_n10965_), .A2(new_n11030_), .ZN(new_n11279_));
  NOR2_X1    g11023(.A1(new_n11279_), .A2(new_n11029_), .ZN(new_n11280_));
  NOR3_X1    g11024(.A1(new_n11278_), .A2(new_n11038_), .A3(new_n11280_), .ZN(new_n11281_));
  OAI21_X1   g11025(.A1(new_n11278_), .A2(new_n11038_), .B(new_n11280_), .ZN(new_n11282_));
  INV_X1     g11026(.I(new_n11282_), .ZN(new_n11283_));
  AOI22_X1   g11027(.A1(new_n7403_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n7408_), .ZN(new_n11284_));
  OAI21_X1   g11028(.A1(new_n941_), .A2(new_n9488_), .B(new_n11284_), .ZN(new_n11285_));
  AOI21_X1   g11029(.A1(new_n1449_), .A2(new_n7414_), .B(new_n11285_), .ZN(new_n11286_));
  XOR2_X1    g11030(.A1(new_n11286_), .A2(new_n7410_), .Z(new_n11287_));
  OAI21_X1   g11031(.A1(new_n10966_), .A2(new_n10689_), .B(new_n11012_), .ZN(new_n11288_));
  OAI22_X1   g11032(.A1(new_n9461_), .A2(new_n852_), .B1(new_n776_), .B2(new_n9462_), .ZN(new_n11289_));
  AOI21_X1   g11033(.A1(\b[9] ), .A2(new_n8575_), .B(new_n11289_), .ZN(new_n11290_));
  OAI21_X1   g11034(.A1(new_n859_), .A2(new_n9460_), .B(new_n11290_), .ZN(new_n11291_));
  XOR2_X1    g11035(.A1(new_n11291_), .A2(\a[50] ), .Z(new_n11292_));
  NAND2_X1   g11036(.A1(new_n10969_), .A2(new_n11003_), .ZN(new_n11293_));
  NAND3_X1   g11037(.A1(new_n10992_), .A2(new_n10970_), .A3(new_n10673_), .ZN(new_n11294_));
  NAND2_X1   g11038(.A1(new_n11294_), .A2(new_n10995_), .ZN(new_n11295_));
  INV_X1     g11039(.I(new_n10399_), .ZN(new_n11296_));
  INV_X1     g11040(.I(new_n10062_), .ZN(new_n11297_));
  INV_X1     g11041(.I(new_n10064_), .ZN(new_n11298_));
  OAI22_X1   g11042(.A1(new_n11298_), .A2(new_n377_), .B1(new_n339_), .B2(new_n11297_), .ZN(new_n11299_));
  AOI21_X1   g11043(.A1(\b[3] ), .A2(new_n11296_), .B(new_n11299_), .ZN(new_n11300_));
  OAI21_X1   g11044(.A1(new_n566_), .A2(new_n10069_), .B(new_n11300_), .ZN(new_n11301_));
  XOR2_X1    g11045(.A1(new_n11301_), .A2(\a[56] ), .Z(new_n11302_));
  AOI22_X1   g11046(.A1(new_n10981_), .A2(\b[2] ), .B1(new_n10979_), .B2(\b[1] ), .ZN(new_n11303_));
  NOR3_X1    g11047(.A1(new_n10667_), .A2(new_n10976_), .A3(\a[59] ), .ZN(new_n11304_));
  NOR3_X1    g11048(.A1(new_n10669_), .A2(\a[58] ), .A3(new_n10989_), .ZN(new_n11305_));
  NOR2_X1    g11049(.A1(new_n11305_), .A2(new_n11304_), .ZN(new_n11306_));
  OAI21_X1   g11050(.A1(new_n258_), .A2(new_n11306_), .B(new_n11303_), .ZN(new_n11307_));
  AOI21_X1   g11051(.A1(new_n554_), .A2(new_n10984_), .B(new_n11307_), .ZN(new_n11308_));
  XOR2_X1    g11052(.A1(new_n11308_), .A2(new_n10989_), .Z(new_n11309_));
  INV_X1     g11053(.I(new_n11309_), .ZN(new_n11310_));
  NOR2_X1    g11054(.A1(new_n11310_), .A2(new_n10988_), .ZN(new_n11311_));
  INV_X1     g11055(.I(new_n10988_), .ZN(new_n11312_));
  NOR2_X1    g11056(.A1(new_n11312_), .A2(new_n11309_), .ZN(new_n11313_));
  NOR2_X1    g11057(.A1(new_n11311_), .A2(new_n11313_), .ZN(new_n11314_));
  OR2_X2     g11058(.A1(new_n11314_), .A2(new_n11302_), .Z(new_n11315_));
  NAND2_X1   g11059(.A1(new_n11314_), .A2(new_n11302_), .ZN(new_n11316_));
  NAND2_X1   g11060(.A1(new_n11315_), .A2(new_n11316_), .ZN(new_n11317_));
  XNOR2_X1   g11061(.A1(new_n11317_), .A2(new_n11295_), .ZN(new_n11318_));
  AOI22_X1   g11062(.A1(new_n9125_), .A2(\b[8] ), .B1(\b[7] ), .B2(new_n9123_), .ZN(new_n11319_));
  OAI21_X1   g11063(.A1(new_n438_), .A2(new_n9470_), .B(new_n11319_), .ZN(new_n11320_));
  AOI21_X1   g11064(.A1(new_n799_), .A2(new_n9129_), .B(new_n11320_), .ZN(new_n11321_));
  XOR2_X1    g11065(.A1(new_n11321_), .A2(new_n9133_), .Z(new_n11322_));
  INV_X1     g11066(.I(new_n11322_), .ZN(new_n11323_));
  OR2_X2     g11067(.A1(new_n11318_), .A2(new_n11323_), .Z(new_n11324_));
  NAND2_X1   g11068(.A1(new_n11318_), .A2(new_n11323_), .ZN(new_n11325_));
  NAND4_X1   g11069(.A1(new_n11324_), .A2(new_n11002_), .A3(new_n11293_), .A4(new_n11325_), .ZN(new_n11326_));
  NAND2_X1   g11070(.A1(new_n11293_), .A2(new_n11002_), .ZN(new_n11327_));
  NAND2_X1   g11071(.A1(new_n11324_), .A2(new_n11325_), .ZN(new_n11328_));
  NAND2_X1   g11072(.A1(new_n11328_), .A2(new_n11327_), .ZN(new_n11329_));
  AND3_X2    g11073(.A1(new_n11329_), .A2(new_n11292_), .A3(new_n11326_), .Z(new_n11330_));
  AOI21_X1   g11074(.A1(new_n11329_), .A2(new_n11326_), .B(new_n11292_), .ZN(new_n11331_));
  NOR2_X1    g11075(.A1(new_n11330_), .A2(new_n11331_), .ZN(new_n11332_));
  NAND3_X1   g11076(.A1(new_n11288_), .A2(new_n11332_), .A3(new_n11016_), .ZN(new_n11333_));
  AOI21_X1   g11077(.A1(new_n11288_), .A2(new_n11016_), .B(new_n11332_), .ZN(new_n11334_));
  INV_X1     g11078(.I(new_n11334_), .ZN(new_n11335_));
  AOI21_X1   g11079(.A1(new_n11335_), .A2(new_n11333_), .B(new_n11287_), .ZN(new_n11336_));
  INV_X1     g11080(.I(new_n11287_), .ZN(new_n11337_));
  INV_X1     g11081(.I(new_n11333_), .ZN(new_n11338_));
  NOR3_X1    g11082(.A1(new_n11338_), .A2(new_n11334_), .A3(new_n11337_), .ZN(new_n11339_));
  NOR2_X1    g11083(.A1(new_n11336_), .A2(new_n11339_), .ZN(new_n11340_));
  OAI22_X1   g11084(.A1(new_n7730_), .A2(new_n1432_), .B1(new_n1296_), .B2(new_n7731_), .ZN(new_n11341_));
  AOI21_X1   g11085(.A1(\b[15] ), .A2(new_n6887_), .B(new_n11341_), .ZN(new_n11342_));
  OAI21_X1   g11086(.A1(new_n1444_), .A2(new_n7728_), .B(new_n11342_), .ZN(new_n11343_));
  XOR2_X1    g11087(.A1(new_n11343_), .A2(\a[44] ), .Z(new_n11344_));
  XNOR2_X1   g11088(.A1(new_n11340_), .A2(new_n11344_), .ZN(new_n11345_));
  INV_X1     g11089(.I(new_n11345_), .ZN(new_n11346_));
  OAI21_X1   g11090(.A1(new_n11283_), .A2(new_n11281_), .B(new_n11346_), .ZN(new_n11347_));
  NOR2_X1    g11091(.A1(new_n11278_), .A2(new_n11038_), .ZN(new_n11348_));
  INV_X1     g11092(.I(new_n11280_), .ZN(new_n11349_));
  NAND2_X1   g11093(.A1(new_n11348_), .A2(new_n11349_), .ZN(new_n11350_));
  NAND3_X1   g11094(.A1(new_n11350_), .A2(new_n11282_), .A3(new_n11345_), .ZN(new_n11351_));
  AOI22_X1   g11095(.A1(new_n6108_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n6111_), .ZN(new_n11352_));
  OAI21_X1   g11096(.A1(new_n1553_), .A2(new_n7708_), .B(new_n11352_), .ZN(new_n11353_));
  AOI21_X1   g11097(.A1(new_n2452_), .A2(new_n6105_), .B(new_n11353_), .ZN(new_n11354_));
  XOR2_X1    g11098(.A1(new_n11354_), .A2(new_n5849_), .Z(new_n11355_));
  AOI21_X1   g11099(.A1(new_n11347_), .A2(new_n11351_), .B(new_n11355_), .ZN(new_n11356_));
  AOI21_X1   g11100(.A1(new_n11350_), .A2(new_n11282_), .B(new_n11345_), .ZN(new_n11357_));
  NOR3_X1    g11101(.A1(new_n11283_), .A2(new_n11281_), .A3(new_n11346_), .ZN(new_n11358_));
  INV_X1     g11102(.I(new_n11355_), .ZN(new_n11359_));
  NOR3_X1    g11103(.A1(new_n11358_), .A2(new_n11357_), .A3(new_n11359_), .ZN(new_n11360_));
  NOR2_X1    g11104(.A1(new_n11360_), .A2(new_n11356_), .ZN(new_n11361_));
  NAND3_X1   g11105(.A1(new_n11361_), .A2(new_n11277_), .A3(new_n11052_), .ZN(new_n11362_));
  NAND2_X1   g11106(.A1(new_n11277_), .A2(new_n11052_), .ZN(new_n11363_));
  OAI21_X1   g11107(.A1(new_n11358_), .A2(new_n11357_), .B(new_n11359_), .ZN(new_n11364_));
  NAND3_X1   g11108(.A1(new_n11347_), .A2(new_n11351_), .A3(new_n11355_), .ZN(new_n11365_));
  NAND2_X1   g11109(.A1(new_n11364_), .A2(new_n11365_), .ZN(new_n11366_));
  NAND2_X1   g11110(.A1(new_n11363_), .A2(new_n11366_), .ZN(new_n11367_));
  AOI22_X1   g11111(.A1(new_n5155_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n5160_), .ZN(new_n11368_));
  OAI21_X1   g11112(.A1(new_n2027_), .A2(new_n6877_), .B(new_n11368_), .ZN(new_n11369_));
  AOI21_X1   g11113(.A1(new_n2470_), .A2(new_n5166_), .B(new_n11369_), .ZN(new_n11370_));
  XOR2_X1    g11114(.A1(new_n11370_), .A2(new_n5162_), .Z(new_n11371_));
  AOI21_X1   g11115(.A1(new_n11367_), .A2(new_n11362_), .B(new_n11371_), .ZN(new_n11372_));
  NOR2_X1    g11116(.A1(new_n11363_), .A2(new_n11366_), .ZN(new_n11373_));
  AOI21_X1   g11117(.A1(new_n11052_), .A2(new_n11277_), .B(new_n11361_), .ZN(new_n11374_));
  INV_X1     g11118(.I(new_n11371_), .ZN(new_n11375_));
  NOR3_X1    g11119(.A1(new_n11374_), .A2(new_n11373_), .A3(new_n11375_), .ZN(new_n11376_));
  NOR2_X1    g11120(.A1(new_n11376_), .A2(new_n11372_), .ZN(new_n11377_));
  AOI21_X1   g11121(.A1(new_n11275_), .A2(new_n11276_), .B(new_n11377_), .ZN(new_n11378_));
  INV_X1     g11122(.I(new_n11058_), .ZN(new_n11379_));
  INV_X1     g11123(.I(new_n11272_), .ZN(new_n11380_));
  NAND3_X1   g11124(.A1(new_n11057_), .A2(new_n11056_), .A3(new_n11055_), .ZN(new_n11381_));
  INV_X1     g11125(.I(new_n11061_), .ZN(new_n11382_));
  NAND2_X1   g11126(.A1(new_n11382_), .A2(new_n11381_), .ZN(new_n11383_));
  AOI21_X1   g11127(.A1(new_n11383_), .A2(new_n11379_), .B(new_n11380_), .ZN(new_n11384_));
  OAI21_X1   g11128(.A1(new_n11374_), .A2(new_n11373_), .B(new_n11375_), .ZN(new_n11385_));
  NAND3_X1   g11129(.A1(new_n11367_), .A2(new_n11362_), .A3(new_n11371_), .ZN(new_n11386_));
  NAND2_X1   g11130(.A1(new_n11385_), .A2(new_n11386_), .ZN(new_n11387_));
  NOR3_X1    g11131(.A1(new_n11384_), .A2(new_n11387_), .A3(new_n11274_), .ZN(new_n11388_));
  NOR2_X1    g11132(.A1(new_n11378_), .A2(new_n11388_), .ZN(new_n11389_));
  INV_X1     g11133(.I(new_n11065_), .ZN(new_n11390_));
  NAND2_X1   g11134(.A1(new_n11266_), .A2(new_n11390_), .ZN(new_n11391_));
  XOR2_X1    g11135(.A1(new_n11059_), .A2(new_n11061_), .Z(new_n11392_));
  OAI21_X1   g11136(.A1(new_n11266_), .A2(new_n11390_), .B(new_n11392_), .ZN(new_n11393_));
  NAND3_X1   g11137(.A1(new_n11389_), .A2(new_n11393_), .A3(new_n11391_), .ZN(new_n11394_));
  OAI21_X1   g11138(.A1(new_n11384_), .A2(new_n11274_), .B(new_n11387_), .ZN(new_n11395_));
  NAND3_X1   g11139(.A1(new_n11275_), .A2(new_n11377_), .A3(new_n11276_), .ZN(new_n11396_));
  NAND2_X1   g11140(.A1(new_n11396_), .A2(new_n11395_), .ZN(new_n11397_));
  NOR2_X1    g11141(.A1(new_n11085_), .A2(new_n10749_), .ZN(new_n11398_));
  NOR2_X1    g11142(.A1(new_n11398_), .A2(new_n11065_), .ZN(new_n11399_));
  XOR2_X1    g11143(.A1(new_n11059_), .A2(new_n11382_), .Z(new_n11400_));
  AOI21_X1   g11144(.A1(new_n11398_), .A2(new_n11065_), .B(new_n11400_), .ZN(new_n11401_));
  OAI21_X1   g11145(.A1(new_n11399_), .A2(new_n11401_), .B(new_n11397_), .ZN(new_n11402_));
  NAND2_X1   g11146(.A1(new_n11402_), .A2(new_n11394_), .ZN(new_n11403_));
  NOR3_X1    g11147(.A1(new_n11268_), .A2(new_n11265_), .A3(new_n11403_), .ZN(new_n11404_));
  NAND2_X1   g11148(.A1(new_n10956_), .A2(new_n11078_), .ZN(new_n11405_));
  XOR2_X1    g11149(.A1(new_n11084_), .A2(new_n11398_), .Z(new_n11406_));
  OAI21_X1   g11150(.A1(new_n10956_), .A2(new_n11078_), .B(new_n11406_), .ZN(new_n11407_));
  NOR3_X1    g11151(.A1(new_n11397_), .A2(new_n11401_), .A3(new_n11399_), .ZN(new_n11408_));
  AOI21_X1   g11152(.A1(new_n11393_), .A2(new_n11391_), .B(new_n11389_), .ZN(new_n11409_));
  NOR2_X1    g11153(.A1(new_n11409_), .A2(new_n11408_), .ZN(new_n11410_));
  AOI21_X1   g11154(.A1(new_n11407_), .A2(new_n11405_), .B(new_n11410_), .ZN(new_n11411_));
  AOI22_X1   g11155(.A1(new_n3267_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n3270_), .ZN(new_n11412_));
  OAI21_X1   g11156(.A1(new_n3624_), .A2(new_n3475_), .B(new_n11412_), .ZN(new_n11413_));
  AOI21_X1   g11157(.A1(new_n4030_), .A2(new_n3273_), .B(new_n11413_), .ZN(new_n11414_));
  XOR2_X1    g11158(.A1(new_n11414_), .A2(new_n3264_), .Z(new_n11415_));
  AOI22_X1   g11159(.A1(new_n3864_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n3869_), .ZN(new_n11416_));
  OAI21_X1   g11160(.A1(new_n3158_), .A2(new_n5410_), .B(new_n11416_), .ZN(new_n11417_));
  AOI21_X1   g11161(.A1(new_n4188_), .A2(new_n3872_), .B(new_n11417_), .ZN(new_n11418_));
  XOR2_X1    g11162(.A1(new_n11418_), .A2(new_n3876_), .Z(new_n11419_));
  INV_X1     g11163(.I(new_n11419_), .ZN(new_n11420_));
  XOR2_X1    g11164(.A1(new_n11415_), .A2(new_n11420_), .Z(new_n11421_));
  INV_X1     g11165(.I(new_n11421_), .ZN(new_n11422_));
  OAI21_X1   g11166(.A1(new_n11404_), .A2(new_n11411_), .B(new_n11422_), .ZN(new_n11423_));
  NAND3_X1   g11167(.A1(new_n11407_), .A2(new_n11405_), .A3(new_n11410_), .ZN(new_n11424_));
  OAI21_X1   g11168(.A1(new_n11268_), .A2(new_n11265_), .B(new_n11403_), .ZN(new_n11425_));
  NAND3_X1   g11169(.A1(new_n11425_), .A2(new_n11424_), .A3(new_n11421_), .ZN(new_n11426_));
  NAND2_X1   g11170(.A1(new_n11423_), .A2(new_n11426_), .ZN(new_n11427_));
  NAND2_X1   g11171(.A1(new_n11264_), .A2(new_n11427_), .ZN(new_n11428_));
  OAI21_X1   g11172(.A1(new_n11114_), .A2(new_n11113_), .B(new_n11107_), .ZN(new_n11429_));
  NAND2_X1   g11173(.A1(new_n11429_), .A2(new_n11106_), .ZN(new_n11430_));
  AOI21_X1   g11174(.A1(new_n11425_), .A2(new_n11424_), .B(new_n11421_), .ZN(new_n11431_));
  NOR3_X1    g11175(.A1(new_n11404_), .A2(new_n11411_), .A3(new_n11422_), .ZN(new_n11432_));
  NOR2_X1    g11176(.A1(new_n11432_), .A2(new_n11431_), .ZN(new_n11433_));
  NAND2_X1   g11177(.A1(new_n11430_), .A2(new_n11433_), .ZN(new_n11434_));
  AOI21_X1   g11178(.A1(new_n11434_), .A2(new_n11428_), .B(new_n11263_), .ZN(new_n11435_));
  INV_X1     g11179(.I(new_n11263_), .ZN(new_n11436_));
  NOR2_X1    g11180(.A1(new_n11430_), .A2(new_n11433_), .ZN(new_n11437_));
  NOR2_X1    g11181(.A1(new_n11264_), .A2(new_n11427_), .ZN(new_n11438_));
  NOR3_X1    g11182(.A1(new_n11437_), .A2(new_n11438_), .A3(new_n11436_), .ZN(new_n11439_));
  NOR2_X1    g11183(.A1(new_n11439_), .A2(new_n11435_), .ZN(new_n11440_));
  AOI21_X1   g11184(.A1(new_n11105_), .A2(new_n11109_), .B(new_n11111_), .ZN(new_n11441_));
  OAI21_X1   g11185(.A1(new_n11127_), .A2(new_n11441_), .B(new_n11440_), .ZN(new_n11442_));
  OAI21_X1   g11186(.A1(new_n11437_), .A2(new_n11438_), .B(new_n11436_), .ZN(new_n11443_));
  NAND3_X1   g11187(.A1(new_n11434_), .A2(new_n11428_), .A3(new_n11263_), .ZN(new_n11444_));
  NAND2_X1   g11188(.A1(new_n11443_), .A2(new_n11444_), .ZN(new_n11445_));
  INV_X1     g11189(.I(new_n11441_), .ZN(new_n11446_));
  NAND3_X1   g11190(.A1(new_n11118_), .A2(new_n11445_), .A3(new_n11446_), .ZN(new_n11447_));
  AOI21_X1   g11191(.A1(new_n11442_), .A2(new_n11447_), .B(new_n11259_), .ZN(new_n11448_));
  INV_X1     g11192(.I(new_n11259_), .ZN(new_n11449_));
  AOI21_X1   g11193(.A1(new_n11118_), .A2(new_n11446_), .B(new_n11445_), .ZN(new_n11450_));
  NOR3_X1    g11194(.A1(new_n11440_), .A2(new_n11127_), .A3(new_n11441_), .ZN(new_n11451_));
  NOR3_X1    g11195(.A1(new_n11450_), .A2(new_n11451_), .A3(new_n11449_), .ZN(new_n11452_));
  NOR2_X1    g11196(.A1(new_n11448_), .A2(new_n11452_), .ZN(new_n11453_));
  OAI21_X1   g11197(.A1(new_n11255_), .A2(new_n11245_), .B(new_n11453_), .ZN(new_n11454_));
  OAI21_X1   g11198(.A1(new_n11450_), .A2(new_n11451_), .B(new_n11449_), .ZN(new_n11455_));
  NAND3_X1   g11199(.A1(new_n11442_), .A2(new_n11447_), .A3(new_n11259_), .ZN(new_n11456_));
  NAND2_X1   g11200(.A1(new_n11455_), .A2(new_n11456_), .ZN(new_n11457_));
  NAND3_X1   g11201(.A1(new_n11248_), .A2(new_n11457_), .A3(new_n11125_), .ZN(new_n11458_));
  NAND3_X1   g11202(.A1(new_n11454_), .A2(new_n11458_), .A3(new_n11253_), .ZN(new_n11459_));
  INV_X1     g11203(.I(new_n11253_), .ZN(new_n11460_));
  AOI21_X1   g11204(.A1(new_n11248_), .A2(new_n11125_), .B(new_n11457_), .ZN(new_n11461_));
  NOR3_X1    g11205(.A1(new_n11255_), .A2(new_n11453_), .A3(new_n11245_), .ZN(new_n11462_));
  OAI21_X1   g11206(.A1(new_n11462_), .A2(new_n11461_), .B(new_n11460_), .ZN(new_n11463_));
  NAND2_X1   g11207(.A1(new_n11463_), .A2(new_n11459_), .ZN(new_n11464_));
  OAI21_X1   g11208(.A1(new_n11249_), .A2(new_n11243_), .B(new_n11464_), .ZN(new_n11465_));
  NAND2_X1   g11209(.A1(new_n10932_), .A2(new_n10943_), .ZN(new_n11466_));
  NAND2_X1   g11210(.A1(new_n11244_), .A2(new_n11248_), .ZN(new_n11467_));
  OAI21_X1   g11211(.A1(new_n10932_), .A2(new_n10943_), .B(new_n11467_), .ZN(new_n11468_));
  NOR3_X1    g11212(.A1(new_n11462_), .A2(new_n11461_), .A3(new_n11460_), .ZN(new_n11469_));
  AOI21_X1   g11213(.A1(new_n11454_), .A2(new_n11458_), .B(new_n11253_), .ZN(new_n11470_));
  NOR2_X1    g11214(.A1(new_n11469_), .A2(new_n11470_), .ZN(new_n11471_));
  NAND3_X1   g11215(.A1(new_n11471_), .A2(new_n11468_), .A3(new_n11466_), .ZN(new_n11472_));
  OAI22_X1   g11216(.A1(new_n1592_), .A2(new_n7074_), .B1(new_n6775_), .B2(new_n1505_), .ZN(new_n11473_));
  AOI21_X1   g11217(.A1(\b[42] ), .A2(new_n1584_), .B(new_n11473_), .ZN(new_n11474_));
  OAI21_X1   g11218(.A1(new_n7081_), .A2(new_n1732_), .B(new_n11474_), .ZN(new_n11475_));
  XOR2_X1    g11219(.A1(new_n11475_), .A2(\a[17] ), .Z(new_n11476_));
  AOI21_X1   g11220(.A1(new_n11465_), .A2(new_n11472_), .B(new_n11476_), .ZN(new_n11477_));
  AOI21_X1   g11221(.A1(new_n11466_), .A2(new_n11468_), .B(new_n11471_), .ZN(new_n11478_));
  NOR3_X1    g11222(.A1(new_n11249_), .A2(new_n11464_), .A3(new_n11243_), .ZN(new_n11479_));
  INV_X1     g11223(.I(new_n11476_), .ZN(new_n11480_));
  NOR3_X1    g11224(.A1(new_n11478_), .A2(new_n11479_), .A3(new_n11480_), .ZN(new_n11481_));
  NOR2_X1    g11225(.A1(new_n11481_), .A2(new_n11477_), .ZN(new_n11482_));
  NOR2_X1    g11226(.A1(new_n11242_), .A2(new_n11482_), .ZN(new_n11483_));
  OAI21_X1   g11227(.A1(new_n10931_), .A2(new_n10835_), .B(new_n11150_), .ZN(new_n11484_));
  OAI21_X1   g11228(.A1(new_n11478_), .A2(new_n11479_), .B(new_n11480_), .ZN(new_n11485_));
  NAND3_X1   g11229(.A1(new_n11465_), .A2(new_n11472_), .A3(new_n11476_), .ZN(new_n11486_));
  NAND2_X1   g11230(.A1(new_n11485_), .A2(new_n11486_), .ZN(new_n11487_));
  AOI21_X1   g11231(.A1(new_n11149_), .A2(new_n11484_), .B(new_n11487_), .ZN(new_n11488_));
  OAI21_X1   g11232(.A1(new_n11483_), .A2(new_n11488_), .B(new_n11241_), .ZN(new_n11489_));
  INV_X1     g11233(.I(new_n11241_), .ZN(new_n11490_));
  NAND3_X1   g11234(.A1(new_n11487_), .A2(new_n11484_), .A3(new_n11149_), .ZN(new_n11491_));
  NAND2_X1   g11235(.A1(new_n11242_), .A2(new_n11482_), .ZN(new_n11492_));
  NAND3_X1   g11236(.A1(new_n11492_), .A2(new_n11491_), .A3(new_n11490_), .ZN(new_n11493_));
  NAND2_X1   g11237(.A1(new_n11489_), .A2(new_n11493_), .ZN(new_n11494_));
  NOR3_X1    g11238(.A1(new_n11236_), .A2(new_n11494_), .A3(new_n11234_), .ZN(new_n11495_));
  AOI21_X1   g11239(.A1(new_n10843_), .A2(new_n10845_), .B(new_n10850_), .ZN(new_n11496_));
  OAI21_X1   g11240(.A1(new_n11496_), .A2(new_n10847_), .B(new_n11155_), .ZN(new_n11497_));
  AOI21_X1   g11241(.A1(new_n11492_), .A2(new_n11491_), .B(new_n11490_), .ZN(new_n11498_));
  NOR3_X1    g11242(.A1(new_n11483_), .A2(new_n11488_), .A3(new_n11241_), .ZN(new_n11499_));
  NOR2_X1    g11243(.A1(new_n11499_), .A2(new_n11498_), .ZN(new_n11500_));
  AOI21_X1   g11244(.A1(new_n11152_), .A2(new_n11497_), .B(new_n11500_), .ZN(new_n11501_));
  OAI21_X1   g11245(.A1(new_n11501_), .A2(new_n11495_), .B(new_n11233_), .ZN(new_n11502_));
  NAND3_X1   g11246(.A1(new_n11497_), .A2(new_n11500_), .A3(new_n11152_), .ZN(new_n11503_));
  OAI21_X1   g11247(.A1(new_n11236_), .A2(new_n11234_), .B(new_n11494_), .ZN(new_n11504_));
  NAND3_X1   g11248(.A1(new_n11504_), .A2(new_n11503_), .A3(new_n11232_), .ZN(new_n11505_));
  NAND2_X1   g11249(.A1(new_n11502_), .A2(new_n11505_), .ZN(new_n11506_));
  AOI21_X1   g11250(.A1(new_n11228_), .A2(new_n11165_), .B(new_n11506_), .ZN(new_n11507_));
  AOI21_X1   g11251(.A1(new_n10922_), .A2(new_n10870_), .B(new_n11173_), .ZN(new_n11508_));
  AOI21_X1   g11252(.A1(new_n11504_), .A2(new_n11503_), .B(new_n11232_), .ZN(new_n11509_));
  NOR3_X1    g11253(.A1(new_n11501_), .A2(new_n11495_), .A3(new_n11233_), .ZN(new_n11510_));
  NOR2_X1    g11254(.A1(new_n11510_), .A2(new_n11509_), .ZN(new_n11511_));
  NOR3_X1    g11255(.A1(new_n11511_), .A2(new_n11508_), .A3(new_n11172_), .ZN(new_n11512_));
  OAI22_X1   g11256(.A1(new_n610_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n612_), .ZN(new_n11513_));
  AOI21_X1   g11257(.A1(\b[51] ), .A2(new_n826_), .B(new_n11513_), .ZN(new_n11514_));
  OAI21_X1   g11258(.A1(new_n9385_), .A2(new_n624_), .B(new_n11514_), .ZN(new_n11515_));
  XOR2_X1    g11259(.A1(new_n11515_), .A2(\a[8] ), .Z(new_n11516_));
  NOR3_X1    g11260(.A1(new_n11507_), .A2(new_n11512_), .A3(new_n11516_), .ZN(new_n11517_));
  OAI21_X1   g11261(.A1(new_n11508_), .A2(new_n11172_), .B(new_n11511_), .ZN(new_n11518_));
  NAND3_X1   g11262(.A1(new_n11506_), .A2(new_n11228_), .A3(new_n11165_), .ZN(new_n11519_));
  INV_X1     g11263(.I(new_n11516_), .ZN(new_n11520_));
  AOI21_X1   g11264(.A1(new_n11518_), .A2(new_n11519_), .B(new_n11520_), .ZN(new_n11521_));
  NOR2_X1    g11265(.A1(new_n11521_), .A2(new_n11517_), .ZN(new_n11522_));
  AOI21_X1   g11266(.A1(new_n10916_), .A2(new_n10917_), .B(new_n11184_), .ZN(new_n11523_));
  INV_X1     g11267(.I(new_n11523_), .ZN(new_n11524_));
  NAND3_X1   g11268(.A1(new_n11524_), .A2(new_n11180_), .A3(new_n11522_), .ZN(new_n11525_));
  NAND3_X1   g11269(.A1(new_n11518_), .A2(new_n11519_), .A3(new_n11520_), .ZN(new_n11526_));
  OAI21_X1   g11270(.A1(new_n11507_), .A2(new_n11512_), .B(new_n11516_), .ZN(new_n11527_));
  NAND2_X1   g11271(.A1(new_n11526_), .A2(new_n11527_), .ZN(new_n11528_));
  OAI21_X1   g11272(.A1(new_n11185_), .A2(new_n11523_), .B(new_n11528_), .ZN(new_n11529_));
  AOI22_X1   g11273(.A1(new_n267_), .A2(\b[59] ), .B1(\b[58] ), .B2(new_n261_), .ZN(new_n11530_));
  OAI21_X1   g11274(.A1(new_n10625_), .A2(new_n284_), .B(new_n11530_), .ZN(new_n11531_));
  NOR3_X1    g11275(.A1(new_n11200_), .A2(\b[57] ), .A3(new_n11195_), .ZN(new_n11532_));
  NOR4_X1    g11276(.A1(new_n11198_), .A2(new_n11199_), .A3(new_n10625_), .A4(\b[58] ), .ZN(new_n11533_));
  OAI21_X1   g11277(.A1(new_n11532_), .A2(new_n11533_), .B(\b[59] ), .ZN(new_n11534_));
  INV_X1     g11278(.I(new_n11534_), .ZN(new_n11535_));
  NOR3_X1    g11279(.A1(new_n11532_), .A2(\b[59] ), .A3(new_n11533_), .ZN(new_n11536_));
  NOR3_X1    g11280(.A1(new_n11535_), .A2(new_n279_), .A3(new_n11536_), .ZN(new_n11537_));
  OAI21_X1   g11281(.A1(new_n11537_), .A2(new_n11531_), .B(\a[2] ), .ZN(new_n11538_));
  INV_X1     g11282(.I(new_n11531_), .ZN(new_n11539_));
  INV_X1     g11283(.I(new_n11536_), .ZN(new_n11540_));
  NAND3_X1   g11284(.A1(new_n11540_), .A2(new_n265_), .A3(new_n11534_), .ZN(new_n11541_));
  NAND3_X1   g11285(.A1(new_n11541_), .A2(new_n270_), .A3(new_n11539_), .ZN(new_n11542_));
  AOI22_X1   g11286(.A1(new_n800_), .A2(\b[55] ), .B1(\b[56] ), .B2(new_n333_), .ZN(new_n11543_));
  OAI21_X1   g11287(.A1(new_n9942_), .A2(new_n392_), .B(new_n11543_), .ZN(new_n11544_));
  AOI21_X1   g11288(.A1(new_n10318_), .A2(new_n330_), .B(new_n11544_), .ZN(new_n11545_));
  XOR2_X1    g11289(.A1(new_n11545_), .A2(new_n312_), .Z(new_n11546_));
  AOI21_X1   g11290(.A1(new_n11538_), .A2(new_n11542_), .B(new_n11546_), .ZN(new_n11547_));
  AOI21_X1   g11291(.A1(new_n11541_), .A2(new_n11539_), .B(new_n270_), .ZN(new_n11548_));
  NOR3_X1    g11292(.A1(new_n11537_), .A2(\a[2] ), .A3(new_n11531_), .ZN(new_n11549_));
  INV_X1     g11293(.I(new_n11546_), .ZN(new_n11550_));
  NOR3_X1    g11294(.A1(new_n11549_), .A2(new_n11548_), .A3(new_n11550_), .ZN(new_n11551_));
  NOR2_X1    g11295(.A1(new_n11551_), .A2(new_n11547_), .ZN(new_n11552_));
  AOI21_X1   g11296(.A1(new_n11525_), .A2(new_n11529_), .B(new_n11552_), .ZN(new_n11553_));
  NOR3_X1    g11297(.A1(new_n11528_), .A2(new_n11523_), .A3(new_n11185_), .ZN(new_n11554_));
  AOI21_X1   g11298(.A1(new_n11524_), .A2(new_n11180_), .B(new_n11522_), .ZN(new_n11555_));
  OAI21_X1   g11299(.A1(new_n11549_), .A2(new_n11548_), .B(new_n11550_), .ZN(new_n11556_));
  NAND3_X1   g11300(.A1(new_n11538_), .A2(new_n11542_), .A3(new_n11546_), .ZN(new_n11557_));
  NAND2_X1   g11301(.A1(new_n11556_), .A2(new_n11557_), .ZN(new_n11558_));
  NOR3_X1    g11302(.A1(new_n11558_), .A2(new_n11555_), .A3(new_n11554_), .ZN(new_n11559_));
  NOR2_X1    g11303(.A1(new_n11553_), .A2(new_n11559_), .ZN(new_n11560_));
  NAND2_X1   g11304(.A1(new_n11190_), .A2(new_n11191_), .ZN(new_n11561_));
  AOI22_X1   g11305(.A1(new_n10909_), .A2(new_n10898_), .B1(new_n10914_), .B2(new_n11561_), .ZN(new_n11562_));
  INV_X1     g11306(.I(new_n11562_), .ZN(new_n11563_));
  NAND3_X1   g11307(.A1(new_n11560_), .A2(new_n11563_), .A3(new_n11192_), .ZN(new_n11564_));
  INV_X1     g11308(.I(new_n11192_), .ZN(new_n11565_));
  OAI21_X1   g11309(.A1(new_n11555_), .A2(new_n11554_), .B(new_n11558_), .ZN(new_n11566_));
  NAND3_X1   g11310(.A1(new_n11552_), .A2(new_n11525_), .A3(new_n11529_), .ZN(new_n11567_));
  NAND2_X1   g11311(.A1(new_n11566_), .A2(new_n11567_), .ZN(new_n11568_));
  OAI21_X1   g11312(.A1(new_n11562_), .A2(new_n11565_), .B(new_n11568_), .ZN(new_n11569_));
  NAND2_X1   g11313(.A1(new_n11569_), .A2(new_n11564_), .ZN(new_n11570_));
  XOR2_X1    g11314(.A1(new_n11226_), .A2(new_n11570_), .Z(\f[59] ));
  NAND2_X1   g11315(.A1(new_n11525_), .A2(new_n11529_), .ZN(new_n11572_));
  AOI21_X1   g11316(.A1(new_n11572_), .A2(new_n11557_), .B(new_n11547_), .ZN(new_n11573_));
  AOI21_X1   g11317(.A1(new_n11228_), .A2(new_n11165_), .B(new_n11510_), .ZN(new_n11574_));
  NOR2_X1    g11318(.A1(new_n11574_), .A2(new_n11509_), .ZN(new_n11575_));
  INV_X1     g11319(.I(new_n11575_), .ZN(new_n11576_));
  INV_X1     g11320(.I(new_n8783_), .ZN(new_n11577_));
  OAI22_X1   g11321(.A1(new_n713_), .A2(new_n8776_), .B1(new_n8500_), .B2(new_n717_), .ZN(new_n11578_));
  AOI21_X1   g11322(.A1(\b[49] ), .A2(new_n1126_), .B(new_n11578_), .ZN(new_n11579_));
  OAI21_X1   g11323(.A1(new_n11577_), .A2(new_n986_), .B(new_n11579_), .ZN(new_n11580_));
  XOR2_X1    g11324(.A1(new_n11580_), .A2(\a[11] ), .Z(new_n11581_));
  INV_X1     g11325(.I(new_n11581_), .ZN(new_n11582_));
  AOI21_X1   g11326(.A1(new_n11242_), .A2(new_n11486_), .B(new_n11477_), .ZN(new_n11583_));
  INV_X1     g11327(.I(new_n11583_), .ZN(new_n11584_));
  OAI22_X1   g11328(.A1(new_n1592_), .A2(new_n7096_), .B1(new_n7074_), .B2(new_n1505_), .ZN(new_n11585_));
  AOI21_X1   g11329(.A1(\b[43] ), .A2(new_n1584_), .B(new_n11585_), .ZN(new_n11586_));
  OAI21_X1   g11330(.A1(new_n7925_), .A2(new_n1732_), .B(new_n11586_), .ZN(new_n11587_));
  XOR2_X1    g11331(.A1(new_n11587_), .A2(\a[17] ), .Z(new_n11588_));
  INV_X1     g11332(.I(new_n11588_), .ZN(new_n11589_));
  AOI21_X1   g11333(.A1(new_n11363_), .A2(new_n11365_), .B(new_n11356_), .ZN(new_n11590_));
  AOI22_X1   g11334(.A1(new_n6108_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n6111_), .ZN(new_n11591_));
  OAI21_X1   g11335(.A1(new_n1859_), .A2(new_n7708_), .B(new_n11591_), .ZN(new_n11592_));
  AOI21_X1   g11336(.A1(new_n2032_), .A2(new_n6105_), .B(new_n11592_), .ZN(new_n11593_));
  XOR2_X1    g11337(.A1(new_n11593_), .A2(new_n5849_), .Z(new_n11594_));
  INV_X1     g11338(.I(new_n11594_), .ZN(new_n11595_));
  NOR2_X1    g11339(.A1(new_n11348_), .A2(new_n11344_), .ZN(new_n11596_));
  OAI21_X1   g11340(.A1(new_n11336_), .A2(new_n11339_), .B(new_n11349_), .ZN(new_n11597_));
  OAI21_X1   g11341(.A1(new_n10964_), .A2(new_n10963_), .B(new_n11027_), .ZN(new_n11598_));
  NAND3_X1   g11342(.A1(new_n11598_), .A2(new_n11024_), .A3(new_n11340_), .ZN(new_n11599_));
  AOI22_X1   g11343(.A1(new_n11348_), .A2(new_n11344_), .B1(new_n11597_), .B2(new_n11599_), .ZN(new_n11600_));
  AOI22_X1   g11344(.A1(new_n6569_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n6574_), .ZN(new_n11601_));
  OAI21_X1   g11345(.A1(new_n1296_), .A2(new_n8565_), .B(new_n11601_), .ZN(new_n11602_));
  AOI21_X1   g11346(.A1(new_n2038_), .A2(new_n6579_), .B(new_n11602_), .ZN(new_n11603_));
  XOR2_X1    g11347(.A1(new_n11603_), .A2(new_n6567_), .Z(new_n11604_));
  NAND2_X1   g11348(.A1(new_n11295_), .A2(new_n11316_), .ZN(new_n11605_));
  NAND2_X1   g11349(.A1(new_n11605_), .A2(new_n11315_), .ZN(new_n11606_));
  INV_X1     g11350(.I(new_n11606_), .ZN(new_n11607_));
  AOI22_X1   g11351(.A1(new_n10064_), .A2(\b[6] ), .B1(\b[5] ), .B2(new_n10062_), .ZN(new_n11608_));
  OAI21_X1   g11352(.A1(new_n339_), .A2(new_n10399_), .B(new_n11608_), .ZN(new_n11609_));
  AOI21_X1   g11353(.A1(new_n916_), .A2(new_n10068_), .B(new_n11609_), .ZN(new_n11610_));
  XOR2_X1    g11354(.A1(new_n11610_), .A2(new_n10057_), .Z(new_n11611_));
  INV_X1     g11355(.I(new_n11611_), .ZN(new_n11612_));
  AOI22_X1   g11356(.A1(new_n10981_), .A2(\b[3] ), .B1(new_n10979_), .B2(\b[2] ), .ZN(new_n11613_));
  OAI21_X1   g11357(.A1(new_n275_), .A2(new_n11306_), .B(new_n11613_), .ZN(new_n11614_));
  AOI21_X1   g11358(.A1(new_n299_), .A2(new_n10984_), .B(new_n11614_), .ZN(new_n11615_));
  XOR2_X1    g11359(.A1(new_n11615_), .A2(\a[59] ), .Z(new_n11616_));
  NAND2_X1   g11360(.A1(\a[59] ), .A2(\a[60] ), .ZN(new_n11617_));
  INV_X1     g11361(.I(new_n11617_), .ZN(new_n11618_));
  NOR2_X1    g11362(.A1(\a[59] ), .A2(\a[60] ), .ZN(new_n11619_));
  NOR2_X1    g11363(.A1(new_n11618_), .A2(new_n11619_), .ZN(new_n11620_));
  INV_X1     g11364(.I(new_n11620_), .ZN(new_n11621_));
  NOR2_X1    g11365(.A1(new_n11621_), .A2(new_n258_), .ZN(new_n11622_));
  INV_X1     g11366(.I(new_n11622_), .ZN(new_n11623_));
  NOR2_X1    g11367(.A1(new_n11616_), .A2(new_n11623_), .ZN(new_n11624_));
  INV_X1     g11368(.I(new_n11624_), .ZN(new_n11625_));
  NAND2_X1   g11369(.A1(new_n11616_), .A2(new_n11623_), .ZN(new_n11626_));
  NAND2_X1   g11370(.A1(new_n11625_), .A2(new_n11626_), .ZN(new_n11627_));
  XOR2_X1    g11371(.A1(new_n11627_), .A2(new_n11311_), .Z(new_n11628_));
  NAND2_X1   g11372(.A1(new_n11628_), .A2(new_n11612_), .ZN(new_n11629_));
  INV_X1     g11373(.I(new_n11629_), .ZN(new_n11630_));
  NOR2_X1    g11374(.A1(new_n11628_), .A2(new_n11612_), .ZN(new_n11631_));
  NOR2_X1    g11375(.A1(new_n11630_), .A2(new_n11631_), .ZN(new_n11632_));
  XOR2_X1    g11376(.A1(new_n11632_), .A2(new_n11607_), .Z(new_n11633_));
  INV_X1     g11377(.I(new_n11633_), .ZN(new_n11634_));
  AOI22_X1   g11378(.A1(new_n9125_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n9123_), .ZN(new_n11635_));
  OAI21_X1   g11379(.A1(new_n471_), .A2(new_n9470_), .B(new_n11635_), .ZN(new_n11636_));
  AOI21_X1   g11380(.A1(new_n676_), .A2(new_n9129_), .B(new_n11636_), .ZN(new_n11637_));
  XOR2_X1    g11381(.A1(new_n11637_), .A2(new_n9133_), .Z(new_n11638_));
  NAND2_X1   g11382(.A1(new_n11326_), .A2(new_n11324_), .ZN(new_n11639_));
  NAND2_X1   g11383(.A1(new_n11639_), .A2(new_n11638_), .ZN(new_n11640_));
  NOR2_X1    g11384(.A1(new_n11639_), .A2(new_n11638_), .ZN(new_n11641_));
  INV_X1     g11385(.I(new_n11641_), .ZN(new_n11642_));
  NAND2_X1   g11386(.A1(new_n11642_), .A2(new_n11640_), .ZN(new_n11643_));
  XOR2_X1    g11387(.A1(new_n11643_), .A2(new_n11634_), .Z(new_n11644_));
  INV_X1     g11388(.I(new_n11644_), .ZN(new_n11645_));
  AOI22_X1   g11389(.A1(new_n8241_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n8246_), .ZN(new_n11646_));
  OAI21_X1   g11390(.A1(new_n776_), .A2(new_n9114_), .B(new_n11646_), .ZN(new_n11647_));
  AOI21_X1   g11391(.A1(new_n1194_), .A2(new_n8252_), .B(new_n11647_), .ZN(new_n11648_));
  XOR2_X1    g11392(.A1(new_n11648_), .A2(new_n8248_), .Z(new_n11649_));
  OAI21_X1   g11393(.A1(new_n11338_), .A2(new_n11330_), .B(new_n11649_), .ZN(new_n11650_));
  INV_X1     g11394(.I(new_n11650_), .ZN(new_n11651_));
  NOR3_X1    g11395(.A1(new_n11338_), .A2(new_n11330_), .A3(new_n11649_), .ZN(new_n11652_));
  NOR3_X1    g11396(.A1(new_n11651_), .A2(new_n11645_), .A3(new_n11652_), .ZN(new_n11653_));
  INV_X1     g11397(.I(new_n11652_), .ZN(new_n11654_));
  AOI21_X1   g11398(.A1(new_n11654_), .A2(new_n11650_), .B(new_n11644_), .ZN(new_n11655_));
  NOR2_X1    g11399(.A1(new_n11655_), .A2(new_n11653_), .ZN(new_n11656_));
  NOR4_X1    g11400(.A1(new_n11279_), .A2(new_n11029_), .A3(new_n11336_), .A4(new_n11339_), .ZN(new_n11657_));
  OAI22_X1   g11401(.A1(new_n1093_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n1268_), .ZN(new_n11658_));
  AOI21_X1   g11402(.A1(\b[13] ), .A2(new_n7719_), .B(new_n11658_), .ZN(new_n11659_));
  OAI21_X1   g11403(.A1(new_n1275_), .A2(new_n8585_), .B(new_n11659_), .ZN(new_n11660_));
  XOR2_X1    g11404(.A1(new_n11660_), .A2(\a[47] ), .Z(new_n11661_));
  OAI21_X1   g11405(.A1(new_n11657_), .A2(new_n11339_), .B(new_n11661_), .ZN(new_n11662_));
  INV_X1     g11406(.I(new_n11339_), .ZN(new_n11663_));
  INV_X1     g11407(.I(new_n11661_), .ZN(new_n11664_));
  NAND3_X1   g11408(.A1(new_n11599_), .A2(new_n11663_), .A3(new_n11664_), .ZN(new_n11665_));
  NAND3_X1   g11409(.A1(new_n11662_), .A2(new_n11665_), .A3(new_n11656_), .ZN(new_n11666_));
  INV_X1     g11410(.I(new_n11656_), .ZN(new_n11667_));
  AOI21_X1   g11411(.A1(new_n11599_), .A2(new_n11663_), .B(new_n11664_), .ZN(new_n11668_));
  NOR3_X1    g11412(.A1(new_n11657_), .A2(new_n11339_), .A3(new_n11661_), .ZN(new_n11669_));
  OAI21_X1   g11413(.A1(new_n11669_), .A2(new_n11668_), .B(new_n11667_), .ZN(new_n11670_));
  AOI21_X1   g11414(.A1(new_n11670_), .A2(new_n11666_), .B(new_n11604_), .ZN(new_n11671_));
  INV_X1     g11415(.I(new_n11604_), .ZN(new_n11672_));
  NOR3_X1    g11416(.A1(new_n11669_), .A2(new_n11667_), .A3(new_n11668_), .ZN(new_n11673_));
  AOI21_X1   g11417(.A1(new_n11662_), .A2(new_n11665_), .B(new_n11656_), .ZN(new_n11674_));
  NOR3_X1    g11418(.A1(new_n11673_), .A2(new_n11674_), .A3(new_n11672_), .ZN(new_n11675_));
  OR4_X2     g11419(.A1(new_n11596_), .A2(new_n11600_), .A3(new_n11671_), .A4(new_n11675_), .Z(new_n11676_));
  OR2_X2     g11420(.A1(new_n11675_), .A2(new_n11671_), .Z(new_n11677_));
  OAI21_X1   g11421(.A1(new_n11596_), .A2(new_n11600_), .B(new_n11677_), .ZN(new_n11678_));
  NAND2_X1   g11422(.A1(new_n11678_), .A2(new_n11676_), .ZN(new_n11679_));
  NAND2_X1   g11423(.A1(new_n11679_), .A2(new_n11595_), .ZN(new_n11680_));
  INV_X1     g11424(.I(new_n11680_), .ZN(new_n11681_));
  NOR2_X1    g11425(.A1(new_n11679_), .A2(new_n11595_), .ZN(new_n11682_));
  NOR2_X1    g11426(.A1(new_n11681_), .A2(new_n11682_), .ZN(new_n11683_));
  XOR2_X1    g11427(.A1(new_n11683_), .A2(new_n11590_), .Z(new_n11684_));
  NOR2_X1    g11428(.A1(new_n11273_), .A2(new_n11058_), .ZN(new_n11685_));
  NAND2_X1   g11429(.A1(new_n11685_), .A2(new_n11386_), .ZN(new_n11686_));
  AOI22_X1   g11430(.A1(new_n5155_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n5160_), .ZN(new_n11687_));
  OAI21_X1   g11431(.A1(new_n2142_), .A2(new_n6877_), .B(new_n11687_), .ZN(new_n11688_));
  AOI21_X1   g11432(.A1(new_n3033_), .A2(new_n5166_), .B(new_n11688_), .ZN(new_n11689_));
  XOR2_X1    g11433(.A1(new_n11689_), .A2(new_n5162_), .Z(new_n11690_));
  AOI21_X1   g11434(.A1(new_n11686_), .A2(new_n11385_), .B(new_n11690_), .ZN(new_n11691_));
  NAND3_X1   g11435(.A1(new_n11686_), .A2(new_n11385_), .A3(new_n11690_), .ZN(new_n11692_));
  INV_X1     g11436(.I(new_n11692_), .ZN(new_n11693_));
  NOR3_X1    g11437(.A1(new_n11693_), .A2(new_n11684_), .A3(new_n11691_), .ZN(new_n11694_));
  INV_X1     g11438(.I(new_n11684_), .ZN(new_n11695_));
  INV_X1     g11439(.I(new_n11691_), .ZN(new_n11696_));
  AOI21_X1   g11440(.A1(new_n11696_), .A2(new_n11692_), .B(new_n11695_), .ZN(new_n11697_));
  NOR2_X1    g11441(.A1(new_n11697_), .A2(new_n11694_), .ZN(new_n11698_));
  INV_X1     g11442(.I(new_n11698_), .ZN(new_n11699_));
  OAI22_X1   g11443(.A1(new_n3158_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n3006_), .ZN(new_n11700_));
  AOI21_X1   g11444(.A1(\b[25] ), .A2(new_n4706_), .B(new_n11700_), .ZN(new_n11701_));
  OAI21_X1   g11445(.A1(new_n3165_), .A2(new_n4458_), .B(new_n11701_), .ZN(new_n11702_));
  XOR2_X1    g11446(.A1(new_n11702_), .A2(\a[35] ), .Z(new_n11703_));
  INV_X1     g11447(.I(new_n11703_), .ZN(new_n11704_));
  XOR2_X1    g11448(.A1(new_n11387_), .A2(new_n11685_), .Z(new_n11705_));
  NAND2_X1   g11449(.A1(new_n11705_), .A2(new_n11272_), .ZN(new_n11706_));
  AOI21_X1   g11450(.A1(new_n11394_), .A2(new_n11706_), .B(new_n11704_), .ZN(new_n11707_));
  NAND3_X1   g11451(.A1(new_n11394_), .A2(new_n11706_), .A3(new_n11704_), .ZN(new_n11708_));
  INV_X1     g11452(.I(new_n11708_), .ZN(new_n11709_));
  NOR3_X1    g11453(.A1(new_n11699_), .A2(new_n11707_), .A3(new_n11709_), .ZN(new_n11710_));
  NOR2_X1    g11454(.A1(new_n11709_), .A2(new_n11707_), .ZN(new_n11711_));
  NOR2_X1    g11455(.A1(new_n11711_), .A2(new_n11698_), .ZN(new_n11712_));
  NOR2_X1    g11456(.A1(new_n11712_), .A2(new_n11710_), .ZN(new_n11713_));
  INV_X1     g11457(.I(new_n11713_), .ZN(new_n11714_));
  AOI22_X1   g11458(.A1(new_n3864_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n3869_), .ZN(new_n11715_));
  OAI21_X1   g11459(.A1(new_n3185_), .A2(new_n5410_), .B(new_n11715_), .ZN(new_n11716_));
  AOI21_X1   g11460(.A1(new_n4230_), .A2(new_n3872_), .B(new_n11716_), .ZN(new_n11717_));
  XOR2_X1    g11461(.A1(new_n11717_), .A2(new_n3876_), .Z(new_n11718_));
  INV_X1     g11462(.I(new_n11718_), .ZN(new_n11719_));
  NOR2_X1    g11463(.A1(new_n11403_), .A2(new_n11420_), .ZN(new_n11720_));
  INV_X1     g11464(.I(new_n11720_), .ZN(new_n11721_));
  NOR2_X1    g11465(.A1(new_n11268_), .A2(new_n11265_), .ZN(new_n11722_));
  NOR2_X1    g11466(.A1(new_n11410_), .A2(new_n11419_), .ZN(new_n11723_));
  NOR2_X1    g11467(.A1(new_n11720_), .A2(new_n11723_), .ZN(new_n11724_));
  NAND2_X1   g11468(.A1(new_n11724_), .A2(new_n11722_), .ZN(new_n11725_));
  AOI21_X1   g11469(.A1(new_n11725_), .A2(new_n11721_), .B(new_n11719_), .ZN(new_n11726_));
  NAND3_X1   g11470(.A1(new_n11725_), .A2(new_n11719_), .A3(new_n11721_), .ZN(new_n11727_));
  INV_X1     g11471(.I(new_n11727_), .ZN(new_n11728_));
  NOR3_X1    g11472(.A1(new_n11728_), .A2(new_n11714_), .A3(new_n11726_), .ZN(new_n11729_));
  INV_X1     g11473(.I(new_n11726_), .ZN(new_n11730_));
  AOI21_X1   g11474(.A1(new_n11730_), .A2(new_n11727_), .B(new_n11713_), .ZN(new_n11731_));
  NOR2_X1    g11475(.A1(new_n11731_), .A2(new_n11729_), .ZN(new_n11732_));
  INV_X1     g11476(.I(new_n11732_), .ZN(new_n11733_));
  AOI22_X1   g11477(.A1(new_n3267_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n3270_), .ZN(new_n11734_));
  OAI21_X1   g11478(.A1(new_n4022_), .A2(new_n3475_), .B(new_n11734_), .ZN(new_n11735_));
  AOI21_X1   g11479(.A1(new_n4223_), .A2(new_n3273_), .B(new_n11735_), .ZN(new_n11736_));
  XOR2_X1    g11480(.A1(new_n11736_), .A2(new_n3264_), .Z(new_n11737_));
  XOR2_X1    g11481(.A1(new_n11724_), .A2(new_n11722_), .Z(new_n11738_));
  NAND2_X1   g11482(.A1(new_n11738_), .A2(new_n11415_), .ZN(new_n11739_));
  NAND2_X1   g11483(.A1(new_n11739_), .A2(new_n11428_), .ZN(new_n11740_));
  NAND2_X1   g11484(.A1(new_n11740_), .A2(new_n11737_), .ZN(new_n11741_));
  INV_X1     g11485(.I(new_n11741_), .ZN(new_n11742_));
  NOR2_X1    g11486(.A1(new_n11740_), .A2(new_n11737_), .ZN(new_n11743_));
  NOR3_X1    g11487(.A1(new_n11742_), .A2(new_n11733_), .A3(new_n11743_), .ZN(new_n11744_));
  INV_X1     g11488(.I(new_n11743_), .ZN(new_n11745_));
  AOI21_X1   g11489(.A1(new_n11745_), .A2(new_n11741_), .B(new_n11732_), .ZN(new_n11746_));
  NOR2_X1    g11490(.A1(new_n11746_), .A2(new_n11744_), .ZN(new_n11747_));
  AOI22_X1   g11491(.A1(new_n2716_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n2719_), .ZN(new_n11748_));
  OAI21_X1   g11492(.A1(new_n4639_), .A2(new_n2924_), .B(new_n11748_), .ZN(new_n11749_));
  AOI21_X1   g11493(.A1(new_n5594_), .A2(new_n2722_), .B(new_n11749_), .ZN(new_n11750_));
  XOR2_X1    g11494(.A1(new_n11750_), .A2(new_n2714_), .Z(new_n11751_));
  NAND2_X1   g11495(.A1(new_n11442_), .A2(new_n11444_), .ZN(new_n11752_));
  NAND2_X1   g11496(.A1(new_n11752_), .A2(new_n11751_), .ZN(new_n11753_));
  OR2_X2     g11497(.A1(new_n11752_), .A2(new_n11751_), .Z(new_n11754_));
  NAND2_X1   g11498(.A1(new_n11754_), .A2(new_n11753_), .ZN(new_n11755_));
  XOR2_X1    g11499(.A1(new_n11755_), .A2(new_n11747_), .Z(new_n11756_));
  INV_X1     g11500(.I(new_n11756_), .ZN(new_n11757_));
  AOI22_X1   g11501(.A1(new_n2202_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n2205_), .ZN(new_n11758_));
  OAI21_X1   g11502(.A1(new_n5312_), .A2(new_n2370_), .B(new_n11758_), .ZN(new_n11759_));
  AOI21_X1   g11503(.A1(new_n6310_), .A2(new_n2208_), .B(new_n11759_), .ZN(new_n11760_));
  XOR2_X1    g11504(.A1(new_n11760_), .A2(\a[23] ), .Z(new_n11761_));
  NOR2_X1    g11505(.A1(new_n11461_), .A2(new_n11452_), .ZN(new_n11762_));
  NOR2_X1    g11506(.A1(new_n11762_), .A2(new_n11761_), .ZN(new_n11763_));
  AND2_X2    g11507(.A1(new_n11762_), .A2(new_n11761_), .Z(new_n11764_));
  NOR2_X1    g11508(.A1(new_n11764_), .A2(new_n11763_), .ZN(new_n11765_));
  XOR2_X1    g11509(.A1(new_n11765_), .A2(new_n11757_), .Z(new_n11766_));
  AOI22_X1   g11510(.A1(new_n1738_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n1743_), .ZN(new_n11767_));
  OAI21_X1   g11511(.A1(new_n6284_), .A2(new_n1931_), .B(new_n11767_), .ZN(new_n11768_));
  AOI21_X1   g11512(.A1(new_n7106_), .A2(new_n1746_), .B(new_n11768_), .ZN(new_n11769_));
  XOR2_X1    g11513(.A1(new_n11769_), .A2(new_n1736_), .Z(new_n11770_));
  NAND2_X1   g11514(.A1(new_n11472_), .A2(new_n11459_), .ZN(new_n11771_));
  NAND2_X1   g11515(.A1(new_n11771_), .A2(new_n11770_), .ZN(new_n11772_));
  INV_X1     g11516(.I(new_n11772_), .ZN(new_n11773_));
  NOR2_X1    g11517(.A1(new_n11771_), .A2(new_n11770_), .ZN(new_n11774_));
  NOR2_X1    g11518(.A1(new_n11773_), .A2(new_n11774_), .ZN(new_n11775_));
  NAND2_X1   g11519(.A1(new_n11775_), .A2(new_n11766_), .ZN(new_n11776_));
  INV_X1     g11520(.I(new_n11766_), .ZN(new_n11777_));
  INV_X1     g11521(.I(new_n11774_), .ZN(new_n11778_));
  NAND2_X1   g11522(.A1(new_n11778_), .A2(new_n11772_), .ZN(new_n11779_));
  NAND2_X1   g11523(.A1(new_n11779_), .A2(new_n11777_), .ZN(new_n11780_));
  NAND3_X1   g11524(.A1(new_n11776_), .A2(new_n11780_), .A3(new_n11589_), .ZN(new_n11781_));
  NOR2_X1    g11525(.A1(new_n11779_), .A2(new_n11777_), .ZN(new_n11782_));
  NOR2_X1    g11526(.A1(new_n11775_), .A2(new_n11766_), .ZN(new_n11783_));
  OAI21_X1   g11527(.A1(new_n11783_), .A2(new_n11782_), .B(new_n11588_), .ZN(new_n11784_));
  AOI21_X1   g11528(.A1(new_n11784_), .A2(new_n11781_), .B(new_n11584_), .ZN(new_n11785_));
  NOR3_X1    g11529(.A1(new_n11783_), .A2(new_n11782_), .A3(new_n11588_), .ZN(new_n11786_));
  AOI21_X1   g11530(.A1(new_n11776_), .A2(new_n11780_), .B(new_n11589_), .ZN(new_n11787_));
  NOR3_X1    g11531(.A1(new_n11787_), .A2(new_n11786_), .A3(new_n11583_), .ZN(new_n11788_));
  OAI22_X1   g11532(.A1(new_n993_), .A2(new_n8127_), .B1(new_n8126_), .B2(new_n997_), .ZN(new_n11789_));
  AOI21_X1   g11533(.A1(\b[46] ), .A2(new_n1486_), .B(new_n11789_), .ZN(new_n11790_));
  OAI21_X1   g11534(.A1(new_n8138_), .A2(new_n1323_), .B(new_n11790_), .ZN(new_n11791_));
  XOR2_X1    g11535(.A1(new_n11791_), .A2(\a[14] ), .Z(new_n11792_));
  INV_X1     g11536(.I(new_n11792_), .ZN(new_n11793_));
  NOR2_X1    g11537(.A1(new_n11495_), .A2(new_n11498_), .ZN(new_n11794_));
  NOR2_X1    g11538(.A1(new_n11794_), .A2(new_n11793_), .ZN(new_n11795_));
  NAND2_X1   g11539(.A1(new_n11503_), .A2(new_n11489_), .ZN(new_n11796_));
  NOR2_X1    g11540(.A1(new_n11796_), .A2(new_n11792_), .ZN(new_n11797_));
  NOR4_X1    g11541(.A1(new_n11795_), .A2(new_n11797_), .A3(new_n11785_), .A4(new_n11788_), .ZN(new_n11798_));
  NOR2_X1    g11542(.A1(new_n11788_), .A2(new_n11785_), .ZN(new_n11799_));
  NAND2_X1   g11543(.A1(new_n11796_), .A2(new_n11792_), .ZN(new_n11800_));
  NAND2_X1   g11544(.A1(new_n11794_), .A2(new_n11793_), .ZN(new_n11801_));
  AOI21_X1   g11545(.A1(new_n11801_), .A2(new_n11800_), .B(new_n11799_), .ZN(new_n11802_));
  NOR2_X1    g11546(.A1(new_n11798_), .A2(new_n11802_), .ZN(new_n11803_));
  NAND2_X1   g11547(.A1(new_n11803_), .A2(new_n11582_), .ZN(new_n11804_));
  OAI21_X1   g11548(.A1(new_n11798_), .A2(new_n11802_), .B(new_n11581_), .ZN(new_n11805_));
  AOI21_X1   g11549(.A1(new_n11804_), .A2(new_n11805_), .B(new_n11576_), .ZN(new_n11806_));
  NOR3_X1    g11550(.A1(new_n11798_), .A2(new_n11802_), .A3(new_n11581_), .ZN(new_n11807_));
  INV_X1     g11551(.I(new_n11805_), .ZN(new_n11808_));
  NOR3_X1    g11552(.A1(new_n11808_), .A2(new_n11575_), .A3(new_n11807_), .ZN(new_n11809_));
  NOR2_X1    g11553(.A1(new_n11806_), .A2(new_n11809_), .ZN(new_n11810_));
  INV_X1     g11554(.I(new_n11810_), .ZN(new_n11811_));
  AOI22_X1   g11555(.A1(new_n518_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n636_), .ZN(new_n11812_));
  OAI21_X1   g11556(.A1(new_n9032_), .A2(new_n917_), .B(new_n11812_), .ZN(new_n11813_));
  AOI21_X1   g11557(.A1(new_n10884_), .A2(new_n618_), .B(new_n11813_), .ZN(new_n11814_));
  XOR2_X1    g11558(.A1(new_n11814_), .A2(new_n488_), .Z(new_n11815_));
  INV_X1     g11559(.I(new_n11815_), .ZN(new_n11816_));
  AOI21_X1   g11560(.A1(new_n11525_), .A2(new_n11527_), .B(new_n11816_), .ZN(new_n11817_));
  NOR3_X1    g11561(.A1(new_n11554_), .A2(new_n11521_), .A3(new_n11815_), .ZN(new_n11818_));
  NOR3_X1    g11562(.A1(new_n11817_), .A2(new_n11811_), .A3(new_n11818_), .ZN(new_n11819_));
  OAI21_X1   g11563(.A1(new_n11554_), .A2(new_n11521_), .B(new_n11815_), .ZN(new_n11820_));
  NAND3_X1   g11564(.A1(new_n11525_), .A2(new_n11527_), .A3(new_n11816_), .ZN(new_n11821_));
  AOI21_X1   g11565(.A1(new_n11821_), .A2(new_n11820_), .B(new_n11810_), .ZN(new_n11822_));
  OAI21_X1   g11566(.A1(new_n11819_), .A2(new_n11822_), .B(new_n11573_), .ZN(new_n11823_));
  OAI21_X1   g11567(.A1(new_n11555_), .A2(new_n11554_), .B(new_n11557_), .ZN(new_n11824_));
  NAND2_X1   g11568(.A1(new_n11824_), .A2(new_n11556_), .ZN(new_n11825_));
  NAND3_X1   g11569(.A1(new_n11821_), .A2(new_n11820_), .A3(new_n11810_), .ZN(new_n11826_));
  OAI21_X1   g11570(.A1(new_n11817_), .A2(new_n11818_), .B(new_n11811_), .ZN(new_n11827_));
  NAND3_X1   g11571(.A1(new_n11827_), .A2(new_n11826_), .A3(new_n11825_), .ZN(new_n11828_));
  AOI22_X1   g11572(.A1(new_n267_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n261_), .ZN(new_n11829_));
  OAI21_X1   g11573(.A1(new_n11195_), .A2(new_n284_), .B(new_n11829_), .ZN(new_n11830_));
  XOR2_X1    g11574(.A1(\b[59] ), .A2(\b[60] ), .Z(new_n11831_));
  OAI21_X1   g11575(.A1(new_n11203_), .A2(new_n10625_), .B(new_n11195_), .ZN(new_n11832_));
  NAND2_X1   g11576(.A1(new_n11832_), .A2(\b[59] ), .ZN(new_n11833_));
  OAI21_X1   g11577(.A1(new_n11200_), .A2(\b[57] ), .B(\b[58] ), .ZN(new_n11834_));
  NAND2_X1   g11578(.A1(new_n11833_), .A2(new_n11834_), .ZN(new_n11835_));
  XOR2_X1    g11579(.A1(new_n11835_), .A2(new_n11831_), .Z(new_n11836_));
  AOI21_X1   g11580(.A1(new_n11836_), .A2(new_n265_), .B(new_n11830_), .ZN(new_n11837_));
  NOR2_X1    g11581(.A1(new_n11837_), .A2(new_n270_), .ZN(new_n11838_));
  INV_X1     g11582(.I(new_n11830_), .ZN(new_n11839_));
  XNOR2_X1   g11583(.A1(new_n11835_), .A2(new_n11831_), .ZN(new_n11840_));
  OAI21_X1   g11584(.A1(new_n11840_), .A2(new_n279_), .B(new_n11839_), .ZN(new_n11841_));
  NOR2_X1    g11585(.A1(new_n11841_), .A2(\a[2] ), .ZN(new_n11842_));
  AOI22_X1   g11586(.A1(new_n800_), .A2(\b[56] ), .B1(\b[57] ), .B2(new_n333_), .ZN(new_n11843_));
  OAI21_X1   g11587(.A1(new_n9972_), .A2(new_n392_), .B(new_n11843_), .ZN(new_n11844_));
  AOI21_X1   g11588(.A1(new_n10631_), .A2(new_n330_), .B(new_n11844_), .ZN(new_n11845_));
  XOR2_X1    g11589(.A1(new_n11845_), .A2(new_n312_), .Z(new_n11846_));
  INV_X1     g11590(.I(new_n11846_), .ZN(new_n11847_));
  OAI21_X1   g11591(.A1(new_n11842_), .A2(new_n11838_), .B(new_n11847_), .ZN(new_n11848_));
  NAND2_X1   g11592(.A1(new_n11841_), .A2(\a[2] ), .ZN(new_n11849_));
  NAND2_X1   g11593(.A1(new_n11837_), .A2(new_n270_), .ZN(new_n11850_));
  NAND3_X1   g11594(.A1(new_n11849_), .A2(new_n11850_), .A3(new_n11846_), .ZN(new_n11851_));
  NAND2_X1   g11595(.A1(new_n11848_), .A2(new_n11851_), .ZN(new_n11852_));
  AOI21_X1   g11596(.A1(new_n11823_), .A2(new_n11828_), .B(new_n11852_), .ZN(new_n11853_));
  AOI21_X1   g11597(.A1(new_n11827_), .A2(new_n11826_), .B(new_n11825_), .ZN(new_n11854_));
  NOR3_X1    g11598(.A1(new_n11819_), .A2(new_n11822_), .A3(new_n11573_), .ZN(new_n11855_));
  AOI21_X1   g11599(.A1(new_n11849_), .A2(new_n11850_), .B(new_n11846_), .ZN(new_n11856_));
  NOR3_X1    g11600(.A1(new_n11842_), .A2(new_n11838_), .A3(new_n11847_), .ZN(new_n11857_));
  NOR2_X1    g11601(.A1(new_n11856_), .A2(new_n11857_), .ZN(new_n11858_));
  NOR3_X1    g11602(.A1(new_n11855_), .A2(new_n11854_), .A3(new_n11858_), .ZN(new_n11859_));
  NOR2_X1    g11603(.A1(new_n11853_), .A2(new_n11859_), .ZN(new_n11860_));
  NOR3_X1    g11604(.A1(new_n11568_), .A2(new_n11565_), .A3(new_n11562_), .ZN(new_n11861_));
  AOI21_X1   g11605(.A1(new_n11192_), .A2(new_n11563_), .B(new_n11560_), .ZN(new_n11862_));
  NOR2_X1    g11606(.A1(new_n11862_), .A2(new_n11861_), .ZN(new_n11863_));
  NAND3_X1   g11607(.A1(new_n11225_), .A2(new_n11223_), .A3(new_n11863_), .ZN(new_n11864_));
  AOI21_X1   g11608(.A1(new_n11864_), .A2(new_n11564_), .B(new_n11860_), .ZN(new_n11865_));
  OAI21_X1   g11609(.A1(new_n11855_), .A2(new_n11854_), .B(new_n11858_), .ZN(new_n11866_));
  NAND3_X1   g11610(.A1(new_n11823_), .A2(new_n11828_), .A3(new_n11852_), .ZN(new_n11867_));
  NAND2_X1   g11611(.A1(new_n11866_), .A2(new_n11867_), .ZN(new_n11868_));
  AOI21_X1   g11612(.A1(new_n11219_), .A2(new_n11208_), .B(new_n11194_), .ZN(new_n11869_));
  NOR3_X1    g11613(.A1(new_n11869_), .A2(new_n11220_), .A3(new_n11570_), .ZN(new_n11870_));
  NOR3_X1    g11614(.A1(new_n11870_), .A2(new_n11861_), .A3(new_n11868_), .ZN(new_n11871_));
  NOR2_X1    g11615(.A1(new_n11871_), .A2(new_n11865_), .ZN(\f[60] ));
  AOI21_X1   g11616(.A1(new_n11576_), .A2(new_n11805_), .B(new_n11807_), .ZN(new_n11873_));
  NAND2_X1   g11617(.A1(new_n11800_), .A2(new_n11799_), .ZN(new_n11874_));
  NAND2_X1   g11618(.A1(new_n11874_), .A2(new_n11801_), .ZN(new_n11875_));
  OAI21_X1   g11619(.A1(new_n11583_), .A2(new_n11787_), .B(new_n11781_), .ZN(new_n11876_));
  NAND2_X1   g11620(.A1(new_n11766_), .A2(new_n11772_), .ZN(new_n11877_));
  NAND2_X1   g11621(.A1(new_n11877_), .A2(new_n11778_), .ZN(new_n11878_));
  NAND2_X1   g11622(.A1(new_n11762_), .A2(new_n11761_), .ZN(new_n11879_));
  OAI21_X1   g11623(.A1(new_n11756_), .A2(new_n11763_), .B(new_n11879_), .ZN(new_n11880_));
  INV_X1     g11624(.I(new_n11880_), .ZN(new_n11881_));
  AOI21_X1   g11625(.A1(new_n11732_), .A2(new_n11741_), .B(new_n11743_), .ZN(new_n11882_));
  INV_X1     g11626(.I(new_n11882_), .ZN(new_n11883_));
  OAI21_X1   g11627(.A1(new_n11714_), .A2(new_n11726_), .B(new_n11727_), .ZN(new_n11884_));
  NOR2_X1    g11628(.A1(new_n11699_), .A2(new_n11707_), .ZN(new_n11885_));
  NOR2_X1    g11629(.A1(new_n11885_), .A2(new_n11709_), .ZN(new_n11886_));
  NOR2_X1    g11630(.A1(new_n11884_), .A2(new_n11886_), .ZN(new_n11887_));
  INV_X1     g11631(.I(new_n11887_), .ZN(new_n11888_));
  NAND2_X1   g11632(.A1(new_n11884_), .A2(new_n11886_), .ZN(new_n11889_));
  AOI22_X1   g11633(.A1(new_n3864_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n3869_), .ZN(new_n11890_));
  OAI21_X1   g11634(.A1(new_n3592_), .A2(new_n5410_), .B(new_n11890_), .ZN(new_n11891_));
  AOI21_X1   g11635(.A1(new_n3796_), .A2(new_n3872_), .B(new_n11891_), .ZN(new_n11892_));
  XOR2_X1    g11636(.A1(new_n11892_), .A2(new_n3876_), .Z(new_n11893_));
  AOI22_X1   g11637(.A1(new_n4918_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n4921_), .ZN(new_n11894_));
  OAI21_X1   g11638(.A1(new_n3006_), .A2(new_n6099_), .B(new_n11894_), .ZN(new_n11895_));
  AOI21_X1   g11639(.A1(new_n3807_), .A2(new_n4699_), .B(new_n11895_), .ZN(new_n11896_));
  XOR2_X1    g11640(.A1(new_n11896_), .A2(new_n4446_), .Z(new_n11897_));
  AOI21_X1   g11641(.A1(new_n11695_), .A2(new_n11692_), .B(new_n11691_), .ZN(new_n11898_));
  OAI22_X1   g11642(.A1(new_n2646_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n2495_), .ZN(new_n11899_));
  AOI21_X1   g11643(.A1(\b[23] ), .A2(new_n5420_), .B(new_n11899_), .ZN(new_n11900_));
  OAI21_X1   g11644(.A1(new_n2655_), .A2(new_n6124_), .B(new_n11900_), .ZN(new_n11901_));
  XOR2_X1    g11645(.A1(new_n11901_), .A2(\a[38] ), .Z(new_n11902_));
  AOI22_X1   g11646(.A1(new_n6108_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n6111_), .ZN(new_n11903_));
  OAI21_X1   g11647(.A1(new_n1860_), .A2(new_n7708_), .B(new_n11903_), .ZN(new_n11904_));
  AOI21_X1   g11648(.A1(new_n2659_), .A2(new_n6105_), .B(new_n11904_), .ZN(new_n11905_));
  XOR2_X1    g11649(.A1(new_n11905_), .A2(new_n5849_), .Z(new_n11906_));
  AOI21_X1   g11650(.A1(new_n11667_), .A2(new_n11662_), .B(new_n11669_), .ZN(new_n11907_));
  AOI21_X1   g11651(.A1(new_n11645_), .A2(new_n11650_), .B(new_n11652_), .ZN(new_n11908_));
  INV_X1     g11652(.I(new_n11908_), .ZN(new_n11909_));
  NAND2_X1   g11653(.A1(new_n11640_), .A2(new_n11634_), .ZN(new_n11910_));
  NAND2_X1   g11654(.A1(new_n11910_), .A2(new_n11642_), .ZN(new_n11911_));
  OAI21_X1   g11655(.A1(new_n11607_), .A2(new_n11631_), .B(new_n11629_), .ZN(new_n11912_));
  AOI21_X1   g11656(.A1(new_n11311_), .A2(new_n11626_), .B(new_n11624_), .ZN(new_n11913_));
  INV_X1     g11657(.I(new_n11913_), .ZN(new_n11914_));
  AOI22_X1   g11658(.A1(new_n10981_), .A2(\b[4] ), .B1(new_n10979_), .B2(\b[3] ), .ZN(new_n11915_));
  OAI21_X1   g11659(.A1(new_n276_), .A2(new_n11306_), .B(new_n11915_), .ZN(new_n11916_));
  AOI21_X1   g11660(.A1(new_n1725_), .A2(new_n10984_), .B(new_n11916_), .ZN(new_n11917_));
  XOR2_X1    g11661(.A1(new_n11917_), .A2(new_n10989_), .Z(new_n11918_));
  INV_X1     g11662(.I(new_n11918_), .ZN(new_n11919_));
  INV_X1     g11663(.I(\a[61] ), .ZN(new_n11920_));
  NOR3_X1    g11664(.A1(new_n11920_), .A2(\a[59] ), .A3(\a[60] ), .ZN(new_n11921_));
  AND3_X2    g11665(.A1(new_n11920_), .A2(\a[59] ), .A3(\a[60] ), .Z(new_n11922_));
  NOR2_X1    g11666(.A1(new_n11922_), .A2(new_n11921_), .ZN(new_n11923_));
  INV_X1     g11667(.I(new_n11923_), .ZN(new_n11924_));
  XOR2_X1    g11668(.A1(\a[61] ), .A2(\a[62] ), .Z(new_n11925_));
  NOR2_X1    g11669(.A1(new_n11621_), .A2(new_n11925_), .ZN(new_n11926_));
  AOI22_X1   g11670(.A1(new_n11926_), .A2(\b[1] ), .B1(new_n11924_), .B2(\b[0] ), .ZN(new_n11927_));
  XNOR2_X1   g11671(.A1(\a[61] ), .A2(\a[62] ), .ZN(new_n11928_));
  NOR2_X1    g11672(.A1(new_n11621_), .A2(new_n11928_), .ZN(new_n11929_));
  INV_X1     g11673(.I(new_n11929_), .ZN(new_n11930_));
  OAI21_X1   g11674(.A1(new_n313_), .A2(new_n11930_), .B(new_n11927_), .ZN(new_n11931_));
  XOR2_X1    g11675(.A1(new_n11931_), .A2(\a[62] ), .Z(new_n11932_));
  NAND2_X1   g11676(.A1(new_n11623_), .A2(\a[62] ), .ZN(new_n11933_));
  XOR2_X1    g11677(.A1(new_n11932_), .A2(new_n11933_), .Z(new_n11934_));
  NOR2_X1    g11678(.A1(new_n11934_), .A2(new_n11919_), .ZN(new_n11935_));
  NAND2_X1   g11679(.A1(new_n11934_), .A2(new_n11919_), .ZN(new_n11936_));
  INV_X1     g11680(.I(new_n11936_), .ZN(new_n11937_));
  NOR2_X1    g11681(.A1(new_n11937_), .A2(new_n11935_), .ZN(new_n11938_));
  XOR2_X1    g11682(.A1(new_n11938_), .A2(new_n11914_), .Z(new_n11939_));
  OAI22_X1   g11683(.A1(new_n11298_), .A2(new_n471_), .B1(new_n438_), .B2(new_n11297_), .ZN(new_n11940_));
  AOI21_X1   g11684(.A1(\b[5] ), .A2(new_n11296_), .B(new_n11940_), .ZN(new_n11941_));
  OAI21_X1   g11685(.A1(new_n485_), .A2(new_n10069_), .B(new_n11941_), .ZN(new_n11942_));
  XOR2_X1    g11686(.A1(new_n11942_), .A2(\a[56] ), .Z(new_n11943_));
  OR2_X2     g11687(.A1(new_n11939_), .A2(new_n11943_), .Z(new_n11944_));
  NAND2_X1   g11688(.A1(new_n11939_), .A2(new_n11943_), .ZN(new_n11945_));
  NAND2_X1   g11689(.A1(new_n11944_), .A2(new_n11945_), .ZN(new_n11946_));
  XNOR2_X1   g11690(.A1(new_n11946_), .A2(new_n11912_), .ZN(new_n11947_));
  AOI22_X1   g11691(.A1(new_n9125_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n9123_), .ZN(new_n11948_));
  OAI21_X1   g11692(.A1(new_n577_), .A2(new_n9470_), .B(new_n11948_), .ZN(new_n11949_));
  AOI21_X1   g11693(.A1(new_n1059_), .A2(new_n9129_), .B(new_n11949_), .ZN(new_n11950_));
  XOR2_X1    g11694(.A1(new_n11950_), .A2(new_n9133_), .Z(new_n11951_));
  INV_X1     g11695(.I(new_n11951_), .ZN(new_n11952_));
  NAND2_X1   g11696(.A1(new_n11947_), .A2(new_n11952_), .ZN(new_n11953_));
  INV_X1     g11697(.I(new_n11947_), .ZN(new_n11954_));
  NAND2_X1   g11698(.A1(new_n11954_), .A2(new_n11951_), .ZN(new_n11955_));
  AND3_X2    g11699(.A1(new_n11911_), .A2(new_n11953_), .A3(new_n11955_), .Z(new_n11956_));
  AOI21_X1   g11700(.A1(new_n11953_), .A2(new_n11955_), .B(new_n11911_), .ZN(new_n11957_));
  NOR2_X1    g11701(.A1(new_n11956_), .A2(new_n11957_), .ZN(new_n11958_));
  OAI22_X1   g11702(.A1(new_n9461_), .A2(new_n1070_), .B1(new_n941_), .B2(new_n9462_), .ZN(new_n11959_));
  AOI21_X1   g11703(.A1(\b[11] ), .A2(new_n8575_), .B(new_n11959_), .ZN(new_n11960_));
  OAI21_X1   g11704(.A1(new_n1082_), .A2(new_n9460_), .B(new_n11960_), .ZN(new_n11961_));
  XOR2_X1    g11705(.A1(new_n11961_), .A2(\a[50] ), .Z(new_n11962_));
  INV_X1     g11706(.I(new_n11962_), .ZN(new_n11963_));
  NAND2_X1   g11707(.A1(new_n11958_), .A2(new_n11963_), .ZN(new_n11964_));
  INV_X1     g11708(.I(new_n11964_), .ZN(new_n11965_));
  NOR2_X1    g11709(.A1(new_n11958_), .A2(new_n11963_), .ZN(new_n11966_));
  OAI21_X1   g11710(.A1(new_n11965_), .A2(new_n11966_), .B(new_n11909_), .ZN(new_n11967_));
  NOR2_X1    g11711(.A1(new_n11965_), .A2(new_n11966_), .ZN(new_n11968_));
  NAND2_X1   g11712(.A1(new_n11968_), .A2(new_n11908_), .ZN(new_n11969_));
  AOI22_X1   g11713(.A1(new_n7403_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n7408_), .ZN(new_n11970_));
  OAI21_X1   g11714(.A1(new_n1093_), .A2(new_n9488_), .B(new_n11970_), .ZN(new_n11971_));
  AOI21_X1   g11715(.A1(new_n1701_), .A2(new_n7414_), .B(new_n11971_), .ZN(new_n11972_));
  XOR2_X1    g11716(.A1(new_n11972_), .A2(new_n7410_), .Z(new_n11973_));
  AOI21_X1   g11717(.A1(new_n11969_), .A2(new_n11967_), .B(new_n11973_), .ZN(new_n11974_));
  AND3_X2    g11718(.A1(new_n11969_), .A2(new_n11967_), .A3(new_n11973_), .Z(new_n11975_));
  NOR2_X1    g11719(.A1(new_n11975_), .A2(new_n11974_), .ZN(new_n11976_));
  XNOR2_X1   g11720(.A1(new_n11976_), .A2(new_n11907_), .ZN(new_n11977_));
  INV_X1     g11721(.I(new_n11977_), .ZN(new_n11978_));
  INV_X1     g11722(.I(new_n11675_), .ZN(new_n11979_));
  AOI22_X1   g11723(.A1(new_n6569_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n6574_), .ZN(new_n11980_));
  OAI21_X1   g11724(.A1(new_n1432_), .A2(new_n8565_), .B(new_n11980_), .ZN(new_n11981_));
  AOI21_X1   g11725(.A1(new_n1695_), .A2(new_n6579_), .B(new_n11981_), .ZN(new_n11982_));
  XOR2_X1    g11726(.A1(new_n11982_), .A2(new_n6567_), .Z(new_n11983_));
  INV_X1     g11727(.I(new_n11983_), .ZN(new_n11984_));
  AOI21_X1   g11728(.A1(new_n11676_), .A2(new_n11979_), .B(new_n11984_), .ZN(new_n11985_));
  NOR3_X1    g11729(.A1(new_n11677_), .A2(new_n11596_), .A3(new_n11600_), .ZN(new_n11986_));
  NOR3_X1    g11730(.A1(new_n11986_), .A2(new_n11675_), .A3(new_n11983_), .ZN(new_n11987_));
  NOR3_X1    g11731(.A1(new_n11987_), .A2(new_n11985_), .A3(new_n11978_), .ZN(new_n11988_));
  OAI21_X1   g11732(.A1(new_n11986_), .A2(new_n11675_), .B(new_n11983_), .ZN(new_n11989_));
  NAND3_X1   g11733(.A1(new_n11676_), .A2(new_n11979_), .A3(new_n11984_), .ZN(new_n11990_));
  AOI21_X1   g11734(.A1(new_n11989_), .A2(new_n11990_), .B(new_n11977_), .ZN(new_n11991_));
  NOR3_X1    g11735(.A1(new_n11988_), .A2(new_n11991_), .A3(new_n11906_), .ZN(new_n11992_));
  INV_X1     g11736(.I(new_n11906_), .ZN(new_n11993_));
  NAND3_X1   g11737(.A1(new_n11989_), .A2(new_n11990_), .A3(new_n11977_), .ZN(new_n11994_));
  OAI21_X1   g11738(.A1(new_n11987_), .A2(new_n11985_), .B(new_n11978_), .ZN(new_n11995_));
  AOI21_X1   g11739(.A1(new_n11995_), .A2(new_n11994_), .B(new_n11993_), .ZN(new_n11996_));
  NOR2_X1    g11740(.A1(new_n11992_), .A2(new_n11996_), .ZN(new_n11997_));
  OAI21_X1   g11741(.A1(new_n11590_), .A2(new_n11682_), .B(new_n11680_), .ZN(new_n11998_));
  NAND2_X1   g11742(.A1(new_n11997_), .A2(new_n11998_), .ZN(new_n11999_));
  NAND3_X1   g11743(.A1(new_n11995_), .A2(new_n11994_), .A3(new_n11993_), .ZN(new_n12000_));
  OAI21_X1   g11744(.A1(new_n11988_), .A2(new_n11991_), .B(new_n11906_), .ZN(new_n12001_));
  NAND2_X1   g11745(.A1(new_n12001_), .A2(new_n12000_), .ZN(new_n12002_));
  INV_X1     g11746(.I(new_n11998_), .ZN(new_n12003_));
  NAND2_X1   g11747(.A1(new_n12002_), .A2(new_n12003_), .ZN(new_n12004_));
  NAND3_X1   g11748(.A1(new_n11999_), .A2(new_n12004_), .A3(new_n11902_), .ZN(new_n12005_));
  AOI21_X1   g11749(.A1(new_n11999_), .A2(new_n12004_), .B(new_n11902_), .ZN(new_n12006_));
  INV_X1     g11750(.I(new_n12006_), .ZN(new_n12007_));
  NAND2_X1   g11751(.A1(new_n12007_), .A2(new_n12005_), .ZN(new_n12008_));
  NAND2_X1   g11752(.A1(new_n12008_), .A2(new_n11898_), .ZN(new_n12009_));
  OAI21_X1   g11753(.A1(new_n11684_), .A2(new_n11693_), .B(new_n11696_), .ZN(new_n12010_));
  INV_X1     g11754(.I(new_n11902_), .ZN(new_n12011_));
  NOR2_X1    g11755(.A1(new_n12002_), .A2(new_n12003_), .ZN(new_n12012_));
  NOR2_X1    g11756(.A1(new_n11997_), .A2(new_n11998_), .ZN(new_n12013_));
  NOR3_X1    g11757(.A1(new_n12013_), .A2(new_n12012_), .A3(new_n12011_), .ZN(new_n12014_));
  NOR2_X1    g11758(.A1(new_n12006_), .A2(new_n12014_), .ZN(new_n12015_));
  NAND2_X1   g11759(.A1(new_n12015_), .A2(new_n12010_), .ZN(new_n12016_));
  NAND3_X1   g11760(.A1(new_n12009_), .A2(new_n11897_), .A3(new_n12016_), .ZN(new_n12017_));
  INV_X1     g11761(.I(new_n11897_), .ZN(new_n12018_));
  NOR2_X1    g11762(.A1(new_n12015_), .A2(new_n12010_), .ZN(new_n12019_));
  NOR2_X1    g11763(.A1(new_n12008_), .A2(new_n11898_), .ZN(new_n12020_));
  OAI21_X1   g11764(.A1(new_n12020_), .A2(new_n12019_), .B(new_n12018_), .ZN(new_n12021_));
  NAND2_X1   g11765(.A1(new_n12021_), .A2(new_n12017_), .ZN(new_n12022_));
  XOR2_X1    g11766(.A1(new_n12022_), .A2(new_n11893_), .Z(new_n12023_));
  AOI21_X1   g11767(.A1(new_n11888_), .A2(new_n11889_), .B(new_n12023_), .ZN(new_n12024_));
  INV_X1     g11768(.I(new_n11889_), .ZN(new_n12025_));
  INV_X1     g11769(.I(new_n12023_), .ZN(new_n12026_));
  NOR3_X1    g11770(.A1(new_n12025_), .A2(new_n11887_), .A3(new_n12026_), .ZN(new_n12027_));
  AOI22_X1   g11771(.A1(new_n3267_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n3270_), .ZN(new_n12028_));
  OAI21_X1   g11772(.A1(new_n4023_), .A2(new_n3475_), .B(new_n12028_), .ZN(new_n12029_));
  AOI21_X1   g11773(.A1(new_n5103_), .A2(new_n3273_), .B(new_n12029_), .ZN(new_n12030_));
  XOR2_X1    g11774(.A1(new_n12030_), .A2(new_n3264_), .Z(new_n12031_));
  INV_X1     g11775(.I(new_n12031_), .ZN(new_n12032_));
  OAI21_X1   g11776(.A1(new_n12024_), .A2(new_n12027_), .B(new_n12032_), .ZN(new_n12033_));
  OAI21_X1   g11777(.A1(new_n12025_), .A2(new_n11887_), .B(new_n12026_), .ZN(new_n12034_));
  NAND3_X1   g11778(.A1(new_n11888_), .A2(new_n11889_), .A3(new_n12023_), .ZN(new_n12035_));
  NAND3_X1   g11779(.A1(new_n12034_), .A2(new_n12035_), .A3(new_n12031_), .ZN(new_n12036_));
  NAND3_X1   g11780(.A1(new_n11883_), .A2(new_n12033_), .A3(new_n12036_), .ZN(new_n12037_));
  AOI21_X1   g11781(.A1(new_n12034_), .A2(new_n12035_), .B(new_n12031_), .ZN(new_n12038_));
  NOR3_X1    g11782(.A1(new_n12024_), .A2(new_n12027_), .A3(new_n12032_), .ZN(new_n12039_));
  OAI21_X1   g11783(.A1(new_n12038_), .A2(new_n12039_), .B(new_n11882_), .ZN(new_n12040_));
  OAI22_X1   g11784(.A1(new_n2703_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n2708_), .ZN(new_n12041_));
  AOI21_X1   g11785(.A1(\b[35] ), .A2(new_n2906_), .B(new_n12041_), .ZN(new_n12042_));
  OAI21_X1   g11786(.A1(new_n5322_), .A2(new_n2711_), .B(new_n12042_), .ZN(new_n12043_));
  XOR2_X1    g11787(.A1(new_n12043_), .A2(\a[26] ), .Z(new_n12044_));
  INV_X1     g11788(.I(new_n12044_), .ZN(new_n12045_));
  NAND3_X1   g11789(.A1(new_n12037_), .A2(new_n12040_), .A3(new_n12045_), .ZN(new_n12046_));
  NOR3_X1    g11790(.A1(new_n12038_), .A2(new_n12039_), .A3(new_n11882_), .ZN(new_n12047_));
  AOI21_X1   g11791(.A1(new_n12033_), .A2(new_n12036_), .B(new_n11883_), .ZN(new_n12048_));
  OAI21_X1   g11792(.A1(new_n12048_), .A2(new_n12047_), .B(new_n12044_), .ZN(new_n12049_));
  NAND2_X1   g11793(.A1(new_n12049_), .A2(new_n12046_), .ZN(new_n12050_));
  NAND2_X1   g11794(.A1(new_n11753_), .A2(new_n11747_), .ZN(new_n12051_));
  AND2_X2    g11795(.A1(new_n12051_), .A2(new_n11754_), .Z(new_n12052_));
  AOI22_X1   g11796(.A1(new_n2202_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n2205_), .ZN(new_n12053_));
  OAI21_X1   g11797(.A1(new_n5341_), .A2(new_n2370_), .B(new_n12053_), .ZN(new_n12054_));
  AOI21_X1   g11798(.A1(new_n5793_), .A2(new_n2208_), .B(new_n12054_), .ZN(new_n12055_));
  XOR2_X1    g11799(.A1(new_n12055_), .A2(new_n2200_), .Z(new_n12056_));
  INV_X1     g11800(.I(new_n12056_), .ZN(new_n12057_));
  NAND2_X1   g11801(.A1(new_n12052_), .A2(new_n12057_), .ZN(new_n12058_));
  NAND2_X1   g11802(.A1(new_n12051_), .A2(new_n11754_), .ZN(new_n12059_));
  NAND2_X1   g11803(.A1(new_n12059_), .A2(new_n12056_), .ZN(new_n12060_));
  AOI21_X1   g11804(.A1(new_n12058_), .A2(new_n12060_), .B(new_n12050_), .ZN(new_n12061_));
  INV_X1     g11805(.I(new_n12050_), .ZN(new_n12062_));
  NOR2_X1    g11806(.A1(new_n12059_), .A2(new_n12056_), .ZN(new_n12063_));
  INV_X1     g11807(.I(new_n12060_), .ZN(new_n12064_));
  NOR3_X1    g11808(.A1(new_n12064_), .A2(new_n12062_), .A3(new_n12063_), .ZN(new_n12065_));
  OR2_X2     g11809(.A1(new_n12065_), .A2(new_n12061_), .Z(new_n12066_));
  NAND2_X1   g11810(.A1(new_n12066_), .A2(new_n11881_), .ZN(new_n12067_));
  NOR2_X1    g11811(.A1(new_n12065_), .A2(new_n12061_), .ZN(new_n12068_));
  NAND2_X1   g11812(.A1(new_n12068_), .A2(new_n11880_), .ZN(new_n12069_));
  OAI22_X1   g11813(.A1(new_n1751_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n1754_), .ZN(new_n12070_));
  AOI21_X1   g11814(.A1(\b[41] ), .A2(new_n1939_), .B(new_n12070_), .ZN(new_n12071_));
  OAI21_X1   g11815(.A1(new_n6785_), .A2(new_n1757_), .B(new_n12071_), .ZN(new_n12072_));
  XOR2_X1    g11816(.A1(new_n12072_), .A2(\a[20] ), .Z(new_n12073_));
  INV_X1     g11817(.I(new_n12073_), .ZN(new_n12074_));
  NAND3_X1   g11818(.A1(new_n12067_), .A2(new_n12069_), .A3(new_n12074_), .ZN(new_n12075_));
  NAND2_X1   g11819(.A1(new_n12067_), .A2(new_n12069_), .ZN(new_n12076_));
  NAND2_X1   g11820(.A1(new_n12076_), .A2(new_n12073_), .ZN(new_n12077_));
  NAND2_X1   g11821(.A1(new_n12077_), .A2(new_n12075_), .ZN(new_n12078_));
  NAND2_X1   g11822(.A1(new_n12078_), .A2(new_n11878_), .ZN(new_n12079_));
  AOI21_X1   g11823(.A1(new_n11766_), .A2(new_n11772_), .B(new_n11774_), .ZN(new_n12080_));
  INV_X1     g11824(.I(new_n12075_), .ZN(new_n12081_));
  AOI21_X1   g11825(.A1(new_n12067_), .A2(new_n12069_), .B(new_n12074_), .ZN(new_n12082_));
  NOR2_X1    g11826(.A1(new_n12081_), .A2(new_n12082_), .ZN(new_n12083_));
  NAND2_X1   g11827(.A1(new_n12083_), .A2(new_n12080_), .ZN(new_n12084_));
  OAI22_X1   g11828(.A1(new_n1592_), .A2(new_n7617_), .B1(new_n7096_), .B2(new_n1505_), .ZN(new_n12085_));
  AOI21_X1   g11829(.A1(\b[44] ), .A2(new_n1584_), .B(new_n12085_), .ZN(new_n12086_));
  OAI21_X1   g11830(.A1(new_n7627_), .A2(new_n1732_), .B(new_n12086_), .ZN(new_n12087_));
  XOR2_X1    g11831(.A1(new_n12087_), .A2(\a[17] ), .Z(new_n12088_));
  AOI21_X1   g11832(.A1(new_n12084_), .A2(new_n12079_), .B(new_n12088_), .ZN(new_n12089_));
  NOR2_X1    g11833(.A1(new_n12083_), .A2(new_n12080_), .ZN(new_n12090_));
  NOR2_X1    g11834(.A1(new_n12078_), .A2(new_n11878_), .ZN(new_n12091_));
  INV_X1     g11835(.I(new_n12088_), .ZN(new_n12092_));
  NOR3_X1    g11836(.A1(new_n12090_), .A2(new_n12091_), .A3(new_n12092_), .ZN(new_n12093_));
  NOR2_X1    g11837(.A1(new_n12089_), .A2(new_n12093_), .ZN(new_n12094_));
  NAND2_X1   g11838(.A1(new_n12094_), .A2(new_n11876_), .ZN(new_n12095_));
  INV_X1     g11839(.I(new_n11876_), .ZN(new_n12096_));
  OAI21_X1   g11840(.A1(new_n12090_), .A2(new_n12091_), .B(new_n12092_), .ZN(new_n12097_));
  NAND3_X1   g11841(.A1(new_n12084_), .A2(new_n12079_), .A3(new_n12088_), .ZN(new_n12098_));
  NAND2_X1   g11842(.A1(new_n12097_), .A2(new_n12098_), .ZN(new_n12099_));
  NAND2_X1   g11843(.A1(new_n12099_), .A2(new_n12096_), .ZN(new_n12100_));
  NAND2_X1   g11844(.A1(new_n12095_), .A2(new_n12100_), .ZN(new_n12101_));
  OAI22_X1   g11845(.A1(new_n993_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n997_), .ZN(new_n12102_));
  AOI21_X1   g11846(.A1(\b[47] ), .A2(new_n1486_), .B(new_n12102_), .ZN(new_n12103_));
  OAI21_X1   g11847(.A1(new_n9050_), .A2(new_n1323_), .B(new_n12103_), .ZN(new_n12104_));
  XOR2_X1    g11848(.A1(new_n12104_), .A2(\a[14] ), .Z(new_n12105_));
  NOR2_X1    g11849(.A1(new_n12101_), .A2(new_n12105_), .ZN(new_n12106_));
  NOR2_X1    g11850(.A1(new_n12099_), .A2(new_n12096_), .ZN(new_n12107_));
  NOR2_X1    g11851(.A1(new_n12094_), .A2(new_n11876_), .ZN(new_n12108_));
  NOR2_X1    g11852(.A1(new_n12108_), .A2(new_n12107_), .ZN(new_n12109_));
  INV_X1     g11853(.I(new_n12105_), .ZN(new_n12110_));
  NOR2_X1    g11854(.A1(new_n12109_), .A2(new_n12110_), .ZN(new_n12111_));
  NOR2_X1    g11855(.A1(new_n12111_), .A2(new_n12106_), .ZN(new_n12112_));
  NAND2_X1   g11856(.A1(new_n12112_), .A2(new_n11875_), .ZN(new_n12113_));
  NAND2_X1   g11857(.A1(new_n12109_), .A2(new_n12110_), .ZN(new_n12114_));
  NAND2_X1   g11858(.A1(new_n12101_), .A2(new_n12105_), .ZN(new_n12115_));
  NAND2_X1   g11859(.A1(new_n12114_), .A2(new_n12115_), .ZN(new_n12116_));
  NAND3_X1   g11860(.A1(new_n12116_), .A2(new_n11801_), .A3(new_n11874_), .ZN(new_n12117_));
  OAI22_X1   g11861(.A1(new_n713_), .A2(new_n9032_), .B1(new_n8776_), .B2(new_n717_), .ZN(new_n12118_));
  AOI21_X1   g11862(.A1(\b[50] ), .A2(new_n1126_), .B(new_n12118_), .ZN(new_n12119_));
  OAI21_X1   g11863(.A1(new_n9043_), .A2(new_n986_), .B(new_n12119_), .ZN(new_n12120_));
  XOR2_X1    g11864(.A1(new_n12120_), .A2(\a[11] ), .Z(new_n12121_));
  INV_X1     g11865(.I(new_n12121_), .ZN(new_n12122_));
  NAND3_X1   g11866(.A1(new_n12117_), .A2(new_n12113_), .A3(new_n12122_), .ZN(new_n12123_));
  AOI21_X1   g11867(.A1(new_n11801_), .A2(new_n11874_), .B(new_n12116_), .ZN(new_n12124_));
  NOR2_X1    g11868(.A1(new_n12112_), .A2(new_n11875_), .ZN(new_n12125_));
  OAI21_X1   g11869(.A1(new_n12124_), .A2(new_n12125_), .B(new_n12121_), .ZN(new_n12126_));
  NAND2_X1   g11870(.A1(new_n12126_), .A2(new_n12123_), .ZN(new_n12127_));
  NOR2_X1    g11871(.A1(new_n12127_), .A2(new_n11873_), .ZN(new_n12128_));
  INV_X1     g11872(.I(new_n11873_), .ZN(new_n12129_));
  NOR3_X1    g11873(.A1(new_n12124_), .A2(new_n12125_), .A3(new_n12121_), .ZN(new_n12130_));
  AOI21_X1   g11874(.A1(new_n12117_), .A2(new_n12113_), .B(new_n12122_), .ZN(new_n12131_));
  NOR2_X1    g11875(.A1(new_n12130_), .A2(new_n12131_), .ZN(new_n12132_));
  NOR2_X1    g11876(.A1(new_n12132_), .A2(new_n12129_), .ZN(new_n12133_));
  AOI22_X1   g11877(.A1(new_n518_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n636_), .ZN(new_n12134_));
  OAI21_X1   g11878(.A1(new_n9376_), .A2(new_n917_), .B(new_n12134_), .ZN(new_n12135_));
  AOI21_X1   g11879(.A1(new_n9979_), .A2(new_n618_), .B(new_n12135_), .ZN(new_n12136_));
  XOR2_X1    g11880(.A1(new_n12136_), .A2(new_n488_), .Z(new_n12137_));
  NOR3_X1    g11881(.A1(new_n12133_), .A2(new_n12128_), .A3(new_n12137_), .ZN(new_n12138_));
  NOR2_X1    g11882(.A1(new_n12133_), .A2(new_n12128_), .ZN(new_n12139_));
  INV_X1     g11883(.I(new_n12137_), .ZN(new_n12140_));
  NOR2_X1    g11884(.A1(new_n12139_), .A2(new_n12140_), .ZN(new_n12141_));
  AOI21_X1   g11885(.A1(new_n11810_), .A2(new_n11820_), .B(new_n11818_), .ZN(new_n12142_));
  NOR3_X1    g11886(.A1(new_n12141_), .A2(new_n12138_), .A3(new_n12142_), .ZN(new_n12143_));
  INV_X1     g11887(.I(new_n12143_), .ZN(new_n12144_));
  OAI21_X1   g11888(.A1(new_n12141_), .A2(new_n12138_), .B(new_n12142_), .ZN(new_n12145_));
  NAND2_X1   g11889(.A1(new_n12144_), .A2(new_n12145_), .ZN(new_n12146_));
  INV_X1     g11890(.I(\b[60] ), .ZN(new_n12147_));
  INV_X1     g11891(.I(\b[61] ), .ZN(new_n12148_));
  OAI22_X1   g11892(.A1(new_n277_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n262_), .ZN(new_n12149_));
  AOI21_X1   g11893(.A1(\b[59] ), .A2(new_n283_), .B(new_n12149_), .ZN(new_n12150_));
  INV_X1     g11894(.I(\b[59] ), .ZN(new_n12151_));
  AOI21_X1   g11895(.A1(new_n11835_), .A2(\b[60] ), .B(new_n12151_), .ZN(new_n12152_));
  NOR2_X1    g11896(.A1(new_n11835_), .A2(\b[60] ), .ZN(new_n12153_));
  NOR2_X1    g11897(.A1(new_n12152_), .A2(new_n12153_), .ZN(new_n12154_));
  NAND3_X1   g11898(.A1(new_n11833_), .A2(new_n11834_), .A3(new_n12148_), .ZN(new_n12155_));
  NAND2_X1   g11899(.A1(new_n11835_), .A2(\b[61] ), .ZN(new_n12156_));
  AND2_X2    g11900(.A1(new_n12156_), .A2(new_n12155_), .Z(new_n12157_));
  OR2_X2     g11901(.A1(new_n12157_), .A2(new_n12154_), .Z(new_n12158_));
  NAND2_X1   g11902(.A1(new_n12157_), .A2(new_n12154_), .ZN(new_n12159_));
  NAND3_X1   g11903(.A1(new_n12158_), .A2(new_n265_), .A3(new_n12159_), .ZN(new_n12160_));
  NAND2_X1   g11904(.A1(new_n12160_), .A2(new_n12150_), .ZN(new_n12161_));
  NAND2_X1   g11905(.A1(new_n12161_), .A2(\a[2] ), .ZN(new_n12162_));
  NAND3_X1   g11906(.A1(new_n12160_), .A2(new_n270_), .A3(new_n12150_), .ZN(new_n12163_));
  INV_X1     g11907(.I(new_n11206_), .ZN(new_n12164_));
  AOI22_X1   g11908(.A1(new_n800_), .A2(\b[57] ), .B1(\b[58] ), .B2(new_n333_), .ZN(new_n12165_));
  OAI21_X1   g11909(.A1(new_n10308_), .A2(new_n392_), .B(new_n12165_), .ZN(new_n12166_));
  AOI21_X1   g11910(.A1(new_n12164_), .A2(new_n330_), .B(new_n12166_), .ZN(new_n12167_));
  XOR2_X1    g11911(.A1(new_n12167_), .A2(new_n312_), .Z(new_n12168_));
  AOI21_X1   g11912(.A1(new_n12162_), .A2(new_n12163_), .B(new_n12168_), .ZN(new_n12169_));
  NAND3_X1   g11913(.A1(new_n12162_), .A2(new_n12163_), .A3(new_n12168_), .ZN(new_n12170_));
  INV_X1     g11914(.I(new_n12170_), .ZN(new_n12171_));
  NOR2_X1    g11915(.A1(new_n12171_), .A2(new_n12169_), .ZN(new_n12172_));
  NAND2_X1   g11916(.A1(new_n12146_), .A2(new_n12172_), .ZN(new_n12173_));
  INV_X1     g11917(.I(new_n12145_), .ZN(new_n12174_));
  NOR2_X1    g11918(.A1(new_n12174_), .A2(new_n12143_), .ZN(new_n12175_));
  INV_X1     g11919(.I(new_n12169_), .ZN(new_n12176_));
  NAND2_X1   g11920(.A1(new_n12176_), .A2(new_n12170_), .ZN(new_n12177_));
  NAND2_X1   g11921(.A1(new_n12175_), .A2(new_n12177_), .ZN(new_n12178_));
  NAND2_X1   g11922(.A1(new_n12178_), .A2(new_n12173_), .ZN(new_n12179_));
  NOR2_X1    g11923(.A1(new_n11819_), .A2(new_n11822_), .ZN(new_n12180_));
  AOI21_X1   g11924(.A1(new_n12180_), .A2(new_n11851_), .B(new_n11856_), .ZN(new_n12181_));
  NAND2_X1   g11925(.A1(new_n12180_), .A2(new_n11858_), .ZN(new_n12182_));
  OAI21_X1   g11926(.A1(new_n11819_), .A2(new_n11822_), .B(new_n11852_), .ZN(new_n12183_));
  AOI21_X1   g11927(.A1(new_n12183_), .A2(new_n12182_), .B(new_n11825_), .ZN(new_n12184_));
  OAI21_X1   g11928(.A1(new_n11865_), .A2(new_n12184_), .B(new_n12181_), .ZN(new_n12185_));
  OAI21_X1   g11929(.A1(new_n11870_), .A2(new_n11861_), .B(new_n11868_), .ZN(new_n12186_));
  INV_X1     g11930(.I(new_n12181_), .ZN(new_n12187_));
  INV_X1     g11931(.I(new_n12184_), .ZN(new_n12188_));
  NAND3_X1   g11932(.A1(new_n12186_), .A2(new_n12187_), .A3(new_n12188_), .ZN(new_n12189_));
  NAND2_X1   g11933(.A1(new_n12185_), .A2(new_n12189_), .ZN(new_n12190_));
  XOR2_X1    g11934(.A1(new_n12190_), .A2(new_n12179_), .Z(\f[61] ));
  NOR2_X1    g11935(.A1(new_n12175_), .A2(new_n12177_), .ZN(new_n12192_));
  NOR2_X1    g11936(.A1(new_n12146_), .A2(new_n12172_), .ZN(new_n12193_));
  NOR2_X1    g11937(.A1(new_n12192_), .A2(new_n12193_), .ZN(new_n12194_));
  AOI21_X1   g11938(.A1(new_n12186_), .A2(new_n12188_), .B(new_n12187_), .ZN(new_n12195_));
  OAI21_X1   g11939(.A1(new_n12194_), .A2(new_n12195_), .B(new_n12189_), .ZN(new_n12196_));
  OAI21_X1   g11940(.A1(new_n12146_), .A2(new_n12171_), .B(new_n12176_), .ZN(new_n12197_));
  INV_X1     g11941(.I(new_n12197_), .ZN(new_n12198_));
  INV_X1     g11942(.I(new_n12138_), .ZN(new_n12199_));
  INV_X1     g11943(.I(new_n12142_), .ZN(new_n12200_));
  OAI21_X1   g11944(.A1(new_n12139_), .A2(new_n12140_), .B(new_n12200_), .ZN(new_n12201_));
  NAND2_X1   g11945(.A1(new_n12201_), .A2(new_n12199_), .ZN(new_n12202_));
  NAND2_X1   g11946(.A1(new_n11540_), .A2(new_n11534_), .ZN(new_n12203_));
  OAI22_X1   g11947(.A1(new_n321_), .A2(new_n12151_), .B1(new_n325_), .B2(new_n11195_), .ZN(new_n12204_));
  AOI21_X1   g11948(.A1(\b[57] ), .A2(new_n602_), .B(new_n12204_), .ZN(new_n12205_));
  OAI21_X1   g11949(.A1(new_n12203_), .A2(new_n318_), .B(new_n12205_), .ZN(new_n12206_));
  XOR2_X1    g11950(.A1(new_n12206_), .A2(new_n312_), .Z(new_n12207_));
  AOI22_X1   g11951(.A1(new_n518_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n636_), .ZN(new_n12208_));
  OAI21_X1   g11952(.A1(new_n9942_), .A2(new_n917_), .B(new_n12208_), .ZN(new_n12209_));
  AOI21_X1   g11953(.A1(new_n10318_), .A2(new_n618_), .B(new_n12209_), .ZN(new_n12210_));
  XOR2_X1    g11954(.A1(new_n12210_), .A2(new_n488_), .Z(new_n12211_));
  INV_X1     g11955(.I(new_n12211_), .ZN(new_n12212_));
  NAND2_X1   g11956(.A1(new_n12207_), .A2(new_n12212_), .ZN(new_n12213_));
  XOR2_X1    g11957(.A1(new_n12206_), .A2(\a[5] ), .Z(new_n12214_));
  NAND2_X1   g11958(.A1(new_n12214_), .A2(new_n12211_), .ZN(new_n12215_));
  NAND2_X1   g11959(.A1(new_n12213_), .A2(new_n12215_), .ZN(new_n12216_));
  INV_X1     g11960(.I(new_n12216_), .ZN(new_n12217_));
  OAI21_X1   g11961(.A1(new_n11873_), .A2(new_n12131_), .B(new_n12123_), .ZN(new_n12218_));
  INV_X1     g11962(.I(new_n12218_), .ZN(new_n12219_));
  OAI22_X1   g11963(.A1(new_n713_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n717_), .ZN(new_n12220_));
  AOI21_X1   g11964(.A1(\b[51] ), .A2(new_n1126_), .B(new_n12220_), .ZN(new_n12221_));
  OAI21_X1   g11965(.A1(new_n9385_), .A2(new_n986_), .B(new_n12221_), .ZN(new_n12222_));
  XOR2_X1    g11966(.A1(new_n12222_), .A2(\a[11] ), .Z(new_n12223_));
  INV_X1     g11967(.I(new_n12223_), .ZN(new_n12224_));
  AOI21_X1   g11968(.A1(new_n11801_), .A2(new_n11874_), .B(new_n12111_), .ZN(new_n12225_));
  OAI22_X1   g11969(.A1(new_n993_), .A2(new_n8500_), .B1(new_n8168_), .B2(new_n997_), .ZN(new_n12226_));
  AOI21_X1   g11970(.A1(\b[48] ), .A2(new_n1486_), .B(new_n12226_), .ZN(new_n12227_));
  OAI21_X1   g11971(.A1(new_n8510_), .A2(new_n1323_), .B(new_n12227_), .ZN(new_n12228_));
  XOR2_X1    g11972(.A1(new_n12228_), .A2(\a[14] ), .Z(new_n12229_));
  INV_X1     g11973(.I(new_n12229_), .ZN(new_n12230_));
  AOI21_X1   g11974(.A1(new_n11876_), .A2(new_n12098_), .B(new_n12089_), .ZN(new_n12231_));
  OAI22_X1   g11975(.A1(new_n1592_), .A2(new_n8126_), .B1(new_n7617_), .B2(new_n1505_), .ZN(new_n12232_));
  AOI21_X1   g11976(.A1(\b[45] ), .A2(new_n1584_), .B(new_n12232_), .ZN(new_n12233_));
  OAI21_X1   g11977(.A1(new_n11237_), .A2(new_n1732_), .B(new_n12233_), .ZN(new_n12234_));
  XOR2_X1    g11978(.A1(new_n12234_), .A2(\a[17] ), .Z(new_n12235_));
  NAND2_X1   g11979(.A1(new_n11878_), .A2(new_n12077_), .ZN(new_n12236_));
  NAND2_X1   g11980(.A1(new_n11880_), .A2(new_n12057_), .ZN(new_n12237_));
  XNOR2_X1   g11981(.A1(new_n12050_), .A2(new_n12059_), .ZN(new_n12238_));
  OAI21_X1   g11982(.A1(new_n11880_), .A2(new_n12057_), .B(new_n12238_), .ZN(new_n12239_));
  OAI22_X1   g11983(.A1(new_n2189_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n2194_), .ZN(new_n12240_));
  AOI21_X1   g11984(.A1(\b[39] ), .A2(new_n2361_), .B(new_n12240_), .ZN(new_n12241_));
  OAI21_X1   g11985(.A1(new_n6299_), .A2(new_n2197_), .B(new_n12241_), .ZN(new_n12242_));
  XOR2_X1    g11986(.A1(new_n12242_), .A2(\a[23] ), .Z(new_n12243_));
  INV_X1     g11987(.I(new_n12243_), .ZN(new_n12244_));
  AOI22_X1   g11988(.A1(new_n2716_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n2719_), .ZN(new_n12245_));
  OAI21_X1   g11989(.A1(new_n4886_), .A2(new_n2924_), .B(new_n12245_), .ZN(new_n12246_));
  AOI21_X1   g11990(.A1(new_n5351_), .A2(new_n2722_), .B(new_n12246_), .ZN(new_n12247_));
  XOR2_X1    g11991(.A1(new_n12247_), .A2(new_n2714_), .Z(new_n12248_));
  INV_X1     g11992(.I(new_n12248_), .ZN(new_n12249_));
  OAI21_X1   g11993(.A1(new_n11883_), .A2(new_n12038_), .B(new_n12036_), .ZN(new_n12250_));
  OAI22_X1   g11994(.A1(new_n4666_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n4639_), .ZN(new_n12251_));
  AOI21_X1   g11995(.A1(\b[33] ), .A2(new_n3456_), .B(new_n12251_), .ZN(new_n12252_));
  OAI21_X1   g11996(.A1(new_n4676_), .A2(new_n3261_), .B(new_n12252_), .ZN(new_n12253_));
  XOR2_X1    g11997(.A1(new_n12253_), .A2(\a[29] ), .Z(new_n12254_));
  INV_X1     g11998(.I(new_n12254_), .ZN(new_n12255_));
  INV_X1     g11999(.I(new_n11893_), .ZN(new_n12256_));
  NAND2_X1   g12000(.A1(new_n11884_), .A2(new_n12256_), .ZN(new_n12257_));
  INV_X1     g12001(.I(new_n12257_), .ZN(new_n12258_));
  NAND3_X1   g12002(.A1(new_n11886_), .A2(new_n12017_), .A3(new_n12021_), .ZN(new_n12259_));
  OAI21_X1   g12003(.A1(new_n11709_), .A2(new_n11885_), .B(new_n12022_), .ZN(new_n12260_));
  NAND2_X1   g12004(.A1(new_n12259_), .A2(new_n12260_), .ZN(new_n12261_));
  OAI21_X1   g12005(.A1(new_n11884_), .A2(new_n12256_), .B(new_n12261_), .ZN(new_n12262_));
  INV_X1     g12006(.I(new_n12262_), .ZN(new_n12263_));
  AOI22_X1   g12007(.A1(new_n3864_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n3869_), .ZN(new_n12264_));
  OAI21_X1   g12008(.A1(new_n3624_), .A2(new_n5410_), .B(new_n12264_), .ZN(new_n12265_));
  AOI21_X1   g12009(.A1(new_n4030_), .A2(new_n3872_), .B(new_n12265_), .ZN(new_n12266_));
  XOR2_X1    g12010(.A1(new_n12266_), .A2(new_n3876_), .Z(new_n12267_));
  INV_X1     g12011(.I(new_n12267_), .ZN(new_n12268_));
  AOI22_X1   g12012(.A1(new_n4918_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n4921_), .ZN(new_n12269_));
  OAI21_X1   g12013(.A1(new_n3158_), .A2(new_n6099_), .B(new_n12269_), .ZN(new_n12270_));
  AOI21_X1   g12014(.A1(new_n4188_), .A2(new_n4699_), .B(new_n12270_), .ZN(new_n12271_));
  XOR2_X1    g12015(.A1(new_n12271_), .A2(new_n4446_), .Z(new_n12272_));
  INV_X1     g12016(.I(new_n12272_), .ZN(new_n12273_));
  AOI22_X1   g12017(.A1(new_n5155_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n5160_), .ZN(new_n12274_));
  OAI21_X1   g12018(.A1(new_n2495_), .A2(new_n6877_), .B(new_n12274_), .ZN(new_n12275_));
  AOI21_X1   g12019(.A1(new_n3407_), .A2(new_n5166_), .B(new_n12275_), .ZN(new_n12276_));
  XOR2_X1    g12020(.A1(new_n12276_), .A2(new_n5162_), .Z(new_n12277_));
  INV_X1     g12021(.I(new_n12277_), .ZN(new_n12278_));
  NAND2_X1   g12022(.A1(new_n12001_), .A2(new_n11998_), .ZN(new_n12279_));
  INV_X1     g12023(.I(new_n12279_), .ZN(new_n12280_));
  AOI22_X1   g12024(.A1(new_n6108_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n6111_), .ZN(new_n12281_));
  OAI21_X1   g12025(.A1(new_n2027_), .A2(new_n7708_), .B(new_n12281_), .ZN(new_n12282_));
  AOI21_X1   g12026(.A1(new_n2470_), .A2(new_n6105_), .B(new_n12282_), .ZN(new_n12283_));
  XOR2_X1    g12027(.A1(new_n12283_), .A2(new_n5849_), .Z(new_n12284_));
  NOR2_X1    g12028(.A1(new_n11985_), .A2(new_n11978_), .ZN(new_n12285_));
  NOR2_X1    g12029(.A1(new_n11975_), .A2(new_n11907_), .ZN(new_n12286_));
  OAI22_X1   g12030(.A1(new_n1296_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n1432_), .ZN(new_n12287_));
  AOI21_X1   g12031(.A1(\b[15] ), .A2(new_n7719_), .B(new_n12287_), .ZN(new_n12288_));
  OAI21_X1   g12032(.A1(new_n1444_), .A2(new_n8585_), .B(new_n12288_), .ZN(new_n12289_));
  XOR2_X1    g12033(.A1(new_n12289_), .A2(\a[47] ), .Z(new_n12290_));
  INV_X1     g12034(.I(new_n12290_), .ZN(new_n12291_));
  NOR2_X1    g12035(.A1(new_n11908_), .A2(new_n11966_), .ZN(new_n12292_));
  AOI22_X1   g12036(.A1(new_n8241_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n8246_), .ZN(new_n12293_));
  OAI21_X1   g12037(.A1(new_n941_), .A2(new_n9114_), .B(new_n12293_), .ZN(new_n12294_));
  AOI21_X1   g12038(.A1(new_n1449_), .A2(new_n8252_), .B(new_n12294_), .ZN(new_n12295_));
  XOR2_X1    g12039(.A1(new_n12295_), .A2(new_n8248_), .Z(new_n12296_));
  INV_X1     g12040(.I(new_n11953_), .ZN(new_n12297_));
  AOI22_X1   g12041(.A1(new_n11910_), .A2(new_n11642_), .B1(new_n11954_), .B2(new_n11951_), .ZN(new_n12298_));
  NOR2_X1    g12042(.A1(new_n12298_), .A2(new_n12297_), .ZN(new_n12299_));
  NAND2_X1   g12043(.A1(new_n11945_), .A2(new_n11912_), .ZN(new_n12300_));
  NAND2_X1   g12044(.A1(new_n12300_), .A2(new_n11944_), .ZN(new_n12301_));
  OAI21_X1   g12045(.A1(new_n11914_), .A2(new_n11935_), .B(new_n11936_), .ZN(new_n12302_));
  INV_X1     g12046(.I(new_n12302_), .ZN(new_n12303_));
  INV_X1     g12047(.I(new_n11306_), .ZN(new_n12304_));
  INV_X1     g12048(.I(new_n10979_), .ZN(new_n12305_));
  INV_X1     g12049(.I(new_n10981_), .ZN(new_n12306_));
  OAI22_X1   g12050(.A1(new_n12306_), .A2(new_n377_), .B1(new_n12305_), .B2(new_n339_), .ZN(new_n12307_));
  AOI21_X1   g12051(.A1(\b[3] ), .A2(new_n12304_), .B(new_n12307_), .ZN(new_n12308_));
  OAI21_X1   g12052(.A1(new_n566_), .A2(new_n10985_), .B(new_n12308_), .ZN(new_n12309_));
  XOR2_X1    g12053(.A1(new_n12309_), .A2(\a[59] ), .Z(new_n12310_));
  NAND3_X1   g12054(.A1(new_n11932_), .A2(\a[62] ), .A3(new_n11623_), .ZN(new_n12311_));
  INV_X1     g12055(.I(\a[62] ), .ZN(new_n12312_));
  AOI22_X1   g12056(.A1(new_n11926_), .A2(\b[2] ), .B1(new_n11924_), .B2(\b[1] ), .ZN(new_n12313_));
  NOR3_X1    g12057(.A1(new_n11617_), .A2(new_n11920_), .A3(\a[62] ), .ZN(new_n12314_));
  NAND3_X1   g12058(.A1(new_n11619_), .A2(new_n11920_), .A3(\a[62] ), .ZN(new_n12315_));
  INV_X1     g12059(.I(new_n12315_), .ZN(new_n12316_));
  NOR2_X1    g12060(.A1(new_n12316_), .A2(new_n12314_), .ZN(new_n12317_));
  OAI21_X1   g12061(.A1(new_n258_), .A2(new_n12317_), .B(new_n12313_), .ZN(new_n12318_));
  AOI21_X1   g12062(.A1(new_n554_), .A2(new_n11929_), .B(new_n12318_), .ZN(new_n12319_));
  XOR2_X1    g12063(.A1(new_n12319_), .A2(new_n12312_), .Z(new_n12320_));
  INV_X1     g12064(.I(new_n12320_), .ZN(new_n12321_));
  NOR2_X1    g12065(.A1(new_n12321_), .A2(new_n12311_), .ZN(new_n12322_));
  INV_X1     g12066(.I(new_n12311_), .ZN(new_n12323_));
  NOR2_X1    g12067(.A1(new_n12323_), .A2(new_n12320_), .ZN(new_n12324_));
  NOR2_X1    g12068(.A1(new_n12322_), .A2(new_n12324_), .ZN(new_n12325_));
  NOR2_X1    g12069(.A1(new_n12325_), .A2(new_n12310_), .ZN(new_n12326_));
  AND2_X2    g12070(.A1(new_n12325_), .A2(new_n12310_), .Z(new_n12327_));
  NOR2_X1    g12071(.A1(new_n12327_), .A2(new_n12326_), .ZN(new_n12328_));
  XOR2_X1    g12072(.A1(new_n12328_), .A2(new_n12303_), .Z(new_n12329_));
  AOI22_X1   g12073(.A1(new_n10064_), .A2(\b[8] ), .B1(\b[7] ), .B2(new_n10062_), .ZN(new_n12330_));
  OAI21_X1   g12074(.A1(new_n438_), .A2(new_n10399_), .B(new_n12330_), .ZN(new_n12331_));
  AOI21_X1   g12075(.A1(new_n799_), .A2(new_n10068_), .B(new_n12331_), .ZN(new_n12332_));
  XOR2_X1    g12076(.A1(new_n12332_), .A2(new_n10057_), .Z(new_n12333_));
  OR2_X2     g12077(.A1(new_n12329_), .A2(new_n12333_), .Z(new_n12334_));
  NAND2_X1   g12078(.A1(new_n12329_), .A2(new_n12333_), .ZN(new_n12335_));
  NAND2_X1   g12079(.A1(new_n12334_), .A2(new_n12335_), .ZN(new_n12336_));
  XOR2_X1    g12080(.A1(new_n12336_), .A2(new_n12301_), .Z(new_n12337_));
  OAI22_X1   g12081(.A1(new_n10390_), .A2(new_n852_), .B1(new_n776_), .B2(new_n10389_), .ZN(new_n12338_));
  AOI21_X1   g12082(.A1(\b[9] ), .A2(new_n9471_), .B(new_n12338_), .ZN(new_n12339_));
  OAI21_X1   g12083(.A1(new_n859_), .A2(new_n10388_), .B(new_n12339_), .ZN(new_n12340_));
  XOR2_X1    g12084(.A1(new_n12340_), .A2(\a[53] ), .Z(new_n12341_));
  NAND2_X1   g12085(.A1(new_n12337_), .A2(new_n12341_), .ZN(new_n12342_));
  INV_X1     g12086(.I(new_n12342_), .ZN(new_n12343_));
  NOR2_X1    g12087(.A1(new_n12337_), .A2(new_n12341_), .ZN(new_n12344_));
  NOR2_X1    g12088(.A1(new_n12343_), .A2(new_n12344_), .ZN(new_n12345_));
  NAND2_X1   g12089(.A1(new_n12345_), .A2(new_n12299_), .ZN(new_n12346_));
  XNOR2_X1   g12090(.A1(new_n12337_), .A2(new_n12341_), .ZN(new_n12347_));
  OAI21_X1   g12091(.A1(new_n12298_), .A2(new_n12297_), .B(new_n12347_), .ZN(new_n12348_));
  AOI21_X1   g12092(.A1(new_n12348_), .A2(new_n12346_), .B(new_n12296_), .ZN(new_n12349_));
  INV_X1     g12093(.I(new_n12296_), .ZN(new_n12350_));
  NOR3_X1    g12094(.A1(new_n12347_), .A2(new_n12297_), .A3(new_n12298_), .ZN(new_n12351_));
  NOR2_X1    g12095(.A1(new_n12345_), .A2(new_n12299_), .ZN(new_n12352_));
  NOR3_X1    g12096(.A1(new_n12351_), .A2(new_n12352_), .A3(new_n12350_), .ZN(new_n12353_));
  NOR4_X1    g12097(.A1(new_n12292_), .A2(new_n11965_), .A3(new_n12349_), .A4(new_n12353_), .ZN(new_n12354_));
  NOR2_X1    g12098(.A1(new_n12292_), .A2(new_n11965_), .ZN(new_n12355_));
  NOR2_X1    g12099(.A1(new_n12349_), .A2(new_n12353_), .ZN(new_n12356_));
  NOR2_X1    g12100(.A1(new_n12355_), .A2(new_n12356_), .ZN(new_n12357_));
  NOR2_X1    g12101(.A1(new_n12357_), .A2(new_n12354_), .ZN(new_n12358_));
  NOR2_X1    g12102(.A1(new_n12358_), .A2(new_n12291_), .ZN(new_n12359_));
  NOR3_X1    g12103(.A1(new_n12357_), .A2(new_n12354_), .A3(new_n12290_), .ZN(new_n12360_));
  NOR2_X1    g12104(.A1(new_n12359_), .A2(new_n12360_), .ZN(new_n12361_));
  OAI21_X1   g12105(.A1(new_n11974_), .A2(new_n12286_), .B(new_n12361_), .ZN(new_n12362_));
  NOR2_X1    g12106(.A1(new_n12286_), .A2(new_n11974_), .ZN(new_n12363_));
  INV_X1     g12107(.I(new_n12361_), .ZN(new_n12364_));
  NAND2_X1   g12108(.A1(new_n12364_), .A2(new_n12363_), .ZN(new_n12365_));
  AOI22_X1   g12109(.A1(new_n6569_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n6574_), .ZN(new_n12366_));
  OAI21_X1   g12110(.A1(new_n1553_), .A2(new_n8565_), .B(new_n12366_), .ZN(new_n12367_));
  AOI21_X1   g12111(.A1(new_n2452_), .A2(new_n6579_), .B(new_n12367_), .ZN(new_n12368_));
  XOR2_X1    g12112(.A1(new_n12368_), .A2(new_n6567_), .Z(new_n12369_));
  AOI21_X1   g12113(.A1(new_n12365_), .A2(new_n12362_), .B(new_n12369_), .ZN(new_n12370_));
  NOR2_X1    g12114(.A1(new_n12364_), .A2(new_n12363_), .ZN(new_n12371_));
  NOR3_X1    g12115(.A1(new_n12361_), .A2(new_n12286_), .A3(new_n11974_), .ZN(new_n12372_));
  INV_X1     g12116(.I(new_n12369_), .ZN(new_n12373_));
  NOR3_X1    g12117(.A1(new_n12371_), .A2(new_n12372_), .A3(new_n12373_), .ZN(new_n12374_));
  NOR2_X1    g12118(.A1(new_n12374_), .A2(new_n12370_), .ZN(new_n12375_));
  NOR3_X1    g12119(.A1(new_n12375_), .A2(new_n12285_), .A3(new_n11987_), .ZN(new_n12376_));
  NAND2_X1   g12120(.A1(new_n11989_), .A2(new_n11977_), .ZN(new_n12377_));
  OAI21_X1   g12121(.A1(new_n12371_), .A2(new_n12372_), .B(new_n12373_), .ZN(new_n12378_));
  NAND3_X1   g12122(.A1(new_n12365_), .A2(new_n12362_), .A3(new_n12369_), .ZN(new_n12379_));
  NAND2_X1   g12123(.A1(new_n12378_), .A2(new_n12379_), .ZN(new_n12380_));
  AOI21_X1   g12124(.A1(new_n12377_), .A2(new_n11990_), .B(new_n12380_), .ZN(new_n12381_));
  OAI21_X1   g12125(.A1(new_n12381_), .A2(new_n12376_), .B(new_n12284_), .ZN(new_n12382_));
  INV_X1     g12126(.I(new_n12284_), .ZN(new_n12383_));
  NAND3_X1   g12127(.A1(new_n12377_), .A2(new_n12380_), .A3(new_n11990_), .ZN(new_n12384_));
  OAI21_X1   g12128(.A1(new_n12285_), .A2(new_n11987_), .B(new_n12375_), .ZN(new_n12385_));
  NAND3_X1   g12129(.A1(new_n12385_), .A2(new_n12384_), .A3(new_n12383_), .ZN(new_n12386_));
  NAND2_X1   g12130(.A1(new_n12382_), .A2(new_n12386_), .ZN(new_n12387_));
  NOR3_X1    g12131(.A1(new_n12387_), .A2(new_n12280_), .A3(new_n11992_), .ZN(new_n12388_));
  AOI21_X1   g12132(.A1(new_n12385_), .A2(new_n12384_), .B(new_n12383_), .ZN(new_n12389_));
  NOR3_X1    g12133(.A1(new_n12381_), .A2(new_n12376_), .A3(new_n12284_), .ZN(new_n12390_));
  NOR2_X1    g12134(.A1(new_n12389_), .A2(new_n12390_), .ZN(new_n12391_));
  AOI21_X1   g12135(.A1(new_n12000_), .A2(new_n12279_), .B(new_n12391_), .ZN(new_n12392_));
  OAI21_X1   g12136(.A1(new_n12392_), .A2(new_n12388_), .B(new_n12278_), .ZN(new_n12393_));
  NAND3_X1   g12137(.A1(new_n12391_), .A2(new_n12000_), .A3(new_n12279_), .ZN(new_n12394_));
  OAI21_X1   g12138(.A1(new_n12280_), .A2(new_n11992_), .B(new_n12387_), .ZN(new_n12395_));
  NAND3_X1   g12139(.A1(new_n12395_), .A2(new_n12394_), .A3(new_n12277_), .ZN(new_n12396_));
  NAND2_X1   g12140(.A1(new_n12393_), .A2(new_n12396_), .ZN(new_n12397_));
  OAI21_X1   g12141(.A1(new_n12013_), .A2(new_n12012_), .B(new_n11902_), .ZN(new_n12398_));
  AOI21_X1   g12142(.A1(new_n12009_), .A2(new_n12398_), .B(new_n12397_), .ZN(new_n12399_));
  AOI21_X1   g12143(.A1(new_n12395_), .A2(new_n12394_), .B(new_n12277_), .ZN(new_n12400_));
  NOR3_X1    g12144(.A1(new_n12392_), .A2(new_n12278_), .A3(new_n12388_), .ZN(new_n12401_));
  NOR2_X1    g12145(.A1(new_n12401_), .A2(new_n12400_), .ZN(new_n12402_));
  OAI21_X1   g12146(.A1(new_n12015_), .A2(new_n12010_), .B(new_n12398_), .ZN(new_n12403_));
  NOR2_X1    g12147(.A1(new_n12402_), .A2(new_n12403_), .ZN(new_n12404_));
  OAI21_X1   g12148(.A1(new_n12399_), .A2(new_n12404_), .B(new_n12273_), .ZN(new_n12405_));
  NAND2_X1   g12149(.A1(new_n12402_), .A2(new_n12403_), .ZN(new_n12406_));
  NAND3_X1   g12150(.A1(new_n12009_), .A2(new_n12397_), .A3(new_n12398_), .ZN(new_n12407_));
  NAND3_X1   g12151(.A1(new_n12407_), .A2(new_n12406_), .A3(new_n12272_), .ZN(new_n12408_));
  NAND2_X1   g12152(.A1(new_n12405_), .A2(new_n12408_), .ZN(new_n12409_));
  AOI21_X1   g12153(.A1(new_n12259_), .A2(new_n12017_), .B(new_n12409_), .ZN(new_n12410_));
  INV_X1     g12154(.I(new_n12017_), .ZN(new_n12411_));
  NOR3_X1    g12155(.A1(new_n12022_), .A2(new_n11885_), .A3(new_n11709_), .ZN(new_n12412_));
  AOI21_X1   g12156(.A1(new_n12407_), .A2(new_n12406_), .B(new_n12272_), .ZN(new_n12413_));
  NOR3_X1    g12157(.A1(new_n12399_), .A2(new_n12404_), .A3(new_n12273_), .ZN(new_n12414_));
  NOR2_X1    g12158(.A1(new_n12414_), .A2(new_n12413_), .ZN(new_n12415_));
  NOR3_X1    g12159(.A1(new_n12415_), .A2(new_n12412_), .A3(new_n12411_), .ZN(new_n12416_));
  NOR3_X1    g12160(.A1(new_n12410_), .A2(new_n12416_), .A3(new_n12268_), .ZN(new_n12417_));
  OAI21_X1   g12161(.A1(new_n12411_), .A2(new_n12412_), .B(new_n12415_), .ZN(new_n12418_));
  NAND3_X1   g12162(.A1(new_n12259_), .A2(new_n12017_), .A3(new_n12409_), .ZN(new_n12419_));
  AOI21_X1   g12163(.A1(new_n12418_), .A2(new_n12419_), .B(new_n12267_), .ZN(new_n12420_));
  NOR2_X1    g12164(.A1(new_n12420_), .A2(new_n12417_), .ZN(new_n12421_));
  NOR3_X1    g12165(.A1(new_n12421_), .A2(new_n12263_), .A3(new_n12258_), .ZN(new_n12422_));
  NAND3_X1   g12166(.A1(new_n12418_), .A2(new_n12419_), .A3(new_n12267_), .ZN(new_n12423_));
  OAI21_X1   g12167(.A1(new_n12410_), .A2(new_n12416_), .B(new_n12268_), .ZN(new_n12424_));
  NAND2_X1   g12168(.A1(new_n12423_), .A2(new_n12424_), .ZN(new_n12425_));
  AOI21_X1   g12169(.A1(new_n12257_), .A2(new_n12262_), .B(new_n12425_), .ZN(new_n12426_));
  NOR3_X1    g12170(.A1(new_n12426_), .A2(new_n12422_), .A3(new_n12255_), .ZN(new_n12427_));
  NAND3_X1   g12171(.A1(new_n12425_), .A2(new_n12257_), .A3(new_n12262_), .ZN(new_n12428_));
  OAI21_X1   g12172(.A1(new_n12263_), .A2(new_n12258_), .B(new_n12421_), .ZN(new_n12429_));
  AOI21_X1   g12173(.A1(new_n12429_), .A2(new_n12428_), .B(new_n12254_), .ZN(new_n12430_));
  NOR2_X1    g12174(.A1(new_n12427_), .A2(new_n12430_), .ZN(new_n12431_));
  NAND2_X1   g12175(.A1(new_n12431_), .A2(new_n12250_), .ZN(new_n12432_));
  AOI21_X1   g12176(.A1(new_n11882_), .A2(new_n12033_), .B(new_n12039_), .ZN(new_n12433_));
  NAND3_X1   g12177(.A1(new_n12429_), .A2(new_n12254_), .A3(new_n12428_), .ZN(new_n12434_));
  OAI21_X1   g12178(.A1(new_n12426_), .A2(new_n12422_), .B(new_n12255_), .ZN(new_n12435_));
  NAND2_X1   g12179(.A1(new_n12435_), .A2(new_n12434_), .ZN(new_n12436_));
  NAND2_X1   g12180(.A1(new_n12436_), .A2(new_n12433_), .ZN(new_n12437_));
  NAND3_X1   g12181(.A1(new_n12437_), .A2(new_n12432_), .A3(new_n12249_), .ZN(new_n12438_));
  NOR2_X1    g12182(.A1(new_n12436_), .A2(new_n12433_), .ZN(new_n12439_));
  NOR2_X1    g12183(.A1(new_n12431_), .A2(new_n12250_), .ZN(new_n12440_));
  OAI21_X1   g12184(.A1(new_n12439_), .A2(new_n12440_), .B(new_n12248_), .ZN(new_n12441_));
  NAND2_X1   g12185(.A1(new_n12441_), .A2(new_n12438_), .ZN(new_n12442_));
  INV_X1     g12186(.I(new_n12049_), .ZN(new_n12443_));
  AOI21_X1   g12187(.A1(new_n12052_), .A2(new_n12046_), .B(new_n12443_), .ZN(new_n12444_));
  NOR2_X1    g12188(.A1(new_n12444_), .A2(new_n12442_), .ZN(new_n12445_));
  NOR3_X1    g12189(.A1(new_n12439_), .A2(new_n12440_), .A3(new_n12248_), .ZN(new_n12446_));
  AOI21_X1   g12190(.A1(new_n12437_), .A2(new_n12432_), .B(new_n12249_), .ZN(new_n12447_));
  NOR2_X1    g12191(.A1(new_n12447_), .A2(new_n12446_), .ZN(new_n12448_));
  OAI21_X1   g12192(.A1(new_n12050_), .A2(new_n12059_), .B(new_n12049_), .ZN(new_n12449_));
  NOR2_X1    g12193(.A1(new_n12448_), .A2(new_n12449_), .ZN(new_n12450_));
  NOR3_X1    g12194(.A1(new_n12445_), .A2(new_n12450_), .A3(new_n12244_), .ZN(new_n12451_));
  NAND2_X1   g12195(.A1(new_n12448_), .A2(new_n12449_), .ZN(new_n12452_));
  NAND2_X1   g12196(.A1(new_n12444_), .A2(new_n12442_), .ZN(new_n12453_));
  AOI21_X1   g12197(.A1(new_n12453_), .A2(new_n12452_), .B(new_n12243_), .ZN(new_n12454_));
  NOR2_X1    g12198(.A1(new_n12451_), .A2(new_n12454_), .ZN(new_n12455_));
  AOI21_X1   g12199(.A1(new_n12237_), .A2(new_n12239_), .B(new_n12455_), .ZN(new_n12456_));
  NAND2_X1   g12200(.A1(new_n12239_), .A2(new_n12237_), .ZN(new_n12457_));
  NAND3_X1   g12201(.A1(new_n12453_), .A2(new_n12452_), .A3(new_n12243_), .ZN(new_n12458_));
  OAI21_X1   g12202(.A1(new_n12445_), .A2(new_n12450_), .B(new_n12244_), .ZN(new_n12459_));
  NAND2_X1   g12203(.A1(new_n12459_), .A2(new_n12458_), .ZN(new_n12460_));
  NOR2_X1    g12204(.A1(new_n12457_), .A2(new_n12460_), .ZN(new_n12461_));
  AOI22_X1   g12205(.A1(new_n1738_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n1743_), .ZN(new_n12462_));
  OAI21_X1   g12206(.A1(new_n6490_), .A2(new_n1931_), .B(new_n12462_), .ZN(new_n12463_));
  AOI21_X1   g12207(.A1(new_n7906_), .A2(new_n1746_), .B(new_n12463_), .ZN(new_n12464_));
  XOR2_X1    g12208(.A1(new_n12464_), .A2(new_n1736_), .Z(new_n12465_));
  INV_X1     g12209(.I(new_n12465_), .ZN(new_n12466_));
  OAI21_X1   g12210(.A1(new_n12456_), .A2(new_n12461_), .B(new_n12466_), .ZN(new_n12467_));
  NAND2_X1   g12211(.A1(new_n12457_), .A2(new_n12460_), .ZN(new_n12468_));
  NAND3_X1   g12212(.A1(new_n12455_), .A2(new_n12239_), .A3(new_n12237_), .ZN(new_n12469_));
  NAND3_X1   g12213(.A1(new_n12468_), .A2(new_n12469_), .A3(new_n12465_), .ZN(new_n12470_));
  NAND2_X1   g12214(.A1(new_n12467_), .A2(new_n12470_), .ZN(new_n12471_));
  NAND3_X1   g12215(.A1(new_n12236_), .A2(new_n12471_), .A3(new_n12075_), .ZN(new_n12472_));
  INV_X1     g12216(.I(new_n12472_), .ZN(new_n12473_));
  AOI21_X1   g12217(.A1(new_n12236_), .A2(new_n12075_), .B(new_n12471_), .ZN(new_n12474_));
  OAI21_X1   g12218(.A1(new_n12473_), .A2(new_n12474_), .B(new_n12235_), .ZN(new_n12475_));
  INV_X1     g12219(.I(new_n12235_), .ZN(new_n12476_));
  NAND2_X1   g12220(.A1(new_n12236_), .A2(new_n12075_), .ZN(new_n12477_));
  INV_X1     g12221(.I(new_n12471_), .ZN(new_n12478_));
  NAND2_X1   g12222(.A1(new_n12477_), .A2(new_n12478_), .ZN(new_n12479_));
  NAND3_X1   g12223(.A1(new_n12479_), .A2(new_n12472_), .A3(new_n12476_), .ZN(new_n12480_));
  NAND3_X1   g12224(.A1(new_n12231_), .A2(new_n12475_), .A3(new_n12480_), .ZN(new_n12481_));
  INV_X1     g12225(.I(new_n12481_), .ZN(new_n12482_));
  AOI21_X1   g12226(.A1(new_n12475_), .A2(new_n12480_), .B(new_n12231_), .ZN(new_n12483_));
  OAI21_X1   g12227(.A1(new_n12482_), .A2(new_n12483_), .B(new_n12230_), .ZN(new_n12484_));
  INV_X1     g12228(.I(new_n12231_), .ZN(new_n12485_));
  NAND2_X1   g12229(.A1(new_n12475_), .A2(new_n12480_), .ZN(new_n12486_));
  NAND2_X1   g12230(.A1(new_n12486_), .A2(new_n12485_), .ZN(new_n12487_));
  NAND3_X1   g12231(.A1(new_n12487_), .A2(new_n12229_), .A3(new_n12481_), .ZN(new_n12488_));
  NAND2_X1   g12232(.A1(new_n12484_), .A2(new_n12488_), .ZN(new_n12489_));
  NOR3_X1    g12233(.A1(new_n12489_), .A2(new_n12225_), .A3(new_n12106_), .ZN(new_n12490_));
  NAND2_X1   g12234(.A1(new_n12115_), .A2(new_n11875_), .ZN(new_n12491_));
  AOI21_X1   g12235(.A1(new_n12487_), .A2(new_n12481_), .B(new_n12229_), .ZN(new_n12492_));
  NOR3_X1    g12236(.A1(new_n12482_), .A2(new_n12483_), .A3(new_n12230_), .ZN(new_n12493_));
  NOR2_X1    g12237(.A1(new_n12492_), .A2(new_n12493_), .ZN(new_n12494_));
  AOI21_X1   g12238(.A1(new_n12114_), .A2(new_n12491_), .B(new_n12494_), .ZN(new_n12495_));
  NOR3_X1    g12239(.A1(new_n12495_), .A2(new_n12490_), .A3(new_n12224_), .ZN(new_n12496_));
  NAND3_X1   g12240(.A1(new_n12494_), .A2(new_n12491_), .A3(new_n12114_), .ZN(new_n12497_));
  OAI21_X1   g12241(.A1(new_n12225_), .A2(new_n12106_), .B(new_n12489_), .ZN(new_n12498_));
  AOI21_X1   g12242(.A1(new_n12498_), .A2(new_n12497_), .B(new_n12223_), .ZN(new_n12499_));
  NOR2_X1    g12243(.A1(new_n12496_), .A2(new_n12499_), .ZN(new_n12500_));
  NAND2_X1   g12244(.A1(new_n12219_), .A2(new_n12500_), .ZN(new_n12501_));
  NAND3_X1   g12245(.A1(new_n12498_), .A2(new_n12497_), .A3(new_n12223_), .ZN(new_n12502_));
  OAI21_X1   g12246(.A1(new_n12495_), .A2(new_n12490_), .B(new_n12224_), .ZN(new_n12503_));
  NAND2_X1   g12247(.A1(new_n12503_), .A2(new_n12502_), .ZN(new_n12504_));
  NAND2_X1   g12248(.A1(new_n12504_), .A2(new_n12218_), .ZN(new_n12505_));
  NAND3_X1   g12249(.A1(new_n12217_), .A2(new_n12501_), .A3(new_n12505_), .ZN(new_n12506_));
  NOR2_X1    g12250(.A1(new_n12504_), .A2(new_n12218_), .ZN(new_n12507_));
  INV_X1     g12251(.I(new_n12505_), .ZN(new_n12508_));
  OAI21_X1   g12252(.A1(new_n12508_), .A2(new_n12507_), .B(new_n12216_), .ZN(new_n12509_));
  AOI22_X1   g12253(.A1(new_n267_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n261_), .ZN(new_n12510_));
  OAI21_X1   g12254(.A1(new_n12147_), .A2(new_n284_), .B(new_n12510_), .ZN(new_n12511_));
  INV_X1     g12255(.I(new_n12511_), .ZN(new_n12512_));
  AOI21_X1   g12256(.A1(new_n12155_), .A2(\b[60] ), .B(\b[59] ), .ZN(new_n12513_));
  INV_X1     g12257(.I(new_n12513_), .ZN(new_n12514_));
  AOI21_X1   g12258(.A1(new_n11835_), .A2(\b[61] ), .B(\b[60] ), .ZN(new_n12515_));
  INV_X1     g12259(.I(new_n12515_), .ZN(new_n12516_));
  XNOR2_X1   g12260(.A1(\b[61] ), .A2(\b[62] ), .ZN(new_n12517_));
  AOI21_X1   g12261(.A1(new_n12514_), .A2(new_n12516_), .B(new_n12517_), .ZN(new_n12518_));
  NAND3_X1   g12262(.A1(new_n12514_), .A2(new_n12516_), .A3(new_n12517_), .ZN(new_n12519_));
  INV_X1     g12263(.I(new_n12519_), .ZN(new_n12520_));
  OAI21_X1   g12264(.A1(new_n12520_), .A2(new_n12518_), .B(new_n265_), .ZN(new_n12521_));
  AOI21_X1   g12265(.A1(new_n12521_), .A2(new_n12512_), .B(new_n270_), .ZN(new_n12522_));
  INV_X1     g12266(.I(new_n12518_), .ZN(new_n12523_));
  AOI21_X1   g12267(.A1(new_n12523_), .A2(new_n12519_), .B(new_n279_), .ZN(new_n12524_));
  NOR3_X1    g12268(.A1(new_n12524_), .A2(\a[2] ), .A3(new_n12511_), .ZN(new_n12525_));
  NOR2_X1    g12269(.A1(new_n12525_), .A2(new_n12522_), .ZN(new_n12526_));
  AOI21_X1   g12270(.A1(new_n12509_), .A2(new_n12506_), .B(new_n12526_), .ZN(new_n12527_));
  INV_X1     g12271(.I(new_n12527_), .ZN(new_n12528_));
  NAND3_X1   g12272(.A1(new_n12509_), .A2(new_n12506_), .A3(new_n12526_), .ZN(new_n12529_));
  NAND3_X1   g12273(.A1(new_n12528_), .A2(new_n12202_), .A3(new_n12529_), .ZN(new_n12530_));
  INV_X1     g12274(.I(new_n12202_), .ZN(new_n12531_));
  NOR3_X1    g12275(.A1(new_n12508_), .A2(new_n12216_), .A3(new_n12507_), .ZN(new_n12532_));
  AOI21_X1   g12276(.A1(new_n12505_), .A2(new_n12501_), .B(new_n12217_), .ZN(new_n12533_));
  NOR4_X1    g12277(.A1(new_n12533_), .A2(new_n12532_), .A3(new_n12522_), .A4(new_n12525_), .ZN(new_n12534_));
  OAI21_X1   g12278(.A1(new_n12527_), .A2(new_n12534_), .B(new_n12531_), .ZN(new_n12535_));
  NAND2_X1   g12279(.A1(new_n12535_), .A2(new_n12530_), .ZN(new_n12536_));
  NAND2_X1   g12280(.A1(new_n12198_), .A2(new_n12536_), .ZN(new_n12537_));
  NAND3_X1   g12281(.A1(new_n12197_), .A2(new_n12530_), .A3(new_n12535_), .ZN(new_n12538_));
  NAND2_X1   g12282(.A1(new_n12537_), .A2(new_n12538_), .ZN(new_n12539_));
  XOR2_X1    g12283(.A1(new_n12539_), .A2(new_n12196_), .Z(\f[62] ));
  INV_X1     g12284(.I(new_n12213_), .ZN(new_n12541_));
  NAND2_X1   g12285(.A1(new_n12501_), .A2(new_n12505_), .ZN(new_n12542_));
  AOI21_X1   g12286(.A1(new_n12542_), .A2(new_n12215_), .B(new_n12541_), .ZN(new_n12543_));
  INV_X1     g12287(.I(new_n12543_), .ZN(new_n12544_));
  AOI22_X1   g12288(.A1(new_n518_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n636_), .ZN(new_n12545_));
  OAI21_X1   g12289(.A1(new_n9972_), .A2(new_n917_), .B(new_n12545_), .ZN(new_n12546_));
  AOI21_X1   g12290(.A1(new_n10631_), .A2(new_n618_), .B(new_n12546_), .ZN(new_n12547_));
  XOR2_X1    g12291(.A1(new_n12547_), .A2(new_n488_), .Z(new_n12548_));
  OAI22_X1   g12292(.A1(new_n713_), .A2(new_n9942_), .B1(new_n9376_), .B2(new_n717_), .ZN(new_n12549_));
  AOI21_X1   g12293(.A1(\b[52] ), .A2(new_n1126_), .B(new_n12549_), .ZN(new_n12550_));
  OAI21_X1   g12294(.A1(new_n9952_), .A2(new_n986_), .B(new_n12550_), .ZN(new_n12551_));
  XOR2_X1    g12295(.A1(new_n12551_), .A2(\a[11] ), .Z(new_n12552_));
  INV_X1     g12296(.I(new_n12552_), .ZN(new_n12553_));
  NAND2_X1   g12297(.A1(new_n12477_), .A2(new_n12470_), .ZN(new_n12554_));
  NAND2_X1   g12298(.A1(new_n12554_), .A2(new_n12467_), .ZN(new_n12555_));
  INV_X1     g12299(.I(new_n12555_), .ZN(new_n12556_));
  AOI22_X1   g12300(.A1(new_n1738_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n1743_), .ZN(new_n12557_));
  OAI21_X1   g12301(.A1(new_n6775_), .A2(new_n1931_), .B(new_n12557_), .ZN(new_n12558_));
  AOI21_X1   g12302(.A1(new_n7926_), .A2(new_n1746_), .B(new_n12558_), .ZN(new_n12559_));
  XOR2_X1    g12303(.A1(new_n12559_), .A2(new_n1736_), .Z(new_n12560_));
  AOI22_X1   g12304(.A1(new_n3864_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n3869_), .ZN(new_n12561_));
  OAI21_X1   g12305(.A1(new_n4022_), .A2(new_n5410_), .B(new_n12561_), .ZN(new_n12562_));
  AOI21_X1   g12306(.A1(new_n4223_), .A2(new_n3872_), .B(new_n12562_), .ZN(new_n12563_));
  XOR2_X1    g12307(.A1(new_n12563_), .A2(new_n3876_), .Z(new_n12564_));
  OAI21_X1   g12308(.A1(new_n12285_), .A2(new_n11987_), .B(new_n12379_), .ZN(new_n12565_));
  NAND2_X1   g12309(.A1(new_n12565_), .A2(new_n12378_), .ZN(new_n12566_));
  AOI22_X1   g12310(.A1(new_n6569_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n6574_), .ZN(new_n12567_));
  OAI21_X1   g12311(.A1(new_n1859_), .A2(new_n8565_), .B(new_n12567_), .ZN(new_n12568_));
  AOI21_X1   g12312(.A1(new_n2032_), .A2(new_n6579_), .B(new_n12568_), .ZN(new_n12569_));
  XOR2_X1    g12313(.A1(new_n12569_), .A2(new_n6567_), .Z(new_n12570_));
  INV_X1     g12314(.I(new_n12570_), .ZN(new_n12571_));
  INV_X1     g12315(.I(new_n12334_), .ZN(new_n12572_));
  AOI21_X1   g12316(.A1(new_n12301_), .A2(new_n12335_), .B(new_n12572_), .ZN(new_n12573_));
  INV_X1     g12317(.I(new_n12573_), .ZN(new_n12574_));
  NOR2_X1    g12318(.A1(new_n12303_), .A2(new_n12327_), .ZN(new_n12575_));
  NOR2_X1    g12319(.A1(new_n12575_), .A2(new_n12326_), .ZN(new_n12576_));
  AOI22_X1   g12320(.A1(new_n11926_), .A2(\b[3] ), .B1(new_n11924_), .B2(\b[2] ), .ZN(new_n12577_));
  OAI21_X1   g12321(.A1(new_n275_), .A2(new_n12317_), .B(new_n12577_), .ZN(new_n12578_));
  AOI21_X1   g12322(.A1(new_n299_), .A2(new_n11929_), .B(new_n12578_), .ZN(new_n12579_));
  XOR2_X1    g12323(.A1(new_n12579_), .A2(new_n12312_), .Z(new_n12580_));
  INV_X1     g12324(.I(\a[63] ), .ZN(new_n12581_));
  NOR2_X1    g12325(.A1(new_n12581_), .A2(\a[62] ), .ZN(new_n12582_));
  NOR2_X1    g12326(.A1(new_n12312_), .A2(\a[63] ), .ZN(new_n12583_));
  NOR2_X1    g12327(.A1(new_n12582_), .A2(new_n12583_), .ZN(new_n12584_));
  NOR2_X1    g12328(.A1(new_n12584_), .A2(new_n258_), .ZN(new_n12585_));
  AND2_X2    g12329(.A1(new_n12580_), .A2(new_n12585_), .Z(new_n12586_));
  NOR2_X1    g12330(.A1(new_n12580_), .A2(new_n12585_), .ZN(new_n12587_));
  NOR2_X1    g12331(.A1(new_n12586_), .A2(new_n12587_), .ZN(new_n12588_));
  XOR2_X1    g12332(.A1(new_n12588_), .A2(new_n12322_), .Z(new_n12589_));
  INV_X1     g12333(.I(new_n12589_), .ZN(new_n12590_));
  AOI22_X1   g12334(.A1(new_n10981_), .A2(\b[6] ), .B1(new_n10979_), .B2(\b[5] ), .ZN(new_n12591_));
  OAI21_X1   g12335(.A1(new_n339_), .A2(new_n11306_), .B(new_n12591_), .ZN(new_n12592_));
  AOI21_X1   g12336(.A1(new_n916_), .A2(new_n10984_), .B(new_n12592_), .ZN(new_n12593_));
  XOR2_X1    g12337(.A1(new_n12593_), .A2(new_n10989_), .Z(new_n12594_));
  INV_X1     g12338(.I(new_n12594_), .ZN(new_n12595_));
  NAND2_X1   g12339(.A1(new_n12590_), .A2(new_n12595_), .ZN(new_n12596_));
  NOR2_X1    g12340(.A1(new_n12590_), .A2(new_n12595_), .ZN(new_n12597_));
  INV_X1     g12341(.I(new_n12597_), .ZN(new_n12598_));
  NAND2_X1   g12342(.A1(new_n12598_), .A2(new_n12596_), .ZN(new_n12599_));
  XOR2_X1    g12343(.A1(new_n12599_), .A2(new_n12576_), .Z(new_n12600_));
  AOI22_X1   g12344(.A1(new_n10064_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n10062_), .ZN(new_n12601_));
  OAI21_X1   g12345(.A1(new_n471_), .A2(new_n10399_), .B(new_n12601_), .ZN(new_n12602_));
  AOI21_X1   g12346(.A1(new_n676_), .A2(new_n10068_), .B(new_n12602_), .ZN(new_n12603_));
  XOR2_X1    g12347(.A1(new_n12603_), .A2(new_n10057_), .Z(new_n12604_));
  INV_X1     g12348(.I(new_n12604_), .ZN(new_n12605_));
  NAND2_X1   g12349(.A1(new_n12600_), .A2(new_n12605_), .ZN(new_n12606_));
  OR2_X2     g12350(.A1(new_n12600_), .A2(new_n12605_), .Z(new_n12607_));
  NAND2_X1   g12351(.A1(new_n12607_), .A2(new_n12606_), .ZN(new_n12608_));
  XOR2_X1    g12352(.A1(new_n12608_), .A2(new_n12574_), .Z(new_n12609_));
  AOI22_X1   g12353(.A1(new_n9125_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n9123_), .ZN(new_n12610_));
  OAI21_X1   g12354(.A1(new_n776_), .A2(new_n9470_), .B(new_n12610_), .ZN(new_n12611_));
  AOI21_X1   g12355(.A1(new_n1194_), .A2(new_n9129_), .B(new_n12611_), .ZN(new_n12612_));
  XOR2_X1    g12356(.A1(new_n12612_), .A2(new_n9133_), .Z(new_n12613_));
  NAND2_X1   g12357(.A1(new_n12346_), .A2(new_n12342_), .ZN(new_n12614_));
  NAND2_X1   g12358(.A1(new_n12614_), .A2(new_n12613_), .ZN(new_n12615_));
  NOR2_X1    g12359(.A1(new_n12614_), .A2(new_n12613_), .ZN(new_n12616_));
  INV_X1     g12360(.I(new_n12616_), .ZN(new_n12617_));
  NAND2_X1   g12361(.A1(new_n12617_), .A2(new_n12615_), .ZN(new_n12618_));
  XOR2_X1    g12362(.A1(new_n12618_), .A2(new_n12609_), .Z(new_n12619_));
  INV_X1     g12363(.I(new_n12619_), .ZN(new_n12620_));
  OAI22_X1   g12364(.A1(new_n9461_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n9462_), .ZN(new_n12621_));
  AOI21_X1   g12365(.A1(\b[13] ), .A2(new_n8575_), .B(new_n12621_), .ZN(new_n12622_));
  OAI21_X1   g12366(.A1(new_n1275_), .A2(new_n9460_), .B(new_n12622_), .ZN(new_n12623_));
  XOR2_X1    g12367(.A1(new_n12623_), .A2(\a[50] ), .Z(new_n12624_));
  OR2_X2     g12368(.A1(new_n12354_), .A2(new_n12353_), .Z(new_n12625_));
  NAND2_X1   g12369(.A1(new_n12625_), .A2(new_n12624_), .ZN(new_n12626_));
  OR2_X2     g12370(.A1(new_n12625_), .A2(new_n12624_), .Z(new_n12627_));
  AND3_X2    g12371(.A1(new_n12627_), .A2(new_n12620_), .A3(new_n12626_), .Z(new_n12628_));
  AOI21_X1   g12372(.A1(new_n12627_), .A2(new_n12626_), .B(new_n12620_), .ZN(new_n12629_));
  NOR2_X1    g12373(.A1(new_n12628_), .A2(new_n12629_), .ZN(new_n12630_));
  AOI22_X1   g12374(.A1(new_n7403_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n7408_), .ZN(new_n12631_));
  OAI21_X1   g12375(.A1(new_n1296_), .A2(new_n9488_), .B(new_n12631_), .ZN(new_n12632_));
  AOI21_X1   g12376(.A1(new_n2038_), .A2(new_n7414_), .B(new_n12632_), .ZN(new_n12633_));
  XOR2_X1    g12377(.A1(new_n12633_), .A2(new_n7410_), .Z(new_n12634_));
  INV_X1     g12378(.I(new_n12634_), .ZN(new_n12635_));
  NAND2_X1   g12379(.A1(new_n12358_), .A2(new_n12290_), .ZN(new_n12636_));
  AOI21_X1   g12380(.A1(new_n12365_), .A2(new_n12636_), .B(new_n12635_), .ZN(new_n12637_));
  INV_X1     g12381(.I(new_n12637_), .ZN(new_n12638_));
  NAND3_X1   g12382(.A1(new_n12365_), .A2(new_n12636_), .A3(new_n12635_), .ZN(new_n12639_));
  NAND3_X1   g12383(.A1(new_n12638_), .A2(new_n12630_), .A3(new_n12639_), .ZN(new_n12640_));
  INV_X1     g12384(.I(new_n12630_), .ZN(new_n12641_));
  INV_X1     g12385(.I(new_n12639_), .ZN(new_n12642_));
  OAI21_X1   g12386(.A1(new_n12642_), .A2(new_n12637_), .B(new_n12641_), .ZN(new_n12643_));
  NAND2_X1   g12387(.A1(new_n12643_), .A2(new_n12640_), .ZN(new_n12644_));
  NAND2_X1   g12388(.A1(new_n12644_), .A2(new_n12571_), .ZN(new_n12645_));
  NAND3_X1   g12389(.A1(new_n12643_), .A2(new_n12640_), .A3(new_n12570_), .ZN(new_n12646_));
  NAND2_X1   g12390(.A1(new_n12645_), .A2(new_n12646_), .ZN(new_n12647_));
  XOR2_X1    g12391(.A1(new_n12647_), .A2(new_n12566_), .Z(new_n12648_));
  AOI22_X1   g12392(.A1(new_n6108_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n6111_), .ZN(new_n12649_));
  OAI21_X1   g12393(.A1(new_n2142_), .A2(new_n7708_), .B(new_n12649_), .ZN(new_n12650_));
  AOI21_X1   g12394(.A1(new_n3033_), .A2(new_n6105_), .B(new_n12650_), .ZN(new_n12651_));
  XOR2_X1    g12395(.A1(new_n12651_), .A2(new_n5849_), .Z(new_n12652_));
  INV_X1     g12396(.I(new_n12652_), .ZN(new_n12653_));
  AOI21_X1   g12397(.A1(new_n12394_), .A2(new_n12382_), .B(new_n12653_), .ZN(new_n12654_));
  NAND3_X1   g12398(.A1(new_n12394_), .A2(new_n12382_), .A3(new_n12653_), .ZN(new_n12655_));
  INV_X1     g12399(.I(new_n12655_), .ZN(new_n12656_));
  NOR3_X1    g12400(.A1(new_n12656_), .A2(new_n12648_), .A3(new_n12654_), .ZN(new_n12657_));
  XNOR2_X1   g12401(.A1(new_n12647_), .A2(new_n12566_), .ZN(new_n12658_));
  INV_X1     g12402(.I(new_n12654_), .ZN(new_n12659_));
  AOI21_X1   g12403(.A1(new_n12659_), .A2(new_n12655_), .B(new_n12658_), .ZN(new_n12660_));
  NOR2_X1    g12404(.A1(new_n12660_), .A2(new_n12657_), .ZN(new_n12661_));
  INV_X1     g12405(.I(new_n12661_), .ZN(new_n12662_));
  OAI22_X1   g12406(.A1(new_n3158_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n3006_), .ZN(new_n12663_));
  AOI21_X1   g12407(.A1(\b[25] ), .A2(new_n5420_), .B(new_n12663_), .ZN(new_n12664_));
  OAI21_X1   g12408(.A1(new_n3165_), .A2(new_n6124_), .B(new_n12664_), .ZN(new_n12665_));
  XOR2_X1    g12409(.A1(new_n12665_), .A2(\a[38] ), .Z(new_n12666_));
  INV_X1     g12410(.I(new_n12666_), .ZN(new_n12667_));
  NOR2_X1    g12411(.A1(new_n12399_), .A2(new_n12401_), .ZN(new_n12668_));
  NOR2_X1    g12412(.A1(new_n12668_), .A2(new_n12667_), .ZN(new_n12669_));
  NAND2_X1   g12413(.A1(new_n12406_), .A2(new_n12396_), .ZN(new_n12670_));
  NOR2_X1    g12414(.A1(new_n12670_), .A2(new_n12666_), .ZN(new_n12671_));
  NOR3_X1    g12415(.A1(new_n12669_), .A2(new_n12662_), .A3(new_n12671_), .ZN(new_n12672_));
  NOR2_X1    g12416(.A1(new_n12669_), .A2(new_n12671_), .ZN(new_n12673_));
  NOR2_X1    g12417(.A1(new_n12673_), .A2(new_n12661_), .ZN(new_n12674_));
  NOR2_X1    g12418(.A1(new_n12674_), .A2(new_n12672_), .ZN(new_n12675_));
  AOI22_X1   g12419(.A1(new_n4918_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n4921_), .ZN(new_n12676_));
  OAI21_X1   g12420(.A1(new_n3185_), .A2(new_n6099_), .B(new_n12676_), .ZN(new_n12677_));
  AOI21_X1   g12421(.A1(new_n4230_), .A2(new_n4699_), .B(new_n12677_), .ZN(new_n12678_));
  XOR2_X1    g12422(.A1(new_n12678_), .A2(new_n4446_), .Z(new_n12679_));
  NAND2_X1   g12423(.A1(new_n12418_), .A2(new_n12408_), .ZN(new_n12680_));
  NAND2_X1   g12424(.A1(new_n12680_), .A2(new_n12679_), .ZN(new_n12681_));
  INV_X1     g12425(.I(new_n12679_), .ZN(new_n12682_));
  NAND3_X1   g12426(.A1(new_n12418_), .A2(new_n12408_), .A3(new_n12682_), .ZN(new_n12683_));
  NAND3_X1   g12427(.A1(new_n12681_), .A2(new_n12675_), .A3(new_n12683_), .ZN(new_n12684_));
  INV_X1     g12428(.I(new_n12675_), .ZN(new_n12685_));
  NAND2_X1   g12429(.A1(new_n12681_), .A2(new_n12683_), .ZN(new_n12686_));
  NAND2_X1   g12430(.A1(new_n12686_), .A2(new_n12685_), .ZN(new_n12687_));
  NAND2_X1   g12431(.A1(new_n12687_), .A2(new_n12684_), .ZN(new_n12688_));
  NOR2_X1    g12432(.A1(new_n12688_), .A2(new_n12564_), .ZN(new_n12689_));
  INV_X1     g12433(.I(new_n12564_), .ZN(new_n12690_));
  AOI21_X1   g12434(.A1(new_n12687_), .A2(new_n12684_), .B(new_n12690_), .ZN(new_n12691_));
  NOR2_X1    g12435(.A1(new_n12689_), .A2(new_n12691_), .ZN(new_n12692_));
  NAND3_X1   g12436(.A1(new_n12421_), .A2(new_n12257_), .A3(new_n12262_), .ZN(new_n12693_));
  NAND2_X1   g12437(.A1(new_n12693_), .A2(new_n12423_), .ZN(new_n12694_));
  XNOR2_X1   g12438(.A1(new_n12692_), .A2(new_n12694_), .ZN(new_n12695_));
  AOI22_X1   g12439(.A1(new_n3267_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n3270_), .ZN(new_n12696_));
  OAI21_X1   g12440(.A1(new_n4639_), .A2(new_n3475_), .B(new_n12696_), .ZN(new_n12697_));
  AOI21_X1   g12441(.A1(new_n5594_), .A2(new_n3273_), .B(new_n12697_), .ZN(new_n12698_));
  XOR2_X1    g12442(.A1(new_n12698_), .A2(new_n3264_), .Z(new_n12699_));
  NAND2_X1   g12443(.A1(new_n12436_), .A2(new_n12250_), .ZN(new_n12700_));
  OAI21_X1   g12444(.A1(new_n12426_), .A2(new_n12422_), .B(new_n12254_), .ZN(new_n12701_));
  NAND2_X1   g12445(.A1(new_n12700_), .A2(new_n12701_), .ZN(new_n12702_));
  NAND2_X1   g12446(.A1(new_n12702_), .A2(new_n12699_), .ZN(new_n12703_));
  INV_X1     g12447(.I(new_n12703_), .ZN(new_n12704_));
  NOR2_X1    g12448(.A1(new_n12702_), .A2(new_n12699_), .ZN(new_n12705_));
  NOR3_X1    g12449(.A1(new_n12704_), .A2(new_n12695_), .A3(new_n12705_), .ZN(new_n12706_));
  XOR2_X1    g12450(.A1(new_n12692_), .A2(new_n12694_), .Z(new_n12707_));
  OR2_X2     g12451(.A1(new_n12702_), .A2(new_n12699_), .Z(new_n12708_));
  AOI21_X1   g12452(.A1(new_n12708_), .A2(new_n12703_), .B(new_n12707_), .ZN(new_n12709_));
  NOR2_X1    g12453(.A1(new_n12706_), .A2(new_n12709_), .ZN(new_n12710_));
  INV_X1     g12454(.I(new_n12710_), .ZN(new_n12711_));
  AOI22_X1   g12455(.A1(new_n2716_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n2719_), .ZN(new_n12712_));
  OAI21_X1   g12456(.A1(new_n5312_), .A2(new_n2924_), .B(new_n12712_), .ZN(new_n12713_));
  AOI21_X1   g12457(.A1(new_n6310_), .A2(new_n2722_), .B(new_n12713_), .ZN(new_n12714_));
  XOR2_X1    g12458(.A1(new_n12714_), .A2(new_n2714_), .Z(new_n12715_));
  INV_X1     g12459(.I(new_n12715_), .ZN(new_n12716_));
  NOR2_X1    g12460(.A1(new_n12445_), .A2(new_n12447_), .ZN(new_n12717_));
  NOR2_X1    g12461(.A1(new_n12717_), .A2(new_n12716_), .ZN(new_n12718_));
  NAND2_X1   g12462(.A1(new_n12452_), .A2(new_n12441_), .ZN(new_n12719_));
  NOR2_X1    g12463(.A1(new_n12719_), .A2(new_n12715_), .ZN(new_n12720_));
  NOR3_X1    g12464(.A1(new_n12711_), .A2(new_n12718_), .A3(new_n12720_), .ZN(new_n12721_));
  NOR2_X1    g12465(.A1(new_n12718_), .A2(new_n12720_), .ZN(new_n12722_));
  NOR2_X1    g12466(.A1(new_n12722_), .A2(new_n12710_), .ZN(new_n12723_));
  NOR2_X1    g12467(.A1(new_n12723_), .A2(new_n12721_), .ZN(new_n12724_));
  AOI22_X1   g12468(.A1(new_n2202_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n2205_), .ZN(new_n12725_));
  OAI21_X1   g12469(.A1(new_n6284_), .A2(new_n2370_), .B(new_n12725_), .ZN(new_n12726_));
  AOI21_X1   g12470(.A1(new_n7106_), .A2(new_n2208_), .B(new_n12726_), .ZN(new_n12727_));
  XOR2_X1    g12471(.A1(new_n12727_), .A2(new_n2200_), .Z(new_n12728_));
  NAND2_X1   g12472(.A1(new_n12469_), .A2(new_n12458_), .ZN(new_n12729_));
  NAND2_X1   g12473(.A1(new_n12729_), .A2(new_n12728_), .ZN(new_n12730_));
  NOR2_X1    g12474(.A1(new_n12729_), .A2(new_n12728_), .ZN(new_n12731_));
  INV_X1     g12475(.I(new_n12731_), .ZN(new_n12732_));
  NAND3_X1   g12476(.A1(new_n12732_), .A2(new_n12730_), .A3(new_n12724_), .ZN(new_n12733_));
  AOI21_X1   g12477(.A1(new_n12732_), .A2(new_n12730_), .B(new_n12724_), .ZN(new_n12734_));
  INV_X1     g12478(.I(new_n12734_), .ZN(new_n12735_));
  AOI21_X1   g12479(.A1(new_n12735_), .A2(new_n12733_), .B(new_n12560_), .ZN(new_n12736_));
  INV_X1     g12480(.I(new_n12560_), .ZN(new_n12737_));
  INV_X1     g12481(.I(new_n12724_), .ZN(new_n12738_));
  INV_X1     g12482(.I(new_n12730_), .ZN(new_n12739_));
  NOR3_X1    g12483(.A1(new_n12739_), .A2(new_n12738_), .A3(new_n12731_), .ZN(new_n12740_));
  NOR3_X1    g12484(.A1(new_n12734_), .A2(new_n12740_), .A3(new_n12737_), .ZN(new_n12741_));
  NOR3_X1    g12485(.A1(new_n12736_), .A2(new_n12556_), .A3(new_n12741_), .ZN(new_n12742_));
  OAI21_X1   g12486(.A1(new_n12734_), .A2(new_n12740_), .B(new_n12737_), .ZN(new_n12743_));
  NAND3_X1   g12487(.A1(new_n12735_), .A2(new_n12733_), .A3(new_n12560_), .ZN(new_n12744_));
  AOI21_X1   g12488(.A1(new_n12743_), .A2(new_n12744_), .B(new_n12555_), .ZN(new_n12745_));
  NOR2_X1    g12489(.A1(new_n12742_), .A2(new_n12745_), .ZN(new_n12746_));
  INV_X1     g12490(.I(new_n12746_), .ZN(new_n12747_));
  OAI22_X1   g12491(.A1(new_n1592_), .A2(new_n8127_), .B1(new_n8126_), .B2(new_n1505_), .ZN(new_n12748_));
  AOI21_X1   g12492(.A1(\b[46] ), .A2(new_n1584_), .B(new_n12748_), .ZN(new_n12749_));
  OAI21_X1   g12493(.A1(new_n8138_), .A2(new_n1732_), .B(new_n12749_), .ZN(new_n12750_));
  XOR2_X1    g12494(.A1(new_n12750_), .A2(\a[17] ), .Z(new_n12751_));
  NAND2_X1   g12495(.A1(new_n12481_), .A2(new_n12475_), .ZN(new_n12752_));
  NAND2_X1   g12496(.A1(new_n12752_), .A2(new_n12751_), .ZN(new_n12753_));
  INV_X1     g12497(.I(new_n12753_), .ZN(new_n12754_));
  NOR2_X1    g12498(.A1(new_n12752_), .A2(new_n12751_), .ZN(new_n12755_));
  NOR3_X1    g12499(.A1(new_n12754_), .A2(new_n12747_), .A3(new_n12755_), .ZN(new_n12756_));
  INV_X1     g12500(.I(new_n12755_), .ZN(new_n12757_));
  AOI21_X1   g12501(.A1(new_n12757_), .A2(new_n12753_), .B(new_n12746_), .ZN(new_n12758_));
  NOR2_X1    g12502(.A1(new_n12758_), .A2(new_n12756_), .ZN(new_n12759_));
  OAI22_X1   g12503(.A1(new_n993_), .A2(new_n8776_), .B1(new_n8500_), .B2(new_n997_), .ZN(new_n12760_));
  AOI21_X1   g12504(.A1(\b[49] ), .A2(new_n1486_), .B(new_n12760_), .ZN(new_n12761_));
  OAI21_X1   g12505(.A1(new_n11577_), .A2(new_n1323_), .B(new_n12761_), .ZN(new_n12762_));
  XOR2_X1    g12506(.A1(new_n12762_), .A2(\a[14] ), .Z(new_n12763_));
  OAI21_X1   g12507(.A1(new_n12490_), .A2(new_n12493_), .B(new_n12763_), .ZN(new_n12764_));
  INV_X1     g12508(.I(new_n12763_), .ZN(new_n12765_));
  NAND3_X1   g12509(.A1(new_n12497_), .A2(new_n12488_), .A3(new_n12765_), .ZN(new_n12766_));
  NAND3_X1   g12510(.A1(new_n12764_), .A2(new_n12766_), .A3(new_n12759_), .ZN(new_n12767_));
  OR2_X2     g12511(.A1(new_n12758_), .A2(new_n12756_), .Z(new_n12768_));
  AOI21_X1   g12512(.A1(new_n12497_), .A2(new_n12488_), .B(new_n12765_), .ZN(new_n12769_));
  NOR3_X1    g12513(.A1(new_n12490_), .A2(new_n12493_), .A3(new_n12763_), .ZN(new_n12770_));
  OAI21_X1   g12514(.A1(new_n12770_), .A2(new_n12769_), .B(new_n12768_), .ZN(new_n12771_));
  NAND3_X1   g12515(.A1(new_n12771_), .A2(new_n12767_), .A3(new_n12553_), .ZN(new_n12772_));
  NOR3_X1    g12516(.A1(new_n12768_), .A2(new_n12770_), .A3(new_n12769_), .ZN(new_n12773_));
  AOI21_X1   g12517(.A1(new_n12764_), .A2(new_n12766_), .B(new_n12759_), .ZN(new_n12774_));
  OAI21_X1   g12518(.A1(new_n12773_), .A2(new_n12774_), .B(new_n12552_), .ZN(new_n12775_));
  NAND2_X1   g12519(.A1(new_n12772_), .A2(new_n12775_), .ZN(new_n12776_));
  NOR2_X1    g12520(.A1(new_n12507_), .A2(new_n12496_), .ZN(new_n12777_));
  NAND2_X1   g12521(.A1(new_n12776_), .A2(new_n12777_), .ZN(new_n12778_));
  NOR3_X1    g12522(.A1(new_n12773_), .A2(new_n12774_), .A3(new_n12552_), .ZN(new_n12779_));
  AOI21_X1   g12523(.A1(new_n12771_), .A2(new_n12767_), .B(new_n12553_), .ZN(new_n12780_));
  NOR2_X1    g12524(.A1(new_n12780_), .A2(new_n12779_), .ZN(new_n12781_));
  NAND2_X1   g12525(.A1(new_n12501_), .A2(new_n12502_), .ZN(new_n12782_));
  NAND2_X1   g12526(.A1(new_n12781_), .A2(new_n12782_), .ZN(new_n12783_));
  NAND3_X1   g12527(.A1(new_n12783_), .A2(new_n12778_), .A3(new_n12548_), .ZN(new_n12784_));
  INV_X1     g12528(.I(new_n12548_), .ZN(new_n12785_));
  NOR2_X1    g12529(.A1(new_n12781_), .A2(new_n12782_), .ZN(new_n12786_));
  NOR2_X1    g12530(.A1(new_n12776_), .A2(new_n12777_), .ZN(new_n12787_));
  OAI21_X1   g12531(.A1(new_n12786_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n12788_));
  NAND3_X1   g12532(.A1(new_n12788_), .A2(new_n12784_), .A3(new_n12544_), .ZN(new_n12789_));
  NOR3_X1    g12533(.A1(new_n12786_), .A2(new_n12787_), .A3(new_n12785_), .ZN(new_n12790_));
  AOI21_X1   g12534(.A1(new_n12783_), .A2(new_n12778_), .B(new_n12548_), .ZN(new_n12791_));
  OAI21_X1   g12535(.A1(new_n12791_), .A2(new_n12790_), .B(new_n12543_), .ZN(new_n12792_));
  NOR2_X1    g12536(.A1(new_n284_), .A2(new_n12148_), .ZN(new_n12793_));
  INV_X1     g12537(.I(new_n12793_), .ZN(new_n12794_));
  AOI22_X1   g12538(.A1(new_n267_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n261_), .ZN(new_n12795_));
  INV_X1     g12539(.I(\b[62] ), .ZN(new_n12796_));
  NAND2_X1   g12540(.A1(new_n12148_), .A2(new_n12796_), .ZN(new_n12797_));
  OAI22_X1   g12541(.A1(new_n12513_), .A2(new_n12515_), .B1(new_n12148_), .B2(new_n12796_), .ZN(new_n12798_));
  NAND2_X1   g12542(.A1(new_n12798_), .A2(new_n12797_), .ZN(new_n12799_));
  INV_X1     g12543(.I(\b[63] ), .ZN(new_n12800_));
  NOR2_X1    g12544(.A1(new_n12800_), .A2(\b[62] ), .ZN(new_n12801_));
  NOR2_X1    g12545(.A1(new_n12796_), .A2(\b[63] ), .ZN(new_n12802_));
  NOR3_X1    g12546(.A1(new_n12799_), .A2(new_n12801_), .A3(new_n12802_), .ZN(new_n12803_));
  INV_X1     g12547(.I(new_n12799_), .ZN(new_n12804_));
  NOR2_X1    g12548(.A1(new_n12801_), .A2(new_n12802_), .ZN(new_n12805_));
  NOR2_X1    g12549(.A1(new_n12804_), .A2(new_n12805_), .ZN(new_n12806_));
  OAI21_X1   g12550(.A1(new_n12806_), .A2(new_n12803_), .B(new_n265_), .ZN(new_n12807_));
  NAND3_X1   g12551(.A1(new_n12807_), .A2(new_n12794_), .A3(new_n12795_), .ZN(new_n12808_));
  NAND2_X1   g12552(.A1(new_n12808_), .A2(\a[2] ), .ZN(new_n12809_));
  INV_X1     g12553(.I(new_n12795_), .ZN(new_n12810_));
  XOR2_X1    g12554(.A1(new_n12799_), .A2(new_n12805_), .Z(new_n12811_));
  AOI21_X1   g12555(.A1(new_n12811_), .A2(new_n265_), .B(new_n12810_), .ZN(new_n12812_));
  NAND3_X1   g12556(.A1(new_n12812_), .A2(new_n270_), .A3(new_n12794_), .ZN(new_n12813_));
  AOI22_X1   g12557(.A1(new_n800_), .A2(\b[59] ), .B1(\b[60] ), .B2(new_n333_), .ZN(new_n12814_));
  OAI21_X1   g12558(.A1(new_n11195_), .A2(new_n392_), .B(new_n12814_), .ZN(new_n12815_));
  AOI21_X1   g12559(.A1(new_n11836_), .A2(new_n330_), .B(new_n12815_), .ZN(new_n12816_));
  XOR2_X1    g12560(.A1(new_n12816_), .A2(new_n312_), .Z(new_n12817_));
  INV_X1     g12561(.I(new_n12817_), .ZN(new_n12818_));
  AOI21_X1   g12562(.A1(new_n12809_), .A2(new_n12813_), .B(new_n12818_), .ZN(new_n12819_));
  AOI21_X1   g12563(.A1(new_n12812_), .A2(new_n12794_), .B(new_n270_), .ZN(new_n12820_));
  NOR2_X1    g12564(.A1(new_n12808_), .A2(\a[2] ), .ZN(new_n12821_));
  NOR3_X1    g12565(.A1(new_n12821_), .A2(new_n12820_), .A3(new_n12817_), .ZN(new_n12822_));
  NOR2_X1    g12566(.A1(new_n12822_), .A2(new_n12819_), .ZN(new_n12823_));
  NAND3_X1   g12567(.A1(new_n12792_), .A2(new_n12789_), .A3(new_n12823_), .ZN(new_n12824_));
  NOR3_X1    g12568(.A1(new_n12791_), .A2(new_n12790_), .A3(new_n12543_), .ZN(new_n12825_));
  AOI21_X1   g12569(.A1(new_n12788_), .A2(new_n12784_), .B(new_n12544_), .ZN(new_n12826_));
  OAI21_X1   g12570(.A1(new_n12821_), .A2(new_n12820_), .B(new_n12817_), .ZN(new_n12827_));
  NAND3_X1   g12571(.A1(new_n12809_), .A2(new_n12813_), .A3(new_n12818_), .ZN(new_n12828_));
  NAND2_X1   g12572(.A1(new_n12827_), .A2(new_n12828_), .ZN(new_n12829_));
  OAI21_X1   g12573(.A1(new_n12825_), .A2(new_n12826_), .B(new_n12829_), .ZN(new_n12830_));
  AOI21_X1   g12574(.A1(new_n12202_), .A2(new_n12529_), .B(new_n12527_), .ZN(new_n12831_));
  AOI21_X1   g12575(.A1(new_n12830_), .A2(new_n12824_), .B(new_n12831_), .ZN(new_n12832_));
  NOR3_X1    g12576(.A1(new_n12825_), .A2(new_n12826_), .A3(new_n12829_), .ZN(new_n12833_));
  AOI21_X1   g12577(.A1(new_n12792_), .A2(new_n12789_), .B(new_n12823_), .ZN(new_n12834_));
  INV_X1     g12578(.I(new_n12831_), .ZN(new_n12835_));
  NOR3_X1    g12579(.A1(new_n12833_), .A2(new_n12834_), .A3(new_n12835_), .ZN(new_n12836_));
  NOR2_X1    g12580(.A1(new_n12832_), .A2(new_n12836_), .ZN(new_n12837_));
  INV_X1     g12581(.I(new_n12538_), .ZN(new_n12838_));
  OAI21_X1   g12582(.A1(new_n12196_), .A2(new_n12838_), .B(new_n12537_), .ZN(new_n12839_));
  XOR2_X1    g12583(.A1(new_n12839_), .A2(new_n12837_), .Z(\f[63] ));
  OAI21_X1   g12584(.A1(new_n12782_), .A2(new_n12780_), .B(new_n12772_), .ZN(new_n12841_));
  AOI22_X1   g12585(.A1(new_n518_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n636_), .ZN(new_n12842_));
  OAI21_X1   g12586(.A1(new_n10308_), .A2(new_n917_), .B(new_n12842_), .ZN(new_n12843_));
  AOI21_X1   g12587(.A1(new_n12164_), .A2(new_n618_), .B(new_n12843_), .ZN(new_n12844_));
  XOR2_X1    g12588(.A1(new_n12844_), .A2(new_n488_), .Z(new_n12845_));
  INV_X1     g12589(.I(new_n12845_), .ZN(new_n12846_));
  NOR2_X1    g12590(.A1(new_n12768_), .A2(new_n12769_), .ZN(new_n12847_));
  OAI22_X1   g12591(.A1(new_n993_), .A2(new_n9032_), .B1(new_n8776_), .B2(new_n997_), .ZN(new_n12848_));
  AOI21_X1   g12592(.A1(\b[50] ), .A2(new_n1486_), .B(new_n12848_), .ZN(new_n12849_));
  OAI21_X1   g12593(.A1(new_n9043_), .A2(new_n1323_), .B(new_n12849_), .ZN(new_n12850_));
  XOR2_X1    g12594(.A1(new_n12850_), .A2(\a[14] ), .Z(new_n12851_));
  NAND2_X1   g12595(.A1(new_n12753_), .A2(new_n12746_), .ZN(new_n12852_));
  OAI22_X1   g12596(.A1(new_n1592_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n1505_), .ZN(new_n12853_));
  AOI21_X1   g12597(.A1(\b[47] ), .A2(new_n1584_), .B(new_n12853_), .ZN(new_n12854_));
  OAI21_X1   g12598(.A1(new_n9050_), .A2(new_n1732_), .B(new_n12854_), .ZN(new_n12855_));
  XOR2_X1    g12599(.A1(new_n12855_), .A2(\a[17] ), .Z(new_n12856_));
  AOI21_X1   g12600(.A1(new_n12555_), .A2(new_n12744_), .B(new_n12736_), .ZN(new_n12857_));
  AOI22_X1   g12601(.A1(new_n1738_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n1743_), .ZN(new_n12858_));
  OAI21_X1   g12602(.A1(new_n7074_), .A2(new_n1931_), .B(new_n12858_), .ZN(new_n12859_));
  AOI21_X1   g12603(.A1(new_n9337_), .A2(new_n1746_), .B(new_n12859_), .ZN(new_n12860_));
  XOR2_X1    g12604(.A1(new_n12860_), .A2(new_n1736_), .Z(new_n12861_));
  AOI21_X1   g12605(.A1(new_n12738_), .A2(new_n12730_), .B(new_n12731_), .ZN(new_n12862_));
  INV_X1     g12606(.I(new_n12862_), .ZN(new_n12863_));
  AOI21_X1   g12607(.A1(new_n12719_), .A2(new_n12715_), .B(new_n12710_), .ZN(new_n12864_));
  AOI21_X1   g12608(.A1(new_n12695_), .A2(new_n12703_), .B(new_n12705_), .ZN(new_n12865_));
  NOR3_X1    g12609(.A1(new_n12864_), .A2(new_n12720_), .A3(new_n12865_), .ZN(new_n12866_));
  OAI21_X1   g12610(.A1(new_n12864_), .A2(new_n12720_), .B(new_n12865_), .ZN(new_n12867_));
  INV_X1     g12611(.I(new_n12867_), .ZN(new_n12868_));
  AOI22_X1   g12612(.A1(new_n2716_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n2719_), .ZN(new_n12869_));
  OAI21_X1   g12613(.A1(new_n5341_), .A2(new_n2924_), .B(new_n12869_), .ZN(new_n12870_));
  AOI21_X1   g12614(.A1(new_n5793_), .A2(new_n2722_), .B(new_n12870_), .ZN(new_n12871_));
  XOR2_X1    g12615(.A1(new_n12871_), .A2(new_n2714_), .Z(new_n12872_));
  OAI22_X1   g12616(.A1(new_n5312_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n4886_), .ZN(new_n12873_));
  AOI21_X1   g12617(.A1(\b[35] ), .A2(new_n3456_), .B(new_n12873_), .ZN(new_n12874_));
  OAI21_X1   g12618(.A1(new_n5322_), .A2(new_n3261_), .B(new_n12874_), .ZN(new_n12875_));
  XOR2_X1    g12619(.A1(new_n12875_), .A2(\a[29] ), .Z(new_n12876_));
  INV_X1     g12620(.I(new_n12691_), .ZN(new_n12877_));
  AOI22_X1   g12621(.A1(new_n3864_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n3869_), .ZN(new_n12878_));
  OAI21_X1   g12622(.A1(new_n4023_), .A2(new_n5410_), .B(new_n12878_), .ZN(new_n12879_));
  AOI21_X1   g12623(.A1(new_n5103_), .A2(new_n3872_), .B(new_n12879_), .ZN(new_n12880_));
  XOR2_X1    g12624(.A1(new_n12880_), .A2(new_n3876_), .Z(new_n12881_));
  NAND2_X1   g12625(.A1(new_n12681_), .A2(new_n12675_), .ZN(new_n12882_));
  AOI21_X1   g12626(.A1(new_n12670_), .A2(new_n12666_), .B(new_n12662_), .ZN(new_n12883_));
  OAI21_X1   g12627(.A1(new_n12648_), .A2(new_n12654_), .B(new_n12655_), .ZN(new_n12884_));
  INV_X1     g12628(.I(new_n12884_), .ZN(new_n12885_));
  NOR3_X1    g12629(.A1(new_n12883_), .A2(new_n12671_), .A3(new_n12885_), .ZN(new_n12886_));
  NAND2_X1   g12630(.A1(new_n12668_), .A2(new_n12667_), .ZN(new_n12887_));
  OAI21_X1   g12631(.A1(new_n12668_), .A2(new_n12667_), .B(new_n12661_), .ZN(new_n12888_));
  AOI21_X1   g12632(.A1(new_n12888_), .A2(new_n12887_), .B(new_n12884_), .ZN(new_n12889_));
  NAND2_X1   g12633(.A1(new_n12566_), .A2(new_n12646_), .ZN(new_n12890_));
  NAND2_X1   g12634(.A1(new_n12890_), .A2(new_n12645_), .ZN(new_n12891_));
  OAI22_X1   g12635(.A1(new_n5852_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n5857_), .ZN(new_n12892_));
  AOI21_X1   g12636(.A1(\b[23] ), .A2(new_n6115_), .B(new_n12892_), .ZN(new_n12893_));
  OAI21_X1   g12637(.A1(new_n2655_), .A2(new_n5861_), .B(new_n12893_), .ZN(new_n12894_));
  XOR2_X1    g12638(.A1(new_n12894_), .A2(\a[41] ), .Z(new_n12895_));
  AOI22_X1   g12639(.A1(new_n6569_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n6574_), .ZN(new_n12896_));
  OAI21_X1   g12640(.A1(new_n1860_), .A2(new_n8565_), .B(new_n12896_), .ZN(new_n12897_));
  AOI21_X1   g12641(.A1(new_n2659_), .A2(new_n6579_), .B(new_n12897_), .ZN(new_n12898_));
  XOR2_X1    g12642(.A1(new_n12898_), .A2(new_n6567_), .Z(new_n12899_));
  NOR2_X1    g12643(.A1(new_n12637_), .A2(new_n12630_), .ZN(new_n12900_));
  NOR2_X1    g12644(.A1(new_n12900_), .A2(new_n12642_), .ZN(new_n12901_));
  NAND2_X1   g12645(.A1(new_n12626_), .A2(new_n12619_), .ZN(new_n12902_));
  NAND2_X1   g12646(.A1(new_n12902_), .A2(new_n12627_), .ZN(new_n12903_));
  AOI21_X1   g12647(.A1(new_n12614_), .A2(new_n12613_), .B(new_n12609_), .ZN(new_n12904_));
  NOR2_X1    g12648(.A1(new_n12904_), .A2(new_n12616_), .ZN(new_n12905_));
  NOR2_X1    g12649(.A1(new_n12903_), .A2(new_n12905_), .ZN(new_n12906_));
  INV_X1     g12650(.I(new_n12905_), .ZN(new_n12907_));
  AOI21_X1   g12651(.A1(new_n12902_), .A2(new_n12627_), .B(new_n12907_), .ZN(new_n12908_));
  AOI22_X1   g12652(.A1(new_n8241_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n8246_), .ZN(new_n12909_));
  OAI21_X1   g12653(.A1(new_n1093_), .A2(new_n9114_), .B(new_n12909_), .ZN(new_n12910_));
  AOI21_X1   g12654(.A1(new_n1701_), .A2(new_n8252_), .B(new_n12910_), .ZN(new_n12911_));
  XOR2_X1    g12655(.A1(new_n12911_), .A2(new_n8248_), .Z(new_n12912_));
  NAND2_X1   g12656(.A1(new_n12607_), .A2(new_n12574_), .ZN(new_n12913_));
  NAND2_X1   g12657(.A1(new_n12913_), .A2(new_n12606_), .ZN(new_n12914_));
  OAI21_X1   g12658(.A1(new_n12576_), .A2(new_n12597_), .B(new_n12596_), .ZN(new_n12915_));
  NOR2_X1    g12659(.A1(new_n12322_), .A2(new_n12586_), .ZN(new_n12916_));
  NOR2_X1    g12660(.A1(new_n12916_), .A2(new_n12587_), .ZN(new_n12917_));
  AOI22_X1   g12661(.A1(new_n11926_), .A2(\b[4] ), .B1(new_n11924_), .B2(\b[3] ), .ZN(new_n12918_));
  OAI21_X1   g12662(.A1(new_n276_), .A2(new_n12317_), .B(new_n12918_), .ZN(new_n12919_));
  AOI21_X1   g12663(.A1(new_n1725_), .A2(new_n11929_), .B(new_n12919_), .ZN(new_n12920_));
  XOR2_X1    g12664(.A1(new_n12920_), .A2(new_n12312_), .Z(new_n12921_));
  INV_X1     g12665(.I(new_n12584_), .ZN(new_n12922_));
  NOR2_X1    g12666(.A1(new_n12312_), .A2(new_n12581_), .ZN(new_n12923_));
  AOI22_X1   g12667(.A1(new_n12922_), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n12923_), .ZN(new_n12924_));
  INV_X1     g12668(.I(new_n12924_), .ZN(new_n12925_));
  NOR2_X1    g12669(.A1(new_n12921_), .A2(new_n12925_), .ZN(new_n12926_));
  NAND2_X1   g12670(.A1(new_n12921_), .A2(new_n12925_), .ZN(new_n12927_));
  INV_X1     g12671(.I(new_n12927_), .ZN(new_n12928_));
  NOR2_X1    g12672(.A1(new_n12928_), .A2(new_n12926_), .ZN(new_n12929_));
  XNOR2_X1   g12673(.A1(new_n12917_), .A2(new_n12929_), .ZN(new_n12930_));
  OAI22_X1   g12674(.A1(new_n12306_), .A2(new_n471_), .B1(new_n12305_), .B2(new_n438_), .ZN(new_n12931_));
  AOI21_X1   g12675(.A1(\b[5] ), .A2(new_n12304_), .B(new_n12931_), .ZN(new_n12932_));
  OAI21_X1   g12676(.A1(new_n485_), .A2(new_n10985_), .B(new_n12932_), .ZN(new_n12933_));
  XOR2_X1    g12677(.A1(new_n12933_), .A2(\a[59] ), .Z(new_n12934_));
  INV_X1     g12678(.I(new_n12934_), .ZN(new_n12935_));
  NAND2_X1   g12679(.A1(new_n12930_), .A2(new_n12935_), .ZN(new_n12936_));
  OR2_X2     g12680(.A1(new_n12930_), .A2(new_n12935_), .Z(new_n12937_));
  NAND2_X1   g12681(.A1(new_n12937_), .A2(new_n12936_), .ZN(new_n12938_));
  XNOR2_X1   g12682(.A1(new_n12938_), .A2(new_n12915_), .ZN(new_n12939_));
  AOI22_X1   g12683(.A1(new_n10064_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n10062_), .ZN(new_n12940_));
  OAI21_X1   g12684(.A1(new_n577_), .A2(new_n10399_), .B(new_n12940_), .ZN(new_n12941_));
  AOI21_X1   g12685(.A1(new_n1059_), .A2(new_n10068_), .B(new_n12941_), .ZN(new_n12942_));
  XOR2_X1    g12686(.A1(new_n12942_), .A2(new_n10057_), .Z(new_n12943_));
  INV_X1     g12687(.I(new_n12943_), .ZN(new_n12944_));
  NAND2_X1   g12688(.A1(new_n12939_), .A2(new_n12944_), .ZN(new_n12945_));
  NOR2_X1    g12689(.A1(new_n12939_), .A2(new_n12944_), .ZN(new_n12946_));
  INV_X1     g12690(.I(new_n12946_), .ZN(new_n12947_));
  NAND2_X1   g12691(.A1(new_n12947_), .A2(new_n12945_), .ZN(new_n12948_));
  XOR2_X1    g12692(.A1(new_n12914_), .A2(new_n12948_), .Z(new_n12949_));
  OAI22_X1   g12693(.A1(new_n10390_), .A2(new_n1070_), .B1(new_n941_), .B2(new_n10389_), .ZN(new_n12950_));
  AOI21_X1   g12694(.A1(\b[11] ), .A2(new_n9471_), .B(new_n12950_), .ZN(new_n12951_));
  OAI21_X1   g12695(.A1(new_n1082_), .A2(new_n10388_), .B(new_n12951_), .ZN(new_n12952_));
  XOR2_X1    g12696(.A1(new_n12952_), .A2(\a[53] ), .Z(new_n12953_));
  NOR2_X1    g12697(.A1(new_n12949_), .A2(new_n12953_), .ZN(new_n12954_));
  AND2_X2    g12698(.A1(new_n12949_), .A2(new_n12953_), .Z(new_n12955_));
  NOR2_X1    g12699(.A1(new_n12955_), .A2(new_n12954_), .ZN(new_n12956_));
  XOR2_X1    g12700(.A1(new_n12956_), .A2(new_n12912_), .Z(new_n12957_));
  INV_X1     g12701(.I(new_n12957_), .ZN(new_n12958_));
  NOR3_X1    g12702(.A1(new_n12906_), .A2(new_n12908_), .A3(new_n12958_), .ZN(new_n12959_));
  INV_X1     g12703(.I(new_n12959_), .ZN(new_n12960_));
  OAI21_X1   g12704(.A1(new_n12906_), .A2(new_n12908_), .B(new_n12958_), .ZN(new_n12961_));
  AOI22_X1   g12705(.A1(new_n7403_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n7408_), .ZN(new_n12962_));
  OAI21_X1   g12706(.A1(new_n1432_), .A2(new_n9488_), .B(new_n12962_), .ZN(new_n12963_));
  AOI21_X1   g12707(.A1(new_n1695_), .A2(new_n7414_), .B(new_n12963_), .ZN(new_n12964_));
  XOR2_X1    g12708(.A1(new_n12964_), .A2(new_n7410_), .Z(new_n12965_));
  INV_X1     g12709(.I(new_n12965_), .ZN(new_n12966_));
  NAND3_X1   g12710(.A1(new_n12960_), .A2(new_n12961_), .A3(new_n12966_), .ZN(new_n12967_));
  INV_X1     g12711(.I(new_n12961_), .ZN(new_n12968_));
  OAI21_X1   g12712(.A1(new_n12968_), .A2(new_n12959_), .B(new_n12965_), .ZN(new_n12969_));
  NAND3_X1   g12713(.A1(new_n12969_), .A2(new_n12967_), .A3(new_n12901_), .ZN(new_n12970_));
  NOR3_X1    g12714(.A1(new_n12968_), .A2(new_n12959_), .A3(new_n12965_), .ZN(new_n12971_));
  AOI21_X1   g12715(.A1(new_n12960_), .A2(new_n12961_), .B(new_n12966_), .ZN(new_n12972_));
  OAI22_X1   g12716(.A1(new_n12972_), .A2(new_n12971_), .B1(new_n12642_), .B2(new_n12900_), .ZN(new_n12973_));
  NAND3_X1   g12717(.A1(new_n12973_), .A2(new_n12970_), .A3(new_n12899_), .ZN(new_n12974_));
  INV_X1     g12718(.I(new_n12899_), .ZN(new_n12975_));
  INV_X1     g12719(.I(new_n12901_), .ZN(new_n12976_));
  NOR3_X1    g12720(.A1(new_n12976_), .A2(new_n12971_), .A3(new_n12972_), .ZN(new_n12977_));
  AOI21_X1   g12721(.A1(new_n12969_), .A2(new_n12967_), .B(new_n12901_), .ZN(new_n12978_));
  OAI21_X1   g12722(.A1(new_n12977_), .A2(new_n12978_), .B(new_n12975_), .ZN(new_n12979_));
  NAND2_X1   g12723(.A1(new_n12979_), .A2(new_n12974_), .ZN(new_n12980_));
  XOR2_X1    g12724(.A1(new_n12980_), .A2(new_n12895_), .Z(new_n12981_));
  NOR2_X1    g12725(.A1(new_n12981_), .A2(new_n12891_), .ZN(new_n12982_));
  INV_X1     g12726(.I(new_n12891_), .ZN(new_n12983_));
  INV_X1     g12727(.I(new_n12895_), .ZN(new_n12984_));
  XOR2_X1    g12728(.A1(new_n12980_), .A2(new_n12984_), .Z(new_n12985_));
  NOR2_X1    g12729(.A1(new_n12985_), .A2(new_n12983_), .ZN(new_n12986_));
  NOR2_X1    g12730(.A1(new_n12982_), .A2(new_n12986_), .ZN(new_n12987_));
  AOI22_X1   g12731(.A1(new_n5155_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n5160_), .ZN(new_n12988_));
  OAI21_X1   g12732(.A1(new_n3006_), .A2(new_n6877_), .B(new_n12988_), .ZN(new_n12989_));
  AOI21_X1   g12733(.A1(new_n3807_), .A2(new_n5166_), .B(new_n12989_), .ZN(new_n12990_));
  XOR2_X1    g12734(.A1(new_n12990_), .A2(new_n5162_), .Z(new_n12991_));
  XOR2_X1    g12735(.A1(new_n12987_), .A2(new_n12991_), .Z(new_n12992_));
  INV_X1     g12736(.I(new_n12992_), .ZN(new_n12993_));
  NOR3_X1    g12737(.A1(new_n12993_), .A2(new_n12886_), .A3(new_n12889_), .ZN(new_n12994_));
  INV_X1     g12738(.I(new_n12994_), .ZN(new_n12995_));
  OAI21_X1   g12739(.A1(new_n12889_), .A2(new_n12886_), .B(new_n12993_), .ZN(new_n12996_));
  AOI22_X1   g12740(.A1(new_n4918_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n4921_), .ZN(new_n12997_));
  OAI21_X1   g12741(.A1(new_n3592_), .A2(new_n6099_), .B(new_n12997_), .ZN(new_n12998_));
  AOI21_X1   g12742(.A1(new_n3796_), .A2(new_n4699_), .B(new_n12998_), .ZN(new_n12999_));
  XOR2_X1    g12743(.A1(new_n12999_), .A2(new_n4446_), .Z(new_n13000_));
  INV_X1     g12744(.I(new_n13000_), .ZN(new_n13001_));
  NAND3_X1   g12745(.A1(new_n12995_), .A2(new_n12996_), .A3(new_n13001_), .ZN(new_n13002_));
  INV_X1     g12746(.I(new_n12996_), .ZN(new_n13003_));
  OAI21_X1   g12747(.A1(new_n13003_), .A2(new_n12994_), .B(new_n13000_), .ZN(new_n13004_));
  NAND4_X1   g12748(.A1(new_n13004_), .A2(new_n13002_), .A3(new_n12882_), .A4(new_n12683_), .ZN(new_n13005_));
  NAND2_X1   g12749(.A1(new_n12882_), .A2(new_n12683_), .ZN(new_n13006_));
  NOR3_X1    g12750(.A1(new_n13003_), .A2(new_n12994_), .A3(new_n13000_), .ZN(new_n13007_));
  AOI21_X1   g12751(.A1(new_n12995_), .A2(new_n12996_), .B(new_n13001_), .ZN(new_n13008_));
  OAI21_X1   g12752(.A1(new_n13007_), .A2(new_n13008_), .B(new_n13006_), .ZN(new_n13009_));
  NAND3_X1   g12753(.A1(new_n13009_), .A2(new_n12881_), .A3(new_n13005_), .ZN(new_n13010_));
  AOI21_X1   g12754(.A1(new_n13009_), .A2(new_n13005_), .B(new_n12881_), .ZN(new_n13011_));
  INV_X1     g12755(.I(new_n13011_), .ZN(new_n13012_));
  NAND2_X1   g12756(.A1(new_n13012_), .A2(new_n13010_), .ZN(new_n13013_));
  OAI21_X1   g12757(.A1(new_n12688_), .A2(new_n12564_), .B(new_n12694_), .ZN(new_n13014_));
  NAND3_X1   g12758(.A1(new_n13013_), .A2(new_n12877_), .A3(new_n13014_), .ZN(new_n13015_));
  INV_X1     g12759(.I(new_n13010_), .ZN(new_n13016_));
  NOR2_X1    g12760(.A1(new_n13016_), .A2(new_n13011_), .ZN(new_n13017_));
  NAND2_X1   g12761(.A1(new_n13014_), .A2(new_n12877_), .ZN(new_n13018_));
  NAND2_X1   g12762(.A1(new_n13017_), .A2(new_n13018_), .ZN(new_n13019_));
  NAND3_X1   g12763(.A1(new_n13015_), .A2(new_n13019_), .A3(new_n12876_), .ZN(new_n13020_));
  INV_X1     g12764(.I(new_n12876_), .ZN(new_n13021_));
  NOR2_X1    g12765(.A1(new_n13017_), .A2(new_n13018_), .ZN(new_n13022_));
  INV_X1     g12766(.I(new_n13019_), .ZN(new_n13023_));
  OAI21_X1   g12767(.A1(new_n13023_), .A2(new_n13022_), .B(new_n13021_), .ZN(new_n13024_));
  NAND2_X1   g12768(.A1(new_n13024_), .A2(new_n13020_), .ZN(new_n13025_));
  XOR2_X1    g12769(.A1(new_n13025_), .A2(new_n12872_), .Z(new_n13026_));
  INV_X1     g12770(.I(new_n13026_), .ZN(new_n13027_));
  OAI21_X1   g12771(.A1(new_n12868_), .A2(new_n12866_), .B(new_n13027_), .ZN(new_n13028_));
  INV_X1     g12772(.I(new_n12866_), .ZN(new_n13029_));
  NAND3_X1   g12773(.A1(new_n13029_), .A2(new_n12867_), .A3(new_n13026_), .ZN(new_n13030_));
  OAI22_X1   g12774(.A1(new_n2189_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n2194_), .ZN(new_n13031_));
  AOI21_X1   g12775(.A1(\b[41] ), .A2(new_n2361_), .B(new_n13031_), .ZN(new_n13032_));
  OAI21_X1   g12776(.A1(new_n6785_), .A2(new_n2197_), .B(new_n13032_), .ZN(new_n13033_));
  XOR2_X1    g12777(.A1(new_n13033_), .A2(\a[23] ), .Z(new_n13034_));
  AOI21_X1   g12778(.A1(new_n13028_), .A2(new_n13030_), .B(new_n13034_), .ZN(new_n13035_));
  AOI21_X1   g12779(.A1(new_n13029_), .A2(new_n12867_), .B(new_n13026_), .ZN(new_n13036_));
  NOR3_X1    g12780(.A1(new_n12868_), .A2(new_n13027_), .A3(new_n12866_), .ZN(new_n13037_));
  INV_X1     g12781(.I(new_n13034_), .ZN(new_n13038_));
  NOR3_X1    g12782(.A1(new_n13036_), .A2(new_n13037_), .A3(new_n13038_), .ZN(new_n13039_));
  NOR2_X1    g12783(.A1(new_n13039_), .A2(new_n13035_), .ZN(new_n13040_));
  NAND2_X1   g12784(.A1(new_n13040_), .A2(new_n12863_), .ZN(new_n13041_));
  OAI21_X1   g12785(.A1(new_n13036_), .A2(new_n13037_), .B(new_n13038_), .ZN(new_n13042_));
  NAND3_X1   g12786(.A1(new_n13028_), .A2(new_n13030_), .A3(new_n13034_), .ZN(new_n13043_));
  NAND2_X1   g12787(.A1(new_n13042_), .A2(new_n13043_), .ZN(new_n13044_));
  NAND2_X1   g12788(.A1(new_n13044_), .A2(new_n12862_), .ZN(new_n13045_));
  NAND3_X1   g12789(.A1(new_n13041_), .A2(new_n13045_), .A3(new_n12861_), .ZN(new_n13046_));
  INV_X1     g12790(.I(new_n12861_), .ZN(new_n13047_));
  NOR2_X1    g12791(.A1(new_n13044_), .A2(new_n12862_), .ZN(new_n13048_));
  NOR2_X1    g12792(.A1(new_n13040_), .A2(new_n12863_), .ZN(new_n13049_));
  OAI21_X1   g12793(.A1(new_n13049_), .A2(new_n13048_), .B(new_n13047_), .ZN(new_n13050_));
  NAND2_X1   g12794(.A1(new_n13050_), .A2(new_n13046_), .ZN(new_n13051_));
  NAND2_X1   g12795(.A1(new_n13051_), .A2(new_n12857_), .ZN(new_n13052_));
  OAI21_X1   g12796(.A1(new_n12556_), .A2(new_n12741_), .B(new_n12743_), .ZN(new_n13053_));
  NOR3_X1    g12797(.A1(new_n13049_), .A2(new_n13048_), .A3(new_n13047_), .ZN(new_n13054_));
  AOI21_X1   g12798(.A1(new_n13041_), .A2(new_n13045_), .B(new_n12861_), .ZN(new_n13055_));
  NOR2_X1    g12799(.A1(new_n13055_), .A2(new_n13054_), .ZN(new_n13056_));
  NAND2_X1   g12800(.A1(new_n13056_), .A2(new_n13053_), .ZN(new_n13057_));
  NAND3_X1   g12801(.A1(new_n13057_), .A2(new_n13052_), .A3(new_n12856_), .ZN(new_n13058_));
  INV_X1     g12802(.I(new_n12856_), .ZN(new_n13059_));
  NOR2_X1    g12803(.A1(new_n13056_), .A2(new_n13053_), .ZN(new_n13060_));
  NOR2_X1    g12804(.A1(new_n13051_), .A2(new_n12857_), .ZN(new_n13061_));
  OAI21_X1   g12805(.A1(new_n13060_), .A2(new_n13061_), .B(new_n13059_), .ZN(new_n13062_));
  NAND4_X1   g12806(.A1(new_n13062_), .A2(new_n13058_), .A3(new_n12852_), .A4(new_n12757_), .ZN(new_n13063_));
  INV_X1     g12807(.I(new_n12852_), .ZN(new_n13064_));
  NOR3_X1    g12808(.A1(new_n13060_), .A2(new_n13061_), .A3(new_n13059_), .ZN(new_n13065_));
  AOI21_X1   g12809(.A1(new_n13057_), .A2(new_n13052_), .B(new_n12856_), .ZN(new_n13066_));
  OAI22_X1   g12810(.A1(new_n13064_), .A2(new_n12755_), .B1(new_n13066_), .B2(new_n13065_), .ZN(new_n13067_));
  AOI21_X1   g12811(.A1(new_n13067_), .A2(new_n13063_), .B(new_n12851_), .ZN(new_n13068_));
  INV_X1     g12812(.I(new_n12851_), .ZN(new_n13069_));
  NOR4_X1    g12813(.A1(new_n13064_), .A2(new_n13065_), .A3(new_n13066_), .A4(new_n12755_), .ZN(new_n13070_));
  AOI22_X1   g12814(.A1(new_n13062_), .A2(new_n13058_), .B1(new_n12757_), .B2(new_n12852_), .ZN(new_n13071_));
  NOR3_X1    g12815(.A1(new_n13070_), .A2(new_n13071_), .A3(new_n13069_), .ZN(new_n13072_));
  NOR2_X1    g12816(.A1(new_n13068_), .A2(new_n13072_), .ZN(new_n13073_));
  OAI21_X1   g12817(.A1(new_n12770_), .A2(new_n12847_), .B(new_n13073_), .ZN(new_n13074_));
  NOR2_X1    g12818(.A1(new_n12847_), .A2(new_n12770_), .ZN(new_n13075_));
  OAI21_X1   g12819(.A1(new_n13070_), .A2(new_n13071_), .B(new_n13069_), .ZN(new_n13076_));
  NAND3_X1   g12820(.A1(new_n13067_), .A2(new_n13063_), .A3(new_n12851_), .ZN(new_n13077_));
  NAND2_X1   g12821(.A1(new_n13077_), .A2(new_n13076_), .ZN(new_n13078_));
  NAND2_X1   g12822(.A1(new_n13075_), .A2(new_n13078_), .ZN(new_n13079_));
  INV_X1     g12823(.I(new_n9979_), .ZN(new_n13080_));
  OAI22_X1   g12824(.A1(new_n713_), .A2(new_n9972_), .B1(new_n9942_), .B2(new_n717_), .ZN(new_n13081_));
  AOI21_X1   g12825(.A1(\b[53] ), .A2(new_n1126_), .B(new_n13081_), .ZN(new_n13082_));
  OAI21_X1   g12826(.A1(new_n13080_), .A2(new_n986_), .B(new_n13082_), .ZN(new_n13083_));
  XOR2_X1    g12827(.A1(new_n13083_), .A2(\a[11] ), .Z(new_n13084_));
  INV_X1     g12828(.I(new_n13084_), .ZN(new_n13085_));
  NAND3_X1   g12829(.A1(new_n13074_), .A2(new_n13079_), .A3(new_n13085_), .ZN(new_n13086_));
  NOR2_X1    g12830(.A1(new_n13075_), .A2(new_n13078_), .ZN(new_n13087_));
  NOR3_X1    g12831(.A1(new_n13073_), .A2(new_n12847_), .A3(new_n12770_), .ZN(new_n13088_));
  OAI21_X1   g12832(.A1(new_n13087_), .A2(new_n13088_), .B(new_n13084_), .ZN(new_n13089_));
  NAND3_X1   g12833(.A1(new_n13086_), .A2(new_n13089_), .A3(new_n12846_), .ZN(new_n13090_));
  NOR3_X1    g12834(.A1(new_n13087_), .A2(new_n13088_), .A3(new_n13084_), .ZN(new_n13091_));
  AOI21_X1   g12835(.A1(new_n13074_), .A2(new_n13079_), .B(new_n13085_), .ZN(new_n13092_));
  OAI21_X1   g12836(.A1(new_n13092_), .A2(new_n13091_), .B(new_n12845_), .ZN(new_n13093_));
  NAND3_X1   g12837(.A1(new_n13093_), .A2(new_n13090_), .A3(new_n12841_), .ZN(new_n13094_));
  AOI21_X1   g12838(.A1(new_n12777_), .A2(new_n12775_), .B(new_n12779_), .ZN(new_n13095_));
  NOR3_X1    g12839(.A1(new_n13092_), .A2(new_n13091_), .A3(new_n12845_), .ZN(new_n13096_));
  AOI21_X1   g12840(.A1(new_n13086_), .A2(new_n13089_), .B(new_n12846_), .ZN(new_n13097_));
  OAI21_X1   g12841(.A1(new_n13097_), .A2(new_n13096_), .B(new_n13095_), .ZN(new_n13098_));
  NAND2_X1   g12842(.A1(new_n13098_), .A2(new_n13094_), .ZN(new_n13099_));
  AOI21_X1   g12843(.A1(new_n12784_), .A2(new_n12818_), .B(new_n12791_), .ZN(new_n13100_));
  NOR2_X1    g12844(.A1(new_n13099_), .A2(new_n13100_), .ZN(new_n13101_));
  NAND2_X1   g12845(.A1(new_n13099_), .A2(new_n13100_), .ZN(new_n13102_));
  INV_X1     g12846(.I(new_n13102_), .ZN(new_n13103_));
  AOI22_X1   g12847(.A1(new_n283_), .A2(\b[62] ), .B1(new_n261_), .B2(\b[63] ), .ZN(new_n13104_));
  NOR3_X1    g12848(.A1(new_n12799_), .A2(new_n12796_), .A3(\b[63] ), .ZN(new_n13105_));
  NOR3_X1    g12849(.A1(new_n12804_), .A2(\b[62] ), .A3(new_n12800_), .ZN(new_n13106_));
  NOR2_X1    g12850(.A1(new_n13106_), .A2(new_n13105_), .ZN(new_n13107_));
  OAI21_X1   g12851(.A1(new_n13107_), .A2(new_n279_), .B(new_n13104_), .ZN(new_n13108_));
  XOR2_X1    g12852(.A1(new_n13108_), .A2(new_n270_), .Z(new_n13109_));
  NAND2_X1   g12853(.A1(new_n12158_), .A2(new_n12159_), .ZN(new_n13110_));
  OAI22_X1   g12854(.A1(new_n321_), .A2(new_n12148_), .B1(new_n325_), .B2(new_n12147_), .ZN(new_n13111_));
  AOI21_X1   g12855(.A1(\b[59] ), .A2(new_n602_), .B(new_n13111_), .ZN(new_n13112_));
  OAI21_X1   g12856(.A1(new_n13110_), .A2(new_n318_), .B(new_n13112_), .ZN(new_n13113_));
  XOR2_X1    g12857(.A1(new_n13113_), .A2(\a[5] ), .Z(new_n13114_));
  INV_X1     g12858(.I(new_n13114_), .ZN(new_n13115_));
  XOR2_X1    g12859(.A1(new_n13109_), .A2(new_n13115_), .Z(new_n13116_));
  INV_X1     g12860(.I(new_n13116_), .ZN(new_n13117_));
  OAI21_X1   g12861(.A1(new_n13103_), .A2(new_n13101_), .B(new_n13117_), .ZN(new_n13118_));
  INV_X1     g12862(.I(new_n13101_), .ZN(new_n13119_));
  NAND3_X1   g12863(.A1(new_n13119_), .A2(new_n13116_), .A3(new_n13102_), .ZN(new_n13120_));
  NAND2_X1   g12864(.A1(new_n13118_), .A2(new_n13120_), .ZN(new_n13121_));
  NOR2_X1    g12865(.A1(new_n12821_), .A2(new_n12820_), .ZN(new_n13122_));
  NOR2_X1    g12866(.A1(new_n13122_), .A2(new_n12543_), .ZN(new_n13123_));
  NAND2_X1   g12867(.A1(new_n13122_), .A2(new_n12543_), .ZN(new_n13124_));
  NAND2_X1   g12868(.A1(new_n12788_), .A2(new_n12784_), .ZN(new_n13125_));
  XOR2_X1    g12869(.A1(new_n13125_), .A2(new_n12817_), .Z(new_n13126_));
  AOI21_X1   g12870(.A1(new_n13126_), .A2(new_n13124_), .B(new_n13123_), .ZN(new_n13127_));
  INV_X1     g12871(.I(new_n13127_), .ZN(new_n13128_));
  AOI21_X1   g12872(.A1(new_n12839_), .A2(new_n12837_), .B(new_n12836_), .ZN(new_n13129_));
  NOR2_X1    g12873(.A1(new_n13129_), .A2(new_n13128_), .ZN(new_n13130_));
  INV_X1     g12874(.I(new_n12836_), .ZN(new_n13131_));
  NOR3_X1    g12875(.A1(new_n11865_), .A2(new_n12181_), .A3(new_n12184_), .ZN(new_n13132_));
  AOI21_X1   g12876(.A1(new_n12179_), .A2(new_n12185_), .B(new_n13132_), .ZN(new_n13133_));
  AOI21_X1   g12877(.A1(new_n12530_), .A2(new_n12535_), .B(new_n12197_), .ZN(new_n13134_));
  AOI21_X1   g12878(.A1(new_n13133_), .A2(new_n12538_), .B(new_n13134_), .ZN(new_n13135_));
  OAI21_X1   g12879(.A1(new_n13135_), .A2(new_n12832_), .B(new_n13131_), .ZN(new_n13136_));
  NOR2_X1    g12880(.A1(new_n13136_), .A2(new_n13127_), .ZN(new_n13137_));
  NOR2_X1    g12881(.A1(new_n13137_), .A2(new_n13130_), .ZN(new_n13138_));
  XOR2_X1    g12882(.A1(new_n13138_), .A2(new_n13121_), .Z(\f[64] ));
  AOI21_X1   g12883(.A1(new_n13136_), .A2(new_n13127_), .B(new_n13121_), .ZN(new_n13140_));
  NOR2_X1    g12884(.A1(new_n13140_), .A2(new_n13137_), .ZN(new_n13141_));
  INV_X1     g12885(.I(new_n13100_), .ZN(new_n13142_));
  NAND2_X1   g12886(.A1(new_n13142_), .A2(new_n13109_), .ZN(new_n13143_));
  INV_X1     g12887(.I(new_n13143_), .ZN(new_n13144_));
  NOR2_X1    g12888(.A1(new_n13142_), .A2(new_n13109_), .ZN(new_n13145_));
  INV_X1     g12889(.I(new_n13145_), .ZN(new_n13146_));
  XOR2_X1    g12890(.A1(new_n13099_), .A2(new_n13114_), .Z(new_n13147_));
  AOI21_X1   g12891(.A1(new_n13147_), .A2(new_n13146_), .B(new_n13144_), .ZN(new_n13148_));
  AOI21_X1   g12892(.A1(new_n12841_), .A2(new_n13089_), .B(new_n13091_), .ZN(new_n13149_));
  INV_X1     g12893(.I(new_n13149_), .ZN(new_n13150_));
  OAI22_X1   g12894(.A1(new_n610_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n612_), .ZN(new_n13151_));
  AOI21_X1   g12895(.A1(\b[57] ), .A2(new_n826_), .B(new_n13151_), .ZN(new_n13152_));
  OAI21_X1   g12896(.A1(new_n12203_), .A2(new_n624_), .B(new_n13152_), .ZN(new_n13153_));
  XOR2_X1    g12897(.A1(new_n13153_), .A2(\a[8] ), .Z(new_n13154_));
  OAI22_X1   g12898(.A1(new_n713_), .A2(new_n10308_), .B1(new_n9972_), .B2(new_n717_), .ZN(new_n13155_));
  AOI21_X1   g12899(.A1(\b[54] ), .A2(new_n1126_), .B(new_n13155_), .ZN(new_n13156_));
  OAI21_X1   g12900(.A1(new_n10319_), .A2(new_n986_), .B(new_n13156_), .ZN(new_n13157_));
  XOR2_X1    g12901(.A1(new_n13157_), .A2(\a[11] ), .Z(new_n13158_));
  NOR2_X1    g12902(.A1(new_n13154_), .A2(new_n13158_), .ZN(new_n13159_));
  NAND2_X1   g12903(.A1(new_n13154_), .A2(new_n13158_), .ZN(new_n13160_));
  INV_X1     g12904(.I(new_n13160_), .ZN(new_n13161_));
  NOR2_X1    g12905(.A1(new_n13161_), .A2(new_n13159_), .ZN(new_n13162_));
  INV_X1     g12906(.I(new_n13162_), .ZN(new_n13163_));
  AOI22_X1   g12907(.A1(new_n1738_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n1743_), .ZN(new_n13164_));
  OAI21_X1   g12908(.A1(new_n7096_), .A2(new_n1931_), .B(new_n13164_), .ZN(new_n13165_));
  AOI21_X1   g12909(.A1(new_n7649_), .A2(new_n1746_), .B(new_n13165_), .ZN(new_n13166_));
  XOR2_X1    g12910(.A1(new_n13166_), .A2(new_n1736_), .Z(new_n13167_));
  INV_X1     g12911(.I(new_n13167_), .ZN(new_n13168_));
  NAND2_X1   g12912(.A1(new_n13042_), .A2(new_n12862_), .ZN(new_n13169_));
  NAND2_X1   g12913(.A1(new_n13169_), .A2(new_n13043_), .ZN(new_n13170_));
  AOI22_X1   g12914(.A1(new_n2202_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n2205_), .ZN(new_n13171_));
  OAI21_X1   g12915(.A1(new_n6490_), .A2(new_n2370_), .B(new_n13171_), .ZN(new_n13172_));
  AOI21_X1   g12916(.A1(new_n7906_), .A2(new_n2208_), .B(new_n13172_), .ZN(new_n13173_));
  XOR2_X1    g12917(.A1(new_n13173_), .A2(new_n2200_), .Z(new_n13174_));
  INV_X1     g12918(.I(new_n13174_), .ZN(new_n13175_));
  INV_X1     g12919(.I(new_n12872_), .ZN(new_n13176_));
  OAI21_X1   g12920(.A1(new_n12864_), .A2(new_n12720_), .B(new_n13176_), .ZN(new_n13177_));
  NOR3_X1    g12921(.A1(new_n12864_), .A2(new_n12720_), .A3(new_n13176_), .ZN(new_n13178_));
  INV_X1     g12922(.I(new_n12865_), .ZN(new_n13179_));
  XOR2_X1    g12923(.A1(new_n13025_), .A2(new_n13179_), .Z(new_n13180_));
  OR2_X2     g12924(.A1(new_n13178_), .A2(new_n13180_), .Z(new_n13181_));
  OAI22_X1   g12925(.A1(new_n2703_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n2708_), .ZN(new_n13182_));
  AOI21_X1   g12926(.A1(\b[39] ), .A2(new_n2906_), .B(new_n13182_), .ZN(new_n13183_));
  OAI21_X1   g12927(.A1(new_n6299_), .A2(new_n2711_), .B(new_n13183_), .ZN(new_n13184_));
  XOR2_X1    g12928(.A1(new_n13184_), .A2(\a[26] ), .Z(new_n13185_));
  AOI22_X1   g12929(.A1(new_n3267_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n3270_), .ZN(new_n13186_));
  OAI21_X1   g12930(.A1(new_n4886_), .A2(new_n3475_), .B(new_n13186_), .ZN(new_n13187_));
  AOI21_X1   g12931(.A1(new_n5351_), .A2(new_n3273_), .B(new_n13187_), .ZN(new_n13188_));
  XOR2_X1    g12932(.A1(new_n13188_), .A2(new_n3264_), .Z(new_n13189_));
  NAND3_X1   g12933(.A1(new_n13010_), .A2(new_n12877_), .A3(new_n13014_), .ZN(new_n13190_));
  NAND2_X1   g12934(.A1(new_n13190_), .A2(new_n13012_), .ZN(new_n13191_));
  NAND2_X1   g12935(.A1(new_n13006_), .A2(new_n13004_), .ZN(new_n13192_));
  INV_X1     g12936(.I(new_n12991_), .ZN(new_n13193_));
  OAI21_X1   g12937(.A1(new_n12883_), .A2(new_n12671_), .B(new_n13193_), .ZN(new_n13194_));
  NAND3_X1   g12938(.A1(new_n12888_), .A2(new_n12887_), .A3(new_n12991_), .ZN(new_n13195_));
  XOR2_X1    g12939(.A1(new_n12987_), .A2(new_n12884_), .Z(new_n13196_));
  NAND2_X1   g12940(.A1(new_n13195_), .A2(new_n13196_), .ZN(new_n13197_));
  NOR2_X1    g12941(.A1(new_n12885_), .A2(new_n12895_), .ZN(new_n13198_));
  XOR2_X1    g12942(.A1(new_n12980_), .A2(new_n12891_), .Z(new_n13199_));
  AOI21_X1   g12943(.A1(new_n12885_), .A2(new_n12895_), .B(new_n13199_), .ZN(new_n13200_));
  NOR2_X1    g12944(.A1(new_n13200_), .A2(new_n13198_), .ZN(new_n13201_));
  AOI21_X1   g12945(.A1(new_n12976_), .A2(new_n12969_), .B(new_n12971_), .ZN(new_n13202_));
  INV_X1     g12946(.I(new_n13202_), .ZN(new_n13203_));
  NAND2_X1   g12947(.A1(new_n12891_), .A2(new_n12974_), .ZN(new_n13204_));
  NAND3_X1   g12948(.A1(new_n13204_), .A2(new_n12979_), .A3(new_n13203_), .ZN(new_n13205_));
  INV_X1     g12949(.I(new_n12979_), .ZN(new_n13206_));
  NOR2_X1    g12950(.A1(new_n12977_), .A2(new_n12978_), .ZN(new_n13207_));
  AOI22_X1   g12951(.A1(new_n13207_), .A2(new_n12899_), .B1(new_n12645_), .B2(new_n12890_), .ZN(new_n13208_));
  OAI21_X1   g12952(.A1(new_n13208_), .A2(new_n13206_), .B(new_n13202_), .ZN(new_n13209_));
  INV_X1     g12953(.I(new_n12912_), .ZN(new_n13210_));
  NAND2_X1   g12954(.A1(new_n12903_), .A2(new_n13210_), .ZN(new_n13211_));
  XNOR2_X1   g12955(.A1(new_n12956_), .A2(new_n12905_), .ZN(new_n13212_));
  OAI21_X1   g12956(.A1(new_n12903_), .A2(new_n13210_), .B(new_n13212_), .ZN(new_n13213_));
  NAND2_X1   g12957(.A1(new_n13213_), .A2(new_n13211_), .ZN(new_n13214_));
  NOR2_X1    g12958(.A1(new_n12905_), .A2(new_n12955_), .ZN(new_n13215_));
  NOR2_X1    g12959(.A1(new_n13215_), .A2(new_n12954_), .ZN(new_n13216_));
  NAND2_X1   g12960(.A1(new_n12914_), .A2(new_n12947_), .ZN(new_n13217_));
  AND2_X2    g12961(.A1(new_n13217_), .A2(new_n12945_), .Z(new_n13218_));
  NAND2_X1   g12962(.A1(new_n12915_), .A2(new_n12937_), .ZN(new_n13219_));
  NAND2_X1   g12963(.A1(new_n13219_), .A2(new_n12936_), .ZN(new_n13220_));
  NOR2_X1    g12964(.A1(new_n12917_), .A2(new_n12928_), .ZN(new_n13221_));
  NOR2_X1    g12965(.A1(new_n13221_), .A2(new_n12926_), .ZN(new_n13222_));
  INV_X1     g12966(.I(new_n12317_), .ZN(new_n13223_));
  INV_X1     g12967(.I(new_n11926_), .ZN(new_n13224_));
  OAI22_X1   g12968(.A1(new_n13224_), .A2(new_n377_), .B1(new_n339_), .B2(new_n11923_), .ZN(new_n13225_));
  AOI21_X1   g12969(.A1(\b[3] ), .A2(new_n13223_), .B(new_n13225_), .ZN(new_n13226_));
  OAI21_X1   g12970(.A1(new_n566_), .A2(new_n11930_), .B(new_n13226_), .ZN(new_n13227_));
  XOR2_X1    g12971(.A1(new_n13227_), .A2(\a[62] ), .Z(new_n13228_));
  AOI22_X1   g12972(.A1(new_n12922_), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n12923_), .ZN(new_n13229_));
  INV_X1     g12973(.I(new_n13229_), .ZN(new_n13230_));
  NOR2_X1    g12974(.A1(new_n13228_), .A2(new_n13230_), .ZN(new_n13231_));
  INV_X1     g12975(.I(new_n13231_), .ZN(new_n13232_));
  NAND2_X1   g12976(.A1(new_n13228_), .A2(new_n13230_), .ZN(new_n13233_));
  NAND2_X1   g12977(.A1(new_n13232_), .A2(new_n13233_), .ZN(new_n13234_));
  XOR2_X1    g12978(.A1(new_n13222_), .A2(new_n13234_), .Z(new_n13235_));
  INV_X1     g12979(.I(new_n13235_), .ZN(new_n13236_));
  AOI22_X1   g12980(.A1(new_n10981_), .A2(\b[8] ), .B1(new_n10979_), .B2(\b[7] ), .ZN(new_n13237_));
  OAI21_X1   g12981(.A1(new_n438_), .A2(new_n11306_), .B(new_n13237_), .ZN(new_n13238_));
  AOI21_X1   g12982(.A1(new_n799_), .A2(new_n10984_), .B(new_n13238_), .ZN(new_n13239_));
  XOR2_X1    g12983(.A1(new_n13239_), .A2(new_n10989_), .Z(new_n13240_));
  NOR2_X1    g12984(.A1(new_n13236_), .A2(new_n13240_), .ZN(new_n13241_));
  INV_X1     g12985(.I(new_n13241_), .ZN(new_n13242_));
  NAND2_X1   g12986(.A1(new_n13236_), .A2(new_n13240_), .ZN(new_n13243_));
  NAND2_X1   g12987(.A1(new_n13242_), .A2(new_n13243_), .ZN(new_n13244_));
  XNOR2_X1   g12988(.A1(new_n13244_), .A2(new_n13220_), .ZN(new_n13245_));
  OAI22_X1   g12989(.A1(new_n11298_), .A2(new_n852_), .B1(new_n776_), .B2(new_n11297_), .ZN(new_n13246_));
  AOI21_X1   g12990(.A1(\b[9] ), .A2(new_n11296_), .B(new_n13246_), .ZN(new_n13247_));
  OAI21_X1   g12991(.A1(new_n859_), .A2(new_n10069_), .B(new_n13247_), .ZN(new_n13248_));
  XOR2_X1    g12992(.A1(new_n13248_), .A2(\a[56] ), .Z(new_n13249_));
  INV_X1     g12993(.I(new_n13249_), .ZN(new_n13250_));
  NAND2_X1   g12994(.A1(new_n13245_), .A2(new_n13250_), .ZN(new_n13251_));
  OR2_X2     g12995(.A1(new_n13245_), .A2(new_n13250_), .Z(new_n13252_));
  NAND2_X1   g12996(.A1(new_n13252_), .A2(new_n13251_), .ZN(new_n13253_));
  XOR2_X1    g12997(.A1(new_n13218_), .A2(new_n13253_), .Z(new_n13254_));
  AOI22_X1   g12998(.A1(new_n9125_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n9123_), .ZN(new_n13255_));
  OAI21_X1   g12999(.A1(new_n941_), .A2(new_n9470_), .B(new_n13255_), .ZN(new_n13256_));
  AOI21_X1   g13000(.A1(new_n1449_), .A2(new_n9129_), .B(new_n13256_), .ZN(new_n13257_));
  XOR2_X1    g13001(.A1(new_n13257_), .A2(new_n9133_), .Z(new_n13258_));
  INV_X1     g13002(.I(new_n13258_), .ZN(new_n13259_));
  NAND2_X1   g13003(.A1(new_n13254_), .A2(new_n13259_), .ZN(new_n13260_));
  OR2_X2     g13004(.A1(new_n13254_), .A2(new_n13259_), .Z(new_n13261_));
  NAND2_X1   g13005(.A1(new_n13261_), .A2(new_n13260_), .ZN(new_n13262_));
  XNOR2_X1   g13006(.A1(new_n13262_), .A2(new_n13216_), .ZN(new_n13263_));
  OAI22_X1   g13007(.A1(new_n9461_), .A2(new_n1432_), .B1(new_n1296_), .B2(new_n9462_), .ZN(new_n13264_));
  AOI21_X1   g13008(.A1(\b[15] ), .A2(new_n8575_), .B(new_n13264_), .ZN(new_n13265_));
  OAI21_X1   g13009(.A1(new_n1444_), .A2(new_n9460_), .B(new_n13265_), .ZN(new_n13266_));
  XOR2_X1    g13010(.A1(new_n13266_), .A2(\a[50] ), .Z(new_n13267_));
  XOR2_X1    g13011(.A1(new_n13263_), .A2(new_n13267_), .Z(new_n13268_));
  XOR2_X1    g13012(.A1(new_n13268_), .A2(new_n13214_), .Z(new_n13269_));
  AOI22_X1   g13013(.A1(new_n7403_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n7408_), .ZN(new_n13270_));
  OAI21_X1   g13014(.A1(new_n1553_), .A2(new_n9488_), .B(new_n13270_), .ZN(new_n13271_));
  AOI21_X1   g13015(.A1(new_n2452_), .A2(new_n7414_), .B(new_n13271_), .ZN(new_n13272_));
  XOR2_X1    g13016(.A1(new_n13272_), .A2(new_n7410_), .Z(new_n13273_));
  INV_X1     g13017(.I(new_n13273_), .ZN(new_n13274_));
  NAND2_X1   g13018(.A1(new_n13269_), .A2(new_n13274_), .ZN(new_n13275_));
  NOR2_X1    g13019(.A1(new_n13269_), .A2(new_n13274_), .ZN(new_n13276_));
  INV_X1     g13020(.I(new_n13276_), .ZN(new_n13277_));
  AOI22_X1   g13021(.A1(new_n6569_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n6574_), .ZN(new_n13278_));
  OAI21_X1   g13022(.A1(new_n2027_), .A2(new_n8565_), .B(new_n13278_), .ZN(new_n13279_));
  AOI21_X1   g13023(.A1(new_n2470_), .A2(new_n6579_), .B(new_n13279_), .ZN(new_n13280_));
  XOR2_X1    g13024(.A1(new_n13280_), .A2(new_n6567_), .Z(new_n13281_));
  AOI21_X1   g13025(.A1(new_n13277_), .A2(new_n13275_), .B(new_n13281_), .ZN(new_n13282_));
  NAND3_X1   g13026(.A1(new_n13277_), .A2(new_n13275_), .A3(new_n13281_), .ZN(new_n13283_));
  INV_X1     g13027(.I(new_n13283_), .ZN(new_n13284_));
  NOR2_X1    g13028(.A1(new_n13284_), .A2(new_n13282_), .ZN(new_n13285_));
  NAND3_X1   g13029(.A1(new_n13285_), .A2(new_n13209_), .A3(new_n13205_), .ZN(new_n13286_));
  NOR3_X1    g13030(.A1(new_n13208_), .A2(new_n13202_), .A3(new_n13206_), .ZN(new_n13287_));
  AOI21_X1   g13031(.A1(new_n13204_), .A2(new_n12979_), .B(new_n13203_), .ZN(new_n13288_));
  INV_X1     g13032(.I(new_n13282_), .ZN(new_n13289_));
  NAND2_X1   g13033(.A1(new_n13289_), .A2(new_n13283_), .ZN(new_n13290_));
  OAI21_X1   g13034(.A1(new_n13287_), .A2(new_n13288_), .B(new_n13290_), .ZN(new_n13291_));
  AOI22_X1   g13035(.A1(new_n6108_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n6111_), .ZN(new_n13292_));
  OAI21_X1   g13036(.A1(new_n2495_), .A2(new_n7708_), .B(new_n13292_), .ZN(new_n13293_));
  AOI21_X1   g13037(.A1(new_n3407_), .A2(new_n6105_), .B(new_n13293_), .ZN(new_n13294_));
  XOR2_X1    g13038(.A1(new_n13294_), .A2(new_n5849_), .Z(new_n13295_));
  INV_X1     g13039(.I(new_n13295_), .ZN(new_n13296_));
  NAND3_X1   g13040(.A1(new_n13291_), .A2(new_n13286_), .A3(new_n13296_), .ZN(new_n13297_));
  NOR3_X1    g13041(.A1(new_n13290_), .A2(new_n13287_), .A3(new_n13288_), .ZN(new_n13298_));
  AOI21_X1   g13042(.A1(new_n13209_), .A2(new_n13205_), .B(new_n13285_), .ZN(new_n13299_));
  OAI21_X1   g13043(.A1(new_n13299_), .A2(new_n13298_), .B(new_n13295_), .ZN(new_n13300_));
  NAND2_X1   g13044(.A1(new_n13300_), .A2(new_n13297_), .ZN(new_n13301_));
  NAND2_X1   g13045(.A1(new_n13201_), .A2(new_n13301_), .ZN(new_n13302_));
  NOR3_X1    g13046(.A1(new_n13299_), .A2(new_n13298_), .A3(new_n13295_), .ZN(new_n13303_));
  AOI21_X1   g13047(.A1(new_n13291_), .A2(new_n13286_), .B(new_n13296_), .ZN(new_n13304_));
  NOR2_X1    g13048(.A1(new_n13303_), .A2(new_n13304_), .ZN(new_n13305_));
  OAI21_X1   g13049(.A1(new_n13198_), .A2(new_n13200_), .B(new_n13305_), .ZN(new_n13306_));
  AOI22_X1   g13050(.A1(new_n5155_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n5160_), .ZN(new_n13307_));
  OAI21_X1   g13051(.A1(new_n3158_), .A2(new_n6877_), .B(new_n13307_), .ZN(new_n13308_));
  AOI21_X1   g13052(.A1(new_n4188_), .A2(new_n5166_), .B(new_n13308_), .ZN(new_n13309_));
  XOR2_X1    g13053(.A1(new_n13309_), .A2(new_n5162_), .Z(new_n13310_));
  INV_X1     g13054(.I(new_n13310_), .ZN(new_n13311_));
  NAND3_X1   g13055(.A1(new_n13306_), .A2(new_n13302_), .A3(new_n13311_), .ZN(new_n13312_));
  NOR3_X1    g13056(.A1(new_n13305_), .A2(new_n13198_), .A3(new_n13200_), .ZN(new_n13313_));
  NOR2_X1    g13057(.A1(new_n13201_), .A2(new_n13301_), .ZN(new_n13314_));
  OAI21_X1   g13058(.A1(new_n13314_), .A2(new_n13313_), .B(new_n13310_), .ZN(new_n13315_));
  NAND2_X1   g13059(.A1(new_n13312_), .A2(new_n13315_), .ZN(new_n13316_));
  AOI21_X1   g13060(.A1(new_n13194_), .A2(new_n13197_), .B(new_n13316_), .ZN(new_n13317_));
  NAND2_X1   g13061(.A1(new_n13197_), .A2(new_n13194_), .ZN(new_n13318_));
  NOR3_X1    g13062(.A1(new_n13314_), .A2(new_n13313_), .A3(new_n13310_), .ZN(new_n13319_));
  AOI21_X1   g13063(.A1(new_n13306_), .A2(new_n13302_), .B(new_n13311_), .ZN(new_n13320_));
  NOR2_X1    g13064(.A1(new_n13320_), .A2(new_n13319_), .ZN(new_n13321_));
  NOR2_X1    g13065(.A1(new_n13318_), .A2(new_n13321_), .ZN(new_n13322_));
  AOI22_X1   g13066(.A1(new_n4918_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n4921_), .ZN(new_n13323_));
  OAI21_X1   g13067(.A1(new_n3624_), .A2(new_n6099_), .B(new_n13323_), .ZN(new_n13324_));
  AOI21_X1   g13068(.A1(new_n4030_), .A2(new_n4699_), .B(new_n13324_), .ZN(new_n13325_));
  XOR2_X1    g13069(.A1(new_n13325_), .A2(new_n4446_), .Z(new_n13326_));
  NOR3_X1    g13070(.A1(new_n13317_), .A2(new_n13322_), .A3(new_n13326_), .ZN(new_n13327_));
  NAND2_X1   g13071(.A1(new_n13318_), .A2(new_n13321_), .ZN(new_n13328_));
  NAND3_X1   g13072(.A1(new_n13316_), .A2(new_n13197_), .A3(new_n13194_), .ZN(new_n13329_));
  INV_X1     g13073(.I(new_n13326_), .ZN(new_n13330_));
  AOI21_X1   g13074(.A1(new_n13328_), .A2(new_n13329_), .B(new_n13330_), .ZN(new_n13331_));
  NOR2_X1    g13075(.A1(new_n13327_), .A2(new_n13331_), .ZN(new_n13332_));
  AOI21_X1   g13076(.A1(new_n13002_), .A2(new_n13192_), .B(new_n13332_), .ZN(new_n13333_));
  AOI21_X1   g13077(.A1(new_n12882_), .A2(new_n12683_), .B(new_n13008_), .ZN(new_n13334_));
  NAND3_X1   g13078(.A1(new_n13328_), .A2(new_n13329_), .A3(new_n13330_), .ZN(new_n13335_));
  OAI21_X1   g13079(.A1(new_n13317_), .A2(new_n13322_), .B(new_n13326_), .ZN(new_n13336_));
  NAND2_X1   g13080(.A1(new_n13336_), .A2(new_n13335_), .ZN(new_n13337_));
  NOR3_X1    g13081(.A1(new_n13337_), .A2(new_n13334_), .A3(new_n13007_), .ZN(new_n13338_));
  OAI22_X1   g13082(.A1(new_n4639_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n4666_), .ZN(new_n13339_));
  AOI21_X1   g13083(.A1(\b[33] ), .A2(new_n4053_), .B(new_n13339_), .ZN(new_n13340_));
  OAI21_X1   g13084(.A1(new_n4676_), .A2(new_n4727_), .B(new_n13340_), .ZN(new_n13341_));
  XOR2_X1    g13085(.A1(new_n13341_), .A2(\a[32] ), .Z(new_n13342_));
  INV_X1     g13086(.I(new_n13342_), .ZN(new_n13343_));
  NOR3_X1    g13087(.A1(new_n13333_), .A2(new_n13338_), .A3(new_n13343_), .ZN(new_n13344_));
  OAI21_X1   g13088(.A1(new_n13007_), .A2(new_n13334_), .B(new_n13337_), .ZN(new_n13345_));
  NAND3_X1   g13089(.A1(new_n13192_), .A2(new_n13332_), .A3(new_n13002_), .ZN(new_n13346_));
  AOI21_X1   g13090(.A1(new_n13345_), .A2(new_n13346_), .B(new_n13342_), .ZN(new_n13347_));
  NOR2_X1    g13091(.A1(new_n13344_), .A2(new_n13347_), .ZN(new_n13348_));
  NOR2_X1    g13092(.A1(new_n13348_), .A2(new_n13191_), .ZN(new_n13349_));
  NAND3_X1   g13093(.A1(new_n13345_), .A2(new_n13346_), .A3(new_n13342_), .ZN(new_n13350_));
  OAI21_X1   g13094(.A1(new_n13333_), .A2(new_n13338_), .B(new_n13343_), .ZN(new_n13351_));
  NAND2_X1   g13095(.A1(new_n13351_), .A2(new_n13350_), .ZN(new_n13352_));
  AOI21_X1   g13096(.A1(new_n13190_), .A2(new_n13012_), .B(new_n13352_), .ZN(new_n13353_));
  NOR3_X1    g13097(.A1(new_n13353_), .A2(new_n13349_), .A3(new_n13189_), .ZN(new_n13354_));
  INV_X1     g13098(.I(new_n13189_), .ZN(new_n13355_));
  NAND3_X1   g13099(.A1(new_n13352_), .A2(new_n13012_), .A3(new_n13190_), .ZN(new_n13356_));
  NAND2_X1   g13100(.A1(new_n13348_), .A2(new_n13191_), .ZN(new_n13357_));
  AOI21_X1   g13101(.A1(new_n13357_), .A2(new_n13356_), .B(new_n13355_), .ZN(new_n13358_));
  NOR2_X1    g13102(.A1(new_n13354_), .A2(new_n13358_), .ZN(new_n13359_));
  NAND2_X1   g13103(.A1(new_n13179_), .A2(new_n13020_), .ZN(new_n13360_));
  NAND3_X1   g13104(.A1(new_n13360_), .A2(new_n13359_), .A3(new_n13024_), .ZN(new_n13361_));
  INV_X1     g13105(.I(new_n13024_), .ZN(new_n13362_));
  NAND3_X1   g13106(.A1(new_n13357_), .A2(new_n13356_), .A3(new_n13355_), .ZN(new_n13363_));
  OAI21_X1   g13107(.A1(new_n13353_), .A2(new_n13349_), .B(new_n13189_), .ZN(new_n13364_));
  NAND2_X1   g13108(.A1(new_n13364_), .A2(new_n13363_), .ZN(new_n13365_));
  NOR2_X1    g13109(.A1(new_n13023_), .A2(new_n13022_), .ZN(new_n13366_));
  AOI21_X1   g13110(.A1(new_n13366_), .A2(new_n12876_), .B(new_n12865_), .ZN(new_n13367_));
  OAI21_X1   g13111(.A1(new_n13367_), .A2(new_n13362_), .B(new_n13365_), .ZN(new_n13368_));
  NAND3_X1   g13112(.A1(new_n13368_), .A2(new_n13361_), .A3(new_n13185_), .ZN(new_n13369_));
  INV_X1     g13113(.I(new_n13185_), .ZN(new_n13370_));
  NOR3_X1    g13114(.A1(new_n13365_), .A2(new_n13367_), .A3(new_n13362_), .ZN(new_n13371_));
  AOI21_X1   g13115(.A1(new_n13360_), .A2(new_n13024_), .B(new_n13359_), .ZN(new_n13372_));
  OAI21_X1   g13116(.A1(new_n13372_), .A2(new_n13371_), .B(new_n13370_), .ZN(new_n13373_));
  NAND2_X1   g13117(.A1(new_n13373_), .A2(new_n13369_), .ZN(new_n13374_));
  AOI21_X1   g13118(.A1(new_n13181_), .A2(new_n13177_), .B(new_n13374_), .ZN(new_n13375_));
  INV_X1     g13119(.I(new_n13177_), .ZN(new_n13376_));
  NOR2_X1    g13120(.A1(new_n13178_), .A2(new_n13180_), .ZN(new_n13377_));
  NOR3_X1    g13121(.A1(new_n13372_), .A2(new_n13371_), .A3(new_n13370_), .ZN(new_n13378_));
  AOI21_X1   g13122(.A1(new_n13368_), .A2(new_n13361_), .B(new_n13185_), .ZN(new_n13379_));
  NOR2_X1    g13123(.A1(new_n13379_), .A2(new_n13378_), .ZN(new_n13380_));
  NOR3_X1    g13124(.A1(new_n13380_), .A2(new_n13377_), .A3(new_n13376_), .ZN(new_n13381_));
  NOR3_X1    g13125(.A1(new_n13375_), .A2(new_n13175_), .A3(new_n13381_), .ZN(new_n13382_));
  OAI21_X1   g13126(.A1(new_n13377_), .A2(new_n13376_), .B(new_n13380_), .ZN(new_n13383_));
  NAND3_X1   g13127(.A1(new_n13181_), .A2(new_n13177_), .A3(new_n13374_), .ZN(new_n13384_));
  AOI21_X1   g13128(.A1(new_n13384_), .A2(new_n13383_), .B(new_n13174_), .ZN(new_n13385_));
  NOR2_X1    g13129(.A1(new_n13382_), .A2(new_n13385_), .ZN(new_n13386_));
  NAND2_X1   g13130(.A1(new_n13170_), .A2(new_n13386_), .ZN(new_n13387_));
  NAND3_X1   g13131(.A1(new_n13384_), .A2(new_n13383_), .A3(new_n13174_), .ZN(new_n13388_));
  OAI21_X1   g13132(.A1(new_n13375_), .A2(new_n13381_), .B(new_n13175_), .ZN(new_n13389_));
  NAND2_X1   g13133(.A1(new_n13389_), .A2(new_n13388_), .ZN(new_n13390_));
  NAND3_X1   g13134(.A1(new_n13390_), .A2(new_n13043_), .A3(new_n13169_), .ZN(new_n13391_));
  NAND3_X1   g13135(.A1(new_n13387_), .A2(new_n13391_), .A3(new_n13168_), .ZN(new_n13392_));
  AOI21_X1   g13136(.A1(new_n13169_), .A2(new_n13043_), .B(new_n13390_), .ZN(new_n13393_));
  NOR2_X1    g13137(.A1(new_n13170_), .A2(new_n13386_), .ZN(new_n13394_));
  OAI21_X1   g13138(.A1(new_n13393_), .A2(new_n13394_), .B(new_n13167_), .ZN(new_n13395_));
  NAND2_X1   g13139(.A1(new_n13395_), .A2(new_n13392_), .ZN(new_n13396_));
  AOI21_X1   g13140(.A1(new_n13041_), .A2(new_n13045_), .B(new_n13047_), .ZN(new_n13397_));
  AOI21_X1   g13141(.A1(new_n13051_), .A2(new_n12857_), .B(new_n13397_), .ZN(new_n13398_));
  NOR2_X1    g13142(.A1(new_n13398_), .A2(new_n13396_), .ZN(new_n13399_));
  NOR3_X1    g13143(.A1(new_n13393_), .A2(new_n13394_), .A3(new_n13167_), .ZN(new_n13400_));
  AOI21_X1   g13144(.A1(new_n13387_), .A2(new_n13391_), .B(new_n13168_), .ZN(new_n13401_));
  NOR2_X1    g13145(.A1(new_n13400_), .A2(new_n13401_), .ZN(new_n13402_));
  NOR3_X1    g13146(.A1(new_n13060_), .A2(new_n13402_), .A3(new_n13397_), .ZN(new_n13403_));
  OAI22_X1   g13147(.A1(new_n1592_), .A2(new_n8500_), .B1(new_n8168_), .B2(new_n1505_), .ZN(new_n13404_));
  AOI21_X1   g13148(.A1(\b[48] ), .A2(new_n1584_), .B(new_n13404_), .ZN(new_n13405_));
  OAI21_X1   g13149(.A1(new_n8510_), .A2(new_n1732_), .B(new_n13405_), .ZN(new_n13406_));
  XOR2_X1    g13150(.A1(new_n13406_), .A2(\a[17] ), .Z(new_n13407_));
  INV_X1     g13151(.I(new_n13407_), .ZN(new_n13408_));
  OAI21_X1   g13152(.A1(new_n13403_), .A2(new_n13399_), .B(new_n13408_), .ZN(new_n13409_));
  OAI21_X1   g13153(.A1(new_n13060_), .A2(new_n13397_), .B(new_n13402_), .ZN(new_n13410_));
  NAND2_X1   g13154(.A1(new_n13398_), .A2(new_n13396_), .ZN(new_n13411_));
  NAND3_X1   g13155(.A1(new_n13410_), .A2(new_n13411_), .A3(new_n13407_), .ZN(new_n13412_));
  NAND4_X1   g13156(.A1(new_n13063_), .A2(new_n13412_), .A3(new_n13409_), .A4(new_n13058_), .ZN(new_n13413_));
  AOI21_X1   g13157(.A1(new_n13410_), .A2(new_n13411_), .B(new_n13407_), .ZN(new_n13414_));
  NOR3_X1    g13158(.A1(new_n13403_), .A2(new_n13399_), .A3(new_n13408_), .ZN(new_n13415_));
  OAI22_X1   g13159(.A1(new_n13070_), .A2(new_n13065_), .B1(new_n13414_), .B2(new_n13415_), .ZN(new_n13416_));
  OAI22_X1   g13160(.A1(new_n993_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n997_), .ZN(new_n13417_));
  AOI21_X1   g13161(.A1(\b[51] ), .A2(new_n1486_), .B(new_n13417_), .ZN(new_n13418_));
  OAI21_X1   g13162(.A1(new_n9385_), .A2(new_n1323_), .B(new_n13418_), .ZN(new_n13419_));
  XOR2_X1    g13163(.A1(new_n13419_), .A2(\a[14] ), .Z(new_n13420_));
  INV_X1     g13164(.I(new_n13420_), .ZN(new_n13421_));
  NAND3_X1   g13165(.A1(new_n13416_), .A2(new_n13413_), .A3(new_n13421_), .ZN(new_n13422_));
  NOR4_X1    g13166(.A1(new_n13070_), .A2(new_n13414_), .A3(new_n13415_), .A4(new_n13065_), .ZN(new_n13423_));
  AOI22_X1   g13167(.A1(new_n13409_), .A2(new_n13412_), .B1(new_n13063_), .B2(new_n13058_), .ZN(new_n13424_));
  OAI21_X1   g13168(.A1(new_n13423_), .A2(new_n13424_), .B(new_n13420_), .ZN(new_n13425_));
  NAND2_X1   g13169(.A1(new_n13425_), .A2(new_n13422_), .ZN(new_n13426_));
  NOR3_X1    g13170(.A1(new_n12847_), .A2(new_n12770_), .A3(new_n13068_), .ZN(new_n13427_));
  INV_X1     g13171(.I(new_n13427_), .ZN(new_n13428_));
  AOI21_X1   g13172(.A1(new_n13428_), .A2(new_n13077_), .B(new_n13426_), .ZN(new_n13429_));
  NOR3_X1    g13173(.A1(new_n13423_), .A2(new_n13424_), .A3(new_n13420_), .ZN(new_n13430_));
  AOI21_X1   g13174(.A1(new_n13416_), .A2(new_n13413_), .B(new_n13421_), .ZN(new_n13431_));
  NOR2_X1    g13175(.A1(new_n13430_), .A2(new_n13431_), .ZN(new_n13432_));
  NOR3_X1    g13176(.A1(new_n13432_), .A2(new_n13072_), .A3(new_n13427_), .ZN(new_n13433_));
  NOR3_X1    g13177(.A1(new_n13429_), .A2(new_n13433_), .A3(new_n13163_), .ZN(new_n13434_));
  OAI21_X1   g13178(.A1(new_n13072_), .A2(new_n13427_), .B(new_n13432_), .ZN(new_n13435_));
  NAND3_X1   g13179(.A1(new_n13426_), .A2(new_n13428_), .A3(new_n13077_), .ZN(new_n13436_));
  AOI21_X1   g13180(.A1(new_n13435_), .A2(new_n13436_), .B(new_n13162_), .ZN(new_n13437_));
  NOR2_X1    g13181(.A1(new_n13437_), .A2(new_n13434_), .ZN(new_n13438_));
  NOR2_X1    g13182(.A1(new_n13438_), .A2(new_n13150_), .ZN(new_n13439_));
  NAND3_X1   g13183(.A1(new_n13435_), .A2(new_n13162_), .A3(new_n13436_), .ZN(new_n13440_));
  OAI21_X1   g13184(.A1(new_n13429_), .A2(new_n13433_), .B(new_n13163_), .ZN(new_n13441_));
  NAND2_X1   g13185(.A1(new_n13441_), .A2(new_n13440_), .ZN(new_n13442_));
  NOR2_X1    g13186(.A1(new_n13442_), .A2(new_n13149_), .ZN(new_n13443_));
  NAND2_X1   g13187(.A1(new_n12523_), .A2(new_n12519_), .ZN(new_n13444_));
  AOI22_X1   g13188(.A1(new_n800_), .A2(\b[61] ), .B1(\b[62] ), .B2(new_n333_), .ZN(new_n13445_));
  OAI21_X1   g13189(.A1(new_n12147_), .A2(new_n392_), .B(new_n13445_), .ZN(new_n13446_));
  AOI21_X1   g13190(.A1(new_n13444_), .A2(new_n330_), .B(new_n13446_), .ZN(new_n13447_));
  XOR2_X1    g13191(.A1(new_n13447_), .A2(new_n312_), .Z(new_n13448_));
  OAI21_X1   g13192(.A1(new_n13439_), .A2(new_n13443_), .B(new_n13448_), .ZN(new_n13449_));
  NAND2_X1   g13193(.A1(new_n13442_), .A2(new_n13149_), .ZN(new_n13450_));
  NAND2_X1   g13194(.A1(new_n13438_), .A2(new_n13150_), .ZN(new_n13451_));
  INV_X1     g13195(.I(new_n13448_), .ZN(new_n13452_));
  NAND3_X1   g13196(.A1(new_n13451_), .A2(new_n13450_), .A3(new_n13452_), .ZN(new_n13453_));
  NAND2_X1   g13197(.A1(new_n13449_), .A2(new_n13453_), .ZN(new_n13454_));
  NOR2_X1    g13198(.A1(new_n13114_), .A2(new_n12845_), .ZN(new_n13455_));
  OAI21_X1   g13199(.A1(new_n13091_), .A2(new_n13092_), .B(new_n12841_), .ZN(new_n13456_));
  NAND3_X1   g13200(.A1(new_n13095_), .A2(new_n13086_), .A3(new_n13089_), .ZN(new_n13457_));
  AOI22_X1   g13201(.A1(new_n13456_), .A2(new_n13457_), .B1(new_n12845_), .B2(new_n13114_), .ZN(new_n13458_));
  NAND2_X1   g13202(.A1(new_n283_), .A2(\b[63] ), .ZN(new_n13459_));
  AOI21_X1   g13203(.A1(new_n12799_), .A2(new_n12796_), .B(new_n12800_), .ZN(new_n13460_));
  AOI21_X1   g13204(.A1(new_n13460_), .A2(new_n265_), .B(new_n270_), .ZN(new_n13461_));
  INV_X1     g13205(.I(new_n13460_), .ZN(new_n13462_));
  NOR3_X1    g13206(.A1(new_n13462_), .A2(\a[2] ), .A3(new_n279_), .ZN(new_n13463_));
  AOI21_X1   g13207(.A1(new_n13461_), .A2(new_n13459_), .B(new_n13463_), .ZN(new_n13464_));
  OAI21_X1   g13208(.A1(new_n13458_), .A2(new_n13455_), .B(new_n13464_), .ZN(new_n13465_));
  INV_X1     g13209(.I(new_n13465_), .ZN(new_n13466_));
  NOR3_X1    g13210(.A1(new_n13458_), .A2(new_n13455_), .A3(new_n13464_), .ZN(new_n13467_));
  NOR2_X1    g13211(.A1(new_n13466_), .A2(new_n13467_), .ZN(new_n13468_));
  NOR2_X1    g13212(.A1(new_n13468_), .A2(new_n13454_), .ZN(new_n13469_));
  NAND2_X1   g13213(.A1(new_n13468_), .A2(new_n13454_), .ZN(new_n13470_));
  INV_X1     g13214(.I(new_n13470_), .ZN(new_n13471_));
  NOR3_X1    g13215(.A1(new_n13471_), .A2(new_n13148_), .A3(new_n13469_), .ZN(new_n13472_));
  XOR2_X1    g13216(.A1(new_n13099_), .A2(new_n13115_), .Z(new_n13473_));
  OAI21_X1   g13217(.A1(new_n13473_), .A2(new_n13145_), .B(new_n13143_), .ZN(new_n13474_));
  INV_X1     g13218(.I(new_n13469_), .ZN(new_n13475_));
  AOI21_X1   g13219(.A1(new_n13475_), .A2(new_n13470_), .B(new_n13474_), .ZN(new_n13476_));
  NOR2_X1    g13220(.A1(new_n13476_), .A2(new_n13472_), .ZN(new_n13477_));
  XOR2_X1    g13221(.A1(new_n13141_), .A2(new_n13477_), .Z(\f[65] ));
  NAND2_X1   g13222(.A1(new_n13129_), .A2(new_n13128_), .ZN(new_n13479_));
  AOI21_X1   g13223(.A1(new_n13119_), .A2(new_n13102_), .B(new_n13116_), .ZN(new_n13480_));
  NOR3_X1    g13224(.A1(new_n13103_), .A2(new_n13117_), .A3(new_n13101_), .ZN(new_n13481_));
  NOR2_X1    g13225(.A1(new_n13480_), .A2(new_n13481_), .ZN(new_n13482_));
  OAI21_X1   g13226(.A1(new_n13129_), .A2(new_n13128_), .B(new_n13482_), .ZN(new_n13483_));
  AOI21_X1   g13227(.A1(new_n13483_), .A2(new_n13479_), .B(new_n13476_), .ZN(new_n13484_));
  NOR2_X1    g13228(.A1(new_n13484_), .A2(new_n13472_), .ZN(new_n13485_));
  INV_X1     g13229(.I(new_n13467_), .ZN(new_n13486_));
  AOI21_X1   g13230(.A1(new_n13454_), .A2(new_n13486_), .B(new_n13466_), .ZN(new_n13487_));
  NOR2_X1    g13231(.A1(new_n13438_), .A2(new_n13448_), .ZN(new_n13488_));
  NAND2_X1   g13232(.A1(new_n13438_), .A2(new_n13448_), .ZN(new_n13489_));
  AOI21_X1   g13233(.A1(new_n13150_), .A2(new_n13489_), .B(new_n13488_), .ZN(new_n13490_));
  AOI22_X1   g13234(.A1(new_n800_), .A2(\b[62] ), .B1(\b[63] ), .B2(new_n333_), .ZN(new_n13491_));
  OAI21_X1   g13235(.A1(new_n12148_), .A2(new_n392_), .B(new_n13491_), .ZN(new_n13492_));
  AOI21_X1   g13236(.A1(new_n12811_), .A2(new_n330_), .B(new_n13492_), .ZN(new_n13493_));
  XOR2_X1    g13237(.A1(new_n13493_), .A2(new_n312_), .Z(new_n13494_));
  INV_X1     g13238(.I(new_n13494_), .ZN(new_n13495_));
  OAI21_X1   g13239(.A1(new_n13334_), .A2(new_n13007_), .B(new_n13336_), .ZN(new_n13496_));
  NAND2_X1   g13240(.A1(new_n13496_), .A2(new_n13335_), .ZN(new_n13497_));
  AOI21_X1   g13241(.A1(new_n13197_), .A2(new_n13194_), .B(new_n13320_), .ZN(new_n13498_));
  NOR2_X1    g13242(.A1(new_n13498_), .A2(new_n13319_), .ZN(new_n13499_));
  INV_X1     g13243(.I(new_n13499_), .ZN(new_n13500_));
  OAI21_X1   g13244(.A1(new_n13201_), .A2(new_n13304_), .B(new_n13297_), .ZN(new_n13501_));
  INV_X1     g13245(.I(new_n13501_), .ZN(new_n13502_));
  NOR2_X1    g13246(.A1(new_n13208_), .A2(new_n13206_), .ZN(new_n13503_));
  NOR2_X1    g13247(.A1(new_n13503_), .A2(new_n13281_), .ZN(new_n13504_));
  NAND2_X1   g13248(.A1(new_n13503_), .A2(new_n13281_), .ZN(new_n13505_));
  NAND2_X1   g13249(.A1(new_n13277_), .A2(new_n13275_), .ZN(new_n13506_));
  XOR2_X1    g13250(.A1(new_n13506_), .A2(new_n13202_), .Z(new_n13507_));
  AOI21_X1   g13251(.A1(new_n13507_), .A2(new_n13505_), .B(new_n13504_), .ZN(new_n13508_));
  NAND2_X1   g13252(.A1(new_n13203_), .A2(new_n13277_), .ZN(new_n13509_));
  NAND2_X1   g13253(.A1(new_n13509_), .A2(new_n13275_), .ZN(new_n13510_));
  NAND2_X1   g13254(.A1(new_n13263_), .A2(new_n13267_), .ZN(new_n13511_));
  NAND2_X1   g13255(.A1(new_n13214_), .A2(new_n13511_), .ZN(new_n13512_));
  OAI21_X1   g13256(.A1(new_n13263_), .A2(new_n13267_), .B(new_n13512_), .ZN(new_n13513_));
  OAI21_X1   g13257(.A1(new_n12954_), .A2(new_n13215_), .B(new_n13261_), .ZN(new_n13514_));
  NAND2_X1   g13258(.A1(new_n13514_), .A2(new_n13260_), .ZN(new_n13515_));
  INV_X1     g13259(.I(new_n13252_), .ZN(new_n13516_));
  OAI21_X1   g13260(.A1(new_n13218_), .A2(new_n13516_), .B(new_n13251_), .ZN(new_n13517_));
  AOI21_X1   g13261(.A1(new_n13220_), .A2(new_n13243_), .B(new_n13241_), .ZN(new_n13518_));
  INV_X1     g13262(.I(new_n13222_), .ZN(new_n13519_));
  AOI21_X1   g13263(.A1(new_n13519_), .A2(new_n13233_), .B(new_n13231_), .ZN(new_n13520_));
  AOI22_X1   g13264(.A1(new_n11926_), .A2(\b[6] ), .B1(new_n11924_), .B2(\b[5] ), .ZN(new_n13521_));
  OAI21_X1   g13265(.A1(new_n339_), .A2(new_n12317_), .B(new_n13521_), .ZN(new_n13522_));
  AOI21_X1   g13266(.A1(new_n916_), .A2(new_n11929_), .B(new_n13522_), .ZN(new_n13523_));
  XOR2_X1    g13267(.A1(new_n13523_), .A2(\a[62] ), .Z(new_n13524_));
  AOI22_X1   g13268(.A1(new_n12922_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n12923_), .ZN(new_n13525_));
  INV_X1     g13269(.I(new_n13525_), .ZN(new_n13526_));
  NAND2_X1   g13270(.A1(new_n13526_), .A2(\a[2] ), .ZN(new_n13527_));
  NOR2_X1    g13271(.A1(new_n13526_), .A2(\a[2] ), .ZN(new_n13528_));
  INV_X1     g13272(.I(new_n13528_), .ZN(new_n13529_));
  NAND2_X1   g13273(.A1(new_n13529_), .A2(new_n13527_), .ZN(new_n13530_));
  XNOR2_X1   g13274(.A1(new_n13524_), .A2(new_n13530_), .ZN(new_n13531_));
  INV_X1     g13275(.I(new_n13531_), .ZN(new_n13532_));
  AOI22_X1   g13276(.A1(new_n10981_), .A2(\b[9] ), .B1(new_n10979_), .B2(\b[8] ), .ZN(new_n13533_));
  OAI21_X1   g13277(.A1(new_n471_), .A2(new_n11306_), .B(new_n13533_), .ZN(new_n13534_));
  AOI21_X1   g13278(.A1(new_n676_), .A2(new_n10984_), .B(new_n13534_), .ZN(new_n13535_));
  XOR2_X1    g13279(.A1(new_n13535_), .A2(new_n10989_), .Z(new_n13536_));
  NOR2_X1    g13280(.A1(new_n13536_), .A2(new_n13532_), .ZN(new_n13537_));
  NAND2_X1   g13281(.A1(new_n13536_), .A2(new_n13532_), .ZN(new_n13538_));
  INV_X1     g13282(.I(new_n13538_), .ZN(new_n13539_));
  NOR2_X1    g13283(.A1(new_n13539_), .A2(new_n13537_), .ZN(new_n13540_));
  XOR2_X1    g13284(.A1(new_n13520_), .A2(new_n13540_), .Z(new_n13541_));
  AOI22_X1   g13285(.A1(new_n10064_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n10062_), .ZN(new_n13542_));
  OAI21_X1   g13286(.A1(new_n776_), .A2(new_n10399_), .B(new_n13542_), .ZN(new_n13543_));
  AOI21_X1   g13287(.A1(new_n1194_), .A2(new_n10068_), .B(new_n13543_), .ZN(new_n13544_));
  XOR2_X1    g13288(.A1(new_n13544_), .A2(new_n10057_), .Z(new_n13545_));
  NOR2_X1    g13289(.A1(new_n13541_), .A2(new_n13545_), .ZN(new_n13546_));
  NAND2_X1   g13290(.A1(new_n13541_), .A2(new_n13545_), .ZN(new_n13547_));
  INV_X1     g13291(.I(new_n13547_), .ZN(new_n13548_));
  NOR2_X1    g13292(.A1(new_n13548_), .A2(new_n13546_), .ZN(new_n13549_));
  XNOR2_X1   g13293(.A1(new_n13549_), .A2(new_n13518_), .ZN(new_n13550_));
  OAI22_X1   g13294(.A1(new_n10390_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n10389_), .ZN(new_n13551_));
  AOI21_X1   g13295(.A1(\b[13] ), .A2(new_n9471_), .B(new_n13551_), .ZN(new_n13552_));
  OAI21_X1   g13296(.A1(new_n1275_), .A2(new_n10388_), .B(new_n13552_), .ZN(new_n13553_));
  XOR2_X1    g13297(.A1(new_n13553_), .A2(\a[53] ), .Z(new_n13554_));
  INV_X1     g13298(.I(new_n13554_), .ZN(new_n13555_));
  NAND2_X1   g13299(.A1(new_n13550_), .A2(new_n13555_), .ZN(new_n13556_));
  INV_X1     g13300(.I(new_n13556_), .ZN(new_n13557_));
  NOR2_X1    g13301(.A1(new_n13550_), .A2(new_n13555_), .ZN(new_n13558_));
  NOR2_X1    g13302(.A1(new_n13557_), .A2(new_n13558_), .ZN(new_n13559_));
  XNOR2_X1   g13303(.A1(new_n13517_), .A2(new_n13559_), .ZN(new_n13560_));
  AOI22_X1   g13304(.A1(new_n8241_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n8246_), .ZN(new_n13561_));
  OAI21_X1   g13305(.A1(new_n1296_), .A2(new_n9114_), .B(new_n13561_), .ZN(new_n13562_));
  AOI21_X1   g13306(.A1(new_n2038_), .A2(new_n8252_), .B(new_n13562_), .ZN(new_n13563_));
  XOR2_X1    g13307(.A1(new_n13563_), .A2(new_n8248_), .Z(new_n13564_));
  NOR2_X1    g13308(.A1(new_n13560_), .A2(new_n13564_), .ZN(new_n13565_));
  INV_X1     g13309(.I(new_n13565_), .ZN(new_n13566_));
  NAND2_X1   g13310(.A1(new_n13560_), .A2(new_n13564_), .ZN(new_n13567_));
  NAND2_X1   g13311(.A1(new_n13566_), .A2(new_n13567_), .ZN(new_n13568_));
  XOR2_X1    g13312(.A1(new_n13515_), .A2(new_n13568_), .Z(new_n13569_));
  AOI22_X1   g13313(.A1(new_n7403_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n7408_), .ZN(new_n13570_));
  OAI21_X1   g13314(.A1(new_n1859_), .A2(new_n9488_), .B(new_n13570_), .ZN(new_n13571_));
  AOI21_X1   g13315(.A1(new_n2032_), .A2(new_n7414_), .B(new_n13571_), .ZN(new_n13572_));
  XOR2_X1    g13316(.A1(new_n13572_), .A2(new_n7410_), .Z(new_n13573_));
  NOR2_X1    g13317(.A1(new_n13569_), .A2(new_n13573_), .ZN(new_n13574_));
  INV_X1     g13318(.I(new_n13574_), .ZN(new_n13575_));
  NAND2_X1   g13319(.A1(new_n13569_), .A2(new_n13573_), .ZN(new_n13576_));
  NAND2_X1   g13320(.A1(new_n13575_), .A2(new_n13576_), .ZN(new_n13577_));
  XOR2_X1    g13321(.A1(new_n13513_), .A2(new_n13577_), .Z(new_n13578_));
  AOI22_X1   g13322(.A1(new_n6569_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n6574_), .ZN(new_n13579_));
  OAI21_X1   g13323(.A1(new_n2142_), .A2(new_n8565_), .B(new_n13579_), .ZN(new_n13580_));
  AOI21_X1   g13324(.A1(new_n3033_), .A2(new_n6579_), .B(new_n13580_), .ZN(new_n13581_));
  XOR2_X1    g13325(.A1(new_n13581_), .A2(new_n6567_), .Z(new_n13582_));
  OR2_X2     g13326(.A1(new_n13578_), .A2(new_n13582_), .Z(new_n13583_));
  NAND2_X1   g13327(.A1(new_n13578_), .A2(new_n13582_), .ZN(new_n13584_));
  NAND2_X1   g13328(.A1(new_n13583_), .A2(new_n13584_), .ZN(new_n13585_));
  XOR2_X1    g13329(.A1(new_n13585_), .A2(new_n13510_), .Z(new_n13586_));
  OAI22_X1   g13330(.A1(new_n5852_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n5857_), .ZN(new_n13587_));
  AOI21_X1   g13331(.A1(\b[25] ), .A2(new_n6115_), .B(new_n13587_), .ZN(new_n13588_));
  OAI21_X1   g13332(.A1(new_n3165_), .A2(new_n5861_), .B(new_n13588_), .ZN(new_n13589_));
  XOR2_X1    g13333(.A1(new_n13589_), .A2(\a[41] ), .Z(new_n13590_));
  NOR2_X1    g13334(.A1(new_n13586_), .A2(new_n13590_), .ZN(new_n13591_));
  XNOR2_X1   g13335(.A1(new_n13585_), .A2(new_n13510_), .ZN(new_n13592_));
  INV_X1     g13336(.I(new_n13590_), .ZN(new_n13593_));
  NOR2_X1    g13337(.A1(new_n13592_), .A2(new_n13593_), .ZN(new_n13594_));
  NOR2_X1    g13338(.A1(new_n13594_), .A2(new_n13591_), .ZN(new_n13595_));
  XNOR2_X1   g13339(.A1(new_n13595_), .A2(new_n13508_), .ZN(new_n13596_));
  AOI22_X1   g13340(.A1(new_n5155_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n5160_), .ZN(new_n13597_));
  OAI21_X1   g13341(.A1(new_n3185_), .A2(new_n6877_), .B(new_n13597_), .ZN(new_n13598_));
  AOI21_X1   g13342(.A1(new_n4230_), .A2(new_n5166_), .B(new_n13598_), .ZN(new_n13599_));
  XOR2_X1    g13343(.A1(new_n13599_), .A2(new_n5162_), .Z(new_n13600_));
  INV_X1     g13344(.I(new_n13600_), .ZN(new_n13601_));
  NAND2_X1   g13345(.A1(new_n13596_), .A2(new_n13601_), .ZN(new_n13602_));
  XOR2_X1    g13346(.A1(new_n13595_), .A2(new_n13508_), .Z(new_n13603_));
  NAND2_X1   g13347(.A1(new_n13603_), .A2(new_n13600_), .ZN(new_n13604_));
  NAND2_X1   g13348(.A1(new_n13602_), .A2(new_n13604_), .ZN(new_n13605_));
  XOR2_X1    g13349(.A1(new_n13605_), .A2(new_n13502_), .Z(new_n13606_));
  AOI22_X1   g13350(.A1(new_n4918_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n4921_), .ZN(new_n13607_));
  OAI21_X1   g13351(.A1(new_n4022_), .A2(new_n6099_), .B(new_n13607_), .ZN(new_n13608_));
  AOI21_X1   g13352(.A1(new_n4223_), .A2(new_n4699_), .B(new_n13608_), .ZN(new_n13609_));
  XOR2_X1    g13353(.A1(new_n13609_), .A2(new_n4446_), .Z(new_n13610_));
  INV_X1     g13354(.I(new_n13610_), .ZN(new_n13611_));
  NAND2_X1   g13355(.A1(new_n13606_), .A2(new_n13611_), .ZN(new_n13612_));
  OR2_X2     g13356(.A1(new_n13606_), .A2(new_n13611_), .Z(new_n13613_));
  NAND2_X1   g13357(.A1(new_n13613_), .A2(new_n13612_), .ZN(new_n13614_));
  XOR2_X1    g13358(.A1(new_n13614_), .A2(new_n13500_), .Z(new_n13615_));
  AOI22_X1   g13359(.A1(new_n3864_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n3869_), .ZN(new_n13616_));
  OAI21_X1   g13360(.A1(new_n4639_), .A2(new_n5410_), .B(new_n13616_), .ZN(new_n13617_));
  AOI21_X1   g13361(.A1(new_n5594_), .A2(new_n3872_), .B(new_n13617_), .ZN(new_n13618_));
  XOR2_X1    g13362(.A1(new_n13618_), .A2(new_n3876_), .Z(new_n13619_));
  XOR2_X1    g13363(.A1(new_n13615_), .A2(new_n13619_), .Z(new_n13620_));
  XOR2_X1    g13364(.A1(new_n13620_), .A2(new_n13497_), .Z(new_n13621_));
  AOI22_X1   g13365(.A1(new_n3267_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n3270_), .ZN(new_n13622_));
  OAI21_X1   g13366(.A1(new_n5312_), .A2(new_n3475_), .B(new_n13622_), .ZN(new_n13623_));
  AOI21_X1   g13367(.A1(new_n6310_), .A2(new_n3273_), .B(new_n13623_), .ZN(new_n13624_));
  XOR2_X1    g13368(.A1(new_n13624_), .A2(new_n3264_), .Z(new_n13625_));
  INV_X1     g13369(.I(new_n13625_), .ZN(new_n13626_));
  OAI21_X1   g13370(.A1(new_n13191_), .A2(new_n13347_), .B(new_n13350_), .ZN(new_n13627_));
  INV_X1     g13371(.I(new_n13627_), .ZN(new_n13628_));
  NOR2_X1    g13372(.A1(new_n13628_), .A2(new_n13626_), .ZN(new_n13629_));
  NOR2_X1    g13373(.A1(new_n13627_), .A2(new_n13625_), .ZN(new_n13630_));
  NOR2_X1    g13374(.A1(new_n13629_), .A2(new_n13630_), .ZN(new_n13631_));
  XOR2_X1    g13375(.A1(new_n13621_), .A2(new_n13631_), .Z(new_n13632_));
  AOI22_X1   g13376(.A1(new_n2716_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n2719_), .ZN(new_n13633_));
  OAI21_X1   g13377(.A1(new_n6284_), .A2(new_n2924_), .B(new_n13633_), .ZN(new_n13634_));
  AOI21_X1   g13378(.A1(new_n7106_), .A2(new_n2722_), .B(new_n13634_), .ZN(new_n13635_));
  XOR2_X1    g13379(.A1(new_n13635_), .A2(new_n2714_), .Z(new_n13636_));
  NAND2_X1   g13380(.A1(new_n13361_), .A2(new_n13364_), .ZN(new_n13637_));
  NAND2_X1   g13381(.A1(new_n13637_), .A2(new_n13636_), .ZN(new_n13638_));
  NOR2_X1    g13382(.A1(new_n13637_), .A2(new_n13636_), .ZN(new_n13639_));
  INV_X1     g13383(.I(new_n13639_), .ZN(new_n13640_));
  NAND2_X1   g13384(.A1(new_n13640_), .A2(new_n13638_), .ZN(new_n13641_));
  XOR2_X1    g13385(.A1(new_n13632_), .A2(new_n13641_), .Z(new_n13642_));
  AOI22_X1   g13386(.A1(new_n2202_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n2205_), .ZN(new_n13643_));
  OAI21_X1   g13387(.A1(new_n6775_), .A2(new_n2370_), .B(new_n13643_), .ZN(new_n13644_));
  AOI21_X1   g13388(.A1(new_n7926_), .A2(new_n2208_), .B(new_n13644_), .ZN(new_n13645_));
  XOR2_X1    g13389(.A1(new_n13645_), .A2(new_n2200_), .Z(new_n13646_));
  INV_X1     g13390(.I(new_n13646_), .ZN(new_n13647_));
  NOR3_X1    g13391(.A1(new_n13374_), .A2(new_n13377_), .A3(new_n13376_), .ZN(new_n13648_));
  NOR2_X1    g13392(.A1(new_n13648_), .A2(new_n13378_), .ZN(new_n13649_));
  NOR2_X1    g13393(.A1(new_n13649_), .A2(new_n13647_), .ZN(new_n13650_));
  NOR3_X1    g13394(.A1(new_n13648_), .A2(new_n13378_), .A3(new_n13646_), .ZN(new_n13651_));
  NOR2_X1    g13395(.A1(new_n13650_), .A2(new_n13651_), .ZN(new_n13652_));
  XOR2_X1    g13396(.A1(new_n13642_), .A2(new_n13652_), .Z(new_n13653_));
  INV_X1     g13397(.I(new_n13653_), .ZN(new_n13654_));
  AOI22_X1   g13398(.A1(new_n1738_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n1743_), .ZN(new_n13655_));
  OAI21_X1   g13399(.A1(new_n7617_), .A2(new_n1931_), .B(new_n13655_), .ZN(new_n13656_));
  AOI21_X1   g13400(.A1(new_n8792_), .A2(new_n1746_), .B(new_n13656_), .ZN(new_n13657_));
  XOR2_X1    g13401(.A1(new_n13657_), .A2(new_n1736_), .Z(new_n13658_));
  INV_X1     g13402(.I(new_n13658_), .ZN(new_n13659_));
  AOI21_X1   g13403(.A1(new_n13043_), .A2(new_n13169_), .B(new_n13386_), .ZN(new_n13660_));
  AOI21_X1   g13404(.A1(new_n13384_), .A2(new_n13383_), .B(new_n13175_), .ZN(new_n13661_));
  NOR2_X1    g13405(.A1(new_n13660_), .A2(new_n13661_), .ZN(new_n13662_));
  NOR2_X1    g13406(.A1(new_n13662_), .A2(new_n13659_), .ZN(new_n13663_));
  NAND2_X1   g13407(.A1(new_n13662_), .A2(new_n13659_), .ZN(new_n13664_));
  INV_X1     g13408(.I(new_n13664_), .ZN(new_n13665_));
  NOR3_X1    g13409(.A1(new_n13665_), .A2(new_n13654_), .A3(new_n13663_), .ZN(new_n13666_));
  INV_X1     g13410(.I(new_n13663_), .ZN(new_n13667_));
  AOI21_X1   g13411(.A1(new_n13667_), .A2(new_n13664_), .B(new_n13653_), .ZN(new_n13668_));
  NOR2_X1    g13412(.A1(new_n13668_), .A2(new_n13666_), .ZN(new_n13669_));
  INV_X1     g13413(.I(new_n13669_), .ZN(new_n13670_));
  OAI22_X1   g13414(.A1(new_n1592_), .A2(new_n8776_), .B1(new_n8500_), .B2(new_n1505_), .ZN(new_n13671_));
  AOI21_X1   g13415(.A1(\b[49] ), .A2(new_n1584_), .B(new_n13671_), .ZN(new_n13672_));
  OAI21_X1   g13416(.A1(new_n11577_), .A2(new_n1732_), .B(new_n13672_), .ZN(new_n13673_));
  XOR2_X1    g13417(.A1(new_n13673_), .A2(\a[17] ), .Z(new_n13674_));
  NAND2_X1   g13418(.A1(new_n13410_), .A2(new_n13395_), .ZN(new_n13675_));
  NAND2_X1   g13419(.A1(new_n13675_), .A2(new_n13674_), .ZN(new_n13676_));
  INV_X1     g13420(.I(new_n13676_), .ZN(new_n13677_));
  NOR2_X1    g13421(.A1(new_n13675_), .A2(new_n13674_), .ZN(new_n13678_));
  NOR3_X1    g13422(.A1(new_n13677_), .A2(new_n13670_), .A3(new_n13678_), .ZN(new_n13679_));
  INV_X1     g13423(.I(new_n13678_), .ZN(new_n13680_));
  AOI21_X1   g13424(.A1(new_n13680_), .A2(new_n13676_), .B(new_n13669_), .ZN(new_n13681_));
  NOR2_X1    g13425(.A1(new_n13681_), .A2(new_n13679_), .ZN(new_n13682_));
  NOR3_X1    g13426(.A1(new_n13070_), .A2(new_n13065_), .A3(new_n13415_), .ZN(new_n13683_));
  OAI22_X1   g13427(.A1(new_n993_), .A2(new_n9942_), .B1(new_n9376_), .B2(new_n997_), .ZN(new_n13684_));
  AOI21_X1   g13428(.A1(\b[52] ), .A2(new_n1486_), .B(new_n13684_), .ZN(new_n13685_));
  OAI21_X1   g13429(.A1(new_n9952_), .A2(new_n1323_), .B(new_n13685_), .ZN(new_n13686_));
  XOR2_X1    g13430(.A1(new_n13686_), .A2(\a[14] ), .Z(new_n13687_));
  INV_X1     g13431(.I(new_n13687_), .ZN(new_n13688_));
  OAI21_X1   g13432(.A1(new_n13683_), .A2(new_n13414_), .B(new_n13688_), .ZN(new_n13689_));
  OR3_X2     g13433(.A1(new_n13683_), .A2(new_n13414_), .A3(new_n13688_), .Z(new_n13690_));
  NAND2_X1   g13434(.A1(new_n13690_), .A2(new_n13689_), .ZN(new_n13691_));
  XNOR2_X1   g13435(.A1(new_n13691_), .A2(new_n13682_), .ZN(new_n13692_));
  INV_X1     g13436(.I(new_n10631_), .ZN(new_n13693_));
  OAI22_X1   g13437(.A1(new_n713_), .A2(new_n10625_), .B1(new_n10308_), .B2(new_n717_), .ZN(new_n13694_));
  AOI21_X1   g13438(.A1(\b[55] ), .A2(new_n1126_), .B(new_n13694_), .ZN(new_n13695_));
  OAI21_X1   g13439(.A1(new_n13693_), .A2(new_n986_), .B(new_n13695_), .ZN(new_n13696_));
  XOR2_X1    g13440(.A1(new_n13696_), .A2(\a[11] ), .Z(new_n13697_));
  OAI21_X1   g13441(.A1(new_n13429_), .A2(new_n13431_), .B(new_n13697_), .ZN(new_n13698_));
  INV_X1     g13442(.I(new_n13697_), .ZN(new_n13699_));
  NAND3_X1   g13443(.A1(new_n13435_), .A2(new_n13425_), .A3(new_n13699_), .ZN(new_n13700_));
  NAND3_X1   g13444(.A1(new_n13692_), .A2(new_n13698_), .A3(new_n13700_), .ZN(new_n13701_));
  XOR2_X1    g13445(.A1(new_n13691_), .A2(new_n13682_), .Z(new_n13702_));
  AOI21_X1   g13446(.A1(new_n13435_), .A2(new_n13425_), .B(new_n13699_), .ZN(new_n13703_));
  NOR3_X1    g13447(.A1(new_n13429_), .A2(new_n13431_), .A3(new_n13697_), .ZN(new_n13704_));
  OAI21_X1   g13448(.A1(new_n13704_), .A2(new_n13703_), .B(new_n13702_), .ZN(new_n13705_));
  AOI21_X1   g13449(.A1(new_n13435_), .A2(new_n13436_), .B(new_n13161_), .ZN(new_n13706_));
  AOI22_X1   g13450(.A1(new_n518_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n636_), .ZN(new_n13707_));
  OAI21_X1   g13451(.A1(new_n11195_), .A2(new_n917_), .B(new_n13707_), .ZN(new_n13708_));
  AOI21_X1   g13452(.A1(new_n11836_), .A2(new_n618_), .B(new_n13708_), .ZN(new_n13709_));
  XOR2_X1    g13453(.A1(new_n13709_), .A2(new_n488_), .Z(new_n13710_));
  INV_X1     g13454(.I(new_n13710_), .ZN(new_n13711_));
  OAI21_X1   g13455(.A1(new_n13706_), .A2(new_n13159_), .B(new_n13711_), .ZN(new_n13712_));
  INV_X1     g13456(.I(new_n13159_), .ZN(new_n13713_));
  OAI21_X1   g13457(.A1(new_n13429_), .A2(new_n13433_), .B(new_n13160_), .ZN(new_n13714_));
  NAND3_X1   g13458(.A1(new_n13714_), .A2(new_n13713_), .A3(new_n13710_), .ZN(new_n13715_));
  AOI22_X1   g13459(.A1(new_n13705_), .A2(new_n13701_), .B1(new_n13712_), .B2(new_n13715_), .ZN(new_n13716_));
  NOR3_X1    g13460(.A1(new_n13702_), .A2(new_n13703_), .A3(new_n13704_), .ZN(new_n13717_));
  AOI21_X1   g13461(.A1(new_n13698_), .A2(new_n13700_), .B(new_n13692_), .ZN(new_n13718_));
  AOI21_X1   g13462(.A1(new_n13714_), .A2(new_n13713_), .B(new_n13710_), .ZN(new_n13719_));
  NOR3_X1    g13463(.A1(new_n13706_), .A2(new_n13159_), .A3(new_n13711_), .ZN(new_n13720_));
  NOR4_X1    g13464(.A1(new_n13718_), .A2(new_n13717_), .A3(new_n13719_), .A4(new_n13720_), .ZN(new_n13721_));
  OAI21_X1   g13465(.A1(new_n13721_), .A2(new_n13716_), .B(new_n13495_), .ZN(new_n13722_));
  OAI22_X1   g13466(.A1(new_n13718_), .A2(new_n13717_), .B1(new_n13719_), .B2(new_n13720_), .ZN(new_n13723_));
  NAND4_X1   g13467(.A1(new_n13705_), .A2(new_n13701_), .A3(new_n13712_), .A4(new_n13715_), .ZN(new_n13724_));
  NAND3_X1   g13468(.A1(new_n13723_), .A2(new_n13724_), .A3(new_n13494_), .ZN(new_n13725_));
  NAND3_X1   g13469(.A1(new_n13722_), .A2(new_n13725_), .A3(new_n13490_), .ZN(new_n13726_));
  INV_X1     g13470(.I(new_n13490_), .ZN(new_n13727_));
  AOI21_X1   g13471(.A1(new_n13723_), .A2(new_n13724_), .B(new_n13494_), .ZN(new_n13728_));
  NOR3_X1    g13472(.A1(new_n13721_), .A2(new_n13716_), .A3(new_n13495_), .ZN(new_n13729_));
  OAI21_X1   g13473(.A1(new_n13729_), .A2(new_n13728_), .B(new_n13727_), .ZN(new_n13730_));
  NAND2_X1   g13474(.A1(new_n13730_), .A2(new_n13726_), .ZN(new_n13731_));
  NAND2_X1   g13475(.A1(new_n13731_), .A2(new_n13487_), .ZN(new_n13732_));
  AND2_X2    g13476(.A1(new_n13449_), .A2(new_n13453_), .Z(new_n13733_));
  OAI21_X1   g13477(.A1(new_n13733_), .A2(new_n13467_), .B(new_n13465_), .ZN(new_n13734_));
  NAND3_X1   g13478(.A1(new_n13734_), .A2(new_n13726_), .A3(new_n13730_), .ZN(new_n13735_));
  NAND2_X1   g13479(.A1(new_n13732_), .A2(new_n13735_), .ZN(new_n13736_));
  XOR2_X1    g13480(.A1(new_n13485_), .A2(new_n13736_), .Z(\f[66] ));
  AOI21_X1   g13481(.A1(new_n13727_), .A2(new_n13725_), .B(new_n13728_), .ZN(new_n13738_));
  INV_X1     g13482(.I(new_n13738_), .ZN(new_n13739_));
  AOI21_X1   g13483(.A1(new_n13702_), .A2(new_n13698_), .B(new_n13704_), .ZN(new_n13740_));
  AOI21_X1   g13484(.A1(new_n13670_), .A2(new_n13676_), .B(new_n13678_), .ZN(new_n13741_));
  INV_X1     g13485(.I(new_n13741_), .ZN(new_n13742_));
  INV_X1     g13486(.I(new_n13651_), .ZN(new_n13743_));
  OAI21_X1   g13487(.A1(new_n13642_), .A2(new_n13650_), .B(new_n13743_), .ZN(new_n13744_));
  AND2_X2    g13488(.A1(new_n13632_), .A2(new_n13638_), .Z(new_n13745_));
  NOR2_X1    g13489(.A1(new_n13745_), .A2(new_n13639_), .ZN(new_n13746_));
  INV_X1     g13490(.I(new_n13746_), .ZN(new_n13747_));
  INV_X1     g13491(.I(new_n13630_), .ZN(new_n13748_));
  OAI21_X1   g13492(.A1(new_n13626_), .A2(new_n13628_), .B(new_n13621_), .ZN(new_n13749_));
  NAND2_X1   g13493(.A1(new_n13749_), .A2(new_n13748_), .ZN(new_n13750_));
  NOR2_X1    g13494(.A1(new_n13615_), .A2(new_n13619_), .ZN(new_n13751_));
  AOI22_X1   g13495(.A1(new_n13615_), .A2(new_n13619_), .B1(new_n13335_), .B2(new_n13496_), .ZN(new_n13752_));
  NAND2_X1   g13496(.A1(new_n13613_), .A2(new_n13500_), .ZN(new_n13753_));
  NAND2_X1   g13497(.A1(new_n13753_), .A2(new_n13612_), .ZN(new_n13754_));
  INV_X1     g13498(.I(new_n13602_), .ZN(new_n13755_));
  AOI21_X1   g13499(.A1(new_n13603_), .A2(new_n13600_), .B(new_n13502_), .ZN(new_n13756_));
  NOR2_X1    g13500(.A1(new_n13755_), .A2(new_n13756_), .ZN(new_n13757_));
  INV_X1     g13501(.I(new_n13591_), .ZN(new_n13758_));
  OAI21_X1   g13502(.A1(new_n13508_), .A2(new_n13594_), .B(new_n13758_), .ZN(new_n13759_));
  NOR2_X1    g13503(.A1(new_n13578_), .A2(new_n13582_), .ZN(new_n13760_));
  AOI21_X1   g13504(.A1(new_n13510_), .A2(new_n13584_), .B(new_n13760_), .ZN(new_n13761_));
  AOI21_X1   g13505(.A1(new_n13513_), .A2(new_n13576_), .B(new_n13574_), .ZN(new_n13762_));
  AOI21_X1   g13506(.A1(new_n13515_), .A2(new_n13567_), .B(new_n13565_), .ZN(new_n13763_));
  INV_X1     g13507(.I(new_n13558_), .ZN(new_n13764_));
  AOI21_X1   g13508(.A1(new_n13517_), .A2(new_n13764_), .B(new_n13557_), .ZN(new_n13765_));
  INV_X1     g13509(.I(new_n13546_), .ZN(new_n13766_));
  OAI21_X1   g13510(.A1(new_n13518_), .A2(new_n13548_), .B(new_n13766_), .ZN(new_n13767_));
  NOR2_X1    g13511(.A1(new_n13520_), .A2(new_n13539_), .ZN(new_n13768_));
  NOR2_X1    g13512(.A1(new_n13768_), .A2(new_n13537_), .ZN(new_n13769_));
  INV_X1     g13513(.I(new_n13769_), .ZN(new_n13770_));
  OAI22_X1   g13514(.A1(new_n13224_), .A2(new_n471_), .B1(new_n438_), .B2(new_n11923_), .ZN(new_n13771_));
  AOI21_X1   g13515(.A1(\b[5] ), .A2(new_n13223_), .B(new_n13771_), .ZN(new_n13772_));
  OAI21_X1   g13516(.A1(new_n485_), .A2(new_n11930_), .B(new_n13772_), .ZN(new_n13773_));
  XOR2_X1    g13517(.A1(new_n13773_), .A2(new_n12312_), .Z(new_n13774_));
  AOI22_X1   g13518(.A1(new_n12922_), .A2(\b[4] ), .B1(\b[3] ), .B2(new_n12923_), .ZN(new_n13775_));
  INV_X1     g13519(.I(new_n13775_), .ZN(new_n13776_));
  NAND2_X1   g13520(.A1(new_n13776_), .A2(\a[2] ), .ZN(new_n13777_));
  NOR2_X1    g13521(.A1(new_n13776_), .A2(\a[2] ), .ZN(new_n13778_));
  INV_X1     g13522(.I(new_n13778_), .ZN(new_n13779_));
  NAND2_X1   g13523(.A1(new_n13779_), .A2(new_n13777_), .ZN(new_n13780_));
  XOR2_X1    g13524(.A1(new_n13774_), .A2(new_n13780_), .Z(new_n13781_));
  INV_X1     g13525(.I(new_n13781_), .ZN(new_n13782_));
  AOI21_X1   g13526(.A1(new_n13524_), .A2(new_n13527_), .B(new_n13528_), .ZN(new_n13783_));
  INV_X1     g13527(.I(new_n13783_), .ZN(new_n13784_));
  AOI22_X1   g13528(.A1(new_n10981_), .A2(\b[10] ), .B1(new_n10979_), .B2(\b[9] ), .ZN(new_n13785_));
  OAI21_X1   g13529(.A1(new_n577_), .A2(new_n11306_), .B(new_n13785_), .ZN(new_n13786_));
  AOI21_X1   g13530(.A1(new_n1059_), .A2(new_n10984_), .B(new_n13786_), .ZN(new_n13787_));
  XOR2_X1    g13531(.A1(new_n13787_), .A2(\a[59] ), .Z(new_n13788_));
  NAND2_X1   g13532(.A1(new_n13788_), .A2(new_n13784_), .ZN(new_n13789_));
  OR2_X2     g13533(.A1(new_n13788_), .A2(new_n13784_), .Z(new_n13790_));
  NAND2_X1   g13534(.A1(new_n13790_), .A2(new_n13789_), .ZN(new_n13791_));
  XOR2_X1    g13535(.A1(new_n13791_), .A2(new_n13782_), .Z(new_n13792_));
  OAI22_X1   g13536(.A1(new_n11298_), .A2(new_n1070_), .B1(new_n941_), .B2(new_n11297_), .ZN(new_n13793_));
  AOI21_X1   g13537(.A1(\b[11] ), .A2(new_n11296_), .B(new_n13793_), .ZN(new_n13794_));
  OAI21_X1   g13538(.A1(new_n1082_), .A2(new_n10069_), .B(new_n13794_), .ZN(new_n13795_));
  XOR2_X1    g13539(.A1(new_n13795_), .A2(\a[56] ), .Z(new_n13796_));
  OR2_X2     g13540(.A1(new_n13792_), .A2(new_n13796_), .Z(new_n13797_));
  NAND2_X1   g13541(.A1(new_n13792_), .A2(new_n13796_), .ZN(new_n13798_));
  NAND2_X1   g13542(.A1(new_n13797_), .A2(new_n13798_), .ZN(new_n13799_));
  XOR2_X1    g13543(.A1(new_n13799_), .A2(new_n13770_), .Z(new_n13800_));
  AOI22_X1   g13544(.A1(new_n9125_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n9123_), .ZN(new_n13801_));
  OAI21_X1   g13545(.A1(new_n1093_), .A2(new_n9470_), .B(new_n13801_), .ZN(new_n13802_));
  AOI21_X1   g13546(.A1(new_n1701_), .A2(new_n9129_), .B(new_n13802_), .ZN(new_n13803_));
  XOR2_X1    g13547(.A1(new_n13803_), .A2(new_n9133_), .Z(new_n13804_));
  OR2_X2     g13548(.A1(new_n13800_), .A2(new_n13804_), .Z(new_n13805_));
  NAND2_X1   g13549(.A1(new_n13800_), .A2(new_n13804_), .ZN(new_n13806_));
  NAND2_X1   g13550(.A1(new_n13805_), .A2(new_n13806_), .ZN(new_n13807_));
  XNOR2_X1   g13551(.A1(new_n13807_), .A2(new_n13767_), .ZN(new_n13808_));
  AOI22_X1   g13552(.A1(new_n8241_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n8246_), .ZN(new_n13809_));
  OAI21_X1   g13553(.A1(new_n1432_), .A2(new_n9114_), .B(new_n13809_), .ZN(new_n13810_));
  AOI21_X1   g13554(.A1(new_n1695_), .A2(new_n8252_), .B(new_n13810_), .ZN(new_n13811_));
  XOR2_X1    g13555(.A1(new_n13811_), .A2(\a[50] ), .Z(new_n13812_));
  NAND2_X1   g13556(.A1(new_n13808_), .A2(new_n13812_), .ZN(new_n13813_));
  INV_X1     g13557(.I(new_n13813_), .ZN(new_n13814_));
  NOR2_X1    g13558(.A1(new_n13808_), .A2(new_n13812_), .ZN(new_n13815_));
  NOR2_X1    g13559(.A1(new_n13814_), .A2(new_n13815_), .ZN(new_n13816_));
  XOR2_X1    g13560(.A1(new_n13816_), .A2(new_n13765_), .Z(new_n13817_));
  AOI22_X1   g13561(.A1(new_n7403_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n7408_), .ZN(new_n13818_));
  OAI21_X1   g13562(.A1(new_n1860_), .A2(new_n9488_), .B(new_n13818_), .ZN(new_n13819_));
  AOI21_X1   g13563(.A1(new_n2659_), .A2(new_n7414_), .B(new_n13819_), .ZN(new_n13820_));
  XOR2_X1    g13564(.A1(new_n13820_), .A2(new_n7410_), .Z(new_n13821_));
  NOR2_X1    g13565(.A1(new_n13817_), .A2(new_n13821_), .ZN(new_n13822_));
  AND2_X2    g13566(.A1(new_n13817_), .A2(new_n13821_), .Z(new_n13823_));
  NOR2_X1    g13567(.A1(new_n13823_), .A2(new_n13822_), .ZN(new_n13824_));
  XNOR2_X1   g13568(.A1(new_n13824_), .A2(new_n13763_), .ZN(new_n13825_));
  OAI22_X1   g13569(.A1(new_n7730_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n7731_), .ZN(new_n13826_));
  AOI21_X1   g13570(.A1(\b[23] ), .A2(new_n6887_), .B(new_n13826_), .ZN(new_n13827_));
  OAI21_X1   g13571(.A1(new_n2655_), .A2(new_n7728_), .B(new_n13827_), .ZN(new_n13828_));
  XOR2_X1    g13572(.A1(new_n13828_), .A2(\a[44] ), .Z(new_n13829_));
  INV_X1     g13573(.I(new_n13829_), .ZN(new_n13830_));
  NAND2_X1   g13574(.A1(new_n13825_), .A2(new_n13830_), .ZN(new_n13831_));
  XOR2_X1    g13575(.A1(new_n13824_), .A2(new_n13763_), .Z(new_n13832_));
  NAND2_X1   g13576(.A1(new_n13832_), .A2(new_n13829_), .ZN(new_n13833_));
  NAND2_X1   g13577(.A1(new_n13831_), .A2(new_n13833_), .ZN(new_n13834_));
  XNOR2_X1   g13578(.A1(new_n13834_), .A2(new_n13762_), .ZN(new_n13835_));
  AOI22_X1   g13579(.A1(new_n6108_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n6111_), .ZN(new_n13836_));
  OAI21_X1   g13580(.A1(new_n3006_), .A2(new_n7708_), .B(new_n13836_), .ZN(new_n13837_));
  AOI21_X1   g13581(.A1(new_n3807_), .A2(new_n6105_), .B(new_n13837_), .ZN(new_n13838_));
  XOR2_X1    g13582(.A1(new_n13838_), .A2(new_n5849_), .Z(new_n13839_));
  NOR2_X1    g13583(.A1(new_n13835_), .A2(new_n13839_), .ZN(new_n13840_));
  XOR2_X1    g13584(.A1(new_n13834_), .A2(new_n13762_), .Z(new_n13841_));
  INV_X1     g13585(.I(new_n13839_), .ZN(new_n13842_));
  NOR2_X1    g13586(.A1(new_n13841_), .A2(new_n13842_), .ZN(new_n13843_));
  NOR2_X1    g13587(.A1(new_n13840_), .A2(new_n13843_), .ZN(new_n13844_));
  XNOR2_X1   g13588(.A1(new_n13844_), .A2(new_n13761_), .ZN(new_n13845_));
  AOI22_X1   g13589(.A1(new_n5155_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n5160_), .ZN(new_n13846_));
  OAI21_X1   g13590(.A1(new_n3592_), .A2(new_n6877_), .B(new_n13846_), .ZN(new_n13847_));
  AOI21_X1   g13591(.A1(new_n3796_), .A2(new_n5166_), .B(new_n13847_), .ZN(new_n13848_));
  XOR2_X1    g13592(.A1(new_n13848_), .A2(new_n5162_), .Z(new_n13849_));
  INV_X1     g13593(.I(new_n13849_), .ZN(new_n13850_));
  NAND2_X1   g13594(.A1(new_n13845_), .A2(new_n13850_), .ZN(new_n13851_));
  XOR2_X1    g13595(.A1(new_n13844_), .A2(new_n13761_), .Z(new_n13852_));
  NAND2_X1   g13596(.A1(new_n13852_), .A2(new_n13849_), .ZN(new_n13853_));
  NAND2_X1   g13597(.A1(new_n13851_), .A2(new_n13853_), .ZN(new_n13854_));
  XOR2_X1    g13598(.A1(new_n13854_), .A2(new_n13759_), .Z(new_n13855_));
  AOI22_X1   g13599(.A1(new_n4918_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n4921_), .ZN(new_n13856_));
  OAI21_X1   g13600(.A1(new_n4023_), .A2(new_n6099_), .B(new_n13856_), .ZN(new_n13857_));
  AOI21_X1   g13601(.A1(new_n5103_), .A2(new_n4699_), .B(new_n13857_), .ZN(new_n13858_));
  XOR2_X1    g13602(.A1(new_n13858_), .A2(new_n4446_), .Z(new_n13859_));
  XOR2_X1    g13603(.A1(new_n13855_), .A2(new_n13859_), .Z(new_n13860_));
  XOR2_X1    g13604(.A1(new_n13860_), .A2(new_n13757_), .Z(new_n13861_));
  OAI22_X1   g13605(.A1(new_n4886_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n5312_), .ZN(new_n13862_));
  AOI21_X1   g13606(.A1(\b[35] ), .A2(new_n4053_), .B(new_n13862_), .ZN(new_n13863_));
  OAI21_X1   g13607(.A1(new_n5322_), .A2(new_n4727_), .B(new_n13863_), .ZN(new_n13864_));
  XOR2_X1    g13608(.A1(new_n13864_), .A2(\a[32] ), .Z(new_n13865_));
  NOR2_X1    g13609(.A1(new_n13861_), .A2(new_n13865_), .ZN(new_n13866_));
  INV_X1     g13610(.I(new_n13757_), .ZN(new_n13867_));
  XOR2_X1    g13611(.A1(new_n13860_), .A2(new_n13867_), .Z(new_n13868_));
  INV_X1     g13612(.I(new_n13865_), .ZN(new_n13869_));
  NOR2_X1    g13613(.A1(new_n13868_), .A2(new_n13869_), .ZN(new_n13870_));
  NOR2_X1    g13614(.A1(new_n13866_), .A2(new_n13870_), .ZN(new_n13871_));
  XNOR2_X1   g13615(.A1(new_n13871_), .A2(new_n13754_), .ZN(new_n13872_));
  AOI22_X1   g13616(.A1(new_n3267_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n3270_), .ZN(new_n13873_));
  OAI21_X1   g13617(.A1(new_n5341_), .A2(new_n3475_), .B(new_n13873_), .ZN(new_n13874_));
  AOI21_X1   g13618(.A1(new_n5793_), .A2(new_n3273_), .B(new_n13874_), .ZN(new_n13875_));
  XOR2_X1    g13619(.A1(new_n13875_), .A2(new_n3264_), .Z(new_n13876_));
  NOR2_X1    g13620(.A1(new_n13872_), .A2(new_n13876_), .ZN(new_n13877_));
  XOR2_X1    g13621(.A1(new_n13871_), .A2(new_n13754_), .Z(new_n13878_));
  INV_X1     g13622(.I(new_n13876_), .ZN(new_n13879_));
  NOR2_X1    g13623(.A1(new_n13878_), .A2(new_n13879_), .ZN(new_n13880_));
  OAI22_X1   g13624(.A1(new_n13877_), .A2(new_n13880_), .B1(new_n13751_), .B2(new_n13752_), .ZN(new_n13881_));
  NOR2_X1    g13625(.A1(new_n13752_), .A2(new_n13751_), .ZN(new_n13882_));
  NOR2_X1    g13626(.A1(new_n13877_), .A2(new_n13880_), .ZN(new_n13883_));
  NAND2_X1   g13627(.A1(new_n13883_), .A2(new_n13882_), .ZN(new_n13884_));
  NAND2_X1   g13628(.A1(new_n13884_), .A2(new_n13881_), .ZN(new_n13885_));
  OAI22_X1   g13629(.A1(new_n2703_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n2708_), .ZN(new_n13886_));
  AOI21_X1   g13630(.A1(\b[41] ), .A2(new_n2906_), .B(new_n13886_), .ZN(new_n13887_));
  OAI21_X1   g13631(.A1(new_n6785_), .A2(new_n2711_), .B(new_n13887_), .ZN(new_n13888_));
  XOR2_X1    g13632(.A1(new_n13888_), .A2(\a[26] ), .Z(new_n13889_));
  INV_X1     g13633(.I(new_n13889_), .ZN(new_n13890_));
  NAND2_X1   g13634(.A1(new_n13885_), .A2(new_n13890_), .ZN(new_n13891_));
  NAND3_X1   g13635(.A1(new_n13884_), .A2(new_n13881_), .A3(new_n13889_), .ZN(new_n13892_));
  NAND2_X1   g13636(.A1(new_n13891_), .A2(new_n13892_), .ZN(new_n13893_));
  XNOR2_X1   g13637(.A1(new_n13893_), .A2(new_n13750_), .ZN(new_n13894_));
  AOI22_X1   g13638(.A1(new_n2202_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n2205_), .ZN(new_n13895_));
  OAI21_X1   g13639(.A1(new_n7074_), .A2(new_n2370_), .B(new_n13895_), .ZN(new_n13896_));
  AOI21_X1   g13640(.A1(new_n9337_), .A2(new_n2208_), .B(new_n13896_), .ZN(new_n13897_));
  XOR2_X1    g13641(.A1(new_n13897_), .A2(new_n2200_), .Z(new_n13898_));
  INV_X1     g13642(.I(new_n13898_), .ZN(new_n13899_));
  NAND2_X1   g13643(.A1(new_n13894_), .A2(new_n13899_), .ZN(new_n13900_));
  XOR2_X1    g13644(.A1(new_n13893_), .A2(new_n13750_), .Z(new_n13901_));
  NAND2_X1   g13645(.A1(new_n13901_), .A2(new_n13898_), .ZN(new_n13902_));
  NAND2_X1   g13646(.A1(new_n13900_), .A2(new_n13902_), .ZN(new_n13903_));
  NOR2_X1    g13647(.A1(new_n13903_), .A2(new_n13747_), .ZN(new_n13904_));
  NOR2_X1    g13648(.A1(new_n13901_), .A2(new_n13898_), .ZN(new_n13905_));
  NOR2_X1    g13649(.A1(new_n13894_), .A2(new_n13899_), .ZN(new_n13906_));
  NOR2_X1    g13650(.A1(new_n13906_), .A2(new_n13905_), .ZN(new_n13907_));
  NOR2_X1    g13651(.A1(new_n13907_), .A2(new_n13746_), .ZN(new_n13908_));
  OAI22_X1   g13652(.A1(new_n1751_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n1754_), .ZN(new_n13909_));
  AOI21_X1   g13653(.A1(\b[47] ), .A2(new_n1939_), .B(new_n13909_), .ZN(new_n13910_));
  OAI21_X1   g13654(.A1(new_n9050_), .A2(new_n1757_), .B(new_n13910_), .ZN(new_n13911_));
  XOR2_X1    g13655(.A1(new_n13911_), .A2(\a[20] ), .Z(new_n13912_));
  INV_X1     g13656(.I(new_n13912_), .ZN(new_n13913_));
  OAI21_X1   g13657(.A1(new_n13908_), .A2(new_n13904_), .B(new_n13913_), .ZN(new_n13914_));
  NAND2_X1   g13658(.A1(new_n13907_), .A2(new_n13746_), .ZN(new_n13915_));
  NAND2_X1   g13659(.A1(new_n13903_), .A2(new_n13747_), .ZN(new_n13916_));
  NAND3_X1   g13660(.A1(new_n13915_), .A2(new_n13916_), .A3(new_n13912_), .ZN(new_n13917_));
  NAND2_X1   g13661(.A1(new_n13914_), .A2(new_n13917_), .ZN(new_n13918_));
  XNOR2_X1   g13662(.A1(new_n13918_), .A2(new_n13744_), .ZN(new_n13919_));
  AOI21_X1   g13663(.A1(new_n13654_), .A2(new_n13667_), .B(new_n13665_), .ZN(new_n13920_));
  OAI22_X1   g13664(.A1(new_n1592_), .A2(new_n9032_), .B1(new_n8776_), .B2(new_n1505_), .ZN(new_n13921_));
  AOI21_X1   g13665(.A1(\b[50] ), .A2(new_n1584_), .B(new_n13921_), .ZN(new_n13922_));
  OAI21_X1   g13666(.A1(new_n9043_), .A2(new_n1732_), .B(new_n13922_), .ZN(new_n13923_));
  XOR2_X1    g13667(.A1(new_n13923_), .A2(\a[17] ), .Z(new_n13924_));
  NOR2_X1    g13668(.A1(new_n13920_), .A2(new_n13924_), .ZN(new_n13925_));
  INV_X1     g13669(.I(new_n13925_), .ZN(new_n13926_));
  NAND2_X1   g13670(.A1(new_n13920_), .A2(new_n13924_), .ZN(new_n13927_));
  NAND2_X1   g13671(.A1(new_n13926_), .A2(new_n13927_), .ZN(new_n13928_));
  NAND2_X1   g13672(.A1(new_n13919_), .A2(new_n13928_), .ZN(new_n13929_));
  XOR2_X1    g13673(.A1(new_n13918_), .A2(new_n13744_), .Z(new_n13930_));
  INV_X1     g13674(.I(new_n13927_), .ZN(new_n13931_));
  NOR2_X1    g13675(.A1(new_n13931_), .A2(new_n13925_), .ZN(new_n13932_));
  NAND2_X1   g13676(.A1(new_n13930_), .A2(new_n13932_), .ZN(new_n13933_));
  OAI22_X1   g13677(.A1(new_n993_), .A2(new_n9972_), .B1(new_n9942_), .B2(new_n997_), .ZN(new_n13934_));
  AOI21_X1   g13678(.A1(\b[53] ), .A2(new_n1486_), .B(new_n13934_), .ZN(new_n13935_));
  OAI21_X1   g13679(.A1(new_n13080_), .A2(new_n1323_), .B(new_n13935_), .ZN(new_n13936_));
  XOR2_X1    g13680(.A1(new_n13936_), .A2(\a[14] ), .Z(new_n13937_));
  AOI21_X1   g13681(.A1(new_n13929_), .A2(new_n13933_), .B(new_n13937_), .ZN(new_n13938_));
  NOR2_X1    g13682(.A1(new_n13930_), .A2(new_n13932_), .ZN(new_n13939_));
  NOR2_X1    g13683(.A1(new_n13919_), .A2(new_n13928_), .ZN(new_n13940_));
  INV_X1     g13684(.I(new_n13937_), .ZN(new_n13941_));
  NOR3_X1    g13685(.A1(new_n13940_), .A2(new_n13939_), .A3(new_n13941_), .ZN(new_n13942_));
  NOR3_X1    g13686(.A1(new_n13942_), .A2(new_n13938_), .A3(new_n13742_), .ZN(new_n13943_));
  OAI21_X1   g13687(.A1(new_n13940_), .A2(new_n13939_), .B(new_n13941_), .ZN(new_n13944_));
  NAND3_X1   g13688(.A1(new_n13929_), .A2(new_n13933_), .A3(new_n13937_), .ZN(new_n13945_));
  AOI21_X1   g13689(.A1(new_n13944_), .A2(new_n13945_), .B(new_n13741_), .ZN(new_n13946_));
  NOR2_X1    g13690(.A1(new_n13943_), .A2(new_n13946_), .ZN(new_n13947_));
  OAI21_X1   g13691(.A1(new_n13679_), .A2(new_n13681_), .B(new_n13690_), .ZN(new_n13948_));
  OAI22_X1   g13692(.A1(new_n713_), .A2(new_n11195_), .B1(new_n10625_), .B2(new_n717_), .ZN(new_n13949_));
  AOI21_X1   g13693(.A1(\b[56] ), .A2(new_n1126_), .B(new_n13949_), .ZN(new_n13950_));
  OAI21_X1   g13694(.A1(new_n11206_), .A2(new_n986_), .B(new_n13950_), .ZN(new_n13951_));
  XOR2_X1    g13695(.A1(new_n13951_), .A2(\a[11] ), .Z(new_n13952_));
  AOI21_X1   g13696(.A1(new_n13948_), .A2(new_n13689_), .B(new_n13952_), .ZN(new_n13953_));
  NAND2_X1   g13697(.A1(new_n13948_), .A2(new_n13689_), .ZN(new_n13954_));
  INV_X1     g13698(.I(new_n13952_), .ZN(new_n13955_));
  NOR2_X1    g13699(.A1(new_n13954_), .A2(new_n13955_), .ZN(new_n13956_));
  NOR2_X1    g13700(.A1(new_n13956_), .A2(new_n13953_), .ZN(new_n13957_));
  NOR2_X1    g13701(.A1(new_n13957_), .A2(new_n13947_), .ZN(new_n13958_));
  INV_X1     g13702(.I(new_n13947_), .ZN(new_n13959_));
  NOR3_X1    g13703(.A1(new_n13959_), .A2(new_n13953_), .A3(new_n13956_), .ZN(new_n13960_));
  OAI22_X1   g13704(.A1(new_n610_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n612_), .ZN(new_n13961_));
  AOI21_X1   g13705(.A1(\b[59] ), .A2(new_n826_), .B(new_n13961_), .ZN(new_n13962_));
  OAI21_X1   g13706(.A1(new_n13110_), .A2(new_n624_), .B(new_n13962_), .ZN(new_n13963_));
  XOR2_X1    g13707(.A1(new_n13963_), .A2(\a[8] ), .Z(new_n13964_));
  INV_X1     g13708(.I(new_n13964_), .ZN(new_n13965_));
  OAI21_X1   g13709(.A1(new_n13960_), .A2(new_n13958_), .B(new_n13965_), .ZN(new_n13966_));
  INV_X1     g13710(.I(new_n13958_), .ZN(new_n13967_));
  NAND2_X1   g13711(.A1(new_n13957_), .A2(new_n13947_), .ZN(new_n13968_));
  NAND3_X1   g13712(.A1(new_n13967_), .A2(new_n13968_), .A3(new_n13964_), .ZN(new_n13969_));
  NAND2_X1   g13713(.A1(new_n13969_), .A2(new_n13966_), .ZN(new_n13970_));
  XOR2_X1    g13714(.A1(new_n13970_), .A2(new_n13740_), .Z(new_n13971_));
  OAI21_X1   g13715(.A1(new_n13718_), .A2(new_n13717_), .B(new_n13715_), .ZN(new_n13972_));
  INV_X1     g13716(.I(new_n13107_), .ZN(new_n13973_));
  OAI22_X1   g13717(.A1(new_n392_), .A2(new_n12796_), .B1(new_n325_), .B2(new_n12800_), .ZN(new_n13974_));
  AOI21_X1   g13718(.A1(new_n13973_), .A2(new_n330_), .B(new_n13974_), .ZN(new_n13975_));
  XOR2_X1    g13719(.A1(new_n13975_), .A2(new_n312_), .Z(new_n13976_));
  AOI21_X1   g13720(.A1(new_n13972_), .A2(new_n13712_), .B(new_n13976_), .ZN(new_n13977_));
  NAND3_X1   g13721(.A1(new_n13972_), .A2(new_n13712_), .A3(new_n13976_), .ZN(new_n13978_));
  INV_X1     g13722(.I(new_n13978_), .ZN(new_n13979_));
  NOR2_X1    g13723(.A1(new_n13979_), .A2(new_n13977_), .ZN(new_n13980_));
  XNOR2_X1   g13724(.A1(new_n13971_), .A2(new_n13980_), .ZN(new_n13981_));
  AOI21_X1   g13725(.A1(new_n13726_), .A2(new_n13730_), .B(new_n13734_), .ZN(new_n13982_));
  INV_X1     g13726(.I(new_n13726_), .ZN(new_n13983_));
  AOI21_X1   g13727(.A1(new_n13722_), .A2(new_n13725_), .B(new_n13490_), .ZN(new_n13984_));
  NOR3_X1    g13728(.A1(new_n13983_), .A2(new_n13487_), .A3(new_n13984_), .ZN(new_n13985_));
  NOR2_X1    g13729(.A1(new_n13982_), .A2(new_n13985_), .ZN(new_n13986_));
  NOR3_X1    g13730(.A1(new_n13484_), .A2(new_n13472_), .A3(new_n13986_), .ZN(new_n13987_));
  NOR2_X1    g13731(.A1(new_n13731_), .A2(new_n13734_), .ZN(new_n13988_));
  OAI21_X1   g13732(.A1(new_n13987_), .A2(new_n13988_), .B(new_n13981_), .ZN(new_n13989_));
  XOR2_X1    g13733(.A1(new_n13971_), .A2(new_n13980_), .Z(new_n13990_));
  INV_X1     g13734(.I(new_n13472_), .ZN(new_n13991_));
  OAI21_X1   g13735(.A1(new_n13471_), .A2(new_n13469_), .B(new_n13148_), .ZN(new_n13992_));
  OAI21_X1   g13736(.A1(new_n13140_), .A2(new_n13137_), .B(new_n13992_), .ZN(new_n13993_));
  NAND3_X1   g13737(.A1(new_n13993_), .A2(new_n13991_), .A3(new_n13736_), .ZN(new_n13994_));
  INV_X1     g13738(.I(new_n13988_), .ZN(new_n13995_));
  NAND3_X1   g13739(.A1(new_n13994_), .A2(new_n13990_), .A3(new_n13995_), .ZN(new_n13996_));
  NAND2_X1   g13740(.A1(new_n13989_), .A2(new_n13996_), .ZN(new_n13997_));
  XOR2_X1    g13741(.A1(new_n13997_), .A2(new_n13739_), .Z(\f[67] ));
  AOI21_X1   g13742(.A1(new_n13994_), .A2(new_n13995_), .B(new_n13990_), .ZN(new_n13999_));
  OAI21_X1   g13743(.A1(new_n13738_), .A2(new_n13999_), .B(new_n13996_), .ZN(new_n14000_));
  AOI21_X1   g13744(.A1(new_n13971_), .A2(new_n13978_), .B(new_n13977_), .ZN(new_n14001_));
  AOI22_X1   g13745(.A1(new_n13460_), .A2(new_n330_), .B1(\b[63] ), .B2(new_n602_), .ZN(new_n14002_));
  XOR2_X1    g13746(.A1(new_n14002_), .A2(new_n312_), .Z(new_n14003_));
  INV_X1     g13747(.I(new_n14003_), .ZN(new_n14004_));
  INV_X1     g13748(.I(new_n13740_), .ZN(new_n14005_));
  NAND2_X1   g13749(.A1(new_n13969_), .A2(new_n14005_), .ZN(new_n14006_));
  NAND2_X1   g13750(.A1(new_n14006_), .A2(new_n13966_), .ZN(new_n14007_));
  INV_X1     g13751(.I(new_n14007_), .ZN(new_n14008_));
  AOI21_X1   g13752(.A1(new_n13742_), .A2(new_n13945_), .B(new_n13938_), .ZN(new_n14009_));
  INV_X1     g13753(.I(new_n14009_), .ZN(new_n14010_));
  OAI21_X1   g13754(.A1(new_n13930_), .A2(new_n13931_), .B(new_n13926_), .ZN(new_n14011_));
  INV_X1     g13755(.I(new_n14011_), .ZN(new_n14012_));
  NAND2_X1   g13756(.A1(new_n13917_), .A2(new_n13744_), .ZN(new_n14013_));
  AOI21_X1   g13757(.A1(new_n13747_), .A2(new_n13902_), .B(new_n13905_), .ZN(new_n14014_));
  NAND2_X1   g13758(.A1(new_n13750_), .A2(new_n13892_), .ZN(new_n14015_));
  NAND2_X1   g13759(.A1(new_n14015_), .A2(new_n13891_), .ZN(new_n14016_));
  NOR2_X1    g13760(.A1(new_n13880_), .A2(new_n13882_), .ZN(new_n14017_));
  NOR2_X1    g13761(.A1(new_n14017_), .A2(new_n13877_), .ZN(new_n14018_));
  INV_X1     g13762(.I(new_n14018_), .ZN(new_n14019_));
  INV_X1     g13763(.I(new_n13870_), .ZN(new_n14020_));
  AOI21_X1   g13764(.A1(new_n14020_), .A2(new_n13754_), .B(new_n13866_), .ZN(new_n14021_));
  NOR2_X1    g13765(.A1(new_n13855_), .A2(new_n13859_), .ZN(new_n14022_));
  NAND2_X1   g13766(.A1(new_n13855_), .A2(new_n13859_), .ZN(new_n14023_));
  AOI21_X1   g13767(.A1(new_n13867_), .A2(new_n14023_), .B(new_n14022_), .ZN(new_n14024_));
  INV_X1     g13768(.I(new_n13851_), .ZN(new_n14025_));
  AOI21_X1   g13769(.A1(new_n13759_), .A2(new_n13853_), .B(new_n14025_), .ZN(new_n14026_));
  INV_X1     g13770(.I(new_n13840_), .ZN(new_n14027_));
  OAI21_X1   g13771(.A1(new_n13761_), .A2(new_n13843_), .B(new_n14027_), .ZN(new_n14028_));
  INV_X1     g13772(.I(new_n13833_), .ZN(new_n14029_));
  OAI21_X1   g13773(.A1(new_n14029_), .A2(new_n13762_), .B(new_n13831_), .ZN(new_n14030_));
  AOI22_X1   g13774(.A1(new_n6569_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n6574_), .ZN(new_n14031_));
  OAI21_X1   g13775(.A1(new_n2495_), .A2(new_n8565_), .B(new_n14031_), .ZN(new_n14032_));
  AOI21_X1   g13776(.A1(new_n3407_), .A2(new_n6579_), .B(new_n14032_), .ZN(new_n14033_));
  XOR2_X1    g13777(.A1(new_n14033_), .A2(new_n6567_), .Z(new_n14034_));
  INV_X1     g13778(.I(new_n14034_), .ZN(new_n14035_));
  INV_X1     g13779(.I(new_n13822_), .ZN(new_n14036_));
  OAI21_X1   g13780(.A1(new_n13763_), .A2(new_n13823_), .B(new_n14036_), .ZN(new_n14037_));
  OAI21_X1   g13781(.A1(new_n13765_), .A2(new_n13815_), .B(new_n13813_), .ZN(new_n14038_));
  INV_X1     g13782(.I(new_n14038_), .ZN(new_n14039_));
  INV_X1     g13783(.I(new_n13805_), .ZN(new_n14040_));
  AOI21_X1   g13784(.A1(new_n13767_), .A2(new_n13806_), .B(new_n14040_), .ZN(new_n14041_));
  NAND2_X1   g13785(.A1(new_n13770_), .A2(new_n13798_), .ZN(new_n14042_));
  AND2_X2    g13786(.A1(new_n14042_), .A2(new_n13797_), .Z(new_n14043_));
  INV_X1     g13787(.I(new_n14043_), .ZN(new_n14044_));
  AOI22_X1   g13788(.A1(new_n10064_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n10062_), .ZN(new_n14045_));
  OAI21_X1   g13789(.A1(new_n941_), .A2(new_n10399_), .B(new_n14045_), .ZN(new_n14046_));
  AOI21_X1   g13790(.A1(new_n1449_), .A2(new_n10068_), .B(new_n14046_), .ZN(new_n14047_));
  XOR2_X1    g13791(.A1(new_n14047_), .A2(new_n10057_), .Z(new_n14048_));
  AOI21_X1   g13792(.A1(new_n13774_), .A2(new_n13777_), .B(new_n13778_), .ZN(new_n14049_));
  INV_X1     g13793(.I(new_n14049_), .ZN(new_n14050_));
  OAI22_X1   g13794(.A1(new_n12306_), .A2(new_n852_), .B1(new_n12305_), .B2(new_n776_), .ZN(new_n14051_));
  AOI21_X1   g13795(.A1(\b[9] ), .A2(new_n12304_), .B(new_n14051_), .ZN(new_n14052_));
  OAI21_X1   g13796(.A1(new_n859_), .A2(new_n10985_), .B(new_n14052_), .ZN(new_n14053_));
  XOR2_X1    g13797(.A1(new_n14053_), .A2(new_n10989_), .Z(new_n14054_));
  NAND2_X1   g13798(.A1(new_n14054_), .A2(new_n14050_), .ZN(new_n14055_));
  XOR2_X1    g13799(.A1(new_n14053_), .A2(\a[59] ), .Z(new_n14056_));
  NAND2_X1   g13800(.A1(new_n14056_), .A2(new_n14049_), .ZN(new_n14057_));
  NAND2_X1   g13801(.A1(new_n14055_), .A2(new_n14057_), .ZN(new_n14058_));
  AOI22_X1   g13802(.A1(new_n11926_), .A2(\b[8] ), .B1(new_n11924_), .B2(\b[7] ), .ZN(new_n14059_));
  OAI21_X1   g13803(.A1(new_n438_), .A2(new_n12317_), .B(new_n14059_), .ZN(new_n14060_));
  AOI21_X1   g13804(.A1(new_n799_), .A2(new_n11929_), .B(new_n14060_), .ZN(new_n14061_));
  XOR2_X1    g13805(.A1(new_n14061_), .A2(\a[62] ), .Z(new_n14062_));
  AOI22_X1   g13806(.A1(new_n12922_), .A2(\b[5] ), .B1(\b[4] ), .B2(new_n12923_), .ZN(new_n14063_));
  INV_X1     g13807(.I(new_n14063_), .ZN(new_n14064_));
  NAND2_X1   g13808(.A1(new_n14064_), .A2(\a[2] ), .ZN(new_n14065_));
  NOR2_X1    g13809(.A1(new_n14064_), .A2(\a[2] ), .ZN(new_n14066_));
  INV_X1     g13810(.I(new_n14066_), .ZN(new_n14067_));
  NAND2_X1   g13811(.A1(new_n14067_), .A2(new_n14065_), .ZN(new_n14068_));
  XOR2_X1    g13812(.A1(new_n14062_), .A2(new_n14068_), .Z(new_n14069_));
  XOR2_X1    g13813(.A1(new_n14058_), .A2(new_n14069_), .Z(new_n14070_));
  NAND2_X1   g13814(.A1(new_n13790_), .A2(new_n13782_), .ZN(new_n14071_));
  NAND2_X1   g13815(.A1(new_n14071_), .A2(new_n13789_), .ZN(new_n14072_));
  NAND2_X1   g13816(.A1(new_n14070_), .A2(new_n14072_), .ZN(new_n14073_));
  INV_X1     g13817(.I(new_n14069_), .ZN(new_n14074_));
  XOR2_X1    g13818(.A1(new_n14058_), .A2(new_n14074_), .Z(new_n14075_));
  NAND3_X1   g13819(.A1(new_n14075_), .A2(new_n13789_), .A3(new_n14071_), .ZN(new_n14076_));
  NAND2_X1   g13820(.A1(new_n14076_), .A2(new_n14073_), .ZN(new_n14077_));
  XOR2_X1    g13821(.A1(new_n14077_), .A2(new_n14048_), .Z(new_n14078_));
  OAI22_X1   g13822(.A1(new_n10390_), .A2(new_n1432_), .B1(new_n1296_), .B2(new_n10389_), .ZN(new_n14079_));
  AOI21_X1   g13823(.A1(\b[15] ), .A2(new_n9471_), .B(new_n14079_), .ZN(new_n14080_));
  OAI21_X1   g13824(.A1(new_n1444_), .A2(new_n10388_), .B(new_n14080_), .ZN(new_n14081_));
  XOR2_X1    g13825(.A1(new_n14081_), .A2(\a[53] ), .Z(new_n14082_));
  INV_X1     g13826(.I(new_n14082_), .ZN(new_n14083_));
  NAND2_X1   g13827(.A1(new_n14078_), .A2(new_n14083_), .ZN(new_n14084_));
  INV_X1     g13828(.I(new_n14048_), .ZN(new_n14085_));
  XOR2_X1    g13829(.A1(new_n14077_), .A2(new_n14085_), .Z(new_n14086_));
  NAND2_X1   g13830(.A1(new_n14086_), .A2(new_n14082_), .ZN(new_n14087_));
  NAND2_X1   g13831(.A1(new_n14084_), .A2(new_n14087_), .ZN(new_n14088_));
  XOR2_X1    g13832(.A1(new_n14088_), .A2(new_n14044_), .Z(new_n14089_));
  AOI22_X1   g13833(.A1(new_n8241_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n8246_), .ZN(new_n14090_));
  OAI21_X1   g13834(.A1(new_n1553_), .A2(new_n9114_), .B(new_n14090_), .ZN(new_n14091_));
  AOI21_X1   g13835(.A1(new_n2452_), .A2(new_n8252_), .B(new_n14091_), .ZN(new_n14092_));
  XOR2_X1    g13836(.A1(new_n14092_), .A2(new_n8248_), .Z(new_n14093_));
  NOR2_X1    g13837(.A1(new_n14089_), .A2(new_n14093_), .ZN(new_n14094_));
  XOR2_X1    g13838(.A1(new_n14088_), .A2(new_n14043_), .Z(new_n14095_));
  INV_X1     g13839(.I(new_n14093_), .ZN(new_n14096_));
  NOR2_X1    g13840(.A1(new_n14095_), .A2(new_n14096_), .ZN(new_n14097_));
  OR2_X2     g13841(.A1(new_n14094_), .A2(new_n14097_), .Z(new_n14098_));
  XOR2_X1    g13842(.A1(new_n14098_), .A2(new_n14041_), .Z(new_n14099_));
  AOI22_X1   g13843(.A1(new_n7403_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n7408_), .ZN(new_n14100_));
  OAI21_X1   g13844(.A1(new_n2027_), .A2(new_n9488_), .B(new_n14100_), .ZN(new_n14101_));
  AOI21_X1   g13845(.A1(new_n2470_), .A2(new_n7414_), .B(new_n14101_), .ZN(new_n14102_));
  XOR2_X1    g13846(.A1(new_n14102_), .A2(new_n7410_), .Z(new_n14103_));
  INV_X1     g13847(.I(new_n14103_), .ZN(new_n14104_));
  NAND2_X1   g13848(.A1(new_n14099_), .A2(new_n14104_), .ZN(new_n14105_));
  XNOR2_X1   g13849(.A1(new_n14098_), .A2(new_n14041_), .ZN(new_n14106_));
  NAND2_X1   g13850(.A1(new_n14106_), .A2(new_n14103_), .ZN(new_n14107_));
  AOI21_X1   g13851(.A1(new_n14107_), .A2(new_n14105_), .B(new_n14039_), .ZN(new_n14108_));
  NAND2_X1   g13852(.A1(new_n14107_), .A2(new_n14105_), .ZN(new_n14109_));
  NOR2_X1    g13853(.A1(new_n14109_), .A2(new_n14038_), .ZN(new_n14110_));
  OAI21_X1   g13854(.A1(new_n14108_), .A2(new_n14110_), .B(new_n14037_), .ZN(new_n14111_));
  OR3_X2     g13855(.A1(new_n14037_), .A2(new_n14108_), .A3(new_n14110_), .Z(new_n14112_));
  NAND2_X1   g13856(.A1(new_n14112_), .A2(new_n14111_), .ZN(new_n14113_));
  XOR2_X1    g13857(.A1(new_n14113_), .A2(new_n14035_), .Z(new_n14114_));
  AOI22_X1   g13858(.A1(new_n6108_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n6111_), .ZN(new_n14115_));
  OAI21_X1   g13859(.A1(new_n3158_), .A2(new_n7708_), .B(new_n14115_), .ZN(new_n14116_));
  AOI21_X1   g13860(.A1(new_n4188_), .A2(new_n6105_), .B(new_n14116_), .ZN(new_n14117_));
  XOR2_X1    g13861(.A1(new_n14117_), .A2(new_n5849_), .Z(new_n14118_));
  OR2_X2     g13862(.A1(new_n14114_), .A2(new_n14118_), .Z(new_n14119_));
  NAND2_X1   g13863(.A1(new_n14114_), .A2(new_n14118_), .ZN(new_n14120_));
  NAND2_X1   g13864(.A1(new_n14119_), .A2(new_n14120_), .ZN(new_n14121_));
  XOR2_X1    g13865(.A1(new_n14121_), .A2(new_n14030_), .Z(new_n14122_));
  AOI22_X1   g13866(.A1(new_n5155_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n5160_), .ZN(new_n14123_));
  OAI21_X1   g13867(.A1(new_n3624_), .A2(new_n6877_), .B(new_n14123_), .ZN(new_n14124_));
  AOI21_X1   g13868(.A1(new_n4030_), .A2(new_n5166_), .B(new_n14124_), .ZN(new_n14125_));
  XOR2_X1    g13869(.A1(new_n14125_), .A2(new_n5162_), .Z(new_n14126_));
  NOR2_X1    g13870(.A1(new_n14122_), .A2(new_n14126_), .ZN(new_n14127_));
  XNOR2_X1   g13871(.A1(new_n14121_), .A2(new_n14030_), .ZN(new_n14128_));
  INV_X1     g13872(.I(new_n14126_), .ZN(new_n14129_));
  NOR2_X1    g13873(.A1(new_n14128_), .A2(new_n14129_), .ZN(new_n14130_));
  NOR2_X1    g13874(.A1(new_n14130_), .A2(new_n14127_), .ZN(new_n14131_));
  XOR2_X1    g13875(.A1(new_n14131_), .A2(new_n14028_), .Z(new_n14132_));
  OAI22_X1   g13876(.A1(new_n4666_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n4639_), .ZN(new_n14133_));
  AOI21_X1   g13877(.A1(\b[33] ), .A2(new_n4706_), .B(new_n14133_), .ZN(new_n14134_));
  OAI21_X1   g13878(.A1(new_n4676_), .A2(new_n4458_), .B(new_n14134_), .ZN(new_n14135_));
  XOR2_X1    g13879(.A1(new_n14135_), .A2(\a[35] ), .Z(new_n14136_));
  INV_X1     g13880(.I(new_n14136_), .ZN(new_n14137_));
  NAND2_X1   g13881(.A1(new_n14132_), .A2(new_n14137_), .ZN(new_n14138_));
  INV_X1     g13882(.I(new_n14028_), .ZN(new_n14139_));
  XOR2_X1    g13883(.A1(new_n14131_), .A2(new_n14139_), .Z(new_n14140_));
  NAND2_X1   g13884(.A1(new_n14140_), .A2(new_n14136_), .ZN(new_n14141_));
  NAND2_X1   g13885(.A1(new_n14138_), .A2(new_n14141_), .ZN(new_n14142_));
  XOR2_X1    g13886(.A1(new_n14142_), .A2(new_n14026_), .Z(new_n14143_));
  AOI22_X1   g13887(.A1(new_n3864_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n3869_), .ZN(new_n14144_));
  OAI21_X1   g13888(.A1(new_n4886_), .A2(new_n5410_), .B(new_n14144_), .ZN(new_n14145_));
  AOI21_X1   g13889(.A1(new_n5351_), .A2(new_n3872_), .B(new_n14145_), .ZN(new_n14146_));
  XOR2_X1    g13890(.A1(new_n14146_), .A2(new_n3876_), .Z(new_n14147_));
  INV_X1     g13891(.I(new_n14147_), .ZN(new_n14148_));
  NAND2_X1   g13892(.A1(new_n14143_), .A2(new_n14148_), .ZN(new_n14149_));
  XNOR2_X1   g13893(.A1(new_n14142_), .A2(new_n14026_), .ZN(new_n14150_));
  NAND2_X1   g13894(.A1(new_n14150_), .A2(new_n14147_), .ZN(new_n14151_));
  NAND2_X1   g13895(.A1(new_n14151_), .A2(new_n14149_), .ZN(new_n14152_));
  XNOR2_X1   g13896(.A1(new_n14152_), .A2(new_n14024_), .ZN(new_n14153_));
  OAI22_X1   g13897(.A1(new_n6285_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n6284_), .ZN(new_n14154_));
  AOI21_X1   g13898(.A1(\b[39] ), .A2(new_n3456_), .B(new_n14154_), .ZN(new_n14155_));
  OAI21_X1   g13899(.A1(new_n6299_), .A2(new_n3261_), .B(new_n14155_), .ZN(new_n14156_));
  XOR2_X1    g13900(.A1(new_n14156_), .A2(\a[29] ), .Z(new_n14157_));
  NOR2_X1    g13901(.A1(new_n14153_), .A2(new_n14157_), .ZN(new_n14158_));
  XOR2_X1    g13902(.A1(new_n14152_), .A2(new_n14024_), .Z(new_n14159_));
  INV_X1     g13903(.I(new_n14157_), .ZN(new_n14160_));
  NOR2_X1    g13904(.A1(new_n14159_), .A2(new_n14160_), .ZN(new_n14161_));
  NOR2_X1    g13905(.A1(new_n14158_), .A2(new_n14161_), .ZN(new_n14162_));
  XOR2_X1    g13906(.A1(new_n14162_), .A2(new_n14021_), .Z(new_n14163_));
  AOI22_X1   g13907(.A1(new_n2716_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n2719_), .ZN(new_n14164_));
  OAI21_X1   g13908(.A1(new_n6490_), .A2(new_n2924_), .B(new_n14164_), .ZN(new_n14165_));
  AOI21_X1   g13909(.A1(new_n7906_), .A2(new_n2722_), .B(new_n14165_), .ZN(new_n14166_));
  XOR2_X1    g13910(.A1(new_n14166_), .A2(new_n2714_), .Z(new_n14167_));
  NOR2_X1    g13911(.A1(new_n14163_), .A2(new_n14167_), .ZN(new_n14168_));
  XNOR2_X1   g13912(.A1(new_n14162_), .A2(new_n14021_), .ZN(new_n14169_));
  INV_X1     g13913(.I(new_n14167_), .ZN(new_n14170_));
  NOR2_X1    g13914(.A1(new_n14169_), .A2(new_n14170_), .ZN(new_n14171_));
  NOR3_X1    g13915(.A1(new_n14171_), .A2(new_n14168_), .A3(new_n14019_), .ZN(new_n14172_));
  NAND2_X1   g13916(.A1(new_n14169_), .A2(new_n14170_), .ZN(new_n14173_));
  NAND2_X1   g13917(.A1(new_n14163_), .A2(new_n14167_), .ZN(new_n14174_));
  AOI21_X1   g13918(.A1(new_n14173_), .A2(new_n14174_), .B(new_n14018_), .ZN(new_n14175_));
  NOR2_X1    g13919(.A1(new_n14172_), .A2(new_n14175_), .ZN(new_n14176_));
  AOI22_X1   g13920(.A1(new_n2202_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n2205_), .ZN(new_n14177_));
  OAI21_X1   g13921(.A1(new_n7096_), .A2(new_n2370_), .B(new_n14177_), .ZN(new_n14178_));
  AOI21_X1   g13922(.A1(new_n7649_), .A2(new_n2208_), .B(new_n14178_), .ZN(new_n14179_));
  XOR2_X1    g13923(.A1(new_n14179_), .A2(new_n2200_), .Z(new_n14180_));
  NOR2_X1    g13924(.A1(new_n14176_), .A2(new_n14180_), .ZN(new_n14181_));
  NAND2_X1   g13925(.A1(new_n14176_), .A2(new_n14180_), .ZN(new_n14182_));
  INV_X1     g13926(.I(new_n14182_), .ZN(new_n14183_));
  NOR3_X1    g13927(.A1(new_n14183_), .A2(new_n14016_), .A3(new_n14181_), .ZN(new_n14184_));
  INV_X1     g13928(.I(new_n14016_), .ZN(new_n14185_));
  INV_X1     g13929(.I(new_n14181_), .ZN(new_n14186_));
  AOI21_X1   g13930(.A1(new_n14186_), .A2(new_n14182_), .B(new_n14185_), .ZN(new_n14187_));
  AOI22_X1   g13931(.A1(new_n1738_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n1743_), .ZN(new_n14188_));
  OAI21_X1   g13932(.A1(new_n8127_), .A2(new_n1931_), .B(new_n14188_), .ZN(new_n14189_));
  AOI21_X1   g13933(.A1(new_n9684_), .A2(new_n1746_), .B(new_n14189_), .ZN(new_n14190_));
  XOR2_X1    g13934(.A1(new_n14190_), .A2(new_n1736_), .Z(new_n14191_));
  INV_X1     g13935(.I(new_n14191_), .ZN(new_n14192_));
  OAI21_X1   g13936(.A1(new_n14187_), .A2(new_n14184_), .B(new_n14192_), .ZN(new_n14193_));
  NAND3_X1   g13937(.A1(new_n14186_), .A2(new_n14185_), .A3(new_n14182_), .ZN(new_n14194_));
  OAI21_X1   g13938(.A1(new_n14183_), .A2(new_n14181_), .B(new_n14016_), .ZN(new_n14195_));
  NAND3_X1   g13939(.A1(new_n14195_), .A2(new_n14194_), .A3(new_n14191_), .ZN(new_n14196_));
  NAND3_X1   g13940(.A1(new_n14193_), .A2(new_n14196_), .A3(new_n14014_), .ZN(new_n14197_));
  OAI21_X1   g13941(.A1(new_n13746_), .A2(new_n13906_), .B(new_n13900_), .ZN(new_n14198_));
  AOI21_X1   g13942(.A1(new_n14195_), .A2(new_n14194_), .B(new_n14191_), .ZN(new_n14199_));
  NOR3_X1    g13943(.A1(new_n14187_), .A2(new_n14184_), .A3(new_n14192_), .ZN(new_n14200_));
  OAI21_X1   g13944(.A1(new_n14199_), .A2(new_n14200_), .B(new_n14198_), .ZN(new_n14201_));
  NAND2_X1   g13945(.A1(new_n14201_), .A2(new_n14197_), .ZN(new_n14202_));
  OAI22_X1   g13946(.A1(new_n1592_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n1505_), .ZN(new_n14203_));
  AOI21_X1   g13947(.A1(\b[51] ), .A2(new_n1584_), .B(new_n14203_), .ZN(new_n14204_));
  OAI21_X1   g13948(.A1(new_n9385_), .A2(new_n1732_), .B(new_n14204_), .ZN(new_n14205_));
  XOR2_X1    g13949(.A1(new_n14205_), .A2(\a[17] ), .Z(new_n14206_));
  INV_X1     g13950(.I(new_n14206_), .ZN(new_n14207_));
  NAND2_X1   g13951(.A1(new_n14202_), .A2(new_n14207_), .ZN(new_n14208_));
  NOR3_X1    g13952(.A1(new_n14199_), .A2(new_n14200_), .A3(new_n14198_), .ZN(new_n14209_));
  AOI21_X1   g13953(.A1(new_n14193_), .A2(new_n14196_), .B(new_n14014_), .ZN(new_n14210_));
  NOR2_X1    g13954(.A1(new_n14209_), .A2(new_n14210_), .ZN(new_n14211_));
  NAND2_X1   g13955(.A1(new_n14211_), .A2(new_n14206_), .ZN(new_n14212_));
  NAND4_X1   g13956(.A1(new_n14212_), .A2(new_n14208_), .A3(new_n13914_), .A4(new_n14013_), .ZN(new_n14213_));
  NAND2_X1   g13957(.A1(new_n14013_), .A2(new_n13914_), .ZN(new_n14214_));
  NAND2_X1   g13958(.A1(new_n14212_), .A2(new_n14208_), .ZN(new_n14215_));
  NAND2_X1   g13959(.A1(new_n14215_), .A2(new_n14214_), .ZN(new_n14216_));
  OAI22_X1   g13960(.A1(new_n993_), .A2(new_n10308_), .B1(new_n9972_), .B2(new_n997_), .ZN(new_n14217_));
  AOI21_X1   g13961(.A1(\b[54] ), .A2(new_n1486_), .B(new_n14217_), .ZN(new_n14218_));
  OAI21_X1   g13962(.A1(new_n10319_), .A2(new_n1323_), .B(new_n14218_), .ZN(new_n14219_));
  XOR2_X1    g13963(.A1(new_n14219_), .A2(\a[14] ), .Z(new_n14220_));
  AOI21_X1   g13964(.A1(new_n14216_), .A2(new_n14213_), .B(new_n14220_), .ZN(new_n14221_));
  NAND2_X1   g13965(.A1(new_n14216_), .A2(new_n14213_), .ZN(new_n14222_));
  INV_X1     g13966(.I(new_n14220_), .ZN(new_n14223_));
  NOR2_X1    g13967(.A1(new_n14222_), .A2(new_n14223_), .ZN(new_n14224_));
  NOR2_X1    g13968(.A1(new_n14224_), .A2(new_n14221_), .ZN(new_n14225_));
  NAND2_X1   g13969(.A1(new_n14225_), .A2(new_n14012_), .ZN(new_n14226_));
  NOR2_X1    g13970(.A1(new_n14225_), .A2(new_n14012_), .ZN(new_n14227_));
  INV_X1     g13971(.I(new_n14227_), .ZN(new_n14228_));
  OAI22_X1   g13972(.A1(new_n713_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n717_), .ZN(new_n14229_));
  AOI21_X1   g13973(.A1(\b[57] ), .A2(new_n1126_), .B(new_n14229_), .ZN(new_n14230_));
  OAI21_X1   g13974(.A1(new_n12203_), .A2(new_n986_), .B(new_n14230_), .ZN(new_n14231_));
  XOR2_X1    g13975(.A1(new_n14231_), .A2(\a[11] ), .Z(new_n14232_));
  AOI21_X1   g13976(.A1(new_n14228_), .A2(new_n14226_), .B(new_n14232_), .ZN(new_n14233_));
  INV_X1     g13977(.I(new_n14226_), .ZN(new_n14234_));
  INV_X1     g13978(.I(new_n14232_), .ZN(new_n14235_));
  NOR3_X1    g13979(.A1(new_n14234_), .A2(new_n14227_), .A3(new_n14235_), .ZN(new_n14236_));
  NOR3_X1    g13980(.A1(new_n14233_), .A2(new_n14236_), .A3(new_n14010_), .ZN(new_n14237_));
  OAI21_X1   g13981(.A1(new_n14234_), .A2(new_n14227_), .B(new_n14235_), .ZN(new_n14238_));
  NAND3_X1   g13982(.A1(new_n14228_), .A2(new_n14226_), .A3(new_n14232_), .ZN(new_n14239_));
  AOI21_X1   g13983(.A1(new_n14238_), .A2(new_n14239_), .B(new_n14009_), .ZN(new_n14240_));
  NOR2_X1    g13984(.A1(new_n14240_), .A2(new_n14237_), .ZN(new_n14241_));
  INV_X1     g13985(.I(new_n13953_), .ZN(new_n14242_));
  OAI21_X1   g13986(.A1(new_n13954_), .A2(new_n13955_), .B(new_n13959_), .ZN(new_n14243_));
  AOI22_X1   g13987(.A1(new_n518_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n636_), .ZN(new_n14244_));
  OAI21_X1   g13988(.A1(new_n12147_), .A2(new_n917_), .B(new_n14244_), .ZN(new_n14245_));
  AOI21_X1   g13989(.A1(new_n13444_), .A2(new_n618_), .B(new_n14245_), .ZN(new_n14246_));
  XOR2_X1    g13990(.A1(new_n14246_), .A2(new_n488_), .Z(new_n14247_));
  AOI21_X1   g13991(.A1(new_n14243_), .A2(new_n14242_), .B(new_n14247_), .ZN(new_n14248_));
  NAND2_X1   g13992(.A1(new_n14243_), .A2(new_n14242_), .ZN(new_n14249_));
  INV_X1     g13993(.I(new_n14247_), .ZN(new_n14250_));
  NOR2_X1    g13994(.A1(new_n14249_), .A2(new_n14250_), .ZN(new_n14251_));
  NOR2_X1    g13995(.A1(new_n14251_), .A2(new_n14248_), .ZN(new_n14252_));
  XOR2_X1    g13996(.A1(new_n14252_), .A2(new_n14241_), .Z(new_n14253_));
  NAND2_X1   g13997(.A1(new_n14253_), .A2(new_n14008_), .ZN(new_n14254_));
  INV_X1     g13998(.I(new_n14241_), .ZN(new_n14255_));
  XOR2_X1    g13999(.A1(new_n14252_), .A2(new_n14255_), .Z(new_n14256_));
  NAND2_X1   g14000(.A1(new_n14256_), .A2(new_n14007_), .ZN(new_n14257_));
  NAND3_X1   g14001(.A1(new_n14257_), .A2(new_n14254_), .A3(new_n14004_), .ZN(new_n14258_));
  NOR2_X1    g14002(.A1(new_n14256_), .A2(new_n14007_), .ZN(new_n14259_));
  NOR2_X1    g14003(.A1(new_n14253_), .A2(new_n14008_), .ZN(new_n14260_));
  OAI21_X1   g14004(.A1(new_n14259_), .A2(new_n14260_), .B(new_n14003_), .ZN(new_n14261_));
  NAND2_X1   g14005(.A1(new_n14261_), .A2(new_n14258_), .ZN(new_n14262_));
  NAND2_X1   g14006(.A1(new_n14262_), .A2(new_n14001_), .ZN(new_n14263_));
  INV_X1     g14007(.I(new_n14001_), .ZN(new_n14264_));
  NOR3_X1    g14008(.A1(new_n14259_), .A2(new_n14260_), .A3(new_n14003_), .ZN(new_n14265_));
  AOI21_X1   g14009(.A1(new_n14257_), .A2(new_n14254_), .B(new_n14004_), .ZN(new_n14266_));
  NOR2_X1    g14010(.A1(new_n14266_), .A2(new_n14265_), .ZN(new_n14267_));
  NAND2_X1   g14011(.A1(new_n14267_), .A2(new_n14264_), .ZN(new_n14268_));
  NAND2_X1   g14012(.A1(new_n14268_), .A2(new_n14263_), .ZN(new_n14269_));
  XOR2_X1    g14013(.A1(new_n14269_), .A2(new_n14000_), .Z(\f[68] ));
  AOI21_X1   g14014(.A1(new_n14004_), .A2(new_n14254_), .B(new_n14260_), .ZN(new_n14271_));
  INV_X1     g14015(.I(new_n14248_), .ZN(new_n14272_));
  OAI21_X1   g14016(.A1(new_n14249_), .A2(new_n14250_), .B(new_n14255_), .ZN(new_n14273_));
  NAND2_X1   g14017(.A1(new_n14273_), .A2(new_n14272_), .ZN(new_n14274_));
  AOI21_X1   g14018(.A1(new_n14010_), .A2(new_n14239_), .B(new_n14233_), .ZN(new_n14275_));
  INV_X1     g14019(.I(new_n14275_), .ZN(new_n14276_));
  NOR2_X1    g14020(.A1(new_n14211_), .A2(new_n14206_), .ZN(new_n14277_));
  AOI21_X1   g14021(.A1(new_n14214_), .A2(new_n14212_), .B(new_n14277_), .ZN(new_n14278_));
  AOI21_X1   g14022(.A1(new_n14198_), .A2(new_n14196_), .B(new_n14199_), .ZN(new_n14279_));
  INV_X1     g14023(.I(new_n14279_), .ZN(new_n14280_));
  AOI21_X1   g14024(.A1(new_n14016_), .A2(new_n14182_), .B(new_n14181_), .ZN(new_n14281_));
  INV_X1     g14025(.I(new_n14281_), .ZN(new_n14282_));
  AOI21_X1   g14026(.A1(new_n14019_), .A2(new_n14174_), .B(new_n14168_), .ZN(new_n14283_));
  NOR2_X1    g14027(.A1(new_n14161_), .A2(new_n14021_), .ZN(new_n14284_));
  NOR2_X1    g14028(.A1(new_n14284_), .A2(new_n14158_), .ZN(new_n14285_));
  INV_X1     g14029(.I(new_n14151_), .ZN(new_n14286_));
  OAI21_X1   g14030(.A1(new_n14286_), .A2(new_n14024_), .B(new_n14149_), .ZN(new_n14287_));
  NOR2_X1    g14031(.A1(new_n14132_), .A2(new_n14137_), .ZN(new_n14288_));
  OAI21_X1   g14032(.A1(new_n14026_), .A2(new_n14288_), .B(new_n14138_), .ZN(new_n14289_));
  NOR2_X1    g14033(.A1(new_n14130_), .A2(new_n14139_), .ZN(new_n14290_));
  NOR2_X1    g14034(.A1(new_n14290_), .A2(new_n14127_), .ZN(new_n14291_));
  XOR2_X1    g14035(.A1(new_n14289_), .A2(new_n14291_), .Z(new_n14292_));
  NAND2_X1   g14036(.A1(new_n14120_), .A2(new_n14030_), .ZN(new_n14293_));
  NAND2_X1   g14037(.A1(new_n14293_), .A2(new_n14119_), .ZN(new_n14294_));
  NAND2_X1   g14038(.A1(new_n14112_), .A2(new_n14035_), .ZN(new_n14295_));
  NAND2_X1   g14039(.A1(new_n14295_), .A2(new_n14111_), .ZN(new_n14296_));
  INV_X1     g14040(.I(new_n14296_), .ZN(new_n14297_));
  INV_X1     g14041(.I(new_n14105_), .ZN(new_n14298_));
  AOI21_X1   g14042(.A1(new_n14038_), .A2(new_n14107_), .B(new_n14298_), .ZN(new_n14299_));
  INV_X1     g14043(.I(new_n14299_), .ZN(new_n14300_));
  INV_X1     g14044(.I(new_n14094_), .ZN(new_n14301_));
  OAI21_X1   g14045(.A1(new_n14041_), .A2(new_n14097_), .B(new_n14301_), .ZN(new_n14302_));
  NOR2_X1    g14046(.A1(new_n14086_), .A2(new_n14082_), .ZN(new_n14303_));
  AOI21_X1   g14047(.A1(new_n14044_), .A2(new_n14087_), .B(new_n14303_), .ZN(new_n14304_));
  INV_X1     g14048(.I(new_n14304_), .ZN(new_n14305_));
  NAND2_X1   g14049(.A1(new_n14076_), .A2(new_n14085_), .ZN(new_n14306_));
  NAND2_X1   g14050(.A1(new_n14306_), .A2(new_n14073_), .ZN(new_n14307_));
  NAND2_X1   g14051(.A1(new_n14057_), .A2(new_n14074_), .ZN(new_n14308_));
  AND2_X2    g14052(.A1(new_n14308_), .A2(new_n14055_), .Z(new_n14309_));
  AOI22_X1   g14053(.A1(new_n10981_), .A2(\b[12] ), .B1(new_n10979_), .B2(\b[11] ), .ZN(new_n14310_));
  OAI21_X1   g14054(.A1(new_n776_), .A2(new_n11306_), .B(new_n14310_), .ZN(new_n14311_));
  AOI21_X1   g14055(.A1(new_n1194_), .A2(new_n10984_), .B(new_n14311_), .ZN(new_n14312_));
  XOR2_X1    g14056(.A1(new_n14312_), .A2(new_n10989_), .Z(new_n14313_));
  INV_X1     g14057(.I(new_n14313_), .ZN(new_n14314_));
  AOI21_X1   g14058(.A1(new_n14062_), .A2(new_n14065_), .B(new_n14066_), .ZN(new_n14315_));
  AOI22_X1   g14059(.A1(new_n11926_), .A2(\b[9] ), .B1(new_n11924_), .B2(\b[8] ), .ZN(new_n14316_));
  OAI21_X1   g14060(.A1(new_n471_), .A2(new_n12317_), .B(new_n14316_), .ZN(new_n14317_));
  AOI21_X1   g14061(.A1(new_n676_), .A2(new_n11929_), .B(new_n14317_), .ZN(new_n14318_));
  XOR2_X1    g14062(.A1(new_n14318_), .A2(new_n12312_), .Z(new_n14319_));
  AOI22_X1   g14063(.A1(new_n12922_), .A2(\b[6] ), .B1(\b[5] ), .B2(new_n12923_), .ZN(new_n14320_));
  XNOR2_X1   g14064(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n14321_));
  XOR2_X1    g14065(.A1(new_n14320_), .A2(new_n14321_), .Z(new_n14322_));
  NAND2_X1   g14066(.A1(new_n14319_), .A2(new_n14322_), .ZN(new_n14323_));
  XOR2_X1    g14067(.A1(new_n14318_), .A2(\a[62] ), .Z(new_n14324_));
  INV_X1     g14068(.I(new_n14322_), .ZN(new_n14325_));
  NAND2_X1   g14069(.A1(new_n14324_), .A2(new_n14325_), .ZN(new_n14326_));
  NAND2_X1   g14070(.A1(new_n14323_), .A2(new_n14326_), .ZN(new_n14327_));
  XOR2_X1    g14071(.A1(new_n14327_), .A2(new_n14315_), .Z(new_n14328_));
  NOR2_X1    g14072(.A1(new_n14328_), .A2(new_n14314_), .ZN(new_n14329_));
  XNOR2_X1   g14073(.A1(new_n14327_), .A2(new_n14315_), .ZN(new_n14330_));
  NOR2_X1    g14074(.A1(new_n14330_), .A2(new_n14313_), .ZN(new_n14331_));
  NOR2_X1    g14075(.A1(new_n14331_), .A2(new_n14329_), .ZN(new_n14332_));
  XNOR2_X1   g14076(.A1(new_n14332_), .A2(new_n14309_), .ZN(new_n14333_));
  OAI22_X1   g14077(.A1(new_n11298_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n11297_), .ZN(new_n14334_));
  AOI21_X1   g14078(.A1(\b[13] ), .A2(new_n11296_), .B(new_n14334_), .ZN(new_n14335_));
  OAI21_X1   g14079(.A1(new_n1275_), .A2(new_n10069_), .B(new_n14335_), .ZN(new_n14336_));
  XOR2_X1    g14080(.A1(new_n14336_), .A2(\a[56] ), .Z(new_n14337_));
  INV_X1     g14081(.I(new_n14337_), .ZN(new_n14338_));
  NAND2_X1   g14082(.A1(new_n14333_), .A2(new_n14338_), .ZN(new_n14339_));
  XOR2_X1    g14083(.A1(new_n14332_), .A2(new_n14309_), .Z(new_n14340_));
  NAND2_X1   g14084(.A1(new_n14340_), .A2(new_n14337_), .ZN(new_n14341_));
  NAND2_X1   g14085(.A1(new_n14339_), .A2(new_n14341_), .ZN(new_n14342_));
  XOR2_X1    g14086(.A1(new_n14342_), .A2(new_n14307_), .Z(new_n14343_));
  AOI22_X1   g14087(.A1(new_n9125_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n9123_), .ZN(new_n14344_));
  OAI21_X1   g14088(.A1(new_n1296_), .A2(new_n9470_), .B(new_n14344_), .ZN(new_n14345_));
  AOI21_X1   g14089(.A1(new_n2038_), .A2(new_n9129_), .B(new_n14345_), .ZN(new_n14346_));
  XOR2_X1    g14090(.A1(new_n14346_), .A2(new_n9133_), .Z(new_n14347_));
  XOR2_X1    g14091(.A1(new_n14343_), .A2(new_n14347_), .Z(new_n14348_));
  XOR2_X1    g14092(.A1(new_n14348_), .A2(new_n14305_), .Z(new_n14349_));
  AOI22_X1   g14093(.A1(new_n8241_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n8246_), .ZN(new_n14350_));
  OAI21_X1   g14094(.A1(new_n1859_), .A2(new_n9114_), .B(new_n14350_), .ZN(new_n14351_));
  AOI21_X1   g14095(.A1(new_n2032_), .A2(new_n8252_), .B(new_n14351_), .ZN(new_n14352_));
  XOR2_X1    g14096(.A1(new_n14352_), .A2(\a[50] ), .Z(new_n14353_));
  NAND2_X1   g14097(.A1(new_n14349_), .A2(new_n14353_), .ZN(new_n14354_));
  OR2_X2     g14098(.A1(new_n14349_), .A2(new_n14353_), .Z(new_n14355_));
  NAND2_X1   g14099(.A1(new_n14355_), .A2(new_n14354_), .ZN(new_n14356_));
  XNOR2_X1   g14100(.A1(new_n14356_), .A2(new_n14302_), .ZN(new_n14357_));
  AOI22_X1   g14101(.A1(new_n7403_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n7408_), .ZN(new_n14358_));
  OAI21_X1   g14102(.A1(new_n2142_), .A2(new_n9488_), .B(new_n14358_), .ZN(new_n14359_));
  AOI21_X1   g14103(.A1(new_n3033_), .A2(new_n7414_), .B(new_n14359_), .ZN(new_n14360_));
  XOR2_X1    g14104(.A1(new_n14360_), .A2(new_n7410_), .Z(new_n14361_));
  INV_X1     g14105(.I(new_n14361_), .ZN(new_n14362_));
  NAND2_X1   g14106(.A1(new_n14357_), .A2(new_n14362_), .ZN(new_n14363_));
  XOR2_X1    g14107(.A1(new_n14356_), .A2(new_n14302_), .Z(new_n14364_));
  NAND2_X1   g14108(.A1(new_n14364_), .A2(new_n14361_), .ZN(new_n14365_));
  NAND2_X1   g14109(.A1(new_n14363_), .A2(new_n14365_), .ZN(new_n14366_));
  XOR2_X1    g14110(.A1(new_n14366_), .A2(new_n14300_), .Z(new_n14367_));
  OAI22_X1   g14111(.A1(new_n7730_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n7731_), .ZN(new_n14368_));
  AOI21_X1   g14112(.A1(\b[25] ), .A2(new_n6887_), .B(new_n14368_), .ZN(new_n14369_));
  OAI21_X1   g14113(.A1(new_n3165_), .A2(new_n7728_), .B(new_n14369_), .ZN(new_n14370_));
  XOR2_X1    g14114(.A1(new_n14370_), .A2(\a[44] ), .Z(new_n14371_));
  NOR2_X1    g14115(.A1(new_n14367_), .A2(new_n14371_), .ZN(new_n14372_));
  XOR2_X1    g14116(.A1(new_n14366_), .A2(new_n14299_), .Z(new_n14373_));
  INV_X1     g14117(.I(new_n14371_), .ZN(new_n14374_));
  NOR2_X1    g14118(.A1(new_n14373_), .A2(new_n14374_), .ZN(new_n14375_));
  NOR2_X1    g14119(.A1(new_n14372_), .A2(new_n14375_), .ZN(new_n14376_));
  XOR2_X1    g14120(.A1(new_n14376_), .A2(new_n14297_), .Z(new_n14377_));
  AOI22_X1   g14121(.A1(new_n6108_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n6111_), .ZN(new_n14378_));
  OAI21_X1   g14122(.A1(new_n3185_), .A2(new_n7708_), .B(new_n14378_), .ZN(new_n14379_));
  AOI21_X1   g14123(.A1(new_n4230_), .A2(new_n6105_), .B(new_n14379_), .ZN(new_n14380_));
  XOR2_X1    g14124(.A1(new_n14380_), .A2(new_n5849_), .Z(new_n14381_));
  NOR2_X1    g14125(.A1(new_n14377_), .A2(new_n14381_), .ZN(new_n14382_));
  INV_X1     g14126(.I(new_n14382_), .ZN(new_n14383_));
  NAND2_X1   g14127(.A1(new_n14377_), .A2(new_n14381_), .ZN(new_n14384_));
  NAND2_X1   g14128(.A1(new_n14383_), .A2(new_n14384_), .ZN(new_n14385_));
  XNOR2_X1   g14129(.A1(new_n14385_), .A2(new_n14294_), .ZN(new_n14386_));
  AOI22_X1   g14130(.A1(new_n5155_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n5160_), .ZN(new_n14387_));
  OAI21_X1   g14131(.A1(new_n4022_), .A2(new_n6877_), .B(new_n14387_), .ZN(new_n14388_));
  AOI21_X1   g14132(.A1(new_n4223_), .A2(new_n5166_), .B(new_n14388_), .ZN(new_n14389_));
  XOR2_X1    g14133(.A1(new_n14389_), .A2(new_n5162_), .Z(new_n14390_));
  INV_X1     g14134(.I(new_n14390_), .ZN(new_n14391_));
  NAND2_X1   g14135(.A1(new_n14386_), .A2(new_n14391_), .ZN(new_n14392_));
  NOR2_X1    g14136(.A1(new_n14386_), .A2(new_n14391_), .ZN(new_n14393_));
  INV_X1     g14137(.I(new_n14393_), .ZN(new_n14394_));
  NAND2_X1   g14138(.A1(new_n14394_), .A2(new_n14392_), .ZN(new_n14395_));
  AOI22_X1   g14139(.A1(new_n4918_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n4921_), .ZN(new_n14396_));
  OAI21_X1   g14140(.A1(new_n4639_), .A2(new_n6099_), .B(new_n14396_), .ZN(new_n14397_));
  AOI21_X1   g14141(.A1(new_n5594_), .A2(new_n4699_), .B(new_n14397_), .ZN(new_n14398_));
  XOR2_X1    g14142(.A1(new_n14398_), .A2(new_n4446_), .Z(new_n14399_));
  INV_X1     g14143(.I(new_n14399_), .ZN(new_n14400_));
  XOR2_X1    g14144(.A1(new_n14395_), .A2(new_n14400_), .Z(new_n14401_));
  XNOR2_X1   g14145(.A1(new_n14292_), .A2(new_n14401_), .ZN(new_n14402_));
  AOI22_X1   g14146(.A1(new_n3864_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n3869_), .ZN(new_n14403_));
  OAI21_X1   g14147(.A1(new_n5312_), .A2(new_n5410_), .B(new_n14403_), .ZN(new_n14404_));
  AOI21_X1   g14148(.A1(new_n6310_), .A2(new_n3872_), .B(new_n14404_), .ZN(new_n14405_));
  XOR2_X1    g14149(.A1(new_n14405_), .A2(new_n3876_), .Z(new_n14406_));
  XNOR2_X1   g14150(.A1(new_n14402_), .A2(new_n14406_), .ZN(new_n14407_));
  XOR2_X1    g14151(.A1(new_n14407_), .A2(new_n14287_), .Z(new_n14408_));
  AOI22_X1   g14152(.A1(new_n3267_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n3270_), .ZN(new_n14409_));
  OAI21_X1   g14153(.A1(new_n6284_), .A2(new_n3475_), .B(new_n14409_), .ZN(new_n14410_));
  AOI21_X1   g14154(.A1(new_n7106_), .A2(new_n3273_), .B(new_n14410_), .ZN(new_n14411_));
  XOR2_X1    g14155(.A1(new_n14411_), .A2(new_n3264_), .Z(new_n14412_));
  NOR2_X1    g14156(.A1(new_n14408_), .A2(new_n14412_), .ZN(new_n14413_));
  AND2_X2    g14157(.A1(new_n14408_), .A2(new_n14412_), .Z(new_n14414_));
  NOR2_X1    g14158(.A1(new_n14414_), .A2(new_n14413_), .ZN(new_n14415_));
  XNOR2_X1   g14159(.A1(new_n14415_), .A2(new_n14285_), .ZN(new_n14416_));
  AOI22_X1   g14160(.A1(new_n2716_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n2719_), .ZN(new_n14417_));
  OAI21_X1   g14161(.A1(new_n6775_), .A2(new_n2924_), .B(new_n14417_), .ZN(new_n14418_));
  AOI21_X1   g14162(.A1(new_n7926_), .A2(new_n2722_), .B(new_n14418_), .ZN(new_n14419_));
  XOR2_X1    g14163(.A1(new_n14419_), .A2(\a[26] ), .Z(new_n14420_));
  NAND2_X1   g14164(.A1(new_n14416_), .A2(new_n14420_), .ZN(new_n14421_));
  OR2_X2     g14165(.A1(new_n14416_), .A2(new_n14420_), .Z(new_n14422_));
  AOI21_X1   g14166(.A1(new_n14422_), .A2(new_n14421_), .B(new_n14283_), .ZN(new_n14423_));
  AND3_X2    g14167(.A1(new_n14422_), .A2(new_n14283_), .A3(new_n14421_), .Z(new_n14424_));
  AOI22_X1   g14168(.A1(new_n2202_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n2205_), .ZN(new_n14425_));
  OAI21_X1   g14169(.A1(new_n7617_), .A2(new_n2370_), .B(new_n14425_), .ZN(new_n14426_));
  AOI21_X1   g14170(.A1(new_n8792_), .A2(new_n2208_), .B(new_n14426_), .ZN(new_n14427_));
  XOR2_X1    g14171(.A1(new_n14427_), .A2(new_n2200_), .Z(new_n14428_));
  INV_X1     g14172(.I(new_n14428_), .ZN(new_n14429_));
  OAI21_X1   g14173(.A1(new_n14424_), .A2(new_n14423_), .B(new_n14429_), .ZN(new_n14430_));
  INV_X1     g14174(.I(new_n14430_), .ZN(new_n14431_));
  NOR3_X1    g14175(.A1(new_n14424_), .A2(new_n14423_), .A3(new_n14429_), .ZN(new_n14432_));
  NOR3_X1    g14176(.A1(new_n14431_), .A2(new_n14282_), .A3(new_n14432_), .ZN(new_n14433_));
  INV_X1     g14177(.I(new_n14433_), .ZN(new_n14434_));
  OAI21_X1   g14178(.A1(new_n14431_), .A2(new_n14432_), .B(new_n14282_), .ZN(new_n14435_));
  AOI22_X1   g14179(.A1(new_n1738_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n1743_), .ZN(new_n14436_));
  OAI21_X1   g14180(.A1(new_n8168_), .A2(new_n1931_), .B(new_n14436_), .ZN(new_n14437_));
  AOI21_X1   g14181(.A1(new_n8783_), .A2(new_n1746_), .B(new_n14437_), .ZN(new_n14438_));
  XOR2_X1    g14182(.A1(new_n14438_), .A2(new_n1736_), .Z(new_n14439_));
  AOI21_X1   g14183(.A1(new_n14434_), .A2(new_n14435_), .B(new_n14439_), .ZN(new_n14440_));
  INV_X1     g14184(.I(new_n14435_), .ZN(new_n14441_));
  INV_X1     g14185(.I(new_n14439_), .ZN(new_n14442_));
  NOR3_X1    g14186(.A1(new_n14441_), .A2(new_n14433_), .A3(new_n14442_), .ZN(new_n14443_));
  NOR3_X1    g14187(.A1(new_n14440_), .A2(new_n14443_), .A3(new_n14280_), .ZN(new_n14444_));
  OAI21_X1   g14188(.A1(new_n14441_), .A2(new_n14433_), .B(new_n14442_), .ZN(new_n14445_));
  NAND3_X1   g14189(.A1(new_n14434_), .A2(new_n14435_), .A3(new_n14439_), .ZN(new_n14446_));
  AOI21_X1   g14190(.A1(new_n14445_), .A2(new_n14446_), .B(new_n14279_), .ZN(new_n14447_));
  OAI22_X1   g14191(.A1(new_n1592_), .A2(new_n9942_), .B1(new_n9376_), .B2(new_n1505_), .ZN(new_n14448_));
  AOI21_X1   g14192(.A1(\b[52] ), .A2(new_n1584_), .B(new_n14448_), .ZN(new_n14449_));
  OAI21_X1   g14193(.A1(new_n9952_), .A2(new_n1732_), .B(new_n14449_), .ZN(new_n14450_));
  XOR2_X1    g14194(.A1(new_n14450_), .A2(\a[17] ), .Z(new_n14451_));
  INV_X1     g14195(.I(new_n14451_), .ZN(new_n14452_));
  OAI21_X1   g14196(.A1(new_n14444_), .A2(new_n14447_), .B(new_n14452_), .ZN(new_n14453_));
  NAND3_X1   g14197(.A1(new_n14445_), .A2(new_n14446_), .A3(new_n14279_), .ZN(new_n14454_));
  OAI21_X1   g14198(.A1(new_n14440_), .A2(new_n14443_), .B(new_n14280_), .ZN(new_n14455_));
  NAND3_X1   g14199(.A1(new_n14455_), .A2(new_n14454_), .A3(new_n14451_), .ZN(new_n14456_));
  NAND2_X1   g14200(.A1(new_n14453_), .A2(new_n14456_), .ZN(new_n14457_));
  XOR2_X1    g14201(.A1(new_n14457_), .A2(new_n14278_), .Z(new_n14458_));
  INV_X1     g14202(.I(new_n14221_), .ZN(new_n14459_));
  OAI21_X1   g14203(.A1(new_n14222_), .A2(new_n14223_), .B(new_n14011_), .ZN(new_n14460_));
  NAND2_X1   g14204(.A1(new_n14460_), .A2(new_n14459_), .ZN(new_n14461_));
  OAI22_X1   g14205(.A1(new_n993_), .A2(new_n10625_), .B1(new_n10308_), .B2(new_n997_), .ZN(new_n14462_));
  AOI21_X1   g14206(.A1(\b[55] ), .A2(new_n1486_), .B(new_n14462_), .ZN(new_n14463_));
  OAI21_X1   g14207(.A1(new_n13693_), .A2(new_n1323_), .B(new_n14463_), .ZN(new_n14464_));
  XOR2_X1    g14208(.A1(new_n14464_), .A2(\a[14] ), .Z(new_n14465_));
  INV_X1     g14209(.I(new_n14465_), .ZN(new_n14466_));
  NAND2_X1   g14210(.A1(new_n14461_), .A2(new_n14466_), .ZN(new_n14467_));
  NOR2_X1    g14211(.A1(new_n14461_), .A2(new_n14466_), .ZN(new_n14468_));
  INV_X1     g14212(.I(new_n14468_), .ZN(new_n14469_));
  NAND2_X1   g14213(.A1(new_n14469_), .A2(new_n14467_), .ZN(new_n14470_));
  NOR2_X1    g14214(.A1(new_n14470_), .A2(new_n14458_), .ZN(new_n14471_));
  INV_X1     g14215(.I(new_n14278_), .ZN(new_n14472_));
  XOR2_X1    g14216(.A1(new_n14457_), .A2(new_n14472_), .Z(new_n14473_));
  AOI21_X1   g14217(.A1(new_n14467_), .A2(new_n14469_), .B(new_n14473_), .ZN(new_n14474_));
  OAI22_X1   g14218(.A1(new_n713_), .A2(new_n12147_), .B1(new_n12151_), .B2(new_n717_), .ZN(new_n14475_));
  AOI21_X1   g14219(.A1(\b[58] ), .A2(new_n1126_), .B(new_n14475_), .ZN(new_n14476_));
  OAI21_X1   g14220(.A1(new_n11840_), .A2(new_n986_), .B(new_n14476_), .ZN(new_n14477_));
  XOR2_X1    g14221(.A1(new_n14477_), .A2(\a[11] ), .Z(new_n14478_));
  INV_X1     g14222(.I(new_n14478_), .ZN(new_n14479_));
  OAI21_X1   g14223(.A1(new_n14474_), .A2(new_n14471_), .B(new_n14479_), .ZN(new_n14480_));
  INV_X1     g14224(.I(new_n14480_), .ZN(new_n14481_));
  NOR3_X1    g14225(.A1(new_n14474_), .A2(new_n14471_), .A3(new_n14479_), .ZN(new_n14482_));
  NOR3_X1    g14226(.A1(new_n14481_), .A2(new_n14482_), .A3(new_n14276_), .ZN(new_n14483_));
  OR3_X2     g14227(.A1(new_n14474_), .A2(new_n14471_), .A3(new_n14479_), .Z(new_n14484_));
  AOI21_X1   g14228(.A1(new_n14484_), .A2(new_n14480_), .B(new_n14275_), .ZN(new_n14485_));
  AOI22_X1   g14229(.A1(new_n518_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n636_), .ZN(new_n14486_));
  OAI21_X1   g14230(.A1(new_n12148_), .A2(new_n917_), .B(new_n14486_), .ZN(new_n14487_));
  AOI21_X1   g14231(.A1(new_n12811_), .A2(new_n618_), .B(new_n14487_), .ZN(new_n14488_));
  XOR2_X1    g14232(.A1(new_n14488_), .A2(new_n488_), .Z(new_n14489_));
  INV_X1     g14233(.I(new_n14489_), .ZN(new_n14490_));
  OAI21_X1   g14234(.A1(new_n14483_), .A2(new_n14485_), .B(new_n14490_), .ZN(new_n14491_));
  NAND3_X1   g14235(.A1(new_n14484_), .A2(new_n14275_), .A3(new_n14480_), .ZN(new_n14492_));
  OAI21_X1   g14236(.A1(new_n14481_), .A2(new_n14482_), .B(new_n14276_), .ZN(new_n14493_));
  NAND3_X1   g14237(.A1(new_n14493_), .A2(new_n14492_), .A3(new_n14489_), .ZN(new_n14494_));
  NAND2_X1   g14238(.A1(new_n14491_), .A2(new_n14494_), .ZN(new_n14495_));
  XOR2_X1    g14239(.A1(new_n14495_), .A2(new_n14274_), .Z(new_n14496_));
  XOR2_X1    g14240(.A1(new_n14496_), .A2(new_n14271_), .Z(new_n14497_));
  NOR2_X1    g14241(.A1(new_n14262_), .A2(new_n14001_), .ZN(new_n14498_));
  AOI21_X1   g14242(.A1(new_n14000_), .A2(new_n14263_), .B(new_n14498_), .ZN(new_n14499_));
  XOR2_X1    g14243(.A1(new_n14499_), .A2(new_n14497_), .Z(\f[69] ));
  AOI21_X1   g14244(.A1(new_n14276_), .A2(new_n14484_), .B(new_n14481_), .ZN(new_n14501_));
  INV_X1     g14245(.I(new_n14467_), .ZN(new_n14502_));
  AOI21_X1   g14246(.A1(new_n14458_), .A2(new_n14469_), .B(new_n14502_), .ZN(new_n14503_));
  INV_X1     g14247(.I(new_n14503_), .ZN(new_n14504_));
  NAND2_X1   g14248(.A1(new_n14456_), .A2(new_n14472_), .ZN(new_n14505_));
  NAND2_X1   g14249(.A1(new_n14505_), .A2(new_n14453_), .ZN(new_n14506_));
  OAI21_X1   g14250(.A1(new_n14279_), .A2(new_n14443_), .B(new_n14445_), .ZN(new_n14507_));
  OAI21_X1   g14251(.A1(new_n14281_), .A2(new_n14432_), .B(new_n14430_), .ZN(new_n14508_));
  INV_X1     g14252(.I(new_n14283_), .ZN(new_n14509_));
  INV_X1     g14253(.I(new_n14421_), .ZN(new_n14510_));
  AOI21_X1   g14254(.A1(new_n14509_), .A2(new_n14422_), .B(new_n14510_), .ZN(new_n14511_));
  NOR2_X1    g14255(.A1(new_n14414_), .A2(new_n14285_), .ZN(new_n14512_));
  NOR2_X1    g14256(.A1(new_n14512_), .A2(new_n14413_), .ZN(new_n14513_));
  NOR2_X1    g14257(.A1(new_n14402_), .A2(new_n14406_), .ZN(new_n14514_));
  NAND2_X1   g14258(.A1(new_n14402_), .A2(new_n14406_), .ZN(new_n14515_));
  AOI21_X1   g14259(.A1(new_n14287_), .A2(new_n14515_), .B(new_n14514_), .ZN(new_n14516_));
  NAND2_X1   g14260(.A1(new_n14289_), .A2(new_n14400_), .ZN(new_n14517_));
  XOR2_X1    g14261(.A1(new_n14395_), .A2(new_n14291_), .Z(new_n14518_));
  OAI21_X1   g14262(.A1(new_n14289_), .A2(new_n14400_), .B(new_n14518_), .ZN(new_n14519_));
  NAND2_X1   g14263(.A1(new_n14519_), .A2(new_n14517_), .ZN(new_n14520_));
  OAI21_X1   g14264(.A1(new_n14291_), .A2(new_n14393_), .B(new_n14392_), .ZN(new_n14521_));
  AOI22_X1   g14265(.A1(new_n5155_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n5160_), .ZN(new_n14522_));
  OAI21_X1   g14266(.A1(new_n4023_), .A2(new_n6877_), .B(new_n14522_), .ZN(new_n14523_));
  AOI21_X1   g14267(.A1(new_n5103_), .A2(new_n5166_), .B(new_n14523_), .ZN(new_n14524_));
  XOR2_X1    g14268(.A1(new_n14524_), .A2(new_n5162_), .Z(new_n14525_));
  AOI21_X1   g14269(.A1(new_n14294_), .A2(new_n14384_), .B(new_n14382_), .ZN(new_n14526_));
  NOR2_X1    g14270(.A1(new_n14375_), .A2(new_n14297_), .ZN(new_n14527_));
  NOR2_X1    g14271(.A1(new_n14527_), .A2(new_n14372_), .ZN(new_n14528_));
  AOI22_X1   g14272(.A1(new_n6569_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n6574_), .ZN(new_n14529_));
  OAI21_X1   g14273(.A1(new_n3006_), .A2(new_n8565_), .B(new_n14529_), .ZN(new_n14530_));
  AOI21_X1   g14274(.A1(new_n3807_), .A2(new_n6579_), .B(new_n14530_), .ZN(new_n14531_));
  XOR2_X1    g14275(.A1(new_n14531_), .A2(new_n6567_), .Z(new_n14532_));
  NAND2_X1   g14276(.A1(new_n14365_), .A2(new_n14300_), .ZN(new_n14533_));
  NAND2_X1   g14277(.A1(new_n14533_), .A2(new_n14363_), .ZN(new_n14534_));
  INV_X1     g14278(.I(new_n14354_), .ZN(new_n14535_));
  AOI21_X1   g14279(.A1(new_n14302_), .A2(new_n14355_), .B(new_n14535_), .ZN(new_n14536_));
  NOR2_X1    g14280(.A1(new_n14343_), .A2(new_n14347_), .ZN(new_n14537_));
  AOI21_X1   g14281(.A1(new_n14343_), .A2(new_n14347_), .B(new_n14304_), .ZN(new_n14538_));
  NOR2_X1    g14282(.A1(new_n14538_), .A2(new_n14537_), .ZN(new_n14539_));
  AOI22_X1   g14283(.A1(new_n8241_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n8246_), .ZN(new_n14540_));
  OAI21_X1   g14284(.A1(new_n1860_), .A2(new_n9114_), .B(new_n14540_), .ZN(new_n14541_));
  AOI21_X1   g14285(.A1(new_n2659_), .A2(new_n8252_), .B(new_n14541_), .ZN(new_n14542_));
  XOR2_X1    g14286(.A1(new_n14542_), .A2(new_n8248_), .Z(new_n14543_));
  AOI22_X1   g14287(.A1(new_n10064_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n10062_), .ZN(new_n14544_));
  OAI21_X1   g14288(.A1(new_n1093_), .A2(new_n10399_), .B(new_n14544_), .ZN(new_n14545_));
  AOI21_X1   g14289(.A1(new_n1701_), .A2(new_n10068_), .B(new_n14545_), .ZN(new_n14546_));
  XOR2_X1    g14290(.A1(new_n14546_), .A2(new_n10057_), .Z(new_n14547_));
  INV_X1     g14291(.I(new_n14323_), .ZN(new_n14548_));
  OAI21_X1   g14292(.A1(new_n14548_), .A2(new_n14315_), .B(new_n14326_), .ZN(new_n14549_));
  AOI22_X1   g14293(.A1(new_n11926_), .A2(\b[10] ), .B1(new_n11924_), .B2(\b[9] ), .ZN(new_n14550_));
  OAI21_X1   g14294(.A1(new_n577_), .A2(new_n12317_), .B(new_n14550_), .ZN(new_n14551_));
  AOI21_X1   g14295(.A1(new_n1059_), .A2(new_n11929_), .B(new_n14551_), .ZN(new_n14552_));
  XOR2_X1    g14296(.A1(new_n14552_), .A2(new_n12312_), .Z(new_n14553_));
  OAI21_X1   g14297(.A1(\a[2] ), .A2(\a[5] ), .B(new_n14320_), .ZN(new_n14554_));
  OAI21_X1   g14298(.A1(new_n270_), .A2(new_n312_), .B(new_n14554_), .ZN(new_n14555_));
  AOI22_X1   g14299(.A1(new_n12922_), .A2(\b[7] ), .B1(\b[6] ), .B2(new_n12923_), .ZN(new_n14556_));
  INV_X1     g14300(.I(new_n14556_), .ZN(new_n14557_));
  NOR2_X1    g14301(.A1(new_n14555_), .A2(new_n14557_), .ZN(new_n14558_));
  NAND2_X1   g14302(.A1(new_n14555_), .A2(new_n14557_), .ZN(new_n14559_));
  INV_X1     g14303(.I(new_n14559_), .ZN(new_n14560_));
  NOR2_X1    g14304(.A1(new_n14560_), .A2(new_n14558_), .ZN(new_n14561_));
  XNOR2_X1   g14305(.A1(new_n14553_), .A2(new_n14561_), .ZN(new_n14562_));
  INV_X1     g14306(.I(new_n14562_), .ZN(new_n14563_));
  OAI22_X1   g14307(.A1(new_n12306_), .A2(new_n1070_), .B1(new_n12305_), .B2(new_n941_), .ZN(new_n14564_));
  AOI21_X1   g14308(.A1(\b[11] ), .A2(new_n12304_), .B(new_n14564_), .ZN(new_n14565_));
  OAI21_X1   g14309(.A1(new_n1082_), .A2(new_n10985_), .B(new_n14565_), .ZN(new_n14566_));
  XOR2_X1    g14310(.A1(new_n14566_), .A2(\a[59] ), .Z(new_n14567_));
  NOR2_X1    g14311(.A1(new_n14567_), .A2(new_n14563_), .ZN(new_n14568_));
  XOR2_X1    g14312(.A1(new_n14566_), .A2(new_n10989_), .Z(new_n14569_));
  NOR2_X1    g14313(.A1(new_n14569_), .A2(new_n14562_), .ZN(new_n14570_));
  OR2_X2     g14314(.A1(new_n14568_), .A2(new_n14570_), .Z(new_n14571_));
  XNOR2_X1   g14315(.A1(new_n14571_), .A2(new_n14549_), .ZN(new_n14572_));
  INV_X1     g14316(.I(new_n14331_), .ZN(new_n14573_));
  OAI21_X1   g14317(.A1(new_n14309_), .A2(new_n14329_), .B(new_n14573_), .ZN(new_n14574_));
  NAND2_X1   g14318(.A1(new_n14572_), .A2(new_n14574_), .ZN(new_n14575_));
  XOR2_X1    g14319(.A1(new_n14571_), .A2(new_n14549_), .Z(new_n14576_));
  INV_X1     g14320(.I(new_n14574_), .ZN(new_n14577_));
  NAND2_X1   g14321(.A1(new_n14576_), .A2(new_n14577_), .ZN(new_n14578_));
  NAND2_X1   g14322(.A1(new_n14575_), .A2(new_n14578_), .ZN(new_n14579_));
  XOR2_X1    g14323(.A1(new_n14579_), .A2(new_n14547_), .Z(new_n14580_));
  NAND2_X1   g14324(.A1(new_n14341_), .A2(new_n14307_), .ZN(new_n14581_));
  NAND2_X1   g14325(.A1(new_n14581_), .A2(new_n14339_), .ZN(new_n14582_));
  AOI22_X1   g14326(.A1(new_n9125_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n9123_), .ZN(new_n14583_));
  OAI21_X1   g14327(.A1(new_n1432_), .A2(new_n9470_), .B(new_n14583_), .ZN(new_n14584_));
  AOI21_X1   g14328(.A1(new_n1695_), .A2(new_n9129_), .B(new_n14584_), .ZN(new_n14585_));
  XOR2_X1    g14329(.A1(new_n14585_), .A2(\a[53] ), .Z(new_n14586_));
  NAND2_X1   g14330(.A1(new_n14582_), .A2(new_n14586_), .ZN(new_n14587_));
  OR2_X2     g14331(.A1(new_n14582_), .A2(new_n14586_), .Z(new_n14588_));
  NAND2_X1   g14332(.A1(new_n14588_), .A2(new_n14587_), .ZN(new_n14589_));
  XOR2_X1    g14333(.A1(new_n14589_), .A2(new_n14580_), .Z(new_n14590_));
  NOR2_X1    g14334(.A1(new_n14590_), .A2(new_n14543_), .ZN(new_n14591_));
  INV_X1     g14335(.I(new_n14543_), .ZN(new_n14592_));
  XNOR2_X1   g14336(.A1(new_n14589_), .A2(new_n14580_), .ZN(new_n14593_));
  NOR2_X1    g14337(.A1(new_n14593_), .A2(new_n14592_), .ZN(new_n14594_));
  NOR2_X1    g14338(.A1(new_n14594_), .A2(new_n14591_), .ZN(new_n14595_));
  NAND2_X1   g14339(.A1(new_n14595_), .A2(new_n14539_), .ZN(new_n14596_));
  OAI22_X1   g14340(.A1(new_n14594_), .A2(new_n14591_), .B1(new_n14537_), .B2(new_n14538_), .ZN(new_n14597_));
  AND2_X2    g14341(.A1(new_n14596_), .A2(new_n14597_), .Z(new_n14598_));
  OAI22_X1   g14342(.A1(new_n2495_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n2646_), .ZN(new_n14599_));
  AOI21_X1   g14343(.A1(\b[23] ), .A2(new_n7719_), .B(new_n14599_), .ZN(new_n14600_));
  OAI21_X1   g14344(.A1(new_n2655_), .A2(new_n8585_), .B(new_n14600_), .ZN(new_n14601_));
  XOR2_X1    g14345(.A1(new_n14601_), .A2(\a[47] ), .Z(new_n14602_));
  NOR2_X1    g14346(.A1(new_n14598_), .A2(new_n14602_), .ZN(new_n14603_));
  AND3_X2    g14347(.A1(new_n14596_), .A2(new_n14597_), .A3(new_n14602_), .Z(new_n14604_));
  NOR2_X1    g14348(.A1(new_n14603_), .A2(new_n14604_), .ZN(new_n14605_));
  XOR2_X1    g14349(.A1(new_n14605_), .A2(new_n14536_), .Z(new_n14606_));
  XOR2_X1    g14350(.A1(new_n14534_), .A2(new_n14606_), .Z(new_n14607_));
  XOR2_X1    g14351(.A1(new_n14607_), .A2(new_n14532_), .Z(new_n14608_));
  AOI22_X1   g14352(.A1(new_n6108_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n6111_), .ZN(new_n14609_));
  OAI21_X1   g14353(.A1(new_n3592_), .A2(new_n7708_), .B(new_n14609_), .ZN(new_n14610_));
  AOI21_X1   g14354(.A1(new_n3796_), .A2(new_n6105_), .B(new_n14610_), .ZN(new_n14611_));
  XOR2_X1    g14355(.A1(new_n14611_), .A2(new_n5849_), .Z(new_n14612_));
  INV_X1     g14356(.I(new_n14612_), .ZN(new_n14613_));
  NAND2_X1   g14357(.A1(new_n14608_), .A2(new_n14613_), .ZN(new_n14614_));
  INV_X1     g14358(.I(new_n14532_), .ZN(new_n14615_));
  XOR2_X1    g14359(.A1(new_n14607_), .A2(new_n14615_), .Z(new_n14616_));
  NAND2_X1   g14360(.A1(new_n14616_), .A2(new_n14612_), .ZN(new_n14617_));
  NAND2_X1   g14361(.A1(new_n14614_), .A2(new_n14617_), .ZN(new_n14618_));
  NOR2_X1    g14362(.A1(new_n14618_), .A2(new_n14528_), .ZN(new_n14619_));
  INV_X1     g14363(.I(new_n14528_), .ZN(new_n14620_));
  AOI21_X1   g14364(.A1(new_n14614_), .A2(new_n14617_), .B(new_n14620_), .ZN(new_n14621_));
  OAI21_X1   g14365(.A1(new_n14619_), .A2(new_n14621_), .B(new_n14526_), .ZN(new_n14622_));
  OR3_X2     g14366(.A1(new_n14526_), .A2(new_n14619_), .A3(new_n14621_), .Z(new_n14623_));
  NAND2_X1   g14367(.A1(new_n14623_), .A2(new_n14622_), .ZN(new_n14624_));
  XOR2_X1    g14368(.A1(new_n14624_), .A2(new_n14525_), .Z(new_n14625_));
  OAI22_X1   g14369(.A1(new_n5312_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n4886_), .ZN(new_n14626_));
  AOI21_X1   g14370(.A1(\b[35] ), .A2(new_n4706_), .B(new_n14626_), .ZN(new_n14627_));
  OAI21_X1   g14371(.A1(new_n5322_), .A2(new_n4458_), .B(new_n14627_), .ZN(new_n14628_));
  XOR2_X1    g14372(.A1(new_n14628_), .A2(\a[35] ), .Z(new_n14629_));
  INV_X1     g14373(.I(new_n14629_), .ZN(new_n14630_));
  NAND2_X1   g14374(.A1(new_n14625_), .A2(new_n14630_), .ZN(new_n14631_));
  INV_X1     g14375(.I(new_n14525_), .ZN(new_n14632_));
  XOR2_X1    g14376(.A1(new_n14624_), .A2(new_n14632_), .Z(new_n14633_));
  NAND2_X1   g14377(.A1(new_n14633_), .A2(new_n14629_), .ZN(new_n14634_));
  NAND2_X1   g14378(.A1(new_n14631_), .A2(new_n14634_), .ZN(new_n14635_));
  XNOR2_X1   g14379(.A1(new_n14635_), .A2(new_n14521_), .ZN(new_n14636_));
  AOI22_X1   g14380(.A1(new_n3864_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n3869_), .ZN(new_n14637_));
  OAI21_X1   g14381(.A1(new_n5341_), .A2(new_n5410_), .B(new_n14637_), .ZN(new_n14638_));
  AOI21_X1   g14382(.A1(new_n5793_), .A2(new_n3872_), .B(new_n14638_), .ZN(new_n14639_));
  XOR2_X1    g14383(.A1(new_n14639_), .A2(new_n3876_), .Z(new_n14640_));
  INV_X1     g14384(.I(new_n14640_), .ZN(new_n14641_));
  NAND2_X1   g14385(.A1(new_n14636_), .A2(new_n14641_), .ZN(new_n14642_));
  XOR2_X1    g14386(.A1(new_n14635_), .A2(new_n14521_), .Z(new_n14643_));
  NAND2_X1   g14387(.A1(new_n14643_), .A2(new_n14640_), .ZN(new_n14644_));
  NAND2_X1   g14388(.A1(new_n14642_), .A2(new_n14644_), .ZN(new_n14645_));
  XOR2_X1    g14389(.A1(new_n14645_), .A2(new_n14520_), .Z(new_n14646_));
  OAI22_X1   g14390(.A1(new_n6775_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n6490_), .ZN(new_n14647_));
  AOI21_X1   g14391(.A1(\b[41] ), .A2(new_n3456_), .B(new_n14647_), .ZN(new_n14648_));
  OAI21_X1   g14392(.A1(new_n6785_), .A2(new_n3261_), .B(new_n14648_), .ZN(new_n14649_));
  XOR2_X1    g14393(.A1(new_n14649_), .A2(\a[29] ), .Z(new_n14650_));
  NOR2_X1    g14394(.A1(new_n14646_), .A2(new_n14650_), .ZN(new_n14651_));
  XNOR2_X1   g14395(.A1(new_n14645_), .A2(new_n14520_), .ZN(new_n14652_));
  INV_X1     g14396(.I(new_n14650_), .ZN(new_n14653_));
  NOR2_X1    g14397(.A1(new_n14652_), .A2(new_n14653_), .ZN(new_n14654_));
  NOR2_X1    g14398(.A1(new_n14654_), .A2(new_n14651_), .ZN(new_n14655_));
  XOR2_X1    g14399(.A1(new_n14655_), .A2(new_n14516_), .Z(new_n14656_));
  AOI22_X1   g14400(.A1(new_n2716_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n2719_), .ZN(new_n14657_));
  OAI21_X1   g14401(.A1(new_n7074_), .A2(new_n2924_), .B(new_n14657_), .ZN(new_n14658_));
  AOI21_X1   g14402(.A1(new_n9337_), .A2(new_n2722_), .B(new_n14658_), .ZN(new_n14659_));
  XOR2_X1    g14403(.A1(new_n14659_), .A2(new_n2714_), .Z(new_n14660_));
  NOR2_X1    g14404(.A1(new_n14656_), .A2(new_n14660_), .ZN(new_n14661_));
  XNOR2_X1   g14405(.A1(new_n14655_), .A2(new_n14516_), .ZN(new_n14662_));
  INV_X1     g14406(.I(new_n14660_), .ZN(new_n14663_));
  NOR2_X1    g14407(.A1(new_n14662_), .A2(new_n14663_), .ZN(new_n14664_));
  NOR2_X1    g14408(.A1(new_n14664_), .A2(new_n14661_), .ZN(new_n14665_));
  XOR2_X1    g14409(.A1(new_n14665_), .A2(new_n14513_), .Z(new_n14666_));
  OAI22_X1   g14410(.A1(new_n2189_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n2194_), .ZN(new_n14667_));
  AOI21_X1   g14411(.A1(\b[47] ), .A2(new_n2361_), .B(new_n14667_), .ZN(new_n14668_));
  OAI21_X1   g14412(.A1(new_n9050_), .A2(new_n2197_), .B(new_n14668_), .ZN(new_n14669_));
  XOR2_X1    g14413(.A1(new_n14669_), .A2(\a[23] ), .Z(new_n14670_));
  NOR2_X1    g14414(.A1(new_n14666_), .A2(new_n14670_), .ZN(new_n14671_));
  XNOR2_X1   g14415(.A1(new_n14665_), .A2(new_n14513_), .ZN(new_n14672_));
  INV_X1     g14416(.I(new_n14670_), .ZN(new_n14673_));
  NOR2_X1    g14417(.A1(new_n14672_), .A2(new_n14673_), .ZN(new_n14674_));
  NOR2_X1    g14418(.A1(new_n14674_), .A2(new_n14671_), .ZN(new_n14675_));
  XNOR2_X1   g14419(.A1(new_n14675_), .A2(new_n14511_), .ZN(new_n14676_));
  AOI22_X1   g14420(.A1(new_n1738_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n1743_), .ZN(new_n14677_));
  OAI21_X1   g14421(.A1(new_n8500_), .A2(new_n1931_), .B(new_n14677_), .ZN(new_n14678_));
  AOI21_X1   g14422(.A1(new_n9987_), .A2(new_n1746_), .B(new_n14678_), .ZN(new_n14679_));
  XOR2_X1    g14423(.A1(new_n14679_), .A2(new_n1736_), .Z(new_n14680_));
  INV_X1     g14424(.I(new_n14680_), .ZN(new_n14681_));
  NAND2_X1   g14425(.A1(new_n14676_), .A2(new_n14681_), .ZN(new_n14682_));
  XOR2_X1    g14426(.A1(new_n14675_), .A2(new_n14511_), .Z(new_n14683_));
  NAND2_X1   g14427(.A1(new_n14683_), .A2(new_n14680_), .ZN(new_n14684_));
  NAND2_X1   g14428(.A1(new_n14682_), .A2(new_n14684_), .ZN(new_n14685_));
  XNOR2_X1   g14429(.A1(new_n14685_), .A2(new_n14508_), .ZN(new_n14686_));
  OAI22_X1   g14430(.A1(new_n1592_), .A2(new_n9972_), .B1(new_n9942_), .B2(new_n1505_), .ZN(new_n14687_));
  AOI21_X1   g14431(.A1(\b[53] ), .A2(new_n1584_), .B(new_n14687_), .ZN(new_n14688_));
  OAI21_X1   g14432(.A1(new_n13080_), .A2(new_n1732_), .B(new_n14688_), .ZN(new_n14689_));
  XOR2_X1    g14433(.A1(new_n14689_), .A2(\a[17] ), .Z(new_n14690_));
  INV_X1     g14434(.I(new_n14690_), .ZN(new_n14691_));
  NAND2_X1   g14435(.A1(new_n14686_), .A2(new_n14691_), .ZN(new_n14692_));
  XOR2_X1    g14436(.A1(new_n14685_), .A2(new_n14508_), .Z(new_n14693_));
  NAND2_X1   g14437(.A1(new_n14693_), .A2(new_n14690_), .ZN(new_n14694_));
  NAND2_X1   g14438(.A1(new_n14692_), .A2(new_n14694_), .ZN(new_n14695_));
  XOR2_X1    g14439(.A1(new_n14695_), .A2(new_n14507_), .Z(new_n14696_));
  OAI22_X1   g14440(.A1(new_n993_), .A2(new_n11195_), .B1(new_n10625_), .B2(new_n997_), .ZN(new_n14697_));
  AOI21_X1   g14441(.A1(\b[56] ), .A2(new_n1486_), .B(new_n14697_), .ZN(new_n14698_));
  OAI21_X1   g14442(.A1(new_n11206_), .A2(new_n1323_), .B(new_n14698_), .ZN(new_n14699_));
  XOR2_X1    g14443(.A1(new_n14699_), .A2(\a[14] ), .Z(new_n14700_));
  OR2_X2     g14444(.A1(new_n14696_), .A2(new_n14700_), .Z(new_n14701_));
  NAND2_X1   g14445(.A1(new_n14696_), .A2(new_n14700_), .ZN(new_n14702_));
  NAND2_X1   g14446(.A1(new_n14701_), .A2(new_n14702_), .ZN(new_n14703_));
  XNOR2_X1   g14447(.A1(new_n14703_), .A2(new_n14506_), .ZN(new_n14704_));
  OAI22_X1   g14448(.A1(new_n713_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n717_), .ZN(new_n14705_));
  AOI21_X1   g14449(.A1(\b[59] ), .A2(new_n1126_), .B(new_n14705_), .ZN(new_n14706_));
  OAI21_X1   g14450(.A1(new_n13110_), .A2(new_n986_), .B(new_n14706_), .ZN(new_n14707_));
  XOR2_X1    g14451(.A1(new_n14707_), .A2(new_n722_), .Z(new_n14708_));
  NAND2_X1   g14452(.A1(new_n14704_), .A2(new_n14708_), .ZN(new_n14709_));
  NOR2_X1    g14453(.A1(new_n14704_), .A2(new_n14708_), .ZN(new_n14710_));
  INV_X1     g14454(.I(new_n14710_), .ZN(new_n14711_));
  NAND3_X1   g14455(.A1(new_n14711_), .A2(new_n14504_), .A3(new_n14709_), .ZN(new_n14712_));
  INV_X1     g14456(.I(new_n14709_), .ZN(new_n14713_));
  OAI21_X1   g14457(.A1(new_n14713_), .A2(new_n14710_), .B(new_n14503_), .ZN(new_n14714_));
  OAI22_X1   g14458(.A1(new_n917_), .A2(new_n12796_), .B1(new_n612_), .B2(new_n12800_), .ZN(new_n14715_));
  AOI21_X1   g14459(.A1(new_n13973_), .A2(new_n618_), .B(new_n14715_), .ZN(new_n14716_));
  XOR2_X1    g14460(.A1(new_n14716_), .A2(new_n488_), .Z(new_n14717_));
  INV_X1     g14461(.I(new_n14717_), .ZN(new_n14718_));
  NAND3_X1   g14462(.A1(new_n14714_), .A2(new_n14712_), .A3(new_n14718_), .ZN(new_n14719_));
  NOR3_X1    g14463(.A1(new_n14713_), .A2(new_n14503_), .A3(new_n14710_), .ZN(new_n14720_));
  AOI21_X1   g14464(.A1(new_n14711_), .A2(new_n14709_), .B(new_n14504_), .ZN(new_n14721_));
  OAI21_X1   g14465(.A1(new_n14721_), .A2(new_n14720_), .B(new_n14717_), .ZN(new_n14722_));
  AOI21_X1   g14466(.A1(new_n14722_), .A2(new_n14719_), .B(new_n14501_), .ZN(new_n14723_));
  INV_X1     g14467(.I(new_n14501_), .ZN(new_n14724_));
  NOR3_X1    g14468(.A1(new_n14721_), .A2(new_n14720_), .A3(new_n14717_), .ZN(new_n14725_));
  AOI21_X1   g14469(.A1(new_n14714_), .A2(new_n14712_), .B(new_n14718_), .ZN(new_n14726_));
  NOR3_X1    g14470(.A1(new_n14726_), .A2(new_n14725_), .A3(new_n14724_), .ZN(new_n14727_));
  NOR2_X1    g14471(.A1(new_n14727_), .A2(new_n14723_), .ZN(new_n14728_));
  NAND2_X1   g14472(.A1(new_n14274_), .A2(new_n14494_), .ZN(new_n14729_));
  NAND2_X1   g14473(.A1(new_n14729_), .A2(new_n14491_), .ZN(new_n14730_));
  NAND2_X1   g14474(.A1(new_n14496_), .A2(new_n14271_), .ZN(new_n14731_));
  INV_X1     g14475(.I(new_n14731_), .ZN(new_n14732_));
  AOI21_X1   g14476(.A1(new_n14499_), .A2(new_n14497_), .B(new_n14732_), .ZN(new_n14733_));
  NOR2_X1    g14477(.A1(new_n14733_), .A2(new_n14730_), .ZN(new_n14734_));
  INV_X1     g14478(.I(new_n14730_), .ZN(new_n14735_));
  XNOR2_X1   g14479(.A1(new_n14496_), .A2(new_n14271_), .ZN(new_n14736_));
  NOR3_X1    g14480(.A1(new_n13987_), .A2(new_n13981_), .A3(new_n13988_), .ZN(new_n14737_));
  AOI21_X1   g14481(.A1(new_n13739_), .A2(new_n13989_), .B(new_n14737_), .ZN(new_n14738_));
  NOR2_X1    g14482(.A1(new_n14267_), .A2(new_n14264_), .ZN(new_n14739_));
  OAI21_X1   g14483(.A1(new_n14738_), .A2(new_n14739_), .B(new_n14268_), .ZN(new_n14740_));
  OAI21_X1   g14484(.A1(new_n14740_), .A2(new_n14736_), .B(new_n14731_), .ZN(new_n14741_));
  NOR2_X1    g14485(.A1(new_n14741_), .A2(new_n14735_), .ZN(new_n14742_));
  NOR2_X1    g14486(.A1(new_n14742_), .A2(new_n14734_), .ZN(new_n14743_));
  XOR2_X1    g14487(.A1(new_n14743_), .A2(new_n14728_), .Z(\f[70] ));
  AOI21_X1   g14488(.A1(new_n14741_), .A2(new_n14735_), .B(new_n14728_), .ZN(new_n14745_));
  NOR2_X1    g14489(.A1(new_n14745_), .A2(new_n14742_), .ZN(new_n14746_));
  AOI21_X1   g14490(.A1(new_n14724_), .A2(new_n14722_), .B(new_n14725_), .ZN(new_n14747_));
  INV_X1     g14491(.I(new_n14747_), .ZN(new_n14748_));
  AOI22_X1   g14492(.A1(new_n13460_), .A2(new_n618_), .B1(\b[63] ), .B2(new_n826_), .ZN(new_n14749_));
  XOR2_X1    g14493(.A1(new_n14749_), .A2(new_n488_), .Z(new_n14750_));
  INV_X1     g14494(.I(new_n14750_), .ZN(new_n14751_));
  OAI21_X1   g14495(.A1(new_n14503_), .A2(new_n14710_), .B(new_n14709_), .ZN(new_n14752_));
  NAND2_X1   g14496(.A1(new_n14694_), .A2(new_n14507_), .ZN(new_n14753_));
  AND2_X2    g14497(.A1(new_n14753_), .A2(new_n14692_), .Z(new_n14754_));
  NAND2_X1   g14498(.A1(new_n14684_), .A2(new_n14508_), .ZN(new_n14755_));
  AND2_X2    g14499(.A1(new_n14755_), .A2(new_n14682_), .Z(new_n14756_));
  INV_X1     g14500(.I(new_n14756_), .ZN(new_n14757_));
  INV_X1     g14501(.I(new_n14671_), .ZN(new_n14758_));
  OAI21_X1   g14502(.A1(new_n14511_), .A2(new_n14674_), .B(new_n14758_), .ZN(new_n14759_));
  NOR2_X1    g14503(.A1(new_n14664_), .A2(new_n14513_), .ZN(new_n14760_));
  NOR2_X1    g14504(.A1(new_n14760_), .A2(new_n14661_), .ZN(new_n14761_));
  INV_X1     g14505(.I(new_n14761_), .ZN(new_n14762_));
  AOI22_X1   g14506(.A1(new_n2202_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n2205_), .ZN(new_n14763_));
  OAI21_X1   g14507(.A1(new_n8127_), .A2(new_n2370_), .B(new_n14763_), .ZN(new_n14764_));
  AOI21_X1   g14508(.A1(new_n9684_), .A2(new_n2208_), .B(new_n14764_), .ZN(new_n14765_));
  XOR2_X1    g14509(.A1(new_n14765_), .A2(new_n2200_), .Z(new_n14766_));
  INV_X1     g14510(.I(new_n14766_), .ZN(new_n14767_));
  INV_X1     g14511(.I(new_n14651_), .ZN(new_n14768_));
  OAI21_X1   g14512(.A1(new_n14516_), .A2(new_n14654_), .B(new_n14768_), .ZN(new_n14769_));
  AOI22_X1   g14513(.A1(new_n2716_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n2719_), .ZN(new_n14770_));
  OAI21_X1   g14514(.A1(new_n7096_), .A2(new_n2924_), .B(new_n14770_), .ZN(new_n14771_));
  AOI21_X1   g14515(.A1(new_n7649_), .A2(new_n2722_), .B(new_n14771_), .ZN(new_n14772_));
  XOR2_X1    g14516(.A1(new_n14772_), .A2(new_n2714_), .Z(new_n14773_));
  INV_X1     g14517(.I(new_n14773_), .ZN(new_n14774_));
  NAND2_X1   g14518(.A1(new_n14634_), .A2(new_n14521_), .ZN(new_n14775_));
  AND2_X2    g14519(.A1(new_n14775_), .A2(new_n14631_), .Z(new_n14776_));
  AOI22_X1   g14520(.A1(new_n4918_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n4921_), .ZN(new_n14777_));
  OAI21_X1   g14521(.A1(new_n4886_), .A2(new_n6099_), .B(new_n14777_), .ZN(new_n14778_));
  AOI21_X1   g14522(.A1(new_n5351_), .A2(new_n4699_), .B(new_n14778_), .ZN(new_n14779_));
  XOR2_X1    g14523(.A1(new_n14779_), .A2(new_n4446_), .Z(new_n14780_));
  INV_X1     g14524(.I(new_n14780_), .ZN(new_n14781_));
  NAND2_X1   g14525(.A1(new_n14622_), .A2(new_n14632_), .ZN(new_n14782_));
  AND2_X2    g14526(.A1(new_n14782_), .A2(new_n14623_), .Z(new_n14783_));
  INV_X1     g14527(.I(new_n14783_), .ZN(new_n14784_));
  INV_X1     g14528(.I(new_n14614_), .ZN(new_n14785_));
  AOI21_X1   g14529(.A1(new_n14620_), .A2(new_n14617_), .B(new_n14785_), .ZN(new_n14786_));
  INV_X1     g14530(.I(new_n14534_), .ZN(new_n14787_));
  NOR2_X1    g14531(.A1(new_n14787_), .A2(new_n14606_), .ZN(new_n14788_));
  NAND2_X1   g14532(.A1(new_n14787_), .A2(new_n14606_), .ZN(new_n14789_));
  AOI21_X1   g14533(.A1(new_n14615_), .A2(new_n14789_), .B(new_n14788_), .ZN(new_n14790_));
  INV_X1     g14534(.I(new_n14603_), .ZN(new_n14791_));
  OAI21_X1   g14535(.A1(new_n14536_), .A2(new_n14604_), .B(new_n14791_), .ZN(new_n14792_));
  INV_X1     g14536(.I(new_n14591_), .ZN(new_n14793_));
  OAI21_X1   g14537(.A1(new_n14539_), .A2(new_n14594_), .B(new_n14793_), .ZN(new_n14794_));
  AOI22_X1   g14538(.A1(new_n7403_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n7408_), .ZN(new_n14795_));
  OAI21_X1   g14539(.A1(new_n2495_), .A2(new_n9488_), .B(new_n14795_), .ZN(new_n14796_));
  AOI21_X1   g14540(.A1(new_n3407_), .A2(new_n7414_), .B(new_n14796_), .ZN(new_n14797_));
  XOR2_X1    g14541(.A1(new_n14797_), .A2(\a[47] ), .Z(new_n14798_));
  AOI22_X1   g14542(.A1(new_n8241_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n8246_), .ZN(new_n14799_));
  OAI21_X1   g14543(.A1(new_n2027_), .A2(new_n9114_), .B(new_n14799_), .ZN(new_n14800_));
  AOI21_X1   g14544(.A1(new_n2470_), .A2(new_n8252_), .B(new_n14800_), .ZN(new_n14801_));
  XOR2_X1    g14545(.A1(new_n14801_), .A2(\a[50] ), .Z(new_n14802_));
  AOI22_X1   g14546(.A1(new_n9125_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n9123_), .ZN(new_n14803_));
  OAI21_X1   g14547(.A1(new_n1553_), .A2(new_n9470_), .B(new_n14803_), .ZN(new_n14804_));
  AOI21_X1   g14548(.A1(new_n2452_), .A2(new_n9129_), .B(new_n14804_), .ZN(new_n14805_));
  XOR2_X1    g14549(.A1(new_n14805_), .A2(new_n9133_), .Z(new_n14806_));
  AOI22_X1   g14550(.A1(new_n10981_), .A2(\b[14] ), .B1(new_n10979_), .B2(\b[13] ), .ZN(new_n14807_));
  OAI21_X1   g14551(.A1(new_n941_), .A2(new_n11306_), .B(new_n14807_), .ZN(new_n14808_));
  AOI21_X1   g14552(.A1(new_n1449_), .A2(new_n10984_), .B(new_n14808_), .ZN(new_n14809_));
  XOR2_X1    g14553(.A1(new_n14809_), .A2(\a[59] ), .Z(new_n14810_));
  OAI22_X1   g14554(.A1(new_n13224_), .A2(new_n852_), .B1(new_n776_), .B2(new_n11923_), .ZN(new_n14811_));
  AOI21_X1   g14555(.A1(\b[9] ), .A2(new_n13223_), .B(new_n14811_), .ZN(new_n14812_));
  OAI21_X1   g14556(.A1(new_n859_), .A2(new_n11930_), .B(new_n14812_), .ZN(new_n14813_));
  XOR2_X1    g14557(.A1(new_n14813_), .A2(\a[62] ), .Z(new_n14814_));
  INV_X1     g14558(.I(new_n14814_), .ZN(new_n14815_));
  NAND2_X1   g14559(.A1(new_n14810_), .A2(new_n14815_), .ZN(new_n14816_));
  OR2_X2     g14560(.A1(new_n14810_), .A2(new_n14815_), .Z(new_n14817_));
  NAND2_X1   g14561(.A1(new_n14817_), .A2(new_n14816_), .ZN(new_n14818_));
  OAI21_X1   g14562(.A1(new_n14553_), .A2(new_n14558_), .B(new_n14559_), .ZN(new_n14819_));
  AOI22_X1   g14563(.A1(new_n12922_), .A2(\b[8] ), .B1(\b[7] ), .B2(new_n12923_), .ZN(new_n14820_));
  INV_X1     g14564(.I(new_n14820_), .ZN(new_n14821_));
  NOR2_X1    g14565(.A1(new_n14821_), .A2(new_n14556_), .ZN(new_n14822_));
  NOR2_X1    g14566(.A1(new_n14557_), .A2(new_n14820_), .ZN(new_n14823_));
  OR2_X2     g14567(.A1(new_n14822_), .A2(new_n14823_), .Z(new_n14824_));
  XOR2_X1    g14568(.A1(new_n14819_), .A2(new_n14824_), .Z(new_n14825_));
  XOR2_X1    g14569(.A1(new_n14818_), .A2(new_n14825_), .Z(new_n14826_));
  OAI22_X1   g14570(.A1(new_n11298_), .A2(new_n1432_), .B1(new_n1296_), .B2(new_n11297_), .ZN(new_n14827_));
  AOI21_X1   g14571(.A1(\b[15] ), .A2(new_n11296_), .B(new_n14827_), .ZN(new_n14828_));
  OAI21_X1   g14572(.A1(new_n1444_), .A2(new_n10069_), .B(new_n14828_), .ZN(new_n14829_));
  XOR2_X1    g14573(.A1(new_n14829_), .A2(\a[56] ), .Z(new_n14830_));
  INV_X1     g14574(.I(new_n14570_), .ZN(new_n14831_));
  AOI21_X1   g14575(.A1(new_n14831_), .A2(new_n14549_), .B(new_n14568_), .ZN(new_n14832_));
  NOR2_X1    g14576(.A1(new_n14830_), .A2(new_n14832_), .ZN(new_n14833_));
  INV_X1     g14577(.I(new_n14833_), .ZN(new_n14834_));
  NAND2_X1   g14578(.A1(new_n14830_), .A2(new_n14832_), .ZN(new_n14835_));
  NAND2_X1   g14579(.A1(new_n14834_), .A2(new_n14835_), .ZN(new_n14836_));
  XNOR2_X1   g14580(.A1(new_n14836_), .A2(new_n14826_), .ZN(new_n14837_));
  NOR2_X1    g14581(.A1(new_n14572_), .A2(new_n14574_), .ZN(new_n14838_));
  OAI21_X1   g14582(.A1(new_n14547_), .A2(new_n14838_), .B(new_n14575_), .ZN(new_n14839_));
  NAND2_X1   g14583(.A1(new_n14837_), .A2(new_n14839_), .ZN(new_n14840_));
  OR2_X2     g14584(.A1(new_n14837_), .A2(new_n14839_), .Z(new_n14841_));
  NAND2_X1   g14585(.A1(new_n14841_), .A2(new_n14840_), .ZN(new_n14842_));
  XOR2_X1    g14586(.A1(new_n14842_), .A2(new_n14806_), .Z(new_n14843_));
  NAND2_X1   g14587(.A1(new_n14580_), .A2(new_n14588_), .ZN(new_n14844_));
  NAND2_X1   g14588(.A1(new_n14844_), .A2(new_n14587_), .ZN(new_n14845_));
  NAND2_X1   g14589(.A1(new_n14843_), .A2(new_n14845_), .ZN(new_n14846_));
  INV_X1     g14590(.I(new_n14806_), .ZN(new_n14847_));
  XOR2_X1    g14591(.A1(new_n14842_), .A2(new_n14847_), .Z(new_n14848_));
  NAND3_X1   g14592(.A1(new_n14848_), .A2(new_n14587_), .A3(new_n14844_), .ZN(new_n14849_));
  NAND2_X1   g14593(.A1(new_n14849_), .A2(new_n14846_), .ZN(new_n14850_));
  XNOR2_X1   g14594(.A1(new_n14850_), .A2(new_n14802_), .ZN(new_n14851_));
  OR2_X2     g14595(.A1(new_n14851_), .A2(new_n14798_), .Z(new_n14852_));
  NAND2_X1   g14596(.A1(new_n14851_), .A2(new_n14798_), .ZN(new_n14853_));
  NAND2_X1   g14597(.A1(new_n14852_), .A2(new_n14853_), .ZN(new_n14854_));
  XOR2_X1    g14598(.A1(new_n14854_), .A2(new_n14794_), .Z(new_n14855_));
  AOI22_X1   g14599(.A1(new_n6569_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n6574_), .ZN(new_n14856_));
  OAI21_X1   g14600(.A1(new_n3158_), .A2(new_n8565_), .B(new_n14856_), .ZN(new_n14857_));
  AOI21_X1   g14601(.A1(new_n4188_), .A2(new_n6579_), .B(new_n14857_), .ZN(new_n14858_));
  XOR2_X1    g14602(.A1(new_n14858_), .A2(new_n6567_), .Z(new_n14859_));
  OR2_X2     g14603(.A1(new_n14855_), .A2(new_n14859_), .Z(new_n14860_));
  NAND2_X1   g14604(.A1(new_n14855_), .A2(new_n14859_), .ZN(new_n14861_));
  NAND2_X1   g14605(.A1(new_n14860_), .A2(new_n14861_), .ZN(new_n14862_));
  XOR2_X1    g14606(.A1(new_n14862_), .A2(new_n14792_), .Z(new_n14863_));
  AOI22_X1   g14607(.A1(new_n6108_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n6111_), .ZN(new_n14864_));
  OAI21_X1   g14608(.A1(new_n3624_), .A2(new_n7708_), .B(new_n14864_), .ZN(new_n14865_));
  AOI21_X1   g14609(.A1(new_n4030_), .A2(new_n6105_), .B(new_n14865_), .ZN(new_n14866_));
  XOR2_X1    g14610(.A1(new_n14866_), .A2(new_n5849_), .Z(new_n14867_));
  NOR2_X1    g14611(.A1(new_n14863_), .A2(new_n14867_), .ZN(new_n14868_));
  XNOR2_X1   g14612(.A1(new_n14862_), .A2(new_n14792_), .ZN(new_n14869_));
  INV_X1     g14613(.I(new_n14867_), .ZN(new_n14870_));
  NOR2_X1    g14614(.A1(new_n14869_), .A2(new_n14870_), .ZN(new_n14871_));
  NOR2_X1    g14615(.A1(new_n14871_), .A2(new_n14868_), .ZN(new_n14872_));
  XNOR2_X1   g14616(.A1(new_n14872_), .A2(new_n14790_), .ZN(new_n14873_));
  OAI22_X1   g14617(.A1(new_n4666_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n4639_), .ZN(new_n14874_));
  AOI21_X1   g14618(.A1(\b[33] ), .A2(new_n5420_), .B(new_n14874_), .ZN(new_n14875_));
  OAI21_X1   g14619(.A1(new_n4676_), .A2(new_n6124_), .B(new_n14875_), .ZN(new_n14876_));
  XOR2_X1    g14620(.A1(new_n14876_), .A2(\a[38] ), .Z(new_n14877_));
  INV_X1     g14621(.I(new_n14877_), .ZN(new_n14878_));
  NAND2_X1   g14622(.A1(new_n14873_), .A2(new_n14878_), .ZN(new_n14879_));
  XOR2_X1    g14623(.A1(new_n14872_), .A2(new_n14790_), .Z(new_n14880_));
  NAND2_X1   g14624(.A1(new_n14880_), .A2(new_n14877_), .ZN(new_n14881_));
  NAND2_X1   g14625(.A1(new_n14879_), .A2(new_n14881_), .ZN(new_n14882_));
  XOR2_X1    g14626(.A1(new_n14882_), .A2(new_n14786_), .Z(new_n14883_));
  NAND2_X1   g14627(.A1(new_n14883_), .A2(new_n14784_), .ZN(new_n14884_));
  INV_X1     g14628(.I(new_n14786_), .ZN(new_n14885_));
  XOR2_X1    g14629(.A1(new_n14882_), .A2(new_n14885_), .Z(new_n14886_));
  NAND2_X1   g14630(.A1(new_n14886_), .A2(new_n14783_), .ZN(new_n14887_));
  NAND2_X1   g14631(.A1(new_n14884_), .A2(new_n14887_), .ZN(new_n14888_));
  XOR2_X1    g14632(.A1(new_n14888_), .A2(new_n14781_), .Z(new_n14889_));
  OAI22_X1   g14633(.A1(new_n6284_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n6285_), .ZN(new_n14890_));
  AOI21_X1   g14634(.A1(\b[39] ), .A2(new_n4053_), .B(new_n14890_), .ZN(new_n14891_));
  OAI21_X1   g14635(.A1(new_n6299_), .A2(new_n4727_), .B(new_n14891_), .ZN(new_n14892_));
  XOR2_X1    g14636(.A1(new_n14892_), .A2(\a[32] ), .Z(new_n14893_));
  OR2_X2     g14637(.A1(new_n14889_), .A2(new_n14893_), .Z(new_n14894_));
  NAND2_X1   g14638(.A1(new_n14889_), .A2(new_n14893_), .ZN(new_n14895_));
  NAND2_X1   g14639(.A1(new_n14894_), .A2(new_n14895_), .ZN(new_n14896_));
  XOR2_X1    g14640(.A1(new_n14896_), .A2(new_n14776_), .Z(new_n14897_));
  NOR2_X1    g14641(.A1(new_n14643_), .A2(new_n14640_), .ZN(new_n14898_));
  AOI21_X1   g14642(.A1(new_n14520_), .A2(new_n14644_), .B(new_n14898_), .ZN(new_n14899_));
  AOI22_X1   g14643(.A1(new_n3267_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n3270_), .ZN(new_n14900_));
  OAI21_X1   g14644(.A1(new_n6490_), .A2(new_n3475_), .B(new_n14900_), .ZN(new_n14901_));
  AOI21_X1   g14645(.A1(new_n7906_), .A2(new_n3273_), .B(new_n14901_), .ZN(new_n14902_));
  XOR2_X1    g14646(.A1(new_n14902_), .A2(new_n3264_), .Z(new_n14903_));
  NAND2_X1   g14647(.A1(new_n14899_), .A2(new_n14903_), .ZN(new_n14904_));
  INV_X1     g14648(.I(new_n14904_), .ZN(new_n14905_));
  NOR2_X1    g14649(.A1(new_n14899_), .A2(new_n14903_), .ZN(new_n14906_));
  NOR2_X1    g14650(.A1(new_n14905_), .A2(new_n14906_), .ZN(new_n14907_));
  XOR2_X1    g14651(.A1(new_n14897_), .A2(new_n14907_), .Z(new_n14908_));
  NAND2_X1   g14652(.A1(new_n14908_), .A2(new_n14774_), .ZN(new_n14909_));
  INV_X1     g14653(.I(new_n14907_), .ZN(new_n14910_));
  XOR2_X1    g14654(.A1(new_n14897_), .A2(new_n14910_), .Z(new_n14911_));
  NAND2_X1   g14655(.A1(new_n14911_), .A2(new_n14773_), .ZN(new_n14912_));
  NAND2_X1   g14656(.A1(new_n14909_), .A2(new_n14912_), .ZN(new_n14913_));
  XNOR2_X1   g14657(.A1(new_n14913_), .A2(new_n14769_), .ZN(new_n14914_));
  NAND2_X1   g14658(.A1(new_n14914_), .A2(new_n14767_), .ZN(new_n14915_));
  XOR2_X1    g14659(.A1(new_n14913_), .A2(new_n14769_), .Z(new_n14916_));
  NAND2_X1   g14660(.A1(new_n14916_), .A2(new_n14766_), .ZN(new_n14917_));
  NAND2_X1   g14661(.A1(new_n14915_), .A2(new_n14917_), .ZN(new_n14918_));
  XOR2_X1    g14662(.A1(new_n14918_), .A2(new_n14762_), .Z(new_n14919_));
  OAI22_X1   g14663(.A1(new_n1751_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n1754_), .ZN(new_n14920_));
  AOI21_X1   g14664(.A1(\b[51] ), .A2(new_n1939_), .B(new_n14920_), .ZN(new_n14921_));
  OAI21_X1   g14665(.A1(new_n9385_), .A2(new_n1757_), .B(new_n14921_), .ZN(new_n14922_));
  XOR2_X1    g14666(.A1(new_n14922_), .A2(\a[20] ), .Z(new_n14923_));
  OR2_X2     g14667(.A1(new_n14919_), .A2(new_n14923_), .Z(new_n14924_));
  NAND2_X1   g14668(.A1(new_n14919_), .A2(new_n14923_), .ZN(new_n14925_));
  NAND2_X1   g14669(.A1(new_n14924_), .A2(new_n14925_), .ZN(new_n14926_));
  XOR2_X1    g14670(.A1(new_n14926_), .A2(new_n14759_), .Z(new_n14927_));
  OAI22_X1   g14671(.A1(new_n1592_), .A2(new_n10308_), .B1(new_n9972_), .B2(new_n1505_), .ZN(new_n14928_));
  AOI21_X1   g14672(.A1(\b[54] ), .A2(new_n1584_), .B(new_n14928_), .ZN(new_n14929_));
  OAI21_X1   g14673(.A1(new_n10319_), .A2(new_n1732_), .B(new_n14929_), .ZN(new_n14930_));
  XOR2_X1    g14674(.A1(new_n14930_), .A2(\a[17] ), .Z(new_n14931_));
  NOR2_X1    g14675(.A1(new_n14927_), .A2(new_n14931_), .ZN(new_n14932_));
  XNOR2_X1   g14676(.A1(new_n14926_), .A2(new_n14759_), .ZN(new_n14933_));
  INV_X1     g14677(.I(new_n14931_), .ZN(new_n14934_));
  NOR2_X1    g14678(.A1(new_n14933_), .A2(new_n14934_), .ZN(new_n14935_));
  NOR2_X1    g14679(.A1(new_n14935_), .A2(new_n14932_), .ZN(new_n14936_));
  XOR2_X1    g14680(.A1(new_n14936_), .A2(new_n14757_), .Z(new_n14937_));
  OAI22_X1   g14681(.A1(new_n993_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n997_), .ZN(new_n14938_));
  AOI21_X1   g14682(.A1(\b[57] ), .A2(new_n1486_), .B(new_n14938_), .ZN(new_n14939_));
  OAI21_X1   g14683(.A1(new_n12203_), .A2(new_n1323_), .B(new_n14939_), .ZN(new_n14940_));
  XOR2_X1    g14684(.A1(new_n14940_), .A2(\a[14] ), .Z(new_n14941_));
  INV_X1     g14685(.I(new_n14941_), .ZN(new_n14942_));
  NAND2_X1   g14686(.A1(new_n14937_), .A2(new_n14942_), .ZN(new_n14943_));
  XOR2_X1    g14687(.A1(new_n14936_), .A2(new_n14756_), .Z(new_n14944_));
  NAND2_X1   g14688(.A1(new_n14944_), .A2(new_n14941_), .ZN(new_n14945_));
  NAND2_X1   g14689(.A1(new_n14945_), .A2(new_n14943_), .ZN(new_n14946_));
  XOR2_X1    g14690(.A1(new_n14946_), .A2(new_n14754_), .Z(new_n14947_));
  NAND2_X1   g14691(.A1(new_n14702_), .A2(new_n14506_), .ZN(new_n14948_));
  AND2_X2    g14692(.A1(new_n14948_), .A2(new_n14701_), .Z(new_n14949_));
  INV_X1     g14693(.I(new_n13444_), .ZN(new_n14950_));
  OAI22_X1   g14694(.A1(new_n713_), .A2(new_n12796_), .B1(new_n12148_), .B2(new_n717_), .ZN(new_n14951_));
  AOI21_X1   g14695(.A1(\b[60] ), .A2(new_n1126_), .B(new_n14951_), .ZN(new_n14952_));
  OAI21_X1   g14696(.A1(new_n14950_), .A2(new_n986_), .B(new_n14952_), .ZN(new_n14953_));
  XOR2_X1    g14697(.A1(new_n14953_), .A2(\a[11] ), .Z(new_n14954_));
  NOR2_X1    g14698(.A1(new_n14949_), .A2(new_n14954_), .ZN(new_n14955_));
  AND3_X2    g14699(.A1(new_n14948_), .A2(new_n14701_), .A3(new_n14954_), .Z(new_n14956_));
  NOR2_X1    g14700(.A1(new_n14955_), .A2(new_n14956_), .ZN(new_n14957_));
  XOR2_X1    g14701(.A1(new_n14947_), .A2(new_n14957_), .Z(new_n14958_));
  NOR2_X1    g14702(.A1(new_n14958_), .A2(new_n14752_), .ZN(new_n14959_));
  INV_X1     g14703(.I(new_n14752_), .ZN(new_n14960_));
  INV_X1     g14704(.I(new_n14754_), .ZN(new_n14961_));
  XOR2_X1    g14705(.A1(new_n14946_), .A2(new_n14961_), .Z(new_n14962_));
  XOR2_X1    g14706(.A1(new_n14962_), .A2(new_n14957_), .Z(new_n14963_));
  NOR2_X1    g14707(.A1(new_n14963_), .A2(new_n14960_), .ZN(new_n14964_));
  NOR2_X1    g14708(.A1(new_n14964_), .A2(new_n14959_), .ZN(new_n14965_));
  NAND2_X1   g14709(.A1(new_n14965_), .A2(new_n14751_), .ZN(new_n14966_));
  NAND2_X1   g14710(.A1(new_n14963_), .A2(new_n14960_), .ZN(new_n14967_));
  NAND2_X1   g14711(.A1(new_n14958_), .A2(new_n14752_), .ZN(new_n14968_));
  NAND2_X1   g14712(.A1(new_n14967_), .A2(new_n14968_), .ZN(new_n14969_));
  NAND2_X1   g14713(.A1(new_n14969_), .A2(new_n14750_), .ZN(new_n14970_));
  AOI21_X1   g14714(.A1(new_n14966_), .A2(new_n14970_), .B(new_n14748_), .ZN(new_n14971_));
  NOR2_X1    g14715(.A1(new_n14969_), .A2(new_n14750_), .ZN(new_n14972_));
  NOR2_X1    g14716(.A1(new_n14965_), .A2(new_n14751_), .ZN(new_n14973_));
  NOR3_X1    g14717(.A1(new_n14973_), .A2(new_n14972_), .A3(new_n14747_), .ZN(new_n14974_));
  NOR2_X1    g14718(.A1(new_n14971_), .A2(new_n14974_), .ZN(new_n14975_));
  XOR2_X1    g14719(.A1(new_n14746_), .A2(new_n14975_), .Z(\f[71] ));
  INV_X1     g14720(.I(new_n14971_), .ZN(new_n14977_));
  AOI21_X1   g14721(.A1(new_n14751_), .A2(new_n14967_), .B(new_n14964_), .ZN(new_n14978_));
  INV_X1     g14722(.I(new_n14978_), .ZN(new_n14979_));
  NOR2_X1    g14723(.A1(new_n14962_), .A2(new_n14956_), .ZN(new_n14980_));
  NOR2_X1    g14724(.A1(new_n14980_), .A2(new_n14955_), .ZN(new_n14981_));
  INV_X1     g14725(.I(new_n14981_), .ZN(new_n14982_));
  NAND2_X1   g14726(.A1(new_n14945_), .A2(new_n14961_), .ZN(new_n14983_));
  NAND2_X1   g14727(.A1(new_n14983_), .A2(new_n14943_), .ZN(new_n14984_));
  NOR2_X1    g14728(.A1(new_n14935_), .A2(new_n14756_), .ZN(new_n14985_));
  NOR2_X1    g14729(.A1(new_n14985_), .A2(new_n14932_), .ZN(new_n14986_));
  NAND2_X1   g14730(.A1(new_n14925_), .A2(new_n14759_), .ZN(new_n14987_));
  NAND2_X1   g14731(.A1(new_n14987_), .A2(new_n14924_), .ZN(new_n14988_));
  NAND2_X1   g14732(.A1(new_n14917_), .A2(new_n14762_), .ZN(new_n14989_));
  AND2_X2    g14733(.A1(new_n14989_), .A2(new_n14915_), .Z(new_n14990_));
  NAND2_X1   g14734(.A1(new_n14912_), .A2(new_n14769_), .ZN(new_n14991_));
  NAND2_X1   g14735(.A1(new_n14991_), .A2(new_n14909_), .ZN(new_n14992_));
  AOI22_X1   g14736(.A1(new_n2716_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n2719_), .ZN(new_n14993_));
  OAI21_X1   g14737(.A1(new_n7617_), .A2(new_n2924_), .B(new_n14993_), .ZN(new_n14994_));
  AOI21_X1   g14738(.A1(new_n8792_), .A2(new_n2722_), .B(new_n14994_), .ZN(new_n14995_));
  XOR2_X1    g14739(.A1(new_n14995_), .A2(new_n2714_), .Z(new_n14996_));
  INV_X1     g14740(.I(new_n14776_), .ZN(new_n14997_));
  NAND2_X1   g14741(.A1(new_n14895_), .A2(new_n14997_), .ZN(new_n14998_));
  NAND2_X1   g14742(.A1(new_n14998_), .A2(new_n14894_), .ZN(new_n14999_));
  NAND2_X1   g14743(.A1(new_n14887_), .A2(new_n14781_), .ZN(new_n15000_));
  NAND2_X1   g14744(.A1(new_n15000_), .A2(new_n14884_), .ZN(new_n15001_));
  NAND2_X1   g14745(.A1(new_n14881_), .A2(new_n14885_), .ZN(new_n15002_));
  AND2_X2    g14746(.A1(new_n15002_), .A2(new_n14879_), .Z(new_n15003_));
  NOR2_X1    g14747(.A1(new_n14871_), .A2(new_n14790_), .ZN(new_n15004_));
  NOR2_X1    g14748(.A1(new_n15004_), .A2(new_n14868_), .ZN(new_n15005_));
  NAND2_X1   g14749(.A1(new_n14861_), .A2(new_n14792_), .ZN(new_n15006_));
  NAND2_X1   g14750(.A1(new_n15006_), .A2(new_n14860_), .ZN(new_n15007_));
  NAND2_X1   g14751(.A1(new_n14852_), .A2(new_n14794_), .ZN(new_n15008_));
  NAND2_X1   g14752(.A1(new_n15008_), .A2(new_n14853_), .ZN(new_n15009_));
  NAND2_X1   g14753(.A1(new_n14849_), .A2(new_n14802_), .ZN(new_n15010_));
  AND2_X2    g14754(.A1(new_n15010_), .A2(new_n14846_), .Z(new_n15011_));
  AOI22_X1   g14755(.A1(new_n8241_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n8246_), .ZN(new_n15012_));
  OAI21_X1   g14756(.A1(new_n2142_), .A2(new_n9114_), .B(new_n15012_), .ZN(new_n15013_));
  AOI21_X1   g14757(.A1(new_n3033_), .A2(new_n8252_), .B(new_n15013_), .ZN(new_n15014_));
  XOR2_X1    g14758(.A1(new_n15014_), .A2(new_n8248_), .Z(new_n15015_));
  INV_X1     g14759(.I(new_n15015_), .ZN(new_n15016_));
  NAND2_X1   g14760(.A1(new_n14841_), .A2(new_n14847_), .ZN(new_n15017_));
  AND2_X2    g14761(.A1(new_n15017_), .A2(new_n14840_), .Z(new_n15018_));
  INV_X1     g14762(.I(new_n14825_), .ZN(new_n15019_));
  NAND2_X1   g14763(.A1(new_n14817_), .A2(new_n15019_), .ZN(new_n15020_));
  AND2_X2    g14764(.A1(new_n15020_), .A2(new_n14816_), .Z(new_n15021_));
  OAI22_X1   g14765(.A1(new_n12306_), .A2(new_n1268_), .B1(new_n12305_), .B2(new_n1093_), .ZN(new_n15022_));
  AOI21_X1   g14766(.A1(\b[13] ), .A2(new_n12304_), .B(new_n15022_), .ZN(new_n15023_));
  OAI21_X1   g14767(.A1(new_n1275_), .A2(new_n10985_), .B(new_n15023_), .ZN(new_n15024_));
  XOR2_X1    g14768(.A1(new_n15024_), .A2(\a[59] ), .Z(new_n15025_));
  INV_X1     g14769(.I(new_n14822_), .ZN(new_n15026_));
  AOI21_X1   g14770(.A1(new_n14819_), .A2(new_n15026_), .B(new_n14823_), .ZN(new_n15027_));
  AOI22_X1   g14771(.A1(new_n11926_), .A2(\b[12] ), .B1(new_n11924_), .B2(\b[11] ), .ZN(new_n15028_));
  OAI21_X1   g14772(.A1(new_n776_), .A2(new_n12317_), .B(new_n15028_), .ZN(new_n15029_));
  AOI21_X1   g14773(.A1(new_n1194_), .A2(new_n11929_), .B(new_n15029_), .ZN(new_n15030_));
  XOR2_X1    g14774(.A1(new_n15030_), .A2(new_n12312_), .Z(new_n15031_));
  AOI22_X1   g14775(.A1(new_n12922_), .A2(\b[9] ), .B1(\b[8] ), .B2(new_n12923_), .ZN(new_n15032_));
  NAND2_X1   g14776(.A1(new_n15032_), .A2(\a[8] ), .ZN(new_n15033_));
  OR2_X2     g14777(.A1(new_n15032_), .A2(\a[8] ), .Z(new_n15034_));
  NAND2_X1   g14778(.A1(new_n15034_), .A2(new_n15033_), .ZN(new_n15035_));
  XOR2_X1    g14779(.A1(new_n15035_), .A2(new_n14821_), .Z(new_n15036_));
  INV_X1     g14780(.I(new_n15036_), .ZN(new_n15037_));
  AND2_X2    g14781(.A1(new_n15031_), .A2(new_n15037_), .Z(new_n15038_));
  NOR2_X1    g14782(.A1(new_n15031_), .A2(new_n15037_), .ZN(new_n15039_));
  NOR2_X1    g14783(.A1(new_n15038_), .A2(new_n15039_), .ZN(new_n15040_));
  XOR2_X1    g14784(.A1(new_n15040_), .A2(new_n15027_), .Z(new_n15041_));
  NOR2_X1    g14785(.A1(new_n15041_), .A2(new_n15025_), .ZN(new_n15042_));
  INV_X1     g14786(.I(new_n15042_), .ZN(new_n15043_));
  NAND2_X1   g14787(.A1(new_n15041_), .A2(new_n15025_), .ZN(new_n15044_));
  NAND2_X1   g14788(.A1(new_n15043_), .A2(new_n15044_), .ZN(new_n15045_));
  XOR2_X1    g14789(.A1(new_n15045_), .A2(new_n15021_), .Z(new_n15046_));
  AOI22_X1   g14790(.A1(new_n10064_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n10062_), .ZN(new_n15047_));
  OAI21_X1   g14791(.A1(new_n1296_), .A2(new_n10399_), .B(new_n15047_), .ZN(new_n15048_));
  AOI21_X1   g14792(.A1(new_n2038_), .A2(new_n10068_), .B(new_n15048_), .ZN(new_n15049_));
  XOR2_X1    g14793(.A1(new_n15049_), .A2(new_n10057_), .Z(new_n15050_));
  AOI21_X1   g14794(.A1(new_n14826_), .A2(new_n14835_), .B(new_n14833_), .ZN(new_n15051_));
  OR2_X2     g14795(.A1(new_n15051_), .A2(new_n15050_), .Z(new_n15052_));
  NAND2_X1   g14796(.A1(new_n15051_), .A2(new_n15050_), .ZN(new_n15053_));
  NAND2_X1   g14797(.A1(new_n15052_), .A2(new_n15053_), .ZN(new_n15054_));
  XNOR2_X1   g14798(.A1(new_n15054_), .A2(new_n15046_), .ZN(new_n15055_));
  AOI22_X1   g14799(.A1(new_n9125_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n9123_), .ZN(new_n15056_));
  OAI21_X1   g14800(.A1(new_n1859_), .A2(new_n9470_), .B(new_n15056_), .ZN(new_n15057_));
  AOI21_X1   g14801(.A1(new_n2032_), .A2(new_n9129_), .B(new_n15057_), .ZN(new_n15058_));
  XOR2_X1    g14802(.A1(new_n15058_), .A2(new_n9133_), .Z(new_n15059_));
  INV_X1     g14803(.I(new_n15059_), .ZN(new_n15060_));
  NAND2_X1   g14804(.A1(new_n15055_), .A2(new_n15060_), .ZN(new_n15061_));
  OR2_X2     g14805(.A1(new_n15055_), .A2(new_n15060_), .Z(new_n15062_));
  NAND2_X1   g14806(.A1(new_n15062_), .A2(new_n15061_), .ZN(new_n15063_));
  XOR2_X1    g14807(.A1(new_n15063_), .A2(new_n15018_), .Z(new_n15064_));
  NOR2_X1    g14808(.A1(new_n15064_), .A2(new_n15016_), .ZN(new_n15065_));
  AND2_X2    g14809(.A1(new_n15064_), .A2(new_n15016_), .Z(new_n15066_));
  NOR2_X1    g14810(.A1(new_n15066_), .A2(new_n15065_), .ZN(new_n15067_));
  XOR2_X1    g14811(.A1(new_n15067_), .A2(new_n15011_), .Z(new_n15068_));
  OAI22_X1   g14812(.A1(new_n3006_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n3158_), .ZN(new_n15069_));
  AOI21_X1   g14813(.A1(\b[25] ), .A2(new_n7719_), .B(new_n15069_), .ZN(new_n15070_));
  OAI21_X1   g14814(.A1(new_n3165_), .A2(new_n8585_), .B(new_n15070_), .ZN(new_n15071_));
  XOR2_X1    g14815(.A1(new_n15071_), .A2(\a[47] ), .Z(new_n15072_));
  OR2_X2     g14816(.A1(new_n15068_), .A2(new_n15072_), .Z(new_n15073_));
  NAND2_X1   g14817(.A1(new_n15068_), .A2(new_n15072_), .ZN(new_n15074_));
  NAND2_X1   g14818(.A1(new_n15073_), .A2(new_n15074_), .ZN(new_n15075_));
  XOR2_X1    g14819(.A1(new_n15075_), .A2(new_n15009_), .Z(new_n15076_));
  AOI22_X1   g14820(.A1(new_n6569_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n6574_), .ZN(new_n15077_));
  OAI21_X1   g14821(.A1(new_n3185_), .A2(new_n8565_), .B(new_n15077_), .ZN(new_n15078_));
  AOI21_X1   g14822(.A1(new_n4230_), .A2(new_n6579_), .B(new_n15078_), .ZN(new_n15079_));
  XOR2_X1    g14823(.A1(new_n15079_), .A2(new_n6567_), .Z(new_n15080_));
  NOR2_X1    g14824(.A1(new_n15076_), .A2(new_n15080_), .ZN(new_n15081_));
  NAND2_X1   g14825(.A1(new_n15076_), .A2(new_n15080_), .ZN(new_n15082_));
  INV_X1     g14826(.I(new_n15082_), .ZN(new_n15083_));
  NOR2_X1    g14827(.A1(new_n15083_), .A2(new_n15081_), .ZN(new_n15084_));
  XOR2_X1    g14828(.A1(new_n15084_), .A2(new_n15007_), .Z(new_n15085_));
  AOI22_X1   g14829(.A1(new_n6108_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n6111_), .ZN(new_n15086_));
  OAI21_X1   g14830(.A1(new_n4022_), .A2(new_n7708_), .B(new_n15086_), .ZN(new_n15087_));
  AOI21_X1   g14831(.A1(new_n4223_), .A2(new_n6105_), .B(new_n15087_), .ZN(new_n15088_));
  XOR2_X1    g14832(.A1(new_n15088_), .A2(\a[41] ), .Z(new_n15089_));
  NAND2_X1   g14833(.A1(new_n15085_), .A2(new_n15089_), .ZN(new_n15090_));
  INV_X1     g14834(.I(new_n15090_), .ZN(new_n15091_));
  NOR2_X1    g14835(.A1(new_n15085_), .A2(new_n15089_), .ZN(new_n15092_));
  NOR2_X1    g14836(.A1(new_n15091_), .A2(new_n15092_), .ZN(new_n15093_));
  XNOR2_X1   g14837(.A1(new_n15093_), .A2(new_n15005_), .ZN(new_n15094_));
  AOI22_X1   g14838(.A1(new_n5155_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n5160_), .ZN(new_n15095_));
  OAI21_X1   g14839(.A1(new_n4639_), .A2(new_n6877_), .B(new_n15095_), .ZN(new_n15096_));
  AOI21_X1   g14840(.A1(new_n5594_), .A2(new_n5166_), .B(new_n15096_), .ZN(new_n15097_));
  XOR2_X1    g14841(.A1(new_n15097_), .A2(new_n5162_), .Z(new_n15098_));
  INV_X1     g14842(.I(new_n15098_), .ZN(new_n15099_));
  NAND2_X1   g14843(.A1(new_n15094_), .A2(new_n15099_), .ZN(new_n15100_));
  XOR2_X1    g14844(.A1(new_n15093_), .A2(new_n15005_), .Z(new_n15101_));
  NAND2_X1   g14845(.A1(new_n15101_), .A2(new_n15098_), .ZN(new_n15102_));
  NAND2_X1   g14846(.A1(new_n15100_), .A2(new_n15102_), .ZN(new_n15103_));
  XOR2_X1    g14847(.A1(new_n15103_), .A2(new_n15003_), .Z(new_n15104_));
  AOI22_X1   g14848(.A1(new_n4918_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n4921_), .ZN(new_n15105_));
  OAI21_X1   g14849(.A1(new_n5312_), .A2(new_n6099_), .B(new_n15105_), .ZN(new_n15106_));
  AOI21_X1   g14850(.A1(new_n6310_), .A2(new_n4699_), .B(new_n15106_), .ZN(new_n15107_));
  XOR2_X1    g14851(.A1(new_n15107_), .A2(new_n4446_), .Z(new_n15108_));
  INV_X1     g14852(.I(new_n15108_), .ZN(new_n15109_));
  NAND2_X1   g14853(.A1(new_n15104_), .A2(new_n15109_), .ZN(new_n15110_));
  INV_X1     g14854(.I(new_n15003_), .ZN(new_n15111_));
  XOR2_X1    g14855(.A1(new_n15103_), .A2(new_n15111_), .Z(new_n15112_));
  NAND2_X1   g14856(.A1(new_n15112_), .A2(new_n15108_), .ZN(new_n15113_));
  NAND2_X1   g14857(.A1(new_n15113_), .A2(new_n15110_), .ZN(new_n15114_));
  XOR2_X1    g14858(.A1(new_n15114_), .A2(new_n15001_), .Z(new_n15115_));
  AOI22_X1   g14859(.A1(new_n3864_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n3869_), .ZN(new_n15116_));
  OAI21_X1   g14860(.A1(new_n6284_), .A2(new_n5410_), .B(new_n15116_), .ZN(new_n15117_));
  AOI21_X1   g14861(.A1(new_n7106_), .A2(new_n3872_), .B(new_n15117_), .ZN(new_n15118_));
  XOR2_X1    g14862(.A1(new_n15118_), .A2(new_n3876_), .Z(new_n15119_));
  OR2_X2     g14863(.A1(new_n15115_), .A2(new_n15119_), .Z(new_n15120_));
  NAND2_X1   g14864(.A1(new_n15115_), .A2(new_n15119_), .ZN(new_n15121_));
  NAND2_X1   g14865(.A1(new_n15120_), .A2(new_n15121_), .ZN(new_n15122_));
  XNOR2_X1   g14866(.A1(new_n15122_), .A2(new_n14999_), .ZN(new_n15123_));
  AOI22_X1   g14867(.A1(new_n3267_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n3270_), .ZN(new_n15124_));
  OAI21_X1   g14868(.A1(new_n6775_), .A2(new_n3475_), .B(new_n15124_), .ZN(new_n15125_));
  AOI21_X1   g14869(.A1(new_n7926_), .A2(new_n3273_), .B(new_n15125_), .ZN(new_n15126_));
  XOR2_X1    g14870(.A1(new_n15126_), .A2(new_n3264_), .Z(new_n15127_));
  OAI21_X1   g14871(.A1(new_n14897_), .A2(new_n14910_), .B(new_n14904_), .ZN(new_n15128_));
  NAND2_X1   g14872(.A1(new_n15128_), .A2(new_n15127_), .ZN(new_n15129_));
  OR2_X2     g14873(.A1(new_n15128_), .A2(new_n15127_), .Z(new_n15130_));
  NAND2_X1   g14874(.A1(new_n15130_), .A2(new_n15129_), .ZN(new_n15131_));
  XOR2_X1    g14875(.A1(new_n15131_), .A2(new_n15123_), .Z(new_n15132_));
  NOR2_X1    g14876(.A1(new_n15132_), .A2(new_n14996_), .ZN(new_n15133_));
  INV_X1     g14877(.I(new_n14996_), .ZN(new_n15134_));
  XOR2_X1    g14878(.A1(new_n15122_), .A2(new_n14999_), .Z(new_n15135_));
  XOR2_X1    g14879(.A1(new_n15131_), .A2(new_n15135_), .Z(new_n15136_));
  NOR2_X1    g14880(.A1(new_n15136_), .A2(new_n15134_), .ZN(new_n15137_));
  NOR2_X1    g14881(.A1(new_n15133_), .A2(new_n15137_), .ZN(new_n15138_));
  XOR2_X1    g14882(.A1(new_n15138_), .A2(new_n14992_), .Z(new_n15139_));
  AOI22_X1   g14883(.A1(new_n2202_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n2205_), .ZN(new_n15140_));
  OAI21_X1   g14884(.A1(new_n8168_), .A2(new_n2370_), .B(new_n15140_), .ZN(new_n15141_));
  AOI21_X1   g14885(.A1(new_n8783_), .A2(new_n2208_), .B(new_n15141_), .ZN(new_n15142_));
  XOR2_X1    g14886(.A1(new_n15142_), .A2(\a[23] ), .Z(new_n15143_));
  AND2_X2    g14887(.A1(new_n15139_), .A2(new_n15143_), .Z(new_n15144_));
  NOR2_X1    g14888(.A1(new_n15139_), .A2(new_n15143_), .ZN(new_n15145_));
  NOR2_X1    g14889(.A1(new_n15144_), .A2(new_n15145_), .ZN(new_n15146_));
  XOR2_X1    g14890(.A1(new_n15146_), .A2(new_n14990_), .Z(new_n15147_));
  AOI22_X1   g14891(.A1(new_n1738_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n1743_), .ZN(new_n15148_));
  OAI21_X1   g14892(.A1(new_n9032_), .A2(new_n1931_), .B(new_n15148_), .ZN(new_n15149_));
  AOI21_X1   g14893(.A1(new_n10884_), .A2(new_n1746_), .B(new_n15149_), .ZN(new_n15150_));
  XOR2_X1    g14894(.A1(new_n15150_), .A2(new_n1736_), .Z(new_n15151_));
  NOR2_X1    g14895(.A1(new_n15147_), .A2(new_n15151_), .ZN(new_n15152_));
  INV_X1     g14896(.I(new_n14990_), .ZN(new_n15153_));
  XOR2_X1    g14897(.A1(new_n15146_), .A2(new_n15153_), .Z(new_n15154_));
  INV_X1     g14898(.I(new_n15151_), .ZN(new_n15155_));
  NOR2_X1    g14899(.A1(new_n15154_), .A2(new_n15155_), .ZN(new_n15156_));
  NOR2_X1    g14900(.A1(new_n15152_), .A2(new_n15156_), .ZN(new_n15157_));
  XOR2_X1    g14901(.A1(new_n15157_), .A2(new_n14988_), .Z(new_n15158_));
  OAI22_X1   g14902(.A1(new_n1592_), .A2(new_n10625_), .B1(new_n10308_), .B2(new_n1505_), .ZN(new_n15159_));
  AOI21_X1   g14903(.A1(\b[55] ), .A2(new_n1584_), .B(new_n15159_), .ZN(new_n15160_));
  OAI21_X1   g14904(.A1(new_n13693_), .A2(new_n1732_), .B(new_n15160_), .ZN(new_n15161_));
  XOR2_X1    g14905(.A1(new_n15161_), .A2(new_n1344_), .Z(new_n15162_));
  NAND2_X1   g14906(.A1(new_n15158_), .A2(new_n15162_), .ZN(new_n15163_));
  OR2_X2     g14907(.A1(new_n15158_), .A2(new_n15162_), .Z(new_n15164_));
  NAND2_X1   g14908(.A1(new_n15164_), .A2(new_n15163_), .ZN(new_n15165_));
  XOR2_X1    g14909(.A1(new_n15165_), .A2(new_n14986_), .Z(new_n15166_));
  OAI22_X1   g14910(.A1(new_n993_), .A2(new_n12147_), .B1(new_n12151_), .B2(new_n997_), .ZN(new_n15167_));
  AOI21_X1   g14911(.A1(\b[58] ), .A2(new_n1486_), .B(new_n15167_), .ZN(new_n15168_));
  OAI21_X1   g14912(.A1(new_n11840_), .A2(new_n1323_), .B(new_n15168_), .ZN(new_n15169_));
  XOR2_X1    g14913(.A1(new_n15169_), .A2(\a[14] ), .Z(new_n15170_));
  INV_X1     g14914(.I(new_n15170_), .ZN(new_n15171_));
  NAND2_X1   g14915(.A1(new_n15166_), .A2(new_n15171_), .ZN(new_n15172_));
  INV_X1     g14916(.I(new_n14986_), .ZN(new_n15173_));
  XOR2_X1    g14917(.A1(new_n15165_), .A2(new_n15173_), .Z(new_n15174_));
  NAND2_X1   g14918(.A1(new_n15174_), .A2(new_n15170_), .ZN(new_n15175_));
  NAND2_X1   g14919(.A1(new_n15172_), .A2(new_n15175_), .ZN(new_n15176_));
  NAND2_X1   g14920(.A1(new_n15176_), .A2(new_n14984_), .ZN(new_n15177_));
  INV_X1     g14921(.I(new_n14984_), .ZN(new_n15178_));
  NOR2_X1    g14922(.A1(new_n15174_), .A2(new_n15170_), .ZN(new_n15179_));
  NOR2_X1    g14923(.A1(new_n15166_), .A2(new_n15171_), .ZN(new_n15180_));
  NOR2_X1    g14924(.A1(new_n15180_), .A2(new_n15179_), .ZN(new_n15181_));
  NAND2_X1   g14925(.A1(new_n15181_), .A2(new_n15178_), .ZN(new_n15182_));
  INV_X1     g14926(.I(new_n12811_), .ZN(new_n15183_));
  OAI22_X1   g14927(.A1(new_n713_), .A2(new_n12800_), .B1(new_n12796_), .B2(new_n717_), .ZN(new_n15184_));
  AOI21_X1   g14928(.A1(\b[61] ), .A2(new_n1126_), .B(new_n15184_), .ZN(new_n15185_));
  OAI21_X1   g14929(.A1(new_n15183_), .A2(new_n986_), .B(new_n15185_), .ZN(new_n15186_));
  XOR2_X1    g14930(.A1(new_n15186_), .A2(\a[11] ), .Z(new_n15187_));
  AOI21_X1   g14931(.A1(new_n15182_), .A2(new_n15177_), .B(new_n15187_), .ZN(new_n15188_));
  NOR2_X1    g14932(.A1(new_n15181_), .A2(new_n15178_), .ZN(new_n15189_));
  NOR2_X1    g14933(.A1(new_n15176_), .A2(new_n14984_), .ZN(new_n15190_));
  INV_X1     g14934(.I(new_n15187_), .ZN(new_n15191_));
  NOR3_X1    g14935(.A1(new_n15189_), .A2(new_n15190_), .A3(new_n15191_), .ZN(new_n15192_));
  NOR3_X1    g14936(.A1(new_n15188_), .A2(new_n15192_), .A3(new_n14982_), .ZN(new_n15193_));
  OAI21_X1   g14937(.A1(new_n15189_), .A2(new_n15190_), .B(new_n15191_), .ZN(new_n15194_));
  NAND3_X1   g14938(.A1(new_n15182_), .A2(new_n15177_), .A3(new_n15187_), .ZN(new_n15195_));
  AOI21_X1   g14939(.A1(new_n15194_), .A2(new_n15195_), .B(new_n14981_), .ZN(new_n15196_));
  OAI21_X1   g14940(.A1(new_n15193_), .A2(new_n15196_), .B(new_n14979_), .ZN(new_n15197_));
  NAND3_X1   g14941(.A1(new_n15194_), .A2(new_n15195_), .A3(new_n14981_), .ZN(new_n15198_));
  OAI21_X1   g14942(.A1(new_n15188_), .A2(new_n15192_), .B(new_n14982_), .ZN(new_n15199_));
  NAND3_X1   g14943(.A1(new_n15199_), .A2(new_n15198_), .A3(new_n14978_), .ZN(new_n15200_));
  NAND2_X1   g14944(.A1(new_n15197_), .A2(new_n15200_), .ZN(new_n15201_));
  NAND2_X1   g14945(.A1(new_n14733_), .A2(new_n14730_), .ZN(new_n15202_));
  OAI21_X1   g14946(.A1(new_n14726_), .A2(new_n14725_), .B(new_n14724_), .ZN(new_n15203_));
  NAND3_X1   g14947(.A1(new_n14722_), .A2(new_n14719_), .A3(new_n14501_), .ZN(new_n15204_));
  NAND2_X1   g14948(.A1(new_n15203_), .A2(new_n15204_), .ZN(new_n15205_));
  OAI21_X1   g14949(.A1(new_n14733_), .A2(new_n14730_), .B(new_n15205_), .ZN(new_n15206_));
  NAND3_X1   g14950(.A1(new_n14966_), .A2(new_n14970_), .A3(new_n14748_), .ZN(new_n15207_));
  NAND3_X1   g14951(.A1(new_n15206_), .A2(new_n15202_), .A3(new_n15207_), .ZN(new_n15208_));
  AOI21_X1   g14952(.A1(new_n15208_), .A2(new_n14977_), .B(new_n15201_), .ZN(new_n15209_));
  AOI21_X1   g14953(.A1(new_n15199_), .A2(new_n15198_), .B(new_n14978_), .ZN(new_n15210_));
  NOR3_X1    g14954(.A1(new_n14979_), .A2(new_n15193_), .A3(new_n15196_), .ZN(new_n15211_));
  NOR2_X1    g14955(.A1(new_n15211_), .A2(new_n15210_), .ZN(new_n15212_));
  NOR3_X1    g14956(.A1(new_n14745_), .A2(new_n14742_), .A3(new_n14974_), .ZN(new_n15213_));
  NOR3_X1    g14957(.A1(new_n15213_), .A2(new_n14971_), .A3(new_n15212_), .ZN(new_n15214_));
  NOR2_X1    g14958(.A1(new_n15214_), .A2(new_n15209_), .ZN(\f[72] ));
  AOI21_X1   g14959(.A1(new_n14982_), .A2(new_n15195_), .B(new_n15188_), .ZN(new_n15216_));
  INV_X1     g14960(.I(new_n15216_), .ZN(new_n15217_));
  AOI21_X1   g14961(.A1(new_n14984_), .A2(new_n15175_), .B(new_n15179_), .ZN(new_n15218_));
  INV_X1     g14962(.I(new_n15218_), .ZN(new_n15219_));
  NAND2_X1   g14963(.A1(new_n15164_), .A2(new_n15173_), .ZN(new_n15220_));
  NAND2_X1   g14964(.A1(new_n15220_), .A2(new_n15163_), .ZN(new_n15221_));
  INV_X1     g14965(.I(new_n15156_), .ZN(new_n15222_));
  AOI21_X1   g14966(.A1(new_n15222_), .A2(new_n14988_), .B(new_n15152_), .ZN(new_n15223_));
  INV_X1     g14967(.I(new_n15223_), .ZN(new_n15224_));
  OAI22_X1   g14968(.A1(new_n1592_), .A2(new_n11195_), .B1(new_n10625_), .B2(new_n1505_), .ZN(new_n15225_));
  AOI21_X1   g14969(.A1(\b[56] ), .A2(new_n1584_), .B(new_n15225_), .ZN(new_n15226_));
  OAI21_X1   g14970(.A1(new_n11206_), .A2(new_n1732_), .B(new_n15226_), .ZN(new_n15227_));
  XOR2_X1    g14971(.A1(new_n15227_), .A2(\a[17] ), .Z(new_n15228_));
  NOR2_X1    g14972(.A1(new_n15145_), .A2(new_n14990_), .ZN(new_n15229_));
  NOR2_X1    g14973(.A1(new_n15229_), .A2(new_n15144_), .ZN(new_n15230_));
  INV_X1     g14974(.I(new_n15230_), .ZN(new_n15231_));
  AOI22_X1   g14975(.A1(new_n1738_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n1743_), .ZN(new_n15232_));
  OAI21_X1   g14976(.A1(new_n9376_), .A2(new_n1931_), .B(new_n15232_), .ZN(new_n15233_));
  AOI21_X1   g14977(.A1(new_n9979_), .A2(new_n1746_), .B(new_n15233_), .ZN(new_n15234_));
  XOR2_X1    g14978(.A1(new_n15234_), .A2(new_n1736_), .Z(new_n15235_));
  INV_X1     g14979(.I(new_n15235_), .ZN(new_n15236_));
  INV_X1     g14980(.I(new_n15137_), .ZN(new_n15237_));
  AOI21_X1   g14981(.A1(new_n15237_), .A2(new_n14992_), .B(new_n15133_), .ZN(new_n15238_));
  INV_X1     g14982(.I(new_n15130_), .ZN(new_n15239_));
  AOI21_X1   g14983(.A1(new_n15123_), .A2(new_n15129_), .B(new_n15239_), .ZN(new_n15240_));
  AOI22_X1   g14984(.A1(new_n3267_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n3270_), .ZN(new_n15241_));
  OAI21_X1   g14985(.A1(new_n7074_), .A2(new_n3475_), .B(new_n15241_), .ZN(new_n15242_));
  AOI21_X1   g14986(.A1(new_n9337_), .A2(new_n3273_), .B(new_n15242_), .ZN(new_n15243_));
  XOR2_X1    g14987(.A1(new_n15243_), .A2(new_n3264_), .Z(new_n15244_));
  INV_X1     g14988(.I(new_n15244_), .ZN(new_n15245_));
  NOR2_X1    g14989(.A1(new_n15115_), .A2(new_n15119_), .ZN(new_n15246_));
  AOI21_X1   g14990(.A1(new_n14999_), .A2(new_n15121_), .B(new_n15246_), .ZN(new_n15247_));
  NAND2_X1   g14991(.A1(new_n15113_), .A2(new_n15001_), .ZN(new_n15248_));
  AND2_X2    g14992(.A1(new_n15248_), .A2(new_n15110_), .Z(new_n15249_));
  NAND2_X1   g14993(.A1(new_n15102_), .A2(new_n15111_), .ZN(new_n15250_));
  AND2_X2    g14994(.A1(new_n15250_), .A2(new_n15100_), .Z(new_n15251_));
  OAI21_X1   g14995(.A1(new_n15005_), .A2(new_n15092_), .B(new_n15090_), .ZN(new_n15252_));
  AOI21_X1   g14996(.A1(new_n15007_), .A2(new_n15082_), .B(new_n15081_), .ZN(new_n15253_));
  AOI22_X1   g14997(.A1(new_n6108_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n6111_), .ZN(new_n15254_));
  OAI21_X1   g14998(.A1(new_n4023_), .A2(new_n7708_), .B(new_n15254_), .ZN(new_n15255_));
  AOI21_X1   g14999(.A1(new_n5103_), .A2(new_n6105_), .B(new_n15255_), .ZN(new_n15256_));
  XOR2_X1    g15000(.A1(new_n15256_), .A2(new_n5849_), .Z(new_n15257_));
  AOI22_X1   g15001(.A1(new_n7403_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n7408_), .ZN(new_n15258_));
  OAI21_X1   g15002(.A1(new_n3006_), .A2(new_n9488_), .B(new_n15258_), .ZN(new_n15259_));
  AOI21_X1   g15003(.A1(new_n3807_), .A2(new_n7414_), .B(new_n15259_), .ZN(new_n15260_));
  XOR2_X1    g15004(.A1(new_n15260_), .A2(new_n7410_), .Z(new_n15261_));
  AOI22_X1   g15005(.A1(new_n9125_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n9123_), .ZN(new_n15262_));
  OAI21_X1   g15006(.A1(new_n1860_), .A2(new_n9470_), .B(new_n15262_), .ZN(new_n15263_));
  AOI21_X1   g15007(.A1(new_n2659_), .A2(new_n9129_), .B(new_n15263_), .ZN(new_n15264_));
  XOR2_X1    g15008(.A1(new_n15264_), .A2(new_n9133_), .Z(new_n15265_));
  INV_X1     g15009(.I(new_n15265_), .ZN(new_n15266_));
  NOR2_X1    g15010(.A1(new_n15038_), .A2(new_n15027_), .ZN(new_n15267_));
  NOR2_X1    g15011(.A1(new_n15267_), .A2(new_n15039_), .ZN(new_n15268_));
  AOI22_X1   g15012(.A1(new_n10981_), .A2(\b[16] ), .B1(new_n10979_), .B2(\b[15] ), .ZN(new_n15269_));
  OAI21_X1   g15013(.A1(new_n1093_), .A2(new_n11306_), .B(new_n15269_), .ZN(new_n15270_));
  AOI21_X1   g15014(.A1(new_n1701_), .A2(new_n10984_), .B(new_n15270_), .ZN(new_n15271_));
  XOR2_X1    g15015(.A1(new_n15271_), .A2(new_n10989_), .Z(new_n15272_));
  OAI22_X1   g15016(.A1(new_n13224_), .A2(new_n1070_), .B1(new_n941_), .B2(new_n11923_), .ZN(new_n15273_));
  AOI21_X1   g15017(.A1(\b[11] ), .A2(new_n13223_), .B(new_n15273_), .ZN(new_n15274_));
  OAI21_X1   g15018(.A1(new_n1082_), .A2(new_n11930_), .B(new_n15274_), .ZN(new_n15275_));
  XOR2_X1    g15019(.A1(new_n15275_), .A2(new_n12312_), .Z(new_n15276_));
  NAND2_X1   g15020(.A1(new_n15034_), .A2(new_n14820_), .ZN(new_n15277_));
  NAND2_X1   g15021(.A1(new_n15277_), .A2(new_n15033_), .ZN(new_n15278_));
  AOI22_X1   g15022(.A1(new_n12922_), .A2(\b[10] ), .B1(\b[9] ), .B2(new_n12923_), .ZN(new_n15279_));
  XOR2_X1    g15023(.A1(new_n15278_), .A2(new_n15279_), .Z(new_n15280_));
  XOR2_X1    g15024(.A1(new_n15276_), .A2(new_n15280_), .Z(new_n15281_));
  NOR2_X1    g15025(.A1(new_n15272_), .A2(new_n15281_), .ZN(new_n15282_));
  NAND2_X1   g15026(.A1(new_n15272_), .A2(new_n15281_), .ZN(new_n15283_));
  INV_X1     g15027(.I(new_n15283_), .ZN(new_n15284_));
  NOR2_X1    g15028(.A1(new_n15284_), .A2(new_n15282_), .ZN(new_n15285_));
  XOR2_X1    g15029(.A1(new_n15285_), .A2(new_n15268_), .Z(new_n15286_));
  INV_X1     g15030(.I(new_n15286_), .ZN(new_n15287_));
  INV_X1     g15031(.I(new_n15021_), .ZN(new_n15288_));
  AOI21_X1   g15032(.A1(new_n15288_), .A2(new_n15044_), .B(new_n15042_), .ZN(new_n15289_));
  AOI22_X1   g15033(.A1(new_n10064_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n10062_), .ZN(new_n15290_));
  OAI21_X1   g15034(.A1(new_n1432_), .A2(new_n10399_), .B(new_n15290_), .ZN(new_n15291_));
  AOI21_X1   g15035(.A1(new_n1695_), .A2(new_n10068_), .B(new_n15291_), .ZN(new_n15292_));
  XOR2_X1    g15036(.A1(new_n15292_), .A2(new_n10057_), .Z(new_n15293_));
  NOR2_X1    g15037(.A1(new_n15289_), .A2(new_n15293_), .ZN(new_n15294_));
  INV_X1     g15038(.I(new_n15294_), .ZN(new_n15295_));
  NAND2_X1   g15039(.A1(new_n15289_), .A2(new_n15293_), .ZN(new_n15296_));
  NAND2_X1   g15040(.A1(new_n15295_), .A2(new_n15296_), .ZN(new_n15297_));
  XOR2_X1    g15041(.A1(new_n15297_), .A2(new_n15287_), .Z(new_n15298_));
  NAND2_X1   g15042(.A1(new_n15046_), .A2(new_n15053_), .ZN(new_n15299_));
  NAND2_X1   g15043(.A1(new_n15299_), .A2(new_n15052_), .ZN(new_n15300_));
  XOR2_X1    g15044(.A1(new_n15298_), .A2(new_n15300_), .Z(new_n15301_));
  XOR2_X1    g15045(.A1(new_n15301_), .A2(new_n15266_), .Z(new_n15302_));
  INV_X1     g15046(.I(new_n15018_), .ZN(new_n15303_));
  INV_X1     g15047(.I(new_n15061_), .ZN(new_n15304_));
  AOI21_X1   g15048(.A1(new_n15303_), .A2(new_n15062_), .B(new_n15304_), .ZN(new_n15305_));
  OAI22_X1   g15049(.A1(new_n9461_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n9462_), .ZN(new_n15306_));
  AOI21_X1   g15050(.A1(\b[23] ), .A2(new_n8575_), .B(new_n15306_), .ZN(new_n15307_));
  OAI21_X1   g15051(.A1(new_n2655_), .A2(new_n9460_), .B(new_n15307_), .ZN(new_n15308_));
  XOR2_X1    g15052(.A1(new_n15308_), .A2(\a[50] ), .Z(new_n15309_));
  OR2_X2     g15053(.A1(new_n15305_), .A2(new_n15309_), .Z(new_n15310_));
  NAND2_X1   g15054(.A1(new_n15305_), .A2(new_n15309_), .ZN(new_n15311_));
  NAND2_X1   g15055(.A1(new_n15310_), .A2(new_n15311_), .ZN(new_n15312_));
  XOR2_X1    g15056(.A1(new_n15312_), .A2(new_n15302_), .Z(new_n15313_));
  NOR2_X1    g15057(.A1(new_n15011_), .A2(new_n15065_), .ZN(new_n15314_));
  NOR2_X1    g15058(.A1(new_n15314_), .A2(new_n15066_), .ZN(new_n15315_));
  INV_X1     g15059(.I(new_n15315_), .ZN(new_n15316_));
  NAND2_X1   g15060(.A1(new_n15316_), .A2(new_n15313_), .ZN(new_n15317_));
  OR2_X2     g15061(.A1(new_n15316_), .A2(new_n15313_), .Z(new_n15318_));
  NAND2_X1   g15062(.A1(new_n15318_), .A2(new_n15317_), .ZN(new_n15319_));
  XOR2_X1    g15063(.A1(new_n15319_), .A2(new_n15261_), .Z(new_n15320_));
  NAND2_X1   g15064(.A1(new_n15074_), .A2(new_n15009_), .ZN(new_n15321_));
  NAND2_X1   g15065(.A1(new_n15321_), .A2(new_n15073_), .ZN(new_n15322_));
  AOI22_X1   g15066(.A1(new_n6569_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n6574_), .ZN(new_n15323_));
  OAI21_X1   g15067(.A1(new_n3592_), .A2(new_n8565_), .B(new_n15323_), .ZN(new_n15324_));
  AOI21_X1   g15068(.A1(new_n3796_), .A2(new_n6579_), .B(new_n15324_), .ZN(new_n15325_));
  XOR2_X1    g15069(.A1(new_n15325_), .A2(new_n6567_), .Z(new_n15326_));
  INV_X1     g15070(.I(new_n15326_), .ZN(new_n15327_));
  NAND2_X1   g15071(.A1(new_n15327_), .A2(new_n15322_), .ZN(new_n15328_));
  NAND3_X1   g15072(.A1(new_n15326_), .A2(new_n15073_), .A3(new_n15321_), .ZN(new_n15329_));
  NAND2_X1   g15073(.A1(new_n15328_), .A2(new_n15329_), .ZN(new_n15330_));
  XOR2_X1    g15074(.A1(new_n15330_), .A2(new_n15320_), .Z(new_n15331_));
  NAND2_X1   g15075(.A1(new_n15331_), .A2(new_n15257_), .ZN(new_n15332_));
  OR2_X2     g15076(.A1(new_n15331_), .A2(new_n15257_), .Z(new_n15333_));
  NAND2_X1   g15077(.A1(new_n15333_), .A2(new_n15332_), .ZN(new_n15334_));
  XOR2_X1    g15078(.A1(new_n15334_), .A2(new_n15253_), .Z(new_n15335_));
  OAI22_X1   g15079(.A1(new_n5312_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n4886_), .ZN(new_n15336_));
  AOI21_X1   g15080(.A1(\b[35] ), .A2(new_n5420_), .B(new_n15336_), .ZN(new_n15337_));
  OAI21_X1   g15081(.A1(new_n5322_), .A2(new_n6124_), .B(new_n15337_), .ZN(new_n15338_));
  XOR2_X1    g15082(.A1(new_n15338_), .A2(\a[38] ), .Z(new_n15339_));
  INV_X1     g15083(.I(new_n15339_), .ZN(new_n15340_));
  AND2_X2    g15084(.A1(new_n15335_), .A2(new_n15340_), .Z(new_n15341_));
  NOR2_X1    g15085(.A1(new_n15335_), .A2(new_n15340_), .ZN(new_n15342_));
  NOR2_X1    g15086(.A1(new_n15341_), .A2(new_n15342_), .ZN(new_n15343_));
  XOR2_X1    g15087(.A1(new_n15343_), .A2(new_n15252_), .Z(new_n15344_));
  AOI22_X1   g15088(.A1(new_n4918_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n4921_), .ZN(new_n15345_));
  OAI21_X1   g15089(.A1(new_n5341_), .A2(new_n6099_), .B(new_n15345_), .ZN(new_n15346_));
  AOI21_X1   g15090(.A1(new_n5793_), .A2(new_n4699_), .B(new_n15346_), .ZN(new_n15347_));
  XOR2_X1    g15091(.A1(new_n15347_), .A2(new_n4446_), .Z(new_n15348_));
  INV_X1     g15092(.I(new_n15348_), .ZN(new_n15349_));
  NAND2_X1   g15093(.A1(new_n15344_), .A2(new_n15349_), .ZN(new_n15350_));
  OR2_X2     g15094(.A1(new_n15344_), .A2(new_n15349_), .Z(new_n15351_));
  NAND2_X1   g15095(.A1(new_n15351_), .A2(new_n15350_), .ZN(new_n15352_));
  XOR2_X1    g15096(.A1(new_n15352_), .A2(new_n15251_), .Z(new_n15353_));
  OAI22_X1   g15097(.A1(new_n6490_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n6775_), .ZN(new_n15354_));
  AOI21_X1   g15098(.A1(\b[41] ), .A2(new_n4053_), .B(new_n15354_), .ZN(new_n15355_));
  OAI21_X1   g15099(.A1(new_n6785_), .A2(new_n4727_), .B(new_n15355_), .ZN(new_n15356_));
  XOR2_X1    g15100(.A1(new_n15356_), .A2(new_n3876_), .Z(new_n15357_));
  NAND2_X1   g15101(.A1(new_n15353_), .A2(new_n15357_), .ZN(new_n15358_));
  OR2_X2     g15102(.A1(new_n15353_), .A2(new_n15357_), .Z(new_n15359_));
  NAND2_X1   g15103(.A1(new_n15359_), .A2(new_n15358_), .ZN(new_n15360_));
  XOR2_X1    g15104(.A1(new_n15360_), .A2(new_n15249_), .Z(new_n15361_));
  XOR2_X1    g15105(.A1(new_n15361_), .A2(new_n15247_), .Z(new_n15362_));
  XOR2_X1    g15106(.A1(new_n15362_), .A2(new_n15245_), .Z(new_n15363_));
  OAI22_X1   g15107(.A1(new_n2703_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n2708_), .ZN(new_n15364_));
  AOI21_X1   g15108(.A1(\b[47] ), .A2(new_n2906_), .B(new_n15364_), .ZN(new_n15365_));
  OAI21_X1   g15109(.A1(new_n9050_), .A2(new_n2711_), .B(new_n15365_), .ZN(new_n15366_));
  XOR2_X1    g15110(.A1(new_n15366_), .A2(\a[26] ), .Z(new_n15367_));
  OR2_X2     g15111(.A1(new_n15363_), .A2(new_n15367_), .Z(new_n15368_));
  NAND2_X1   g15112(.A1(new_n15363_), .A2(new_n15367_), .ZN(new_n15369_));
  NAND2_X1   g15113(.A1(new_n15368_), .A2(new_n15369_), .ZN(new_n15370_));
  XOR2_X1    g15114(.A1(new_n15370_), .A2(new_n15240_), .Z(new_n15371_));
  XOR2_X1    g15115(.A1(new_n15371_), .A2(new_n15238_), .Z(new_n15372_));
  AOI22_X1   g15116(.A1(new_n2202_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n2205_), .ZN(new_n15373_));
  OAI21_X1   g15117(.A1(new_n8500_), .A2(new_n2370_), .B(new_n15373_), .ZN(new_n15374_));
  AOI21_X1   g15118(.A1(new_n9987_), .A2(new_n2208_), .B(new_n15374_), .ZN(new_n15375_));
  XOR2_X1    g15119(.A1(new_n15375_), .A2(new_n2200_), .Z(new_n15376_));
  XOR2_X1    g15120(.A1(new_n15372_), .A2(new_n15376_), .Z(new_n15377_));
  NAND2_X1   g15121(.A1(new_n15377_), .A2(new_n15236_), .ZN(new_n15378_));
  INV_X1     g15122(.I(new_n15376_), .ZN(new_n15379_));
  XOR2_X1    g15123(.A1(new_n15372_), .A2(new_n15379_), .Z(new_n15380_));
  NAND2_X1   g15124(.A1(new_n15380_), .A2(new_n15235_), .ZN(new_n15381_));
  NAND2_X1   g15125(.A1(new_n15378_), .A2(new_n15381_), .ZN(new_n15382_));
  XOR2_X1    g15126(.A1(new_n15382_), .A2(new_n15231_), .Z(new_n15383_));
  NOR2_X1    g15127(.A1(new_n15383_), .A2(new_n15228_), .ZN(new_n15384_));
  INV_X1     g15128(.I(new_n15228_), .ZN(new_n15385_));
  XOR2_X1    g15129(.A1(new_n15382_), .A2(new_n15230_), .Z(new_n15386_));
  NOR2_X1    g15130(.A1(new_n15386_), .A2(new_n15385_), .ZN(new_n15387_));
  NOR2_X1    g15131(.A1(new_n15387_), .A2(new_n15384_), .ZN(new_n15388_));
  XOR2_X1    g15132(.A1(new_n15388_), .A2(new_n15224_), .Z(new_n15389_));
  OAI22_X1   g15133(.A1(new_n993_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n997_), .ZN(new_n15390_));
  AOI21_X1   g15134(.A1(\b[59] ), .A2(new_n1486_), .B(new_n15390_), .ZN(new_n15391_));
  OAI21_X1   g15135(.A1(new_n13110_), .A2(new_n1323_), .B(new_n15391_), .ZN(new_n15392_));
  XOR2_X1    g15136(.A1(new_n15392_), .A2(\a[14] ), .Z(new_n15393_));
  INV_X1     g15137(.I(new_n15393_), .ZN(new_n15394_));
  NAND2_X1   g15138(.A1(new_n15389_), .A2(new_n15394_), .ZN(new_n15395_));
  XOR2_X1    g15139(.A1(new_n15388_), .A2(new_n15223_), .Z(new_n15396_));
  NAND2_X1   g15140(.A1(new_n15396_), .A2(new_n15393_), .ZN(new_n15397_));
  NAND2_X1   g15141(.A1(new_n15397_), .A2(new_n15395_), .ZN(new_n15398_));
  XNOR2_X1   g15142(.A1(new_n15398_), .A2(new_n15221_), .ZN(new_n15399_));
  AOI22_X1   g15143(.A1(new_n1126_), .A2(\b[62] ), .B1(\b[63] ), .B2(new_n732_), .ZN(new_n15400_));
  OAI21_X1   g15144(.A1(new_n13107_), .A2(new_n986_), .B(new_n15400_), .ZN(new_n15401_));
  XOR2_X1    g15145(.A1(new_n15401_), .A2(\a[11] ), .Z(new_n15402_));
  INV_X1     g15146(.I(new_n15402_), .ZN(new_n15403_));
  NAND2_X1   g15147(.A1(new_n15399_), .A2(new_n15403_), .ZN(new_n15404_));
  XOR2_X1    g15148(.A1(new_n15398_), .A2(new_n15221_), .Z(new_n15405_));
  NAND2_X1   g15149(.A1(new_n15405_), .A2(new_n15402_), .ZN(new_n15406_));
  NAND2_X1   g15150(.A1(new_n15404_), .A2(new_n15406_), .ZN(new_n15407_));
  XOR2_X1    g15151(.A1(new_n15407_), .A2(new_n15219_), .Z(new_n15408_));
  OAI21_X1   g15152(.A1(new_n15209_), .A2(new_n15211_), .B(new_n15408_), .ZN(new_n15409_));
  OAI21_X1   g15153(.A1(new_n15213_), .A2(new_n14971_), .B(new_n15212_), .ZN(new_n15410_));
  XOR2_X1    g15154(.A1(new_n15407_), .A2(new_n15218_), .Z(new_n15411_));
  NAND3_X1   g15155(.A1(new_n15410_), .A2(new_n15200_), .A3(new_n15411_), .ZN(new_n15412_));
  NAND2_X1   g15156(.A1(new_n15412_), .A2(new_n15409_), .ZN(new_n15413_));
  XOR2_X1    g15157(.A1(new_n15413_), .A2(new_n15217_), .Z(\f[73] ));
  AOI21_X1   g15158(.A1(new_n15410_), .A2(new_n15200_), .B(new_n15411_), .ZN(new_n15415_));
  OAI21_X1   g15159(.A1(new_n15216_), .A2(new_n15415_), .B(new_n15412_), .ZN(new_n15416_));
  NAND2_X1   g15160(.A1(new_n15406_), .A2(new_n15219_), .ZN(new_n15417_));
  NAND2_X1   g15161(.A1(new_n15417_), .A2(new_n15404_), .ZN(new_n15418_));
  OAI22_X1   g15162(.A1(new_n13462_), .A2(new_n986_), .B1(new_n12800_), .B2(new_n1127_), .ZN(new_n15419_));
  XOR2_X1    g15163(.A1(new_n15419_), .A2(\a[11] ), .Z(new_n15420_));
  NAND2_X1   g15164(.A1(new_n15397_), .A2(new_n15221_), .ZN(new_n15421_));
  NAND2_X1   g15165(.A1(new_n15421_), .A2(new_n15395_), .ZN(new_n15422_));
  NOR2_X1    g15166(.A1(new_n15387_), .A2(new_n15223_), .ZN(new_n15423_));
  NOR2_X1    g15167(.A1(new_n15423_), .A2(new_n15384_), .ZN(new_n15424_));
  NAND2_X1   g15168(.A1(new_n15381_), .A2(new_n15231_), .ZN(new_n15425_));
  AND2_X2    g15169(.A1(new_n15425_), .A2(new_n15378_), .Z(new_n15426_));
  INV_X1     g15170(.I(new_n15426_), .ZN(new_n15427_));
  AOI22_X1   g15171(.A1(new_n1738_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n1743_), .ZN(new_n15428_));
  OAI21_X1   g15172(.A1(new_n9942_), .A2(new_n1931_), .B(new_n15428_), .ZN(new_n15429_));
  AOI21_X1   g15173(.A1(new_n10318_), .A2(new_n1746_), .B(new_n15429_), .ZN(new_n15430_));
  XOR2_X1    g15174(.A1(new_n15430_), .A2(new_n1736_), .Z(new_n15431_));
  INV_X1     g15175(.I(new_n15431_), .ZN(new_n15432_));
  INV_X1     g15176(.I(new_n15371_), .ZN(new_n15433_));
  NOR2_X1    g15177(.A1(new_n15433_), .A2(new_n15238_), .ZN(new_n15434_));
  NAND2_X1   g15178(.A1(new_n15433_), .A2(new_n15238_), .ZN(new_n15435_));
  AOI21_X1   g15179(.A1(new_n15379_), .A2(new_n15435_), .B(new_n15434_), .ZN(new_n15436_));
  INV_X1     g15180(.I(new_n15369_), .ZN(new_n15437_));
  OAI21_X1   g15181(.A1(new_n15437_), .A2(new_n15240_), .B(new_n15368_), .ZN(new_n15438_));
  INV_X1     g15182(.I(new_n15361_), .ZN(new_n15439_));
  NOR2_X1    g15183(.A1(new_n15439_), .A2(new_n15247_), .ZN(new_n15440_));
  NAND2_X1   g15184(.A1(new_n15439_), .A2(new_n15247_), .ZN(new_n15441_));
  AOI21_X1   g15185(.A1(new_n15245_), .A2(new_n15441_), .B(new_n15440_), .ZN(new_n15442_));
  INV_X1     g15186(.I(new_n15249_), .ZN(new_n15443_));
  INV_X1     g15187(.I(new_n15358_), .ZN(new_n15444_));
  AOI21_X1   g15188(.A1(new_n15443_), .A2(new_n15359_), .B(new_n15444_), .ZN(new_n15445_));
  AOI22_X1   g15189(.A1(new_n3864_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n3869_), .ZN(new_n15446_));
  OAI21_X1   g15190(.A1(new_n6490_), .A2(new_n5410_), .B(new_n15446_), .ZN(new_n15447_));
  AOI21_X1   g15191(.A1(new_n7906_), .A2(new_n3872_), .B(new_n15447_), .ZN(new_n15448_));
  XOR2_X1    g15192(.A1(new_n15448_), .A2(new_n3876_), .Z(new_n15449_));
  INV_X1     g15193(.I(new_n15449_), .ZN(new_n15450_));
  INV_X1     g15194(.I(new_n15351_), .ZN(new_n15451_));
  OAI21_X1   g15195(.A1(new_n15451_), .A2(new_n15251_), .B(new_n15350_), .ZN(new_n15452_));
  INV_X1     g15196(.I(new_n15252_), .ZN(new_n15453_));
  NOR2_X1    g15197(.A1(new_n15342_), .A2(new_n15453_), .ZN(new_n15454_));
  NOR2_X1    g15198(.A1(new_n15454_), .A2(new_n15341_), .ZN(new_n15455_));
  OAI22_X1   g15199(.A1(new_n6285_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n6284_), .ZN(new_n15456_));
  AOI21_X1   g15200(.A1(\b[39] ), .A2(new_n4706_), .B(new_n15456_), .ZN(new_n15457_));
  OAI21_X1   g15201(.A1(new_n6299_), .A2(new_n4458_), .B(new_n15457_), .ZN(new_n15458_));
  XOR2_X1    g15202(.A1(new_n15458_), .A2(\a[35] ), .Z(new_n15459_));
  INV_X1     g15203(.I(new_n15459_), .ZN(new_n15460_));
  INV_X1     g15204(.I(new_n15253_), .ZN(new_n15461_));
  INV_X1     g15205(.I(new_n15333_), .ZN(new_n15462_));
  AOI21_X1   g15206(.A1(new_n15461_), .A2(new_n15332_), .B(new_n15462_), .ZN(new_n15463_));
  AOI22_X1   g15207(.A1(new_n5155_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n5160_), .ZN(new_n15464_));
  OAI21_X1   g15208(.A1(new_n4886_), .A2(new_n6877_), .B(new_n15464_), .ZN(new_n15465_));
  AOI21_X1   g15209(.A1(new_n5351_), .A2(new_n5166_), .B(new_n15465_), .ZN(new_n15466_));
  XOR2_X1    g15210(.A1(new_n15466_), .A2(new_n5162_), .Z(new_n15467_));
  AOI22_X1   g15211(.A1(new_n6569_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n6574_), .ZN(new_n15468_));
  OAI21_X1   g15212(.A1(new_n3624_), .A2(new_n8565_), .B(new_n15468_), .ZN(new_n15469_));
  AOI21_X1   g15213(.A1(new_n4030_), .A2(new_n6579_), .B(new_n15469_), .ZN(new_n15470_));
  XOR2_X1    g15214(.A1(new_n15470_), .A2(new_n6567_), .Z(new_n15471_));
  AOI22_X1   g15215(.A1(new_n8241_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n8246_), .ZN(new_n15472_));
  OAI21_X1   g15216(.A1(new_n2495_), .A2(new_n9114_), .B(new_n15472_), .ZN(new_n15473_));
  AOI21_X1   g15217(.A1(new_n3407_), .A2(new_n8252_), .B(new_n15473_), .ZN(new_n15474_));
  XOR2_X1    g15218(.A1(new_n15474_), .A2(new_n8248_), .Z(new_n15475_));
  INV_X1     g15219(.I(new_n15300_), .ZN(new_n15476_));
  NOR2_X1    g15220(.A1(new_n15298_), .A2(new_n15476_), .ZN(new_n15477_));
  NAND2_X1   g15221(.A1(new_n15298_), .A2(new_n15476_), .ZN(new_n15478_));
  AOI21_X1   g15222(.A1(new_n15266_), .A2(new_n15478_), .B(new_n15477_), .ZN(new_n15479_));
  INV_X1     g15223(.I(new_n15479_), .ZN(new_n15480_));
  AOI22_X1   g15224(.A1(new_n9125_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n9123_), .ZN(new_n15481_));
  OAI21_X1   g15225(.A1(new_n2027_), .A2(new_n9470_), .B(new_n15481_), .ZN(new_n15482_));
  AOI21_X1   g15226(.A1(new_n2470_), .A2(new_n9129_), .B(new_n15482_), .ZN(new_n15483_));
  XOR2_X1    g15227(.A1(new_n15483_), .A2(\a[53] ), .Z(new_n15484_));
  AOI22_X1   g15228(.A1(new_n10064_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n10062_), .ZN(new_n15485_));
  OAI21_X1   g15229(.A1(new_n1553_), .A2(new_n10399_), .B(new_n15485_), .ZN(new_n15486_));
  AOI21_X1   g15230(.A1(new_n2452_), .A2(new_n10068_), .B(new_n15486_), .ZN(new_n15487_));
  XOR2_X1    g15231(.A1(new_n15487_), .A2(new_n10057_), .Z(new_n15488_));
  INV_X1     g15232(.I(new_n15279_), .ZN(new_n15489_));
  NAND2_X1   g15233(.A1(new_n15278_), .A2(new_n15489_), .ZN(new_n15490_));
  OAI21_X1   g15234(.A1(new_n15278_), .A2(new_n15489_), .B(new_n15276_), .ZN(new_n15491_));
  NAND2_X1   g15235(.A1(new_n15491_), .A2(new_n15490_), .ZN(new_n15492_));
  AOI22_X1   g15236(.A1(new_n12922_), .A2(\b[11] ), .B1(\b[10] ), .B2(new_n12923_), .ZN(new_n15493_));
  INV_X1     g15237(.I(new_n15493_), .ZN(new_n15494_));
  NOR2_X1    g15238(.A1(new_n15494_), .A2(new_n15279_), .ZN(new_n15495_));
  NOR2_X1    g15239(.A1(new_n15489_), .A2(new_n15493_), .ZN(new_n15496_));
  NOR2_X1    g15240(.A1(new_n15495_), .A2(new_n15496_), .ZN(new_n15497_));
  XOR2_X1    g15241(.A1(new_n15492_), .A2(new_n15497_), .Z(new_n15498_));
  OAI22_X1   g15242(.A1(new_n12306_), .A2(new_n1432_), .B1(new_n12305_), .B2(new_n1296_), .ZN(new_n15499_));
  AOI21_X1   g15243(.A1(\b[15] ), .A2(new_n12304_), .B(new_n15499_), .ZN(new_n15500_));
  OAI21_X1   g15244(.A1(new_n1444_), .A2(new_n10985_), .B(new_n15500_), .ZN(new_n15501_));
  XOR2_X1    g15245(.A1(new_n15501_), .A2(\a[59] ), .Z(new_n15502_));
  AOI22_X1   g15246(.A1(new_n11926_), .A2(\b[14] ), .B1(new_n11924_), .B2(\b[13] ), .ZN(new_n15503_));
  OAI21_X1   g15247(.A1(new_n941_), .A2(new_n12317_), .B(new_n15503_), .ZN(new_n15504_));
  AOI21_X1   g15248(.A1(new_n1449_), .A2(new_n11929_), .B(new_n15504_), .ZN(new_n15505_));
  XOR2_X1    g15249(.A1(new_n15505_), .A2(new_n12312_), .Z(new_n15506_));
  NOR2_X1    g15250(.A1(new_n15502_), .A2(new_n15506_), .ZN(new_n15507_));
  INV_X1     g15251(.I(new_n15507_), .ZN(new_n15508_));
  NAND2_X1   g15252(.A1(new_n15502_), .A2(new_n15506_), .ZN(new_n15509_));
  NAND2_X1   g15253(.A1(new_n15508_), .A2(new_n15509_), .ZN(new_n15510_));
  XOR2_X1    g15254(.A1(new_n15510_), .A2(new_n15498_), .Z(new_n15511_));
  NOR2_X1    g15255(.A1(new_n15284_), .A2(new_n15268_), .ZN(new_n15512_));
  NOR2_X1    g15256(.A1(new_n15512_), .A2(new_n15282_), .ZN(new_n15513_));
  NOR2_X1    g15257(.A1(new_n15511_), .A2(new_n15513_), .ZN(new_n15514_));
  INV_X1     g15258(.I(new_n15514_), .ZN(new_n15515_));
  NAND2_X1   g15259(.A1(new_n15511_), .A2(new_n15513_), .ZN(new_n15516_));
  NAND2_X1   g15260(.A1(new_n15515_), .A2(new_n15516_), .ZN(new_n15517_));
  XOR2_X1    g15261(.A1(new_n15517_), .A2(new_n15488_), .Z(new_n15518_));
  AOI21_X1   g15262(.A1(new_n15287_), .A2(new_n15296_), .B(new_n15294_), .ZN(new_n15519_));
  INV_X1     g15263(.I(new_n15519_), .ZN(new_n15520_));
  NAND2_X1   g15264(.A1(new_n15518_), .A2(new_n15520_), .ZN(new_n15521_));
  OR2_X2     g15265(.A1(new_n15518_), .A2(new_n15520_), .Z(new_n15522_));
  NAND2_X1   g15266(.A1(new_n15522_), .A2(new_n15521_), .ZN(new_n15523_));
  XNOR2_X1   g15267(.A1(new_n15523_), .A2(new_n15484_), .ZN(new_n15524_));
  NOR2_X1    g15268(.A1(new_n15524_), .A2(new_n15480_), .ZN(new_n15525_));
  INV_X1     g15269(.I(new_n15525_), .ZN(new_n15526_));
  NAND2_X1   g15270(.A1(new_n15524_), .A2(new_n15480_), .ZN(new_n15527_));
  NAND2_X1   g15271(.A1(new_n15526_), .A2(new_n15527_), .ZN(new_n15528_));
  XOR2_X1    g15272(.A1(new_n15528_), .A2(new_n15475_), .Z(new_n15529_));
  AOI22_X1   g15273(.A1(new_n7403_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n7408_), .ZN(new_n15530_));
  OAI21_X1   g15274(.A1(new_n3158_), .A2(new_n9488_), .B(new_n15530_), .ZN(new_n15531_));
  AOI21_X1   g15275(.A1(new_n4188_), .A2(new_n7414_), .B(new_n15531_), .ZN(new_n15532_));
  XOR2_X1    g15276(.A1(new_n15532_), .A2(new_n7410_), .Z(new_n15533_));
  INV_X1     g15277(.I(new_n15302_), .ZN(new_n15534_));
  INV_X1     g15278(.I(new_n15310_), .ZN(new_n15535_));
  AOI21_X1   g15279(.A1(new_n15534_), .A2(new_n15311_), .B(new_n15535_), .ZN(new_n15536_));
  OR2_X2     g15280(.A1(new_n15533_), .A2(new_n15536_), .Z(new_n15537_));
  NAND2_X1   g15281(.A1(new_n15533_), .A2(new_n15536_), .ZN(new_n15538_));
  NAND2_X1   g15282(.A1(new_n15537_), .A2(new_n15538_), .ZN(new_n15539_));
  XOR2_X1    g15283(.A1(new_n15529_), .A2(new_n15539_), .Z(new_n15540_));
  INV_X1     g15284(.I(new_n15261_), .ZN(new_n15541_));
  INV_X1     g15285(.I(new_n15317_), .ZN(new_n15542_));
  AOI21_X1   g15286(.A1(new_n15541_), .A2(new_n15318_), .B(new_n15542_), .ZN(new_n15543_));
  NOR2_X1    g15287(.A1(new_n15540_), .A2(new_n15543_), .ZN(new_n15544_));
  INV_X1     g15288(.I(new_n15544_), .ZN(new_n15545_));
  NAND2_X1   g15289(.A1(new_n15540_), .A2(new_n15543_), .ZN(new_n15546_));
  NAND2_X1   g15290(.A1(new_n15545_), .A2(new_n15546_), .ZN(new_n15547_));
  XOR2_X1    g15291(.A1(new_n15547_), .A2(new_n15471_), .Z(new_n15548_));
  OAI22_X1   g15292(.A1(new_n5852_), .A2(new_n4666_), .B1(new_n4639_), .B2(new_n5857_), .ZN(new_n15549_));
  AOI21_X1   g15293(.A1(\b[33] ), .A2(new_n6115_), .B(new_n15549_), .ZN(new_n15550_));
  OAI21_X1   g15294(.A1(new_n4676_), .A2(new_n5861_), .B(new_n15550_), .ZN(new_n15551_));
  XOR2_X1    g15295(.A1(new_n15551_), .A2(\a[41] ), .Z(new_n15552_));
  INV_X1     g15296(.I(new_n15328_), .ZN(new_n15553_));
  AOI21_X1   g15297(.A1(new_n15320_), .A2(new_n15329_), .B(new_n15553_), .ZN(new_n15554_));
  NOR2_X1    g15298(.A1(new_n15552_), .A2(new_n15554_), .ZN(new_n15555_));
  INV_X1     g15299(.I(new_n15555_), .ZN(new_n15556_));
  NAND2_X1   g15300(.A1(new_n15552_), .A2(new_n15554_), .ZN(new_n15557_));
  NAND2_X1   g15301(.A1(new_n15556_), .A2(new_n15557_), .ZN(new_n15558_));
  XOR2_X1    g15302(.A1(new_n15548_), .A2(new_n15558_), .Z(new_n15559_));
  NOR2_X1    g15303(.A1(new_n15559_), .A2(new_n15467_), .ZN(new_n15560_));
  AND2_X2    g15304(.A1(new_n15559_), .A2(new_n15467_), .Z(new_n15561_));
  OR2_X2     g15305(.A1(new_n15561_), .A2(new_n15560_), .Z(new_n15562_));
  XOR2_X1    g15306(.A1(new_n15562_), .A2(new_n15463_), .Z(new_n15563_));
  NOR2_X1    g15307(.A1(new_n15563_), .A2(new_n15460_), .ZN(new_n15564_));
  AND2_X2    g15308(.A1(new_n15563_), .A2(new_n15460_), .Z(new_n15565_));
  NOR2_X1    g15309(.A1(new_n15565_), .A2(new_n15564_), .ZN(new_n15566_));
  XNOR2_X1   g15310(.A1(new_n15566_), .A2(new_n15455_), .ZN(new_n15567_));
  NAND2_X1   g15311(.A1(new_n15567_), .A2(new_n15452_), .ZN(new_n15568_));
  OR2_X2     g15312(.A1(new_n15567_), .A2(new_n15452_), .Z(new_n15569_));
  NAND2_X1   g15313(.A1(new_n15569_), .A2(new_n15568_), .ZN(new_n15570_));
  XOR2_X1    g15314(.A1(new_n15570_), .A2(new_n15450_), .Z(new_n15571_));
  AOI22_X1   g15315(.A1(new_n3267_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n3270_), .ZN(new_n15572_));
  OAI21_X1   g15316(.A1(new_n7096_), .A2(new_n3475_), .B(new_n15572_), .ZN(new_n15573_));
  AOI21_X1   g15317(.A1(new_n7649_), .A2(new_n3273_), .B(new_n15573_), .ZN(new_n15574_));
  XOR2_X1    g15318(.A1(new_n15574_), .A2(new_n3264_), .Z(new_n15575_));
  NOR2_X1    g15319(.A1(new_n15571_), .A2(new_n15575_), .ZN(new_n15576_));
  XOR2_X1    g15320(.A1(new_n15570_), .A2(new_n15449_), .Z(new_n15577_));
  INV_X1     g15321(.I(new_n15575_), .ZN(new_n15578_));
  NOR2_X1    g15322(.A1(new_n15577_), .A2(new_n15578_), .ZN(new_n15579_));
  NOR2_X1    g15323(.A1(new_n15576_), .A2(new_n15579_), .ZN(new_n15580_));
  XOR2_X1    g15324(.A1(new_n15580_), .A2(new_n15445_), .Z(new_n15581_));
  NAND2_X1   g15325(.A1(new_n15581_), .A2(new_n15442_), .ZN(new_n15582_));
  OR2_X2     g15326(.A1(new_n15581_), .A2(new_n15442_), .Z(new_n15583_));
  NAND2_X1   g15327(.A1(new_n15583_), .A2(new_n15582_), .ZN(new_n15584_));
  AOI22_X1   g15328(.A1(new_n2716_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n2719_), .ZN(new_n15585_));
  OAI21_X1   g15329(.A1(new_n8127_), .A2(new_n2924_), .B(new_n15585_), .ZN(new_n15586_));
  AOI21_X1   g15330(.A1(new_n9684_), .A2(new_n2722_), .B(new_n15586_), .ZN(new_n15587_));
  XOR2_X1    g15331(.A1(new_n15587_), .A2(new_n2714_), .Z(new_n15588_));
  INV_X1     g15332(.I(new_n15588_), .ZN(new_n15589_));
  XOR2_X1    g15333(.A1(new_n15584_), .A2(new_n15589_), .Z(new_n15590_));
  OAI22_X1   g15334(.A1(new_n2189_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n2194_), .ZN(new_n15591_));
  AOI21_X1   g15335(.A1(\b[51] ), .A2(new_n2361_), .B(new_n15591_), .ZN(new_n15592_));
  OAI21_X1   g15336(.A1(new_n9385_), .A2(new_n2197_), .B(new_n15592_), .ZN(new_n15593_));
  XOR2_X1    g15337(.A1(new_n15593_), .A2(\a[23] ), .Z(new_n15594_));
  OR2_X2     g15338(.A1(new_n15590_), .A2(new_n15594_), .Z(new_n15595_));
  NAND2_X1   g15339(.A1(new_n15590_), .A2(new_n15594_), .ZN(new_n15596_));
  NAND2_X1   g15340(.A1(new_n15595_), .A2(new_n15596_), .ZN(new_n15597_));
  XOR2_X1    g15341(.A1(new_n15597_), .A2(new_n15438_), .Z(new_n15598_));
  XOR2_X1    g15342(.A1(new_n15598_), .A2(new_n15436_), .Z(new_n15599_));
  XOR2_X1    g15343(.A1(new_n15599_), .A2(new_n15432_), .Z(new_n15600_));
  OAI22_X1   g15344(.A1(new_n1592_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n1505_), .ZN(new_n15601_));
  AOI21_X1   g15345(.A1(\b[57] ), .A2(new_n1584_), .B(new_n15601_), .ZN(new_n15602_));
  OAI21_X1   g15346(.A1(new_n12203_), .A2(new_n1732_), .B(new_n15602_), .ZN(new_n15603_));
  XOR2_X1    g15347(.A1(new_n15603_), .A2(\a[17] ), .Z(new_n15604_));
  INV_X1     g15348(.I(new_n15604_), .ZN(new_n15605_));
  NAND2_X1   g15349(.A1(new_n15600_), .A2(new_n15605_), .ZN(new_n15606_));
  XOR2_X1    g15350(.A1(new_n15599_), .A2(new_n15431_), .Z(new_n15607_));
  NAND2_X1   g15351(.A1(new_n15607_), .A2(new_n15604_), .ZN(new_n15608_));
  NAND2_X1   g15352(.A1(new_n15606_), .A2(new_n15608_), .ZN(new_n15609_));
  XOR2_X1    g15353(.A1(new_n15609_), .A2(new_n15427_), .Z(new_n15610_));
  NAND2_X1   g15354(.A1(new_n15610_), .A2(new_n15424_), .ZN(new_n15611_));
  XOR2_X1    g15355(.A1(new_n15609_), .A2(new_n15426_), .Z(new_n15612_));
  OAI21_X1   g15356(.A1(new_n15384_), .A2(new_n15423_), .B(new_n15612_), .ZN(new_n15613_));
  NAND2_X1   g15357(.A1(new_n15613_), .A2(new_n15611_), .ZN(new_n15614_));
  OAI22_X1   g15358(.A1(new_n993_), .A2(new_n12796_), .B1(new_n12148_), .B2(new_n997_), .ZN(new_n15615_));
  AOI21_X1   g15359(.A1(\b[60] ), .A2(new_n1486_), .B(new_n15615_), .ZN(new_n15616_));
  OAI21_X1   g15360(.A1(new_n14950_), .A2(new_n1323_), .B(new_n15616_), .ZN(new_n15617_));
  XOR2_X1    g15361(.A1(new_n15617_), .A2(\a[14] ), .Z(new_n15618_));
  XOR2_X1    g15362(.A1(new_n15614_), .A2(new_n15618_), .Z(new_n15619_));
  NAND2_X1   g15363(.A1(new_n15619_), .A2(new_n15422_), .ZN(new_n15620_));
  INV_X1     g15364(.I(new_n15422_), .ZN(new_n15621_));
  INV_X1     g15365(.I(new_n15618_), .ZN(new_n15622_));
  XOR2_X1    g15366(.A1(new_n15614_), .A2(new_n15622_), .Z(new_n15623_));
  NAND2_X1   g15367(.A1(new_n15623_), .A2(new_n15621_), .ZN(new_n15624_));
  NAND2_X1   g15368(.A1(new_n15620_), .A2(new_n15624_), .ZN(new_n15625_));
  XOR2_X1    g15369(.A1(new_n15625_), .A2(new_n15420_), .Z(new_n15626_));
  NAND2_X1   g15370(.A1(new_n15626_), .A2(new_n15418_), .ZN(new_n15627_));
  INV_X1     g15371(.I(new_n15418_), .ZN(new_n15628_));
  INV_X1     g15372(.I(new_n15420_), .ZN(new_n15629_));
  XOR2_X1    g15373(.A1(new_n15625_), .A2(new_n15629_), .Z(new_n15630_));
  NAND2_X1   g15374(.A1(new_n15630_), .A2(new_n15628_), .ZN(new_n15631_));
  NAND2_X1   g15375(.A1(new_n15627_), .A2(new_n15631_), .ZN(new_n15632_));
  XOR2_X1    g15376(.A1(new_n15632_), .A2(new_n15416_), .Z(\f[74] ));
  INV_X1     g15377(.I(new_n15620_), .ZN(new_n15634_));
  AOI21_X1   g15378(.A1(new_n15629_), .A2(new_n15624_), .B(new_n15634_), .ZN(new_n15635_));
  NAND2_X1   g15379(.A1(new_n15611_), .A2(new_n15622_), .ZN(new_n15636_));
  NAND2_X1   g15380(.A1(new_n15636_), .A2(new_n15613_), .ZN(new_n15637_));
  NAND2_X1   g15381(.A1(new_n15608_), .A2(new_n15427_), .ZN(new_n15638_));
  NAND2_X1   g15382(.A1(new_n15638_), .A2(new_n15606_), .ZN(new_n15639_));
  NOR2_X1    g15383(.A1(new_n15598_), .A2(new_n15436_), .ZN(new_n15640_));
  NAND2_X1   g15384(.A1(new_n15598_), .A2(new_n15436_), .ZN(new_n15641_));
  AOI21_X1   g15385(.A1(new_n15432_), .A2(new_n15641_), .B(new_n15640_), .ZN(new_n15642_));
  NAND2_X1   g15386(.A1(new_n15596_), .A2(new_n15438_), .ZN(new_n15643_));
  NAND2_X1   g15387(.A1(new_n15643_), .A2(new_n15595_), .ZN(new_n15644_));
  INV_X1     g15388(.I(new_n15583_), .ZN(new_n15645_));
  AOI21_X1   g15389(.A1(new_n15582_), .A2(new_n15589_), .B(new_n15645_), .ZN(new_n15646_));
  NOR2_X1    g15390(.A1(new_n15579_), .A2(new_n15445_), .ZN(new_n15647_));
  NOR2_X1    g15391(.A1(new_n15647_), .A2(new_n15576_), .ZN(new_n15648_));
  NAND2_X1   g15392(.A1(new_n15569_), .A2(new_n15450_), .ZN(new_n15649_));
  AND2_X2    g15393(.A1(new_n15649_), .A2(new_n15568_), .Z(new_n15650_));
  INV_X1     g15394(.I(new_n15650_), .ZN(new_n15651_));
  NOR2_X1    g15395(.A1(new_n15564_), .A2(new_n15455_), .ZN(new_n15652_));
  NOR2_X1    g15396(.A1(new_n15652_), .A2(new_n15565_), .ZN(new_n15653_));
  INV_X1     g15397(.I(new_n15560_), .ZN(new_n15654_));
  OAI21_X1   g15398(.A1(new_n15463_), .A2(new_n15561_), .B(new_n15654_), .ZN(new_n15655_));
  AOI21_X1   g15399(.A1(new_n15548_), .A2(new_n15557_), .B(new_n15555_), .ZN(new_n15656_));
  INV_X1     g15400(.I(new_n15471_), .ZN(new_n15657_));
  AOI21_X1   g15401(.A1(new_n15657_), .A2(new_n15546_), .B(new_n15544_), .ZN(new_n15658_));
  NAND2_X1   g15402(.A1(new_n15529_), .A2(new_n15538_), .ZN(new_n15659_));
  NAND2_X1   g15403(.A1(new_n15659_), .A2(new_n15537_), .ZN(new_n15660_));
  OAI21_X1   g15404(.A1(new_n15475_), .A2(new_n15525_), .B(new_n15527_), .ZN(new_n15661_));
  NAND2_X1   g15405(.A1(new_n15522_), .A2(new_n15484_), .ZN(new_n15662_));
  AND2_X2    g15406(.A1(new_n15662_), .A2(new_n15521_), .Z(new_n15663_));
  AOI22_X1   g15407(.A1(new_n9125_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n9123_), .ZN(new_n15664_));
  OAI21_X1   g15408(.A1(new_n2142_), .A2(new_n9470_), .B(new_n15664_), .ZN(new_n15665_));
  AOI21_X1   g15409(.A1(new_n3033_), .A2(new_n9129_), .B(new_n15665_), .ZN(new_n15666_));
  XOR2_X1    g15410(.A1(new_n15666_), .A2(new_n9133_), .Z(new_n15667_));
  INV_X1     g15411(.I(new_n15667_), .ZN(new_n15668_));
  INV_X1     g15412(.I(new_n15488_), .ZN(new_n15669_));
  AOI21_X1   g15413(.A1(new_n15669_), .A2(new_n15516_), .B(new_n15514_), .ZN(new_n15670_));
  AOI22_X1   g15414(.A1(new_n10981_), .A2(\b[18] ), .B1(new_n10979_), .B2(\b[17] ), .ZN(new_n15671_));
  OAI21_X1   g15415(.A1(new_n1296_), .A2(new_n11306_), .B(new_n15671_), .ZN(new_n15672_));
  AOI21_X1   g15416(.A1(new_n2038_), .A2(new_n10984_), .B(new_n15672_), .ZN(new_n15673_));
  XOR2_X1    g15417(.A1(new_n15673_), .A2(new_n10989_), .Z(new_n15674_));
  AOI21_X1   g15418(.A1(new_n15498_), .A2(new_n15509_), .B(new_n15507_), .ZN(new_n15675_));
  OR2_X2     g15419(.A1(new_n15675_), .A2(new_n15674_), .Z(new_n15676_));
  NAND2_X1   g15420(.A1(new_n15675_), .A2(new_n15674_), .ZN(new_n15677_));
  NAND2_X1   g15421(.A1(new_n15676_), .A2(new_n15677_), .ZN(new_n15678_));
  INV_X1     g15422(.I(new_n15496_), .ZN(new_n15679_));
  AOI21_X1   g15423(.A1(new_n15492_), .A2(new_n15679_), .B(new_n15495_), .ZN(new_n15680_));
  OAI22_X1   g15424(.A1(new_n13224_), .A2(new_n1268_), .B1(new_n1093_), .B2(new_n11923_), .ZN(new_n15681_));
  AOI21_X1   g15425(.A1(\b[13] ), .A2(new_n13223_), .B(new_n15681_), .ZN(new_n15682_));
  OAI21_X1   g15426(.A1(new_n1275_), .A2(new_n11930_), .B(new_n15682_), .ZN(new_n15683_));
  XOR2_X1    g15427(.A1(new_n15683_), .A2(\a[62] ), .Z(new_n15684_));
  AOI22_X1   g15428(.A1(new_n12922_), .A2(\b[12] ), .B1(\b[11] ), .B2(new_n12923_), .ZN(new_n15685_));
  INV_X1     g15429(.I(new_n15685_), .ZN(new_n15686_));
  NOR2_X1    g15430(.A1(new_n15686_), .A2(new_n722_), .ZN(new_n15687_));
  NOR2_X1    g15431(.A1(new_n15685_), .A2(\a[11] ), .ZN(new_n15688_));
  NOR2_X1    g15432(.A1(new_n15687_), .A2(new_n15688_), .ZN(new_n15689_));
  XOR2_X1    g15433(.A1(new_n15689_), .A2(new_n15279_), .Z(new_n15690_));
  INV_X1     g15434(.I(new_n15690_), .ZN(new_n15691_));
  NAND2_X1   g15435(.A1(new_n15684_), .A2(new_n15691_), .ZN(new_n15692_));
  NOR2_X1    g15436(.A1(new_n15684_), .A2(new_n15691_), .ZN(new_n15693_));
  INV_X1     g15437(.I(new_n15693_), .ZN(new_n15694_));
  NAND2_X1   g15438(.A1(new_n15694_), .A2(new_n15692_), .ZN(new_n15695_));
  XOR2_X1    g15439(.A1(new_n15695_), .A2(new_n15680_), .Z(new_n15696_));
  XNOR2_X1   g15440(.A1(new_n15678_), .A2(new_n15696_), .ZN(new_n15697_));
  AOI22_X1   g15441(.A1(new_n10064_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n10062_), .ZN(new_n15698_));
  OAI21_X1   g15442(.A1(new_n1859_), .A2(new_n10399_), .B(new_n15698_), .ZN(new_n15699_));
  AOI21_X1   g15443(.A1(new_n2032_), .A2(new_n10068_), .B(new_n15699_), .ZN(new_n15700_));
  XOR2_X1    g15444(.A1(new_n15700_), .A2(new_n10057_), .Z(new_n15701_));
  INV_X1     g15445(.I(new_n15701_), .ZN(new_n15702_));
  NAND2_X1   g15446(.A1(new_n15697_), .A2(new_n15702_), .ZN(new_n15703_));
  OR2_X2     g15447(.A1(new_n15697_), .A2(new_n15702_), .Z(new_n15704_));
  NAND2_X1   g15448(.A1(new_n15704_), .A2(new_n15703_), .ZN(new_n15705_));
  XOR2_X1    g15449(.A1(new_n15705_), .A2(new_n15670_), .Z(new_n15706_));
  NOR2_X1    g15450(.A1(new_n15706_), .A2(new_n15668_), .ZN(new_n15707_));
  AND2_X2    g15451(.A1(new_n15706_), .A2(new_n15668_), .Z(new_n15708_));
  NOR2_X1    g15452(.A1(new_n15708_), .A2(new_n15707_), .ZN(new_n15709_));
  XOR2_X1    g15453(.A1(new_n15709_), .A2(new_n15663_), .Z(new_n15710_));
  OAI22_X1   g15454(.A1(new_n9461_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n9462_), .ZN(new_n15711_));
  AOI21_X1   g15455(.A1(\b[25] ), .A2(new_n8575_), .B(new_n15711_), .ZN(new_n15712_));
  OAI21_X1   g15456(.A1(new_n3165_), .A2(new_n9460_), .B(new_n15712_), .ZN(new_n15713_));
  XOR2_X1    g15457(.A1(new_n15713_), .A2(\a[50] ), .Z(new_n15714_));
  OR2_X2     g15458(.A1(new_n15710_), .A2(new_n15714_), .Z(new_n15715_));
  NAND2_X1   g15459(.A1(new_n15710_), .A2(new_n15714_), .ZN(new_n15716_));
  NAND2_X1   g15460(.A1(new_n15715_), .A2(new_n15716_), .ZN(new_n15717_));
  XOR2_X1    g15461(.A1(new_n15717_), .A2(new_n15661_), .Z(new_n15718_));
  AOI22_X1   g15462(.A1(new_n7403_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n7408_), .ZN(new_n15719_));
  OAI21_X1   g15463(.A1(new_n3185_), .A2(new_n9488_), .B(new_n15719_), .ZN(new_n15720_));
  AOI21_X1   g15464(.A1(new_n4230_), .A2(new_n7414_), .B(new_n15720_), .ZN(new_n15721_));
  XOR2_X1    g15465(.A1(new_n15721_), .A2(new_n7410_), .Z(new_n15722_));
  NOR2_X1    g15466(.A1(new_n15718_), .A2(new_n15722_), .ZN(new_n15723_));
  AND2_X2    g15467(.A1(new_n15718_), .A2(new_n15722_), .Z(new_n15724_));
  NOR2_X1    g15468(.A1(new_n15724_), .A2(new_n15723_), .ZN(new_n15725_));
  XOR2_X1    g15469(.A1(new_n15725_), .A2(new_n15660_), .Z(new_n15726_));
  AOI22_X1   g15470(.A1(new_n6569_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n6574_), .ZN(new_n15727_));
  OAI21_X1   g15471(.A1(new_n4022_), .A2(new_n8565_), .B(new_n15727_), .ZN(new_n15728_));
  AOI21_X1   g15472(.A1(new_n4223_), .A2(new_n6579_), .B(new_n15728_), .ZN(new_n15729_));
  XOR2_X1    g15473(.A1(new_n15729_), .A2(\a[44] ), .Z(new_n15730_));
  NAND2_X1   g15474(.A1(new_n15726_), .A2(new_n15730_), .ZN(new_n15731_));
  OR2_X2     g15475(.A1(new_n15726_), .A2(new_n15730_), .Z(new_n15732_));
  NAND2_X1   g15476(.A1(new_n15732_), .A2(new_n15731_), .ZN(new_n15733_));
  XOR2_X1    g15477(.A1(new_n15733_), .A2(new_n15658_), .Z(new_n15734_));
  AOI22_X1   g15478(.A1(new_n6108_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n6111_), .ZN(new_n15735_));
  OAI21_X1   g15479(.A1(new_n4639_), .A2(new_n7708_), .B(new_n15735_), .ZN(new_n15736_));
  AOI21_X1   g15480(.A1(new_n5594_), .A2(new_n6105_), .B(new_n15736_), .ZN(new_n15737_));
  XOR2_X1    g15481(.A1(new_n15737_), .A2(new_n5849_), .Z(new_n15738_));
  INV_X1     g15482(.I(new_n15738_), .ZN(new_n15739_));
  NAND2_X1   g15483(.A1(new_n15734_), .A2(new_n15739_), .ZN(new_n15740_));
  INV_X1     g15484(.I(new_n15658_), .ZN(new_n15741_));
  XOR2_X1    g15485(.A1(new_n15733_), .A2(new_n15741_), .Z(new_n15742_));
  NAND2_X1   g15486(.A1(new_n15742_), .A2(new_n15738_), .ZN(new_n15743_));
  NAND2_X1   g15487(.A1(new_n15740_), .A2(new_n15743_), .ZN(new_n15744_));
  XOR2_X1    g15488(.A1(new_n15744_), .A2(new_n15656_), .Z(new_n15745_));
  AOI22_X1   g15489(.A1(new_n5155_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n5160_), .ZN(new_n15746_));
  OAI21_X1   g15490(.A1(new_n5312_), .A2(new_n6877_), .B(new_n15746_), .ZN(new_n15747_));
  AOI21_X1   g15491(.A1(new_n6310_), .A2(new_n5166_), .B(new_n15747_), .ZN(new_n15748_));
  XOR2_X1    g15492(.A1(new_n15748_), .A2(new_n5162_), .Z(new_n15749_));
  INV_X1     g15493(.I(new_n15749_), .ZN(new_n15750_));
  NAND2_X1   g15494(.A1(new_n15745_), .A2(new_n15750_), .ZN(new_n15751_));
  INV_X1     g15495(.I(new_n15656_), .ZN(new_n15752_));
  XOR2_X1    g15496(.A1(new_n15744_), .A2(new_n15752_), .Z(new_n15753_));
  NAND2_X1   g15497(.A1(new_n15753_), .A2(new_n15749_), .ZN(new_n15754_));
  NAND2_X1   g15498(.A1(new_n15751_), .A2(new_n15754_), .ZN(new_n15755_));
  XNOR2_X1   g15499(.A1(new_n15755_), .A2(new_n15655_), .ZN(new_n15756_));
  AOI22_X1   g15500(.A1(new_n4918_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n4921_), .ZN(new_n15757_));
  OAI21_X1   g15501(.A1(new_n6284_), .A2(new_n6099_), .B(new_n15757_), .ZN(new_n15758_));
  AOI21_X1   g15502(.A1(new_n7106_), .A2(new_n4699_), .B(new_n15758_), .ZN(new_n15759_));
  XOR2_X1    g15503(.A1(new_n15759_), .A2(new_n4446_), .Z(new_n15760_));
  INV_X1     g15504(.I(new_n15760_), .ZN(new_n15761_));
  NAND2_X1   g15505(.A1(new_n15756_), .A2(new_n15761_), .ZN(new_n15762_));
  XOR2_X1    g15506(.A1(new_n15755_), .A2(new_n15655_), .Z(new_n15763_));
  NAND2_X1   g15507(.A1(new_n15763_), .A2(new_n15760_), .ZN(new_n15764_));
  NAND2_X1   g15508(.A1(new_n15762_), .A2(new_n15764_), .ZN(new_n15765_));
  XOR2_X1    g15509(.A1(new_n15765_), .A2(new_n15653_), .Z(new_n15766_));
  AOI22_X1   g15510(.A1(new_n3864_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n3869_), .ZN(new_n15767_));
  OAI21_X1   g15511(.A1(new_n6775_), .A2(new_n5410_), .B(new_n15767_), .ZN(new_n15768_));
  AOI21_X1   g15512(.A1(new_n7926_), .A2(new_n3872_), .B(new_n15768_), .ZN(new_n15769_));
  XOR2_X1    g15513(.A1(new_n15769_), .A2(new_n3876_), .Z(new_n15770_));
  INV_X1     g15514(.I(new_n15770_), .ZN(new_n15771_));
  NAND2_X1   g15515(.A1(new_n15766_), .A2(new_n15771_), .ZN(new_n15772_));
  INV_X1     g15516(.I(new_n15653_), .ZN(new_n15773_));
  XOR2_X1    g15517(.A1(new_n15765_), .A2(new_n15773_), .Z(new_n15774_));
  NAND2_X1   g15518(.A1(new_n15774_), .A2(new_n15770_), .ZN(new_n15775_));
  NAND2_X1   g15519(.A1(new_n15772_), .A2(new_n15775_), .ZN(new_n15776_));
  XOR2_X1    g15520(.A1(new_n15776_), .A2(new_n15651_), .Z(new_n15777_));
  AOI22_X1   g15521(.A1(new_n3267_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n3270_), .ZN(new_n15778_));
  OAI21_X1   g15522(.A1(new_n7617_), .A2(new_n3475_), .B(new_n15778_), .ZN(new_n15779_));
  AOI21_X1   g15523(.A1(new_n8792_), .A2(new_n3273_), .B(new_n15779_), .ZN(new_n15780_));
  XOR2_X1    g15524(.A1(new_n15780_), .A2(new_n3264_), .Z(new_n15781_));
  NOR2_X1    g15525(.A1(new_n15777_), .A2(new_n15781_), .ZN(new_n15782_));
  XOR2_X1    g15526(.A1(new_n15776_), .A2(new_n15650_), .Z(new_n15783_));
  INV_X1     g15527(.I(new_n15781_), .ZN(new_n15784_));
  NOR2_X1    g15528(.A1(new_n15783_), .A2(new_n15784_), .ZN(new_n15785_));
  NOR2_X1    g15529(.A1(new_n15782_), .A2(new_n15785_), .ZN(new_n15786_));
  XOR2_X1    g15530(.A1(new_n15786_), .A2(new_n15648_), .Z(new_n15787_));
  AOI22_X1   g15531(.A1(new_n2716_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n2719_), .ZN(new_n15788_));
  OAI21_X1   g15532(.A1(new_n8168_), .A2(new_n2924_), .B(new_n15788_), .ZN(new_n15789_));
  AOI21_X1   g15533(.A1(new_n8783_), .A2(new_n2722_), .B(new_n15789_), .ZN(new_n15790_));
  XOR2_X1    g15534(.A1(new_n15790_), .A2(new_n2714_), .Z(new_n15791_));
  NOR2_X1    g15535(.A1(new_n15787_), .A2(new_n15791_), .ZN(new_n15792_));
  XNOR2_X1   g15536(.A1(new_n15786_), .A2(new_n15648_), .ZN(new_n15793_));
  INV_X1     g15537(.I(new_n15791_), .ZN(new_n15794_));
  NOR2_X1    g15538(.A1(new_n15793_), .A2(new_n15794_), .ZN(new_n15795_));
  NOR2_X1    g15539(.A1(new_n15795_), .A2(new_n15792_), .ZN(new_n15796_));
  XOR2_X1    g15540(.A1(new_n15796_), .A2(new_n15646_), .Z(new_n15797_));
  AOI22_X1   g15541(.A1(new_n2202_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n2205_), .ZN(new_n15798_));
  OAI21_X1   g15542(.A1(new_n9032_), .A2(new_n2370_), .B(new_n15798_), .ZN(new_n15799_));
  AOI21_X1   g15543(.A1(new_n10884_), .A2(new_n2208_), .B(new_n15799_), .ZN(new_n15800_));
  XOR2_X1    g15544(.A1(new_n15800_), .A2(new_n2200_), .Z(new_n15801_));
  NOR2_X1    g15545(.A1(new_n15797_), .A2(new_n15801_), .ZN(new_n15802_));
  AND2_X2    g15546(.A1(new_n15797_), .A2(new_n15801_), .Z(new_n15803_));
  NOR2_X1    g15547(.A1(new_n15803_), .A2(new_n15802_), .ZN(new_n15804_));
  XOR2_X1    g15548(.A1(new_n15804_), .A2(new_n15644_), .Z(new_n15805_));
  AOI22_X1   g15549(.A1(new_n1738_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n1743_), .ZN(new_n15806_));
  OAI21_X1   g15550(.A1(new_n9972_), .A2(new_n1931_), .B(new_n15806_), .ZN(new_n15807_));
  AOI21_X1   g15551(.A1(new_n10631_), .A2(new_n1746_), .B(new_n15807_), .ZN(new_n15808_));
  XOR2_X1    g15552(.A1(new_n15808_), .A2(\a[20] ), .Z(new_n15809_));
  NAND2_X1   g15553(.A1(new_n15805_), .A2(new_n15809_), .ZN(new_n15810_));
  OR2_X2     g15554(.A1(new_n15805_), .A2(new_n15809_), .Z(new_n15811_));
  NAND2_X1   g15555(.A1(new_n15811_), .A2(new_n15810_), .ZN(new_n15812_));
  XOR2_X1    g15556(.A1(new_n15812_), .A2(new_n15642_), .Z(new_n15813_));
  OAI22_X1   g15557(.A1(new_n1592_), .A2(new_n12147_), .B1(new_n12151_), .B2(new_n1505_), .ZN(new_n15814_));
  AOI21_X1   g15558(.A1(\b[58] ), .A2(new_n1584_), .B(new_n15814_), .ZN(new_n15815_));
  OAI21_X1   g15559(.A1(new_n11840_), .A2(new_n1732_), .B(new_n15815_), .ZN(new_n15816_));
  XOR2_X1    g15560(.A1(new_n15816_), .A2(\a[17] ), .Z(new_n15817_));
  INV_X1     g15561(.I(new_n15817_), .ZN(new_n15818_));
  NAND2_X1   g15562(.A1(new_n15813_), .A2(new_n15818_), .ZN(new_n15819_));
  INV_X1     g15563(.I(new_n15642_), .ZN(new_n15820_));
  XOR2_X1    g15564(.A1(new_n15812_), .A2(new_n15820_), .Z(new_n15821_));
  NAND2_X1   g15565(.A1(new_n15821_), .A2(new_n15817_), .ZN(new_n15822_));
  NAND2_X1   g15566(.A1(new_n15822_), .A2(new_n15819_), .ZN(new_n15823_));
  XNOR2_X1   g15567(.A1(new_n15823_), .A2(new_n15639_), .ZN(new_n15824_));
  OAI22_X1   g15568(.A1(new_n993_), .A2(new_n12800_), .B1(new_n12796_), .B2(new_n997_), .ZN(new_n15825_));
  AOI21_X1   g15569(.A1(\b[61] ), .A2(new_n1486_), .B(new_n15825_), .ZN(new_n15826_));
  OAI21_X1   g15570(.A1(new_n15183_), .A2(new_n1323_), .B(new_n15826_), .ZN(new_n15827_));
  XOR2_X1    g15571(.A1(new_n15827_), .A2(\a[14] ), .Z(new_n15828_));
  INV_X1     g15572(.I(new_n15828_), .ZN(new_n15829_));
  NAND2_X1   g15573(.A1(new_n15824_), .A2(new_n15829_), .ZN(new_n15830_));
  XOR2_X1    g15574(.A1(new_n15823_), .A2(new_n15639_), .Z(new_n15831_));
  NAND2_X1   g15575(.A1(new_n15831_), .A2(new_n15828_), .ZN(new_n15832_));
  NAND2_X1   g15576(.A1(new_n15830_), .A2(new_n15832_), .ZN(new_n15833_));
  XOR2_X1    g15577(.A1(new_n15833_), .A2(new_n15637_), .Z(new_n15834_));
  XNOR2_X1   g15578(.A1(new_n15834_), .A2(new_n15635_), .ZN(new_n15835_));
  NOR3_X1    g15579(.A1(new_n15209_), .A2(new_n15408_), .A3(new_n15211_), .ZN(new_n15836_));
  AOI21_X1   g15580(.A1(new_n15217_), .A2(new_n15409_), .B(new_n15836_), .ZN(new_n15837_));
  NOR2_X1    g15581(.A1(new_n15626_), .A2(new_n15418_), .ZN(new_n15838_));
  AOI21_X1   g15582(.A1(new_n15837_), .A2(new_n15627_), .B(new_n15838_), .ZN(new_n15839_));
  XOR2_X1    g15583(.A1(new_n15839_), .A2(new_n15835_), .Z(\f[75] ));
  NAND2_X1   g15584(.A1(new_n15832_), .A2(new_n15637_), .ZN(new_n15841_));
  AND2_X2    g15585(.A1(new_n15841_), .A2(new_n15830_), .Z(new_n15842_));
  NAND2_X1   g15586(.A1(new_n15822_), .A2(new_n15639_), .ZN(new_n15843_));
  AND2_X2    g15587(.A1(new_n15843_), .A2(new_n15819_), .Z(new_n15844_));
  NAND2_X1   g15588(.A1(new_n15811_), .A2(new_n15820_), .ZN(new_n15845_));
  AND2_X2    g15589(.A1(new_n15845_), .A2(new_n15810_), .Z(new_n15846_));
  INV_X1     g15590(.I(new_n15846_), .ZN(new_n15847_));
  AOI22_X1   g15591(.A1(new_n1738_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n1743_), .ZN(new_n15848_));
  OAI21_X1   g15592(.A1(new_n10308_), .A2(new_n1931_), .B(new_n15848_), .ZN(new_n15849_));
  AOI21_X1   g15593(.A1(new_n12164_), .A2(new_n1746_), .B(new_n15849_), .ZN(new_n15850_));
  XOR2_X1    g15594(.A1(new_n15850_), .A2(new_n1736_), .Z(new_n15851_));
  INV_X1     g15595(.I(new_n15803_), .ZN(new_n15852_));
  AOI21_X1   g15596(.A1(new_n15852_), .A2(new_n15644_), .B(new_n15802_), .ZN(new_n15853_));
  NOR2_X1    g15597(.A1(new_n15795_), .A2(new_n15646_), .ZN(new_n15854_));
  NOR2_X1    g15598(.A1(new_n15854_), .A2(new_n15792_), .ZN(new_n15855_));
  INV_X1     g15599(.I(new_n15855_), .ZN(new_n15856_));
  NOR2_X1    g15600(.A1(new_n15785_), .A2(new_n15648_), .ZN(new_n15857_));
  NOR2_X1    g15601(.A1(new_n15857_), .A2(new_n15782_), .ZN(new_n15858_));
  INV_X1     g15602(.I(new_n15858_), .ZN(new_n15859_));
  NAND2_X1   g15603(.A1(new_n15775_), .A2(new_n15651_), .ZN(new_n15860_));
  AND2_X2    g15604(.A1(new_n15860_), .A2(new_n15772_), .Z(new_n15861_));
  INV_X1     g15605(.I(new_n15861_), .ZN(new_n15862_));
  INV_X1     g15606(.I(new_n15762_), .ZN(new_n15863_));
  AOI21_X1   g15607(.A1(new_n15773_), .A2(new_n15764_), .B(new_n15863_), .ZN(new_n15864_));
  AOI22_X1   g15608(.A1(new_n3864_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n3869_), .ZN(new_n15865_));
  OAI21_X1   g15609(.A1(new_n7074_), .A2(new_n5410_), .B(new_n15865_), .ZN(new_n15866_));
  AOI21_X1   g15610(.A1(new_n9337_), .A2(new_n3872_), .B(new_n15866_), .ZN(new_n15867_));
  XOR2_X1    g15611(.A1(new_n15864_), .A2(new_n15867_), .Z(new_n15868_));
  INV_X1     g15612(.I(new_n15751_), .ZN(new_n15869_));
  AOI21_X1   g15613(.A1(new_n15655_), .A2(new_n15754_), .B(new_n15869_), .ZN(new_n15870_));
  AOI22_X1   g15614(.A1(new_n5155_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n5160_), .ZN(new_n15871_));
  OAI21_X1   g15615(.A1(new_n5341_), .A2(new_n6877_), .B(new_n15871_), .ZN(new_n15872_));
  AOI21_X1   g15616(.A1(new_n5793_), .A2(new_n5166_), .B(new_n15872_), .ZN(new_n15873_));
  XOR2_X1    g15617(.A1(new_n15873_), .A2(new_n5162_), .Z(new_n15874_));
  INV_X1     g15618(.I(new_n15740_), .ZN(new_n15875_));
  AOI21_X1   g15619(.A1(new_n15752_), .A2(new_n15743_), .B(new_n15875_), .ZN(new_n15876_));
  OAI22_X1   g15620(.A1(new_n5852_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n5857_), .ZN(new_n15877_));
  AOI21_X1   g15621(.A1(\b[35] ), .A2(new_n6115_), .B(new_n15877_), .ZN(new_n15878_));
  OAI21_X1   g15622(.A1(new_n5322_), .A2(new_n5861_), .B(new_n15878_), .ZN(new_n15879_));
  XOR2_X1    g15623(.A1(new_n15879_), .A2(new_n5849_), .Z(new_n15880_));
  NAND2_X1   g15624(.A1(new_n15732_), .A2(new_n15741_), .ZN(new_n15881_));
  AND2_X2    g15625(.A1(new_n15881_), .A2(new_n15731_), .Z(new_n15882_));
  AOI22_X1   g15626(.A1(new_n6569_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n6574_), .ZN(new_n15883_));
  OAI21_X1   g15627(.A1(new_n4023_), .A2(new_n8565_), .B(new_n15883_), .ZN(new_n15884_));
  AOI21_X1   g15628(.A1(new_n5103_), .A2(new_n6579_), .B(new_n15884_), .ZN(new_n15885_));
  XOR2_X1    g15629(.A1(new_n15885_), .A2(new_n6567_), .Z(new_n15886_));
  INV_X1     g15630(.I(new_n15724_), .ZN(new_n15887_));
  AOI21_X1   g15631(.A1(new_n15887_), .A2(new_n15660_), .B(new_n15723_), .ZN(new_n15888_));
  INV_X1     g15632(.I(new_n15888_), .ZN(new_n15889_));
  AOI22_X1   g15633(.A1(new_n7403_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n7408_), .ZN(new_n15890_));
  OAI21_X1   g15634(.A1(new_n3592_), .A2(new_n9488_), .B(new_n15890_), .ZN(new_n15891_));
  AOI21_X1   g15635(.A1(new_n3796_), .A2(new_n7414_), .B(new_n15891_), .ZN(new_n15892_));
  XOR2_X1    g15636(.A1(new_n15892_), .A2(\a[47] ), .Z(new_n15893_));
  INV_X1     g15637(.I(new_n15715_), .ZN(new_n15894_));
  AOI21_X1   g15638(.A1(new_n15661_), .A2(new_n15716_), .B(new_n15894_), .ZN(new_n15895_));
  AOI22_X1   g15639(.A1(new_n8241_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n8246_), .ZN(new_n15896_));
  OAI21_X1   g15640(.A1(new_n3006_), .A2(new_n9114_), .B(new_n15896_), .ZN(new_n15897_));
  AOI21_X1   g15641(.A1(new_n3807_), .A2(new_n8252_), .B(new_n15897_), .ZN(new_n15898_));
  XOR2_X1    g15642(.A1(new_n15898_), .A2(new_n8248_), .Z(new_n15899_));
  AOI22_X1   g15643(.A1(new_n10064_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n10062_), .ZN(new_n15900_));
  OAI21_X1   g15644(.A1(new_n1860_), .A2(new_n10399_), .B(new_n15900_), .ZN(new_n15901_));
  AOI21_X1   g15645(.A1(new_n2659_), .A2(new_n10068_), .B(new_n15901_), .ZN(new_n15902_));
  XOR2_X1    g15646(.A1(new_n15902_), .A2(new_n10057_), .Z(new_n15903_));
  INV_X1     g15647(.I(new_n15903_), .ZN(new_n15904_));
  AOI22_X1   g15648(.A1(new_n11926_), .A2(\b[16] ), .B1(new_n11924_), .B2(\b[15] ), .ZN(new_n15905_));
  OAI21_X1   g15649(.A1(new_n1093_), .A2(new_n12317_), .B(new_n15905_), .ZN(new_n15906_));
  AOI21_X1   g15650(.A1(new_n1701_), .A2(new_n11929_), .B(new_n15906_), .ZN(new_n15907_));
  XOR2_X1    g15651(.A1(new_n15907_), .A2(\a[62] ), .Z(new_n15908_));
  NOR2_X1    g15652(.A1(new_n15688_), .A2(new_n15489_), .ZN(new_n15909_));
  NOR2_X1    g15653(.A1(new_n15909_), .A2(new_n15687_), .ZN(new_n15910_));
  AOI22_X1   g15654(.A1(new_n12922_), .A2(\b[13] ), .B1(\b[12] ), .B2(new_n12923_), .ZN(new_n15911_));
  INV_X1     g15655(.I(new_n15911_), .ZN(new_n15912_));
  XOR2_X1    g15656(.A1(new_n15910_), .A2(new_n15912_), .Z(new_n15913_));
  XOR2_X1    g15657(.A1(new_n15908_), .A2(new_n15913_), .Z(new_n15914_));
  INV_X1     g15658(.I(new_n15914_), .ZN(new_n15915_));
  INV_X1     g15659(.I(new_n15680_), .ZN(new_n15916_));
  AOI21_X1   g15660(.A1(new_n15916_), .A2(new_n15692_), .B(new_n15693_), .ZN(new_n15917_));
  AOI22_X1   g15661(.A1(new_n10981_), .A2(\b[19] ), .B1(new_n10979_), .B2(\b[18] ), .ZN(new_n15918_));
  OAI21_X1   g15662(.A1(new_n1432_), .A2(new_n11306_), .B(new_n15918_), .ZN(new_n15919_));
  AOI21_X1   g15663(.A1(new_n1695_), .A2(new_n10984_), .B(new_n15919_), .ZN(new_n15920_));
  XOR2_X1    g15664(.A1(new_n15920_), .A2(new_n10989_), .Z(new_n15921_));
  NOR2_X1    g15665(.A1(new_n15921_), .A2(new_n15917_), .ZN(new_n15922_));
  INV_X1     g15666(.I(new_n15922_), .ZN(new_n15923_));
  NAND2_X1   g15667(.A1(new_n15921_), .A2(new_n15917_), .ZN(new_n15924_));
  NAND2_X1   g15668(.A1(new_n15923_), .A2(new_n15924_), .ZN(new_n15925_));
  XOR2_X1    g15669(.A1(new_n15925_), .A2(new_n15915_), .Z(new_n15926_));
  NAND2_X1   g15670(.A1(new_n15696_), .A2(new_n15677_), .ZN(new_n15927_));
  NAND2_X1   g15671(.A1(new_n15927_), .A2(new_n15676_), .ZN(new_n15928_));
  INV_X1     g15672(.I(new_n15928_), .ZN(new_n15929_));
  NOR2_X1    g15673(.A1(new_n15926_), .A2(new_n15929_), .ZN(new_n15930_));
  INV_X1     g15674(.I(new_n15930_), .ZN(new_n15931_));
  NAND2_X1   g15675(.A1(new_n15926_), .A2(new_n15929_), .ZN(new_n15932_));
  NAND2_X1   g15676(.A1(new_n15931_), .A2(new_n15932_), .ZN(new_n15933_));
  XOR2_X1    g15677(.A1(new_n15933_), .A2(new_n15904_), .Z(new_n15934_));
  INV_X1     g15678(.I(new_n15934_), .ZN(new_n15935_));
  INV_X1     g15679(.I(new_n15670_), .ZN(new_n15936_));
  INV_X1     g15680(.I(new_n15703_), .ZN(new_n15937_));
  AOI21_X1   g15681(.A1(new_n15936_), .A2(new_n15704_), .B(new_n15937_), .ZN(new_n15938_));
  OAI22_X1   g15682(.A1(new_n10390_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n10389_), .ZN(new_n15939_));
  AOI21_X1   g15683(.A1(\b[23] ), .A2(new_n9471_), .B(new_n15939_), .ZN(new_n15940_));
  OAI21_X1   g15684(.A1(new_n2655_), .A2(new_n10388_), .B(new_n15940_), .ZN(new_n15941_));
  XOR2_X1    g15685(.A1(new_n15941_), .A2(\a[53] ), .Z(new_n15942_));
  NOR2_X1    g15686(.A1(new_n15938_), .A2(new_n15942_), .ZN(new_n15943_));
  INV_X1     g15687(.I(new_n15943_), .ZN(new_n15944_));
  NAND2_X1   g15688(.A1(new_n15938_), .A2(new_n15942_), .ZN(new_n15945_));
  NAND2_X1   g15689(.A1(new_n15944_), .A2(new_n15945_), .ZN(new_n15946_));
  XOR2_X1    g15690(.A1(new_n15946_), .A2(new_n15935_), .Z(new_n15947_));
  NOR2_X1    g15691(.A1(new_n15663_), .A2(new_n15707_), .ZN(new_n15948_));
  NOR2_X1    g15692(.A1(new_n15948_), .A2(new_n15708_), .ZN(new_n15949_));
  NOR2_X1    g15693(.A1(new_n15949_), .A2(new_n15947_), .ZN(new_n15950_));
  INV_X1     g15694(.I(new_n15950_), .ZN(new_n15951_));
  NAND2_X1   g15695(.A1(new_n15949_), .A2(new_n15947_), .ZN(new_n15952_));
  NAND2_X1   g15696(.A1(new_n15951_), .A2(new_n15952_), .ZN(new_n15953_));
  XOR2_X1    g15697(.A1(new_n15953_), .A2(new_n15899_), .Z(new_n15954_));
  INV_X1     g15698(.I(new_n15954_), .ZN(new_n15955_));
  NAND2_X1   g15699(.A1(new_n15955_), .A2(new_n15895_), .ZN(new_n15956_));
  NOR2_X1    g15700(.A1(new_n15955_), .A2(new_n15895_), .ZN(new_n15957_));
  INV_X1     g15701(.I(new_n15957_), .ZN(new_n15958_));
  NAND2_X1   g15702(.A1(new_n15958_), .A2(new_n15956_), .ZN(new_n15959_));
  XNOR2_X1   g15703(.A1(new_n15959_), .A2(new_n15893_), .ZN(new_n15960_));
  NOR2_X1    g15704(.A1(new_n15960_), .A2(new_n15889_), .ZN(new_n15961_));
  NAND2_X1   g15705(.A1(new_n15960_), .A2(new_n15889_), .ZN(new_n15962_));
  INV_X1     g15706(.I(new_n15962_), .ZN(new_n15963_));
  NOR2_X1    g15707(.A1(new_n15963_), .A2(new_n15961_), .ZN(new_n15964_));
  XOR2_X1    g15708(.A1(new_n15964_), .A2(new_n15886_), .Z(new_n15965_));
  NAND2_X1   g15709(.A1(new_n15965_), .A2(new_n15882_), .ZN(new_n15966_));
  OR2_X2     g15710(.A1(new_n15965_), .A2(new_n15882_), .Z(new_n15967_));
  NAND2_X1   g15711(.A1(new_n15967_), .A2(new_n15966_), .ZN(new_n15968_));
  XOR2_X1    g15712(.A1(new_n15968_), .A2(new_n15880_), .Z(new_n15969_));
  NAND2_X1   g15713(.A1(new_n15969_), .A2(new_n15876_), .ZN(new_n15970_));
  OR2_X2     g15714(.A1(new_n15969_), .A2(new_n15876_), .Z(new_n15971_));
  NAND2_X1   g15715(.A1(new_n15971_), .A2(new_n15970_), .ZN(new_n15972_));
  XOR2_X1    g15716(.A1(new_n15972_), .A2(new_n15874_), .Z(new_n15973_));
  OAI22_X1   g15717(.A1(new_n6775_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n6490_), .ZN(new_n15974_));
  AOI21_X1   g15718(.A1(\b[41] ), .A2(new_n4706_), .B(new_n15974_), .ZN(new_n15975_));
  OAI21_X1   g15719(.A1(new_n6785_), .A2(new_n4458_), .B(new_n15975_), .ZN(new_n15976_));
  XOR2_X1    g15720(.A1(new_n15976_), .A2(\a[35] ), .Z(new_n15977_));
  XOR2_X1    g15721(.A1(new_n15973_), .A2(new_n15977_), .Z(new_n15978_));
  XOR2_X1    g15722(.A1(new_n15978_), .A2(new_n15870_), .Z(new_n15979_));
  XOR2_X1    g15723(.A1(new_n15979_), .A2(new_n3876_), .Z(new_n15980_));
  XOR2_X1    g15724(.A1(new_n15980_), .A2(new_n15868_), .Z(new_n15981_));
  OAI22_X1   g15725(.A1(new_n8168_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n8127_), .ZN(new_n15982_));
  AOI21_X1   g15726(.A1(\b[47] ), .A2(new_n3456_), .B(new_n15982_), .ZN(new_n15983_));
  OAI21_X1   g15727(.A1(new_n9050_), .A2(new_n3261_), .B(new_n15983_), .ZN(new_n15984_));
  XOR2_X1    g15728(.A1(new_n15984_), .A2(\a[29] ), .Z(new_n15985_));
  INV_X1     g15729(.I(new_n15985_), .ZN(new_n15986_));
  NAND2_X1   g15730(.A1(new_n15981_), .A2(new_n15986_), .ZN(new_n15987_));
  OR2_X2     g15731(.A1(new_n15981_), .A2(new_n15986_), .Z(new_n15988_));
  NAND2_X1   g15732(.A1(new_n15988_), .A2(new_n15987_), .ZN(new_n15989_));
  XOR2_X1    g15733(.A1(new_n15989_), .A2(new_n15862_), .Z(new_n15990_));
  AOI22_X1   g15734(.A1(new_n2716_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n2719_), .ZN(new_n15991_));
  OAI21_X1   g15735(.A1(new_n8500_), .A2(new_n2924_), .B(new_n15991_), .ZN(new_n15992_));
  AOI21_X1   g15736(.A1(new_n9987_), .A2(new_n2722_), .B(new_n15992_), .ZN(new_n15993_));
  XOR2_X1    g15737(.A1(new_n15993_), .A2(new_n2714_), .Z(new_n15994_));
  OR2_X2     g15738(.A1(new_n15990_), .A2(new_n15994_), .Z(new_n15995_));
  NAND2_X1   g15739(.A1(new_n15990_), .A2(new_n15994_), .ZN(new_n15996_));
  NAND2_X1   g15740(.A1(new_n15995_), .A2(new_n15996_), .ZN(new_n15997_));
  XOR2_X1    g15741(.A1(new_n15997_), .A2(new_n15859_), .Z(new_n15998_));
  AOI22_X1   g15742(.A1(new_n2202_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n2205_), .ZN(new_n15999_));
  OAI21_X1   g15743(.A1(new_n9376_), .A2(new_n2370_), .B(new_n15999_), .ZN(new_n16000_));
  AOI21_X1   g15744(.A1(new_n9979_), .A2(new_n2208_), .B(new_n16000_), .ZN(new_n16001_));
  XOR2_X1    g15745(.A1(new_n16001_), .A2(new_n2200_), .Z(new_n16002_));
  OR2_X2     g15746(.A1(new_n15998_), .A2(new_n16002_), .Z(new_n16003_));
  NAND2_X1   g15747(.A1(new_n15998_), .A2(new_n16002_), .ZN(new_n16004_));
  NAND2_X1   g15748(.A1(new_n16003_), .A2(new_n16004_), .ZN(new_n16005_));
  XOR2_X1    g15749(.A1(new_n16005_), .A2(new_n15856_), .Z(new_n16006_));
  XOR2_X1    g15750(.A1(new_n16006_), .A2(new_n15853_), .Z(new_n16007_));
  XOR2_X1    g15751(.A1(new_n16007_), .A2(new_n15851_), .Z(new_n16008_));
  OAI22_X1   g15752(.A1(new_n1592_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n1505_), .ZN(new_n16009_));
  AOI21_X1   g15753(.A1(\b[59] ), .A2(new_n1584_), .B(new_n16009_), .ZN(new_n16010_));
  OAI21_X1   g15754(.A1(new_n13110_), .A2(new_n1732_), .B(new_n16010_), .ZN(new_n16011_));
  XOR2_X1    g15755(.A1(new_n16011_), .A2(\a[17] ), .Z(new_n16012_));
  OR2_X2     g15756(.A1(new_n16008_), .A2(new_n16012_), .Z(new_n16013_));
  NAND2_X1   g15757(.A1(new_n16008_), .A2(new_n16012_), .ZN(new_n16014_));
  NAND2_X1   g15758(.A1(new_n16013_), .A2(new_n16014_), .ZN(new_n16015_));
  XOR2_X1    g15759(.A1(new_n16015_), .A2(new_n15847_), .Z(new_n16016_));
  AOI22_X1   g15760(.A1(new_n1486_), .A2(\b[62] ), .B1(\b[63] ), .B2(new_n1009_), .ZN(new_n16017_));
  OAI21_X1   g15761(.A1(new_n13107_), .A2(new_n1323_), .B(new_n16017_), .ZN(new_n16018_));
  XOR2_X1    g15762(.A1(new_n16018_), .A2(\a[14] ), .Z(new_n16019_));
  OR2_X2     g15763(.A1(new_n16016_), .A2(new_n16019_), .Z(new_n16020_));
  NAND2_X1   g15764(.A1(new_n16016_), .A2(new_n16019_), .ZN(new_n16021_));
  NAND2_X1   g15765(.A1(new_n16020_), .A2(new_n16021_), .ZN(new_n16022_));
  XOR2_X1    g15766(.A1(new_n16022_), .A2(new_n15844_), .Z(new_n16023_));
  OR2_X2     g15767(.A1(new_n15834_), .A2(new_n15635_), .Z(new_n16024_));
  NAND2_X1   g15768(.A1(new_n15834_), .A2(new_n15635_), .ZN(new_n16025_));
  INV_X1     g15769(.I(new_n16025_), .ZN(new_n16026_));
  NOR2_X1    g15770(.A1(new_n15630_), .A2(new_n15628_), .ZN(new_n16027_));
  OAI21_X1   g15771(.A1(new_n15416_), .A2(new_n16027_), .B(new_n15631_), .ZN(new_n16028_));
  AOI21_X1   g15772(.A1(new_n16028_), .A2(new_n16024_), .B(new_n16026_), .ZN(new_n16029_));
  NOR2_X1    g15773(.A1(new_n16029_), .A2(new_n16023_), .ZN(new_n16030_));
  INV_X1     g15774(.I(new_n15844_), .ZN(new_n16031_));
  XOR2_X1    g15775(.A1(new_n16022_), .A2(new_n16031_), .Z(new_n16032_));
  OAI21_X1   g15776(.A1(new_n15839_), .A2(new_n15835_), .B(new_n16025_), .ZN(new_n16033_));
  NOR2_X1    g15777(.A1(new_n16033_), .A2(new_n16032_), .ZN(new_n16034_));
  NOR2_X1    g15778(.A1(new_n16030_), .A2(new_n16034_), .ZN(new_n16035_));
  XOR2_X1    g15779(.A1(new_n16035_), .A2(new_n15842_), .Z(\f[76] ));
  NAND2_X1   g15780(.A1(new_n16029_), .A2(new_n16023_), .ZN(new_n16037_));
  INV_X1     g15781(.I(new_n15842_), .ZN(new_n16038_));
  OAI21_X1   g15782(.A1(new_n16029_), .A2(new_n16023_), .B(new_n16038_), .ZN(new_n16039_));
  NAND2_X1   g15783(.A1(new_n16039_), .A2(new_n16037_), .ZN(new_n16040_));
  NAND2_X1   g15784(.A1(new_n16021_), .A2(new_n16031_), .ZN(new_n16041_));
  NAND2_X1   g15785(.A1(new_n16041_), .A2(new_n16020_), .ZN(new_n16042_));
  OAI22_X1   g15786(.A1(new_n13462_), .A2(new_n1323_), .B1(new_n12800_), .B2(new_n1481_), .ZN(new_n16043_));
  XOR2_X1    g15787(.A1(new_n16043_), .A2(\a[14] ), .Z(new_n16044_));
  NAND2_X1   g15788(.A1(new_n16014_), .A2(new_n15847_), .ZN(new_n16045_));
  NAND2_X1   g15789(.A1(new_n16045_), .A2(new_n16013_), .ZN(new_n16046_));
  INV_X1     g15790(.I(new_n16046_), .ZN(new_n16047_));
  OAI22_X1   g15791(.A1(new_n1592_), .A2(new_n12796_), .B1(new_n12148_), .B2(new_n1505_), .ZN(new_n16048_));
  AOI21_X1   g15792(.A1(\b[60] ), .A2(new_n1584_), .B(new_n16048_), .ZN(new_n16049_));
  OAI21_X1   g15793(.A1(new_n14950_), .A2(new_n1732_), .B(new_n16049_), .ZN(new_n16050_));
  XOR2_X1    g15794(.A1(new_n16050_), .A2(new_n1344_), .Z(new_n16051_));
  INV_X1     g15795(.I(new_n15851_), .ZN(new_n16052_));
  NOR2_X1    g15796(.A1(new_n16006_), .A2(new_n15853_), .ZN(new_n16053_));
  NAND2_X1   g15797(.A1(new_n16006_), .A2(new_n15853_), .ZN(new_n16054_));
  AOI21_X1   g15798(.A1(new_n16052_), .A2(new_n16054_), .B(new_n16053_), .ZN(new_n16055_));
  INV_X1     g15799(.I(new_n16003_), .ZN(new_n16056_));
  AOI21_X1   g15800(.A1(new_n15856_), .A2(new_n16004_), .B(new_n16056_), .ZN(new_n16057_));
  OAI22_X1   g15801(.A1(new_n1751_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n1754_), .ZN(new_n16058_));
  AOI21_X1   g15802(.A1(\b[57] ), .A2(new_n1939_), .B(new_n16058_), .ZN(new_n16059_));
  OAI21_X1   g15803(.A1(new_n12203_), .A2(new_n1757_), .B(new_n16059_), .ZN(new_n16060_));
  XOR2_X1    g15804(.A1(new_n16060_), .A2(\a[20] ), .Z(new_n16061_));
  INV_X1     g15805(.I(new_n16061_), .ZN(new_n16062_));
  NAND2_X1   g15806(.A1(new_n15996_), .A2(new_n15859_), .ZN(new_n16063_));
  AND2_X2    g15807(.A1(new_n16063_), .A2(new_n15995_), .Z(new_n16064_));
  NAND2_X1   g15808(.A1(new_n15988_), .A2(new_n15862_), .ZN(new_n16065_));
  AND2_X2    g15809(.A1(new_n16065_), .A2(new_n15987_), .Z(new_n16066_));
  OAI22_X1   g15810(.A1(new_n2703_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n2708_), .ZN(new_n16067_));
  AOI21_X1   g15811(.A1(\b[51] ), .A2(new_n2906_), .B(new_n16067_), .ZN(new_n16068_));
  OAI21_X1   g15812(.A1(new_n9385_), .A2(new_n2711_), .B(new_n16068_), .ZN(new_n16069_));
  XOR2_X1    g15813(.A1(new_n16069_), .A2(\a[26] ), .Z(new_n16070_));
  INV_X1     g15814(.I(new_n16070_), .ZN(new_n16071_));
  INV_X1     g15815(.I(new_n15979_), .ZN(new_n16072_));
  NOR2_X1    g15816(.A1(new_n16072_), .A2(new_n15864_), .ZN(new_n16073_));
  NAND2_X1   g15817(.A1(new_n16072_), .A2(new_n15864_), .ZN(new_n16074_));
  XOR2_X1    g15818(.A1(new_n15867_), .A2(new_n3876_), .Z(new_n16075_));
  INV_X1     g15819(.I(new_n16075_), .ZN(new_n16076_));
  AOI21_X1   g15820(.A1(new_n16074_), .A2(new_n16076_), .B(new_n16073_), .ZN(new_n16077_));
  AOI22_X1   g15821(.A1(new_n3267_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n3270_), .ZN(new_n16078_));
  OAI21_X1   g15822(.A1(new_n8127_), .A2(new_n3475_), .B(new_n16078_), .ZN(new_n16079_));
  NOR2_X1    g15823(.A1(new_n8510_), .A2(new_n3261_), .ZN(new_n16080_));
  NOR2_X1    g15824(.A1(new_n16080_), .A2(new_n16079_), .ZN(new_n16081_));
  XNOR2_X1   g15825(.A1(new_n16077_), .A2(new_n16081_), .ZN(new_n16082_));
  AOI22_X1   g15826(.A1(new_n3864_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n3869_), .ZN(new_n16083_));
  OAI21_X1   g15827(.A1(new_n7096_), .A2(new_n5410_), .B(new_n16083_), .ZN(new_n16084_));
  AOI21_X1   g15828(.A1(new_n7649_), .A2(new_n3872_), .B(new_n16084_), .ZN(new_n16085_));
  XOR2_X1    g15829(.A1(new_n16085_), .A2(new_n3876_), .Z(new_n16086_));
  INV_X1     g15830(.I(new_n16086_), .ZN(new_n16087_));
  INV_X1     g15831(.I(new_n15977_), .ZN(new_n16088_));
  NAND2_X1   g15832(.A1(new_n15973_), .A2(new_n16088_), .ZN(new_n16089_));
  NOR2_X1    g15833(.A1(new_n15973_), .A2(new_n16088_), .ZN(new_n16090_));
  OAI21_X1   g15834(.A1(new_n15870_), .A2(new_n16090_), .B(new_n16089_), .ZN(new_n16091_));
  AOI22_X1   g15835(.A1(new_n4918_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n4921_), .ZN(new_n16092_));
  OAI21_X1   g15836(.A1(new_n6490_), .A2(new_n6099_), .B(new_n16092_), .ZN(new_n16093_));
  AOI21_X1   g15837(.A1(new_n7906_), .A2(new_n4699_), .B(new_n16093_), .ZN(new_n16094_));
  XOR2_X1    g15838(.A1(new_n16094_), .A2(new_n4446_), .Z(new_n16095_));
  INV_X1     g15839(.I(new_n15970_), .ZN(new_n16096_));
  OAI21_X1   g15840(.A1(new_n15874_), .A2(new_n16096_), .B(new_n15971_), .ZN(new_n16097_));
  OAI22_X1   g15841(.A1(new_n6285_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n6284_), .ZN(new_n16098_));
  AOI21_X1   g15842(.A1(\b[39] ), .A2(new_n5420_), .B(new_n16098_), .ZN(new_n16099_));
  OAI21_X1   g15843(.A1(new_n6299_), .A2(new_n6124_), .B(new_n16099_), .ZN(new_n16100_));
  XOR2_X1    g15844(.A1(new_n16100_), .A2(new_n5162_), .Z(new_n16101_));
  AOI22_X1   g15845(.A1(new_n6108_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n6111_), .ZN(new_n16102_));
  OAI21_X1   g15846(.A1(new_n4886_), .A2(new_n7708_), .B(new_n16102_), .ZN(new_n16103_));
  AOI21_X1   g15847(.A1(new_n5351_), .A2(new_n6105_), .B(new_n16103_), .ZN(new_n16104_));
  XOR2_X1    g15848(.A1(new_n16104_), .A2(new_n5849_), .Z(new_n16105_));
  AOI22_X1   g15849(.A1(new_n7403_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n7408_), .ZN(new_n16106_));
  OAI21_X1   g15850(.A1(new_n3624_), .A2(new_n9488_), .B(new_n16106_), .ZN(new_n16107_));
  AOI21_X1   g15851(.A1(new_n4030_), .A2(new_n7414_), .B(new_n16107_), .ZN(new_n16108_));
  XOR2_X1    g15852(.A1(new_n16108_), .A2(new_n7410_), .Z(new_n16109_));
  AOI22_X1   g15853(.A1(new_n9125_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n9123_), .ZN(new_n16110_));
  OAI21_X1   g15854(.A1(new_n2495_), .A2(new_n9470_), .B(new_n16110_), .ZN(new_n16111_));
  AOI21_X1   g15855(.A1(new_n3407_), .A2(new_n9129_), .B(new_n16111_), .ZN(new_n16112_));
  XOR2_X1    g15856(.A1(new_n16112_), .A2(new_n9133_), .Z(new_n16113_));
  AOI21_X1   g15857(.A1(new_n15904_), .A2(new_n15932_), .B(new_n15930_), .ZN(new_n16114_));
  INV_X1     g15858(.I(new_n16114_), .ZN(new_n16115_));
  AOI22_X1   g15859(.A1(new_n10064_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n10062_), .ZN(new_n16116_));
  OAI21_X1   g15860(.A1(new_n2027_), .A2(new_n10399_), .B(new_n16116_), .ZN(new_n16117_));
  AOI21_X1   g15861(.A1(new_n2470_), .A2(new_n10068_), .B(new_n16117_), .ZN(new_n16118_));
  XOR2_X1    g15862(.A1(new_n16118_), .A2(new_n10057_), .Z(new_n16119_));
  AOI21_X1   g15863(.A1(new_n15915_), .A2(new_n15924_), .B(new_n15922_), .ZN(new_n16120_));
  NOR2_X1    g15864(.A1(new_n16119_), .A2(new_n16120_), .ZN(new_n16121_));
  INV_X1     g15865(.I(new_n16121_), .ZN(new_n16122_));
  NAND2_X1   g15866(.A1(new_n16119_), .A2(new_n16120_), .ZN(new_n16123_));
  NAND2_X1   g15867(.A1(new_n16122_), .A2(new_n16123_), .ZN(new_n16124_));
  AOI22_X1   g15868(.A1(new_n10981_), .A2(\b[20] ), .B1(new_n10979_), .B2(\b[19] ), .ZN(new_n16125_));
  OAI21_X1   g15869(.A1(new_n1553_), .A2(new_n11306_), .B(new_n16125_), .ZN(new_n16126_));
  AOI21_X1   g15870(.A1(new_n2452_), .A2(new_n10984_), .B(new_n16126_), .ZN(new_n16127_));
  XOR2_X1    g15871(.A1(new_n16127_), .A2(new_n10989_), .Z(new_n16128_));
  NOR2_X1    g15872(.A1(new_n15910_), .A2(new_n15911_), .ZN(new_n16129_));
  NAND2_X1   g15873(.A1(new_n15910_), .A2(new_n15911_), .ZN(new_n16130_));
  AOI21_X1   g15874(.A1(new_n15908_), .A2(new_n16130_), .B(new_n16129_), .ZN(new_n16131_));
  INV_X1     g15875(.I(new_n16131_), .ZN(new_n16132_));
  OAI22_X1   g15876(.A1(new_n13224_), .A2(new_n1432_), .B1(new_n1296_), .B2(new_n11923_), .ZN(new_n16133_));
  AOI21_X1   g15877(.A1(\b[15] ), .A2(new_n13223_), .B(new_n16133_), .ZN(new_n16134_));
  OAI21_X1   g15878(.A1(new_n1444_), .A2(new_n11930_), .B(new_n16134_), .ZN(new_n16135_));
  XOR2_X1    g15879(.A1(new_n16135_), .A2(\a[62] ), .Z(new_n16136_));
  AOI22_X1   g15880(.A1(new_n12922_), .A2(\b[14] ), .B1(\b[13] ), .B2(new_n12923_), .ZN(new_n16137_));
  INV_X1     g15881(.I(new_n16137_), .ZN(new_n16138_));
  NOR2_X1    g15882(.A1(new_n16138_), .A2(new_n15911_), .ZN(new_n16139_));
  NOR2_X1    g15883(.A1(new_n15912_), .A2(new_n16137_), .ZN(new_n16140_));
  NOR2_X1    g15884(.A1(new_n16139_), .A2(new_n16140_), .ZN(new_n16141_));
  XNOR2_X1   g15885(.A1(new_n16136_), .A2(new_n16141_), .ZN(new_n16142_));
  NOR2_X1    g15886(.A1(new_n16142_), .A2(new_n16132_), .ZN(new_n16143_));
  INV_X1     g15887(.I(new_n16143_), .ZN(new_n16144_));
  NAND2_X1   g15888(.A1(new_n16142_), .A2(new_n16132_), .ZN(new_n16145_));
  NAND2_X1   g15889(.A1(new_n16144_), .A2(new_n16145_), .ZN(new_n16146_));
  XOR2_X1    g15890(.A1(new_n16146_), .A2(new_n16128_), .Z(new_n16147_));
  XNOR2_X1   g15891(.A1(new_n16124_), .A2(new_n16147_), .ZN(new_n16148_));
  NOR2_X1    g15892(.A1(new_n16148_), .A2(new_n16115_), .ZN(new_n16149_));
  INV_X1     g15893(.I(new_n16149_), .ZN(new_n16150_));
  NAND2_X1   g15894(.A1(new_n16148_), .A2(new_n16115_), .ZN(new_n16151_));
  NAND2_X1   g15895(.A1(new_n16150_), .A2(new_n16151_), .ZN(new_n16152_));
  XOR2_X1    g15896(.A1(new_n16152_), .A2(new_n16113_), .Z(new_n16153_));
  AOI22_X1   g15897(.A1(new_n8241_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n8246_), .ZN(new_n16154_));
  OAI21_X1   g15898(.A1(new_n3158_), .A2(new_n9114_), .B(new_n16154_), .ZN(new_n16155_));
  AOI21_X1   g15899(.A1(new_n4188_), .A2(new_n8252_), .B(new_n16155_), .ZN(new_n16156_));
  XOR2_X1    g15900(.A1(new_n16156_), .A2(new_n8248_), .Z(new_n16157_));
  AOI21_X1   g15901(.A1(new_n15935_), .A2(new_n15945_), .B(new_n15943_), .ZN(new_n16158_));
  NOR2_X1    g15902(.A1(new_n16157_), .A2(new_n16158_), .ZN(new_n16159_));
  INV_X1     g15903(.I(new_n16159_), .ZN(new_n16160_));
  NAND2_X1   g15904(.A1(new_n16157_), .A2(new_n16158_), .ZN(new_n16161_));
  NAND2_X1   g15905(.A1(new_n16160_), .A2(new_n16161_), .ZN(new_n16162_));
  XOR2_X1    g15906(.A1(new_n16162_), .A2(new_n16153_), .Z(new_n16163_));
  INV_X1     g15907(.I(new_n16163_), .ZN(new_n16164_));
  INV_X1     g15908(.I(new_n15899_), .ZN(new_n16165_));
  AOI21_X1   g15909(.A1(new_n16165_), .A2(new_n15952_), .B(new_n15950_), .ZN(new_n16166_));
  INV_X1     g15910(.I(new_n16166_), .ZN(new_n16167_));
  NAND2_X1   g15911(.A1(new_n16164_), .A2(new_n16167_), .ZN(new_n16168_));
  NOR2_X1    g15912(.A1(new_n16164_), .A2(new_n16167_), .ZN(new_n16169_));
  INV_X1     g15913(.I(new_n16169_), .ZN(new_n16170_));
  NAND2_X1   g15914(.A1(new_n16170_), .A2(new_n16168_), .ZN(new_n16171_));
  XNOR2_X1   g15915(.A1(new_n16171_), .A2(new_n16109_), .ZN(new_n16172_));
  INV_X1     g15916(.I(new_n16172_), .ZN(new_n16173_));
  OAI22_X1   g15917(.A1(new_n7730_), .A2(new_n4666_), .B1(new_n4639_), .B2(new_n7731_), .ZN(new_n16174_));
  AOI21_X1   g15918(.A1(\b[33] ), .A2(new_n6887_), .B(new_n16174_), .ZN(new_n16175_));
  OAI21_X1   g15919(.A1(new_n4676_), .A2(new_n7728_), .B(new_n16175_), .ZN(new_n16176_));
  XOR2_X1    g15920(.A1(new_n16176_), .A2(\a[44] ), .Z(new_n16177_));
  AOI21_X1   g15921(.A1(new_n15893_), .A2(new_n15956_), .B(new_n15957_), .ZN(new_n16178_));
  NOR2_X1    g15922(.A1(new_n16177_), .A2(new_n16178_), .ZN(new_n16179_));
  INV_X1     g15923(.I(new_n16179_), .ZN(new_n16180_));
  NAND2_X1   g15924(.A1(new_n16177_), .A2(new_n16178_), .ZN(new_n16181_));
  NAND2_X1   g15925(.A1(new_n16180_), .A2(new_n16181_), .ZN(new_n16182_));
  XOR2_X1    g15926(.A1(new_n16182_), .A2(new_n16173_), .Z(new_n16183_));
  OAI21_X1   g15927(.A1(new_n15886_), .A2(new_n15961_), .B(new_n15962_), .ZN(new_n16184_));
  INV_X1     g15928(.I(new_n16184_), .ZN(new_n16185_));
  NOR2_X1    g15929(.A1(new_n16185_), .A2(new_n16183_), .ZN(new_n16186_));
  INV_X1     g15930(.I(new_n16186_), .ZN(new_n16187_));
  NAND2_X1   g15931(.A1(new_n16185_), .A2(new_n16183_), .ZN(new_n16188_));
  NAND2_X1   g15932(.A1(new_n16187_), .A2(new_n16188_), .ZN(new_n16189_));
  XOR2_X1    g15933(.A1(new_n16189_), .A2(new_n16105_), .Z(new_n16190_));
  INV_X1     g15934(.I(new_n16190_), .ZN(new_n16191_));
  INV_X1     g15935(.I(new_n15967_), .ZN(new_n16192_));
  AOI21_X1   g15936(.A1(new_n15880_), .A2(new_n15966_), .B(new_n16192_), .ZN(new_n16193_));
  NOR2_X1    g15937(.A1(new_n16193_), .A2(new_n16191_), .ZN(new_n16194_));
  INV_X1     g15938(.I(new_n16194_), .ZN(new_n16195_));
  NAND2_X1   g15939(.A1(new_n16193_), .A2(new_n16191_), .ZN(new_n16196_));
  NAND2_X1   g15940(.A1(new_n16195_), .A2(new_n16196_), .ZN(new_n16197_));
  XNOR2_X1   g15941(.A1(new_n16197_), .A2(new_n16101_), .ZN(new_n16198_));
  OR2_X2     g15942(.A1(new_n16198_), .A2(new_n16097_), .Z(new_n16199_));
  NAND2_X1   g15943(.A1(new_n16198_), .A2(new_n16097_), .ZN(new_n16200_));
  NAND2_X1   g15944(.A1(new_n16199_), .A2(new_n16200_), .ZN(new_n16201_));
  XOR2_X1    g15945(.A1(new_n16201_), .A2(new_n16095_), .Z(new_n16202_));
  NAND2_X1   g15946(.A1(new_n16202_), .A2(new_n16091_), .ZN(new_n16203_));
  OR2_X2     g15947(.A1(new_n16202_), .A2(new_n16091_), .Z(new_n16204_));
  NAND2_X1   g15948(.A1(new_n16204_), .A2(new_n16203_), .ZN(new_n16205_));
  XOR2_X1    g15949(.A1(new_n16205_), .A2(new_n16087_), .Z(new_n16206_));
  XOR2_X1    g15950(.A1(new_n16206_), .A2(new_n3264_), .Z(new_n16207_));
  XOR2_X1    g15951(.A1(new_n16207_), .A2(new_n16082_), .Z(new_n16208_));
  NAND2_X1   g15952(.A1(new_n16208_), .A2(new_n16071_), .ZN(new_n16209_));
  OR2_X2     g15953(.A1(new_n16208_), .A2(new_n16071_), .Z(new_n16210_));
  NAND2_X1   g15954(.A1(new_n16210_), .A2(new_n16209_), .ZN(new_n16211_));
  XOR2_X1    g15955(.A1(new_n16211_), .A2(new_n16066_), .Z(new_n16212_));
  XOR2_X1    g15956(.A1(new_n16212_), .A2(new_n16064_), .Z(new_n16213_));
  AOI22_X1   g15957(.A1(new_n2202_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n2205_), .ZN(new_n16214_));
  OAI21_X1   g15958(.A1(new_n9942_), .A2(new_n2370_), .B(new_n16214_), .ZN(new_n16215_));
  AOI21_X1   g15959(.A1(new_n10318_), .A2(new_n2208_), .B(new_n16215_), .ZN(new_n16216_));
  XOR2_X1    g15960(.A1(new_n16216_), .A2(new_n2200_), .Z(new_n16217_));
  XOR2_X1    g15961(.A1(new_n16213_), .A2(new_n16217_), .Z(new_n16218_));
  AND2_X2    g15962(.A1(new_n16218_), .A2(new_n16062_), .Z(new_n16219_));
  NOR2_X1    g15963(.A1(new_n16218_), .A2(new_n16062_), .ZN(new_n16220_));
  NOR2_X1    g15964(.A1(new_n16219_), .A2(new_n16220_), .ZN(new_n16221_));
  XOR2_X1    g15965(.A1(new_n16221_), .A2(new_n16057_), .Z(new_n16222_));
  OR2_X2     g15966(.A1(new_n16222_), .A2(new_n16055_), .Z(new_n16223_));
  NAND2_X1   g15967(.A1(new_n16222_), .A2(new_n16055_), .ZN(new_n16224_));
  NAND2_X1   g15968(.A1(new_n16223_), .A2(new_n16224_), .ZN(new_n16225_));
  XNOR2_X1   g15969(.A1(new_n16225_), .A2(new_n16051_), .ZN(new_n16226_));
  XOR2_X1    g15970(.A1(new_n16226_), .A2(new_n16047_), .Z(new_n16227_));
  XOR2_X1    g15971(.A1(new_n16227_), .A2(new_n16044_), .Z(new_n16228_));
  NOR2_X1    g15972(.A1(new_n16228_), .A2(new_n16042_), .ZN(new_n16229_));
  INV_X1     g15973(.I(new_n16229_), .ZN(new_n16230_));
  NAND2_X1   g15974(.A1(new_n16228_), .A2(new_n16042_), .ZN(new_n16231_));
  NAND2_X1   g15975(.A1(new_n16230_), .A2(new_n16231_), .ZN(new_n16232_));
  XOR2_X1    g15976(.A1(new_n16040_), .A2(new_n16232_), .Z(\f[77] ));
  INV_X1     g15977(.I(new_n16231_), .ZN(new_n16234_));
  AOI21_X1   g15978(.A1(new_n16039_), .A2(new_n16037_), .B(new_n16229_), .ZN(new_n16235_));
  NOR2_X1    g15979(.A1(new_n16235_), .A2(new_n16234_), .ZN(new_n16236_));
  INV_X1     g15980(.I(new_n16226_), .ZN(new_n16237_));
  AOI21_X1   g15981(.A1(new_n16237_), .A2(new_n16047_), .B(new_n16044_), .ZN(new_n16238_));
  AOI21_X1   g15982(.A1(new_n16046_), .A2(new_n16226_), .B(new_n16238_), .ZN(new_n16239_));
  INV_X1     g15983(.I(new_n16223_), .ZN(new_n16240_));
  AOI21_X1   g15984(.A1(new_n16051_), .A2(new_n16224_), .B(new_n16240_), .ZN(new_n16241_));
  NOR2_X1    g15985(.A1(new_n16220_), .A2(new_n16057_), .ZN(new_n16242_));
  NOR2_X1    g15986(.A1(new_n16242_), .A2(new_n16219_), .ZN(new_n16243_));
  INV_X1     g15987(.I(new_n16243_), .ZN(new_n16244_));
  INV_X1     g15988(.I(new_n16064_), .ZN(new_n16245_));
  NAND2_X1   g15989(.A1(new_n16212_), .A2(new_n16245_), .ZN(new_n16246_));
  NOR2_X1    g15990(.A1(new_n16212_), .A2(new_n16245_), .ZN(new_n16247_));
  OAI21_X1   g15991(.A1(new_n16217_), .A2(new_n16247_), .B(new_n16246_), .ZN(new_n16248_));
  INV_X1     g15992(.I(new_n16066_), .ZN(new_n16249_));
  NAND2_X1   g15993(.A1(new_n16210_), .A2(new_n16249_), .ZN(new_n16250_));
  AND2_X2    g15994(.A1(new_n16250_), .A2(new_n16209_), .Z(new_n16251_));
  AOI22_X1   g15995(.A1(new_n2716_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n2719_), .ZN(new_n16252_));
  OAI21_X1   g15996(.A1(new_n9032_), .A2(new_n2924_), .B(new_n16252_), .ZN(new_n16253_));
  AOI21_X1   g15997(.A1(new_n10884_), .A2(new_n2722_), .B(new_n16253_), .ZN(new_n16254_));
  XOR2_X1    g15998(.A1(new_n16254_), .A2(new_n2714_), .Z(new_n16255_));
  INV_X1     g15999(.I(new_n16255_), .ZN(new_n16256_));
  INV_X1     g16000(.I(new_n16077_), .ZN(new_n16257_));
  INV_X1     g16001(.I(new_n16206_), .ZN(new_n16258_));
  NAND2_X1   g16002(.A1(new_n16258_), .A2(new_n16257_), .ZN(new_n16259_));
  NOR2_X1    g16003(.A1(new_n16258_), .A2(new_n16257_), .ZN(new_n16260_));
  XOR2_X1    g16004(.A1(new_n16081_), .A2(new_n3264_), .Z(new_n16261_));
  OAI21_X1   g16005(.A1(new_n16260_), .A2(new_n16261_), .B(new_n16259_), .ZN(new_n16262_));
  AOI22_X1   g16006(.A1(new_n3267_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n3270_), .ZN(new_n16263_));
  OAI21_X1   g16007(.A1(new_n8168_), .A2(new_n3475_), .B(new_n16263_), .ZN(new_n16264_));
  AOI21_X1   g16008(.A1(new_n8783_), .A2(new_n3273_), .B(new_n16264_), .ZN(new_n16265_));
  XOR2_X1    g16009(.A1(new_n16265_), .A2(\a[29] ), .Z(new_n16266_));
  INV_X1     g16010(.I(new_n16199_), .ZN(new_n16267_));
  OAI21_X1   g16011(.A1(new_n16267_), .A2(new_n16095_), .B(new_n16200_), .ZN(new_n16268_));
  AOI21_X1   g16012(.A1(new_n16101_), .A2(new_n16196_), .B(new_n16194_), .ZN(new_n16269_));
  INV_X1     g16013(.I(new_n16269_), .ZN(new_n16270_));
  INV_X1     g16014(.I(new_n16105_), .ZN(new_n16271_));
  AOI21_X1   g16015(.A1(new_n16271_), .A2(new_n16188_), .B(new_n16186_), .ZN(new_n16272_));
  AOI21_X1   g16016(.A1(new_n16173_), .A2(new_n16181_), .B(new_n16179_), .ZN(new_n16273_));
  INV_X1     g16017(.I(new_n16273_), .ZN(new_n16274_));
  AOI22_X1   g16018(.A1(new_n6569_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n6574_), .ZN(new_n16275_));
  OAI21_X1   g16019(.A1(new_n4639_), .A2(new_n8565_), .B(new_n16275_), .ZN(new_n16276_));
  AOI21_X1   g16020(.A1(new_n5594_), .A2(new_n6579_), .B(new_n16276_), .ZN(new_n16277_));
  XOR2_X1    g16021(.A1(new_n16277_), .A2(new_n6567_), .Z(new_n16278_));
  OAI21_X1   g16022(.A1(new_n16109_), .A2(new_n16169_), .B(new_n16168_), .ZN(new_n16279_));
  OAI21_X1   g16023(.A1(new_n16113_), .A2(new_n16149_), .B(new_n16151_), .ZN(new_n16280_));
  AOI21_X1   g16024(.A1(new_n16123_), .A2(new_n16147_), .B(new_n16121_), .ZN(new_n16281_));
  OAI21_X1   g16025(.A1(new_n16128_), .A2(new_n16143_), .B(new_n16145_), .ZN(new_n16282_));
  AOI22_X1   g16026(.A1(new_n11926_), .A2(\b[18] ), .B1(new_n11924_), .B2(\b[17] ), .ZN(new_n16283_));
  OAI21_X1   g16027(.A1(new_n1296_), .A2(new_n12317_), .B(new_n16283_), .ZN(new_n16284_));
  AOI21_X1   g16028(.A1(new_n2038_), .A2(new_n11929_), .B(new_n16284_), .ZN(new_n16285_));
  XOR2_X1    g16029(.A1(new_n16285_), .A2(new_n12312_), .Z(new_n16286_));
  NOR2_X1    g16030(.A1(new_n16136_), .A2(new_n16140_), .ZN(new_n16287_));
  NOR2_X1    g16031(.A1(new_n16287_), .A2(new_n16139_), .ZN(new_n16288_));
  AOI22_X1   g16032(.A1(new_n12922_), .A2(\b[15] ), .B1(\b[14] ), .B2(new_n12923_), .ZN(new_n16289_));
  XOR2_X1    g16033(.A1(new_n16289_), .A2(new_n1002_), .Z(new_n16290_));
  XOR2_X1    g16034(.A1(new_n16290_), .A2(new_n15911_), .Z(new_n16291_));
  NOR2_X1    g16035(.A1(new_n16288_), .A2(new_n16291_), .ZN(new_n16292_));
  INV_X1     g16036(.I(new_n16292_), .ZN(new_n16293_));
  NAND2_X1   g16037(.A1(new_n16288_), .A2(new_n16291_), .ZN(new_n16294_));
  NAND2_X1   g16038(.A1(new_n16293_), .A2(new_n16294_), .ZN(new_n16295_));
  XOR2_X1    g16039(.A1(new_n16295_), .A2(new_n16286_), .Z(new_n16296_));
  INV_X1     g16040(.I(new_n16296_), .ZN(new_n16297_));
  AOI22_X1   g16041(.A1(new_n10981_), .A2(\b[21] ), .B1(new_n10979_), .B2(\b[20] ), .ZN(new_n16298_));
  OAI21_X1   g16042(.A1(new_n1859_), .A2(new_n11306_), .B(new_n16298_), .ZN(new_n16299_));
  AOI21_X1   g16043(.A1(new_n2032_), .A2(new_n10984_), .B(new_n16299_), .ZN(new_n16300_));
  XOR2_X1    g16044(.A1(new_n16300_), .A2(new_n10989_), .Z(new_n16301_));
  NOR2_X1    g16045(.A1(new_n16297_), .A2(new_n16301_), .ZN(new_n16302_));
  NAND2_X1   g16046(.A1(new_n16297_), .A2(new_n16301_), .ZN(new_n16303_));
  INV_X1     g16047(.I(new_n16303_), .ZN(new_n16304_));
  NOR2_X1    g16048(.A1(new_n16304_), .A2(new_n16302_), .ZN(new_n16305_));
  XOR2_X1    g16049(.A1(new_n16305_), .A2(new_n16282_), .Z(new_n16306_));
  INV_X1     g16050(.I(new_n16306_), .ZN(new_n16307_));
  AOI22_X1   g16051(.A1(new_n10064_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n10062_), .ZN(new_n16308_));
  OAI21_X1   g16052(.A1(new_n2142_), .A2(new_n10399_), .B(new_n16308_), .ZN(new_n16309_));
  AOI21_X1   g16053(.A1(new_n3033_), .A2(new_n10068_), .B(new_n16309_), .ZN(new_n16310_));
  XOR2_X1    g16054(.A1(new_n16310_), .A2(new_n10057_), .Z(new_n16311_));
  NOR2_X1    g16055(.A1(new_n16307_), .A2(new_n16311_), .ZN(new_n16312_));
  NAND2_X1   g16056(.A1(new_n16307_), .A2(new_n16311_), .ZN(new_n16313_));
  INV_X1     g16057(.I(new_n16313_), .ZN(new_n16314_));
  NOR2_X1    g16058(.A1(new_n16314_), .A2(new_n16312_), .ZN(new_n16315_));
  XOR2_X1    g16059(.A1(new_n16315_), .A2(new_n16281_), .Z(new_n16316_));
  OAI22_X1   g16060(.A1(new_n10390_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n10389_), .ZN(new_n16317_));
  AOI21_X1   g16061(.A1(\b[25] ), .A2(new_n9471_), .B(new_n16317_), .ZN(new_n16318_));
  OAI21_X1   g16062(.A1(new_n3165_), .A2(new_n10388_), .B(new_n16318_), .ZN(new_n16319_));
  XOR2_X1    g16063(.A1(new_n16319_), .A2(\a[53] ), .Z(new_n16320_));
  NOR2_X1    g16064(.A1(new_n16316_), .A2(new_n16320_), .ZN(new_n16321_));
  NAND2_X1   g16065(.A1(new_n16316_), .A2(new_n16320_), .ZN(new_n16322_));
  INV_X1     g16066(.I(new_n16322_), .ZN(new_n16323_));
  NOR2_X1    g16067(.A1(new_n16323_), .A2(new_n16321_), .ZN(new_n16324_));
  XOR2_X1    g16068(.A1(new_n16324_), .A2(new_n16280_), .Z(new_n16325_));
  AOI22_X1   g16069(.A1(new_n8241_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n8246_), .ZN(new_n16326_));
  OAI21_X1   g16070(.A1(new_n3185_), .A2(new_n9114_), .B(new_n16326_), .ZN(new_n16327_));
  AOI21_X1   g16071(.A1(new_n4230_), .A2(new_n8252_), .B(new_n16327_), .ZN(new_n16328_));
  XOR2_X1    g16072(.A1(new_n16328_), .A2(new_n8248_), .Z(new_n16329_));
  INV_X1     g16073(.I(new_n16329_), .ZN(new_n16330_));
  NAND2_X1   g16074(.A1(new_n16153_), .A2(new_n16161_), .ZN(new_n16331_));
  NAND2_X1   g16075(.A1(new_n16331_), .A2(new_n16160_), .ZN(new_n16332_));
  NAND2_X1   g16076(.A1(new_n16332_), .A2(new_n16330_), .ZN(new_n16333_));
  NAND3_X1   g16077(.A1(new_n16331_), .A2(new_n16160_), .A3(new_n16329_), .ZN(new_n16334_));
  NAND2_X1   g16078(.A1(new_n16333_), .A2(new_n16334_), .ZN(new_n16335_));
  XNOR2_X1   g16079(.A1(new_n16325_), .A2(new_n16335_), .ZN(new_n16336_));
  INV_X1     g16080(.I(new_n16336_), .ZN(new_n16337_));
  AOI22_X1   g16081(.A1(new_n7403_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n7408_), .ZN(new_n16338_));
  OAI21_X1   g16082(.A1(new_n4022_), .A2(new_n9488_), .B(new_n16338_), .ZN(new_n16339_));
  AOI21_X1   g16083(.A1(new_n4223_), .A2(new_n7414_), .B(new_n16339_), .ZN(new_n16340_));
  XOR2_X1    g16084(.A1(new_n16340_), .A2(new_n7410_), .Z(new_n16341_));
  NOR2_X1    g16085(.A1(new_n16337_), .A2(new_n16341_), .ZN(new_n16342_));
  INV_X1     g16086(.I(new_n16342_), .ZN(new_n16343_));
  NAND2_X1   g16087(.A1(new_n16337_), .A2(new_n16341_), .ZN(new_n16344_));
  NAND2_X1   g16088(.A1(new_n16343_), .A2(new_n16344_), .ZN(new_n16345_));
  XOR2_X1    g16089(.A1(new_n16345_), .A2(new_n16279_), .Z(new_n16346_));
  NOR2_X1    g16090(.A1(new_n16346_), .A2(new_n16278_), .ZN(new_n16347_));
  NAND2_X1   g16091(.A1(new_n16346_), .A2(new_n16278_), .ZN(new_n16348_));
  INV_X1     g16092(.I(new_n16348_), .ZN(new_n16349_));
  NOR2_X1    g16093(.A1(new_n16349_), .A2(new_n16347_), .ZN(new_n16350_));
  XOR2_X1    g16094(.A1(new_n16350_), .A2(new_n16274_), .Z(new_n16351_));
  INV_X1     g16095(.I(new_n16351_), .ZN(new_n16352_));
  AOI22_X1   g16096(.A1(new_n6108_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n6111_), .ZN(new_n16353_));
  OAI21_X1   g16097(.A1(new_n5312_), .A2(new_n7708_), .B(new_n16353_), .ZN(new_n16354_));
  AOI21_X1   g16098(.A1(new_n6310_), .A2(new_n6105_), .B(new_n16354_), .ZN(new_n16355_));
  XOR2_X1    g16099(.A1(new_n16355_), .A2(new_n5849_), .Z(new_n16356_));
  NOR2_X1    g16100(.A1(new_n16352_), .A2(new_n16356_), .ZN(new_n16357_));
  NAND2_X1   g16101(.A1(new_n16352_), .A2(new_n16356_), .ZN(new_n16358_));
  INV_X1     g16102(.I(new_n16358_), .ZN(new_n16359_));
  NOR2_X1    g16103(.A1(new_n16359_), .A2(new_n16357_), .ZN(new_n16360_));
  XOR2_X1    g16104(.A1(new_n16360_), .A2(new_n16272_), .Z(new_n16361_));
  AOI22_X1   g16105(.A1(new_n5155_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n5160_), .ZN(new_n16362_));
  OAI21_X1   g16106(.A1(new_n6284_), .A2(new_n6877_), .B(new_n16362_), .ZN(new_n16363_));
  AOI21_X1   g16107(.A1(new_n7106_), .A2(new_n5166_), .B(new_n16363_), .ZN(new_n16364_));
  XOR2_X1    g16108(.A1(new_n16364_), .A2(new_n5162_), .Z(new_n16365_));
  NOR2_X1    g16109(.A1(new_n16361_), .A2(new_n16365_), .ZN(new_n16366_));
  NAND2_X1   g16110(.A1(new_n16361_), .A2(new_n16365_), .ZN(new_n16367_));
  INV_X1     g16111(.I(new_n16367_), .ZN(new_n16368_));
  NOR2_X1    g16112(.A1(new_n16368_), .A2(new_n16366_), .ZN(new_n16369_));
  XOR2_X1    g16113(.A1(new_n16369_), .A2(new_n16270_), .Z(new_n16370_));
  AOI22_X1   g16114(.A1(new_n4918_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n4921_), .ZN(new_n16371_));
  OAI21_X1   g16115(.A1(new_n6775_), .A2(new_n6099_), .B(new_n16371_), .ZN(new_n16372_));
  AOI21_X1   g16116(.A1(new_n7926_), .A2(new_n4699_), .B(new_n16372_), .ZN(new_n16373_));
  XOR2_X1    g16117(.A1(new_n16373_), .A2(new_n4446_), .Z(new_n16374_));
  INV_X1     g16118(.I(new_n16374_), .ZN(new_n16375_));
  AND2_X2    g16119(.A1(new_n16370_), .A2(new_n16375_), .Z(new_n16376_));
  NOR2_X1    g16120(.A1(new_n16370_), .A2(new_n16375_), .ZN(new_n16377_));
  NOR2_X1    g16121(.A1(new_n16376_), .A2(new_n16377_), .ZN(new_n16378_));
  XNOR2_X1   g16122(.A1(new_n16378_), .A2(new_n16268_), .ZN(new_n16379_));
  NAND2_X1   g16123(.A1(new_n16204_), .A2(new_n16087_), .ZN(new_n16380_));
  NAND2_X1   g16124(.A1(new_n16380_), .A2(new_n16203_), .ZN(new_n16381_));
  AOI22_X1   g16125(.A1(new_n3864_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n3869_), .ZN(new_n16382_));
  OAI21_X1   g16126(.A1(new_n7617_), .A2(new_n5410_), .B(new_n16382_), .ZN(new_n16383_));
  AOI21_X1   g16127(.A1(new_n8792_), .A2(new_n3872_), .B(new_n16383_), .ZN(new_n16384_));
  XOR2_X1    g16128(.A1(new_n16384_), .A2(new_n3876_), .Z(new_n16385_));
  INV_X1     g16129(.I(new_n16385_), .ZN(new_n16386_));
  NAND2_X1   g16130(.A1(new_n16381_), .A2(new_n16386_), .ZN(new_n16387_));
  NAND3_X1   g16131(.A1(new_n16380_), .A2(new_n16203_), .A3(new_n16385_), .ZN(new_n16388_));
  NAND2_X1   g16132(.A1(new_n16387_), .A2(new_n16388_), .ZN(new_n16389_));
  XOR2_X1    g16133(.A1(new_n16379_), .A2(new_n16389_), .Z(new_n16390_));
  OR2_X2     g16134(.A1(new_n16390_), .A2(new_n16266_), .Z(new_n16391_));
  NAND2_X1   g16135(.A1(new_n16390_), .A2(new_n16266_), .ZN(new_n16392_));
  NAND2_X1   g16136(.A1(new_n16391_), .A2(new_n16392_), .ZN(new_n16393_));
  XNOR2_X1   g16137(.A1(new_n16393_), .A2(new_n16262_), .ZN(new_n16394_));
  NAND2_X1   g16138(.A1(new_n16394_), .A2(new_n16256_), .ZN(new_n16395_));
  OR2_X2     g16139(.A1(new_n16394_), .A2(new_n16256_), .Z(new_n16396_));
  NAND2_X1   g16140(.A1(new_n16396_), .A2(new_n16395_), .ZN(new_n16397_));
  XOR2_X1    g16141(.A1(new_n16397_), .A2(new_n16251_), .Z(new_n16398_));
  AOI22_X1   g16142(.A1(new_n2202_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n2205_), .ZN(new_n16399_));
  OAI21_X1   g16143(.A1(new_n9972_), .A2(new_n2370_), .B(new_n16399_), .ZN(new_n16400_));
  AOI21_X1   g16144(.A1(new_n10631_), .A2(new_n2208_), .B(new_n16400_), .ZN(new_n16401_));
  XOR2_X1    g16145(.A1(new_n16401_), .A2(\a[23] ), .Z(new_n16402_));
  NAND2_X1   g16146(.A1(new_n16398_), .A2(new_n16402_), .ZN(new_n16403_));
  OR2_X2     g16147(.A1(new_n16398_), .A2(new_n16402_), .Z(new_n16404_));
  NAND2_X1   g16148(.A1(new_n16404_), .A2(new_n16403_), .ZN(new_n16405_));
  XNOR2_X1   g16149(.A1(new_n16405_), .A2(new_n16248_), .ZN(new_n16406_));
  AOI22_X1   g16150(.A1(new_n1738_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n1743_), .ZN(new_n16407_));
  OAI21_X1   g16151(.A1(new_n11195_), .A2(new_n1931_), .B(new_n16407_), .ZN(new_n16408_));
  AOI21_X1   g16152(.A1(new_n11836_), .A2(new_n1746_), .B(new_n16408_), .ZN(new_n16409_));
  XOR2_X1    g16153(.A1(new_n16409_), .A2(new_n1736_), .Z(new_n16410_));
  INV_X1     g16154(.I(new_n16410_), .ZN(new_n16411_));
  NAND2_X1   g16155(.A1(new_n16406_), .A2(new_n16411_), .ZN(new_n16412_));
  OR2_X2     g16156(.A1(new_n16406_), .A2(new_n16411_), .Z(new_n16413_));
  NAND2_X1   g16157(.A1(new_n16413_), .A2(new_n16412_), .ZN(new_n16414_));
  XOR2_X1    g16158(.A1(new_n16414_), .A2(new_n16244_), .Z(new_n16415_));
  OAI22_X1   g16159(.A1(new_n1592_), .A2(new_n12800_), .B1(new_n12796_), .B2(new_n1505_), .ZN(new_n16416_));
  AOI21_X1   g16160(.A1(\b[61] ), .A2(new_n1584_), .B(new_n16416_), .ZN(new_n16417_));
  OAI21_X1   g16161(.A1(new_n15183_), .A2(new_n1732_), .B(new_n16417_), .ZN(new_n16418_));
  XOR2_X1    g16162(.A1(new_n16418_), .A2(\a[17] ), .Z(new_n16419_));
  NOR2_X1    g16163(.A1(new_n16415_), .A2(new_n16419_), .ZN(new_n16420_));
  AND2_X2    g16164(.A1(new_n16415_), .A2(new_n16419_), .Z(new_n16421_));
  NOR2_X1    g16165(.A1(new_n16421_), .A2(new_n16420_), .ZN(new_n16422_));
  XOR2_X1    g16166(.A1(new_n16422_), .A2(new_n16241_), .Z(new_n16423_));
  NAND2_X1   g16167(.A1(new_n16423_), .A2(new_n16239_), .ZN(new_n16424_));
  INV_X1     g16168(.I(new_n16424_), .ZN(new_n16425_));
  NOR2_X1    g16169(.A1(new_n16423_), .A2(new_n16239_), .ZN(new_n16426_));
  NOR2_X1    g16170(.A1(new_n16425_), .A2(new_n16426_), .ZN(new_n16427_));
  XOR2_X1    g16171(.A1(new_n16236_), .A2(new_n16427_), .Z(\f[78] ));
  NOR2_X1    g16172(.A1(new_n16421_), .A2(new_n16241_), .ZN(new_n16429_));
  NOR2_X1    g16173(.A1(new_n16429_), .A2(new_n16420_), .ZN(new_n16430_));
  INV_X1     g16174(.I(new_n16430_), .ZN(new_n16431_));
  NAND2_X1   g16175(.A1(new_n16413_), .A2(new_n16244_), .ZN(new_n16432_));
  AND2_X2    g16176(.A1(new_n16432_), .A2(new_n16412_), .Z(new_n16433_));
  INV_X1     g16177(.I(new_n16433_), .ZN(new_n16434_));
  NAND2_X1   g16178(.A1(new_n16404_), .A2(new_n16248_), .ZN(new_n16435_));
  AND2_X2    g16179(.A1(new_n16435_), .A2(new_n16403_), .Z(new_n16436_));
  OAI22_X1   g16180(.A1(new_n1751_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n1754_), .ZN(new_n16437_));
  AOI21_X1   g16181(.A1(\b[59] ), .A2(new_n1939_), .B(new_n16437_), .ZN(new_n16438_));
  OAI21_X1   g16182(.A1(new_n13110_), .A2(new_n1757_), .B(new_n16438_), .ZN(new_n16439_));
  XOR2_X1    g16183(.A1(new_n16439_), .A2(\a[20] ), .Z(new_n16440_));
  AOI22_X1   g16184(.A1(new_n2202_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n2205_), .ZN(new_n16441_));
  OAI21_X1   g16185(.A1(new_n10308_), .A2(new_n2370_), .B(new_n16441_), .ZN(new_n16442_));
  AOI21_X1   g16186(.A1(new_n12164_), .A2(new_n2208_), .B(new_n16442_), .ZN(new_n16443_));
  XOR2_X1    g16187(.A1(new_n16443_), .A2(new_n2200_), .Z(new_n16444_));
  INV_X1     g16188(.I(new_n16444_), .ZN(new_n16445_));
  INV_X1     g16189(.I(new_n16251_), .ZN(new_n16446_));
  INV_X1     g16190(.I(new_n16395_), .ZN(new_n16447_));
  AOI21_X1   g16191(.A1(new_n16446_), .A2(new_n16396_), .B(new_n16447_), .ZN(new_n16448_));
  INV_X1     g16192(.I(new_n16448_), .ZN(new_n16449_));
  AOI22_X1   g16193(.A1(new_n2716_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n2719_), .ZN(new_n16450_));
  OAI21_X1   g16194(.A1(new_n9376_), .A2(new_n2924_), .B(new_n16450_), .ZN(new_n16451_));
  AOI21_X1   g16195(.A1(new_n9979_), .A2(new_n2722_), .B(new_n16451_), .ZN(new_n16452_));
  XOR2_X1    g16196(.A1(new_n16452_), .A2(new_n2714_), .Z(new_n16453_));
  INV_X1     g16197(.I(new_n16453_), .ZN(new_n16454_));
  INV_X1     g16198(.I(new_n16392_), .ZN(new_n16455_));
  AOI21_X1   g16199(.A1(new_n16262_), .A2(new_n16391_), .B(new_n16455_), .ZN(new_n16456_));
  AOI22_X1   g16200(.A1(new_n3267_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n3270_), .ZN(new_n16457_));
  OAI21_X1   g16201(.A1(new_n8500_), .A2(new_n3475_), .B(new_n16457_), .ZN(new_n16458_));
  AOI21_X1   g16202(.A1(new_n9987_), .A2(new_n3273_), .B(new_n16458_), .ZN(new_n16459_));
  XOR2_X1    g16203(.A1(new_n16459_), .A2(new_n3264_), .Z(new_n16460_));
  INV_X1     g16204(.I(new_n16379_), .ZN(new_n16461_));
  INV_X1     g16205(.I(new_n16387_), .ZN(new_n16462_));
  AOI21_X1   g16206(.A1(new_n16461_), .A2(new_n16388_), .B(new_n16462_), .ZN(new_n16463_));
  OAI22_X1   g16207(.A1(new_n8127_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n8168_), .ZN(new_n16464_));
  AOI21_X1   g16208(.A1(\b[47] ), .A2(new_n4053_), .B(new_n16464_), .ZN(new_n16465_));
  OAI21_X1   g16209(.A1(new_n9050_), .A2(new_n4727_), .B(new_n16465_), .ZN(new_n16466_));
  XOR2_X1    g16210(.A1(new_n16466_), .A2(new_n3876_), .Z(new_n16467_));
  INV_X1     g16211(.I(new_n16377_), .ZN(new_n16468_));
  AOI21_X1   g16212(.A1(new_n16268_), .A2(new_n16468_), .B(new_n16376_), .ZN(new_n16469_));
  AOI22_X1   g16213(.A1(new_n4918_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n4921_), .ZN(new_n16470_));
  OAI21_X1   g16214(.A1(new_n7074_), .A2(new_n6099_), .B(new_n16470_), .ZN(new_n16471_));
  AOI21_X1   g16215(.A1(new_n9337_), .A2(new_n4699_), .B(new_n16471_), .ZN(new_n16472_));
  XOR2_X1    g16216(.A1(new_n16472_), .A2(new_n4446_), .Z(new_n16473_));
  INV_X1     g16217(.I(new_n16473_), .ZN(new_n16474_));
  NOR2_X1    g16218(.A1(new_n16359_), .A2(new_n16272_), .ZN(new_n16475_));
  NOR2_X1    g16219(.A1(new_n16475_), .A2(new_n16357_), .ZN(new_n16476_));
  AOI22_X1   g16220(.A1(new_n6108_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n6111_), .ZN(new_n16477_));
  OAI21_X1   g16221(.A1(new_n5341_), .A2(new_n7708_), .B(new_n16477_), .ZN(new_n16478_));
  AOI21_X1   g16222(.A1(new_n5793_), .A2(new_n6105_), .B(new_n16478_), .ZN(new_n16479_));
  XOR2_X1    g16223(.A1(new_n16479_), .A2(new_n5849_), .Z(new_n16480_));
  AOI21_X1   g16224(.A1(new_n16274_), .A2(new_n16348_), .B(new_n16347_), .ZN(new_n16481_));
  INV_X1     g16225(.I(new_n16481_), .ZN(new_n16482_));
  OAI22_X1   g16226(.A1(new_n7730_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n7731_), .ZN(new_n16483_));
  AOI21_X1   g16227(.A1(\b[35] ), .A2(new_n6887_), .B(new_n16483_), .ZN(new_n16484_));
  OAI21_X1   g16228(.A1(new_n5322_), .A2(new_n7728_), .B(new_n16484_), .ZN(new_n16485_));
  XOR2_X1    g16229(.A1(new_n16485_), .A2(\a[44] ), .Z(new_n16486_));
  AOI21_X1   g16230(.A1(new_n16279_), .A2(new_n16344_), .B(new_n16342_), .ZN(new_n16487_));
  AOI22_X1   g16231(.A1(new_n7403_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n7408_), .ZN(new_n16488_));
  OAI21_X1   g16232(.A1(new_n4023_), .A2(new_n9488_), .B(new_n16488_), .ZN(new_n16489_));
  AOI21_X1   g16233(.A1(new_n5103_), .A2(new_n7414_), .B(new_n16489_), .ZN(new_n16490_));
  XOR2_X1    g16234(.A1(new_n16490_), .A2(new_n7410_), .Z(new_n16491_));
  INV_X1     g16235(.I(new_n16491_), .ZN(new_n16492_));
  AOI22_X1   g16236(.A1(new_n9125_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n9123_), .ZN(new_n16493_));
  OAI21_X1   g16237(.A1(new_n3006_), .A2(new_n9470_), .B(new_n16493_), .ZN(new_n16494_));
  AOI21_X1   g16238(.A1(new_n3807_), .A2(new_n9129_), .B(new_n16494_), .ZN(new_n16495_));
  XOR2_X1    g16239(.A1(new_n16495_), .A2(new_n9133_), .Z(new_n16496_));
  NOR2_X1    g16240(.A1(new_n16314_), .A2(new_n16281_), .ZN(new_n16497_));
  NOR2_X1    g16241(.A1(new_n16497_), .A2(new_n16312_), .ZN(new_n16498_));
  AOI22_X1   g16242(.A1(new_n10981_), .A2(\b[22] ), .B1(new_n10979_), .B2(\b[21] ), .ZN(new_n16499_));
  OAI21_X1   g16243(.A1(new_n1860_), .A2(new_n11306_), .B(new_n16499_), .ZN(new_n16500_));
  AOI21_X1   g16244(.A1(new_n2659_), .A2(new_n10984_), .B(new_n16500_), .ZN(new_n16501_));
  XOR2_X1    g16245(.A1(new_n16501_), .A2(new_n10989_), .Z(new_n16502_));
  INV_X1     g16246(.I(new_n16286_), .ZN(new_n16503_));
  AOI21_X1   g16247(.A1(new_n16503_), .A2(new_n16294_), .B(new_n16292_), .ZN(new_n16504_));
  INV_X1     g16248(.I(new_n16504_), .ZN(new_n16505_));
  AOI22_X1   g16249(.A1(new_n11926_), .A2(\b[19] ), .B1(new_n11924_), .B2(\b[18] ), .ZN(new_n16506_));
  OAI21_X1   g16250(.A1(new_n1432_), .A2(new_n12317_), .B(new_n16506_), .ZN(new_n16507_));
  AOI21_X1   g16251(.A1(new_n1695_), .A2(new_n11929_), .B(new_n16507_), .ZN(new_n16508_));
  XOR2_X1    g16252(.A1(new_n16508_), .A2(\a[62] ), .Z(new_n16509_));
  NOR2_X1    g16253(.A1(new_n16289_), .A2(\a[14] ), .ZN(new_n16510_));
  NOR2_X1    g16254(.A1(new_n16510_), .A2(new_n15912_), .ZN(new_n16511_));
  AOI21_X1   g16255(.A1(\a[14] ), .A2(new_n16289_), .B(new_n16511_), .ZN(new_n16512_));
  AOI22_X1   g16256(.A1(new_n12922_), .A2(\b[16] ), .B1(\b[15] ), .B2(new_n12923_), .ZN(new_n16513_));
  NAND2_X1   g16257(.A1(new_n16512_), .A2(new_n16513_), .ZN(new_n16514_));
  NOR2_X1    g16258(.A1(new_n16512_), .A2(new_n16513_), .ZN(new_n16515_));
  INV_X1     g16259(.I(new_n16515_), .ZN(new_n16516_));
  NAND2_X1   g16260(.A1(new_n16516_), .A2(new_n16514_), .ZN(new_n16517_));
  XNOR2_X1   g16261(.A1(new_n16509_), .A2(new_n16517_), .ZN(new_n16518_));
  NOR2_X1    g16262(.A1(new_n16505_), .A2(new_n16518_), .ZN(new_n16519_));
  NAND2_X1   g16263(.A1(new_n16505_), .A2(new_n16518_), .ZN(new_n16520_));
  INV_X1     g16264(.I(new_n16520_), .ZN(new_n16521_));
  NOR2_X1    g16265(.A1(new_n16521_), .A2(new_n16519_), .ZN(new_n16522_));
  XOR2_X1    g16266(.A1(new_n16522_), .A2(new_n16502_), .Z(new_n16523_));
  INV_X1     g16267(.I(new_n16523_), .ZN(new_n16524_));
  AOI21_X1   g16268(.A1(new_n16282_), .A2(new_n16303_), .B(new_n16302_), .ZN(new_n16525_));
  OAI22_X1   g16269(.A1(new_n11298_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n11297_), .ZN(new_n16526_));
  AOI21_X1   g16270(.A1(\b[23] ), .A2(new_n11296_), .B(new_n16526_), .ZN(new_n16527_));
  OAI21_X1   g16271(.A1(new_n2655_), .A2(new_n10069_), .B(new_n16527_), .ZN(new_n16528_));
  XOR2_X1    g16272(.A1(new_n16528_), .A2(\a[56] ), .Z(new_n16529_));
  NOR2_X1    g16273(.A1(new_n16529_), .A2(new_n16525_), .ZN(new_n16530_));
  INV_X1     g16274(.I(new_n16530_), .ZN(new_n16531_));
  NAND2_X1   g16275(.A1(new_n16529_), .A2(new_n16525_), .ZN(new_n16532_));
  NAND2_X1   g16276(.A1(new_n16531_), .A2(new_n16532_), .ZN(new_n16533_));
  XOR2_X1    g16277(.A1(new_n16533_), .A2(new_n16524_), .Z(new_n16534_));
  NOR2_X1    g16278(.A1(new_n16498_), .A2(new_n16534_), .ZN(new_n16535_));
  INV_X1     g16279(.I(new_n16535_), .ZN(new_n16536_));
  NAND2_X1   g16280(.A1(new_n16498_), .A2(new_n16534_), .ZN(new_n16537_));
  NAND2_X1   g16281(.A1(new_n16536_), .A2(new_n16537_), .ZN(new_n16538_));
  XOR2_X1    g16282(.A1(new_n16538_), .A2(new_n16496_), .Z(new_n16539_));
  AOI21_X1   g16283(.A1(new_n16280_), .A2(new_n16322_), .B(new_n16321_), .ZN(new_n16540_));
  AOI22_X1   g16284(.A1(new_n8241_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n8246_), .ZN(new_n16541_));
  OAI21_X1   g16285(.A1(new_n3592_), .A2(new_n9114_), .B(new_n16541_), .ZN(new_n16542_));
  AOI21_X1   g16286(.A1(new_n3796_), .A2(new_n8252_), .B(new_n16542_), .ZN(new_n16543_));
  XOR2_X1    g16287(.A1(new_n16543_), .A2(new_n8248_), .Z(new_n16544_));
  NOR2_X1    g16288(.A1(new_n16540_), .A2(new_n16544_), .ZN(new_n16545_));
  INV_X1     g16289(.I(new_n16545_), .ZN(new_n16546_));
  NAND2_X1   g16290(.A1(new_n16540_), .A2(new_n16544_), .ZN(new_n16547_));
  NAND2_X1   g16291(.A1(new_n16546_), .A2(new_n16547_), .ZN(new_n16548_));
  XOR2_X1    g16292(.A1(new_n16548_), .A2(new_n16539_), .Z(new_n16549_));
  NAND2_X1   g16293(.A1(new_n16325_), .A2(new_n16334_), .ZN(new_n16550_));
  NAND2_X1   g16294(.A1(new_n16550_), .A2(new_n16333_), .ZN(new_n16551_));
  INV_X1     g16295(.I(new_n16551_), .ZN(new_n16552_));
  NOR2_X1    g16296(.A1(new_n16552_), .A2(new_n16549_), .ZN(new_n16553_));
  INV_X1     g16297(.I(new_n16553_), .ZN(new_n16554_));
  NAND2_X1   g16298(.A1(new_n16552_), .A2(new_n16549_), .ZN(new_n16555_));
  NAND2_X1   g16299(.A1(new_n16554_), .A2(new_n16555_), .ZN(new_n16556_));
  XOR2_X1    g16300(.A1(new_n16556_), .A2(new_n16492_), .Z(new_n16557_));
  NAND2_X1   g16301(.A1(new_n16557_), .A2(new_n16487_), .ZN(new_n16558_));
  NOR2_X1    g16302(.A1(new_n16557_), .A2(new_n16487_), .ZN(new_n16559_));
  INV_X1     g16303(.I(new_n16559_), .ZN(new_n16560_));
  NAND2_X1   g16304(.A1(new_n16560_), .A2(new_n16558_), .ZN(new_n16561_));
  XOR2_X1    g16305(.A1(new_n16561_), .A2(new_n16486_), .Z(new_n16562_));
  NOR2_X1    g16306(.A1(new_n16562_), .A2(new_n16482_), .ZN(new_n16563_));
  INV_X1     g16307(.I(new_n16563_), .ZN(new_n16564_));
  NAND2_X1   g16308(.A1(new_n16562_), .A2(new_n16482_), .ZN(new_n16565_));
  NAND2_X1   g16309(.A1(new_n16564_), .A2(new_n16565_), .ZN(new_n16566_));
  XOR2_X1    g16310(.A1(new_n16566_), .A2(new_n16480_), .Z(new_n16567_));
  INV_X1     g16311(.I(new_n16567_), .ZN(new_n16568_));
  OAI22_X1   g16312(.A1(new_n6775_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n6490_), .ZN(new_n16569_));
  AOI21_X1   g16313(.A1(\b[41] ), .A2(new_n5420_), .B(new_n16569_), .ZN(new_n16570_));
  OAI21_X1   g16314(.A1(new_n6785_), .A2(new_n6124_), .B(new_n16570_), .ZN(new_n16571_));
  XOR2_X1    g16315(.A1(new_n16571_), .A2(\a[38] ), .Z(new_n16572_));
  NOR2_X1    g16316(.A1(new_n16568_), .A2(new_n16572_), .ZN(new_n16573_));
  NAND2_X1   g16317(.A1(new_n16568_), .A2(new_n16572_), .ZN(new_n16574_));
  INV_X1     g16318(.I(new_n16574_), .ZN(new_n16575_));
  NOR2_X1    g16319(.A1(new_n16575_), .A2(new_n16573_), .ZN(new_n16576_));
  XOR2_X1    g16320(.A1(new_n16576_), .A2(new_n16476_), .Z(new_n16577_));
  AOI21_X1   g16321(.A1(new_n16270_), .A2(new_n16367_), .B(new_n16366_), .ZN(new_n16578_));
  NOR2_X1    g16322(.A1(new_n16577_), .A2(new_n16578_), .ZN(new_n16579_));
  INV_X1     g16323(.I(new_n16579_), .ZN(new_n16580_));
  NAND2_X1   g16324(.A1(new_n16577_), .A2(new_n16578_), .ZN(new_n16581_));
  NAND2_X1   g16325(.A1(new_n16580_), .A2(new_n16581_), .ZN(new_n16582_));
  XOR2_X1    g16326(.A1(new_n16582_), .A2(new_n16474_), .Z(new_n16583_));
  NOR2_X1    g16327(.A1(new_n16583_), .A2(new_n16469_), .ZN(new_n16584_));
  INV_X1     g16328(.I(new_n16584_), .ZN(new_n16585_));
  NAND2_X1   g16329(.A1(new_n16583_), .A2(new_n16469_), .ZN(new_n16586_));
  NAND2_X1   g16330(.A1(new_n16585_), .A2(new_n16586_), .ZN(new_n16587_));
  XNOR2_X1   g16331(.A1(new_n16587_), .A2(new_n16467_), .ZN(new_n16588_));
  INV_X1     g16332(.I(new_n16588_), .ZN(new_n16589_));
  NOR2_X1    g16333(.A1(new_n16589_), .A2(new_n16463_), .ZN(new_n16590_));
  INV_X1     g16334(.I(new_n16590_), .ZN(new_n16591_));
  NAND2_X1   g16335(.A1(new_n16589_), .A2(new_n16463_), .ZN(new_n16592_));
  NAND2_X1   g16336(.A1(new_n16591_), .A2(new_n16592_), .ZN(new_n16593_));
  XOR2_X1    g16337(.A1(new_n16593_), .A2(new_n16460_), .Z(new_n16594_));
  INV_X1     g16338(.I(new_n16594_), .ZN(new_n16595_));
  NOR2_X1    g16339(.A1(new_n16595_), .A2(new_n16456_), .ZN(new_n16596_));
  NAND2_X1   g16340(.A1(new_n16595_), .A2(new_n16456_), .ZN(new_n16597_));
  INV_X1     g16341(.I(new_n16597_), .ZN(new_n16598_));
  NOR2_X1    g16342(.A1(new_n16598_), .A2(new_n16596_), .ZN(new_n16599_));
  XOR2_X1    g16343(.A1(new_n16599_), .A2(new_n16454_), .Z(new_n16600_));
  NAND2_X1   g16344(.A1(new_n16600_), .A2(new_n16449_), .ZN(new_n16601_));
  OR2_X2     g16345(.A1(new_n16600_), .A2(new_n16449_), .Z(new_n16602_));
  NAND2_X1   g16346(.A1(new_n16602_), .A2(new_n16601_), .ZN(new_n16603_));
  XOR2_X1    g16347(.A1(new_n16603_), .A2(new_n16445_), .Z(new_n16604_));
  OR2_X2     g16348(.A1(new_n16604_), .A2(new_n16440_), .Z(new_n16605_));
  NAND2_X1   g16349(.A1(new_n16604_), .A2(new_n16440_), .ZN(new_n16606_));
  NAND2_X1   g16350(.A1(new_n16605_), .A2(new_n16606_), .ZN(new_n16607_));
  XOR2_X1    g16351(.A1(new_n16607_), .A2(new_n16436_), .Z(new_n16608_));
  AOI22_X1   g16352(.A1(new_n1584_), .A2(\b[62] ), .B1(\b[63] ), .B2(new_n1495_), .ZN(new_n16609_));
  OAI21_X1   g16353(.A1(new_n13107_), .A2(new_n1732_), .B(new_n16609_), .ZN(new_n16610_));
  XOR2_X1    g16354(.A1(new_n16610_), .A2(\a[17] ), .Z(new_n16611_));
  INV_X1     g16355(.I(new_n16611_), .ZN(new_n16612_));
  NAND2_X1   g16356(.A1(new_n16608_), .A2(new_n16612_), .ZN(new_n16613_));
  OR2_X2     g16357(.A1(new_n16608_), .A2(new_n16612_), .Z(new_n16614_));
  NAND2_X1   g16358(.A1(new_n16614_), .A2(new_n16613_), .ZN(new_n16615_));
  XOR2_X1    g16359(.A1(new_n16615_), .A2(new_n16434_), .Z(new_n16616_));
  INV_X1     g16360(.I(new_n16427_), .ZN(new_n16617_));
  NOR3_X1    g16361(.A1(new_n16235_), .A2(new_n16234_), .A3(new_n16617_), .ZN(new_n16618_));
  OAI21_X1   g16362(.A1(new_n16618_), .A2(new_n16425_), .B(new_n16616_), .ZN(new_n16619_));
  INV_X1     g16363(.I(new_n16616_), .ZN(new_n16620_));
  AOI21_X1   g16364(.A1(new_n16033_), .A2(new_n16032_), .B(new_n15842_), .ZN(new_n16621_));
  OAI21_X1   g16365(.A1(new_n16621_), .A2(new_n16034_), .B(new_n16230_), .ZN(new_n16622_));
  NAND3_X1   g16366(.A1(new_n16622_), .A2(new_n16231_), .A3(new_n16427_), .ZN(new_n16623_));
  NAND3_X1   g16367(.A1(new_n16623_), .A2(new_n16424_), .A3(new_n16620_), .ZN(new_n16624_));
  NAND2_X1   g16368(.A1(new_n16619_), .A2(new_n16624_), .ZN(new_n16625_));
  XOR2_X1    g16369(.A1(new_n16625_), .A2(new_n16431_), .Z(\f[79] ));
  AOI21_X1   g16370(.A1(new_n16623_), .A2(new_n16424_), .B(new_n16620_), .ZN(new_n16627_));
  OAI21_X1   g16371(.A1(new_n16430_), .A2(new_n16627_), .B(new_n16624_), .ZN(new_n16628_));
  INV_X1     g16372(.I(new_n16613_), .ZN(new_n16629_));
  AOI21_X1   g16373(.A1(new_n16434_), .A2(new_n16614_), .B(new_n16629_), .ZN(new_n16630_));
  OAI22_X1   g16374(.A1(new_n13462_), .A2(new_n1732_), .B1(new_n12800_), .B2(new_n1917_), .ZN(new_n16631_));
  XOR2_X1    g16375(.A1(new_n16631_), .A2(\a[17] ), .Z(new_n16632_));
  INV_X1     g16376(.I(new_n16436_), .ZN(new_n16633_));
  INV_X1     g16377(.I(new_n16605_), .ZN(new_n16634_));
  AOI21_X1   g16378(.A1(new_n16633_), .A2(new_n16606_), .B(new_n16634_), .ZN(new_n16635_));
  AOI22_X1   g16379(.A1(new_n1738_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n1743_), .ZN(new_n16636_));
  OAI21_X1   g16380(.A1(new_n12147_), .A2(new_n1931_), .B(new_n16636_), .ZN(new_n16637_));
  AOI21_X1   g16381(.A1(new_n13444_), .A2(new_n1746_), .B(new_n16637_), .ZN(new_n16638_));
  XOR2_X1    g16382(.A1(new_n16638_), .A2(new_n1736_), .Z(new_n16639_));
  INV_X1     g16383(.I(new_n16639_), .ZN(new_n16640_));
  INV_X1     g16384(.I(new_n16601_), .ZN(new_n16641_));
  AOI21_X1   g16385(.A1(new_n16445_), .A2(new_n16602_), .B(new_n16641_), .ZN(new_n16642_));
  OAI22_X1   g16386(.A1(new_n2189_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n2194_), .ZN(new_n16643_));
  AOI21_X1   g16387(.A1(\b[57] ), .A2(new_n2361_), .B(new_n16643_), .ZN(new_n16644_));
  OAI21_X1   g16388(.A1(new_n12203_), .A2(new_n2197_), .B(new_n16644_), .ZN(new_n16645_));
  XOR2_X1    g16389(.A1(new_n16645_), .A2(\a[23] ), .Z(new_n16646_));
  INV_X1     g16390(.I(new_n16646_), .ZN(new_n16647_));
  AOI21_X1   g16391(.A1(new_n16454_), .A2(new_n16597_), .B(new_n16596_), .ZN(new_n16648_));
  AOI22_X1   g16392(.A1(new_n2716_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n2719_), .ZN(new_n16649_));
  OAI21_X1   g16393(.A1(new_n9942_), .A2(new_n2924_), .B(new_n16649_), .ZN(new_n16650_));
  AOI21_X1   g16394(.A1(new_n10318_), .A2(new_n2722_), .B(new_n16650_), .ZN(new_n16651_));
  XOR2_X1    g16395(.A1(new_n16651_), .A2(new_n2714_), .Z(new_n16652_));
  INV_X1     g16396(.I(new_n16460_), .ZN(new_n16653_));
  AOI21_X1   g16397(.A1(new_n16653_), .A2(new_n16592_), .B(new_n16590_), .ZN(new_n16654_));
  OAI22_X1   g16398(.A1(new_n9376_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n9032_), .ZN(new_n16655_));
  AOI21_X1   g16399(.A1(\b[51] ), .A2(new_n3456_), .B(new_n16655_), .ZN(new_n16656_));
  OAI21_X1   g16400(.A1(new_n9385_), .A2(new_n3261_), .B(new_n16656_), .ZN(new_n16657_));
  XOR2_X1    g16401(.A1(new_n16657_), .A2(new_n3264_), .Z(new_n16658_));
  AOI22_X1   g16402(.A1(new_n3864_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n3869_), .ZN(new_n16659_));
  OAI21_X1   g16403(.A1(new_n8127_), .A2(new_n5410_), .B(new_n16659_), .ZN(new_n16660_));
  AOI21_X1   g16404(.A1(new_n9684_), .A2(new_n3872_), .B(new_n16660_), .ZN(new_n16661_));
  XOR2_X1    g16405(.A1(new_n16661_), .A2(new_n3876_), .Z(new_n16662_));
  AOI21_X1   g16406(.A1(new_n16474_), .A2(new_n16581_), .B(new_n16579_), .ZN(new_n16663_));
  AOI22_X1   g16407(.A1(new_n5155_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n5160_), .ZN(new_n16664_));
  OAI21_X1   g16408(.A1(new_n6490_), .A2(new_n6877_), .B(new_n16664_), .ZN(new_n16665_));
  AOI21_X1   g16409(.A1(new_n7906_), .A2(new_n5166_), .B(new_n16665_), .ZN(new_n16666_));
  XOR2_X1    g16410(.A1(new_n16666_), .A2(new_n5162_), .Z(new_n16667_));
  OAI21_X1   g16411(.A1(new_n16480_), .A2(new_n16563_), .B(new_n16565_), .ZN(new_n16668_));
  OAI22_X1   g16412(.A1(new_n5852_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n5857_), .ZN(new_n16669_));
  AOI21_X1   g16413(.A1(\b[39] ), .A2(new_n6115_), .B(new_n16669_), .ZN(new_n16670_));
  OAI21_X1   g16414(.A1(new_n6299_), .A2(new_n5861_), .B(new_n16670_), .ZN(new_n16671_));
  XOR2_X1    g16415(.A1(new_n16671_), .A2(new_n5849_), .Z(new_n16672_));
  AOI22_X1   g16416(.A1(new_n6569_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n6574_), .ZN(new_n16673_));
  OAI21_X1   g16417(.A1(new_n4886_), .A2(new_n8565_), .B(new_n16673_), .ZN(new_n16674_));
  AOI21_X1   g16418(.A1(new_n5351_), .A2(new_n6579_), .B(new_n16674_), .ZN(new_n16675_));
  XOR2_X1    g16419(.A1(new_n16675_), .A2(new_n6567_), .Z(new_n16676_));
  AOI22_X1   g16420(.A1(new_n8241_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n8246_), .ZN(new_n16677_));
  OAI21_X1   g16421(.A1(new_n3624_), .A2(new_n9114_), .B(new_n16677_), .ZN(new_n16678_));
  AOI21_X1   g16422(.A1(new_n4030_), .A2(new_n8252_), .B(new_n16678_), .ZN(new_n16679_));
  XOR2_X1    g16423(.A1(new_n16679_), .A2(new_n8248_), .Z(new_n16680_));
  INV_X1     g16424(.I(new_n16680_), .ZN(new_n16681_));
  AOI22_X1   g16425(.A1(new_n10064_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n10062_), .ZN(new_n16682_));
  OAI21_X1   g16426(.A1(new_n2495_), .A2(new_n10399_), .B(new_n16682_), .ZN(new_n16683_));
  AOI21_X1   g16427(.A1(new_n3407_), .A2(new_n10068_), .B(new_n16683_), .ZN(new_n16684_));
  XOR2_X1    g16428(.A1(new_n16684_), .A2(new_n10057_), .Z(new_n16685_));
  OAI21_X1   g16429(.A1(new_n16502_), .A2(new_n16519_), .B(new_n16520_), .ZN(new_n16686_));
  AOI22_X1   g16430(.A1(new_n10981_), .A2(\b[23] ), .B1(new_n10979_), .B2(\b[22] ), .ZN(new_n16687_));
  OAI21_X1   g16431(.A1(new_n2027_), .A2(new_n11306_), .B(new_n16687_), .ZN(new_n16688_));
  AOI21_X1   g16432(.A1(new_n2470_), .A2(new_n10984_), .B(new_n16688_), .ZN(new_n16689_));
  XOR2_X1    g16433(.A1(new_n16689_), .A2(new_n10989_), .Z(new_n16690_));
  AOI21_X1   g16434(.A1(new_n16509_), .A2(new_n16514_), .B(new_n16515_), .ZN(new_n16691_));
  NOR2_X1    g16435(.A1(new_n16690_), .A2(new_n16691_), .ZN(new_n16692_));
  INV_X1     g16436(.I(new_n16692_), .ZN(new_n16693_));
  NAND2_X1   g16437(.A1(new_n16690_), .A2(new_n16691_), .ZN(new_n16694_));
  NAND2_X1   g16438(.A1(new_n16693_), .A2(new_n16694_), .ZN(new_n16695_));
  AOI22_X1   g16439(.A1(new_n11926_), .A2(\b[20] ), .B1(new_n11924_), .B2(\b[19] ), .ZN(new_n16696_));
  OAI21_X1   g16440(.A1(new_n1553_), .A2(new_n12317_), .B(new_n16696_), .ZN(new_n16697_));
  AOI21_X1   g16441(.A1(new_n2452_), .A2(new_n11929_), .B(new_n16697_), .ZN(new_n16698_));
  XOR2_X1    g16442(.A1(new_n16698_), .A2(new_n12312_), .Z(new_n16699_));
  AOI22_X1   g16443(.A1(new_n12922_), .A2(\b[17] ), .B1(\b[16] ), .B2(new_n12923_), .ZN(new_n16700_));
  INV_X1     g16444(.I(new_n16700_), .ZN(new_n16701_));
  NOR2_X1    g16445(.A1(new_n16701_), .A2(new_n16513_), .ZN(new_n16702_));
  INV_X1     g16446(.I(new_n16702_), .ZN(new_n16703_));
  NAND2_X1   g16447(.A1(new_n16701_), .A2(new_n16513_), .ZN(new_n16704_));
  NAND2_X1   g16448(.A1(new_n16703_), .A2(new_n16704_), .ZN(new_n16705_));
  XNOR2_X1   g16449(.A1(new_n16699_), .A2(new_n16705_), .ZN(new_n16706_));
  XOR2_X1    g16450(.A1(new_n16695_), .A2(new_n16706_), .Z(new_n16707_));
  NOR2_X1    g16451(.A1(new_n16707_), .A2(new_n16686_), .ZN(new_n16708_));
  INV_X1     g16452(.I(new_n16708_), .ZN(new_n16709_));
  NAND2_X1   g16453(.A1(new_n16707_), .A2(new_n16686_), .ZN(new_n16710_));
  NAND2_X1   g16454(.A1(new_n16709_), .A2(new_n16710_), .ZN(new_n16711_));
  XOR2_X1    g16455(.A1(new_n16711_), .A2(new_n16685_), .Z(new_n16712_));
  AOI22_X1   g16456(.A1(new_n9125_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n9123_), .ZN(new_n16713_));
  OAI21_X1   g16457(.A1(new_n3158_), .A2(new_n9470_), .B(new_n16713_), .ZN(new_n16714_));
  AOI21_X1   g16458(.A1(new_n4188_), .A2(new_n9129_), .B(new_n16714_), .ZN(new_n16715_));
  XOR2_X1    g16459(.A1(new_n16715_), .A2(new_n9133_), .Z(new_n16716_));
  AOI21_X1   g16460(.A1(new_n16524_), .A2(new_n16532_), .B(new_n16530_), .ZN(new_n16717_));
  NOR2_X1    g16461(.A1(new_n16716_), .A2(new_n16717_), .ZN(new_n16718_));
  INV_X1     g16462(.I(new_n16718_), .ZN(new_n16719_));
  NAND2_X1   g16463(.A1(new_n16716_), .A2(new_n16717_), .ZN(new_n16720_));
  NAND2_X1   g16464(.A1(new_n16719_), .A2(new_n16720_), .ZN(new_n16721_));
  XOR2_X1    g16465(.A1(new_n16721_), .A2(new_n16712_), .Z(new_n16722_));
  INV_X1     g16466(.I(new_n16496_), .ZN(new_n16723_));
  AOI21_X1   g16467(.A1(new_n16723_), .A2(new_n16537_), .B(new_n16535_), .ZN(new_n16724_));
  NOR2_X1    g16468(.A1(new_n16722_), .A2(new_n16724_), .ZN(new_n16725_));
  INV_X1     g16469(.I(new_n16725_), .ZN(new_n16726_));
  NAND2_X1   g16470(.A1(new_n16722_), .A2(new_n16724_), .ZN(new_n16727_));
  NAND2_X1   g16471(.A1(new_n16726_), .A2(new_n16727_), .ZN(new_n16728_));
  XOR2_X1    g16472(.A1(new_n16728_), .A2(new_n16681_), .Z(new_n16729_));
  INV_X1     g16473(.I(new_n16729_), .ZN(new_n16730_));
  OAI22_X1   g16474(.A1(new_n4639_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n4666_), .ZN(new_n16731_));
  AOI21_X1   g16475(.A1(\b[33] ), .A2(new_n7719_), .B(new_n16731_), .ZN(new_n16732_));
  OAI21_X1   g16476(.A1(new_n4676_), .A2(new_n8585_), .B(new_n16732_), .ZN(new_n16733_));
  XOR2_X1    g16477(.A1(new_n16733_), .A2(\a[47] ), .Z(new_n16734_));
  AOI21_X1   g16478(.A1(new_n16539_), .A2(new_n16547_), .B(new_n16545_), .ZN(new_n16735_));
  NOR2_X1    g16479(.A1(new_n16734_), .A2(new_n16735_), .ZN(new_n16736_));
  INV_X1     g16480(.I(new_n16736_), .ZN(new_n16737_));
  NAND2_X1   g16481(.A1(new_n16734_), .A2(new_n16735_), .ZN(new_n16738_));
  NAND2_X1   g16482(.A1(new_n16737_), .A2(new_n16738_), .ZN(new_n16739_));
  XOR2_X1    g16483(.A1(new_n16739_), .A2(new_n16730_), .Z(new_n16740_));
  AOI21_X1   g16484(.A1(new_n16492_), .A2(new_n16555_), .B(new_n16553_), .ZN(new_n16741_));
  XOR2_X1    g16485(.A1(new_n16740_), .A2(new_n16741_), .Z(new_n16742_));
  XOR2_X1    g16486(.A1(new_n16742_), .A2(new_n16676_), .Z(new_n16743_));
  INV_X1     g16487(.I(new_n16486_), .ZN(new_n16744_));
  AOI21_X1   g16488(.A1(new_n16744_), .A2(new_n16558_), .B(new_n16559_), .ZN(new_n16745_));
  NOR2_X1    g16489(.A1(new_n16743_), .A2(new_n16745_), .ZN(new_n16746_));
  INV_X1     g16490(.I(new_n16746_), .ZN(new_n16747_));
  NAND2_X1   g16491(.A1(new_n16743_), .A2(new_n16745_), .ZN(new_n16748_));
  NAND2_X1   g16492(.A1(new_n16747_), .A2(new_n16748_), .ZN(new_n16749_));
  XNOR2_X1   g16493(.A1(new_n16749_), .A2(new_n16672_), .ZN(new_n16750_));
  NOR2_X1    g16494(.A1(new_n16750_), .A2(new_n16668_), .ZN(new_n16751_));
  NAND2_X1   g16495(.A1(new_n16750_), .A2(new_n16668_), .ZN(new_n16752_));
  INV_X1     g16496(.I(new_n16752_), .ZN(new_n16753_));
  NOR2_X1    g16497(.A1(new_n16753_), .A2(new_n16751_), .ZN(new_n16754_));
  XOR2_X1    g16498(.A1(new_n16754_), .A2(new_n16667_), .Z(new_n16755_));
  AOI22_X1   g16499(.A1(new_n4918_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n4921_), .ZN(new_n16756_));
  OAI21_X1   g16500(.A1(new_n7096_), .A2(new_n6099_), .B(new_n16756_), .ZN(new_n16757_));
  AOI21_X1   g16501(.A1(new_n7649_), .A2(new_n4699_), .B(new_n16757_), .ZN(new_n16758_));
  XOR2_X1    g16502(.A1(new_n16758_), .A2(new_n4446_), .Z(new_n16759_));
  NOR2_X1    g16503(.A1(new_n16575_), .A2(new_n16476_), .ZN(new_n16760_));
  NOR2_X1    g16504(.A1(new_n16760_), .A2(new_n16573_), .ZN(new_n16761_));
  NOR2_X1    g16505(.A1(new_n16761_), .A2(new_n16759_), .ZN(new_n16762_));
  AND2_X2    g16506(.A1(new_n16761_), .A2(new_n16759_), .Z(new_n16763_));
  NOR2_X1    g16507(.A1(new_n16763_), .A2(new_n16762_), .ZN(new_n16764_));
  XOR2_X1    g16508(.A1(new_n16764_), .A2(new_n16755_), .Z(new_n16765_));
  NOR2_X1    g16509(.A1(new_n16765_), .A2(new_n16663_), .ZN(new_n16766_));
  INV_X1     g16510(.I(new_n16766_), .ZN(new_n16767_));
  NAND2_X1   g16511(.A1(new_n16765_), .A2(new_n16663_), .ZN(new_n16768_));
  NAND2_X1   g16512(.A1(new_n16767_), .A2(new_n16768_), .ZN(new_n16769_));
  XOR2_X1    g16513(.A1(new_n16769_), .A2(new_n16662_), .Z(new_n16770_));
  AOI21_X1   g16514(.A1(new_n16467_), .A2(new_n16586_), .B(new_n16584_), .ZN(new_n16771_));
  INV_X1     g16515(.I(new_n16771_), .ZN(new_n16772_));
  NAND2_X1   g16516(.A1(new_n16770_), .A2(new_n16772_), .ZN(new_n16773_));
  OR2_X2     g16517(.A1(new_n16770_), .A2(new_n16772_), .Z(new_n16774_));
  NAND2_X1   g16518(.A1(new_n16774_), .A2(new_n16773_), .ZN(new_n16775_));
  XOR2_X1    g16519(.A1(new_n16775_), .A2(new_n16658_), .Z(new_n16776_));
  XOR2_X1    g16520(.A1(new_n16776_), .A2(new_n16654_), .Z(new_n16777_));
  XOR2_X1    g16521(.A1(new_n16777_), .A2(new_n16652_), .Z(new_n16778_));
  OR2_X2     g16522(.A1(new_n16648_), .A2(new_n16778_), .Z(new_n16779_));
  NAND2_X1   g16523(.A1(new_n16648_), .A2(new_n16778_), .ZN(new_n16780_));
  NAND2_X1   g16524(.A1(new_n16779_), .A2(new_n16780_), .ZN(new_n16781_));
  XOR2_X1    g16525(.A1(new_n16781_), .A2(new_n16647_), .Z(new_n16782_));
  XOR2_X1    g16526(.A1(new_n16642_), .A2(new_n16782_), .Z(new_n16783_));
  XOR2_X1    g16527(.A1(new_n16783_), .A2(new_n16640_), .Z(new_n16784_));
  INV_X1     g16528(.I(new_n16784_), .ZN(new_n16785_));
  XOR2_X1    g16529(.A1(new_n16635_), .A2(new_n16785_), .Z(new_n16786_));
  XOR2_X1    g16530(.A1(new_n16786_), .A2(new_n16632_), .Z(new_n16787_));
  NAND2_X1   g16531(.A1(new_n16787_), .A2(new_n16630_), .ZN(new_n16788_));
  INV_X1     g16532(.I(new_n16788_), .ZN(new_n16789_));
  NOR2_X1    g16533(.A1(new_n16787_), .A2(new_n16630_), .ZN(new_n16790_));
  NOR2_X1    g16534(.A1(new_n16789_), .A2(new_n16790_), .ZN(new_n16791_));
  INV_X1     g16535(.I(new_n16791_), .ZN(new_n16792_));
  XOR2_X1    g16536(.A1(new_n16628_), .A2(new_n16792_), .Z(\f[80] ));
  NOR2_X1    g16537(.A1(new_n16635_), .A2(new_n16785_), .ZN(new_n16794_));
  AOI21_X1   g16538(.A1(new_n16635_), .A2(new_n16785_), .B(new_n16632_), .ZN(new_n16795_));
  NOR2_X1    g16539(.A1(new_n16795_), .A2(new_n16794_), .ZN(new_n16796_));
  NOR2_X1    g16540(.A1(new_n16642_), .A2(new_n16782_), .ZN(new_n16797_));
  NAND2_X1   g16541(.A1(new_n16642_), .A2(new_n16782_), .ZN(new_n16798_));
  AOI21_X1   g16542(.A1(new_n16640_), .A2(new_n16798_), .B(new_n16797_), .ZN(new_n16799_));
  INV_X1     g16543(.I(new_n16799_), .ZN(new_n16800_));
  AOI22_X1   g16544(.A1(new_n1738_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n1743_), .ZN(new_n16801_));
  OAI21_X1   g16545(.A1(new_n12148_), .A2(new_n1931_), .B(new_n16801_), .ZN(new_n16802_));
  AOI21_X1   g16546(.A1(new_n12811_), .A2(new_n1746_), .B(new_n16802_), .ZN(new_n16803_));
  XOR2_X1    g16547(.A1(new_n16803_), .A2(new_n1736_), .Z(new_n16804_));
  AOI22_X1   g16548(.A1(new_n2202_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n2205_), .ZN(new_n16805_));
  OAI21_X1   g16549(.A1(new_n11195_), .A2(new_n2370_), .B(new_n16805_), .ZN(new_n16806_));
  AOI21_X1   g16550(.A1(new_n11836_), .A2(new_n2208_), .B(new_n16806_), .ZN(new_n16807_));
  XOR2_X1    g16551(.A1(new_n16807_), .A2(\a[23] ), .Z(new_n16808_));
  NAND2_X1   g16552(.A1(new_n16780_), .A2(new_n16647_), .ZN(new_n16809_));
  NAND2_X1   g16553(.A1(new_n16809_), .A2(new_n16779_), .ZN(new_n16810_));
  INV_X1     g16554(.I(new_n16652_), .ZN(new_n16811_));
  NOR2_X1    g16555(.A1(new_n16776_), .A2(new_n16654_), .ZN(new_n16812_));
  NAND2_X1   g16556(.A1(new_n16776_), .A2(new_n16654_), .ZN(new_n16813_));
  AOI21_X1   g16557(.A1(new_n16811_), .A2(new_n16813_), .B(new_n16812_), .ZN(new_n16814_));
  INV_X1     g16558(.I(new_n16814_), .ZN(new_n16815_));
  AOI22_X1   g16559(.A1(new_n3267_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n3270_), .ZN(new_n16816_));
  OAI21_X1   g16560(.A1(new_n9032_), .A2(new_n3475_), .B(new_n16816_), .ZN(new_n16817_));
  AOI21_X1   g16561(.A1(new_n10884_), .A2(new_n3273_), .B(new_n16817_), .ZN(new_n16818_));
  XOR2_X1    g16562(.A1(new_n16818_), .A2(new_n3264_), .Z(new_n16819_));
  NAND2_X1   g16563(.A1(new_n16774_), .A2(new_n16658_), .ZN(new_n16820_));
  NAND2_X1   g16564(.A1(new_n16820_), .A2(new_n16773_), .ZN(new_n16821_));
  INV_X1     g16565(.I(new_n16821_), .ZN(new_n16822_));
  INV_X1     g16566(.I(new_n16662_), .ZN(new_n16823_));
  AOI21_X1   g16567(.A1(new_n16823_), .A2(new_n16768_), .B(new_n16766_), .ZN(new_n16824_));
  INV_X1     g16568(.I(new_n16824_), .ZN(new_n16825_));
  OAI21_X1   g16569(.A1(new_n16667_), .A2(new_n16751_), .B(new_n16752_), .ZN(new_n16826_));
  AOI21_X1   g16570(.A1(new_n16672_), .A2(new_n16748_), .B(new_n16746_), .ZN(new_n16827_));
  INV_X1     g16571(.I(new_n16827_), .ZN(new_n16828_));
  INV_X1     g16572(.I(new_n16676_), .ZN(new_n16829_));
  NOR2_X1    g16573(.A1(new_n16740_), .A2(new_n16741_), .ZN(new_n16830_));
  NAND2_X1   g16574(.A1(new_n16740_), .A2(new_n16741_), .ZN(new_n16831_));
  AOI21_X1   g16575(.A1(new_n16829_), .A2(new_n16831_), .B(new_n16830_), .ZN(new_n16832_));
  AOI21_X1   g16576(.A1(new_n16730_), .A2(new_n16738_), .B(new_n16736_), .ZN(new_n16833_));
  INV_X1     g16577(.I(new_n16833_), .ZN(new_n16834_));
  AOI22_X1   g16578(.A1(new_n7403_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n7408_), .ZN(new_n16835_));
  OAI21_X1   g16579(.A1(new_n4639_), .A2(new_n9488_), .B(new_n16835_), .ZN(new_n16836_));
  AOI21_X1   g16580(.A1(new_n5594_), .A2(new_n7414_), .B(new_n16836_), .ZN(new_n16837_));
  XOR2_X1    g16581(.A1(new_n16837_), .A2(new_n7410_), .Z(new_n16838_));
  AOI21_X1   g16582(.A1(new_n16681_), .A2(new_n16727_), .B(new_n16725_), .ZN(new_n16839_));
  INV_X1     g16583(.I(new_n16839_), .ZN(new_n16840_));
  OAI21_X1   g16584(.A1(new_n16685_), .A2(new_n16708_), .B(new_n16710_), .ZN(new_n16841_));
  INV_X1     g16585(.I(new_n16706_), .ZN(new_n16842_));
  AOI21_X1   g16586(.A1(new_n16694_), .A2(new_n16842_), .B(new_n16692_), .ZN(new_n16843_));
  AOI22_X1   g16587(.A1(new_n10981_), .A2(\b[24] ), .B1(new_n10979_), .B2(\b[23] ), .ZN(new_n16844_));
  OAI21_X1   g16588(.A1(new_n2142_), .A2(new_n11306_), .B(new_n16844_), .ZN(new_n16845_));
  AOI21_X1   g16589(.A1(new_n3033_), .A2(new_n10984_), .B(new_n16845_), .ZN(new_n16846_));
  XOR2_X1    g16590(.A1(new_n16846_), .A2(new_n10989_), .Z(new_n16847_));
  OAI21_X1   g16591(.A1(new_n16699_), .A2(new_n16702_), .B(new_n16704_), .ZN(new_n16848_));
  INV_X1     g16592(.I(new_n16848_), .ZN(new_n16849_));
  AOI22_X1   g16593(.A1(new_n11926_), .A2(\b[21] ), .B1(new_n11924_), .B2(\b[20] ), .ZN(new_n16850_));
  OAI21_X1   g16594(.A1(new_n1859_), .A2(new_n12317_), .B(new_n16850_), .ZN(new_n16851_));
  AOI21_X1   g16595(.A1(new_n2032_), .A2(new_n11929_), .B(new_n16851_), .ZN(new_n16852_));
  XOR2_X1    g16596(.A1(new_n16852_), .A2(new_n12312_), .Z(new_n16853_));
  INV_X1     g16597(.I(new_n16853_), .ZN(new_n16854_));
  AOI22_X1   g16598(.A1(new_n12922_), .A2(\b[18] ), .B1(\b[17] ), .B2(new_n12923_), .ZN(new_n16855_));
  INV_X1     g16599(.I(new_n16855_), .ZN(new_n16856_));
  NOR2_X1    g16600(.A1(new_n16856_), .A2(new_n1344_), .ZN(new_n16857_));
  NOR2_X1    g16601(.A1(new_n16855_), .A2(\a[17] ), .ZN(new_n16858_));
  NOR2_X1    g16602(.A1(new_n16857_), .A2(new_n16858_), .ZN(new_n16859_));
  XOR2_X1    g16603(.A1(new_n16859_), .A2(new_n16700_), .Z(new_n16860_));
  NOR2_X1    g16604(.A1(new_n16854_), .A2(new_n16860_), .ZN(new_n16861_));
  NAND2_X1   g16605(.A1(new_n16854_), .A2(new_n16860_), .ZN(new_n16862_));
  INV_X1     g16606(.I(new_n16862_), .ZN(new_n16863_));
  NOR2_X1    g16607(.A1(new_n16863_), .A2(new_n16861_), .ZN(new_n16864_));
  XOR2_X1    g16608(.A1(new_n16864_), .A2(new_n16849_), .Z(new_n16865_));
  NOR2_X1    g16609(.A1(new_n16865_), .A2(new_n16847_), .ZN(new_n16866_));
  INV_X1     g16610(.I(new_n16866_), .ZN(new_n16867_));
  NAND2_X1   g16611(.A1(new_n16865_), .A2(new_n16847_), .ZN(new_n16868_));
  NAND2_X1   g16612(.A1(new_n16867_), .A2(new_n16868_), .ZN(new_n16869_));
  XOR2_X1    g16613(.A1(new_n16869_), .A2(new_n16843_), .Z(new_n16870_));
  OAI22_X1   g16614(.A1(new_n11298_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n11297_), .ZN(new_n16871_));
  AOI21_X1   g16615(.A1(\b[25] ), .A2(new_n11296_), .B(new_n16871_), .ZN(new_n16872_));
  OAI21_X1   g16616(.A1(new_n3165_), .A2(new_n10069_), .B(new_n16872_), .ZN(new_n16873_));
  XOR2_X1    g16617(.A1(new_n16873_), .A2(new_n10057_), .Z(new_n16874_));
  NAND2_X1   g16618(.A1(new_n16870_), .A2(new_n16874_), .ZN(new_n16875_));
  OR2_X2     g16619(.A1(new_n16870_), .A2(new_n16874_), .Z(new_n16876_));
  NAND2_X1   g16620(.A1(new_n16876_), .A2(new_n16875_), .ZN(new_n16877_));
  XNOR2_X1   g16621(.A1(new_n16877_), .A2(new_n16841_), .ZN(new_n16878_));
  AOI22_X1   g16622(.A1(new_n9125_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n9123_), .ZN(new_n16879_));
  OAI21_X1   g16623(.A1(new_n3185_), .A2(new_n9470_), .B(new_n16879_), .ZN(new_n16880_));
  AOI21_X1   g16624(.A1(new_n4230_), .A2(new_n9129_), .B(new_n16880_), .ZN(new_n16881_));
  XOR2_X1    g16625(.A1(new_n16881_), .A2(new_n9133_), .Z(new_n16882_));
  INV_X1     g16626(.I(new_n16882_), .ZN(new_n16883_));
  NAND2_X1   g16627(.A1(new_n16712_), .A2(new_n16720_), .ZN(new_n16884_));
  NAND2_X1   g16628(.A1(new_n16884_), .A2(new_n16719_), .ZN(new_n16885_));
  NAND2_X1   g16629(.A1(new_n16885_), .A2(new_n16883_), .ZN(new_n16886_));
  NAND3_X1   g16630(.A1(new_n16884_), .A2(new_n16719_), .A3(new_n16882_), .ZN(new_n16887_));
  NAND2_X1   g16631(.A1(new_n16886_), .A2(new_n16887_), .ZN(new_n16888_));
  XNOR2_X1   g16632(.A1(new_n16878_), .A2(new_n16888_), .ZN(new_n16889_));
  INV_X1     g16633(.I(new_n16889_), .ZN(new_n16890_));
  AOI22_X1   g16634(.A1(new_n8241_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n8246_), .ZN(new_n16891_));
  OAI21_X1   g16635(.A1(new_n4022_), .A2(new_n9114_), .B(new_n16891_), .ZN(new_n16892_));
  AOI21_X1   g16636(.A1(new_n4223_), .A2(new_n8252_), .B(new_n16892_), .ZN(new_n16893_));
  XOR2_X1    g16637(.A1(new_n16893_), .A2(new_n8248_), .Z(new_n16894_));
  NOR2_X1    g16638(.A1(new_n16890_), .A2(new_n16894_), .ZN(new_n16895_));
  INV_X1     g16639(.I(new_n16895_), .ZN(new_n16896_));
  NAND2_X1   g16640(.A1(new_n16890_), .A2(new_n16894_), .ZN(new_n16897_));
  NAND2_X1   g16641(.A1(new_n16896_), .A2(new_n16897_), .ZN(new_n16898_));
  XOR2_X1    g16642(.A1(new_n16898_), .A2(new_n16840_), .Z(new_n16899_));
  NOR2_X1    g16643(.A1(new_n16899_), .A2(new_n16838_), .ZN(new_n16900_));
  NAND2_X1   g16644(.A1(new_n16899_), .A2(new_n16838_), .ZN(new_n16901_));
  INV_X1     g16645(.I(new_n16901_), .ZN(new_n16902_));
  NOR2_X1    g16646(.A1(new_n16902_), .A2(new_n16900_), .ZN(new_n16903_));
  XOR2_X1    g16647(.A1(new_n16903_), .A2(new_n16834_), .Z(new_n16904_));
  INV_X1     g16648(.I(new_n16904_), .ZN(new_n16905_));
  AOI22_X1   g16649(.A1(new_n6569_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n6574_), .ZN(new_n16906_));
  OAI21_X1   g16650(.A1(new_n5312_), .A2(new_n8565_), .B(new_n16906_), .ZN(new_n16907_));
  AOI21_X1   g16651(.A1(new_n6310_), .A2(new_n6579_), .B(new_n16907_), .ZN(new_n16908_));
  XOR2_X1    g16652(.A1(new_n16908_), .A2(new_n6567_), .Z(new_n16909_));
  NOR2_X1    g16653(.A1(new_n16905_), .A2(new_n16909_), .ZN(new_n16910_));
  NAND2_X1   g16654(.A1(new_n16905_), .A2(new_n16909_), .ZN(new_n16911_));
  INV_X1     g16655(.I(new_n16911_), .ZN(new_n16912_));
  NOR2_X1    g16656(.A1(new_n16912_), .A2(new_n16910_), .ZN(new_n16913_));
  XOR2_X1    g16657(.A1(new_n16913_), .A2(new_n16832_), .Z(new_n16914_));
  AOI22_X1   g16658(.A1(new_n6108_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n6111_), .ZN(new_n16915_));
  OAI21_X1   g16659(.A1(new_n6284_), .A2(new_n7708_), .B(new_n16915_), .ZN(new_n16916_));
  AOI21_X1   g16660(.A1(new_n7106_), .A2(new_n6105_), .B(new_n16916_), .ZN(new_n16917_));
  XOR2_X1    g16661(.A1(new_n16917_), .A2(new_n5849_), .Z(new_n16918_));
  NOR2_X1    g16662(.A1(new_n16914_), .A2(new_n16918_), .ZN(new_n16919_));
  NAND2_X1   g16663(.A1(new_n16914_), .A2(new_n16918_), .ZN(new_n16920_));
  INV_X1     g16664(.I(new_n16920_), .ZN(new_n16921_));
  NOR2_X1    g16665(.A1(new_n16921_), .A2(new_n16919_), .ZN(new_n16922_));
  XOR2_X1    g16666(.A1(new_n16922_), .A2(new_n16828_), .Z(new_n16923_));
  INV_X1     g16667(.I(new_n16923_), .ZN(new_n16924_));
  AOI22_X1   g16668(.A1(new_n5155_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n5160_), .ZN(new_n16925_));
  OAI21_X1   g16669(.A1(new_n6775_), .A2(new_n6877_), .B(new_n16925_), .ZN(new_n16926_));
  AOI21_X1   g16670(.A1(new_n7926_), .A2(new_n5166_), .B(new_n16926_), .ZN(new_n16927_));
  XOR2_X1    g16671(.A1(new_n16927_), .A2(new_n5162_), .Z(new_n16928_));
  NOR2_X1    g16672(.A1(new_n16924_), .A2(new_n16928_), .ZN(new_n16929_));
  NAND2_X1   g16673(.A1(new_n16924_), .A2(new_n16928_), .ZN(new_n16930_));
  INV_X1     g16674(.I(new_n16930_), .ZN(new_n16931_));
  NOR2_X1    g16675(.A1(new_n16931_), .A2(new_n16929_), .ZN(new_n16932_));
  XOR2_X1    g16676(.A1(new_n16932_), .A2(new_n16826_), .Z(new_n16933_));
  AOI22_X1   g16677(.A1(new_n4918_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n4921_), .ZN(new_n16934_));
  OAI21_X1   g16678(.A1(new_n7617_), .A2(new_n6099_), .B(new_n16934_), .ZN(new_n16935_));
  AOI21_X1   g16679(.A1(new_n8792_), .A2(new_n4699_), .B(new_n16935_), .ZN(new_n16936_));
  XOR2_X1    g16680(.A1(new_n16936_), .A2(\a[35] ), .Z(new_n16937_));
  INV_X1     g16681(.I(new_n16762_), .ZN(new_n16938_));
  OAI21_X1   g16682(.A1(new_n16755_), .A2(new_n16763_), .B(new_n16938_), .ZN(new_n16939_));
  NAND2_X1   g16683(.A1(new_n16939_), .A2(new_n16937_), .ZN(new_n16940_));
  OR2_X2     g16684(.A1(new_n16939_), .A2(new_n16937_), .Z(new_n16941_));
  NAND2_X1   g16685(.A1(new_n16941_), .A2(new_n16940_), .ZN(new_n16942_));
  XNOR2_X1   g16686(.A1(new_n16933_), .A2(new_n16942_), .ZN(new_n16943_));
  INV_X1     g16687(.I(new_n16943_), .ZN(new_n16944_));
  AOI22_X1   g16688(.A1(new_n3864_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n3869_), .ZN(new_n16945_));
  OAI21_X1   g16689(.A1(new_n8168_), .A2(new_n5410_), .B(new_n16945_), .ZN(new_n16946_));
  AOI21_X1   g16690(.A1(new_n8783_), .A2(new_n3872_), .B(new_n16946_), .ZN(new_n16947_));
  XOR2_X1    g16691(.A1(new_n16947_), .A2(new_n3876_), .Z(new_n16948_));
  NOR2_X1    g16692(.A1(new_n16944_), .A2(new_n16948_), .ZN(new_n16949_));
  INV_X1     g16693(.I(new_n16949_), .ZN(new_n16950_));
  NAND2_X1   g16694(.A1(new_n16944_), .A2(new_n16948_), .ZN(new_n16951_));
  NAND2_X1   g16695(.A1(new_n16950_), .A2(new_n16951_), .ZN(new_n16952_));
  XOR2_X1    g16696(.A1(new_n16952_), .A2(new_n16825_), .Z(new_n16953_));
  NOR2_X1    g16697(.A1(new_n16822_), .A2(new_n16953_), .ZN(new_n16954_));
  NAND2_X1   g16698(.A1(new_n16822_), .A2(new_n16953_), .ZN(new_n16955_));
  INV_X1     g16699(.I(new_n16955_), .ZN(new_n16956_));
  NOR2_X1    g16700(.A1(new_n16956_), .A2(new_n16954_), .ZN(new_n16957_));
  XOR2_X1    g16701(.A1(new_n16957_), .A2(new_n16819_), .Z(new_n16958_));
  AOI22_X1   g16702(.A1(new_n2716_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n2719_), .ZN(new_n16959_));
  OAI21_X1   g16703(.A1(new_n9972_), .A2(new_n2924_), .B(new_n16959_), .ZN(new_n16960_));
  AOI21_X1   g16704(.A1(new_n10631_), .A2(new_n2722_), .B(new_n16960_), .ZN(new_n16961_));
  XOR2_X1    g16705(.A1(new_n16961_), .A2(new_n2714_), .Z(new_n16962_));
  NOR2_X1    g16706(.A1(new_n16958_), .A2(new_n16962_), .ZN(new_n16963_));
  NAND2_X1   g16707(.A1(new_n16958_), .A2(new_n16962_), .ZN(new_n16964_));
  INV_X1     g16708(.I(new_n16964_), .ZN(new_n16965_));
  NOR2_X1    g16709(.A1(new_n16965_), .A2(new_n16963_), .ZN(new_n16966_));
  XOR2_X1    g16710(.A1(new_n16966_), .A2(new_n16815_), .Z(new_n16967_));
  XNOR2_X1   g16711(.A1(new_n16967_), .A2(new_n16810_), .ZN(new_n16968_));
  XOR2_X1    g16712(.A1(new_n16968_), .A2(new_n16808_), .Z(new_n16969_));
  NOR2_X1    g16713(.A1(new_n16969_), .A2(new_n16804_), .ZN(new_n16970_));
  INV_X1     g16714(.I(new_n16970_), .ZN(new_n16971_));
  NAND2_X1   g16715(.A1(new_n16969_), .A2(new_n16804_), .ZN(new_n16972_));
  NAND2_X1   g16716(.A1(new_n16971_), .A2(new_n16972_), .ZN(new_n16973_));
  XOR2_X1    g16717(.A1(new_n16973_), .A2(new_n16800_), .Z(new_n16974_));
  NOR2_X1    g16718(.A1(new_n16974_), .A2(new_n16796_), .ZN(new_n16975_));
  NAND2_X1   g16719(.A1(new_n16974_), .A2(new_n16796_), .ZN(new_n16976_));
  INV_X1     g16720(.I(new_n16976_), .ZN(new_n16977_));
  NOR2_X1    g16721(.A1(new_n16977_), .A2(new_n16975_), .ZN(new_n16978_));
  OAI21_X1   g16722(.A1(new_n16628_), .A2(new_n16792_), .B(new_n16788_), .ZN(new_n16979_));
  XOR2_X1    g16723(.A1(new_n16979_), .A2(new_n16978_), .Z(\f[81] ));
  AOI21_X1   g16724(.A1(new_n16800_), .A2(new_n16972_), .B(new_n16970_), .ZN(new_n16981_));
  OAI22_X1   g16725(.A1(new_n1931_), .A2(new_n12796_), .B1(new_n12800_), .B2(new_n1754_), .ZN(new_n16982_));
  AOI21_X1   g16726(.A1(new_n13973_), .A2(new_n1746_), .B(new_n16982_), .ZN(new_n16983_));
  XOR2_X1    g16727(.A1(new_n16983_), .A2(new_n1736_), .Z(new_n16984_));
  NAND2_X1   g16728(.A1(new_n16967_), .A2(new_n16810_), .ZN(new_n16985_));
  OAI21_X1   g16729(.A1(new_n16967_), .A2(new_n16810_), .B(new_n16808_), .ZN(new_n16986_));
  NAND2_X1   g16730(.A1(new_n16986_), .A2(new_n16985_), .ZN(new_n16987_));
  OAI22_X1   g16731(.A1(new_n2189_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n2194_), .ZN(new_n16988_));
  AOI21_X1   g16732(.A1(\b[59] ), .A2(new_n2361_), .B(new_n16988_), .ZN(new_n16989_));
  OAI21_X1   g16733(.A1(new_n13110_), .A2(new_n2197_), .B(new_n16989_), .ZN(new_n16990_));
  XOR2_X1    g16734(.A1(new_n16990_), .A2(new_n2200_), .Z(new_n16991_));
  AOI21_X1   g16735(.A1(new_n16815_), .A2(new_n16964_), .B(new_n16963_), .ZN(new_n16992_));
  AOI22_X1   g16736(.A1(new_n2716_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n2719_), .ZN(new_n16993_));
  OAI21_X1   g16737(.A1(new_n10308_), .A2(new_n2924_), .B(new_n16993_), .ZN(new_n16994_));
  AOI21_X1   g16738(.A1(new_n12164_), .A2(new_n2722_), .B(new_n16994_), .ZN(new_n16995_));
  XOR2_X1    g16739(.A1(new_n16995_), .A2(new_n2714_), .Z(new_n16996_));
  NOR2_X1    g16740(.A1(new_n16956_), .A2(new_n16819_), .ZN(new_n16997_));
  NOR2_X1    g16741(.A1(new_n16997_), .A2(new_n16954_), .ZN(new_n16998_));
  AOI22_X1   g16742(.A1(new_n3267_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n3270_), .ZN(new_n16999_));
  OAI21_X1   g16743(.A1(new_n9376_), .A2(new_n3475_), .B(new_n16999_), .ZN(new_n17000_));
  AOI21_X1   g16744(.A1(new_n9979_), .A2(new_n3273_), .B(new_n17000_), .ZN(new_n17001_));
  XOR2_X1    g16745(.A1(new_n17001_), .A2(new_n3264_), .Z(new_n17002_));
  AOI21_X1   g16746(.A1(new_n16825_), .A2(new_n16951_), .B(new_n16949_), .ZN(new_n17003_));
  INV_X1     g16747(.I(new_n17003_), .ZN(new_n17004_));
  AOI22_X1   g16748(.A1(new_n3864_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n3869_), .ZN(new_n17005_));
  OAI21_X1   g16749(.A1(new_n8500_), .A2(new_n5410_), .B(new_n17005_), .ZN(new_n17006_));
  AOI21_X1   g16750(.A1(new_n9987_), .A2(new_n3872_), .B(new_n17006_), .ZN(new_n17007_));
  XOR2_X1    g16751(.A1(new_n17007_), .A2(new_n3876_), .Z(new_n17008_));
  INV_X1     g16752(.I(new_n16940_), .ZN(new_n17009_));
  AOI21_X1   g16753(.A1(new_n16933_), .A2(new_n16941_), .B(new_n17009_), .ZN(new_n17010_));
  AOI22_X1   g16754(.A1(new_n5155_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n5160_), .ZN(new_n17011_));
  OAI21_X1   g16755(.A1(new_n7074_), .A2(new_n6877_), .B(new_n17011_), .ZN(new_n17012_));
  AOI21_X1   g16756(.A1(new_n9337_), .A2(new_n5166_), .B(new_n17012_), .ZN(new_n17013_));
  XOR2_X1    g16757(.A1(new_n17013_), .A2(new_n5162_), .Z(new_n17014_));
  INV_X1     g16758(.I(new_n17014_), .ZN(new_n17015_));
  NOR2_X1    g16759(.A1(new_n16912_), .A2(new_n16832_), .ZN(new_n17016_));
  NOR2_X1    g16760(.A1(new_n17016_), .A2(new_n16910_), .ZN(new_n17017_));
  AOI22_X1   g16761(.A1(new_n6569_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n6574_), .ZN(new_n17018_));
  OAI21_X1   g16762(.A1(new_n5341_), .A2(new_n8565_), .B(new_n17018_), .ZN(new_n17019_));
  AOI21_X1   g16763(.A1(new_n5793_), .A2(new_n6579_), .B(new_n17019_), .ZN(new_n17020_));
  XOR2_X1    g16764(.A1(new_n17020_), .A2(new_n6567_), .Z(new_n17021_));
  AOI21_X1   g16765(.A1(new_n16834_), .A2(new_n16901_), .B(new_n16900_), .ZN(new_n17022_));
  INV_X1     g16766(.I(new_n17022_), .ZN(new_n17023_));
  AOI22_X1   g16767(.A1(new_n8241_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n8246_), .ZN(new_n17024_));
  OAI21_X1   g16768(.A1(new_n4023_), .A2(new_n9114_), .B(new_n17024_), .ZN(new_n17025_));
  AOI21_X1   g16769(.A1(new_n5103_), .A2(new_n8252_), .B(new_n17025_), .ZN(new_n17026_));
  XOR2_X1    g16770(.A1(new_n17026_), .A2(new_n8248_), .Z(new_n17027_));
  INV_X1     g16771(.I(new_n17027_), .ZN(new_n17028_));
  AOI22_X1   g16772(.A1(new_n10064_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n10062_), .ZN(new_n17029_));
  OAI21_X1   g16773(.A1(new_n3006_), .A2(new_n10399_), .B(new_n17029_), .ZN(new_n17030_));
  AOI21_X1   g16774(.A1(new_n3807_), .A2(new_n10068_), .B(new_n17030_), .ZN(new_n17031_));
  XOR2_X1    g16775(.A1(new_n17031_), .A2(new_n10057_), .Z(new_n17032_));
  INV_X1     g16776(.I(new_n16843_), .ZN(new_n17033_));
  AOI21_X1   g16777(.A1(new_n17033_), .A2(new_n16868_), .B(new_n16866_), .ZN(new_n17034_));
  AOI22_X1   g16778(.A1(new_n11926_), .A2(\b[22] ), .B1(new_n11924_), .B2(\b[21] ), .ZN(new_n17035_));
  OAI21_X1   g16779(.A1(new_n1860_), .A2(new_n12317_), .B(new_n17035_), .ZN(new_n17036_));
  AOI21_X1   g16780(.A1(new_n2659_), .A2(new_n11929_), .B(new_n17036_), .ZN(new_n17037_));
  XOR2_X1    g16781(.A1(new_n17037_), .A2(\a[62] ), .Z(new_n17038_));
  NOR2_X1    g16782(.A1(new_n16858_), .A2(new_n16701_), .ZN(new_n17039_));
  NOR2_X1    g16783(.A1(new_n17039_), .A2(new_n16857_), .ZN(new_n17040_));
  AOI22_X1   g16784(.A1(new_n12922_), .A2(\b[19] ), .B1(\b[18] ), .B2(new_n12923_), .ZN(new_n17041_));
  NAND2_X1   g16785(.A1(new_n17040_), .A2(new_n17041_), .ZN(new_n17042_));
  NOR2_X1    g16786(.A1(new_n17040_), .A2(new_n17041_), .ZN(new_n17043_));
  INV_X1     g16787(.I(new_n17043_), .ZN(new_n17044_));
  NAND2_X1   g16788(.A1(new_n17044_), .A2(new_n17042_), .ZN(new_n17045_));
  XNOR2_X1   g16789(.A1(new_n17038_), .A2(new_n17045_), .ZN(new_n17046_));
  OAI21_X1   g16790(.A1(new_n16849_), .A2(new_n16861_), .B(new_n16862_), .ZN(new_n17047_));
  INV_X1     g16791(.I(new_n17047_), .ZN(new_n17048_));
  OAI22_X1   g16792(.A1(new_n12306_), .A2(new_n2646_), .B1(new_n12305_), .B2(new_n2495_), .ZN(new_n17049_));
  AOI21_X1   g16793(.A1(\b[23] ), .A2(new_n12304_), .B(new_n17049_), .ZN(new_n17050_));
  OAI21_X1   g16794(.A1(new_n2655_), .A2(new_n10985_), .B(new_n17050_), .ZN(new_n17051_));
  XOR2_X1    g16795(.A1(new_n17051_), .A2(\a[59] ), .Z(new_n17052_));
  NOR2_X1    g16796(.A1(new_n17052_), .A2(new_n17048_), .ZN(new_n17053_));
  INV_X1     g16797(.I(new_n17053_), .ZN(new_n17054_));
  NAND2_X1   g16798(.A1(new_n17052_), .A2(new_n17048_), .ZN(new_n17055_));
  NAND2_X1   g16799(.A1(new_n17054_), .A2(new_n17055_), .ZN(new_n17056_));
  XOR2_X1    g16800(.A1(new_n17056_), .A2(new_n17046_), .Z(new_n17057_));
  NOR2_X1    g16801(.A1(new_n17057_), .A2(new_n17034_), .ZN(new_n17058_));
  INV_X1     g16802(.I(new_n17058_), .ZN(new_n17059_));
  NAND2_X1   g16803(.A1(new_n17057_), .A2(new_n17034_), .ZN(new_n17060_));
  NAND2_X1   g16804(.A1(new_n17059_), .A2(new_n17060_), .ZN(new_n17061_));
  XOR2_X1    g16805(.A1(new_n17061_), .A2(new_n17032_), .Z(new_n17062_));
  INV_X1     g16806(.I(new_n16875_), .ZN(new_n17063_));
  AOI21_X1   g16807(.A1(new_n16841_), .A2(new_n16876_), .B(new_n17063_), .ZN(new_n17064_));
  AOI22_X1   g16808(.A1(new_n9125_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n9123_), .ZN(new_n17065_));
  OAI21_X1   g16809(.A1(new_n3592_), .A2(new_n9470_), .B(new_n17065_), .ZN(new_n17066_));
  AOI21_X1   g16810(.A1(new_n3796_), .A2(new_n9129_), .B(new_n17066_), .ZN(new_n17067_));
  XOR2_X1    g16811(.A1(new_n17067_), .A2(new_n9133_), .Z(new_n17068_));
  NOR2_X1    g16812(.A1(new_n17068_), .A2(new_n17064_), .ZN(new_n17069_));
  INV_X1     g16813(.I(new_n17069_), .ZN(new_n17070_));
  NAND2_X1   g16814(.A1(new_n17068_), .A2(new_n17064_), .ZN(new_n17071_));
  NAND2_X1   g16815(.A1(new_n17070_), .A2(new_n17071_), .ZN(new_n17072_));
  XOR2_X1    g16816(.A1(new_n17072_), .A2(new_n17062_), .Z(new_n17073_));
  NAND2_X1   g16817(.A1(new_n16878_), .A2(new_n16887_), .ZN(new_n17074_));
  NAND2_X1   g16818(.A1(new_n17074_), .A2(new_n16886_), .ZN(new_n17075_));
  INV_X1     g16819(.I(new_n17075_), .ZN(new_n17076_));
  NOR2_X1    g16820(.A1(new_n17073_), .A2(new_n17076_), .ZN(new_n17077_));
  INV_X1     g16821(.I(new_n17077_), .ZN(new_n17078_));
  NAND2_X1   g16822(.A1(new_n17073_), .A2(new_n17076_), .ZN(new_n17079_));
  NAND2_X1   g16823(.A1(new_n17078_), .A2(new_n17079_), .ZN(new_n17080_));
  XOR2_X1    g16824(.A1(new_n17080_), .A2(new_n17028_), .Z(new_n17081_));
  AOI21_X1   g16825(.A1(new_n16840_), .A2(new_n16897_), .B(new_n16895_), .ZN(new_n17082_));
  OAI22_X1   g16826(.A1(new_n4886_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n5312_), .ZN(new_n17083_));
  AOI21_X1   g16827(.A1(\b[35] ), .A2(new_n7719_), .B(new_n17083_), .ZN(new_n17084_));
  OAI21_X1   g16828(.A1(new_n5322_), .A2(new_n8585_), .B(new_n17084_), .ZN(new_n17085_));
  XOR2_X1    g16829(.A1(new_n17085_), .A2(\a[47] ), .Z(new_n17086_));
  NOR2_X1    g16830(.A1(new_n17086_), .A2(new_n17082_), .ZN(new_n17087_));
  INV_X1     g16831(.I(new_n17087_), .ZN(new_n17088_));
  NAND2_X1   g16832(.A1(new_n17086_), .A2(new_n17082_), .ZN(new_n17089_));
  NAND2_X1   g16833(.A1(new_n17088_), .A2(new_n17089_), .ZN(new_n17090_));
  XOR2_X1    g16834(.A1(new_n17090_), .A2(new_n17081_), .Z(new_n17091_));
  NOR2_X1    g16835(.A1(new_n17023_), .A2(new_n17091_), .ZN(new_n17092_));
  INV_X1     g16836(.I(new_n17092_), .ZN(new_n17093_));
  NAND2_X1   g16837(.A1(new_n17023_), .A2(new_n17091_), .ZN(new_n17094_));
  NAND2_X1   g16838(.A1(new_n17093_), .A2(new_n17094_), .ZN(new_n17095_));
  XOR2_X1    g16839(.A1(new_n17095_), .A2(new_n17021_), .Z(new_n17096_));
  INV_X1     g16840(.I(new_n17096_), .ZN(new_n17097_));
  OAI22_X1   g16841(.A1(new_n5852_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n5857_), .ZN(new_n17098_));
  AOI21_X1   g16842(.A1(\b[41] ), .A2(new_n6115_), .B(new_n17098_), .ZN(new_n17099_));
  OAI21_X1   g16843(.A1(new_n6785_), .A2(new_n5861_), .B(new_n17099_), .ZN(new_n17100_));
  XOR2_X1    g16844(.A1(new_n17100_), .A2(\a[41] ), .Z(new_n17101_));
  NOR2_X1    g16845(.A1(new_n17097_), .A2(new_n17101_), .ZN(new_n17102_));
  NAND2_X1   g16846(.A1(new_n17097_), .A2(new_n17101_), .ZN(new_n17103_));
  INV_X1     g16847(.I(new_n17103_), .ZN(new_n17104_));
  NOR2_X1    g16848(.A1(new_n17104_), .A2(new_n17102_), .ZN(new_n17105_));
  XOR2_X1    g16849(.A1(new_n17105_), .A2(new_n17017_), .Z(new_n17106_));
  AOI21_X1   g16850(.A1(new_n16828_), .A2(new_n16920_), .B(new_n16919_), .ZN(new_n17107_));
  NOR2_X1    g16851(.A1(new_n17106_), .A2(new_n17107_), .ZN(new_n17108_));
  INV_X1     g16852(.I(new_n17108_), .ZN(new_n17109_));
  NAND2_X1   g16853(.A1(new_n17106_), .A2(new_n17107_), .ZN(new_n17110_));
  NAND2_X1   g16854(.A1(new_n17109_), .A2(new_n17110_), .ZN(new_n17111_));
  XOR2_X1    g16855(.A1(new_n17111_), .A2(new_n17015_), .Z(new_n17112_));
  AOI21_X1   g16856(.A1(new_n16826_), .A2(new_n16930_), .B(new_n16929_), .ZN(new_n17113_));
  OAI22_X1   g16857(.A1(new_n8168_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n8127_), .ZN(new_n17114_));
  AOI21_X1   g16858(.A1(\b[47] ), .A2(new_n4706_), .B(new_n17114_), .ZN(new_n17115_));
  OAI21_X1   g16859(.A1(new_n9050_), .A2(new_n4458_), .B(new_n17115_), .ZN(new_n17116_));
  XOR2_X1    g16860(.A1(new_n17116_), .A2(\a[35] ), .Z(new_n17117_));
  NOR2_X1    g16861(.A1(new_n17113_), .A2(new_n17117_), .ZN(new_n17118_));
  NAND2_X1   g16862(.A1(new_n17113_), .A2(new_n17117_), .ZN(new_n17119_));
  INV_X1     g16863(.I(new_n17119_), .ZN(new_n17120_));
  NOR2_X1    g16864(.A1(new_n17120_), .A2(new_n17118_), .ZN(new_n17121_));
  XOR2_X1    g16865(.A1(new_n17121_), .A2(new_n17112_), .Z(new_n17122_));
  NOR2_X1    g16866(.A1(new_n17122_), .A2(new_n17010_), .ZN(new_n17123_));
  INV_X1     g16867(.I(new_n17123_), .ZN(new_n17124_));
  NAND2_X1   g16868(.A1(new_n17122_), .A2(new_n17010_), .ZN(new_n17125_));
  NAND2_X1   g16869(.A1(new_n17124_), .A2(new_n17125_), .ZN(new_n17126_));
  XOR2_X1    g16870(.A1(new_n17126_), .A2(new_n17008_), .Z(new_n17127_));
  NOR2_X1    g16871(.A1(new_n17127_), .A2(new_n17004_), .ZN(new_n17128_));
  NAND2_X1   g16872(.A1(new_n17127_), .A2(new_n17004_), .ZN(new_n17129_));
  INV_X1     g16873(.I(new_n17129_), .ZN(new_n17130_));
  NOR2_X1    g16874(.A1(new_n17130_), .A2(new_n17128_), .ZN(new_n17131_));
  XOR2_X1    g16875(.A1(new_n17131_), .A2(new_n17002_), .Z(new_n17132_));
  NOR2_X1    g16876(.A1(new_n17132_), .A2(new_n16998_), .ZN(new_n17133_));
  INV_X1     g16877(.I(new_n17133_), .ZN(new_n17134_));
  NAND2_X1   g16878(.A1(new_n17132_), .A2(new_n16998_), .ZN(new_n17135_));
  NAND2_X1   g16879(.A1(new_n17134_), .A2(new_n17135_), .ZN(new_n17136_));
  XOR2_X1    g16880(.A1(new_n17136_), .A2(new_n16996_), .Z(new_n17137_));
  INV_X1     g16881(.I(new_n17137_), .ZN(new_n17138_));
  NAND2_X1   g16882(.A1(new_n17138_), .A2(new_n16992_), .ZN(new_n17139_));
  NOR2_X1    g16883(.A1(new_n17138_), .A2(new_n16992_), .ZN(new_n17140_));
  INV_X1     g16884(.I(new_n17140_), .ZN(new_n17141_));
  NAND2_X1   g16885(.A1(new_n17141_), .A2(new_n17139_), .ZN(new_n17142_));
  XNOR2_X1   g16886(.A1(new_n17142_), .A2(new_n16991_), .ZN(new_n17143_));
  NAND2_X1   g16887(.A1(new_n17143_), .A2(new_n16987_), .ZN(new_n17144_));
  NOR2_X1    g16888(.A1(new_n17143_), .A2(new_n16987_), .ZN(new_n17145_));
  INV_X1     g16889(.I(new_n17145_), .ZN(new_n17146_));
  NAND2_X1   g16890(.A1(new_n17146_), .A2(new_n17144_), .ZN(new_n17147_));
  XOR2_X1    g16891(.A1(new_n17147_), .A2(new_n16984_), .Z(new_n17148_));
  AOI21_X1   g16892(.A1(new_n16979_), .A2(new_n16978_), .B(new_n16977_), .ZN(new_n17149_));
  NOR2_X1    g16893(.A1(new_n17149_), .A2(new_n17148_), .ZN(new_n17150_));
  INV_X1     g16894(.I(new_n17148_), .ZN(new_n17151_));
  NOR3_X1    g16895(.A1(new_n16618_), .A2(new_n16425_), .A3(new_n16616_), .ZN(new_n17152_));
  AOI21_X1   g16896(.A1(new_n16431_), .A2(new_n16619_), .B(new_n17152_), .ZN(new_n17153_));
  AOI21_X1   g16897(.A1(new_n17153_), .A2(new_n16791_), .B(new_n16789_), .ZN(new_n17154_));
  OAI21_X1   g16898(.A1(new_n17154_), .A2(new_n16975_), .B(new_n16976_), .ZN(new_n17155_));
  NOR2_X1    g16899(.A1(new_n17155_), .A2(new_n17151_), .ZN(new_n17156_));
  NOR2_X1    g16900(.A1(new_n17156_), .A2(new_n17150_), .ZN(new_n17157_));
  XOR2_X1    g16901(.A1(new_n17157_), .A2(new_n16981_), .Z(\f[82] ));
  NAND2_X1   g16902(.A1(new_n17149_), .A2(new_n17148_), .ZN(new_n17159_));
  INV_X1     g16903(.I(new_n16981_), .ZN(new_n17160_));
  OAI21_X1   g16904(.A1(new_n17149_), .A2(new_n17148_), .B(new_n17160_), .ZN(new_n17161_));
  NAND2_X1   g16905(.A1(new_n17161_), .A2(new_n17159_), .ZN(new_n17162_));
  OAI21_X1   g16906(.A1(new_n16984_), .A2(new_n17145_), .B(new_n17144_), .ZN(new_n17163_));
  AOI22_X1   g16907(.A1(new_n13460_), .A2(new_n1746_), .B1(\b[63] ), .B2(new_n1939_), .ZN(new_n17164_));
  XOR2_X1    g16908(.A1(new_n17164_), .A2(new_n1736_), .Z(new_n17165_));
  OAI22_X1   g16909(.A1(new_n2703_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n2708_), .ZN(new_n17166_));
  AOI21_X1   g16910(.A1(\b[57] ), .A2(new_n2906_), .B(new_n17166_), .ZN(new_n17167_));
  OAI21_X1   g16911(.A1(new_n12203_), .A2(new_n2711_), .B(new_n17167_), .ZN(new_n17168_));
  XOR2_X1    g16912(.A1(new_n17168_), .A2(\a[26] ), .Z(new_n17169_));
  INV_X1     g16913(.I(new_n17169_), .ZN(new_n17170_));
  AOI22_X1   g16914(.A1(new_n3267_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n3270_), .ZN(new_n17171_));
  OAI21_X1   g16915(.A1(new_n9942_), .A2(new_n3475_), .B(new_n17171_), .ZN(new_n17172_));
  AOI21_X1   g16916(.A1(new_n10318_), .A2(new_n3273_), .B(new_n17172_), .ZN(new_n17173_));
  XOR2_X1    g16917(.A1(new_n17173_), .A2(new_n3264_), .Z(new_n17174_));
  INV_X1     g16918(.I(new_n17174_), .ZN(new_n17175_));
  INV_X1     g16919(.I(new_n17008_), .ZN(new_n17176_));
  AOI21_X1   g16920(.A1(new_n17176_), .A2(new_n17125_), .B(new_n17123_), .ZN(new_n17177_));
  OAI22_X1   g16921(.A1(new_n9032_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n9376_), .ZN(new_n17178_));
  AOI21_X1   g16922(.A1(\b[51] ), .A2(new_n4053_), .B(new_n17178_), .ZN(new_n17179_));
  OAI21_X1   g16923(.A1(new_n9385_), .A2(new_n4727_), .B(new_n17179_), .ZN(new_n17180_));
  XOR2_X1    g16924(.A1(new_n17180_), .A2(\a[32] ), .Z(new_n17181_));
  INV_X1     g16925(.I(new_n17181_), .ZN(new_n17182_));
  AOI22_X1   g16926(.A1(new_n4918_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n4921_), .ZN(new_n17183_));
  OAI21_X1   g16927(.A1(new_n8127_), .A2(new_n6099_), .B(new_n17183_), .ZN(new_n17184_));
  AOI21_X1   g16928(.A1(new_n9684_), .A2(new_n4699_), .B(new_n17184_), .ZN(new_n17185_));
  XOR2_X1    g16929(.A1(new_n17185_), .A2(new_n4446_), .Z(new_n17186_));
  AOI22_X1   g16930(.A1(new_n6108_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n6111_), .ZN(new_n17187_));
  OAI21_X1   g16931(.A1(new_n6490_), .A2(new_n7708_), .B(new_n17187_), .ZN(new_n17188_));
  AOI21_X1   g16932(.A1(new_n7906_), .A2(new_n6105_), .B(new_n17188_), .ZN(new_n17189_));
  XOR2_X1    g16933(.A1(new_n17189_), .A2(new_n5849_), .Z(new_n17190_));
  OAI21_X1   g16934(.A1(new_n17021_), .A2(new_n17092_), .B(new_n17094_), .ZN(new_n17191_));
  OAI22_X1   g16935(.A1(new_n7730_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n7731_), .ZN(new_n17192_));
  AOI21_X1   g16936(.A1(\b[39] ), .A2(new_n6887_), .B(new_n17192_), .ZN(new_n17193_));
  OAI21_X1   g16937(.A1(new_n6299_), .A2(new_n7728_), .B(new_n17193_), .ZN(new_n17194_));
  XOR2_X1    g16938(.A1(new_n17194_), .A2(\a[44] ), .Z(new_n17195_));
  AOI22_X1   g16939(.A1(new_n7403_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n7408_), .ZN(new_n17196_));
  OAI21_X1   g16940(.A1(new_n4886_), .A2(new_n9488_), .B(new_n17196_), .ZN(new_n17197_));
  AOI21_X1   g16941(.A1(new_n5351_), .A2(new_n7414_), .B(new_n17197_), .ZN(new_n17198_));
  XOR2_X1    g16942(.A1(new_n17198_), .A2(new_n7410_), .Z(new_n17199_));
  AOI21_X1   g16943(.A1(new_n17028_), .A2(new_n17079_), .B(new_n17077_), .ZN(new_n17200_));
  INV_X1     g16944(.I(new_n17200_), .ZN(new_n17201_));
  OAI22_X1   g16945(.A1(new_n9461_), .A2(new_n4666_), .B1(new_n4639_), .B2(new_n9462_), .ZN(new_n17202_));
  AOI21_X1   g16946(.A1(\b[33] ), .A2(new_n8575_), .B(new_n17202_), .ZN(new_n17203_));
  OAI21_X1   g16947(.A1(new_n4676_), .A2(new_n9460_), .B(new_n17203_), .ZN(new_n17204_));
  XOR2_X1    g16948(.A1(new_n17204_), .A2(new_n8248_), .Z(new_n17205_));
  AOI22_X1   g16949(.A1(new_n9125_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n9123_), .ZN(new_n17206_));
  OAI21_X1   g16950(.A1(new_n3624_), .A2(new_n9470_), .B(new_n17206_), .ZN(new_n17207_));
  AOI21_X1   g16951(.A1(new_n4030_), .A2(new_n9129_), .B(new_n17207_), .ZN(new_n17208_));
  XOR2_X1    g16952(.A1(new_n17208_), .A2(new_n9133_), .Z(new_n17209_));
  INV_X1     g16953(.I(new_n17209_), .ZN(new_n17210_));
  AOI22_X1   g16954(.A1(new_n10981_), .A2(\b[26] ), .B1(new_n10979_), .B2(\b[25] ), .ZN(new_n17211_));
  OAI21_X1   g16955(.A1(new_n2495_), .A2(new_n11306_), .B(new_n17211_), .ZN(new_n17212_));
  AOI21_X1   g16956(.A1(new_n3407_), .A2(new_n10984_), .B(new_n17212_), .ZN(new_n17213_));
  XOR2_X1    g16957(.A1(new_n17213_), .A2(new_n10989_), .Z(new_n17214_));
  AOI21_X1   g16958(.A1(new_n17038_), .A2(new_n17042_), .B(new_n17043_), .ZN(new_n17215_));
  INV_X1     g16959(.I(new_n17215_), .ZN(new_n17216_));
  AOI22_X1   g16960(.A1(new_n11926_), .A2(\b[23] ), .B1(new_n11924_), .B2(\b[22] ), .ZN(new_n17217_));
  OAI21_X1   g16961(.A1(new_n2027_), .A2(new_n12317_), .B(new_n17217_), .ZN(new_n17218_));
  AOI21_X1   g16962(.A1(new_n2470_), .A2(new_n11929_), .B(new_n17218_), .ZN(new_n17219_));
  XOR2_X1    g16963(.A1(new_n17219_), .A2(new_n12312_), .Z(new_n17220_));
  AOI22_X1   g16964(.A1(new_n12922_), .A2(\b[20] ), .B1(\b[19] ), .B2(new_n12923_), .ZN(new_n17221_));
  INV_X1     g16965(.I(new_n17221_), .ZN(new_n17222_));
  NOR2_X1    g16966(.A1(new_n17222_), .A2(new_n17041_), .ZN(new_n17223_));
  INV_X1     g16967(.I(new_n17223_), .ZN(new_n17224_));
  NAND2_X1   g16968(.A1(new_n17222_), .A2(new_n17041_), .ZN(new_n17225_));
  NAND2_X1   g16969(.A1(new_n17224_), .A2(new_n17225_), .ZN(new_n17226_));
  XOR2_X1    g16970(.A1(new_n17220_), .A2(new_n17226_), .Z(new_n17227_));
  NOR2_X1    g16971(.A1(new_n17227_), .A2(new_n17216_), .ZN(new_n17228_));
  INV_X1     g16972(.I(new_n17228_), .ZN(new_n17229_));
  NAND2_X1   g16973(.A1(new_n17227_), .A2(new_n17216_), .ZN(new_n17230_));
  NAND2_X1   g16974(.A1(new_n17229_), .A2(new_n17230_), .ZN(new_n17231_));
  XOR2_X1    g16975(.A1(new_n17231_), .A2(new_n17214_), .Z(new_n17232_));
  AOI22_X1   g16976(.A1(new_n10064_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n10062_), .ZN(new_n17233_));
  OAI21_X1   g16977(.A1(new_n3158_), .A2(new_n10399_), .B(new_n17233_), .ZN(new_n17234_));
  AOI21_X1   g16978(.A1(new_n4188_), .A2(new_n10068_), .B(new_n17234_), .ZN(new_n17235_));
  XOR2_X1    g16979(.A1(new_n17235_), .A2(new_n10057_), .Z(new_n17236_));
  AOI21_X1   g16980(.A1(new_n17046_), .A2(new_n17055_), .B(new_n17053_), .ZN(new_n17237_));
  NOR2_X1    g16981(.A1(new_n17236_), .A2(new_n17237_), .ZN(new_n17238_));
  INV_X1     g16982(.I(new_n17238_), .ZN(new_n17239_));
  NAND2_X1   g16983(.A1(new_n17236_), .A2(new_n17237_), .ZN(new_n17240_));
  NAND2_X1   g16984(.A1(new_n17239_), .A2(new_n17240_), .ZN(new_n17241_));
  XOR2_X1    g16985(.A1(new_n17241_), .A2(new_n17232_), .Z(new_n17242_));
  INV_X1     g16986(.I(new_n17032_), .ZN(new_n17243_));
  AOI21_X1   g16987(.A1(new_n17243_), .A2(new_n17060_), .B(new_n17058_), .ZN(new_n17244_));
  NOR2_X1    g16988(.A1(new_n17242_), .A2(new_n17244_), .ZN(new_n17245_));
  INV_X1     g16989(.I(new_n17245_), .ZN(new_n17246_));
  NAND2_X1   g16990(.A1(new_n17242_), .A2(new_n17244_), .ZN(new_n17247_));
  NAND2_X1   g16991(.A1(new_n17246_), .A2(new_n17247_), .ZN(new_n17248_));
  XOR2_X1    g16992(.A1(new_n17248_), .A2(new_n17210_), .Z(new_n17249_));
  AOI21_X1   g16993(.A1(new_n17062_), .A2(new_n17071_), .B(new_n17069_), .ZN(new_n17250_));
  NOR2_X1    g16994(.A1(new_n17249_), .A2(new_n17250_), .ZN(new_n17251_));
  INV_X1     g16995(.I(new_n17251_), .ZN(new_n17252_));
  NAND2_X1   g16996(.A1(new_n17249_), .A2(new_n17250_), .ZN(new_n17253_));
  NAND2_X1   g16997(.A1(new_n17252_), .A2(new_n17253_), .ZN(new_n17254_));
  XNOR2_X1   g16998(.A1(new_n17254_), .A2(new_n17205_), .ZN(new_n17255_));
  NOR2_X1    g16999(.A1(new_n17255_), .A2(new_n17201_), .ZN(new_n17256_));
  INV_X1     g17000(.I(new_n17256_), .ZN(new_n17257_));
  NAND2_X1   g17001(.A1(new_n17255_), .A2(new_n17201_), .ZN(new_n17258_));
  NAND2_X1   g17002(.A1(new_n17257_), .A2(new_n17258_), .ZN(new_n17259_));
  XOR2_X1    g17003(.A1(new_n17259_), .A2(new_n17199_), .Z(new_n17260_));
  INV_X1     g17004(.I(new_n17081_), .ZN(new_n17261_));
  AOI21_X1   g17005(.A1(new_n17261_), .A2(new_n17089_), .B(new_n17087_), .ZN(new_n17262_));
  XOR2_X1    g17006(.A1(new_n17260_), .A2(new_n17262_), .Z(new_n17263_));
  XOR2_X1    g17007(.A1(new_n17263_), .A2(new_n17195_), .Z(new_n17264_));
  NOR2_X1    g17008(.A1(new_n17264_), .A2(new_n17191_), .ZN(new_n17265_));
  INV_X1     g17009(.I(new_n17265_), .ZN(new_n17266_));
  NAND2_X1   g17010(.A1(new_n17264_), .A2(new_n17191_), .ZN(new_n17267_));
  NAND2_X1   g17011(.A1(new_n17266_), .A2(new_n17267_), .ZN(new_n17268_));
  XNOR2_X1   g17012(.A1(new_n17268_), .A2(new_n17190_), .ZN(new_n17269_));
  AOI22_X1   g17013(.A1(new_n5155_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n5160_), .ZN(new_n17270_));
  OAI21_X1   g17014(.A1(new_n7096_), .A2(new_n6877_), .B(new_n17270_), .ZN(new_n17271_));
  AOI21_X1   g17015(.A1(new_n7649_), .A2(new_n5166_), .B(new_n17271_), .ZN(new_n17272_));
  XOR2_X1    g17016(.A1(new_n17272_), .A2(new_n5162_), .Z(new_n17273_));
  NOR2_X1    g17017(.A1(new_n17104_), .A2(new_n17017_), .ZN(new_n17274_));
  NOR2_X1    g17018(.A1(new_n17274_), .A2(new_n17102_), .ZN(new_n17275_));
  NOR2_X1    g17019(.A1(new_n17275_), .A2(new_n17273_), .ZN(new_n17276_));
  AND2_X2    g17020(.A1(new_n17275_), .A2(new_n17273_), .Z(new_n17277_));
  NOR2_X1    g17021(.A1(new_n17277_), .A2(new_n17276_), .ZN(new_n17278_));
  XOR2_X1    g17022(.A1(new_n17269_), .A2(new_n17278_), .Z(new_n17279_));
  AOI21_X1   g17023(.A1(new_n17015_), .A2(new_n17110_), .B(new_n17108_), .ZN(new_n17280_));
  NOR2_X1    g17024(.A1(new_n17279_), .A2(new_n17280_), .ZN(new_n17281_));
  INV_X1     g17025(.I(new_n17281_), .ZN(new_n17282_));
  NAND2_X1   g17026(.A1(new_n17279_), .A2(new_n17280_), .ZN(new_n17283_));
  NAND2_X1   g17027(.A1(new_n17282_), .A2(new_n17283_), .ZN(new_n17284_));
  XOR2_X1    g17028(.A1(new_n17284_), .A2(new_n17186_), .Z(new_n17285_));
  INV_X1     g17029(.I(new_n17285_), .ZN(new_n17286_));
  NOR2_X1    g17030(.A1(new_n17120_), .A2(new_n17112_), .ZN(new_n17287_));
  NOR2_X1    g17031(.A1(new_n17287_), .A2(new_n17118_), .ZN(new_n17288_));
  NOR2_X1    g17032(.A1(new_n17286_), .A2(new_n17288_), .ZN(new_n17289_));
  INV_X1     g17033(.I(new_n17289_), .ZN(new_n17290_));
  NAND2_X1   g17034(.A1(new_n17286_), .A2(new_n17288_), .ZN(new_n17291_));
  NAND2_X1   g17035(.A1(new_n17290_), .A2(new_n17291_), .ZN(new_n17292_));
  XOR2_X1    g17036(.A1(new_n17292_), .A2(new_n17182_), .Z(new_n17293_));
  NOR2_X1    g17037(.A1(new_n17293_), .A2(new_n17177_), .ZN(new_n17294_));
  INV_X1     g17038(.I(new_n17294_), .ZN(new_n17295_));
  NAND2_X1   g17039(.A1(new_n17293_), .A2(new_n17177_), .ZN(new_n17296_));
  NAND2_X1   g17040(.A1(new_n17295_), .A2(new_n17296_), .ZN(new_n17297_));
  XOR2_X1    g17041(.A1(new_n17297_), .A2(new_n17175_), .Z(new_n17298_));
  OAI21_X1   g17042(.A1(new_n17002_), .A2(new_n17128_), .B(new_n17129_), .ZN(new_n17299_));
  INV_X1     g17043(.I(new_n17299_), .ZN(new_n17300_));
  OR2_X2     g17044(.A1(new_n17298_), .A2(new_n17300_), .Z(new_n17301_));
  NAND2_X1   g17045(.A1(new_n17298_), .A2(new_n17300_), .ZN(new_n17302_));
  NAND2_X1   g17046(.A1(new_n17301_), .A2(new_n17302_), .ZN(new_n17303_));
  XOR2_X1    g17047(.A1(new_n17303_), .A2(new_n17170_), .Z(new_n17304_));
  XOR2_X1    g17048(.A1(new_n17304_), .A2(new_n2200_), .Z(new_n17305_));
  AOI22_X1   g17049(.A1(new_n2202_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n2205_), .ZN(new_n17306_));
  OAI21_X1   g17050(.A1(new_n12147_), .A2(new_n2370_), .B(new_n17306_), .ZN(new_n17307_));
  AOI21_X1   g17051(.A1(new_n13444_), .A2(new_n2208_), .B(new_n17307_), .ZN(new_n17308_));
  INV_X1     g17052(.I(new_n16996_), .ZN(new_n17309_));
  AOI21_X1   g17053(.A1(new_n17309_), .A2(new_n17135_), .B(new_n17133_), .ZN(new_n17310_));
  XOR2_X1    g17054(.A1(new_n17310_), .A2(new_n17308_), .Z(new_n17311_));
  XOR2_X1    g17055(.A1(new_n17305_), .A2(new_n17311_), .Z(new_n17312_));
  AOI21_X1   g17056(.A1(new_n16991_), .A2(new_n17139_), .B(new_n17140_), .ZN(new_n17313_));
  INV_X1     g17057(.I(new_n17313_), .ZN(new_n17314_));
  XOR2_X1    g17058(.A1(new_n17312_), .A2(new_n17314_), .Z(new_n17315_));
  XNOR2_X1   g17059(.A1(new_n17315_), .A2(new_n17165_), .ZN(new_n17316_));
  INV_X1     g17060(.I(new_n17316_), .ZN(new_n17317_));
  NOR2_X1    g17061(.A1(new_n17317_), .A2(new_n17163_), .ZN(new_n17318_));
  INV_X1     g17062(.I(new_n17318_), .ZN(new_n17319_));
  NAND2_X1   g17063(.A1(new_n17317_), .A2(new_n17163_), .ZN(new_n17320_));
  NAND2_X1   g17064(.A1(new_n17319_), .A2(new_n17320_), .ZN(new_n17321_));
  XOR2_X1    g17065(.A1(new_n17162_), .A2(new_n17321_), .Z(\f[83] ));
  INV_X1     g17066(.I(new_n17320_), .ZN(new_n17323_));
  AOI21_X1   g17067(.A1(new_n17161_), .A2(new_n17159_), .B(new_n17318_), .ZN(new_n17324_));
  NOR2_X1    g17068(.A1(new_n17324_), .A2(new_n17323_), .ZN(new_n17325_));
  NOR2_X1    g17069(.A1(new_n17304_), .A2(new_n17310_), .ZN(new_n17326_));
  NAND2_X1   g17070(.A1(new_n17304_), .A2(new_n17310_), .ZN(new_n17327_));
  XOR2_X1    g17071(.A1(new_n17308_), .A2(new_n2200_), .Z(new_n17328_));
  INV_X1     g17072(.I(new_n17328_), .ZN(new_n17329_));
  AOI21_X1   g17073(.A1(new_n17327_), .A2(new_n17329_), .B(new_n17326_), .ZN(new_n17330_));
  INV_X1     g17074(.I(new_n17330_), .ZN(new_n17331_));
  AOI22_X1   g17075(.A1(new_n2202_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n2205_), .ZN(new_n17332_));
  OAI21_X1   g17076(.A1(new_n12148_), .A2(new_n2370_), .B(new_n17332_), .ZN(new_n17333_));
  AOI21_X1   g17077(.A1(new_n12811_), .A2(new_n2208_), .B(new_n17333_), .ZN(new_n17334_));
  XOR2_X1    g17078(.A1(new_n17334_), .A2(new_n2200_), .Z(new_n17335_));
  AOI22_X1   g17079(.A1(new_n2716_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n2719_), .ZN(new_n17336_));
  OAI21_X1   g17080(.A1(new_n11195_), .A2(new_n2924_), .B(new_n17336_), .ZN(new_n17337_));
  AOI21_X1   g17081(.A1(new_n11836_), .A2(new_n2722_), .B(new_n17337_), .ZN(new_n17338_));
  XOR2_X1    g17082(.A1(new_n17338_), .A2(new_n2714_), .Z(new_n17339_));
  INV_X1     g17083(.I(new_n17339_), .ZN(new_n17340_));
  NAND2_X1   g17084(.A1(new_n17302_), .A2(new_n17170_), .ZN(new_n17341_));
  NAND2_X1   g17085(.A1(new_n17341_), .A2(new_n17301_), .ZN(new_n17342_));
  INV_X1     g17086(.I(new_n17342_), .ZN(new_n17343_));
  AOI21_X1   g17087(.A1(new_n17175_), .A2(new_n17296_), .B(new_n17294_), .ZN(new_n17344_));
  AOI22_X1   g17088(.A1(new_n3267_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n3270_), .ZN(new_n17345_));
  OAI21_X1   g17089(.A1(new_n9972_), .A2(new_n3475_), .B(new_n17345_), .ZN(new_n17346_));
  AOI21_X1   g17090(.A1(new_n10631_), .A2(new_n3273_), .B(new_n17346_), .ZN(new_n17347_));
  XOR2_X1    g17091(.A1(new_n17347_), .A2(new_n3264_), .Z(new_n17348_));
  INV_X1     g17092(.I(new_n17348_), .ZN(new_n17349_));
  AOI22_X1   g17093(.A1(new_n3864_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n3869_), .ZN(new_n17350_));
  OAI21_X1   g17094(.A1(new_n9032_), .A2(new_n5410_), .B(new_n17350_), .ZN(new_n17351_));
  AOI21_X1   g17095(.A1(new_n10884_), .A2(new_n3872_), .B(new_n17351_), .ZN(new_n17352_));
  XOR2_X1    g17096(.A1(new_n17352_), .A2(new_n3876_), .Z(new_n17353_));
  NAND2_X1   g17097(.A1(new_n17291_), .A2(new_n17182_), .ZN(new_n17354_));
  NAND2_X1   g17098(.A1(new_n17354_), .A2(new_n17290_), .ZN(new_n17355_));
  INV_X1     g17099(.I(new_n17355_), .ZN(new_n17356_));
  INV_X1     g17100(.I(new_n17186_), .ZN(new_n17357_));
  AOI21_X1   g17101(.A1(new_n17357_), .A2(new_n17283_), .B(new_n17281_), .ZN(new_n17358_));
  INV_X1     g17102(.I(new_n17358_), .ZN(new_n17359_));
  OAI21_X1   g17103(.A1(new_n17190_), .A2(new_n17265_), .B(new_n17267_), .ZN(new_n17360_));
  OAI21_X1   g17104(.A1(new_n17199_), .A2(new_n17256_), .B(new_n17258_), .ZN(new_n17361_));
  AOI21_X1   g17105(.A1(new_n17205_), .A2(new_n17253_), .B(new_n17251_), .ZN(new_n17362_));
  INV_X1     g17106(.I(new_n17362_), .ZN(new_n17363_));
  AOI22_X1   g17107(.A1(new_n8241_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n8246_), .ZN(new_n17364_));
  OAI21_X1   g17108(.A1(new_n4639_), .A2(new_n9114_), .B(new_n17364_), .ZN(new_n17365_));
  AOI21_X1   g17109(.A1(new_n5594_), .A2(new_n8252_), .B(new_n17365_), .ZN(new_n17366_));
  XOR2_X1    g17110(.A1(new_n17366_), .A2(new_n8248_), .Z(new_n17367_));
  AOI21_X1   g17111(.A1(new_n17210_), .A2(new_n17247_), .B(new_n17245_), .ZN(new_n17368_));
  INV_X1     g17112(.I(new_n17368_), .ZN(new_n17369_));
  OAI21_X1   g17113(.A1(new_n17214_), .A2(new_n17228_), .B(new_n17230_), .ZN(new_n17370_));
  INV_X1     g17114(.I(new_n17370_), .ZN(new_n17371_));
  OAI22_X1   g17115(.A1(new_n12306_), .A2(new_n3158_), .B1(new_n12305_), .B2(new_n3006_), .ZN(new_n17372_));
  AOI21_X1   g17116(.A1(\b[25] ), .A2(new_n12304_), .B(new_n17372_), .ZN(new_n17373_));
  OAI21_X1   g17117(.A1(new_n3165_), .A2(new_n10985_), .B(new_n17373_), .ZN(new_n17374_));
  XOR2_X1    g17118(.A1(new_n17374_), .A2(new_n10989_), .Z(new_n17375_));
  AOI22_X1   g17119(.A1(new_n11926_), .A2(\b[24] ), .B1(new_n11924_), .B2(\b[23] ), .ZN(new_n17376_));
  OAI21_X1   g17120(.A1(new_n2142_), .A2(new_n12317_), .B(new_n17376_), .ZN(new_n17377_));
  AOI21_X1   g17121(.A1(new_n3033_), .A2(new_n11929_), .B(new_n17377_), .ZN(new_n17378_));
  XOR2_X1    g17122(.A1(new_n17378_), .A2(new_n12312_), .Z(new_n17379_));
  OAI21_X1   g17123(.A1(new_n17220_), .A2(new_n17223_), .B(new_n17225_), .ZN(new_n17380_));
  AOI22_X1   g17124(.A1(new_n12922_), .A2(\b[21] ), .B1(\b[20] ), .B2(new_n12923_), .ZN(new_n17381_));
  INV_X1     g17125(.I(new_n17381_), .ZN(new_n17382_));
  NOR2_X1    g17126(.A1(new_n17382_), .A2(new_n1736_), .ZN(new_n17383_));
  NOR2_X1    g17127(.A1(new_n17381_), .A2(\a[20] ), .ZN(new_n17384_));
  NOR2_X1    g17128(.A1(new_n17383_), .A2(new_n17384_), .ZN(new_n17385_));
  XOR2_X1    g17129(.A1(new_n17385_), .A2(new_n17221_), .Z(new_n17386_));
  NOR2_X1    g17130(.A1(new_n17380_), .A2(new_n17386_), .ZN(new_n17387_));
  INV_X1     g17131(.I(new_n17387_), .ZN(new_n17388_));
  NAND2_X1   g17132(.A1(new_n17380_), .A2(new_n17386_), .ZN(new_n17389_));
  NAND2_X1   g17133(.A1(new_n17388_), .A2(new_n17389_), .ZN(new_n17390_));
  XOR2_X1    g17134(.A1(new_n17390_), .A2(new_n17379_), .Z(new_n17391_));
  NAND2_X1   g17135(.A1(new_n17375_), .A2(new_n17391_), .ZN(new_n17392_));
  NOR2_X1    g17136(.A1(new_n17375_), .A2(new_n17391_), .ZN(new_n17393_));
  INV_X1     g17137(.I(new_n17393_), .ZN(new_n17394_));
  NAND2_X1   g17138(.A1(new_n17394_), .A2(new_n17392_), .ZN(new_n17395_));
  XOR2_X1    g17139(.A1(new_n17395_), .A2(new_n17371_), .Z(new_n17396_));
  AOI22_X1   g17140(.A1(new_n10064_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n10062_), .ZN(new_n17397_));
  OAI21_X1   g17141(.A1(new_n3185_), .A2(new_n10399_), .B(new_n17397_), .ZN(new_n17398_));
  AOI21_X1   g17142(.A1(new_n4230_), .A2(new_n10068_), .B(new_n17398_), .ZN(new_n17399_));
  XOR2_X1    g17143(.A1(new_n17399_), .A2(new_n10057_), .Z(new_n17400_));
  INV_X1     g17144(.I(new_n17400_), .ZN(new_n17401_));
  NAND2_X1   g17145(.A1(new_n17240_), .A2(new_n17232_), .ZN(new_n17402_));
  NAND2_X1   g17146(.A1(new_n17402_), .A2(new_n17239_), .ZN(new_n17403_));
  NAND2_X1   g17147(.A1(new_n17403_), .A2(new_n17401_), .ZN(new_n17404_));
  NAND3_X1   g17148(.A1(new_n17402_), .A2(new_n17239_), .A3(new_n17400_), .ZN(new_n17405_));
  NAND2_X1   g17149(.A1(new_n17404_), .A2(new_n17405_), .ZN(new_n17406_));
  XNOR2_X1   g17150(.A1(new_n17406_), .A2(new_n17396_), .ZN(new_n17407_));
  INV_X1     g17151(.I(new_n17407_), .ZN(new_n17408_));
  AOI22_X1   g17152(.A1(new_n9125_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n9123_), .ZN(new_n17409_));
  OAI21_X1   g17153(.A1(new_n4022_), .A2(new_n9470_), .B(new_n17409_), .ZN(new_n17410_));
  AOI21_X1   g17154(.A1(new_n4223_), .A2(new_n9129_), .B(new_n17410_), .ZN(new_n17411_));
  XOR2_X1    g17155(.A1(new_n17411_), .A2(new_n9133_), .Z(new_n17412_));
  NOR2_X1    g17156(.A1(new_n17408_), .A2(new_n17412_), .ZN(new_n17413_));
  INV_X1     g17157(.I(new_n17413_), .ZN(new_n17414_));
  NAND2_X1   g17158(.A1(new_n17408_), .A2(new_n17412_), .ZN(new_n17415_));
  NAND2_X1   g17159(.A1(new_n17414_), .A2(new_n17415_), .ZN(new_n17416_));
  XOR2_X1    g17160(.A1(new_n17416_), .A2(new_n17369_), .Z(new_n17417_));
  NOR2_X1    g17161(.A1(new_n17417_), .A2(new_n17367_), .ZN(new_n17418_));
  NAND2_X1   g17162(.A1(new_n17417_), .A2(new_n17367_), .ZN(new_n17419_));
  INV_X1     g17163(.I(new_n17419_), .ZN(new_n17420_));
  NOR2_X1    g17164(.A1(new_n17420_), .A2(new_n17418_), .ZN(new_n17421_));
  XOR2_X1    g17165(.A1(new_n17421_), .A2(new_n17363_), .Z(new_n17422_));
  INV_X1     g17166(.I(new_n17422_), .ZN(new_n17423_));
  AOI22_X1   g17167(.A1(new_n7403_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n7408_), .ZN(new_n17424_));
  OAI21_X1   g17168(.A1(new_n5312_), .A2(new_n9488_), .B(new_n17424_), .ZN(new_n17425_));
  AOI21_X1   g17169(.A1(new_n6310_), .A2(new_n7414_), .B(new_n17425_), .ZN(new_n17426_));
  XOR2_X1    g17170(.A1(new_n17426_), .A2(new_n7410_), .Z(new_n17427_));
  NOR2_X1    g17171(.A1(new_n17423_), .A2(new_n17427_), .ZN(new_n17428_));
  NAND2_X1   g17172(.A1(new_n17423_), .A2(new_n17427_), .ZN(new_n17429_));
  INV_X1     g17173(.I(new_n17429_), .ZN(new_n17430_));
  NOR2_X1    g17174(.A1(new_n17430_), .A2(new_n17428_), .ZN(new_n17431_));
  XOR2_X1    g17175(.A1(new_n17431_), .A2(new_n17361_), .Z(new_n17432_));
  AOI22_X1   g17176(.A1(new_n6569_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n6574_), .ZN(new_n17433_));
  OAI21_X1   g17177(.A1(new_n6284_), .A2(new_n8565_), .B(new_n17433_), .ZN(new_n17434_));
  AOI21_X1   g17178(.A1(new_n7106_), .A2(new_n6579_), .B(new_n17434_), .ZN(new_n17435_));
  XOR2_X1    g17179(.A1(new_n17435_), .A2(new_n6567_), .Z(new_n17436_));
  INV_X1     g17180(.I(new_n17260_), .ZN(new_n17437_));
  NOR2_X1    g17181(.A1(new_n17437_), .A2(new_n17262_), .ZN(new_n17438_));
  AOI21_X1   g17182(.A1(new_n17437_), .A2(new_n17262_), .B(new_n17195_), .ZN(new_n17439_));
  NOR2_X1    g17183(.A1(new_n17439_), .A2(new_n17438_), .ZN(new_n17440_));
  NOR2_X1    g17184(.A1(new_n17440_), .A2(new_n17436_), .ZN(new_n17441_));
  NAND2_X1   g17185(.A1(new_n17440_), .A2(new_n17436_), .ZN(new_n17442_));
  INV_X1     g17186(.I(new_n17442_), .ZN(new_n17443_));
  NOR2_X1    g17187(.A1(new_n17443_), .A2(new_n17441_), .ZN(new_n17444_));
  XOR2_X1    g17188(.A1(new_n17444_), .A2(new_n17432_), .Z(new_n17445_));
  AOI22_X1   g17189(.A1(new_n6108_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n6111_), .ZN(new_n17446_));
  OAI21_X1   g17190(.A1(new_n6775_), .A2(new_n7708_), .B(new_n17446_), .ZN(new_n17447_));
  AOI21_X1   g17191(.A1(new_n7926_), .A2(new_n6105_), .B(new_n17447_), .ZN(new_n17448_));
  XOR2_X1    g17192(.A1(new_n17448_), .A2(\a[41] ), .Z(new_n17449_));
  NAND2_X1   g17193(.A1(new_n17445_), .A2(new_n17449_), .ZN(new_n17450_));
  OR2_X2     g17194(.A1(new_n17445_), .A2(new_n17449_), .Z(new_n17451_));
  NAND2_X1   g17195(.A1(new_n17451_), .A2(new_n17450_), .ZN(new_n17452_));
  XNOR2_X1   g17196(.A1(new_n17452_), .A2(new_n17360_), .ZN(new_n17453_));
  AOI22_X1   g17197(.A1(new_n5155_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n5160_), .ZN(new_n17454_));
  OAI21_X1   g17198(.A1(new_n7617_), .A2(new_n6877_), .B(new_n17454_), .ZN(new_n17455_));
  AOI21_X1   g17199(.A1(new_n8792_), .A2(new_n5166_), .B(new_n17455_), .ZN(new_n17456_));
  XOR2_X1    g17200(.A1(new_n17456_), .A2(\a[38] ), .Z(new_n17457_));
  INV_X1     g17201(.I(new_n17276_), .ZN(new_n17458_));
  OAI21_X1   g17202(.A1(new_n17269_), .A2(new_n17277_), .B(new_n17458_), .ZN(new_n17459_));
  NAND2_X1   g17203(.A1(new_n17459_), .A2(new_n17457_), .ZN(new_n17460_));
  OR2_X2     g17204(.A1(new_n17459_), .A2(new_n17457_), .Z(new_n17461_));
  NAND2_X1   g17205(.A1(new_n17461_), .A2(new_n17460_), .ZN(new_n17462_));
  XNOR2_X1   g17206(.A1(new_n17462_), .A2(new_n17453_), .ZN(new_n17463_));
  INV_X1     g17207(.I(new_n17463_), .ZN(new_n17464_));
  AOI22_X1   g17208(.A1(new_n4918_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n4921_), .ZN(new_n17465_));
  OAI21_X1   g17209(.A1(new_n8168_), .A2(new_n6099_), .B(new_n17465_), .ZN(new_n17466_));
  AOI21_X1   g17210(.A1(new_n8783_), .A2(new_n4699_), .B(new_n17466_), .ZN(new_n17467_));
  XOR2_X1    g17211(.A1(new_n17467_), .A2(new_n4446_), .Z(new_n17468_));
  NOR2_X1    g17212(.A1(new_n17464_), .A2(new_n17468_), .ZN(new_n17469_));
  INV_X1     g17213(.I(new_n17469_), .ZN(new_n17470_));
  NAND2_X1   g17214(.A1(new_n17464_), .A2(new_n17468_), .ZN(new_n17471_));
  NAND2_X1   g17215(.A1(new_n17470_), .A2(new_n17471_), .ZN(new_n17472_));
  XOR2_X1    g17216(.A1(new_n17472_), .A2(new_n17359_), .Z(new_n17473_));
  NOR2_X1    g17217(.A1(new_n17473_), .A2(new_n17356_), .ZN(new_n17474_));
  INV_X1     g17218(.I(new_n17474_), .ZN(new_n17475_));
  NAND2_X1   g17219(.A1(new_n17473_), .A2(new_n17356_), .ZN(new_n17476_));
  NAND2_X1   g17220(.A1(new_n17475_), .A2(new_n17476_), .ZN(new_n17477_));
  XOR2_X1    g17221(.A1(new_n17477_), .A2(new_n17353_), .Z(new_n17478_));
  NOR2_X1    g17222(.A1(new_n17478_), .A2(new_n17349_), .ZN(new_n17479_));
  NAND2_X1   g17223(.A1(new_n17478_), .A2(new_n17349_), .ZN(new_n17480_));
  INV_X1     g17224(.I(new_n17480_), .ZN(new_n17481_));
  NOR2_X1    g17225(.A1(new_n17481_), .A2(new_n17479_), .ZN(new_n17482_));
  XOR2_X1    g17226(.A1(new_n17482_), .A2(new_n17344_), .Z(new_n17483_));
  NOR2_X1    g17227(.A1(new_n17483_), .A2(new_n17343_), .ZN(new_n17484_));
  INV_X1     g17228(.I(new_n17484_), .ZN(new_n17485_));
  NAND2_X1   g17229(.A1(new_n17483_), .A2(new_n17343_), .ZN(new_n17486_));
  NAND2_X1   g17230(.A1(new_n17485_), .A2(new_n17486_), .ZN(new_n17487_));
  XOR2_X1    g17231(.A1(new_n17487_), .A2(new_n17340_), .Z(new_n17488_));
  NAND2_X1   g17232(.A1(new_n17488_), .A2(new_n17335_), .ZN(new_n17489_));
  NOR2_X1    g17233(.A1(new_n17488_), .A2(new_n17335_), .ZN(new_n17490_));
  INV_X1     g17234(.I(new_n17490_), .ZN(new_n17491_));
  NAND2_X1   g17235(.A1(new_n17491_), .A2(new_n17489_), .ZN(new_n17492_));
  XOR2_X1    g17236(.A1(new_n17492_), .A2(new_n17331_), .Z(new_n17493_));
  INV_X1     g17237(.I(new_n17493_), .ZN(new_n17494_));
  INV_X1     g17238(.I(new_n17312_), .ZN(new_n17495_));
  NAND2_X1   g17239(.A1(new_n17495_), .A2(new_n17314_), .ZN(new_n17496_));
  NOR2_X1    g17240(.A1(new_n17495_), .A2(new_n17314_), .ZN(new_n17497_));
  OAI21_X1   g17241(.A1(new_n17165_), .A2(new_n17497_), .B(new_n17496_), .ZN(new_n17498_));
  NOR2_X1    g17242(.A1(new_n17494_), .A2(new_n17498_), .ZN(new_n17499_));
  INV_X1     g17243(.I(new_n17499_), .ZN(new_n17500_));
  NAND2_X1   g17244(.A1(new_n17494_), .A2(new_n17498_), .ZN(new_n17501_));
  AND2_X2    g17245(.A1(new_n17500_), .A2(new_n17501_), .Z(new_n17502_));
  XOR2_X1    g17246(.A1(new_n17325_), .A2(new_n17502_), .Z(\f[84] ));
  OAI22_X1   g17247(.A1(new_n2370_), .A2(new_n12796_), .B1(new_n12800_), .B2(new_n2194_), .ZN(new_n17504_));
  AOI21_X1   g17248(.A1(new_n13973_), .A2(new_n2208_), .B(new_n17504_), .ZN(new_n17505_));
  XOR2_X1    g17249(.A1(new_n17505_), .A2(new_n2200_), .Z(new_n17506_));
  INV_X1     g17250(.I(new_n17506_), .ZN(new_n17507_));
  AOI21_X1   g17251(.A1(new_n17340_), .A2(new_n17486_), .B(new_n17484_), .ZN(new_n17508_));
  INV_X1     g17252(.I(new_n17508_), .ZN(new_n17509_));
  OAI22_X1   g17253(.A1(new_n2703_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n2708_), .ZN(new_n17510_));
  AOI21_X1   g17254(.A1(\b[59] ), .A2(new_n2906_), .B(new_n17510_), .ZN(new_n17511_));
  OAI21_X1   g17255(.A1(new_n13110_), .A2(new_n2711_), .B(new_n17511_), .ZN(new_n17512_));
  XOR2_X1    g17256(.A1(new_n17512_), .A2(new_n2714_), .Z(new_n17513_));
  OAI21_X1   g17257(.A1(new_n17344_), .A2(new_n17479_), .B(new_n17480_), .ZN(new_n17514_));
  INV_X1     g17258(.I(new_n17514_), .ZN(new_n17515_));
  AOI22_X1   g17259(.A1(new_n3267_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n3270_), .ZN(new_n17516_));
  OAI21_X1   g17260(.A1(new_n10308_), .A2(new_n3475_), .B(new_n17516_), .ZN(new_n17517_));
  AOI21_X1   g17261(.A1(new_n12164_), .A2(new_n3273_), .B(new_n17517_), .ZN(new_n17518_));
  XOR2_X1    g17262(.A1(new_n17518_), .A2(new_n3264_), .Z(new_n17519_));
  INV_X1     g17263(.I(new_n17353_), .ZN(new_n17520_));
  AOI21_X1   g17264(.A1(new_n17520_), .A2(new_n17476_), .B(new_n17474_), .ZN(new_n17521_));
  INV_X1     g17265(.I(new_n17521_), .ZN(new_n17522_));
  AOI21_X1   g17266(.A1(new_n17359_), .A2(new_n17471_), .B(new_n17469_), .ZN(new_n17523_));
  AOI22_X1   g17267(.A1(new_n3864_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n3869_), .ZN(new_n17524_));
  OAI21_X1   g17268(.A1(new_n9376_), .A2(new_n5410_), .B(new_n17524_), .ZN(new_n17525_));
  AOI21_X1   g17269(.A1(new_n9979_), .A2(new_n3872_), .B(new_n17525_), .ZN(new_n17526_));
  XOR2_X1    g17270(.A1(new_n17526_), .A2(new_n3876_), .Z(new_n17527_));
  AOI22_X1   g17271(.A1(new_n4918_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n4921_), .ZN(new_n17528_));
  OAI21_X1   g17272(.A1(new_n8500_), .A2(new_n6099_), .B(new_n17528_), .ZN(new_n17529_));
  AOI21_X1   g17273(.A1(new_n9987_), .A2(new_n4699_), .B(new_n17529_), .ZN(new_n17530_));
  XOR2_X1    g17274(.A1(new_n17530_), .A2(new_n4446_), .Z(new_n17531_));
  AOI22_X1   g17275(.A1(new_n6108_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n6111_), .ZN(new_n17532_));
  OAI21_X1   g17276(.A1(new_n7074_), .A2(new_n7708_), .B(new_n17532_), .ZN(new_n17533_));
  AOI21_X1   g17277(.A1(new_n9337_), .A2(new_n6105_), .B(new_n17533_), .ZN(new_n17534_));
  XOR2_X1    g17278(.A1(new_n17534_), .A2(new_n5849_), .Z(new_n17535_));
  INV_X1     g17279(.I(new_n17535_), .ZN(new_n17536_));
  AOI21_X1   g17280(.A1(new_n17361_), .A2(new_n17429_), .B(new_n17428_), .ZN(new_n17537_));
  AOI22_X1   g17281(.A1(new_n7403_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n7408_), .ZN(new_n17538_));
  OAI21_X1   g17282(.A1(new_n5341_), .A2(new_n9488_), .B(new_n17538_), .ZN(new_n17539_));
  AOI21_X1   g17283(.A1(new_n5793_), .A2(new_n7414_), .B(new_n17539_), .ZN(new_n17540_));
  XOR2_X1    g17284(.A1(new_n17540_), .A2(new_n7410_), .Z(new_n17541_));
  AOI21_X1   g17285(.A1(new_n17363_), .A2(new_n17419_), .B(new_n17418_), .ZN(new_n17542_));
  INV_X1     g17286(.I(new_n17542_), .ZN(new_n17543_));
  AOI22_X1   g17287(.A1(new_n9125_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n9123_), .ZN(new_n17544_));
  OAI21_X1   g17288(.A1(new_n4023_), .A2(new_n9470_), .B(new_n17544_), .ZN(new_n17545_));
  AOI21_X1   g17289(.A1(new_n5103_), .A2(new_n9129_), .B(new_n17545_), .ZN(new_n17546_));
  XOR2_X1    g17290(.A1(new_n17546_), .A2(new_n9133_), .Z(new_n17547_));
  INV_X1     g17291(.I(new_n17547_), .ZN(new_n17548_));
  OAI21_X1   g17292(.A1(new_n17371_), .A2(new_n17393_), .B(new_n17392_), .ZN(new_n17549_));
  AOI22_X1   g17293(.A1(new_n10981_), .A2(\b[28] ), .B1(new_n10979_), .B2(\b[27] ), .ZN(new_n17550_));
  OAI21_X1   g17294(.A1(new_n3006_), .A2(new_n11306_), .B(new_n17550_), .ZN(new_n17551_));
  AOI21_X1   g17295(.A1(new_n3807_), .A2(new_n10984_), .B(new_n17551_), .ZN(new_n17552_));
  XOR2_X1    g17296(.A1(new_n17552_), .A2(new_n10989_), .Z(new_n17553_));
  OAI21_X1   g17297(.A1(new_n17379_), .A2(new_n17387_), .B(new_n17389_), .ZN(new_n17554_));
  OAI22_X1   g17298(.A1(new_n13224_), .A2(new_n2646_), .B1(new_n2495_), .B2(new_n11923_), .ZN(new_n17555_));
  AOI21_X1   g17299(.A1(\b[23] ), .A2(new_n13223_), .B(new_n17555_), .ZN(new_n17556_));
  OAI21_X1   g17300(.A1(new_n2655_), .A2(new_n11930_), .B(new_n17556_), .ZN(new_n17557_));
  XOR2_X1    g17301(.A1(new_n17557_), .A2(new_n12312_), .Z(new_n17558_));
  NOR2_X1    g17302(.A1(new_n17384_), .A2(new_n17222_), .ZN(new_n17559_));
  NOR2_X1    g17303(.A1(new_n17559_), .A2(new_n17383_), .ZN(new_n17560_));
  AOI22_X1   g17304(.A1(new_n12922_), .A2(\b[22] ), .B1(\b[21] ), .B2(new_n12923_), .ZN(new_n17561_));
  NAND2_X1   g17305(.A1(new_n17560_), .A2(new_n17561_), .ZN(new_n17562_));
  NOR2_X1    g17306(.A1(new_n17560_), .A2(new_n17561_), .ZN(new_n17563_));
  INV_X1     g17307(.I(new_n17563_), .ZN(new_n17564_));
  NAND2_X1   g17308(.A1(new_n17564_), .A2(new_n17562_), .ZN(new_n17565_));
  XNOR2_X1   g17309(.A1(new_n17558_), .A2(new_n17565_), .ZN(new_n17566_));
  NOR2_X1    g17310(.A1(new_n17566_), .A2(new_n17554_), .ZN(new_n17567_));
  INV_X1     g17311(.I(new_n17567_), .ZN(new_n17568_));
  NAND2_X1   g17312(.A1(new_n17566_), .A2(new_n17554_), .ZN(new_n17569_));
  NAND2_X1   g17313(.A1(new_n17568_), .A2(new_n17569_), .ZN(new_n17570_));
  XOR2_X1    g17314(.A1(new_n17570_), .A2(new_n17553_), .Z(new_n17571_));
  INV_X1     g17315(.I(new_n17571_), .ZN(new_n17572_));
  AOI22_X1   g17316(.A1(new_n10064_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n10062_), .ZN(new_n17573_));
  OAI21_X1   g17317(.A1(new_n3592_), .A2(new_n10399_), .B(new_n17573_), .ZN(new_n17574_));
  AOI21_X1   g17318(.A1(new_n3796_), .A2(new_n10068_), .B(new_n17574_), .ZN(new_n17575_));
  XOR2_X1    g17319(.A1(new_n17575_), .A2(new_n10057_), .Z(new_n17576_));
  NOR2_X1    g17320(.A1(new_n17576_), .A2(new_n17572_), .ZN(new_n17577_));
  NAND2_X1   g17321(.A1(new_n17576_), .A2(new_n17572_), .ZN(new_n17578_));
  INV_X1     g17322(.I(new_n17578_), .ZN(new_n17579_));
  NOR2_X1    g17323(.A1(new_n17579_), .A2(new_n17577_), .ZN(new_n17580_));
  XNOR2_X1   g17324(.A1(new_n17580_), .A2(new_n17549_), .ZN(new_n17581_));
  NAND2_X1   g17325(.A1(new_n17396_), .A2(new_n17405_), .ZN(new_n17582_));
  NAND2_X1   g17326(.A1(new_n17582_), .A2(new_n17404_), .ZN(new_n17583_));
  INV_X1     g17327(.I(new_n17583_), .ZN(new_n17584_));
  NOR2_X1    g17328(.A1(new_n17581_), .A2(new_n17584_), .ZN(new_n17585_));
  INV_X1     g17329(.I(new_n17585_), .ZN(new_n17586_));
  NAND2_X1   g17330(.A1(new_n17581_), .A2(new_n17584_), .ZN(new_n17587_));
  NAND2_X1   g17331(.A1(new_n17586_), .A2(new_n17587_), .ZN(new_n17588_));
  XOR2_X1    g17332(.A1(new_n17588_), .A2(new_n17548_), .Z(new_n17589_));
  AOI21_X1   g17333(.A1(new_n17369_), .A2(new_n17415_), .B(new_n17413_), .ZN(new_n17590_));
  OAI22_X1   g17334(.A1(new_n9461_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n9462_), .ZN(new_n17591_));
  AOI21_X1   g17335(.A1(\b[35] ), .A2(new_n8575_), .B(new_n17591_), .ZN(new_n17592_));
  OAI21_X1   g17336(.A1(new_n5322_), .A2(new_n9460_), .B(new_n17592_), .ZN(new_n17593_));
  XOR2_X1    g17337(.A1(new_n17593_), .A2(\a[50] ), .Z(new_n17594_));
  NOR2_X1    g17338(.A1(new_n17594_), .A2(new_n17590_), .ZN(new_n17595_));
  INV_X1     g17339(.I(new_n17595_), .ZN(new_n17596_));
  NAND2_X1   g17340(.A1(new_n17594_), .A2(new_n17590_), .ZN(new_n17597_));
  NAND2_X1   g17341(.A1(new_n17596_), .A2(new_n17597_), .ZN(new_n17598_));
  XOR2_X1    g17342(.A1(new_n17589_), .A2(new_n17598_), .Z(new_n17599_));
  NOR2_X1    g17343(.A1(new_n17599_), .A2(new_n17543_), .ZN(new_n17600_));
  INV_X1     g17344(.I(new_n17600_), .ZN(new_n17601_));
  NAND2_X1   g17345(.A1(new_n17599_), .A2(new_n17543_), .ZN(new_n17602_));
  NAND2_X1   g17346(.A1(new_n17601_), .A2(new_n17602_), .ZN(new_n17603_));
  XOR2_X1    g17347(.A1(new_n17603_), .A2(new_n17541_), .Z(new_n17604_));
  INV_X1     g17348(.I(new_n17604_), .ZN(new_n17605_));
  OAI22_X1   g17349(.A1(new_n7730_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n7731_), .ZN(new_n17606_));
  AOI21_X1   g17350(.A1(\b[41] ), .A2(new_n6887_), .B(new_n17606_), .ZN(new_n17607_));
  OAI21_X1   g17351(.A1(new_n6785_), .A2(new_n7728_), .B(new_n17607_), .ZN(new_n17608_));
  XOR2_X1    g17352(.A1(new_n17608_), .A2(\a[44] ), .Z(new_n17609_));
  NOR2_X1    g17353(.A1(new_n17605_), .A2(new_n17609_), .ZN(new_n17610_));
  NAND2_X1   g17354(.A1(new_n17605_), .A2(new_n17609_), .ZN(new_n17611_));
  INV_X1     g17355(.I(new_n17611_), .ZN(new_n17612_));
  NOR2_X1    g17356(.A1(new_n17612_), .A2(new_n17610_), .ZN(new_n17613_));
  XOR2_X1    g17357(.A1(new_n17613_), .A2(new_n17537_), .Z(new_n17614_));
  AOI21_X1   g17358(.A1(new_n17432_), .A2(new_n17442_), .B(new_n17441_), .ZN(new_n17615_));
  NOR2_X1    g17359(.A1(new_n17614_), .A2(new_n17615_), .ZN(new_n17616_));
  INV_X1     g17360(.I(new_n17616_), .ZN(new_n17617_));
  NAND2_X1   g17361(.A1(new_n17614_), .A2(new_n17615_), .ZN(new_n17618_));
  NAND2_X1   g17362(.A1(new_n17617_), .A2(new_n17618_), .ZN(new_n17619_));
  XOR2_X1    g17363(.A1(new_n17619_), .A2(new_n17536_), .Z(new_n17620_));
  INV_X1     g17364(.I(new_n17620_), .ZN(new_n17621_));
  INV_X1     g17365(.I(new_n17450_), .ZN(new_n17622_));
  AOI21_X1   g17366(.A1(new_n17360_), .A2(new_n17451_), .B(new_n17622_), .ZN(new_n17623_));
  OAI22_X1   g17367(.A1(new_n8168_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n8127_), .ZN(new_n17624_));
  AOI21_X1   g17368(.A1(\b[47] ), .A2(new_n5420_), .B(new_n17624_), .ZN(new_n17625_));
  OAI21_X1   g17369(.A1(new_n9050_), .A2(new_n6124_), .B(new_n17625_), .ZN(new_n17626_));
  XOR2_X1    g17370(.A1(new_n17626_), .A2(\a[38] ), .Z(new_n17627_));
  NOR2_X1    g17371(.A1(new_n17623_), .A2(new_n17627_), .ZN(new_n17628_));
  INV_X1     g17372(.I(new_n17628_), .ZN(new_n17629_));
  NAND2_X1   g17373(.A1(new_n17623_), .A2(new_n17627_), .ZN(new_n17630_));
  NAND2_X1   g17374(.A1(new_n17629_), .A2(new_n17630_), .ZN(new_n17631_));
  XOR2_X1    g17375(.A1(new_n17631_), .A2(new_n17621_), .Z(new_n17632_));
  NAND2_X1   g17376(.A1(new_n17453_), .A2(new_n17461_), .ZN(new_n17633_));
  AND2_X2    g17377(.A1(new_n17633_), .A2(new_n17460_), .Z(new_n17634_));
  XOR2_X1    g17378(.A1(new_n17632_), .A2(new_n17634_), .Z(new_n17635_));
  XOR2_X1    g17379(.A1(new_n17635_), .A2(new_n17531_), .Z(new_n17636_));
  NOR2_X1    g17380(.A1(new_n17636_), .A2(new_n17527_), .ZN(new_n17637_));
  NAND2_X1   g17381(.A1(new_n17636_), .A2(new_n17527_), .ZN(new_n17638_));
  INV_X1     g17382(.I(new_n17638_), .ZN(new_n17639_));
  NOR2_X1    g17383(.A1(new_n17639_), .A2(new_n17637_), .ZN(new_n17640_));
  XNOR2_X1   g17384(.A1(new_n17640_), .A2(new_n17523_), .ZN(new_n17641_));
  NOR2_X1    g17385(.A1(new_n17641_), .A2(new_n17522_), .ZN(new_n17642_));
  NAND2_X1   g17386(.A1(new_n17641_), .A2(new_n17522_), .ZN(new_n17643_));
  INV_X1     g17387(.I(new_n17643_), .ZN(new_n17644_));
  NOR2_X1    g17388(.A1(new_n17644_), .A2(new_n17642_), .ZN(new_n17645_));
  XOR2_X1    g17389(.A1(new_n17645_), .A2(new_n17519_), .Z(new_n17646_));
  OR2_X2     g17390(.A1(new_n17646_), .A2(new_n17515_), .Z(new_n17647_));
  NAND2_X1   g17391(.A1(new_n17646_), .A2(new_n17515_), .ZN(new_n17648_));
  NAND2_X1   g17392(.A1(new_n17647_), .A2(new_n17648_), .ZN(new_n17649_));
  XNOR2_X1   g17393(.A1(new_n17649_), .A2(new_n17513_), .ZN(new_n17650_));
  NOR2_X1    g17394(.A1(new_n17650_), .A2(new_n17509_), .ZN(new_n17651_));
  INV_X1     g17395(.I(new_n17651_), .ZN(new_n17652_));
  NAND2_X1   g17396(.A1(new_n17650_), .A2(new_n17509_), .ZN(new_n17653_));
  NAND2_X1   g17397(.A1(new_n17652_), .A2(new_n17653_), .ZN(new_n17654_));
  XOR2_X1    g17398(.A1(new_n17654_), .A2(new_n17507_), .Z(new_n17655_));
  INV_X1     g17399(.I(new_n17655_), .ZN(new_n17656_));
  AOI21_X1   g17400(.A1(new_n17331_), .A2(new_n17489_), .B(new_n17490_), .ZN(new_n17657_));
  INV_X1     g17401(.I(new_n17502_), .ZN(new_n17658_));
  NOR3_X1    g17402(.A1(new_n17324_), .A2(new_n17323_), .A3(new_n17658_), .ZN(new_n17659_));
  OAI21_X1   g17403(.A1(new_n17659_), .A2(new_n17499_), .B(new_n17657_), .ZN(new_n17660_));
  INV_X1     g17404(.I(new_n17657_), .ZN(new_n17661_));
  AOI21_X1   g17405(.A1(new_n17155_), .A2(new_n17151_), .B(new_n16981_), .ZN(new_n17662_));
  OAI21_X1   g17406(.A1(new_n17662_), .A2(new_n17156_), .B(new_n17319_), .ZN(new_n17663_));
  NAND3_X1   g17407(.A1(new_n17663_), .A2(new_n17320_), .A3(new_n17502_), .ZN(new_n17664_));
  NAND3_X1   g17408(.A1(new_n17664_), .A2(new_n17500_), .A3(new_n17661_), .ZN(new_n17665_));
  NAND2_X1   g17409(.A1(new_n17665_), .A2(new_n17660_), .ZN(new_n17666_));
  XOR2_X1    g17410(.A1(new_n17666_), .A2(new_n17656_), .Z(\f[85] ));
  NOR3_X1    g17411(.A1(new_n17659_), .A2(new_n17499_), .A3(new_n17657_), .ZN(new_n17668_));
  AOI21_X1   g17412(.A1(new_n17656_), .A2(new_n17660_), .B(new_n17668_), .ZN(new_n17669_));
  OAI21_X1   g17413(.A1(new_n17506_), .A2(new_n17651_), .B(new_n17653_), .ZN(new_n17670_));
  AOI22_X1   g17414(.A1(new_n13460_), .A2(new_n2208_), .B1(\b[63] ), .B2(new_n2361_), .ZN(new_n17671_));
  OAI22_X1   g17415(.A1(new_n12151_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n11195_), .ZN(new_n17672_));
  AOI21_X1   g17416(.A1(\b[57] ), .A2(new_n3456_), .B(new_n17672_), .ZN(new_n17673_));
  OAI21_X1   g17417(.A1(new_n12203_), .A2(new_n3261_), .B(new_n17673_), .ZN(new_n17674_));
  XOR2_X1    g17418(.A1(new_n17674_), .A2(new_n3264_), .Z(new_n17675_));
  AOI22_X1   g17419(.A1(new_n3864_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n3869_), .ZN(new_n17676_));
  OAI21_X1   g17420(.A1(new_n9942_), .A2(new_n5410_), .B(new_n17676_), .ZN(new_n17677_));
  AOI21_X1   g17421(.A1(new_n10318_), .A2(new_n3872_), .B(new_n17677_), .ZN(new_n17678_));
  XOR2_X1    g17422(.A1(new_n17678_), .A2(new_n3876_), .Z(new_n17679_));
  INV_X1     g17423(.I(new_n17679_), .ZN(new_n17680_));
  INV_X1     g17424(.I(new_n17531_), .ZN(new_n17681_));
  NOR2_X1    g17425(.A1(new_n17632_), .A2(new_n17634_), .ZN(new_n17682_));
  NAND2_X1   g17426(.A1(new_n17632_), .A2(new_n17634_), .ZN(new_n17683_));
  AOI21_X1   g17427(.A1(new_n17681_), .A2(new_n17683_), .B(new_n17682_), .ZN(new_n17684_));
  OAI22_X1   g17428(.A1(new_n9376_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n9032_), .ZN(new_n17685_));
  AOI21_X1   g17429(.A1(\b[51] ), .A2(new_n4706_), .B(new_n17685_), .ZN(new_n17686_));
  OAI21_X1   g17430(.A1(new_n9385_), .A2(new_n4458_), .B(new_n17686_), .ZN(new_n17687_));
  XOR2_X1    g17431(.A1(new_n17687_), .A2(new_n4446_), .Z(new_n17688_));
  AOI22_X1   g17432(.A1(new_n5155_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n5160_), .ZN(new_n17689_));
  OAI21_X1   g17433(.A1(new_n8127_), .A2(new_n6877_), .B(new_n17689_), .ZN(new_n17690_));
  AOI21_X1   g17434(.A1(new_n9684_), .A2(new_n5166_), .B(new_n17690_), .ZN(new_n17691_));
  XOR2_X1    g17435(.A1(new_n17691_), .A2(new_n5162_), .Z(new_n17692_));
  AOI22_X1   g17436(.A1(new_n6569_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n6574_), .ZN(new_n17693_));
  OAI21_X1   g17437(.A1(new_n6490_), .A2(new_n8565_), .B(new_n17693_), .ZN(new_n17694_));
  AOI21_X1   g17438(.A1(new_n7906_), .A2(new_n6579_), .B(new_n17694_), .ZN(new_n17695_));
  XOR2_X1    g17439(.A1(new_n17695_), .A2(new_n6567_), .Z(new_n17696_));
  INV_X1     g17440(.I(new_n17696_), .ZN(new_n17697_));
  OAI21_X1   g17441(.A1(new_n17541_), .A2(new_n17600_), .B(new_n17602_), .ZN(new_n17698_));
  INV_X1     g17442(.I(new_n17698_), .ZN(new_n17699_));
  AOI22_X1   g17443(.A1(new_n8241_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n8246_), .ZN(new_n17700_));
  OAI21_X1   g17444(.A1(new_n4886_), .A2(new_n9114_), .B(new_n17700_), .ZN(new_n17701_));
  AOI21_X1   g17445(.A1(new_n5351_), .A2(new_n8252_), .B(new_n17701_), .ZN(new_n17702_));
  XOR2_X1    g17446(.A1(new_n17702_), .A2(new_n8248_), .Z(new_n17703_));
  AOI21_X1   g17447(.A1(new_n17548_), .A2(new_n17587_), .B(new_n17585_), .ZN(new_n17704_));
  INV_X1     g17448(.I(new_n17704_), .ZN(new_n17705_));
  OAI22_X1   g17449(.A1(new_n10390_), .A2(new_n4666_), .B1(new_n4639_), .B2(new_n10389_), .ZN(new_n17706_));
  AOI21_X1   g17450(.A1(\b[33] ), .A2(new_n9471_), .B(new_n17706_), .ZN(new_n17707_));
  OAI21_X1   g17451(.A1(new_n4676_), .A2(new_n10388_), .B(new_n17707_), .ZN(new_n17708_));
  XOR2_X1    g17452(.A1(new_n17708_), .A2(\a[53] ), .Z(new_n17709_));
  AOI22_X1   g17453(.A1(new_n10064_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n10062_), .ZN(new_n17710_));
  OAI21_X1   g17454(.A1(new_n3624_), .A2(new_n10399_), .B(new_n17710_), .ZN(new_n17711_));
  AOI21_X1   g17455(.A1(new_n4030_), .A2(new_n10068_), .B(new_n17711_), .ZN(new_n17712_));
  XOR2_X1    g17456(.A1(new_n17712_), .A2(new_n10057_), .Z(new_n17713_));
  AOI22_X1   g17457(.A1(new_n11926_), .A2(\b[26] ), .B1(new_n11924_), .B2(\b[25] ), .ZN(new_n17714_));
  OAI21_X1   g17458(.A1(new_n2495_), .A2(new_n12317_), .B(new_n17714_), .ZN(new_n17715_));
  AOI21_X1   g17459(.A1(new_n3407_), .A2(new_n11929_), .B(new_n17715_), .ZN(new_n17716_));
  XOR2_X1    g17460(.A1(new_n17716_), .A2(new_n12312_), .Z(new_n17717_));
  AOI22_X1   g17461(.A1(new_n12922_), .A2(\b[23] ), .B1(\b[22] ), .B2(new_n12923_), .ZN(new_n17718_));
  INV_X1     g17462(.I(new_n17718_), .ZN(new_n17719_));
  NOR2_X1    g17463(.A1(new_n17719_), .A2(new_n17561_), .ZN(new_n17720_));
  INV_X1     g17464(.I(new_n17720_), .ZN(new_n17721_));
  NAND2_X1   g17465(.A1(new_n17719_), .A2(new_n17561_), .ZN(new_n17722_));
  NAND2_X1   g17466(.A1(new_n17721_), .A2(new_n17722_), .ZN(new_n17723_));
  XOR2_X1    g17467(.A1(new_n17717_), .A2(new_n17723_), .Z(new_n17724_));
  AOI22_X1   g17468(.A1(new_n10981_), .A2(\b[29] ), .B1(new_n10979_), .B2(\b[28] ), .ZN(new_n17725_));
  OAI21_X1   g17469(.A1(new_n3158_), .A2(new_n11306_), .B(new_n17725_), .ZN(new_n17726_));
  AOI21_X1   g17470(.A1(new_n4188_), .A2(new_n10984_), .B(new_n17726_), .ZN(new_n17727_));
  XOR2_X1    g17471(.A1(new_n17727_), .A2(new_n10989_), .Z(new_n17728_));
  AOI21_X1   g17472(.A1(new_n17558_), .A2(new_n17562_), .B(new_n17563_), .ZN(new_n17729_));
  NOR2_X1    g17473(.A1(new_n17728_), .A2(new_n17729_), .ZN(new_n17730_));
  INV_X1     g17474(.I(new_n17730_), .ZN(new_n17731_));
  NAND2_X1   g17475(.A1(new_n17728_), .A2(new_n17729_), .ZN(new_n17732_));
  NAND2_X1   g17476(.A1(new_n17731_), .A2(new_n17732_), .ZN(new_n17733_));
  XOR2_X1    g17477(.A1(new_n17733_), .A2(new_n17724_), .Z(new_n17734_));
  INV_X1     g17478(.I(new_n17734_), .ZN(new_n17735_));
  OAI21_X1   g17479(.A1(new_n17553_), .A2(new_n17567_), .B(new_n17569_), .ZN(new_n17736_));
  NAND2_X1   g17480(.A1(new_n17735_), .A2(new_n17736_), .ZN(new_n17737_));
  NOR2_X1    g17481(.A1(new_n17735_), .A2(new_n17736_), .ZN(new_n17738_));
  INV_X1     g17482(.I(new_n17738_), .ZN(new_n17739_));
  NAND2_X1   g17483(.A1(new_n17739_), .A2(new_n17737_), .ZN(new_n17740_));
  XOR2_X1    g17484(.A1(new_n17740_), .A2(new_n17713_), .Z(new_n17741_));
  AOI21_X1   g17485(.A1(new_n17549_), .A2(new_n17578_), .B(new_n17577_), .ZN(new_n17742_));
  XOR2_X1    g17486(.A1(new_n17741_), .A2(new_n17742_), .Z(new_n17743_));
  XOR2_X1    g17487(.A1(new_n17743_), .A2(new_n17709_), .Z(new_n17744_));
  NOR2_X1    g17488(.A1(new_n17744_), .A2(new_n17705_), .ZN(new_n17745_));
  INV_X1     g17489(.I(new_n17745_), .ZN(new_n17746_));
  NAND2_X1   g17490(.A1(new_n17744_), .A2(new_n17705_), .ZN(new_n17747_));
  NAND2_X1   g17491(.A1(new_n17746_), .A2(new_n17747_), .ZN(new_n17748_));
  XNOR2_X1   g17492(.A1(new_n17748_), .A2(new_n17703_), .ZN(new_n17749_));
  OAI22_X1   g17493(.A1(new_n6284_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n6285_), .ZN(new_n17750_));
  AOI21_X1   g17494(.A1(\b[39] ), .A2(new_n7719_), .B(new_n17750_), .ZN(new_n17751_));
  OAI21_X1   g17495(.A1(new_n6299_), .A2(new_n8585_), .B(new_n17751_), .ZN(new_n17752_));
  XOR2_X1    g17496(.A1(new_n17752_), .A2(\a[47] ), .Z(new_n17753_));
  INV_X1     g17497(.I(new_n17589_), .ZN(new_n17754_));
  AOI21_X1   g17498(.A1(new_n17754_), .A2(new_n17597_), .B(new_n17595_), .ZN(new_n17755_));
  NOR2_X1    g17499(.A1(new_n17753_), .A2(new_n17755_), .ZN(new_n17756_));
  INV_X1     g17500(.I(new_n17756_), .ZN(new_n17757_));
  NAND2_X1   g17501(.A1(new_n17753_), .A2(new_n17755_), .ZN(new_n17758_));
  NAND2_X1   g17502(.A1(new_n17757_), .A2(new_n17758_), .ZN(new_n17759_));
  XNOR2_X1   g17503(.A1(new_n17749_), .A2(new_n17759_), .ZN(new_n17760_));
  NOR2_X1    g17504(.A1(new_n17760_), .A2(new_n17699_), .ZN(new_n17761_));
  INV_X1     g17505(.I(new_n17761_), .ZN(new_n17762_));
  NAND2_X1   g17506(.A1(new_n17760_), .A2(new_n17699_), .ZN(new_n17763_));
  NAND2_X1   g17507(.A1(new_n17762_), .A2(new_n17763_), .ZN(new_n17764_));
  XOR2_X1    g17508(.A1(new_n17764_), .A2(new_n17697_), .Z(new_n17765_));
  AOI22_X1   g17509(.A1(new_n6108_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n6111_), .ZN(new_n17766_));
  OAI21_X1   g17510(.A1(new_n7096_), .A2(new_n7708_), .B(new_n17766_), .ZN(new_n17767_));
  AOI21_X1   g17511(.A1(new_n7649_), .A2(new_n6105_), .B(new_n17767_), .ZN(new_n17768_));
  XOR2_X1    g17512(.A1(new_n17768_), .A2(new_n5849_), .Z(new_n17769_));
  NOR2_X1    g17513(.A1(new_n17612_), .A2(new_n17537_), .ZN(new_n17770_));
  NOR2_X1    g17514(.A1(new_n17770_), .A2(new_n17610_), .ZN(new_n17771_));
  NOR2_X1    g17515(.A1(new_n17771_), .A2(new_n17769_), .ZN(new_n17772_));
  AND2_X2    g17516(.A1(new_n17771_), .A2(new_n17769_), .Z(new_n17773_));
  NOR2_X1    g17517(.A1(new_n17773_), .A2(new_n17772_), .ZN(new_n17774_));
  XOR2_X1    g17518(.A1(new_n17774_), .A2(new_n17765_), .Z(new_n17775_));
  AOI21_X1   g17519(.A1(new_n17536_), .A2(new_n17618_), .B(new_n17616_), .ZN(new_n17776_));
  NOR2_X1    g17520(.A1(new_n17775_), .A2(new_n17776_), .ZN(new_n17777_));
  INV_X1     g17521(.I(new_n17777_), .ZN(new_n17778_));
  NAND2_X1   g17522(.A1(new_n17775_), .A2(new_n17776_), .ZN(new_n17779_));
  NAND2_X1   g17523(.A1(new_n17778_), .A2(new_n17779_), .ZN(new_n17780_));
  XOR2_X1    g17524(.A1(new_n17780_), .A2(new_n17692_), .Z(new_n17781_));
  INV_X1     g17525(.I(new_n17781_), .ZN(new_n17782_));
  AOI21_X1   g17526(.A1(new_n17621_), .A2(new_n17630_), .B(new_n17628_), .ZN(new_n17783_));
  NOR2_X1    g17527(.A1(new_n17782_), .A2(new_n17783_), .ZN(new_n17784_));
  INV_X1     g17528(.I(new_n17784_), .ZN(new_n17785_));
  NAND2_X1   g17529(.A1(new_n17782_), .A2(new_n17783_), .ZN(new_n17786_));
  NAND2_X1   g17530(.A1(new_n17785_), .A2(new_n17786_), .ZN(new_n17787_));
  XOR2_X1    g17531(.A1(new_n17787_), .A2(new_n17688_), .Z(new_n17788_));
  NOR2_X1    g17532(.A1(new_n17788_), .A2(new_n17684_), .ZN(new_n17789_));
  INV_X1     g17533(.I(new_n17789_), .ZN(new_n17790_));
  NAND2_X1   g17534(.A1(new_n17788_), .A2(new_n17684_), .ZN(new_n17791_));
  NAND2_X1   g17535(.A1(new_n17790_), .A2(new_n17791_), .ZN(new_n17792_));
  XOR2_X1    g17536(.A1(new_n17792_), .A2(new_n17680_), .Z(new_n17793_));
  NOR2_X1    g17537(.A1(new_n17639_), .A2(new_n17523_), .ZN(new_n17794_));
  NOR2_X1    g17538(.A1(new_n17794_), .A2(new_n17637_), .ZN(new_n17795_));
  NOR2_X1    g17539(.A1(new_n17793_), .A2(new_n17795_), .ZN(new_n17796_));
  INV_X1     g17540(.I(new_n17796_), .ZN(new_n17797_));
  NAND2_X1   g17541(.A1(new_n17793_), .A2(new_n17795_), .ZN(new_n17798_));
  NAND2_X1   g17542(.A1(new_n17797_), .A2(new_n17798_), .ZN(new_n17799_));
  XOR2_X1    g17543(.A1(new_n17799_), .A2(new_n17675_), .Z(new_n17800_));
  XOR2_X1    g17544(.A1(new_n17800_), .A2(new_n2714_), .Z(new_n17801_));
  AOI22_X1   g17545(.A1(new_n2716_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n2719_), .ZN(new_n17802_));
  OAI21_X1   g17546(.A1(new_n12147_), .A2(new_n2924_), .B(new_n17802_), .ZN(new_n17803_));
  NOR2_X1    g17547(.A1(new_n14950_), .A2(new_n2711_), .ZN(new_n17804_));
  NOR2_X1    g17548(.A1(new_n17804_), .A2(new_n17803_), .ZN(new_n17805_));
  OAI21_X1   g17549(.A1(new_n17519_), .A2(new_n17642_), .B(new_n17643_), .ZN(new_n17806_));
  XNOR2_X1   g17550(.A1(new_n17806_), .A2(new_n17805_), .ZN(new_n17807_));
  XOR2_X1    g17551(.A1(new_n17801_), .A2(new_n17807_), .Z(new_n17808_));
  XOR2_X1    g17552(.A1(new_n17808_), .A2(new_n17671_), .Z(new_n17809_));
  NAND2_X1   g17553(.A1(new_n17648_), .A2(new_n17513_), .ZN(new_n17810_));
  NAND2_X1   g17554(.A1(new_n17810_), .A2(new_n17647_), .ZN(new_n17811_));
  XOR2_X1    g17555(.A1(new_n17811_), .A2(\a[23] ), .Z(new_n17812_));
  XOR2_X1    g17556(.A1(new_n17809_), .A2(new_n17812_), .Z(new_n17813_));
  INV_X1     g17557(.I(new_n17813_), .ZN(new_n17814_));
  NAND2_X1   g17558(.A1(new_n17814_), .A2(new_n17670_), .ZN(new_n17815_));
  NOR2_X1    g17559(.A1(new_n17814_), .A2(new_n17670_), .ZN(new_n17816_));
  INV_X1     g17560(.I(new_n17816_), .ZN(new_n17817_));
  AND2_X2    g17561(.A1(new_n17817_), .A2(new_n17815_), .Z(new_n17818_));
  XOR2_X1    g17562(.A1(new_n17669_), .A2(new_n17818_), .Z(\f[86] ));
  INV_X1     g17563(.I(new_n17811_), .ZN(new_n17820_));
  NOR2_X1    g17564(.A1(new_n17808_), .A2(new_n17820_), .ZN(new_n17821_));
  XOR2_X1    g17565(.A1(new_n17671_), .A2(new_n2200_), .Z(new_n17822_));
  AOI21_X1   g17566(.A1(new_n17808_), .A2(new_n17820_), .B(new_n17822_), .ZN(new_n17823_));
  NOR2_X1    g17567(.A1(new_n17823_), .A2(new_n17821_), .ZN(new_n17824_));
  INV_X1     g17568(.I(new_n17824_), .ZN(new_n17825_));
  INV_X1     g17569(.I(new_n17800_), .ZN(new_n17826_));
  INV_X1     g17570(.I(new_n17806_), .ZN(new_n17827_));
  XOR2_X1    g17571(.A1(new_n17805_), .A2(new_n2714_), .Z(new_n17828_));
  AOI21_X1   g17572(.A1(new_n17800_), .A2(new_n17827_), .B(new_n17828_), .ZN(new_n17829_));
  AOI21_X1   g17573(.A1(new_n17826_), .A2(new_n17806_), .B(new_n17829_), .ZN(new_n17830_));
  INV_X1     g17574(.I(new_n17830_), .ZN(new_n17831_));
  AOI22_X1   g17575(.A1(new_n2716_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n2719_), .ZN(new_n17832_));
  OAI21_X1   g17576(.A1(new_n12148_), .A2(new_n2924_), .B(new_n17832_), .ZN(new_n17833_));
  AOI21_X1   g17577(.A1(new_n12811_), .A2(new_n2722_), .B(new_n17833_), .ZN(new_n17834_));
  XOR2_X1    g17578(.A1(new_n17834_), .A2(new_n2714_), .Z(new_n17835_));
  AOI21_X1   g17579(.A1(new_n17675_), .A2(new_n17798_), .B(new_n17796_), .ZN(new_n17836_));
  AOI22_X1   g17580(.A1(new_n3267_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n3270_), .ZN(new_n17837_));
  OAI21_X1   g17581(.A1(new_n11195_), .A2(new_n3475_), .B(new_n17837_), .ZN(new_n17838_));
  AOI21_X1   g17582(.A1(new_n11836_), .A2(new_n3273_), .B(new_n17838_), .ZN(new_n17839_));
  XOR2_X1    g17583(.A1(new_n17839_), .A2(new_n3264_), .Z(new_n17840_));
  INV_X1     g17584(.I(new_n17840_), .ZN(new_n17841_));
  AOI21_X1   g17585(.A1(new_n17680_), .A2(new_n17791_), .B(new_n17789_), .ZN(new_n17842_));
  AOI22_X1   g17586(.A1(new_n3864_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n3869_), .ZN(new_n17843_));
  OAI21_X1   g17587(.A1(new_n9972_), .A2(new_n5410_), .B(new_n17843_), .ZN(new_n17844_));
  AOI21_X1   g17588(.A1(new_n10631_), .A2(new_n3872_), .B(new_n17844_), .ZN(new_n17845_));
  XOR2_X1    g17589(.A1(new_n17845_), .A2(new_n3876_), .Z(new_n17846_));
  INV_X1     g17590(.I(new_n17846_), .ZN(new_n17847_));
  AOI21_X1   g17591(.A1(new_n17688_), .A2(new_n17786_), .B(new_n17784_), .ZN(new_n17848_));
  INV_X1     g17592(.I(new_n17848_), .ZN(new_n17849_));
  AOI22_X1   g17593(.A1(new_n4918_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n4921_), .ZN(new_n17850_));
  OAI21_X1   g17594(.A1(new_n9032_), .A2(new_n6099_), .B(new_n17850_), .ZN(new_n17851_));
  AOI21_X1   g17595(.A1(new_n10884_), .A2(new_n4699_), .B(new_n17851_), .ZN(new_n17852_));
  XOR2_X1    g17596(.A1(new_n17852_), .A2(new_n4446_), .Z(new_n17853_));
  INV_X1     g17597(.I(new_n17692_), .ZN(new_n17854_));
  AOI21_X1   g17598(.A1(new_n17854_), .A2(new_n17779_), .B(new_n17777_), .ZN(new_n17855_));
  INV_X1     g17599(.I(new_n17855_), .ZN(new_n17856_));
  AOI21_X1   g17600(.A1(new_n17697_), .A2(new_n17763_), .B(new_n17761_), .ZN(new_n17857_));
  INV_X1     g17601(.I(new_n17857_), .ZN(new_n17858_));
  INV_X1     g17602(.I(new_n17749_), .ZN(new_n17859_));
  AOI21_X1   g17603(.A1(new_n17859_), .A2(new_n17758_), .B(new_n17756_), .ZN(new_n17860_));
  OAI21_X1   g17604(.A1(new_n17703_), .A2(new_n17745_), .B(new_n17747_), .ZN(new_n17861_));
  OAI21_X1   g17605(.A1(new_n17713_), .A2(new_n17738_), .B(new_n17737_), .ZN(new_n17862_));
  AOI21_X1   g17606(.A1(new_n17724_), .A2(new_n17732_), .B(new_n17730_), .ZN(new_n17863_));
  AOI22_X1   g17607(.A1(new_n10981_), .A2(\b[30] ), .B1(new_n10979_), .B2(\b[29] ), .ZN(new_n17864_));
  OAI21_X1   g17608(.A1(new_n3185_), .A2(new_n11306_), .B(new_n17864_), .ZN(new_n17865_));
  AOI21_X1   g17609(.A1(new_n4230_), .A2(new_n10984_), .B(new_n17865_), .ZN(new_n17866_));
  XOR2_X1    g17610(.A1(new_n17866_), .A2(new_n10989_), .Z(new_n17867_));
  OAI21_X1   g17611(.A1(new_n17717_), .A2(new_n17720_), .B(new_n17722_), .ZN(new_n17868_));
  INV_X1     g17612(.I(new_n17868_), .ZN(new_n17869_));
  OAI22_X1   g17613(.A1(new_n13224_), .A2(new_n3158_), .B1(new_n3006_), .B2(new_n11923_), .ZN(new_n17870_));
  AOI21_X1   g17614(.A1(\b[25] ), .A2(new_n13223_), .B(new_n17870_), .ZN(new_n17871_));
  OAI21_X1   g17615(.A1(new_n3165_), .A2(new_n11930_), .B(new_n17871_), .ZN(new_n17872_));
  XOR2_X1    g17616(.A1(new_n17872_), .A2(\a[62] ), .Z(new_n17873_));
  INV_X1     g17617(.I(new_n17873_), .ZN(new_n17874_));
  AOI22_X1   g17618(.A1(new_n12922_), .A2(\b[24] ), .B1(\b[23] ), .B2(new_n12923_), .ZN(new_n17875_));
  INV_X1     g17619(.I(new_n17875_), .ZN(new_n17876_));
  NOR2_X1    g17620(.A1(new_n17876_), .A2(new_n2200_), .ZN(new_n17877_));
  NOR2_X1    g17621(.A1(new_n17875_), .A2(\a[23] ), .ZN(new_n17878_));
  NOR2_X1    g17622(.A1(new_n17877_), .A2(new_n17878_), .ZN(new_n17879_));
  XOR2_X1    g17623(.A1(new_n17879_), .A2(new_n17718_), .Z(new_n17880_));
  NOR2_X1    g17624(.A1(new_n17874_), .A2(new_n17880_), .ZN(new_n17881_));
  NAND2_X1   g17625(.A1(new_n17874_), .A2(new_n17880_), .ZN(new_n17882_));
  INV_X1     g17626(.I(new_n17882_), .ZN(new_n17883_));
  NOR2_X1    g17627(.A1(new_n17883_), .A2(new_n17881_), .ZN(new_n17884_));
  XOR2_X1    g17628(.A1(new_n17884_), .A2(new_n17869_), .Z(new_n17885_));
  NOR2_X1    g17629(.A1(new_n17885_), .A2(new_n17867_), .ZN(new_n17886_));
  INV_X1     g17630(.I(new_n17886_), .ZN(new_n17887_));
  NAND2_X1   g17631(.A1(new_n17885_), .A2(new_n17867_), .ZN(new_n17888_));
  NAND2_X1   g17632(.A1(new_n17887_), .A2(new_n17888_), .ZN(new_n17889_));
  XOR2_X1    g17633(.A1(new_n17889_), .A2(new_n17863_), .Z(new_n17890_));
  AOI22_X1   g17634(.A1(new_n10064_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n10062_), .ZN(new_n17891_));
  OAI21_X1   g17635(.A1(new_n4022_), .A2(new_n10399_), .B(new_n17891_), .ZN(new_n17892_));
  AOI21_X1   g17636(.A1(new_n4223_), .A2(new_n10068_), .B(new_n17892_), .ZN(new_n17893_));
  XOR2_X1    g17637(.A1(new_n17893_), .A2(\a[56] ), .Z(new_n17894_));
  NAND2_X1   g17638(.A1(new_n17890_), .A2(new_n17894_), .ZN(new_n17895_));
  OR2_X2     g17639(.A1(new_n17890_), .A2(new_n17894_), .Z(new_n17896_));
  NAND2_X1   g17640(.A1(new_n17896_), .A2(new_n17895_), .ZN(new_n17897_));
  XNOR2_X1   g17641(.A1(new_n17897_), .A2(new_n17862_), .ZN(new_n17898_));
  AOI22_X1   g17642(.A1(new_n9125_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n9123_), .ZN(new_n17899_));
  OAI21_X1   g17643(.A1(new_n4639_), .A2(new_n9470_), .B(new_n17899_), .ZN(new_n17900_));
  AOI21_X1   g17644(.A1(new_n5594_), .A2(new_n9129_), .B(new_n17900_), .ZN(new_n17901_));
  XOR2_X1    g17645(.A1(new_n17901_), .A2(new_n9133_), .Z(new_n17902_));
  INV_X1     g17646(.I(new_n17741_), .ZN(new_n17903_));
  NOR2_X1    g17647(.A1(new_n17903_), .A2(new_n17742_), .ZN(new_n17904_));
  AOI21_X1   g17648(.A1(new_n17903_), .A2(new_n17742_), .B(new_n17709_), .ZN(new_n17905_));
  NOR2_X1    g17649(.A1(new_n17905_), .A2(new_n17904_), .ZN(new_n17906_));
  NOR2_X1    g17650(.A1(new_n17906_), .A2(new_n17902_), .ZN(new_n17907_));
  NAND2_X1   g17651(.A1(new_n17906_), .A2(new_n17902_), .ZN(new_n17908_));
  INV_X1     g17652(.I(new_n17908_), .ZN(new_n17909_));
  NOR2_X1    g17653(.A1(new_n17909_), .A2(new_n17907_), .ZN(new_n17910_));
  XOR2_X1    g17654(.A1(new_n17910_), .A2(new_n17898_), .Z(new_n17911_));
  AOI22_X1   g17655(.A1(new_n8241_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n8246_), .ZN(new_n17912_));
  OAI21_X1   g17656(.A1(new_n5312_), .A2(new_n9114_), .B(new_n17912_), .ZN(new_n17913_));
  AOI21_X1   g17657(.A1(new_n6310_), .A2(new_n8252_), .B(new_n17913_), .ZN(new_n17914_));
  XOR2_X1    g17658(.A1(new_n17914_), .A2(\a[50] ), .Z(new_n17915_));
  NAND2_X1   g17659(.A1(new_n17911_), .A2(new_n17915_), .ZN(new_n17916_));
  OR2_X2     g17660(.A1(new_n17911_), .A2(new_n17915_), .Z(new_n17917_));
  NAND2_X1   g17661(.A1(new_n17917_), .A2(new_n17916_), .ZN(new_n17918_));
  XNOR2_X1   g17662(.A1(new_n17918_), .A2(new_n17861_), .ZN(new_n17919_));
  INV_X1     g17663(.I(new_n17919_), .ZN(new_n17920_));
  AOI22_X1   g17664(.A1(new_n7403_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n7408_), .ZN(new_n17921_));
  OAI21_X1   g17665(.A1(new_n6284_), .A2(new_n9488_), .B(new_n17921_), .ZN(new_n17922_));
  AOI21_X1   g17666(.A1(new_n7106_), .A2(new_n7414_), .B(new_n17922_), .ZN(new_n17923_));
  XOR2_X1    g17667(.A1(new_n17923_), .A2(new_n7410_), .Z(new_n17924_));
  NOR2_X1    g17668(.A1(new_n17920_), .A2(new_n17924_), .ZN(new_n17925_));
  NAND2_X1   g17669(.A1(new_n17920_), .A2(new_n17924_), .ZN(new_n17926_));
  INV_X1     g17670(.I(new_n17926_), .ZN(new_n17927_));
  NOR2_X1    g17671(.A1(new_n17927_), .A2(new_n17925_), .ZN(new_n17928_));
  XOR2_X1    g17672(.A1(new_n17928_), .A2(new_n17860_), .Z(new_n17929_));
  AOI22_X1   g17673(.A1(new_n6569_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n6574_), .ZN(new_n17930_));
  OAI21_X1   g17674(.A1(new_n6775_), .A2(new_n8565_), .B(new_n17930_), .ZN(new_n17931_));
  AOI21_X1   g17675(.A1(new_n7926_), .A2(new_n6579_), .B(new_n17931_), .ZN(new_n17932_));
  XOR2_X1    g17676(.A1(new_n17932_), .A2(new_n6567_), .Z(new_n17933_));
  NOR2_X1    g17677(.A1(new_n17929_), .A2(new_n17933_), .ZN(new_n17934_));
  NAND2_X1   g17678(.A1(new_n17929_), .A2(new_n17933_), .ZN(new_n17935_));
  INV_X1     g17679(.I(new_n17935_), .ZN(new_n17936_));
  NOR2_X1    g17680(.A1(new_n17936_), .A2(new_n17934_), .ZN(new_n17937_));
  XOR2_X1    g17681(.A1(new_n17937_), .A2(new_n17858_), .Z(new_n17938_));
  AOI22_X1   g17682(.A1(new_n6108_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n6111_), .ZN(new_n17939_));
  OAI21_X1   g17683(.A1(new_n7617_), .A2(new_n7708_), .B(new_n17939_), .ZN(new_n17940_));
  AOI21_X1   g17684(.A1(new_n8792_), .A2(new_n6105_), .B(new_n17940_), .ZN(new_n17941_));
  XOR2_X1    g17685(.A1(new_n17941_), .A2(\a[41] ), .Z(new_n17942_));
  INV_X1     g17686(.I(new_n17772_), .ZN(new_n17943_));
  OAI21_X1   g17687(.A1(new_n17765_), .A2(new_n17773_), .B(new_n17943_), .ZN(new_n17944_));
  NAND2_X1   g17688(.A1(new_n17944_), .A2(new_n17942_), .ZN(new_n17945_));
  OR2_X2     g17689(.A1(new_n17944_), .A2(new_n17942_), .Z(new_n17946_));
  NAND2_X1   g17690(.A1(new_n17946_), .A2(new_n17945_), .ZN(new_n17947_));
  XNOR2_X1   g17691(.A1(new_n17938_), .A2(new_n17947_), .ZN(new_n17948_));
  INV_X1     g17692(.I(new_n17948_), .ZN(new_n17949_));
  AOI22_X1   g17693(.A1(new_n5155_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n5160_), .ZN(new_n17950_));
  OAI21_X1   g17694(.A1(new_n8168_), .A2(new_n6877_), .B(new_n17950_), .ZN(new_n17951_));
  AOI21_X1   g17695(.A1(new_n8783_), .A2(new_n5166_), .B(new_n17951_), .ZN(new_n17952_));
  XOR2_X1    g17696(.A1(new_n17952_), .A2(new_n5162_), .Z(new_n17953_));
  NOR2_X1    g17697(.A1(new_n17949_), .A2(new_n17953_), .ZN(new_n17954_));
  INV_X1     g17698(.I(new_n17954_), .ZN(new_n17955_));
  NAND2_X1   g17699(.A1(new_n17949_), .A2(new_n17953_), .ZN(new_n17956_));
  NAND2_X1   g17700(.A1(new_n17955_), .A2(new_n17956_), .ZN(new_n17957_));
  XOR2_X1    g17701(.A1(new_n17957_), .A2(new_n17856_), .Z(new_n17958_));
  NOR2_X1    g17702(.A1(new_n17958_), .A2(new_n17853_), .ZN(new_n17959_));
  NAND2_X1   g17703(.A1(new_n17958_), .A2(new_n17853_), .ZN(new_n17960_));
  INV_X1     g17704(.I(new_n17960_), .ZN(new_n17961_));
  NOR2_X1    g17705(.A1(new_n17961_), .A2(new_n17959_), .ZN(new_n17962_));
  XOR2_X1    g17706(.A1(new_n17962_), .A2(new_n17849_), .Z(new_n17963_));
  NOR2_X1    g17707(.A1(new_n17963_), .A2(new_n17847_), .ZN(new_n17964_));
  NAND2_X1   g17708(.A1(new_n17963_), .A2(new_n17847_), .ZN(new_n17965_));
  INV_X1     g17709(.I(new_n17965_), .ZN(new_n17966_));
  NOR2_X1    g17710(.A1(new_n17966_), .A2(new_n17964_), .ZN(new_n17967_));
  XNOR2_X1   g17711(.A1(new_n17967_), .A2(new_n17842_), .ZN(new_n17968_));
  NOR2_X1    g17712(.A1(new_n17968_), .A2(new_n17841_), .ZN(new_n17969_));
  INV_X1     g17713(.I(new_n17969_), .ZN(new_n17970_));
  NAND2_X1   g17714(.A1(new_n17968_), .A2(new_n17841_), .ZN(new_n17971_));
  NAND2_X1   g17715(.A1(new_n17970_), .A2(new_n17971_), .ZN(new_n17972_));
  XNOR2_X1   g17716(.A1(new_n17972_), .A2(new_n17836_), .ZN(new_n17973_));
  NOR2_X1    g17717(.A1(new_n17973_), .A2(new_n17835_), .ZN(new_n17974_));
  INV_X1     g17718(.I(new_n17974_), .ZN(new_n17975_));
  NAND2_X1   g17719(.A1(new_n17973_), .A2(new_n17835_), .ZN(new_n17976_));
  NAND2_X1   g17720(.A1(new_n17975_), .A2(new_n17976_), .ZN(new_n17977_));
  XOR2_X1    g17721(.A1(new_n17977_), .A2(new_n17831_), .Z(new_n17978_));
  INV_X1     g17722(.I(new_n17978_), .ZN(new_n17979_));
  NAND2_X1   g17723(.A1(new_n17979_), .A2(new_n17825_), .ZN(new_n17980_));
  NOR2_X1    g17724(.A1(new_n17979_), .A2(new_n17825_), .ZN(new_n17981_));
  INV_X1     g17725(.I(new_n17981_), .ZN(new_n17982_));
  AND2_X2    g17726(.A1(new_n17982_), .A2(new_n17980_), .Z(new_n17983_));
  INV_X1     g17727(.I(new_n17983_), .ZN(new_n17984_));
  AOI21_X1   g17728(.A1(new_n17669_), .A2(new_n17818_), .B(new_n17816_), .ZN(new_n17985_));
  XOR2_X1    g17729(.A1(new_n17985_), .A2(new_n17984_), .Z(\f[87] ));
  AOI21_X1   g17730(.A1(new_n17831_), .A2(new_n17976_), .B(new_n17974_), .ZN(new_n17987_));
  OAI22_X1   g17731(.A1(new_n2924_), .A2(new_n12796_), .B1(new_n12800_), .B2(new_n2708_), .ZN(new_n17988_));
  AOI21_X1   g17732(.A1(new_n13973_), .A2(new_n2722_), .B(new_n17988_), .ZN(new_n17989_));
  XOR2_X1    g17733(.A1(new_n17989_), .A2(new_n2714_), .Z(new_n17990_));
  OAI21_X1   g17734(.A1(new_n17836_), .A2(new_n17969_), .B(new_n17971_), .ZN(new_n17991_));
  OAI22_X1   g17735(.A1(new_n12148_), .A2(new_n3253_), .B1(new_n3258_), .B2(new_n12147_), .ZN(new_n17992_));
  AOI21_X1   g17736(.A1(\b[59] ), .A2(new_n3456_), .B(new_n17992_), .ZN(new_n17993_));
  OAI21_X1   g17737(.A1(new_n13110_), .A2(new_n3261_), .B(new_n17993_), .ZN(new_n17994_));
  XOR2_X1    g17738(.A1(new_n17994_), .A2(new_n3264_), .Z(new_n17995_));
  OAI21_X1   g17739(.A1(new_n17842_), .A2(new_n17964_), .B(new_n17965_), .ZN(new_n17996_));
  AOI22_X1   g17740(.A1(new_n3864_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n3869_), .ZN(new_n17997_));
  OAI21_X1   g17741(.A1(new_n10308_), .A2(new_n5410_), .B(new_n17997_), .ZN(new_n17998_));
  AOI21_X1   g17742(.A1(new_n12164_), .A2(new_n3872_), .B(new_n17998_), .ZN(new_n17999_));
  XOR2_X1    g17743(.A1(new_n17999_), .A2(new_n3876_), .Z(new_n18000_));
  AOI21_X1   g17744(.A1(new_n17849_), .A2(new_n17960_), .B(new_n17959_), .ZN(new_n18001_));
  INV_X1     g17745(.I(new_n18001_), .ZN(new_n18002_));
  AOI21_X1   g17746(.A1(new_n17856_), .A2(new_n17956_), .B(new_n17954_), .ZN(new_n18003_));
  INV_X1     g17747(.I(new_n18003_), .ZN(new_n18004_));
  AOI22_X1   g17748(.A1(new_n5155_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n5160_), .ZN(new_n18005_));
  OAI21_X1   g17749(.A1(new_n8500_), .A2(new_n6877_), .B(new_n18005_), .ZN(new_n18006_));
  AOI21_X1   g17750(.A1(new_n9987_), .A2(new_n5166_), .B(new_n18006_), .ZN(new_n18007_));
  XOR2_X1    g17751(.A1(new_n18007_), .A2(new_n5162_), .Z(new_n18008_));
  AOI22_X1   g17752(.A1(new_n6569_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n6574_), .ZN(new_n18009_));
  OAI21_X1   g17753(.A1(new_n7074_), .A2(new_n8565_), .B(new_n18009_), .ZN(new_n18010_));
  AOI21_X1   g17754(.A1(new_n9337_), .A2(new_n6579_), .B(new_n18010_), .ZN(new_n18011_));
  XOR2_X1    g17755(.A1(new_n18011_), .A2(new_n6567_), .Z(new_n18012_));
  INV_X1     g17756(.I(new_n18012_), .ZN(new_n18013_));
  INV_X1     g17757(.I(new_n17916_), .ZN(new_n18014_));
  AOI21_X1   g17758(.A1(new_n17861_), .A2(new_n17917_), .B(new_n18014_), .ZN(new_n18015_));
  AOI22_X1   g17759(.A1(new_n8241_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n8246_), .ZN(new_n18016_));
  OAI21_X1   g17760(.A1(new_n5341_), .A2(new_n9114_), .B(new_n18016_), .ZN(new_n18017_));
  AOI21_X1   g17761(.A1(new_n5793_), .A2(new_n8252_), .B(new_n18017_), .ZN(new_n18018_));
  XOR2_X1    g17762(.A1(new_n18018_), .A2(new_n8248_), .Z(new_n18019_));
  AOI21_X1   g17763(.A1(new_n17898_), .A2(new_n17908_), .B(new_n17907_), .ZN(new_n18020_));
  INV_X1     g17764(.I(new_n18020_), .ZN(new_n18021_));
  AOI22_X1   g17765(.A1(new_n10064_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n10062_), .ZN(new_n18022_));
  OAI21_X1   g17766(.A1(new_n4023_), .A2(new_n10399_), .B(new_n18022_), .ZN(new_n18023_));
  AOI21_X1   g17767(.A1(new_n5103_), .A2(new_n10068_), .B(new_n18023_), .ZN(new_n18024_));
  XOR2_X1    g17768(.A1(new_n18024_), .A2(new_n10057_), .Z(new_n18025_));
  INV_X1     g17769(.I(new_n18025_), .ZN(new_n18026_));
  OAI21_X1   g17770(.A1(new_n17869_), .A2(new_n17881_), .B(new_n17882_), .ZN(new_n18027_));
  AOI22_X1   g17771(.A1(new_n11926_), .A2(\b[28] ), .B1(new_n11924_), .B2(\b[27] ), .ZN(new_n18028_));
  OAI21_X1   g17772(.A1(new_n3006_), .A2(new_n12317_), .B(new_n18028_), .ZN(new_n18029_));
  AOI21_X1   g17773(.A1(new_n3807_), .A2(new_n11929_), .B(new_n18029_), .ZN(new_n18030_));
  XOR2_X1    g17774(.A1(new_n18030_), .A2(\a[62] ), .Z(new_n18031_));
  NOR2_X1    g17775(.A1(new_n17878_), .A2(new_n17719_), .ZN(new_n18032_));
  NOR2_X1    g17776(.A1(new_n18032_), .A2(new_n17877_), .ZN(new_n18033_));
  AOI22_X1   g17777(.A1(new_n12922_), .A2(\b[25] ), .B1(\b[24] ), .B2(new_n12923_), .ZN(new_n18034_));
  NAND2_X1   g17778(.A1(new_n18033_), .A2(new_n18034_), .ZN(new_n18035_));
  NOR2_X1    g17779(.A1(new_n18033_), .A2(new_n18034_), .ZN(new_n18036_));
  INV_X1     g17780(.I(new_n18036_), .ZN(new_n18037_));
  NAND2_X1   g17781(.A1(new_n18037_), .A2(new_n18035_), .ZN(new_n18038_));
  XNOR2_X1   g17782(.A1(new_n18031_), .A2(new_n18038_), .ZN(new_n18039_));
  INV_X1     g17783(.I(new_n18039_), .ZN(new_n18040_));
  AOI22_X1   g17784(.A1(new_n10981_), .A2(\b[31] ), .B1(new_n10979_), .B2(\b[30] ), .ZN(new_n18041_));
  OAI21_X1   g17785(.A1(new_n3592_), .A2(new_n11306_), .B(new_n18041_), .ZN(new_n18042_));
  AOI21_X1   g17786(.A1(new_n3796_), .A2(new_n10984_), .B(new_n18042_), .ZN(new_n18043_));
  XOR2_X1    g17787(.A1(new_n18043_), .A2(new_n10989_), .Z(new_n18044_));
  NOR2_X1    g17788(.A1(new_n18044_), .A2(new_n18040_), .ZN(new_n18045_));
  NAND2_X1   g17789(.A1(new_n18044_), .A2(new_n18040_), .ZN(new_n18046_));
  INV_X1     g17790(.I(new_n18046_), .ZN(new_n18047_));
  NOR2_X1    g17791(.A1(new_n18047_), .A2(new_n18045_), .ZN(new_n18048_));
  XNOR2_X1   g17792(.A1(new_n18048_), .A2(new_n18027_), .ZN(new_n18049_));
  INV_X1     g17793(.I(new_n17863_), .ZN(new_n18050_));
  AOI21_X1   g17794(.A1(new_n18050_), .A2(new_n17888_), .B(new_n17886_), .ZN(new_n18051_));
  NOR2_X1    g17795(.A1(new_n18049_), .A2(new_n18051_), .ZN(new_n18052_));
  INV_X1     g17796(.I(new_n18052_), .ZN(new_n18053_));
  NAND2_X1   g17797(.A1(new_n18049_), .A2(new_n18051_), .ZN(new_n18054_));
  NAND2_X1   g17798(.A1(new_n18053_), .A2(new_n18054_), .ZN(new_n18055_));
  XOR2_X1    g17799(.A1(new_n18055_), .A2(new_n18026_), .Z(new_n18056_));
  INV_X1     g17800(.I(new_n17895_), .ZN(new_n18057_));
  AOI21_X1   g17801(.A1(new_n17862_), .A2(new_n17896_), .B(new_n18057_), .ZN(new_n18058_));
  OAI22_X1   g17802(.A1(new_n10390_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n10389_), .ZN(new_n18059_));
  AOI21_X1   g17803(.A1(\b[35] ), .A2(new_n9471_), .B(new_n18059_), .ZN(new_n18060_));
  OAI21_X1   g17804(.A1(new_n5322_), .A2(new_n10388_), .B(new_n18060_), .ZN(new_n18061_));
  XOR2_X1    g17805(.A1(new_n18061_), .A2(\a[53] ), .Z(new_n18062_));
  NOR2_X1    g17806(.A1(new_n18058_), .A2(new_n18062_), .ZN(new_n18063_));
  INV_X1     g17807(.I(new_n18063_), .ZN(new_n18064_));
  NAND2_X1   g17808(.A1(new_n18058_), .A2(new_n18062_), .ZN(new_n18065_));
  NAND2_X1   g17809(.A1(new_n18064_), .A2(new_n18065_), .ZN(new_n18066_));
  XOR2_X1    g17810(.A1(new_n18066_), .A2(new_n18056_), .Z(new_n18067_));
  NOR2_X1    g17811(.A1(new_n18067_), .A2(new_n18021_), .ZN(new_n18068_));
  INV_X1     g17812(.I(new_n18068_), .ZN(new_n18069_));
  NAND2_X1   g17813(.A1(new_n18067_), .A2(new_n18021_), .ZN(new_n18070_));
  NAND2_X1   g17814(.A1(new_n18069_), .A2(new_n18070_), .ZN(new_n18071_));
  XOR2_X1    g17815(.A1(new_n18071_), .A2(new_n18019_), .Z(new_n18072_));
  INV_X1     g17816(.I(new_n18072_), .ZN(new_n18073_));
  OAI22_X1   g17817(.A1(new_n6490_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n6775_), .ZN(new_n18074_));
  AOI21_X1   g17818(.A1(\b[41] ), .A2(new_n7719_), .B(new_n18074_), .ZN(new_n18075_));
  OAI21_X1   g17819(.A1(new_n6785_), .A2(new_n8585_), .B(new_n18075_), .ZN(new_n18076_));
  XOR2_X1    g17820(.A1(new_n18076_), .A2(\a[47] ), .Z(new_n18077_));
  NOR2_X1    g17821(.A1(new_n18073_), .A2(new_n18077_), .ZN(new_n18078_));
  NAND2_X1   g17822(.A1(new_n18073_), .A2(new_n18077_), .ZN(new_n18079_));
  INV_X1     g17823(.I(new_n18079_), .ZN(new_n18080_));
  NOR2_X1    g17824(.A1(new_n18080_), .A2(new_n18078_), .ZN(new_n18081_));
  XOR2_X1    g17825(.A1(new_n18081_), .A2(new_n18015_), .Z(new_n18082_));
  NOR2_X1    g17826(.A1(new_n17927_), .A2(new_n17860_), .ZN(new_n18083_));
  NOR2_X1    g17827(.A1(new_n18083_), .A2(new_n17925_), .ZN(new_n18084_));
  NOR2_X1    g17828(.A1(new_n18084_), .A2(new_n18082_), .ZN(new_n18085_));
  INV_X1     g17829(.I(new_n18085_), .ZN(new_n18086_));
  NAND2_X1   g17830(.A1(new_n18084_), .A2(new_n18082_), .ZN(new_n18087_));
  NAND2_X1   g17831(.A1(new_n18086_), .A2(new_n18087_), .ZN(new_n18088_));
  XOR2_X1    g17832(.A1(new_n18088_), .A2(new_n18013_), .Z(new_n18089_));
  AOI21_X1   g17833(.A1(new_n17858_), .A2(new_n17935_), .B(new_n17934_), .ZN(new_n18090_));
  OAI22_X1   g17834(.A1(new_n5852_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n5857_), .ZN(new_n18091_));
  AOI21_X1   g17835(.A1(\b[47] ), .A2(new_n6115_), .B(new_n18091_), .ZN(new_n18092_));
  OAI21_X1   g17836(.A1(new_n9050_), .A2(new_n5861_), .B(new_n18092_), .ZN(new_n18093_));
  XOR2_X1    g17837(.A1(new_n18093_), .A2(\a[41] ), .Z(new_n18094_));
  NOR2_X1    g17838(.A1(new_n18090_), .A2(new_n18094_), .ZN(new_n18095_));
  NAND2_X1   g17839(.A1(new_n18090_), .A2(new_n18094_), .ZN(new_n18096_));
  INV_X1     g17840(.I(new_n18096_), .ZN(new_n18097_));
  NOR2_X1    g17841(.A1(new_n18097_), .A2(new_n18095_), .ZN(new_n18098_));
  XOR2_X1    g17842(.A1(new_n18098_), .A2(new_n18089_), .Z(new_n18099_));
  INV_X1     g17843(.I(new_n17945_), .ZN(new_n18100_));
  AOI21_X1   g17844(.A1(new_n17938_), .A2(new_n17946_), .B(new_n18100_), .ZN(new_n18101_));
  XOR2_X1    g17845(.A1(new_n18099_), .A2(new_n18101_), .Z(new_n18102_));
  XOR2_X1    g17846(.A1(new_n18102_), .A2(new_n18008_), .Z(new_n18103_));
  AOI22_X1   g17847(.A1(new_n4918_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n4921_), .ZN(new_n18104_));
  OAI21_X1   g17848(.A1(new_n9376_), .A2(new_n6099_), .B(new_n18104_), .ZN(new_n18105_));
  AOI21_X1   g17849(.A1(new_n9979_), .A2(new_n4699_), .B(new_n18105_), .ZN(new_n18106_));
  XOR2_X1    g17850(.A1(new_n18106_), .A2(new_n4446_), .Z(new_n18107_));
  NOR2_X1    g17851(.A1(new_n18103_), .A2(new_n18107_), .ZN(new_n18108_));
  NAND2_X1   g17852(.A1(new_n18103_), .A2(new_n18107_), .ZN(new_n18109_));
  INV_X1     g17853(.I(new_n18109_), .ZN(new_n18110_));
  NOR2_X1    g17854(.A1(new_n18110_), .A2(new_n18108_), .ZN(new_n18111_));
  XOR2_X1    g17855(.A1(new_n18111_), .A2(new_n18004_), .Z(new_n18112_));
  NOR2_X1    g17856(.A1(new_n18112_), .A2(new_n18002_), .ZN(new_n18113_));
  INV_X1     g17857(.I(new_n18113_), .ZN(new_n18114_));
  NAND2_X1   g17858(.A1(new_n18112_), .A2(new_n18002_), .ZN(new_n18115_));
  NAND2_X1   g17859(.A1(new_n18114_), .A2(new_n18115_), .ZN(new_n18116_));
  XOR2_X1    g17860(.A1(new_n18116_), .A2(new_n18000_), .Z(new_n18117_));
  OR2_X2     g17861(.A1(new_n18117_), .A2(new_n17996_), .Z(new_n18118_));
  NAND2_X1   g17862(.A1(new_n18117_), .A2(new_n17996_), .ZN(new_n18119_));
  NAND2_X1   g17863(.A1(new_n18118_), .A2(new_n18119_), .ZN(new_n18120_));
  XNOR2_X1   g17864(.A1(new_n18120_), .A2(new_n17995_), .ZN(new_n18121_));
  NAND2_X1   g17865(.A1(new_n18121_), .A2(new_n17991_), .ZN(new_n18122_));
  NOR2_X1    g17866(.A1(new_n18121_), .A2(new_n17991_), .ZN(new_n18123_));
  INV_X1     g17867(.I(new_n18123_), .ZN(new_n18124_));
  NAND2_X1   g17868(.A1(new_n18124_), .A2(new_n18122_), .ZN(new_n18125_));
  XOR2_X1    g17869(.A1(new_n18125_), .A2(new_n17990_), .Z(new_n18126_));
  AOI21_X1   g17870(.A1(new_n17664_), .A2(new_n17500_), .B(new_n17661_), .ZN(new_n18127_));
  OAI21_X1   g17871(.A1(new_n17655_), .A2(new_n18127_), .B(new_n17665_), .ZN(new_n18128_));
  INV_X1     g17872(.I(new_n17818_), .ZN(new_n18129_));
  OAI21_X1   g17873(.A1(new_n18128_), .A2(new_n18129_), .B(new_n17817_), .ZN(new_n18130_));
  AOI21_X1   g17874(.A1(new_n18130_), .A2(new_n17983_), .B(new_n17981_), .ZN(new_n18131_));
  NOR2_X1    g17875(.A1(new_n18131_), .A2(new_n18126_), .ZN(new_n18132_));
  INV_X1     g17876(.I(new_n18126_), .ZN(new_n18133_));
  OAI21_X1   g17877(.A1(new_n17985_), .A2(new_n17984_), .B(new_n17982_), .ZN(new_n18134_));
  NOR2_X1    g17878(.A1(new_n18134_), .A2(new_n18133_), .ZN(new_n18135_));
  NOR2_X1    g17879(.A1(new_n18132_), .A2(new_n18135_), .ZN(new_n18136_));
  XOR2_X1    g17880(.A1(new_n18136_), .A2(new_n17987_), .Z(\f[88] ));
  AOI21_X1   g17881(.A1(new_n18134_), .A2(new_n18133_), .B(new_n17987_), .ZN(new_n18138_));
  NOR2_X1    g17882(.A1(new_n18138_), .A2(new_n18135_), .ZN(new_n18139_));
  OAI21_X1   g17883(.A1(new_n17990_), .A2(new_n18123_), .B(new_n18122_), .ZN(new_n18140_));
  AOI22_X1   g17884(.A1(new_n13460_), .A2(new_n2722_), .B1(\b[63] ), .B2(new_n2906_), .ZN(new_n18141_));
  AOI22_X1   g17885(.A1(new_n3267_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n3270_), .ZN(new_n18142_));
  OAI21_X1   g17886(.A1(new_n12147_), .A2(new_n3475_), .B(new_n18142_), .ZN(new_n18143_));
  AOI21_X1   g17887(.A1(new_n13444_), .A2(new_n3273_), .B(new_n18143_), .ZN(new_n18144_));
  XOR2_X1    g17888(.A1(new_n18144_), .A2(new_n3264_), .Z(new_n18145_));
  OAI21_X1   g17889(.A1(new_n18000_), .A2(new_n18113_), .B(new_n18115_), .ZN(new_n18146_));
  INV_X1     g17890(.I(new_n18146_), .ZN(new_n18147_));
  OAI22_X1   g17891(.A1(new_n11195_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n12151_), .ZN(new_n18148_));
  AOI21_X1   g17892(.A1(\b[57] ), .A2(new_n4053_), .B(new_n18148_), .ZN(new_n18149_));
  OAI21_X1   g17893(.A1(new_n12203_), .A2(new_n4727_), .B(new_n18149_), .ZN(new_n18150_));
  XOR2_X1    g17894(.A1(new_n18150_), .A2(\a[32] ), .Z(new_n18151_));
  AOI21_X1   g17895(.A1(new_n18004_), .A2(new_n18109_), .B(new_n18108_), .ZN(new_n18152_));
  AOI22_X1   g17896(.A1(new_n4918_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n4921_), .ZN(new_n18153_));
  OAI21_X1   g17897(.A1(new_n9942_), .A2(new_n6099_), .B(new_n18153_), .ZN(new_n18154_));
  AOI21_X1   g17898(.A1(new_n10318_), .A2(new_n4699_), .B(new_n18154_), .ZN(new_n18155_));
  XOR2_X1    g17899(.A1(new_n18155_), .A2(new_n4446_), .Z(new_n18156_));
  INV_X1     g17900(.I(new_n18008_), .ZN(new_n18157_));
  NOR2_X1    g17901(.A1(new_n18099_), .A2(new_n18101_), .ZN(new_n18158_));
  NAND2_X1   g17902(.A1(new_n18099_), .A2(new_n18101_), .ZN(new_n18159_));
  AOI21_X1   g17903(.A1(new_n18157_), .A2(new_n18159_), .B(new_n18158_), .ZN(new_n18160_));
  INV_X1     g17904(.I(new_n18160_), .ZN(new_n18161_));
  OAI22_X1   g17905(.A1(new_n9376_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n9032_), .ZN(new_n18162_));
  AOI21_X1   g17906(.A1(\b[51] ), .A2(new_n5420_), .B(new_n18162_), .ZN(new_n18163_));
  OAI21_X1   g17907(.A1(new_n9385_), .A2(new_n6124_), .B(new_n18163_), .ZN(new_n18164_));
  XOR2_X1    g17908(.A1(new_n18164_), .A2(new_n5162_), .Z(new_n18165_));
  AOI22_X1   g17909(.A1(new_n6108_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n6111_), .ZN(new_n18166_));
  OAI21_X1   g17910(.A1(new_n8127_), .A2(new_n7708_), .B(new_n18166_), .ZN(new_n18167_));
  AOI21_X1   g17911(.A1(new_n9684_), .A2(new_n6105_), .B(new_n18167_), .ZN(new_n18168_));
  XOR2_X1    g17912(.A1(new_n18168_), .A2(new_n5849_), .Z(new_n18169_));
  AOI22_X1   g17913(.A1(new_n7403_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n7408_), .ZN(new_n18170_));
  OAI21_X1   g17914(.A1(new_n6490_), .A2(new_n9488_), .B(new_n18170_), .ZN(new_n18171_));
  AOI21_X1   g17915(.A1(new_n7906_), .A2(new_n7414_), .B(new_n18171_), .ZN(new_n18172_));
  XOR2_X1    g17916(.A1(new_n18172_), .A2(new_n7410_), .Z(new_n18173_));
  INV_X1     g17917(.I(new_n18173_), .ZN(new_n18174_));
  OAI21_X1   g17918(.A1(new_n18019_), .A2(new_n18068_), .B(new_n18070_), .ZN(new_n18175_));
  INV_X1     g17919(.I(new_n18175_), .ZN(new_n18176_));
  AOI22_X1   g17920(.A1(new_n9125_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n9123_), .ZN(new_n18177_));
  OAI21_X1   g17921(.A1(new_n4886_), .A2(new_n9470_), .B(new_n18177_), .ZN(new_n18178_));
  AOI21_X1   g17922(.A1(new_n5351_), .A2(new_n9129_), .B(new_n18178_), .ZN(new_n18179_));
  XOR2_X1    g17923(.A1(new_n18179_), .A2(new_n9133_), .Z(new_n18180_));
  AOI21_X1   g17924(.A1(new_n18026_), .A2(new_n18054_), .B(new_n18052_), .ZN(new_n18181_));
  INV_X1     g17925(.I(new_n18181_), .ZN(new_n18182_));
  OAI22_X1   g17926(.A1(new_n11298_), .A2(new_n4666_), .B1(new_n4639_), .B2(new_n11297_), .ZN(new_n18183_));
  AOI21_X1   g17927(.A1(\b[33] ), .A2(new_n11296_), .B(new_n18183_), .ZN(new_n18184_));
  OAI21_X1   g17928(.A1(new_n4676_), .A2(new_n10069_), .B(new_n18184_), .ZN(new_n18185_));
  XOR2_X1    g17929(.A1(new_n18185_), .A2(\a[56] ), .Z(new_n18186_));
  AOI22_X1   g17930(.A1(new_n10981_), .A2(\b[32] ), .B1(new_n10979_), .B2(\b[31] ), .ZN(new_n18187_));
  OAI21_X1   g17931(.A1(new_n3624_), .A2(new_n11306_), .B(new_n18187_), .ZN(new_n18188_));
  AOI21_X1   g17932(.A1(new_n4030_), .A2(new_n10984_), .B(new_n18188_), .ZN(new_n18189_));
  XOR2_X1    g17933(.A1(new_n18189_), .A2(new_n10989_), .Z(new_n18190_));
  AOI21_X1   g17934(.A1(new_n18031_), .A2(new_n18035_), .B(new_n18036_), .ZN(new_n18191_));
  INV_X1     g17935(.I(new_n18191_), .ZN(new_n18192_));
  AOI22_X1   g17936(.A1(new_n11926_), .A2(\b[29] ), .B1(new_n11924_), .B2(\b[28] ), .ZN(new_n18193_));
  OAI21_X1   g17937(.A1(new_n3158_), .A2(new_n12317_), .B(new_n18193_), .ZN(new_n18194_));
  AOI21_X1   g17938(.A1(new_n4188_), .A2(new_n11929_), .B(new_n18194_), .ZN(new_n18195_));
  XOR2_X1    g17939(.A1(new_n18195_), .A2(\a[62] ), .Z(new_n18196_));
  INV_X1     g17940(.I(new_n18034_), .ZN(new_n18197_));
  AOI22_X1   g17941(.A1(new_n12922_), .A2(\b[26] ), .B1(\b[25] ), .B2(new_n12923_), .ZN(new_n18198_));
  NAND2_X1   g17942(.A1(new_n18197_), .A2(new_n18198_), .ZN(new_n18199_));
  INV_X1     g17943(.I(new_n18198_), .ZN(new_n18200_));
  NAND2_X1   g17944(.A1(new_n18200_), .A2(new_n18034_), .ZN(new_n18201_));
  NAND2_X1   g17945(.A1(new_n18199_), .A2(new_n18201_), .ZN(new_n18202_));
  XNOR2_X1   g17946(.A1(new_n18196_), .A2(new_n18202_), .ZN(new_n18203_));
  NOR2_X1    g17947(.A1(new_n18203_), .A2(new_n18192_), .ZN(new_n18204_));
  INV_X1     g17948(.I(new_n18204_), .ZN(new_n18205_));
  NAND2_X1   g17949(.A1(new_n18203_), .A2(new_n18192_), .ZN(new_n18206_));
  NAND2_X1   g17950(.A1(new_n18205_), .A2(new_n18206_), .ZN(new_n18207_));
  XOR2_X1    g17951(.A1(new_n18207_), .A2(new_n18190_), .Z(new_n18208_));
  AOI21_X1   g17952(.A1(new_n18027_), .A2(new_n18046_), .B(new_n18045_), .ZN(new_n18209_));
  XOR2_X1    g17953(.A1(new_n18208_), .A2(new_n18209_), .Z(new_n18210_));
  XOR2_X1    g17954(.A1(new_n18210_), .A2(new_n18186_), .Z(new_n18211_));
  NOR2_X1    g17955(.A1(new_n18182_), .A2(new_n18211_), .ZN(new_n18212_));
  INV_X1     g17956(.I(new_n18212_), .ZN(new_n18213_));
  NAND2_X1   g17957(.A1(new_n18182_), .A2(new_n18211_), .ZN(new_n18214_));
  NAND2_X1   g17958(.A1(new_n18213_), .A2(new_n18214_), .ZN(new_n18215_));
  XNOR2_X1   g17959(.A1(new_n18215_), .A2(new_n18180_), .ZN(new_n18216_));
  INV_X1     g17960(.I(new_n18216_), .ZN(new_n18217_));
  OAI22_X1   g17961(.A1(new_n9461_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n9462_), .ZN(new_n18218_));
  AOI21_X1   g17962(.A1(\b[39] ), .A2(new_n8575_), .B(new_n18218_), .ZN(new_n18219_));
  OAI21_X1   g17963(.A1(new_n6299_), .A2(new_n9460_), .B(new_n18219_), .ZN(new_n18220_));
  XOR2_X1    g17964(.A1(new_n18220_), .A2(\a[50] ), .Z(new_n18221_));
  INV_X1     g17965(.I(new_n18056_), .ZN(new_n18222_));
  AOI21_X1   g17966(.A1(new_n18222_), .A2(new_n18065_), .B(new_n18063_), .ZN(new_n18223_));
  NOR2_X1    g17967(.A1(new_n18221_), .A2(new_n18223_), .ZN(new_n18224_));
  INV_X1     g17968(.I(new_n18224_), .ZN(new_n18225_));
  NAND2_X1   g17969(.A1(new_n18221_), .A2(new_n18223_), .ZN(new_n18226_));
  NAND2_X1   g17970(.A1(new_n18225_), .A2(new_n18226_), .ZN(new_n18227_));
  XOR2_X1    g17971(.A1(new_n18227_), .A2(new_n18217_), .Z(new_n18228_));
  NOR2_X1    g17972(.A1(new_n18228_), .A2(new_n18176_), .ZN(new_n18229_));
  INV_X1     g17973(.I(new_n18229_), .ZN(new_n18230_));
  NAND2_X1   g17974(.A1(new_n18228_), .A2(new_n18176_), .ZN(new_n18231_));
  NAND2_X1   g17975(.A1(new_n18230_), .A2(new_n18231_), .ZN(new_n18232_));
  XOR2_X1    g17976(.A1(new_n18232_), .A2(new_n18174_), .Z(new_n18233_));
  AOI22_X1   g17977(.A1(new_n6569_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n6574_), .ZN(new_n18234_));
  OAI21_X1   g17978(.A1(new_n7096_), .A2(new_n8565_), .B(new_n18234_), .ZN(new_n18235_));
  AOI21_X1   g17979(.A1(new_n7649_), .A2(new_n6579_), .B(new_n18235_), .ZN(new_n18236_));
  XOR2_X1    g17980(.A1(new_n18236_), .A2(new_n6567_), .Z(new_n18237_));
  NOR2_X1    g17981(.A1(new_n18080_), .A2(new_n18015_), .ZN(new_n18238_));
  NOR2_X1    g17982(.A1(new_n18238_), .A2(new_n18078_), .ZN(new_n18239_));
  NOR2_X1    g17983(.A1(new_n18239_), .A2(new_n18237_), .ZN(new_n18240_));
  AND2_X2    g17984(.A1(new_n18239_), .A2(new_n18237_), .Z(new_n18241_));
  NOR2_X1    g17985(.A1(new_n18241_), .A2(new_n18240_), .ZN(new_n18242_));
  XOR2_X1    g17986(.A1(new_n18242_), .A2(new_n18233_), .Z(new_n18243_));
  AOI21_X1   g17987(.A1(new_n18013_), .A2(new_n18087_), .B(new_n18085_), .ZN(new_n18244_));
  NOR2_X1    g17988(.A1(new_n18243_), .A2(new_n18244_), .ZN(new_n18245_));
  INV_X1     g17989(.I(new_n18245_), .ZN(new_n18246_));
  NAND2_X1   g17990(.A1(new_n18243_), .A2(new_n18244_), .ZN(new_n18247_));
  NAND2_X1   g17991(.A1(new_n18246_), .A2(new_n18247_), .ZN(new_n18248_));
  XOR2_X1    g17992(.A1(new_n18248_), .A2(new_n18169_), .Z(new_n18249_));
  INV_X1     g17993(.I(new_n18249_), .ZN(new_n18250_));
  NOR2_X1    g17994(.A1(new_n18097_), .A2(new_n18089_), .ZN(new_n18251_));
  NOR2_X1    g17995(.A1(new_n18251_), .A2(new_n18095_), .ZN(new_n18252_));
  NOR2_X1    g17996(.A1(new_n18250_), .A2(new_n18252_), .ZN(new_n18253_));
  INV_X1     g17997(.I(new_n18253_), .ZN(new_n18254_));
  NAND2_X1   g17998(.A1(new_n18250_), .A2(new_n18252_), .ZN(new_n18255_));
  NAND2_X1   g17999(.A1(new_n18254_), .A2(new_n18255_), .ZN(new_n18256_));
  XNOR2_X1   g18000(.A1(new_n18256_), .A2(new_n18165_), .ZN(new_n18257_));
  NOR2_X1    g18001(.A1(new_n18257_), .A2(new_n18161_), .ZN(new_n18258_));
  NAND2_X1   g18002(.A1(new_n18257_), .A2(new_n18161_), .ZN(new_n18259_));
  INV_X1     g18003(.I(new_n18259_), .ZN(new_n18260_));
  NOR2_X1    g18004(.A1(new_n18260_), .A2(new_n18258_), .ZN(new_n18261_));
  XOR2_X1    g18005(.A1(new_n18261_), .A2(new_n18156_), .Z(new_n18262_));
  NOR2_X1    g18006(.A1(new_n18262_), .A2(new_n18152_), .ZN(new_n18263_));
  NAND2_X1   g18007(.A1(new_n18262_), .A2(new_n18152_), .ZN(new_n18264_));
  INV_X1     g18008(.I(new_n18264_), .ZN(new_n18265_));
  NOR2_X1    g18009(.A1(new_n18265_), .A2(new_n18263_), .ZN(new_n18266_));
  XOR2_X1    g18010(.A1(new_n18266_), .A2(new_n18151_), .Z(new_n18267_));
  NOR2_X1    g18011(.A1(new_n18267_), .A2(new_n18147_), .ZN(new_n18268_));
  INV_X1     g18012(.I(new_n18268_), .ZN(new_n18269_));
  NAND2_X1   g18013(.A1(new_n18267_), .A2(new_n18147_), .ZN(new_n18270_));
  NAND2_X1   g18014(.A1(new_n18269_), .A2(new_n18270_), .ZN(new_n18271_));
  XOR2_X1    g18015(.A1(new_n18271_), .A2(new_n18145_), .Z(new_n18272_));
  XOR2_X1    g18016(.A1(new_n18272_), .A2(new_n18141_), .Z(new_n18273_));
  NAND2_X1   g18017(.A1(new_n18118_), .A2(new_n17995_), .ZN(new_n18274_));
  NAND2_X1   g18018(.A1(new_n18274_), .A2(new_n18119_), .ZN(new_n18275_));
  XOR2_X1    g18019(.A1(new_n18275_), .A2(\a[26] ), .Z(new_n18276_));
  XOR2_X1    g18020(.A1(new_n18273_), .A2(new_n18276_), .Z(new_n18277_));
  NOR2_X1    g18021(.A1(new_n18277_), .A2(new_n18140_), .ZN(new_n18278_));
  NAND2_X1   g18022(.A1(new_n18277_), .A2(new_n18140_), .ZN(new_n18279_));
  INV_X1     g18023(.I(new_n18279_), .ZN(new_n18280_));
  NOR2_X1    g18024(.A1(new_n18280_), .A2(new_n18278_), .ZN(new_n18281_));
  XOR2_X1    g18025(.A1(new_n18139_), .A2(new_n18281_), .Z(\f[89] ));
  NAND2_X1   g18026(.A1(new_n18131_), .A2(new_n18126_), .ZN(new_n18283_));
  INV_X1     g18027(.I(new_n17987_), .ZN(new_n18284_));
  OAI21_X1   g18028(.A1(new_n18131_), .A2(new_n18126_), .B(new_n18284_), .ZN(new_n18285_));
  AOI21_X1   g18029(.A1(new_n18285_), .A2(new_n18283_), .B(new_n18278_), .ZN(new_n18286_));
  NOR2_X1    g18030(.A1(new_n18272_), .A2(new_n18275_), .ZN(new_n18287_));
  XOR2_X1    g18031(.A1(new_n18141_), .A2(new_n2714_), .Z(new_n18288_));
  NOR2_X1    g18032(.A1(new_n18287_), .A2(new_n18288_), .ZN(new_n18289_));
  AOI21_X1   g18033(.A1(new_n18272_), .A2(new_n18275_), .B(new_n18289_), .ZN(new_n18290_));
  INV_X1     g18034(.I(new_n18290_), .ZN(new_n18291_));
  INV_X1     g18035(.I(new_n18145_), .ZN(new_n18292_));
  AOI21_X1   g18036(.A1(new_n18292_), .A2(new_n18270_), .B(new_n18268_), .ZN(new_n18293_));
  INV_X1     g18037(.I(new_n18293_), .ZN(new_n18294_));
  AOI22_X1   g18038(.A1(new_n3267_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n3270_), .ZN(new_n18295_));
  OAI21_X1   g18039(.A1(new_n12148_), .A2(new_n3475_), .B(new_n18295_), .ZN(new_n18296_));
  AOI21_X1   g18040(.A1(new_n12811_), .A2(new_n3273_), .B(new_n18296_), .ZN(new_n18297_));
  XOR2_X1    g18041(.A1(new_n18297_), .A2(new_n3264_), .Z(new_n18298_));
  OAI21_X1   g18042(.A1(new_n18156_), .A2(new_n18258_), .B(new_n18259_), .ZN(new_n18299_));
  AOI21_X1   g18043(.A1(new_n18165_), .A2(new_n18255_), .B(new_n18253_), .ZN(new_n18300_));
  INV_X1     g18044(.I(new_n18300_), .ZN(new_n18301_));
  AOI22_X1   g18045(.A1(new_n5155_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n5160_), .ZN(new_n18302_));
  OAI21_X1   g18046(.A1(new_n9032_), .A2(new_n6877_), .B(new_n18302_), .ZN(new_n18303_));
  AOI21_X1   g18047(.A1(new_n10884_), .A2(new_n5166_), .B(new_n18303_), .ZN(new_n18304_));
  XOR2_X1    g18048(.A1(new_n18304_), .A2(new_n5162_), .Z(new_n18305_));
  INV_X1     g18049(.I(new_n18169_), .ZN(new_n18306_));
  AOI21_X1   g18050(.A1(new_n18306_), .A2(new_n18247_), .B(new_n18245_), .ZN(new_n18307_));
  INV_X1     g18051(.I(new_n18307_), .ZN(new_n18308_));
  AOI21_X1   g18052(.A1(new_n18174_), .A2(new_n18231_), .B(new_n18229_), .ZN(new_n18309_));
  AOI21_X1   g18053(.A1(new_n18217_), .A2(new_n18226_), .B(new_n18224_), .ZN(new_n18310_));
  OAI21_X1   g18054(.A1(new_n18180_), .A2(new_n18212_), .B(new_n18214_), .ZN(new_n18311_));
  OAI21_X1   g18055(.A1(new_n18190_), .A2(new_n18204_), .B(new_n18206_), .ZN(new_n18312_));
  AOI22_X1   g18056(.A1(new_n10981_), .A2(\b[33] ), .B1(new_n10979_), .B2(\b[32] ), .ZN(new_n18313_));
  OAI21_X1   g18057(.A1(new_n4022_), .A2(new_n11306_), .B(new_n18313_), .ZN(new_n18314_));
  AOI21_X1   g18058(.A1(new_n4223_), .A2(new_n10984_), .B(new_n18314_), .ZN(new_n18315_));
  XOR2_X1    g18059(.A1(new_n18315_), .A2(new_n10989_), .Z(new_n18316_));
  NAND2_X1   g18060(.A1(new_n18196_), .A2(new_n18199_), .ZN(new_n18317_));
  NAND2_X1   g18061(.A1(new_n18317_), .A2(new_n18201_), .ZN(new_n18318_));
  INV_X1     g18062(.I(new_n18318_), .ZN(new_n18319_));
  AOI22_X1   g18063(.A1(new_n11926_), .A2(\b[30] ), .B1(new_n11924_), .B2(\b[29] ), .ZN(new_n18320_));
  OAI21_X1   g18064(.A1(new_n3185_), .A2(new_n12317_), .B(new_n18320_), .ZN(new_n18321_));
  AOI21_X1   g18065(.A1(new_n4230_), .A2(new_n11929_), .B(new_n18321_), .ZN(new_n18322_));
  XOR2_X1    g18066(.A1(new_n18322_), .A2(new_n12312_), .Z(new_n18323_));
  INV_X1     g18067(.I(new_n18323_), .ZN(new_n18324_));
  AOI22_X1   g18068(.A1(new_n12922_), .A2(\b[27] ), .B1(\b[26] ), .B2(new_n12923_), .ZN(new_n18325_));
  INV_X1     g18069(.I(new_n18325_), .ZN(new_n18326_));
  NOR2_X1    g18070(.A1(new_n18326_), .A2(new_n2714_), .ZN(new_n18327_));
  NOR2_X1    g18071(.A1(new_n18325_), .A2(\a[26] ), .ZN(new_n18328_));
  NOR2_X1    g18072(.A1(new_n18327_), .A2(new_n18328_), .ZN(new_n18329_));
  XOR2_X1    g18073(.A1(new_n18329_), .A2(new_n18198_), .Z(new_n18330_));
  NOR2_X1    g18074(.A1(new_n18324_), .A2(new_n18330_), .ZN(new_n18331_));
  NAND2_X1   g18075(.A1(new_n18324_), .A2(new_n18330_), .ZN(new_n18332_));
  INV_X1     g18076(.I(new_n18332_), .ZN(new_n18333_));
  NOR2_X1    g18077(.A1(new_n18333_), .A2(new_n18331_), .ZN(new_n18334_));
  XOR2_X1    g18078(.A1(new_n18334_), .A2(new_n18319_), .Z(new_n18335_));
  NOR2_X1    g18079(.A1(new_n18335_), .A2(new_n18316_), .ZN(new_n18336_));
  NAND2_X1   g18080(.A1(new_n18335_), .A2(new_n18316_), .ZN(new_n18337_));
  INV_X1     g18081(.I(new_n18337_), .ZN(new_n18338_));
  NOR2_X1    g18082(.A1(new_n18338_), .A2(new_n18336_), .ZN(new_n18339_));
  XOR2_X1    g18083(.A1(new_n18339_), .A2(new_n18312_), .Z(new_n18340_));
  AOI22_X1   g18084(.A1(new_n10064_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n10062_), .ZN(new_n18341_));
  OAI21_X1   g18085(.A1(new_n4639_), .A2(new_n10399_), .B(new_n18341_), .ZN(new_n18342_));
  AOI21_X1   g18086(.A1(new_n5594_), .A2(new_n10068_), .B(new_n18342_), .ZN(new_n18343_));
  XOR2_X1    g18087(.A1(new_n18343_), .A2(new_n10057_), .Z(new_n18344_));
  INV_X1     g18088(.I(new_n18208_), .ZN(new_n18345_));
  NOR2_X1    g18089(.A1(new_n18345_), .A2(new_n18209_), .ZN(new_n18346_));
  AOI21_X1   g18090(.A1(new_n18345_), .A2(new_n18209_), .B(new_n18186_), .ZN(new_n18347_));
  NOR2_X1    g18091(.A1(new_n18347_), .A2(new_n18346_), .ZN(new_n18348_));
  NOR2_X1    g18092(.A1(new_n18348_), .A2(new_n18344_), .ZN(new_n18349_));
  NAND2_X1   g18093(.A1(new_n18348_), .A2(new_n18344_), .ZN(new_n18350_));
  INV_X1     g18094(.I(new_n18350_), .ZN(new_n18351_));
  NOR2_X1    g18095(.A1(new_n18351_), .A2(new_n18349_), .ZN(new_n18352_));
  XOR2_X1    g18096(.A1(new_n18352_), .A2(new_n18340_), .Z(new_n18353_));
  AOI22_X1   g18097(.A1(new_n9125_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n9123_), .ZN(new_n18354_));
  OAI21_X1   g18098(.A1(new_n5312_), .A2(new_n9470_), .B(new_n18354_), .ZN(new_n18355_));
  AOI21_X1   g18099(.A1(new_n6310_), .A2(new_n9129_), .B(new_n18355_), .ZN(new_n18356_));
  XOR2_X1    g18100(.A1(new_n18356_), .A2(\a[53] ), .Z(new_n18357_));
  NAND2_X1   g18101(.A1(new_n18353_), .A2(new_n18357_), .ZN(new_n18358_));
  OR2_X2     g18102(.A1(new_n18353_), .A2(new_n18357_), .Z(new_n18359_));
  NAND2_X1   g18103(.A1(new_n18359_), .A2(new_n18358_), .ZN(new_n18360_));
  XNOR2_X1   g18104(.A1(new_n18360_), .A2(new_n18311_), .ZN(new_n18361_));
  INV_X1     g18105(.I(new_n18361_), .ZN(new_n18362_));
  AOI22_X1   g18106(.A1(new_n8241_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n8246_), .ZN(new_n18363_));
  OAI21_X1   g18107(.A1(new_n6284_), .A2(new_n9114_), .B(new_n18363_), .ZN(new_n18364_));
  AOI21_X1   g18108(.A1(new_n7106_), .A2(new_n8252_), .B(new_n18364_), .ZN(new_n18365_));
  XOR2_X1    g18109(.A1(new_n18365_), .A2(new_n8248_), .Z(new_n18366_));
  NOR2_X1    g18110(.A1(new_n18362_), .A2(new_n18366_), .ZN(new_n18367_));
  NAND2_X1   g18111(.A1(new_n18362_), .A2(new_n18366_), .ZN(new_n18368_));
  INV_X1     g18112(.I(new_n18368_), .ZN(new_n18369_));
  NOR2_X1    g18113(.A1(new_n18369_), .A2(new_n18367_), .ZN(new_n18370_));
  XOR2_X1    g18114(.A1(new_n18370_), .A2(new_n18310_), .Z(new_n18371_));
  AOI22_X1   g18115(.A1(new_n7403_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n7408_), .ZN(new_n18372_));
  OAI21_X1   g18116(.A1(new_n6775_), .A2(new_n9488_), .B(new_n18372_), .ZN(new_n18373_));
  AOI21_X1   g18117(.A1(new_n7926_), .A2(new_n7414_), .B(new_n18373_), .ZN(new_n18374_));
  XOR2_X1    g18118(.A1(new_n18374_), .A2(new_n7410_), .Z(new_n18375_));
  NOR2_X1    g18119(.A1(new_n18371_), .A2(new_n18375_), .ZN(new_n18376_));
  INV_X1     g18120(.I(new_n18376_), .ZN(new_n18377_));
  NAND2_X1   g18121(.A1(new_n18371_), .A2(new_n18375_), .ZN(new_n18378_));
  NAND2_X1   g18122(.A1(new_n18377_), .A2(new_n18378_), .ZN(new_n18379_));
  XOR2_X1    g18123(.A1(new_n18379_), .A2(new_n18309_), .Z(new_n18380_));
  AOI22_X1   g18124(.A1(new_n6569_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n6574_), .ZN(new_n18381_));
  OAI21_X1   g18125(.A1(new_n7617_), .A2(new_n8565_), .B(new_n18381_), .ZN(new_n18382_));
  AOI21_X1   g18126(.A1(new_n8792_), .A2(new_n6579_), .B(new_n18382_), .ZN(new_n18383_));
  XOR2_X1    g18127(.A1(new_n18383_), .A2(\a[44] ), .Z(new_n18384_));
  INV_X1     g18128(.I(new_n18240_), .ZN(new_n18385_));
  OAI21_X1   g18129(.A1(new_n18233_), .A2(new_n18241_), .B(new_n18385_), .ZN(new_n18386_));
  NAND2_X1   g18130(.A1(new_n18386_), .A2(new_n18384_), .ZN(new_n18387_));
  OR2_X2     g18131(.A1(new_n18386_), .A2(new_n18384_), .Z(new_n18388_));
  NAND2_X1   g18132(.A1(new_n18388_), .A2(new_n18387_), .ZN(new_n18389_));
  XNOR2_X1   g18133(.A1(new_n18380_), .A2(new_n18389_), .ZN(new_n18390_));
  INV_X1     g18134(.I(new_n18390_), .ZN(new_n18391_));
  AOI22_X1   g18135(.A1(new_n6108_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n6111_), .ZN(new_n18392_));
  OAI21_X1   g18136(.A1(new_n8168_), .A2(new_n7708_), .B(new_n18392_), .ZN(new_n18393_));
  AOI21_X1   g18137(.A1(new_n8783_), .A2(new_n6105_), .B(new_n18393_), .ZN(new_n18394_));
  XOR2_X1    g18138(.A1(new_n18394_), .A2(new_n5849_), .Z(new_n18395_));
  NOR2_X1    g18139(.A1(new_n18391_), .A2(new_n18395_), .ZN(new_n18396_));
  INV_X1     g18140(.I(new_n18396_), .ZN(new_n18397_));
  NAND2_X1   g18141(.A1(new_n18391_), .A2(new_n18395_), .ZN(new_n18398_));
  NAND2_X1   g18142(.A1(new_n18397_), .A2(new_n18398_), .ZN(new_n18399_));
  XOR2_X1    g18143(.A1(new_n18399_), .A2(new_n18308_), .Z(new_n18400_));
  NOR2_X1    g18144(.A1(new_n18400_), .A2(new_n18305_), .ZN(new_n18401_));
  NAND2_X1   g18145(.A1(new_n18400_), .A2(new_n18305_), .ZN(new_n18402_));
  INV_X1     g18146(.I(new_n18402_), .ZN(new_n18403_));
  NOR2_X1    g18147(.A1(new_n18403_), .A2(new_n18401_), .ZN(new_n18404_));
  XOR2_X1    g18148(.A1(new_n18404_), .A2(new_n18301_), .Z(new_n18405_));
  INV_X1     g18149(.I(new_n18405_), .ZN(new_n18406_));
  AOI22_X1   g18150(.A1(new_n4918_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n4921_), .ZN(new_n18407_));
  OAI21_X1   g18151(.A1(new_n9972_), .A2(new_n6099_), .B(new_n18407_), .ZN(new_n18408_));
  AOI21_X1   g18152(.A1(new_n10631_), .A2(new_n4699_), .B(new_n18408_), .ZN(new_n18409_));
  XOR2_X1    g18153(.A1(new_n18409_), .A2(new_n4446_), .Z(new_n18410_));
  NOR2_X1    g18154(.A1(new_n18406_), .A2(new_n18410_), .ZN(new_n18411_));
  NAND2_X1   g18155(.A1(new_n18406_), .A2(new_n18410_), .ZN(new_n18412_));
  INV_X1     g18156(.I(new_n18412_), .ZN(new_n18413_));
  NOR2_X1    g18157(.A1(new_n18413_), .A2(new_n18411_), .ZN(new_n18414_));
  XOR2_X1    g18158(.A1(new_n18414_), .A2(new_n18299_), .Z(new_n18415_));
  AOI22_X1   g18159(.A1(new_n3864_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n3869_), .ZN(new_n18416_));
  OAI21_X1   g18160(.A1(new_n11195_), .A2(new_n5410_), .B(new_n18416_), .ZN(new_n18417_));
  AOI21_X1   g18161(.A1(new_n11836_), .A2(new_n3872_), .B(new_n18417_), .ZN(new_n18418_));
  XOR2_X1    g18162(.A1(new_n18418_), .A2(new_n3876_), .Z(new_n18419_));
  NOR2_X1    g18163(.A1(new_n18265_), .A2(new_n18151_), .ZN(new_n18420_));
  NOR2_X1    g18164(.A1(new_n18420_), .A2(new_n18263_), .ZN(new_n18421_));
  NOR2_X1    g18165(.A1(new_n18421_), .A2(new_n18419_), .ZN(new_n18422_));
  INV_X1     g18166(.I(new_n18422_), .ZN(new_n18423_));
  NAND2_X1   g18167(.A1(new_n18421_), .A2(new_n18419_), .ZN(new_n18424_));
  NAND2_X1   g18168(.A1(new_n18423_), .A2(new_n18424_), .ZN(new_n18425_));
  XOR2_X1    g18169(.A1(new_n18425_), .A2(new_n18415_), .Z(new_n18426_));
  NOR2_X1    g18170(.A1(new_n18426_), .A2(new_n18298_), .ZN(new_n18427_));
  NAND2_X1   g18171(.A1(new_n18426_), .A2(new_n18298_), .ZN(new_n18428_));
  INV_X1     g18172(.I(new_n18428_), .ZN(new_n18429_));
  NOR2_X1    g18173(.A1(new_n18429_), .A2(new_n18427_), .ZN(new_n18430_));
  XOR2_X1    g18174(.A1(new_n18430_), .A2(new_n18294_), .Z(new_n18431_));
  NOR2_X1    g18175(.A1(new_n18291_), .A2(new_n18431_), .ZN(new_n18432_));
  INV_X1     g18176(.I(new_n18432_), .ZN(new_n18433_));
  NAND2_X1   g18177(.A1(new_n18291_), .A2(new_n18431_), .ZN(new_n18434_));
  AND2_X2    g18178(.A1(new_n18433_), .A2(new_n18434_), .Z(new_n18435_));
  INV_X1     g18179(.I(new_n18435_), .ZN(new_n18436_));
  NOR3_X1    g18180(.A1(new_n18286_), .A2(new_n18280_), .A3(new_n18436_), .ZN(new_n18437_));
  INV_X1     g18181(.I(new_n18278_), .ZN(new_n18438_));
  OAI21_X1   g18182(.A1(new_n18138_), .A2(new_n18135_), .B(new_n18438_), .ZN(new_n18439_));
  AOI21_X1   g18183(.A1(new_n18439_), .A2(new_n18279_), .B(new_n18435_), .ZN(new_n18440_));
  NOR2_X1    g18184(.A1(new_n18437_), .A2(new_n18440_), .ZN(\f[90] ));
  OAI22_X1   g18185(.A1(new_n3475_), .A2(new_n12796_), .B1(new_n3258_), .B2(new_n12800_), .ZN(new_n18442_));
  AOI21_X1   g18186(.A1(new_n13973_), .A2(new_n3273_), .B(new_n18442_), .ZN(new_n18443_));
  XOR2_X1    g18187(.A1(new_n18443_), .A2(new_n3264_), .Z(new_n18444_));
  INV_X1     g18188(.I(new_n18444_), .ZN(new_n18445_));
  AOI21_X1   g18189(.A1(new_n18415_), .A2(new_n18424_), .B(new_n18422_), .ZN(new_n18446_));
  INV_X1     g18190(.I(new_n18446_), .ZN(new_n18447_));
  OAI22_X1   g18191(.A1(new_n12147_), .A2(new_n4730_), .B1(new_n4729_), .B2(new_n12148_), .ZN(new_n18448_));
  AOI21_X1   g18192(.A1(\b[59] ), .A2(new_n4053_), .B(new_n18448_), .ZN(new_n18449_));
  OAI21_X1   g18193(.A1(new_n13110_), .A2(new_n4727_), .B(new_n18449_), .ZN(new_n18450_));
  XOR2_X1    g18194(.A1(new_n18450_), .A2(new_n3876_), .Z(new_n18451_));
  AOI21_X1   g18195(.A1(new_n18299_), .A2(new_n18412_), .B(new_n18411_), .ZN(new_n18452_));
  AOI22_X1   g18196(.A1(new_n4918_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n4921_), .ZN(new_n18453_));
  OAI21_X1   g18197(.A1(new_n10308_), .A2(new_n6099_), .B(new_n18453_), .ZN(new_n18454_));
  AOI21_X1   g18198(.A1(new_n12164_), .A2(new_n4699_), .B(new_n18454_), .ZN(new_n18455_));
  XOR2_X1    g18199(.A1(new_n18455_), .A2(new_n4446_), .Z(new_n18456_));
  AOI21_X1   g18200(.A1(new_n18301_), .A2(new_n18402_), .B(new_n18401_), .ZN(new_n18457_));
  INV_X1     g18201(.I(new_n18457_), .ZN(new_n18458_));
  AOI21_X1   g18202(.A1(new_n18308_), .A2(new_n18398_), .B(new_n18396_), .ZN(new_n18459_));
  INV_X1     g18203(.I(new_n18459_), .ZN(new_n18460_));
  AOI22_X1   g18204(.A1(new_n6108_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n6111_), .ZN(new_n18461_));
  OAI21_X1   g18205(.A1(new_n8500_), .A2(new_n7708_), .B(new_n18461_), .ZN(new_n18462_));
  AOI21_X1   g18206(.A1(new_n9987_), .A2(new_n6105_), .B(new_n18462_), .ZN(new_n18463_));
  XOR2_X1    g18207(.A1(new_n18463_), .A2(new_n5849_), .Z(new_n18464_));
  AOI22_X1   g18208(.A1(new_n7403_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n7408_), .ZN(new_n18465_));
  OAI21_X1   g18209(.A1(new_n7074_), .A2(new_n9488_), .B(new_n18465_), .ZN(new_n18466_));
  AOI21_X1   g18210(.A1(new_n9337_), .A2(new_n7414_), .B(new_n18466_), .ZN(new_n18467_));
  XOR2_X1    g18211(.A1(new_n18467_), .A2(new_n7410_), .Z(new_n18468_));
  INV_X1     g18212(.I(new_n18468_), .ZN(new_n18469_));
  INV_X1     g18213(.I(new_n18358_), .ZN(new_n18470_));
  AOI21_X1   g18214(.A1(new_n18311_), .A2(new_n18359_), .B(new_n18470_), .ZN(new_n18471_));
  AOI22_X1   g18215(.A1(new_n9125_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n9123_), .ZN(new_n18472_));
  OAI21_X1   g18216(.A1(new_n5341_), .A2(new_n9470_), .B(new_n18472_), .ZN(new_n18473_));
  AOI21_X1   g18217(.A1(new_n5793_), .A2(new_n9129_), .B(new_n18473_), .ZN(new_n18474_));
  XOR2_X1    g18218(.A1(new_n18474_), .A2(new_n9133_), .Z(new_n18475_));
  AOI21_X1   g18219(.A1(new_n18340_), .A2(new_n18350_), .B(new_n18349_), .ZN(new_n18476_));
  AOI22_X1   g18220(.A1(new_n10981_), .A2(\b[34] ), .B1(new_n10979_), .B2(\b[33] ), .ZN(new_n18477_));
  OAI21_X1   g18221(.A1(new_n4023_), .A2(new_n11306_), .B(new_n18477_), .ZN(new_n18478_));
  AOI21_X1   g18222(.A1(new_n5103_), .A2(new_n10984_), .B(new_n18478_), .ZN(new_n18479_));
  XOR2_X1    g18223(.A1(new_n18479_), .A2(new_n10989_), .Z(new_n18480_));
  AOI22_X1   g18224(.A1(new_n11926_), .A2(\b[31] ), .B1(new_n11924_), .B2(\b[30] ), .ZN(new_n18481_));
  OAI21_X1   g18225(.A1(new_n3592_), .A2(new_n12317_), .B(new_n18481_), .ZN(new_n18482_));
  AOI21_X1   g18226(.A1(new_n3796_), .A2(new_n11929_), .B(new_n18482_), .ZN(new_n18483_));
  XOR2_X1    g18227(.A1(new_n18483_), .A2(new_n12312_), .Z(new_n18484_));
  INV_X1     g18228(.I(new_n18328_), .ZN(new_n18485_));
  AOI21_X1   g18229(.A1(new_n18198_), .A2(new_n18485_), .B(new_n18327_), .ZN(new_n18486_));
  AOI22_X1   g18230(.A1(new_n12922_), .A2(\b[28] ), .B1(\b[27] ), .B2(new_n12923_), .ZN(new_n18487_));
  AND2_X2    g18231(.A1(new_n18486_), .A2(new_n18487_), .Z(new_n18488_));
  NOR2_X1    g18232(.A1(new_n18486_), .A2(new_n18487_), .ZN(new_n18489_));
  NOR2_X1    g18233(.A1(new_n18488_), .A2(new_n18489_), .ZN(new_n18490_));
  XNOR2_X1   g18234(.A1(new_n18484_), .A2(new_n18490_), .ZN(new_n18491_));
  INV_X1     g18235(.I(new_n18491_), .ZN(new_n18492_));
  OAI21_X1   g18236(.A1(new_n18319_), .A2(new_n18331_), .B(new_n18332_), .ZN(new_n18493_));
  INV_X1     g18237(.I(new_n18493_), .ZN(new_n18494_));
  NOR2_X1    g18238(.A1(new_n18492_), .A2(new_n18494_), .ZN(new_n18495_));
  NOR2_X1    g18239(.A1(new_n18491_), .A2(new_n18493_), .ZN(new_n18496_));
  NOR2_X1    g18240(.A1(new_n18495_), .A2(new_n18496_), .ZN(new_n18497_));
  XOR2_X1    g18241(.A1(new_n18497_), .A2(new_n18480_), .Z(new_n18498_));
  INV_X1     g18242(.I(new_n18498_), .ZN(new_n18499_));
  AOI21_X1   g18243(.A1(new_n18312_), .A2(new_n18337_), .B(new_n18336_), .ZN(new_n18500_));
  OAI22_X1   g18244(.A1(new_n11298_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n11297_), .ZN(new_n18501_));
  AOI21_X1   g18245(.A1(\b[35] ), .A2(new_n11296_), .B(new_n18501_), .ZN(new_n18502_));
  OAI21_X1   g18246(.A1(new_n5322_), .A2(new_n10069_), .B(new_n18502_), .ZN(new_n18503_));
  XOR2_X1    g18247(.A1(new_n18503_), .A2(\a[56] ), .Z(new_n18504_));
  NOR2_X1    g18248(.A1(new_n18504_), .A2(new_n18500_), .ZN(new_n18505_));
  INV_X1     g18249(.I(new_n18505_), .ZN(new_n18506_));
  NAND2_X1   g18250(.A1(new_n18504_), .A2(new_n18500_), .ZN(new_n18507_));
  NAND2_X1   g18251(.A1(new_n18506_), .A2(new_n18507_), .ZN(new_n18508_));
  XOR2_X1    g18252(.A1(new_n18508_), .A2(new_n18499_), .Z(new_n18509_));
  NOR2_X1    g18253(.A1(new_n18509_), .A2(new_n18476_), .ZN(new_n18510_));
  INV_X1     g18254(.I(new_n18510_), .ZN(new_n18511_));
  NAND2_X1   g18255(.A1(new_n18509_), .A2(new_n18476_), .ZN(new_n18512_));
  NAND2_X1   g18256(.A1(new_n18511_), .A2(new_n18512_), .ZN(new_n18513_));
  XOR2_X1    g18257(.A1(new_n18513_), .A2(new_n18475_), .Z(new_n18514_));
  INV_X1     g18258(.I(new_n18514_), .ZN(new_n18515_));
  OAI22_X1   g18259(.A1(new_n9461_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n9462_), .ZN(new_n18516_));
  AOI21_X1   g18260(.A1(\b[41] ), .A2(new_n8575_), .B(new_n18516_), .ZN(new_n18517_));
  OAI21_X1   g18261(.A1(new_n6785_), .A2(new_n9460_), .B(new_n18517_), .ZN(new_n18518_));
  XOR2_X1    g18262(.A1(new_n18518_), .A2(\a[50] ), .Z(new_n18519_));
  NOR2_X1    g18263(.A1(new_n18515_), .A2(new_n18519_), .ZN(new_n18520_));
  NAND2_X1   g18264(.A1(new_n18515_), .A2(new_n18519_), .ZN(new_n18521_));
  INV_X1     g18265(.I(new_n18521_), .ZN(new_n18522_));
  NOR2_X1    g18266(.A1(new_n18522_), .A2(new_n18520_), .ZN(new_n18523_));
  XOR2_X1    g18267(.A1(new_n18523_), .A2(new_n18471_), .Z(new_n18524_));
  NOR2_X1    g18268(.A1(new_n18369_), .A2(new_n18310_), .ZN(new_n18525_));
  NOR2_X1    g18269(.A1(new_n18525_), .A2(new_n18367_), .ZN(new_n18526_));
  NOR2_X1    g18270(.A1(new_n18524_), .A2(new_n18526_), .ZN(new_n18527_));
  INV_X1     g18271(.I(new_n18527_), .ZN(new_n18528_));
  NAND2_X1   g18272(.A1(new_n18524_), .A2(new_n18526_), .ZN(new_n18529_));
  NAND2_X1   g18273(.A1(new_n18528_), .A2(new_n18529_), .ZN(new_n18530_));
  XOR2_X1    g18274(.A1(new_n18530_), .A2(new_n18469_), .Z(new_n18531_));
  INV_X1     g18275(.I(new_n18309_), .ZN(new_n18532_));
  AOI21_X1   g18276(.A1(new_n18532_), .A2(new_n18378_), .B(new_n18376_), .ZN(new_n18533_));
  OAI22_X1   g18277(.A1(new_n7730_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n7731_), .ZN(new_n18534_));
  AOI21_X1   g18278(.A1(\b[47] ), .A2(new_n6887_), .B(new_n18534_), .ZN(new_n18535_));
  OAI21_X1   g18279(.A1(new_n9050_), .A2(new_n7728_), .B(new_n18535_), .ZN(new_n18536_));
  XOR2_X1    g18280(.A1(new_n18536_), .A2(\a[44] ), .Z(new_n18537_));
  NOR2_X1    g18281(.A1(new_n18533_), .A2(new_n18537_), .ZN(new_n18538_));
  NAND2_X1   g18282(.A1(new_n18533_), .A2(new_n18537_), .ZN(new_n18539_));
  INV_X1     g18283(.I(new_n18539_), .ZN(new_n18540_));
  NOR2_X1    g18284(.A1(new_n18540_), .A2(new_n18538_), .ZN(new_n18541_));
  XOR2_X1    g18285(.A1(new_n18541_), .A2(new_n18531_), .Z(new_n18542_));
  INV_X1     g18286(.I(new_n18387_), .ZN(new_n18543_));
  AOI21_X1   g18287(.A1(new_n18380_), .A2(new_n18388_), .B(new_n18543_), .ZN(new_n18544_));
  XOR2_X1    g18288(.A1(new_n18542_), .A2(new_n18544_), .Z(new_n18545_));
  XOR2_X1    g18289(.A1(new_n18545_), .A2(new_n18464_), .Z(new_n18546_));
  AOI22_X1   g18290(.A1(new_n5155_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n5160_), .ZN(new_n18547_));
  OAI21_X1   g18291(.A1(new_n9376_), .A2(new_n6877_), .B(new_n18547_), .ZN(new_n18548_));
  AOI21_X1   g18292(.A1(new_n9979_), .A2(new_n5166_), .B(new_n18548_), .ZN(new_n18549_));
  XOR2_X1    g18293(.A1(new_n18549_), .A2(new_n5162_), .Z(new_n18550_));
  NOR2_X1    g18294(.A1(new_n18546_), .A2(new_n18550_), .ZN(new_n18551_));
  NAND2_X1   g18295(.A1(new_n18546_), .A2(new_n18550_), .ZN(new_n18552_));
  INV_X1     g18296(.I(new_n18552_), .ZN(new_n18553_));
  NOR2_X1    g18297(.A1(new_n18553_), .A2(new_n18551_), .ZN(new_n18554_));
  XOR2_X1    g18298(.A1(new_n18554_), .A2(new_n18460_), .Z(new_n18555_));
  NOR2_X1    g18299(.A1(new_n18555_), .A2(new_n18458_), .ZN(new_n18556_));
  NAND2_X1   g18300(.A1(new_n18555_), .A2(new_n18458_), .ZN(new_n18557_));
  INV_X1     g18301(.I(new_n18557_), .ZN(new_n18558_));
  NOR2_X1    g18302(.A1(new_n18558_), .A2(new_n18556_), .ZN(new_n18559_));
  XOR2_X1    g18303(.A1(new_n18559_), .A2(new_n18456_), .Z(new_n18560_));
  OR2_X2     g18304(.A1(new_n18560_), .A2(new_n18452_), .Z(new_n18561_));
  NAND2_X1   g18305(.A1(new_n18560_), .A2(new_n18452_), .ZN(new_n18562_));
  NAND2_X1   g18306(.A1(new_n18561_), .A2(new_n18562_), .ZN(new_n18563_));
  XNOR2_X1   g18307(.A1(new_n18563_), .A2(new_n18451_), .ZN(new_n18564_));
  NOR2_X1    g18308(.A1(new_n18564_), .A2(new_n18447_), .ZN(new_n18565_));
  INV_X1     g18309(.I(new_n18565_), .ZN(new_n18566_));
  NAND2_X1   g18310(.A1(new_n18564_), .A2(new_n18447_), .ZN(new_n18567_));
  NAND2_X1   g18311(.A1(new_n18566_), .A2(new_n18567_), .ZN(new_n18568_));
  XOR2_X1    g18312(.A1(new_n18568_), .A2(new_n18445_), .Z(new_n18569_));
  INV_X1     g18313(.I(new_n18569_), .ZN(new_n18570_));
  AOI21_X1   g18314(.A1(new_n18294_), .A2(new_n18428_), .B(new_n18427_), .ZN(new_n18571_));
  OAI21_X1   g18315(.A1(new_n18437_), .A2(new_n18432_), .B(new_n18571_), .ZN(new_n18572_));
  NAND3_X1   g18316(.A1(new_n18439_), .A2(new_n18279_), .A3(new_n18435_), .ZN(new_n18573_));
  INV_X1     g18317(.I(new_n18571_), .ZN(new_n18574_));
  NAND3_X1   g18318(.A1(new_n18573_), .A2(new_n18433_), .A3(new_n18574_), .ZN(new_n18575_));
  NAND2_X1   g18319(.A1(new_n18572_), .A2(new_n18575_), .ZN(new_n18576_));
  XOR2_X1    g18320(.A1(new_n18576_), .A2(new_n18570_), .Z(\f[91] ));
  AOI21_X1   g18321(.A1(new_n18573_), .A2(new_n18433_), .B(new_n18574_), .ZN(new_n18578_));
  OAI21_X1   g18322(.A1(new_n18569_), .A2(new_n18578_), .B(new_n18575_), .ZN(new_n18579_));
  OAI21_X1   g18323(.A1(new_n18444_), .A2(new_n18565_), .B(new_n18567_), .ZN(new_n18580_));
  AOI22_X1   g18324(.A1(new_n13460_), .A2(new_n3273_), .B1(\b[63] ), .B2(new_n3456_), .ZN(new_n18581_));
  AOI22_X1   g18325(.A1(new_n3864_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n3869_), .ZN(new_n18582_));
  OAI21_X1   g18326(.A1(new_n12147_), .A2(new_n5410_), .B(new_n18582_), .ZN(new_n18583_));
  AOI21_X1   g18327(.A1(new_n13444_), .A2(new_n3872_), .B(new_n18583_), .ZN(new_n18584_));
  XOR2_X1    g18328(.A1(new_n18584_), .A2(new_n3876_), .Z(new_n18585_));
  OAI21_X1   g18329(.A1(new_n18456_), .A2(new_n18556_), .B(new_n18557_), .ZN(new_n18586_));
  INV_X1     g18330(.I(new_n18586_), .ZN(new_n18587_));
  AOI22_X1   g18331(.A1(new_n5155_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n5160_), .ZN(new_n18588_));
  OAI21_X1   g18332(.A1(new_n9942_), .A2(new_n6877_), .B(new_n18588_), .ZN(new_n18589_));
  AOI21_X1   g18333(.A1(new_n10318_), .A2(new_n5166_), .B(new_n18589_), .ZN(new_n18590_));
  XOR2_X1    g18334(.A1(new_n18590_), .A2(new_n5162_), .Z(new_n18591_));
  INV_X1     g18335(.I(new_n18464_), .ZN(new_n18592_));
  NOR2_X1    g18336(.A1(new_n18542_), .A2(new_n18544_), .ZN(new_n18593_));
  NAND2_X1   g18337(.A1(new_n18542_), .A2(new_n18544_), .ZN(new_n18594_));
  AOI21_X1   g18338(.A1(new_n18592_), .A2(new_n18594_), .B(new_n18593_), .ZN(new_n18595_));
  INV_X1     g18339(.I(new_n18595_), .ZN(new_n18596_));
  OAI22_X1   g18340(.A1(new_n5852_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n5857_), .ZN(new_n18597_));
  AOI21_X1   g18341(.A1(\b[51] ), .A2(new_n6115_), .B(new_n18597_), .ZN(new_n18598_));
  OAI21_X1   g18342(.A1(new_n9385_), .A2(new_n5861_), .B(new_n18598_), .ZN(new_n18599_));
  XOR2_X1    g18343(.A1(new_n18599_), .A2(new_n5849_), .Z(new_n18600_));
  AOI22_X1   g18344(.A1(new_n6569_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n6574_), .ZN(new_n18601_));
  OAI21_X1   g18345(.A1(new_n8127_), .A2(new_n8565_), .B(new_n18601_), .ZN(new_n18602_));
  AOI21_X1   g18346(.A1(new_n9684_), .A2(new_n6579_), .B(new_n18602_), .ZN(new_n18603_));
  XOR2_X1    g18347(.A1(new_n18603_), .A2(new_n6567_), .Z(new_n18604_));
  AOI22_X1   g18348(.A1(new_n8241_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n8246_), .ZN(new_n18605_));
  OAI21_X1   g18349(.A1(new_n6490_), .A2(new_n9114_), .B(new_n18605_), .ZN(new_n18606_));
  AOI21_X1   g18350(.A1(new_n7906_), .A2(new_n8252_), .B(new_n18606_), .ZN(new_n18607_));
  XOR2_X1    g18351(.A1(new_n18607_), .A2(new_n8248_), .Z(new_n18608_));
  INV_X1     g18352(.I(new_n18608_), .ZN(new_n18609_));
  INV_X1     g18353(.I(new_n18475_), .ZN(new_n18610_));
  AOI21_X1   g18354(.A1(new_n18610_), .A2(new_n18512_), .B(new_n18510_), .ZN(new_n18611_));
  AOI22_X1   g18355(.A1(new_n10064_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n10062_), .ZN(new_n18612_));
  OAI21_X1   g18356(.A1(new_n4886_), .A2(new_n10399_), .B(new_n18612_), .ZN(new_n18613_));
  AOI21_X1   g18357(.A1(new_n5351_), .A2(new_n10068_), .B(new_n18613_), .ZN(new_n18614_));
  XOR2_X1    g18358(.A1(new_n18614_), .A2(new_n10057_), .Z(new_n18615_));
  NOR2_X1    g18359(.A1(new_n18480_), .A2(new_n18496_), .ZN(new_n18616_));
  NOR2_X1    g18360(.A1(new_n18616_), .A2(new_n18495_), .ZN(new_n18617_));
  INV_X1     g18361(.I(new_n18617_), .ZN(new_n18618_));
  OAI22_X1   g18362(.A1(new_n12306_), .A2(new_n4666_), .B1(new_n12305_), .B2(new_n4639_), .ZN(new_n18619_));
  AOI21_X1   g18363(.A1(\b[33] ), .A2(new_n12304_), .B(new_n18619_), .ZN(new_n18620_));
  OAI21_X1   g18364(.A1(new_n4676_), .A2(new_n10985_), .B(new_n18620_), .ZN(new_n18621_));
  XOR2_X1    g18365(.A1(new_n18621_), .A2(new_n10989_), .Z(new_n18622_));
  AOI22_X1   g18366(.A1(new_n11926_), .A2(\b[32] ), .B1(new_n11924_), .B2(\b[31] ), .ZN(new_n18623_));
  OAI21_X1   g18367(.A1(new_n3624_), .A2(new_n12317_), .B(new_n18623_), .ZN(new_n18624_));
  AOI21_X1   g18368(.A1(new_n4030_), .A2(new_n11929_), .B(new_n18624_), .ZN(new_n18625_));
  XOR2_X1    g18369(.A1(new_n18625_), .A2(new_n12312_), .Z(new_n18626_));
  NOR2_X1    g18370(.A1(new_n18484_), .A2(new_n18488_), .ZN(new_n18627_));
  NOR2_X1    g18371(.A1(new_n18627_), .A2(new_n18489_), .ZN(new_n18628_));
  AOI22_X1   g18372(.A1(new_n12922_), .A2(\b[29] ), .B1(\b[28] ), .B2(new_n12923_), .ZN(new_n18629_));
  INV_X1     g18373(.I(new_n18629_), .ZN(new_n18630_));
  NOR2_X1    g18374(.A1(new_n18630_), .A2(new_n18487_), .ZN(new_n18631_));
  INV_X1     g18375(.I(new_n18487_), .ZN(new_n18632_));
  NOR2_X1    g18376(.A1(new_n18632_), .A2(new_n18629_), .ZN(new_n18633_));
  NOR2_X1    g18377(.A1(new_n18631_), .A2(new_n18633_), .ZN(new_n18634_));
  XOR2_X1    g18378(.A1(new_n18628_), .A2(new_n18634_), .Z(new_n18635_));
  NOR2_X1    g18379(.A1(new_n18635_), .A2(new_n18626_), .ZN(new_n18636_));
  INV_X1     g18380(.I(new_n18636_), .ZN(new_n18637_));
  NAND2_X1   g18381(.A1(new_n18635_), .A2(new_n18626_), .ZN(new_n18638_));
  NAND2_X1   g18382(.A1(new_n18637_), .A2(new_n18638_), .ZN(new_n18639_));
  XNOR2_X1   g18383(.A1(new_n18639_), .A2(new_n18622_), .ZN(new_n18640_));
  NOR2_X1    g18384(.A1(new_n18640_), .A2(new_n18618_), .ZN(new_n18641_));
  NAND2_X1   g18385(.A1(new_n18640_), .A2(new_n18618_), .ZN(new_n18642_));
  INV_X1     g18386(.I(new_n18642_), .ZN(new_n18643_));
  NOR2_X1    g18387(.A1(new_n18643_), .A2(new_n18641_), .ZN(new_n18644_));
  XOR2_X1    g18388(.A1(new_n18644_), .A2(new_n18615_), .Z(new_n18645_));
  INV_X1     g18389(.I(new_n18645_), .ZN(new_n18646_));
  OAI22_X1   g18390(.A1(new_n10390_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n10389_), .ZN(new_n18647_));
  AOI21_X1   g18391(.A1(\b[39] ), .A2(new_n9471_), .B(new_n18647_), .ZN(new_n18648_));
  OAI21_X1   g18392(.A1(new_n6299_), .A2(new_n10388_), .B(new_n18648_), .ZN(new_n18649_));
  XOR2_X1    g18393(.A1(new_n18649_), .A2(\a[53] ), .Z(new_n18650_));
  AOI21_X1   g18394(.A1(new_n18499_), .A2(new_n18507_), .B(new_n18505_), .ZN(new_n18651_));
  OR2_X2     g18395(.A1(new_n18650_), .A2(new_n18651_), .Z(new_n18652_));
  NAND2_X1   g18396(.A1(new_n18650_), .A2(new_n18651_), .ZN(new_n18653_));
  NAND2_X1   g18397(.A1(new_n18652_), .A2(new_n18653_), .ZN(new_n18654_));
  XOR2_X1    g18398(.A1(new_n18654_), .A2(new_n18646_), .Z(new_n18655_));
  NOR2_X1    g18399(.A1(new_n18655_), .A2(new_n18611_), .ZN(new_n18656_));
  INV_X1     g18400(.I(new_n18656_), .ZN(new_n18657_));
  NAND2_X1   g18401(.A1(new_n18655_), .A2(new_n18611_), .ZN(new_n18658_));
  NAND2_X1   g18402(.A1(new_n18657_), .A2(new_n18658_), .ZN(new_n18659_));
  XOR2_X1    g18403(.A1(new_n18659_), .A2(new_n18609_), .Z(new_n18660_));
  AOI22_X1   g18404(.A1(new_n7403_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n7408_), .ZN(new_n18661_));
  OAI21_X1   g18405(.A1(new_n7096_), .A2(new_n9488_), .B(new_n18661_), .ZN(new_n18662_));
  AOI21_X1   g18406(.A1(new_n7649_), .A2(new_n7414_), .B(new_n18662_), .ZN(new_n18663_));
  XOR2_X1    g18407(.A1(new_n18663_), .A2(new_n7410_), .Z(new_n18664_));
  NOR2_X1    g18408(.A1(new_n18522_), .A2(new_n18471_), .ZN(new_n18665_));
  NOR2_X1    g18409(.A1(new_n18665_), .A2(new_n18520_), .ZN(new_n18666_));
  NOR2_X1    g18410(.A1(new_n18666_), .A2(new_n18664_), .ZN(new_n18667_));
  AND2_X2    g18411(.A1(new_n18666_), .A2(new_n18664_), .Z(new_n18668_));
  NOR2_X1    g18412(.A1(new_n18668_), .A2(new_n18667_), .ZN(new_n18669_));
  XOR2_X1    g18413(.A1(new_n18669_), .A2(new_n18660_), .Z(new_n18670_));
  AOI21_X1   g18414(.A1(new_n18469_), .A2(new_n18529_), .B(new_n18527_), .ZN(new_n18671_));
  NOR2_X1    g18415(.A1(new_n18670_), .A2(new_n18671_), .ZN(new_n18672_));
  INV_X1     g18416(.I(new_n18672_), .ZN(new_n18673_));
  NAND2_X1   g18417(.A1(new_n18670_), .A2(new_n18671_), .ZN(new_n18674_));
  NAND2_X1   g18418(.A1(new_n18673_), .A2(new_n18674_), .ZN(new_n18675_));
  XOR2_X1    g18419(.A1(new_n18675_), .A2(new_n18604_), .Z(new_n18676_));
  INV_X1     g18420(.I(new_n18676_), .ZN(new_n18677_));
  NOR2_X1    g18421(.A1(new_n18531_), .A2(new_n18540_), .ZN(new_n18678_));
  NOR2_X1    g18422(.A1(new_n18678_), .A2(new_n18538_), .ZN(new_n18679_));
  NOR2_X1    g18423(.A1(new_n18677_), .A2(new_n18679_), .ZN(new_n18680_));
  INV_X1     g18424(.I(new_n18680_), .ZN(new_n18681_));
  NAND2_X1   g18425(.A1(new_n18677_), .A2(new_n18679_), .ZN(new_n18682_));
  NAND2_X1   g18426(.A1(new_n18681_), .A2(new_n18682_), .ZN(new_n18683_));
  XNOR2_X1   g18427(.A1(new_n18683_), .A2(new_n18600_), .ZN(new_n18684_));
  NOR2_X1    g18428(.A1(new_n18684_), .A2(new_n18596_), .ZN(new_n18685_));
  NAND2_X1   g18429(.A1(new_n18684_), .A2(new_n18596_), .ZN(new_n18686_));
  INV_X1     g18430(.I(new_n18686_), .ZN(new_n18687_));
  NOR2_X1    g18431(.A1(new_n18687_), .A2(new_n18685_), .ZN(new_n18688_));
  XOR2_X1    g18432(.A1(new_n18688_), .A2(new_n18591_), .Z(new_n18689_));
  OAI22_X1   g18433(.A1(new_n12151_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n11195_), .ZN(new_n18690_));
  AOI21_X1   g18434(.A1(\b[57] ), .A2(new_n4706_), .B(new_n18690_), .ZN(new_n18691_));
  OAI21_X1   g18435(.A1(new_n12203_), .A2(new_n4458_), .B(new_n18691_), .ZN(new_n18692_));
  XOR2_X1    g18436(.A1(new_n18692_), .A2(\a[35] ), .Z(new_n18693_));
  AOI21_X1   g18437(.A1(new_n18460_), .A2(new_n18552_), .B(new_n18551_), .ZN(new_n18694_));
  NOR2_X1    g18438(.A1(new_n18694_), .A2(new_n18693_), .ZN(new_n18695_));
  AND2_X2    g18439(.A1(new_n18694_), .A2(new_n18693_), .Z(new_n18696_));
  NOR2_X1    g18440(.A1(new_n18696_), .A2(new_n18695_), .ZN(new_n18697_));
  XOR2_X1    g18441(.A1(new_n18689_), .A2(new_n18697_), .Z(new_n18698_));
  NOR2_X1    g18442(.A1(new_n18698_), .A2(new_n18587_), .ZN(new_n18699_));
  INV_X1     g18443(.I(new_n18699_), .ZN(new_n18700_));
  NAND2_X1   g18444(.A1(new_n18698_), .A2(new_n18587_), .ZN(new_n18701_));
  NAND2_X1   g18445(.A1(new_n18700_), .A2(new_n18701_), .ZN(new_n18702_));
  XOR2_X1    g18446(.A1(new_n18702_), .A2(new_n18585_), .Z(new_n18703_));
  XOR2_X1    g18447(.A1(new_n18703_), .A2(new_n18581_), .Z(new_n18704_));
  NAND2_X1   g18448(.A1(new_n18562_), .A2(new_n18451_), .ZN(new_n18705_));
  NAND2_X1   g18449(.A1(new_n18705_), .A2(new_n18561_), .ZN(new_n18706_));
  XOR2_X1    g18450(.A1(new_n18706_), .A2(\a[29] ), .Z(new_n18707_));
  XOR2_X1    g18451(.A1(new_n18704_), .A2(new_n18707_), .Z(new_n18708_));
  NOR2_X1    g18452(.A1(new_n18708_), .A2(new_n18580_), .ZN(new_n18709_));
  INV_X1     g18453(.I(new_n18709_), .ZN(new_n18710_));
  NAND2_X1   g18454(.A1(new_n18708_), .A2(new_n18580_), .ZN(new_n18711_));
  AND2_X2    g18455(.A1(new_n18710_), .A2(new_n18711_), .Z(new_n18712_));
  INV_X1     g18456(.I(new_n18712_), .ZN(new_n18713_));
  XOR2_X1    g18457(.A1(new_n18579_), .A2(new_n18713_), .Z(\f[92] ));
  OAI21_X1   g18458(.A1(new_n18579_), .A2(new_n18713_), .B(new_n18710_), .ZN(new_n18715_));
  NOR2_X1    g18459(.A1(new_n18703_), .A2(new_n18706_), .ZN(new_n18716_));
  XOR2_X1    g18460(.A1(new_n18581_), .A2(new_n3264_), .Z(new_n18717_));
  NOR2_X1    g18461(.A1(new_n18716_), .A2(new_n18717_), .ZN(new_n18718_));
  AOI21_X1   g18462(.A1(new_n18703_), .A2(new_n18706_), .B(new_n18718_), .ZN(new_n18719_));
  INV_X1     g18463(.I(new_n18719_), .ZN(new_n18720_));
  INV_X1     g18464(.I(new_n18585_), .ZN(new_n18721_));
  AOI21_X1   g18465(.A1(new_n18721_), .A2(new_n18701_), .B(new_n18699_), .ZN(new_n18722_));
  AOI22_X1   g18466(.A1(new_n3864_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n3869_), .ZN(new_n18723_));
  OAI21_X1   g18467(.A1(new_n12148_), .A2(new_n5410_), .B(new_n18723_), .ZN(new_n18724_));
  AOI21_X1   g18468(.A1(new_n12811_), .A2(new_n3872_), .B(new_n18724_), .ZN(new_n18725_));
  XOR2_X1    g18469(.A1(new_n18725_), .A2(new_n3876_), .Z(new_n18726_));
  INV_X1     g18470(.I(new_n18726_), .ZN(new_n18727_));
  OAI21_X1   g18471(.A1(new_n18591_), .A2(new_n18685_), .B(new_n18686_), .ZN(new_n18728_));
  AOI21_X1   g18472(.A1(new_n18600_), .A2(new_n18682_), .B(new_n18680_), .ZN(new_n18729_));
  INV_X1     g18473(.I(new_n18729_), .ZN(new_n18730_));
  AOI22_X1   g18474(.A1(new_n6108_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n6111_), .ZN(new_n18731_));
  OAI21_X1   g18475(.A1(new_n9032_), .A2(new_n7708_), .B(new_n18731_), .ZN(new_n18732_));
  AOI21_X1   g18476(.A1(new_n10884_), .A2(new_n6105_), .B(new_n18732_), .ZN(new_n18733_));
  XOR2_X1    g18477(.A1(new_n18733_), .A2(new_n5849_), .Z(new_n18734_));
  INV_X1     g18478(.I(new_n18604_), .ZN(new_n18735_));
  AOI21_X1   g18479(.A1(new_n18735_), .A2(new_n18674_), .B(new_n18672_), .ZN(new_n18736_));
  INV_X1     g18480(.I(new_n18736_), .ZN(new_n18737_));
  AOI21_X1   g18481(.A1(new_n18609_), .A2(new_n18658_), .B(new_n18656_), .ZN(new_n18738_));
  NAND2_X1   g18482(.A1(new_n18646_), .A2(new_n18653_), .ZN(new_n18739_));
  NAND2_X1   g18483(.A1(new_n18739_), .A2(new_n18652_), .ZN(new_n18740_));
  OAI21_X1   g18484(.A1(new_n18615_), .A2(new_n18641_), .B(new_n18642_), .ZN(new_n18741_));
  AOI21_X1   g18485(.A1(new_n18622_), .A2(new_n18638_), .B(new_n18636_), .ZN(new_n18742_));
  INV_X1     g18486(.I(new_n18742_), .ZN(new_n18743_));
  INV_X1     g18487(.I(new_n18633_), .ZN(new_n18744_));
  OAI21_X1   g18488(.A1(new_n18628_), .A2(new_n18631_), .B(new_n18744_), .ZN(new_n18745_));
  AOI22_X1   g18489(.A1(new_n11926_), .A2(\b[33] ), .B1(new_n11924_), .B2(\b[32] ), .ZN(new_n18746_));
  OAI21_X1   g18490(.A1(new_n4022_), .A2(new_n12317_), .B(new_n18746_), .ZN(new_n18747_));
  AOI21_X1   g18491(.A1(new_n4223_), .A2(new_n11929_), .B(new_n18747_), .ZN(new_n18748_));
  XOR2_X1    g18492(.A1(new_n18748_), .A2(new_n12312_), .Z(new_n18749_));
  AOI22_X1   g18493(.A1(new_n12922_), .A2(\b[30] ), .B1(\b[29] ), .B2(new_n12923_), .ZN(new_n18750_));
  XOR2_X1    g18494(.A1(new_n18750_), .A2(new_n3264_), .Z(new_n18751_));
  XOR2_X1    g18495(.A1(new_n18751_), .A2(new_n18629_), .Z(new_n18752_));
  NOR2_X1    g18496(.A1(new_n18749_), .A2(new_n18752_), .ZN(new_n18753_));
  INV_X1     g18497(.I(new_n18753_), .ZN(new_n18754_));
  NAND2_X1   g18498(.A1(new_n18749_), .A2(new_n18752_), .ZN(new_n18755_));
  NAND2_X1   g18499(.A1(new_n18754_), .A2(new_n18755_), .ZN(new_n18756_));
  XOR2_X1    g18500(.A1(new_n18756_), .A2(new_n18745_), .Z(new_n18757_));
  AOI22_X1   g18501(.A1(new_n10981_), .A2(\b[36] ), .B1(new_n10979_), .B2(\b[35] ), .ZN(new_n18758_));
  OAI21_X1   g18502(.A1(new_n4639_), .A2(new_n11306_), .B(new_n18758_), .ZN(new_n18759_));
  AOI21_X1   g18503(.A1(new_n5594_), .A2(new_n10984_), .B(new_n18759_), .ZN(new_n18760_));
  XOR2_X1    g18504(.A1(new_n18760_), .A2(new_n10989_), .Z(new_n18761_));
  NOR2_X1    g18505(.A1(new_n18757_), .A2(new_n18761_), .ZN(new_n18762_));
  NAND2_X1   g18506(.A1(new_n18757_), .A2(new_n18761_), .ZN(new_n18763_));
  INV_X1     g18507(.I(new_n18763_), .ZN(new_n18764_));
  NOR2_X1    g18508(.A1(new_n18764_), .A2(new_n18762_), .ZN(new_n18765_));
  XOR2_X1    g18509(.A1(new_n18765_), .A2(new_n18743_), .Z(new_n18766_));
  INV_X1     g18510(.I(new_n18766_), .ZN(new_n18767_));
  AOI22_X1   g18511(.A1(new_n10064_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n10062_), .ZN(new_n18768_));
  OAI21_X1   g18512(.A1(new_n5312_), .A2(new_n10399_), .B(new_n18768_), .ZN(new_n18769_));
  AOI21_X1   g18513(.A1(new_n6310_), .A2(new_n10068_), .B(new_n18769_), .ZN(new_n18770_));
  XOR2_X1    g18514(.A1(new_n18770_), .A2(new_n10057_), .Z(new_n18771_));
  NOR2_X1    g18515(.A1(new_n18767_), .A2(new_n18771_), .ZN(new_n18772_));
  INV_X1     g18516(.I(new_n18772_), .ZN(new_n18773_));
  NAND2_X1   g18517(.A1(new_n18767_), .A2(new_n18771_), .ZN(new_n18774_));
  NAND2_X1   g18518(.A1(new_n18773_), .A2(new_n18774_), .ZN(new_n18775_));
  XOR2_X1    g18519(.A1(new_n18775_), .A2(new_n18741_), .Z(new_n18776_));
  AOI22_X1   g18520(.A1(new_n9125_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n9123_), .ZN(new_n18777_));
  OAI21_X1   g18521(.A1(new_n6284_), .A2(new_n9470_), .B(new_n18777_), .ZN(new_n18778_));
  AOI21_X1   g18522(.A1(new_n7106_), .A2(new_n9129_), .B(new_n18778_), .ZN(new_n18779_));
  XOR2_X1    g18523(.A1(new_n18779_), .A2(new_n9133_), .Z(new_n18780_));
  NOR2_X1    g18524(.A1(new_n18776_), .A2(new_n18780_), .ZN(new_n18781_));
  NAND2_X1   g18525(.A1(new_n18776_), .A2(new_n18780_), .ZN(new_n18782_));
  INV_X1     g18526(.I(new_n18782_), .ZN(new_n18783_));
  NOR2_X1    g18527(.A1(new_n18783_), .A2(new_n18781_), .ZN(new_n18784_));
  XOR2_X1    g18528(.A1(new_n18784_), .A2(new_n18740_), .Z(new_n18785_));
  AOI22_X1   g18529(.A1(new_n8241_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n8246_), .ZN(new_n18786_));
  OAI21_X1   g18530(.A1(new_n6775_), .A2(new_n9114_), .B(new_n18786_), .ZN(new_n18787_));
  AOI21_X1   g18531(.A1(new_n7926_), .A2(new_n8252_), .B(new_n18787_), .ZN(new_n18788_));
  XOR2_X1    g18532(.A1(new_n18788_), .A2(\a[50] ), .Z(new_n18789_));
  NAND2_X1   g18533(.A1(new_n18785_), .A2(new_n18789_), .ZN(new_n18790_));
  NOR2_X1    g18534(.A1(new_n18785_), .A2(new_n18789_), .ZN(new_n18791_));
  INV_X1     g18535(.I(new_n18791_), .ZN(new_n18792_));
  NAND2_X1   g18536(.A1(new_n18792_), .A2(new_n18790_), .ZN(new_n18793_));
  XOR2_X1    g18537(.A1(new_n18793_), .A2(new_n18738_), .Z(new_n18794_));
  AOI22_X1   g18538(.A1(new_n7403_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n7408_), .ZN(new_n18795_));
  OAI21_X1   g18539(.A1(new_n7617_), .A2(new_n9488_), .B(new_n18795_), .ZN(new_n18796_));
  AOI21_X1   g18540(.A1(new_n8792_), .A2(new_n7414_), .B(new_n18796_), .ZN(new_n18797_));
  XOR2_X1    g18541(.A1(new_n18797_), .A2(\a[47] ), .Z(new_n18798_));
  INV_X1     g18542(.I(new_n18667_), .ZN(new_n18799_));
  OAI21_X1   g18543(.A1(new_n18660_), .A2(new_n18668_), .B(new_n18799_), .ZN(new_n18800_));
  NAND2_X1   g18544(.A1(new_n18800_), .A2(new_n18798_), .ZN(new_n18801_));
  OR2_X2     g18545(.A1(new_n18800_), .A2(new_n18798_), .Z(new_n18802_));
  NAND2_X1   g18546(.A1(new_n18802_), .A2(new_n18801_), .ZN(new_n18803_));
  XNOR2_X1   g18547(.A1(new_n18794_), .A2(new_n18803_), .ZN(new_n18804_));
  INV_X1     g18548(.I(new_n18804_), .ZN(new_n18805_));
  AOI22_X1   g18549(.A1(new_n6569_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n6574_), .ZN(new_n18806_));
  OAI21_X1   g18550(.A1(new_n8168_), .A2(new_n8565_), .B(new_n18806_), .ZN(new_n18807_));
  AOI21_X1   g18551(.A1(new_n8783_), .A2(new_n6579_), .B(new_n18807_), .ZN(new_n18808_));
  XOR2_X1    g18552(.A1(new_n18808_), .A2(new_n6567_), .Z(new_n18809_));
  NOR2_X1    g18553(.A1(new_n18805_), .A2(new_n18809_), .ZN(new_n18810_));
  INV_X1     g18554(.I(new_n18810_), .ZN(new_n18811_));
  NAND2_X1   g18555(.A1(new_n18805_), .A2(new_n18809_), .ZN(new_n18812_));
  NAND2_X1   g18556(.A1(new_n18811_), .A2(new_n18812_), .ZN(new_n18813_));
  XOR2_X1    g18557(.A1(new_n18813_), .A2(new_n18737_), .Z(new_n18814_));
  NOR2_X1    g18558(.A1(new_n18814_), .A2(new_n18734_), .ZN(new_n18815_));
  NAND2_X1   g18559(.A1(new_n18814_), .A2(new_n18734_), .ZN(new_n18816_));
  INV_X1     g18560(.I(new_n18816_), .ZN(new_n18817_));
  NOR2_X1    g18561(.A1(new_n18817_), .A2(new_n18815_), .ZN(new_n18818_));
  XOR2_X1    g18562(.A1(new_n18818_), .A2(new_n18730_), .Z(new_n18819_));
  INV_X1     g18563(.I(new_n18819_), .ZN(new_n18820_));
  AOI22_X1   g18564(.A1(new_n5155_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n5160_), .ZN(new_n18821_));
  OAI21_X1   g18565(.A1(new_n9972_), .A2(new_n6877_), .B(new_n18821_), .ZN(new_n18822_));
  AOI21_X1   g18566(.A1(new_n10631_), .A2(new_n5166_), .B(new_n18822_), .ZN(new_n18823_));
  XOR2_X1    g18567(.A1(new_n18823_), .A2(new_n5162_), .Z(new_n18824_));
  NOR2_X1    g18568(.A1(new_n18820_), .A2(new_n18824_), .ZN(new_n18825_));
  INV_X1     g18569(.I(new_n18825_), .ZN(new_n18826_));
  NAND2_X1   g18570(.A1(new_n18820_), .A2(new_n18824_), .ZN(new_n18827_));
  NAND2_X1   g18571(.A1(new_n18826_), .A2(new_n18827_), .ZN(new_n18828_));
  XNOR2_X1   g18572(.A1(new_n18828_), .A2(new_n18728_), .ZN(new_n18829_));
  AOI22_X1   g18573(.A1(new_n4918_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n4921_), .ZN(new_n18830_));
  OAI21_X1   g18574(.A1(new_n11195_), .A2(new_n6099_), .B(new_n18830_), .ZN(new_n18831_));
  AOI21_X1   g18575(.A1(new_n11836_), .A2(new_n4699_), .B(new_n18831_), .ZN(new_n18832_));
  XOR2_X1    g18576(.A1(new_n18832_), .A2(\a[35] ), .Z(new_n18833_));
  INV_X1     g18577(.I(new_n18695_), .ZN(new_n18834_));
  OAI21_X1   g18578(.A1(new_n18689_), .A2(new_n18696_), .B(new_n18834_), .ZN(new_n18835_));
  NAND2_X1   g18579(.A1(new_n18835_), .A2(new_n18833_), .ZN(new_n18836_));
  OR2_X2     g18580(.A1(new_n18835_), .A2(new_n18833_), .Z(new_n18837_));
  NAND2_X1   g18581(.A1(new_n18837_), .A2(new_n18836_), .ZN(new_n18838_));
  XNOR2_X1   g18582(.A1(new_n18829_), .A2(new_n18838_), .ZN(new_n18839_));
  NOR2_X1    g18583(.A1(new_n18839_), .A2(new_n18727_), .ZN(new_n18840_));
  NAND2_X1   g18584(.A1(new_n18839_), .A2(new_n18727_), .ZN(new_n18841_));
  INV_X1     g18585(.I(new_n18841_), .ZN(new_n18842_));
  NOR2_X1    g18586(.A1(new_n18842_), .A2(new_n18840_), .ZN(new_n18843_));
  XNOR2_X1   g18587(.A1(new_n18843_), .A2(new_n18722_), .ZN(new_n18844_));
  NOR2_X1    g18588(.A1(new_n18844_), .A2(new_n18720_), .ZN(new_n18845_));
  INV_X1     g18589(.I(new_n18845_), .ZN(new_n18846_));
  NAND2_X1   g18590(.A1(new_n18844_), .A2(new_n18720_), .ZN(new_n18847_));
  AND2_X2    g18591(.A1(new_n18846_), .A2(new_n18847_), .Z(new_n18848_));
  XOR2_X1    g18592(.A1(new_n18715_), .A2(new_n18848_), .Z(\f[93] ));
  OAI22_X1   g18593(.A1(new_n5410_), .A2(new_n12796_), .B1(new_n12800_), .B2(new_n4730_), .ZN(new_n18850_));
  AOI21_X1   g18594(.A1(new_n13973_), .A2(new_n3872_), .B(new_n18850_), .ZN(new_n18851_));
  XOR2_X1    g18595(.A1(new_n18851_), .A2(new_n3876_), .Z(new_n18852_));
  INV_X1     g18596(.I(new_n18852_), .ZN(new_n18853_));
  INV_X1     g18597(.I(new_n18836_), .ZN(new_n18854_));
  AOI21_X1   g18598(.A1(new_n18829_), .A2(new_n18837_), .B(new_n18854_), .ZN(new_n18855_));
  INV_X1     g18599(.I(new_n18855_), .ZN(new_n18856_));
  AOI21_X1   g18600(.A1(new_n18728_), .A2(new_n18827_), .B(new_n18825_), .ZN(new_n18857_));
  OAI22_X1   g18601(.A1(new_n12148_), .A2(new_n4449_), .B1(new_n4454_), .B2(new_n12147_), .ZN(new_n18858_));
  AOI21_X1   g18602(.A1(\b[59] ), .A2(new_n4706_), .B(new_n18858_), .ZN(new_n18859_));
  OAI21_X1   g18603(.A1(new_n13110_), .A2(new_n4458_), .B(new_n18859_), .ZN(new_n18860_));
  XOR2_X1    g18604(.A1(new_n18860_), .A2(\a[35] ), .Z(new_n18861_));
  NOR2_X1    g18605(.A1(new_n18857_), .A2(new_n18861_), .ZN(new_n18862_));
  INV_X1     g18606(.I(new_n18862_), .ZN(new_n18863_));
  NAND2_X1   g18607(.A1(new_n18857_), .A2(new_n18861_), .ZN(new_n18864_));
  NAND2_X1   g18608(.A1(new_n18863_), .A2(new_n18864_), .ZN(new_n18865_));
  AOI22_X1   g18609(.A1(new_n5155_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n5160_), .ZN(new_n18866_));
  OAI21_X1   g18610(.A1(new_n10308_), .A2(new_n6877_), .B(new_n18866_), .ZN(new_n18867_));
  AOI21_X1   g18611(.A1(new_n12164_), .A2(new_n5166_), .B(new_n18867_), .ZN(new_n18868_));
  XOR2_X1    g18612(.A1(new_n18868_), .A2(new_n5162_), .Z(new_n18869_));
  INV_X1     g18613(.I(new_n18869_), .ZN(new_n18870_));
  AOI21_X1   g18614(.A1(new_n18730_), .A2(new_n18816_), .B(new_n18815_), .ZN(new_n18871_));
  INV_X1     g18615(.I(new_n18871_), .ZN(new_n18872_));
  AOI21_X1   g18616(.A1(new_n18737_), .A2(new_n18812_), .B(new_n18810_), .ZN(new_n18873_));
  INV_X1     g18617(.I(new_n18873_), .ZN(new_n18874_));
  AOI22_X1   g18618(.A1(new_n6569_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n6574_), .ZN(new_n18875_));
  OAI21_X1   g18619(.A1(new_n8500_), .A2(new_n8565_), .B(new_n18875_), .ZN(new_n18876_));
  AOI21_X1   g18620(.A1(new_n9987_), .A2(new_n6579_), .B(new_n18876_), .ZN(new_n18877_));
  XOR2_X1    g18621(.A1(new_n18877_), .A2(new_n6567_), .Z(new_n18878_));
  AOI22_X1   g18622(.A1(new_n8241_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n8246_), .ZN(new_n18879_));
  OAI21_X1   g18623(.A1(new_n7074_), .A2(new_n9114_), .B(new_n18879_), .ZN(new_n18880_));
  AOI21_X1   g18624(.A1(new_n9337_), .A2(new_n8252_), .B(new_n18880_), .ZN(new_n18881_));
  XOR2_X1    g18625(.A1(new_n18881_), .A2(new_n8248_), .Z(new_n18882_));
  INV_X1     g18626(.I(new_n18882_), .ZN(new_n18883_));
  AOI21_X1   g18627(.A1(new_n18741_), .A2(new_n18774_), .B(new_n18772_), .ZN(new_n18884_));
  AOI22_X1   g18628(.A1(new_n10064_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n10062_), .ZN(new_n18885_));
  OAI21_X1   g18629(.A1(new_n5341_), .A2(new_n10399_), .B(new_n18885_), .ZN(new_n18886_));
  AOI21_X1   g18630(.A1(new_n5793_), .A2(new_n10068_), .B(new_n18886_), .ZN(new_n18887_));
  XOR2_X1    g18631(.A1(new_n18887_), .A2(new_n10057_), .Z(new_n18888_));
  AOI21_X1   g18632(.A1(new_n18743_), .A2(new_n18763_), .B(new_n18762_), .ZN(new_n18889_));
  INV_X1     g18633(.I(new_n18889_), .ZN(new_n18890_));
  OAI22_X1   g18634(.A1(new_n12306_), .A2(new_n5312_), .B1(new_n12305_), .B2(new_n4886_), .ZN(new_n18891_));
  AOI21_X1   g18635(.A1(\b[35] ), .A2(new_n12304_), .B(new_n18891_), .ZN(new_n18892_));
  OAI21_X1   g18636(.A1(new_n5322_), .A2(new_n10985_), .B(new_n18892_), .ZN(new_n18893_));
  XOR2_X1    g18637(.A1(new_n18893_), .A2(new_n10989_), .Z(new_n18894_));
  AOI21_X1   g18638(.A1(new_n18745_), .A2(new_n18755_), .B(new_n18753_), .ZN(new_n18895_));
  AOI22_X1   g18639(.A1(new_n11926_), .A2(\b[34] ), .B1(new_n11924_), .B2(\b[33] ), .ZN(new_n18896_));
  OAI21_X1   g18640(.A1(new_n4023_), .A2(new_n12317_), .B(new_n18896_), .ZN(new_n18897_));
  AOI21_X1   g18641(.A1(new_n5103_), .A2(new_n11929_), .B(new_n18897_), .ZN(new_n18898_));
  XOR2_X1    g18642(.A1(new_n18898_), .A2(new_n12312_), .Z(new_n18899_));
  NOR2_X1    g18643(.A1(new_n18750_), .A2(\a[29] ), .ZN(new_n18900_));
  NOR2_X1    g18644(.A1(new_n18900_), .A2(new_n18630_), .ZN(new_n18901_));
  AOI21_X1   g18645(.A1(\a[29] ), .A2(new_n18750_), .B(new_n18901_), .ZN(new_n18902_));
  AOI22_X1   g18646(.A1(new_n12922_), .A2(\b[31] ), .B1(\b[30] ), .B2(new_n12923_), .ZN(new_n18903_));
  AND2_X2    g18647(.A1(new_n18902_), .A2(new_n18903_), .Z(new_n18904_));
  NOR2_X1    g18648(.A1(new_n18902_), .A2(new_n18903_), .ZN(new_n18905_));
  NOR2_X1    g18649(.A1(new_n18904_), .A2(new_n18905_), .ZN(new_n18906_));
  XNOR2_X1   g18650(.A1(new_n18899_), .A2(new_n18906_), .ZN(new_n18907_));
  INV_X1     g18651(.I(new_n18907_), .ZN(new_n18908_));
  NAND2_X1   g18652(.A1(new_n18908_), .A2(new_n18895_), .ZN(new_n18909_));
  NOR2_X1    g18653(.A1(new_n18908_), .A2(new_n18895_), .ZN(new_n18910_));
  INV_X1     g18654(.I(new_n18910_), .ZN(new_n18911_));
  NAND2_X1   g18655(.A1(new_n18911_), .A2(new_n18909_), .ZN(new_n18912_));
  XNOR2_X1   g18656(.A1(new_n18912_), .A2(new_n18894_), .ZN(new_n18913_));
  NOR2_X1    g18657(.A1(new_n18913_), .A2(new_n18890_), .ZN(new_n18914_));
  INV_X1     g18658(.I(new_n18914_), .ZN(new_n18915_));
  NAND2_X1   g18659(.A1(new_n18913_), .A2(new_n18890_), .ZN(new_n18916_));
  NAND2_X1   g18660(.A1(new_n18915_), .A2(new_n18916_), .ZN(new_n18917_));
  XOR2_X1    g18661(.A1(new_n18917_), .A2(new_n18888_), .Z(new_n18918_));
  INV_X1     g18662(.I(new_n18918_), .ZN(new_n18919_));
  OAI22_X1   g18663(.A1(new_n10390_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n10389_), .ZN(new_n18920_));
  AOI21_X1   g18664(.A1(\b[41] ), .A2(new_n9471_), .B(new_n18920_), .ZN(new_n18921_));
  OAI21_X1   g18665(.A1(new_n6785_), .A2(new_n10388_), .B(new_n18921_), .ZN(new_n18922_));
  XOR2_X1    g18666(.A1(new_n18922_), .A2(\a[53] ), .Z(new_n18923_));
  NOR2_X1    g18667(.A1(new_n18919_), .A2(new_n18923_), .ZN(new_n18924_));
  NAND2_X1   g18668(.A1(new_n18919_), .A2(new_n18923_), .ZN(new_n18925_));
  INV_X1     g18669(.I(new_n18925_), .ZN(new_n18926_));
  NOR2_X1    g18670(.A1(new_n18926_), .A2(new_n18924_), .ZN(new_n18927_));
  XOR2_X1    g18671(.A1(new_n18927_), .A2(new_n18884_), .Z(new_n18928_));
  AOI21_X1   g18672(.A1(new_n18740_), .A2(new_n18782_), .B(new_n18781_), .ZN(new_n18929_));
  NOR2_X1    g18673(.A1(new_n18928_), .A2(new_n18929_), .ZN(new_n18930_));
  INV_X1     g18674(.I(new_n18930_), .ZN(new_n18931_));
  NAND2_X1   g18675(.A1(new_n18928_), .A2(new_n18929_), .ZN(new_n18932_));
  NAND2_X1   g18676(.A1(new_n18931_), .A2(new_n18932_), .ZN(new_n18933_));
  XOR2_X1    g18677(.A1(new_n18933_), .A2(new_n18883_), .Z(new_n18934_));
  OAI21_X1   g18678(.A1(new_n18738_), .A2(new_n18791_), .B(new_n18790_), .ZN(new_n18935_));
  INV_X1     g18679(.I(new_n18935_), .ZN(new_n18936_));
  OAI22_X1   g18680(.A1(new_n8127_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n8168_), .ZN(new_n18937_));
  AOI21_X1   g18681(.A1(\b[47] ), .A2(new_n7719_), .B(new_n18937_), .ZN(new_n18938_));
  OAI21_X1   g18682(.A1(new_n9050_), .A2(new_n8585_), .B(new_n18938_), .ZN(new_n18939_));
  XOR2_X1    g18683(.A1(new_n18939_), .A2(\a[47] ), .Z(new_n18940_));
  NOR2_X1    g18684(.A1(new_n18936_), .A2(new_n18940_), .ZN(new_n18941_));
  NAND2_X1   g18685(.A1(new_n18936_), .A2(new_n18940_), .ZN(new_n18942_));
  INV_X1     g18686(.I(new_n18942_), .ZN(new_n18943_));
  NOR2_X1    g18687(.A1(new_n18943_), .A2(new_n18941_), .ZN(new_n18944_));
  XOR2_X1    g18688(.A1(new_n18944_), .A2(new_n18934_), .Z(new_n18945_));
  INV_X1     g18689(.I(new_n18801_), .ZN(new_n18946_));
  AOI21_X1   g18690(.A1(new_n18794_), .A2(new_n18802_), .B(new_n18946_), .ZN(new_n18947_));
  XOR2_X1    g18691(.A1(new_n18945_), .A2(new_n18947_), .Z(new_n18948_));
  XOR2_X1    g18692(.A1(new_n18948_), .A2(new_n18878_), .Z(new_n18949_));
  AOI22_X1   g18693(.A1(new_n6108_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n6111_), .ZN(new_n18950_));
  OAI21_X1   g18694(.A1(new_n9376_), .A2(new_n7708_), .B(new_n18950_), .ZN(new_n18951_));
  AOI21_X1   g18695(.A1(new_n9979_), .A2(new_n6105_), .B(new_n18951_), .ZN(new_n18952_));
  XOR2_X1    g18696(.A1(new_n18952_), .A2(new_n5849_), .Z(new_n18953_));
  NOR2_X1    g18697(.A1(new_n18949_), .A2(new_n18953_), .ZN(new_n18954_));
  NAND2_X1   g18698(.A1(new_n18949_), .A2(new_n18953_), .ZN(new_n18955_));
  INV_X1     g18699(.I(new_n18955_), .ZN(new_n18956_));
  NOR2_X1    g18700(.A1(new_n18956_), .A2(new_n18954_), .ZN(new_n18957_));
  XOR2_X1    g18701(.A1(new_n18957_), .A2(new_n18874_), .Z(new_n18958_));
  NOR2_X1    g18702(.A1(new_n18958_), .A2(new_n18872_), .ZN(new_n18959_));
  INV_X1     g18703(.I(new_n18959_), .ZN(new_n18960_));
  NAND2_X1   g18704(.A1(new_n18958_), .A2(new_n18872_), .ZN(new_n18961_));
  NAND2_X1   g18705(.A1(new_n18960_), .A2(new_n18961_), .ZN(new_n18962_));
  XOR2_X1    g18706(.A1(new_n18962_), .A2(new_n18870_), .Z(new_n18963_));
  XOR2_X1    g18707(.A1(new_n18865_), .A2(new_n18963_), .Z(new_n18964_));
  NOR2_X1    g18708(.A1(new_n18964_), .A2(new_n18856_), .ZN(new_n18965_));
  INV_X1     g18709(.I(new_n18965_), .ZN(new_n18966_));
  NAND2_X1   g18710(.A1(new_n18964_), .A2(new_n18856_), .ZN(new_n18967_));
  NAND2_X1   g18711(.A1(new_n18966_), .A2(new_n18967_), .ZN(new_n18968_));
  XOR2_X1    g18712(.A1(new_n18968_), .A2(new_n18853_), .Z(new_n18969_));
  OAI21_X1   g18713(.A1(new_n18722_), .A2(new_n18840_), .B(new_n18841_), .ZN(new_n18970_));
  AOI21_X1   g18714(.A1(new_n18715_), .A2(new_n18848_), .B(new_n18845_), .ZN(new_n18971_));
  NOR2_X1    g18715(.A1(new_n18971_), .A2(new_n18970_), .ZN(new_n18972_));
  INV_X1     g18716(.I(new_n18970_), .ZN(new_n18973_));
  NOR3_X1    g18717(.A1(new_n18437_), .A2(new_n18432_), .A3(new_n18571_), .ZN(new_n18974_));
  AOI21_X1   g18718(.A1(new_n18570_), .A2(new_n18572_), .B(new_n18974_), .ZN(new_n18975_));
  AOI21_X1   g18719(.A1(new_n18975_), .A2(new_n18712_), .B(new_n18709_), .ZN(new_n18976_));
  INV_X1     g18720(.I(new_n18848_), .ZN(new_n18977_));
  OAI21_X1   g18721(.A1(new_n18976_), .A2(new_n18977_), .B(new_n18846_), .ZN(new_n18978_));
  NOR2_X1    g18722(.A1(new_n18978_), .A2(new_n18973_), .ZN(new_n18979_));
  NOR2_X1    g18723(.A1(new_n18979_), .A2(new_n18972_), .ZN(new_n18980_));
  XOR2_X1    g18724(.A1(new_n18980_), .A2(new_n18969_), .Z(\f[94] ));
  NAND2_X1   g18725(.A1(new_n18971_), .A2(new_n18970_), .ZN(new_n18982_));
  INV_X1     g18726(.I(new_n18969_), .ZN(new_n18983_));
  OAI21_X1   g18727(.A1(new_n18971_), .A2(new_n18970_), .B(new_n18983_), .ZN(new_n18984_));
  NAND2_X1   g18728(.A1(new_n18984_), .A2(new_n18982_), .ZN(new_n18985_));
  OAI21_X1   g18729(.A1(new_n18852_), .A2(new_n18965_), .B(new_n18967_), .ZN(new_n18986_));
  AOI22_X1   g18730(.A1(new_n13460_), .A2(new_n3872_), .B1(\b[63] ), .B2(new_n4053_), .ZN(new_n18987_));
  AOI22_X1   g18731(.A1(new_n4918_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n4921_), .ZN(new_n18988_));
  OAI21_X1   g18732(.A1(new_n12147_), .A2(new_n6099_), .B(new_n18988_), .ZN(new_n18989_));
  AOI21_X1   g18733(.A1(new_n13444_), .A2(new_n4699_), .B(new_n18989_), .ZN(new_n18990_));
  XOR2_X1    g18734(.A1(new_n18990_), .A2(new_n4446_), .Z(new_n18991_));
  INV_X1     g18735(.I(new_n18991_), .ZN(new_n18992_));
  AOI22_X1   g18736(.A1(new_n6108_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n6111_), .ZN(new_n18993_));
  OAI21_X1   g18737(.A1(new_n9942_), .A2(new_n7708_), .B(new_n18993_), .ZN(new_n18994_));
  AOI21_X1   g18738(.A1(new_n10318_), .A2(new_n6105_), .B(new_n18994_), .ZN(new_n18995_));
  XOR2_X1    g18739(.A1(new_n18995_), .A2(new_n5849_), .Z(new_n18996_));
  INV_X1     g18740(.I(new_n18878_), .ZN(new_n18997_));
  NOR2_X1    g18741(.A1(new_n18945_), .A2(new_n18947_), .ZN(new_n18998_));
  NAND2_X1   g18742(.A1(new_n18945_), .A2(new_n18947_), .ZN(new_n18999_));
  AOI21_X1   g18743(.A1(new_n18997_), .A2(new_n18999_), .B(new_n18998_), .ZN(new_n19000_));
  INV_X1     g18744(.I(new_n19000_), .ZN(new_n19001_));
  OAI22_X1   g18745(.A1(new_n7730_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n7731_), .ZN(new_n19002_));
  AOI21_X1   g18746(.A1(\b[51] ), .A2(new_n6887_), .B(new_n19002_), .ZN(new_n19003_));
  OAI21_X1   g18747(.A1(new_n9385_), .A2(new_n7728_), .B(new_n19003_), .ZN(new_n19004_));
  XOR2_X1    g18748(.A1(new_n19004_), .A2(new_n6567_), .Z(new_n19005_));
  AOI22_X1   g18749(.A1(new_n7403_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n7408_), .ZN(new_n19006_));
  OAI21_X1   g18750(.A1(new_n8127_), .A2(new_n9488_), .B(new_n19006_), .ZN(new_n19007_));
  AOI21_X1   g18751(.A1(new_n9684_), .A2(new_n7414_), .B(new_n19007_), .ZN(new_n19008_));
  XOR2_X1    g18752(.A1(new_n19008_), .A2(new_n7410_), .Z(new_n19009_));
  AOI22_X1   g18753(.A1(new_n9125_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n9123_), .ZN(new_n19010_));
  OAI21_X1   g18754(.A1(new_n6490_), .A2(new_n9470_), .B(new_n19010_), .ZN(new_n19011_));
  AOI21_X1   g18755(.A1(new_n7906_), .A2(new_n9129_), .B(new_n19011_), .ZN(new_n19012_));
  XOR2_X1    g18756(.A1(new_n19012_), .A2(new_n9133_), .Z(new_n19013_));
  OAI21_X1   g18757(.A1(new_n18888_), .A2(new_n18914_), .B(new_n18916_), .ZN(new_n19014_));
  OAI22_X1   g18758(.A1(new_n11298_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n11297_), .ZN(new_n19015_));
  AOI21_X1   g18759(.A1(\b[39] ), .A2(new_n11296_), .B(new_n19015_), .ZN(new_n19016_));
  OAI21_X1   g18760(.A1(new_n6299_), .A2(new_n10069_), .B(new_n19016_), .ZN(new_n19017_));
  XOR2_X1    g18761(.A1(new_n19017_), .A2(\a[56] ), .Z(new_n19018_));
  INV_X1     g18762(.I(new_n18905_), .ZN(new_n19019_));
  OAI21_X1   g18763(.A1(new_n18899_), .A2(new_n18904_), .B(new_n19019_), .ZN(new_n19020_));
  INV_X1     g18764(.I(new_n18903_), .ZN(new_n19021_));
  AOI22_X1   g18765(.A1(new_n12922_), .A2(\b[32] ), .B1(\b[31] ), .B2(new_n12923_), .ZN(new_n19022_));
  NAND2_X1   g18766(.A1(new_n19021_), .A2(new_n19022_), .ZN(new_n19023_));
  NOR2_X1    g18767(.A1(new_n19021_), .A2(new_n19022_), .ZN(new_n19024_));
  INV_X1     g18768(.I(new_n19024_), .ZN(new_n19025_));
  NAND2_X1   g18769(.A1(new_n19025_), .A2(new_n19023_), .ZN(new_n19026_));
  XOR2_X1    g18770(.A1(new_n19020_), .A2(new_n19026_), .Z(new_n19027_));
  INV_X1     g18771(.I(new_n19027_), .ZN(new_n19028_));
  AOI22_X1   g18772(.A1(new_n10981_), .A2(\b[38] ), .B1(new_n10979_), .B2(\b[37] ), .ZN(new_n19029_));
  OAI21_X1   g18773(.A1(new_n4886_), .A2(new_n11306_), .B(new_n19029_), .ZN(new_n19030_));
  AOI21_X1   g18774(.A1(new_n5351_), .A2(new_n10984_), .B(new_n19030_), .ZN(new_n19031_));
  XOR2_X1    g18775(.A1(new_n19031_), .A2(new_n10989_), .Z(new_n19032_));
  OAI22_X1   g18776(.A1(new_n13224_), .A2(new_n4666_), .B1(new_n4639_), .B2(new_n11923_), .ZN(new_n19033_));
  AOI21_X1   g18777(.A1(\b[33] ), .A2(new_n13223_), .B(new_n19033_), .ZN(new_n19034_));
  OAI21_X1   g18778(.A1(new_n4676_), .A2(new_n11930_), .B(new_n19034_), .ZN(new_n19035_));
  XOR2_X1    g18779(.A1(new_n19035_), .A2(\a[62] ), .Z(new_n19036_));
  NOR2_X1    g18780(.A1(new_n19032_), .A2(new_n19036_), .ZN(new_n19037_));
  INV_X1     g18781(.I(new_n19037_), .ZN(new_n19038_));
  NAND2_X1   g18782(.A1(new_n19032_), .A2(new_n19036_), .ZN(new_n19039_));
  NAND2_X1   g18783(.A1(new_n19038_), .A2(new_n19039_), .ZN(new_n19040_));
  XOR2_X1    g18784(.A1(new_n19040_), .A2(new_n19028_), .Z(new_n19041_));
  AOI21_X1   g18785(.A1(new_n18894_), .A2(new_n18909_), .B(new_n18910_), .ZN(new_n19042_));
  XNOR2_X1   g18786(.A1(new_n19041_), .A2(new_n19042_), .ZN(new_n19043_));
  XOR2_X1    g18787(.A1(new_n19043_), .A2(new_n19018_), .Z(new_n19044_));
  NOR2_X1    g18788(.A1(new_n19044_), .A2(new_n19014_), .ZN(new_n19045_));
  INV_X1     g18789(.I(new_n19045_), .ZN(new_n19046_));
  NAND2_X1   g18790(.A1(new_n19044_), .A2(new_n19014_), .ZN(new_n19047_));
  NAND2_X1   g18791(.A1(new_n19046_), .A2(new_n19047_), .ZN(new_n19048_));
  XNOR2_X1   g18792(.A1(new_n19048_), .A2(new_n19013_), .ZN(new_n19049_));
  AOI22_X1   g18793(.A1(new_n8241_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n8246_), .ZN(new_n19050_));
  OAI21_X1   g18794(.A1(new_n7096_), .A2(new_n9114_), .B(new_n19050_), .ZN(new_n19051_));
  AOI21_X1   g18795(.A1(new_n7649_), .A2(new_n8252_), .B(new_n19051_), .ZN(new_n19052_));
  XOR2_X1    g18796(.A1(new_n19052_), .A2(new_n8248_), .Z(new_n19053_));
  NOR2_X1    g18797(.A1(new_n18926_), .A2(new_n18884_), .ZN(new_n19054_));
  NOR2_X1    g18798(.A1(new_n19054_), .A2(new_n18924_), .ZN(new_n19055_));
  NOR2_X1    g18799(.A1(new_n19055_), .A2(new_n19053_), .ZN(new_n19056_));
  AND2_X2    g18800(.A1(new_n19055_), .A2(new_n19053_), .Z(new_n19057_));
  NOR2_X1    g18801(.A1(new_n19057_), .A2(new_n19056_), .ZN(new_n19058_));
  XOR2_X1    g18802(.A1(new_n19058_), .A2(new_n19049_), .Z(new_n19059_));
  AOI21_X1   g18803(.A1(new_n18883_), .A2(new_n18932_), .B(new_n18930_), .ZN(new_n19060_));
  NOR2_X1    g18804(.A1(new_n19059_), .A2(new_n19060_), .ZN(new_n19061_));
  INV_X1     g18805(.I(new_n19061_), .ZN(new_n19062_));
  NAND2_X1   g18806(.A1(new_n19059_), .A2(new_n19060_), .ZN(new_n19063_));
  NAND2_X1   g18807(.A1(new_n19062_), .A2(new_n19063_), .ZN(new_n19064_));
  XOR2_X1    g18808(.A1(new_n19064_), .A2(new_n19009_), .Z(new_n19065_));
  INV_X1     g18809(.I(new_n19065_), .ZN(new_n19066_));
  INV_X1     g18810(.I(new_n18934_), .ZN(new_n19067_));
  AOI21_X1   g18811(.A1(new_n19067_), .A2(new_n18942_), .B(new_n18941_), .ZN(new_n19068_));
  NOR2_X1    g18812(.A1(new_n19066_), .A2(new_n19068_), .ZN(new_n19069_));
  INV_X1     g18813(.I(new_n19069_), .ZN(new_n19070_));
  NAND2_X1   g18814(.A1(new_n19066_), .A2(new_n19068_), .ZN(new_n19071_));
  NAND2_X1   g18815(.A1(new_n19070_), .A2(new_n19071_), .ZN(new_n19072_));
  XNOR2_X1   g18816(.A1(new_n19072_), .A2(new_n19005_), .ZN(new_n19073_));
  NOR2_X1    g18817(.A1(new_n19073_), .A2(new_n19001_), .ZN(new_n19074_));
  NAND2_X1   g18818(.A1(new_n19073_), .A2(new_n19001_), .ZN(new_n19075_));
  INV_X1     g18819(.I(new_n19075_), .ZN(new_n19076_));
  NOR2_X1    g18820(.A1(new_n19076_), .A2(new_n19074_), .ZN(new_n19077_));
  XOR2_X1    g18821(.A1(new_n19077_), .A2(new_n18996_), .Z(new_n19078_));
  OAI22_X1   g18822(.A1(new_n12151_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n11195_), .ZN(new_n19079_));
  AOI21_X1   g18823(.A1(\b[57] ), .A2(new_n5420_), .B(new_n19079_), .ZN(new_n19080_));
  OAI21_X1   g18824(.A1(new_n12203_), .A2(new_n6124_), .B(new_n19080_), .ZN(new_n19081_));
  XOR2_X1    g18825(.A1(new_n19081_), .A2(\a[38] ), .Z(new_n19082_));
  AOI21_X1   g18826(.A1(new_n18874_), .A2(new_n18955_), .B(new_n18954_), .ZN(new_n19083_));
  NOR2_X1    g18827(.A1(new_n19083_), .A2(new_n19082_), .ZN(new_n19084_));
  AND2_X2    g18828(.A1(new_n19083_), .A2(new_n19082_), .Z(new_n19085_));
  NOR2_X1    g18829(.A1(new_n19085_), .A2(new_n19084_), .ZN(new_n19086_));
  XOR2_X1    g18830(.A1(new_n19078_), .A2(new_n19086_), .Z(new_n19087_));
  OAI21_X1   g18831(.A1(new_n18869_), .A2(new_n18959_), .B(new_n18961_), .ZN(new_n19088_));
  INV_X1     g18832(.I(new_n19088_), .ZN(new_n19089_));
  NOR2_X1    g18833(.A1(new_n19087_), .A2(new_n19089_), .ZN(new_n19090_));
  INV_X1     g18834(.I(new_n19090_), .ZN(new_n19091_));
  NAND2_X1   g18835(.A1(new_n19087_), .A2(new_n19089_), .ZN(new_n19092_));
  NAND2_X1   g18836(.A1(new_n19091_), .A2(new_n19092_), .ZN(new_n19093_));
  XOR2_X1    g18837(.A1(new_n19093_), .A2(new_n18992_), .Z(new_n19094_));
  XOR2_X1    g18838(.A1(new_n19094_), .A2(new_n18987_), .Z(new_n19095_));
  INV_X1     g18839(.I(new_n18963_), .ZN(new_n19096_));
  NAND2_X1   g18840(.A1(new_n19096_), .A2(new_n18864_), .ZN(new_n19097_));
  NAND2_X1   g18841(.A1(new_n19097_), .A2(new_n18863_), .ZN(new_n19098_));
  XOR2_X1    g18842(.A1(new_n19098_), .A2(\a[32] ), .Z(new_n19099_));
  XOR2_X1    g18843(.A1(new_n19095_), .A2(new_n19099_), .Z(new_n19100_));
  INV_X1     g18844(.I(new_n19100_), .ZN(new_n19101_));
  NAND2_X1   g18845(.A1(new_n19101_), .A2(new_n18986_), .ZN(new_n19102_));
  NOR2_X1    g18846(.A1(new_n19101_), .A2(new_n18986_), .ZN(new_n19103_));
  INV_X1     g18847(.I(new_n19103_), .ZN(new_n19104_));
  AND2_X2    g18848(.A1(new_n19104_), .A2(new_n19102_), .Z(new_n19105_));
  INV_X1     g18849(.I(new_n19105_), .ZN(new_n19106_));
  XOR2_X1    g18850(.A1(new_n18985_), .A2(new_n19106_), .Z(\f[95] ));
  NAND3_X1   g18851(.A1(new_n18984_), .A2(new_n18982_), .A3(new_n19105_), .ZN(new_n19108_));
  INV_X1     g18852(.I(new_n19094_), .ZN(new_n19109_));
  INV_X1     g18853(.I(new_n19098_), .ZN(new_n19110_));
  XOR2_X1    g18854(.A1(new_n18987_), .A2(new_n3876_), .Z(new_n19111_));
  AOI21_X1   g18855(.A1(new_n19110_), .A2(new_n19094_), .B(new_n19111_), .ZN(new_n19112_));
  AOI21_X1   g18856(.A1(new_n19109_), .A2(new_n19098_), .B(new_n19112_), .ZN(new_n19113_));
  INV_X1     g18857(.I(new_n19113_), .ZN(new_n19114_));
  AOI21_X1   g18858(.A1(new_n18992_), .A2(new_n19092_), .B(new_n19090_), .ZN(new_n19115_));
  AOI22_X1   g18859(.A1(new_n4918_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n4921_), .ZN(new_n19116_));
  OAI21_X1   g18860(.A1(new_n12148_), .A2(new_n6099_), .B(new_n19116_), .ZN(new_n19117_));
  AOI21_X1   g18861(.A1(new_n12811_), .A2(new_n4699_), .B(new_n19117_), .ZN(new_n19118_));
  XOR2_X1    g18862(.A1(new_n19118_), .A2(new_n4446_), .Z(new_n19119_));
  INV_X1     g18863(.I(new_n19119_), .ZN(new_n19120_));
  OAI21_X1   g18864(.A1(new_n18996_), .A2(new_n19074_), .B(new_n19075_), .ZN(new_n19121_));
  AOI21_X1   g18865(.A1(new_n19005_), .A2(new_n19071_), .B(new_n19069_), .ZN(new_n19122_));
  INV_X1     g18866(.I(new_n19122_), .ZN(new_n19123_));
  AOI22_X1   g18867(.A1(new_n6569_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n6574_), .ZN(new_n19124_));
  OAI21_X1   g18868(.A1(new_n9032_), .A2(new_n8565_), .B(new_n19124_), .ZN(new_n19125_));
  AOI21_X1   g18869(.A1(new_n10884_), .A2(new_n6579_), .B(new_n19125_), .ZN(new_n19126_));
  XOR2_X1    g18870(.A1(new_n19126_), .A2(new_n6567_), .Z(new_n19127_));
  INV_X1     g18871(.I(new_n19009_), .ZN(new_n19128_));
  AOI21_X1   g18872(.A1(new_n19128_), .A2(new_n19063_), .B(new_n19061_), .ZN(new_n19129_));
  INV_X1     g18873(.I(new_n19129_), .ZN(new_n19130_));
  OAI21_X1   g18874(.A1(new_n19013_), .A2(new_n19045_), .B(new_n19047_), .ZN(new_n19131_));
  AOI21_X1   g18875(.A1(new_n19028_), .A2(new_n19039_), .B(new_n19037_), .ZN(new_n19132_));
  AOI21_X1   g18876(.A1(new_n19020_), .A2(new_n19023_), .B(new_n19024_), .ZN(new_n19133_));
  AOI22_X1   g18877(.A1(new_n11926_), .A2(\b[36] ), .B1(new_n11924_), .B2(\b[35] ), .ZN(new_n19134_));
  OAI21_X1   g18878(.A1(new_n4639_), .A2(new_n12317_), .B(new_n19134_), .ZN(new_n19135_));
  AOI21_X1   g18879(.A1(new_n5594_), .A2(new_n11929_), .B(new_n19135_), .ZN(new_n19136_));
  XOR2_X1    g18880(.A1(new_n19136_), .A2(new_n12312_), .Z(new_n19137_));
  AOI22_X1   g18881(.A1(new_n12922_), .A2(\b[33] ), .B1(\b[32] ), .B2(new_n12923_), .ZN(new_n19138_));
  XOR2_X1    g18882(.A1(new_n19138_), .A2(new_n3876_), .Z(new_n19139_));
  XOR2_X1    g18883(.A1(new_n19139_), .A2(new_n19022_), .Z(new_n19140_));
  NOR2_X1    g18884(.A1(new_n19137_), .A2(new_n19140_), .ZN(new_n19141_));
  NAND2_X1   g18885(.A1(new_n19137_), .A2(new_n19140_), .ZN(new_n19142_));
  INV_X1     g18886(.I(new_n19142_), .ZN(new_n19143_));
  NOR2_X1    g18887(.A1(new_n19143_), .A2(new_n19141_), .ZN(new_n19144_));
  XOR2_X1    g18888(.A1(new_n19144_), .A2(new_n19133_), .Z(new_n19145_));
  AOI22_X1   g18889(.A1(new_n10981_), .A2(\b[39] ), .B1(new_n10979_), .B2(\b[38] ), .ZN(new_n19146_));
  OAI21_X1   g18890(.A1(new_n5312_), .A2(new_n11306_), .B(new_n19146_), .ZN(new_n19147_));
  AOI21_X1   g18891(.A1(new_n6310_), .A2(new_n10984_), .B(new_n19147_), .ZN(new_n19148_));
  XOR2_X1    g18892(.A1(new_n19148_), .A2(new_n10989_), .Z(new_n19149_));
  NOR2_X1    g18893(.A1(new_n19145_), .A2(new_n19149_), .ZN(new_n19150_));
  INV_X1     g18894(.I(new_n19150_), .ZN(new_n19151_));
  NAND2_X1   g18895(.A1(new_n19145_), .A2(new_n19149_), .ZN(new_n19152_));
  NAND2_X1   g18896(.A1(new_n19151_), .A2(new_n19152_), .ZN(new_n19153_));
  XOR2_X1    g18897(.A1(new_n19153_), .A2(new_n19132_), .Z(new_n19154_));
  AOI22_X1   g18898(.A1(new_n10064_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n10062_), .ZN(new_n19155_));
  OAI21_X1   g18899(.A1(new_n6284_), .A2(new_n10399_), .B(new_n19155_), .ZN(new_n19156_));
  AOI21_X1   g18900(.A1(new_n7106_), .A2(new_n10068_), .B(new_n19156_), .ZN(new_n19157_));
  XOR2_X1    g18901(.A1(new_n19157_), .A2(new_n10057_), .Z(new_n19158_));
  NOR2_X1    g18902(.A1(new_n19041_), .A2(new_n19042_), .ZN(new_n19159_));
  AOI21_X1   g18903(.A1(new_n19041_), .A2(new_n19042_), .B(new_n19018_), .ZN(new_n19160_));
  NOR2_X1    g18904(.A1(new_n19160_), .A2(new_n19159_), .ZN(new_n19161_));
  NOR2_X1    g18905(.A1(new_n19161_), .A2(new_n19158_), .ZN(new_n19162_));
  NAND2_X1   g18906(.A1(new_n19161_), .A2(new_n19158_), .ZN(new_n19163_));
  INV_X1     g18907(.I(new_n19163_), .ZN(new_n19164_));
  NOR2_X1    g18908(.A1(new_n19164_), .A2(new_n19162_), .ZN(new_n19165_));
  XOR2_X1    g18909(.A1(new_n19165_), .A2(new_n19154_), .Z(new_n19166_));
  AOI22_X1   g18910(.A1(new_n9125_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n9123_), .ZN(new_n19167_));
  OAI21_X1   g18911(.A1(new_n6775_), .A2(new_n9470_), .B(new_n19167_), .ZN(new_n19168_));
  AOI21_X1   g18912(.A1(new_n7926_), .A2(new_n9129_), .B(new_n19168_), .ZN(new_n19169_));
  XOR2_X1    g18913(.A1(new_n19169_), .A2(\a[53] ), .Z(new_n19170_));
  NAND2_X1   g18914(.A1(new_n19166_), .A2(new_n19170_), .ZN(new_n19171_));
  OR2_X2     g18915(.A1(new_n19166_), .A2(new_n19170_), .Z(new_n19172_));
  NAND2_X1   g18916(.A1(new_n19172_), .A2(new_n19171_), .ZN(new_n19173_));
  XNOR2_X1   g18917(.A1(new_n19173_), .A2(new_n19131_), .ZN(new_n19174_));
  AOI22_X1   g18918(.A1(new_n8241_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n8246_), .ZN(new_n19175_));
  OAI21_X1   g18919(.A1(new_n7617_), .A2(new_n9114_), .B(new_n19175_), .ZN(new_n19176_));
  AOI21_X1   g18920(.A1(new_n8792_), .A2(new_n8252_), .B(new_n19176_), .ZN(new_n19177_));
  XOR2_X1    g18921(.A1(new_n19177_), .A2(\a[50] ), .Z(new_n19178_));
  INV_X1     g18922(.I(new_n19056_), .ZN(new_n19179_));
  OAI21_X1   g18923(.A1(new_n19049_), .A2(new_n19057_), .B(new_n19179_), .ZN(new_n19180_));
  NAND2_X1   g18924(.A1(new_n19180_), .A2(new_n19178_), .ZN(new_n19181_));
  OR2_X2     g18925(.A1(new_n19180_), .A2(new_n19178_), .Z(new_n19182_));
  NAND2_X1   g18926(.A1(new_n19182_), .A2(new_n19181_), .ZN(new_n19183_));
  XNOR2_X1   g18927(.A1(new_n19183_), .A2(new_n19174_), .ZN(new_n19184_));
  INV_X1     g18928(.I(new_n19184_), .ZN(new_n19185_));
  AOI22_X1   g18929(.A1(new_n7403_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n7408_), .ZN(new_n19186_));
  OAI21_X1   g18930(.A1(new_n8168_), .A2(new_n9488_), .B(new_n19186_), .ZN(new_n19187_));
  AOI21_X1   g18931(.A1(new_n8783_), .A2(new_n7414_), .B(new_n19187_), .ZN(new_n19188_));
  XOR2_X1    g18932(.A1(new_n19188_), .A2(new_n7410_), .Z(new_n19189_));
  NOR2_X1    g18933(.A1(new_n19185_), .A2(new_n19189_), .ZN(new_n19190_));
  INV_X1     g18934(.I(new_n19190_), .ZN(new_n19191_));
  NAND2_X1   g18935(.A1(new_n19185_), .A2(new_n19189_), .ZN(new_n19192_));
  NAND2_X1   g18936(.A1(new_n19191_), .A2(new_n19192_), .ZN(new_n19193_));
  XOR2_X1    g18937(.A1(new_n19193_), .A2(new_n19130_), .Z(new_n19194_));
  NOR2_X1    g18938(.A1(new_n19194_), .A2(new_n19127_), .ZN(new_n19195_));
  NAND2_X1   g18939(.A1(new_n19194_), .A2(new_n19127_), .ZN(new_n19196_));
  INV_X1     g18940(.I(new_n19196_), .ZN(new_n19197_));
  NOR2_X1    g18941(.A1(new_n19197_), .A2(new_n19195_), .ZN(new_n19198_));
  XOR2_X1    g18942(.A1(new_n19198_), .A2(new_n19123_), .Z(new_n19199_));
  INV_X1     g18943(.I(new_n19199_), .ZN(new_n19200_));
  AOI22_X1   g18944(.A1(new_n6108_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n6111_), .ZN(new_n19201_));
  OAI21_X1   g18945(.A1(new_n9972_), .A2(new_n7708_), .B(new_n19201_), .ZN(new_n19202_));
  AOI21_X1   g18946(.A1(new_n10631_), .A2(new_n6105_), .B(new_n19202_), .ZN(new_n19203_));
  XOR2_X1    g18947(.A1(new_n19203_), .A2(new_n5849_), .Z(new_n19204_));
  NOR2_X1    g18948(.A1(new_n19200_), .A2(new_n19204_), .ZN(new_n19205_));
  INV_X1     g18949(.I(new_n19205_), .ZN(new_n19206_));
  NAND2_X1   g18950(.A1(new_n19200_), .A2(new_n19204_), .ZN(new_n19207_));
  NAND2_X1   g18951(.A1(new_n19206_), .A2(new_n19207_), .ZN(new_n19208_));
  XNOR2_X1   g18952(.A1(new_n19208_), .A2(new_n19121_), .ZN(new_n19209_));
  AOI22_X1   g18953(.A1(new_n5155_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n5160_), .ZN(new_n19210_));
  OAI21_X1   g18954(.A1(new_n11195_), .A2(new_n6877_), .B(new_n19210_), .ZN(new_n19211_));
  AOI21_X1   g18955(.A1(new_n11836_), .A2(new_n5166_), .B(new_n19211_), .ZN(new_n19212_));
  XOR2_X1    g18956(.A1(new_n19212_), .A2(\a[38] ), .Z(new_n19213_));
  INV_X1     g18957(.I(new_n19084_), .ZN(new_n19214_));
  OAI21_X1   g18958(.A1(new_n19078_), .A2(new_n19085_), .B(new_n19214_), .ZN(new_n19215_));
  NAND2_X1   g18959(.A1(new_n19215_), .A2(new_n19213_), .ZN(new_n19216_));
  OR2_X2     g18960(.A1(new_n19215_), .A2(new_n19213_), .Z(new_n19217_));
  NAND2_X1   g18961(.A1(new_n19217_), .A2(new_n19216_), .ZN(new_n19218_));
  XNOR2_X1   g18962(.A1(new_n19209_), .A2(new_n19218_), .ZN(new_n19219_));
  NOR2_X1    g18963(.A1(new_n19219_), .A2(new_n19120_), .ZN(new_n19220_));
  NAND2_X1   g18964(.A1(new_n19219_), .A2(new_n19120_), .ZN(new_n19221_));
  INV_X1     g18965(.I(new_n19221_), .ZN(new_n19222_));
  NOR2_X1    g18966(.A1(new_n19222_), .A2(new_n19220_), .ZN(new_n19223_));
  XNOR2_X1   g18967(.A1(new_n19223_), .A2(new_n19115_), .ZN(new_n19224_));
  NOR2_X1    g18968(.A1(new_n19224_), .A2(new_n19114_), .ZN(new_n19225_));
  INV_X1     g18969(.I(new_n19225_), .ZN(new_n19226_));
  NAND2_X1   g18970(.A1(new_n19224_), .A2(new_n19114_), .ZN(new_n19227_));
  AND2_X2    g18971(.A1(new_n19226_), .A2(new_n19227_), .Z(new_n19228_));
  INV_X1     g18972(.I(new_n19228_), .ZN(new_n19229_));
  AOI21_X1   g18973(.A1(new_n19108_), .A2(new_n19104_), .B(new_n19229_), .ZN(new_n19230_));
  AOI21_X1   g18974(.A1(new_n18978_), .A2(new_n18973_), .B(new_n18969_), .ZN(new_n19231_));
  NOR3_X1    g18975(.A1(new_n19231_), .A2(new_n18979_), .A3(new_n19106_), .ZN(new_n19232_));
  NOR3_X1    g18976(.A1(new_n19232_), .A2(new_n19103_), .A3(new_n19228_), .ZN(new_n19233_));
  NOR2_X1    g18977(.A1(new_n19233_), .A2(new_n19230_), .ZN(\f[96] ));
  OAI22_X1   g18978(.A1(new_n6099_), .A2(new_n12796_), .B1(new_n12800_), .B2(new_n4454_), .ZN(new_n19235_));
  AOI21_X1   g18979(.A1(new_n13973_), .A2(new_n4699_), .B(new_n19235_), .ZN(new_n19236_));
  XOR2_X1    g18980(.A1(new_n19236_), .A2(new_n4446_), .Z(new_n19237_));
  INV_X1     g18981(.I(new_n19237_), .ZN(new_n19238_));
  INV_X1     g18982(.I(new_n19216_), .ZN(new_n19239_));
  AOI21_X1   g18983(.A1(new_n19209_), .A2(new_n19217_), .B(new_n19239_), .ZN(new_n19240_));
  INV_X1     g18984(.I(new_n19240_), .ZN(new_n19241_));
  AOI21_X1   g18985(.A1(new_n19121_), .A2(new_n19207_), .B(new_n19205_), .ZN(new_n19242_));
  OAI22_X1   g18986(.A1(new_n12148_), .A2(new_n6126_), .B1(new_n6129_), .B2(new_n12147_), .ZN(new_n19243_));
  AOI21_X1   g18987(.A1(\b[59] ), .A2(new_n5420_), .B(new_n19243_), .ZN(new_n19244_));
  OAI21_X1   g18988(.A1(new_n13110_), .A2(new_n6124_), .B(new_n19244_), .ZN(new_n19245_));
  XOR2_X1    g18989(.A1(new_n19245_), .A2(\a[38] ), .Z(new_n19246_));
  NOR2_X1    g18990(.A1(new_n19242_), .A2(new_n19246_), .ZN(new_n19247_));
  INV_X1     g18991(.I(new_n19247_), .ZN(new_n19248_));
  NAND2_X1   g18992(.A1(new_n19242_), .A2(new_n19246_), .ZN(new_n19249_));
  NAND2_X1   g18993(.A1(new_n19248_), .A2(new_n19249_), .ZN(new_n19250_));
  AOI22_X1   g18994(.A1(new_n6108_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n6111_), .ZN(new_n19251_));
  OAI21_X1   g18995(.A1(new_n10308_), .A2(new_n7708_), .B(new_n19251_), .ZN(new_n19252_));
  AOI21_X1   g18996(.A1(new_n12164_), .A2(new_n6105_), .B(new_n19252_), .ZN(new_n19253_));
  XOR2_X1    g18997(.A1(new_n19253_), .A2(new_n5849_), .Z(new_n19254_));
  INV_X1     g18998(.I(new_n19254_), .ZN(new_n19255_));
  AOI21_X1   g18999(.A1(new_n19123_), .A2(new_n19196_), .B(new_n19195_), .ZN(new_n19256_));
  INV_X1     g19000(.I(new_n19256_), .ZN(new_n19257_));
  AOI21_X1   g19001(.A1(new_n19130_), .A2(new_n19192_), .B(new_n19190_), .ZN(new_n19258_));
  INV_X1     g19002(.I(new_n19258_), .ZN(new_n19259_));
  AOI22_X1   g19003(.A1(new_n7403_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n7408_), .ZN(new_n19260_));
  OAI21_X1   g19004(.A1(new_n8500_), .A2(new_n9488_), .B(new_n19260_), .ZN(new_n19261_));
  AOI21_X1   g19005(.A1(new_n9987_), .A2(new_n7414_), .B(new_n19261_), .ZN(new_n19262_));
  XOR2_X1    g19006(.A1(new_n19262_), .A2(new_n7410_), .Z(new_n19263_));
  AOI22_X1   g19007(.A1(new_n9125_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n9123_), .ZN(new_n19264_));
  OAI21_X1   g19008(.A1(new_n7074_), .A2(new_n9470_), .B(new_n19264_), .ZN(new_n19265_));
  AOI21_X1   g19009(.A1(new_n9337_), .A2(new_n9129_), .B(new_n19265_), .ZN(new_n19266_));
  XOR2_X1    g19010(.A1(new_n19266_), .A2(new_n9133_), .Z(new_n19267_));
  INV_X1     g19011(.I(new_n19267_), .ZN(new_n19268_));
  INV_X1     g19012(.I(new_n19132_), .ZN(new_n19269_));
  AOI21_X1   g19013(.A1(new_n19269_), .A2(new_n19152_), .B(new_n19150_), .ZN(new_n19270_));
  INV_X1     g19014(.I(new_n19270_), .ZN(new_n19271_));
  AOI22_X1   g19015(.A1(new_n10981_), .A2(\b[40] ), .B1(new_n10979_), .B2(\b[39] ), .ZN(new_n19272_));
  OAI21_X1   g19016(.A1(new_n5341_), .A2(new_n11306_), .B(new_n19272_), .ZN(new_n19273_));
  AOI21_X1   g19017(.A1(new_n5793_), .A2(new_n10984_), .B(new_n19273_), .ZN(new_n19274_));
  XOR2_X1    g19018(.A1(new_n19274_), .A2(new_n10989_), .Z(new_n19275_));
  NOR2_X1    g19019(.A1(new_n19143_), .A2(new_n19133_), .ZN(new_n19276_));
  NOR2_X1    g19020(.A1(new_n19276_), .A2(new_n19141_), .ZN(new_n19277_));
  INV_X1     g19021(.I(new_n19277_), .ZN(new_n19278_));
  OAI22_X1   g19022(.A1(new_n13224_), .A2(new_n5312_), .B1(new_n4886_), .B2(new_n11923_), .ZN(new_n19279_));
  AOI21_X1   g19023(.A1(\b[35] ), .A2(new_n13223_), .B(new_n19279_), .ZN(new_n19280_));
  OAI21_X1   g19024(.A1(new_n5322_), .A2(new_n11930_), .B(new_n19280_), .ZN(new_n19281_));
  XOR2_X1    g19025(.A1(new_n19281_), .A2(new_n12312_), .Z(new_n19282_));
  OAI21_X1   g19026(.A1(\a[32] ), .A2(new_n19138_), .B(new_n19022_), .ZN(new_n19283_));
  INV_X1     g19027(.I(new_n19283_), .ZN(new_n19284_));
  AOI21_X1   g19028(.A1(\a[32] ), .A2(new_n19138_), .B(new_n19284_), .ZN(new_n19285_));
  AOI22_X1   g19029(.A1(new_n12922_), .A2(\b[34] ), .B1(\b[33] ), .B2(new_n12923_), .ZN(new_n19286_));
  NAND2_X1   g19030(.A1(new_n19285_), .A2(new_n19286_), .ZN(new_n19287_));
  OR2_X2     g19031(.A1(new_n19285_), .A2(new_n19286_), .Z(new_n19288_));
  NAND2_X1   g19032(.A1(new_n19288_), .A2(new_n19287_), .ZN(new_n19289_));
  XNOR2_X1   g19033(.A1(new_n19282_), .A2(new_n19289_), .ZN(new_n19290_));
  NOR2_X1    g19034(.A1(new_n19278_), .A2(new_n19290_), .ZN(new_n19291_));
  INV_X1     g19035(.I(new_n19291_), .ZN(new_n19292_));
  NAND2_X1   g19036(.A1(new_n19278_), .A2(new_n19290_), .ZN(new_n19293_));
  NAND2_X1   g19037(.A1(new_n19292_), .A2(new_n19293_), .ZN(new_n19294_));
  XOR2_X1    g19038(.A1(new_n19294_), .A2(new_n19275_), .Z(new_n19295_));
  INV_X1     g19039(.I(new_n19295_), .ZN(new_n19296_));
  OAI22_X1   g19040(.A1(new_n11298_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n11297_), .ZN(new_n19297_));
  AOI21_X1   g19041(.A1(\b[41] ), .A2(new_n11296_), .B(new_n19297_), .ZN(new_n19298_));
  OAI21_X1   g19042(.A1(new_n6785_), .A2(new_n10069_), .B(new_n19298_), .ZN(new_n19299_));
  XOR2_X1    g19043(.A1(new_n19299_), .A2(\a[56] ), .Z(new_n19300_));
  NOR2_X1    g19044(.A1(new_n19296_), .A2(new_n19300_), .ZN(new_n19301_));
  INV_X1     g19045(.I(new_n19301_), .ZN(new_n19302_));
  NAND2_X1   g19046(.A1(new_n19296_), .A2(new_n19300_), .ZN(new_n19303_));
  NAND2_X1   g19047(.A1(new_n19302_), .A2(new_n19303_), .ZN(new_n19304_));
  XOR2_X1    g19048(.A1(new_n19304_), .A2(new_n19271_), .Z(new_n19305_));
  AOI21_X1   g19049(.A1(new_n19154_), .A2(new_n19163_), .B(new_n19162_), .ZN(new_n19306_));
  NOR2_X1    g19050(.A1(new_n19305_), .A2(new_n19306_), .ZN(new_n19307_));
  INV_X1     g19051(.I(new_n19307_), .ZN(new_n19308_));
  NAND2_X1   g19052(.A1(new_n19305_), .A2(new_n19306_), .ZN(new_n19309_));
  NAND2_X1   g19053(.A1(new_n19308_), .A2(new_n19309_), .ZN(new_n19310_));
  XOR2_X1    g19054(.A1(new_n19310_), .A2(new_n19268_), .Z(new_n19311_));
  INV_X1     g19055(.I(new_n19171_), .ZN(new_n19312_));
  AOI21_X1   g19056(.A1(new_n19131_), .A2(new_n19172_), .B(new_n19312_), .ZN(new_n19313_));
  OAI22_X1   g19057(.A1(new_n9461_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n9462_), .ZN(new_n19314_));
  AOI21_X1   g19058(.A1(\b[47] ), .A2(new_n8575_), .B(new_n19314_), .ZN(new_n19315_));
  OAI21_X1   g19059(.A1(new_n9050_), .A2(new_n9460_), .B(new_n19315_), .ZN(new_n19316_));
  XOR2_X1    g19060(.A1(new_n19316_), .A2(\a[50] ), .Z(new_n19317_));
  NOR2_X1    g19061(.A1(new_n19313_), .A2(new_n19317_), .ZN(new_n19318_));
  NAND2_X1   g19062(.A1(new_n19313_), .A2(new_n19317_), .ZN(new_n19319_));
  INV_X1     g19063(.I(new_n19319_), .ZN(new_n19320_));
  NOR2_X1    g19064(.A1(new_n19320_), .A2(new_n19318_), .ZN(new_n19321_));
  XOR2_X1    g19065(.A1(new_n19321_), .A2(new_n19311_), .Z(new_n19322_));
  NAND2_X1   g19066(.A1(new_n19182_), .A2(new_n19174_), .ZN(new_n19323_));
  AND2_X2    g19067(.A1(new_n19323_), .A2(new_n19181_), .Z(new_n19324_));
  XOR2_X1    g19068(.A1(new_n19322_), .A2(new_n19324_), .Z(new_n19325_));
  XOR2_X1    g19069(.A1(new_n19325_), .A2(new_n19263_), .Z(new_n19326_));
  AOI22_X1   g19070(.A1(new_n6569_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n6574_), .ZN(new_n19327_));
  OAI21_X1   g19071(.A1(new_n9376_), .A2(new_n8565_), .B(new_n19327_), .ZN(new_n19328_));
  AOI21_X1   g19072(.A1(new_n9979_), .A2(new_n6579_), .B(new_n19328_), .ZN(new_n19329_));
  XOR2_X1    g19073(.A1(new_n19329_), .A2(new_n6567_), .Z(new_n19330_));
  NOR2_X1    g19074(.A1(new_n19326_), .A2(new_n19330_), .ZN(new_n19331_));
  NAND2_X1   g19075(.A1(new_n19326_), .A2(new_n19330_), .ZN(new_n19332_));
  INV_X1     g19076(.I(new_n19332_), .ZN(new_n19333_));
  NOR2_X1    g19077(.A1(new_n19333_), .A2(new_n19331_), .ZN(new_n19334_));
  XOR2_X1    g19078(.A1(new_n19334_), .A2(new_n19259_), .Z(new_n19335_));
  NOR2_X1    g19079(.A1(new_n19335_), .A2(new_n19257_), .ZN(new_n19336_));
  INV_X1     g19080(.I(new_n19336_), .ZN(new_n19337_));
  NAND2_X1   g19081(.A1(new_n19335_), .A2(new_n19257_), .ZN(new_n19338_));
  NAND2_X1   g19082(.A1(new_n19337_), .A2(new_n19338_), .ZN(new_n19339_));
  XOR2_X1    g19083(.A1(new_n19339_), .A2(new_n19255_), .Z(new_n19340_));
  XOR2_X1    g19084(.A1(new_n19250_), .A2(new_n19340_), .Z(new_n19341_));
  NOR2_X1    g19085(.A1(new_n19341_), .A2(new_n19241_), .ZN(new_n19342_));
  INV_X1     g19086(.I(new_n19342_), .ZN(new_n19343_));
  NAND2_X1   g19087(.A1(new_n19341_), .A2(new_n19241_), .ZN(new_n19344_));
  NAND2_X1   g19088(.A1(new_n19343_), .A2(new_n19344_), .ZN(new_n19345_));
  XOR2_X1    g19089(.A1(new_n19345_), .A2(new_n19238_), .Z(new_n19346_));
  INV_X1     g19090(.I(new_n19346_), .ZN(new_n19347_));
  OAI21_X1   g19091(.A1(new_n19115_), .A2(new_n19220_), .B(new_n19221_), .ZN(new_n19348_));
  INV_X1     g19092(.I(new_n19348_), .ZN(new_n19349_));
  OAI21_X1   g19093(.A1(new_n19230_), .A2(new_n19225_), .B(new_n19349_), .ZN(new_n19350_));
  OAI21_X1   g19094(.A1(new_n19232_), .A2(new_n19103_), .B(new_n19228_), .ZN(new_n19351_));
  NAND3_X1   g19095(.A1(new_n19351_), .A2(new_n19226_), .A3(new_n19348_), .ZN(new_n19352_));
  NAND2_X1   g19096(.A1(new_n19352_), .A2(new_n19350_), .ZN(new_n19353_));
  XOR2_X1    g19097(.A1(new_n19353_), .A2(new_n19347_), .Z(\f[97] ));
  NOR3_X1    g19098(.A1(new_n19230_), .A2(new_n19225_), .A3(new_n19349_), .ZN(new_n19355_));
  AOI21_X1   g19099(.A1(new_n19347_), .A2(new_n19350_), .B(new_n19355_), .ZN(new_n19356_));
  OAI21_X1   g19100(.A1(new_n19237_), .A2(new_n19342_), .B(new_n19344_), .ZN(new_n19357_));
  INV_X1     g19101(.I(new_n19357_), .ZN(new_n19358_));
  AOI22_X1   g19102(.A1(new_n13460_), .A2(new_n4699_), .B1(\b[63] ), .B2(new_n4706_), .ZN(new_n19359_));
  AOI22_X1   g19103(.A1(new_n5155_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n5160_), .ZN(new_n19360_));
  OAI21_X1   g19104(.A1(new_n12147_), .A2(new_n6877_), .B(new_n19360_), .ZN(new_n19361_));
  AOI21_X1   g19105(.A1(new_n13444_), .A2(new_n5166_), .B(new_n19361_), .ZN(new_n19362_));
  XOR2_X1    g19106(.A1(new_n19362_), .A2(new_n5162_), .Z(new_n19363_));
  INV_X1     g19107(.I(new_n19363_), .ZN(new_n19364_));
  AOI22_X1   g19108(.A1(new_n6569_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n6574_), .ZN(new_n19365_));
  OAI21_X1   g19109(.A1(new_n9942_), .A2(new_n8565_), .B(new_n19365_), .ZN(new_n19366_));
  AOI21_X1   g19110(.A1(new_n10318_), .A2(new_n6579_), .B(new_n19366_), .ZN(new_n19367_));
  XOR2_X1    g19111(.A1(new_n19367_), .A2(new_n6567_), .Z(new_n19368_));
  INV_X1     g19112(.I(new_n19263_), .ZN(new_n19369_));
  NOR2_X1    g19113(.A1(new_n19322_), .A2(new_n19324_), .ZN(new_n19370_));
  NAND2_X1   g19114(.A1(new_n19322_), .A2(new_n19324_), .ZN(new_n19371_));
  AOI21_X1   g19115(.A1(new_n19369_), .A2(new_n19371_), .B(new_n19370_), .ZN(new_n19372_));
  INV_X1     g19116(.I(new_n19372_), .ZN(new_n19373_));
  OAI22_X1   g19117(.A1(new_n9032_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n9376_), .ZN(new_n19374_));
  AOI21_X1   g19118(.A1(\b[51] ), .A2(new_n7719_), .B(new_n19374_), .ZN(new_n19375_));
  OAI21_X1   g19119(.A1(new_n9385_), .A2(new_n8585_), .B(new_n19375_), .ZN(new_n19376_));
  XOR2_X1    g19120(.A1(new_n19376_), .A2(new_n7410_), .Z(new_n19377_));
  AOI22_X1   g19121(.A1(new_n8241_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n8246_), .ZN(new_n19378_));
  OAI21_X1   g19122(.A1(new_n8127_), .A2(new_n9114_), .B(new_n19378_), .ZN(new_n19379_));
  AOI21_X1   g19123(.A1(new_n9684_), .A2(new_n8252_), .B(new_n19379_), .ZN(new_n19380_));
  XOR2_X1    g19124(.A1(new_n19380_), .A2(new_n8248_), .Z(new_n19381_));
  AOI22_X1   g19125(.A1(new_n10064_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n10062_), .ZN(new_n19382_));
  OAI21_X1   g19126(.A1(new_n6490_), .A2(new_n10399_), .B(new_n19382_), .ZN(new_n19383_));
  AOI21_X1   g19127(.A1(new_n7906_), .A2(new_n10068_), .B(new_n19383_), .ZN(new_n19384_));
  XOR2_X1    g19128(.A1(new_n19384_), .A2(new_n10057_), .Z(new_n19385_));
  INV_X1     g19129(.I(new_n19385_), .ZN(new_n19386_));
  OAI21_X1   g19130(.A1(new_n19275_), .A2(new_n19291_), .B(new_n19293_), .ZN(new_n19387_));
  INV_X1     g19131(.I(new_n19387_), .ZN(new_n19388_));
  NAND2_X1   g19132(.A1(new_n19282_), .A2(new_n19287_), .ZN(new_n19389_));
  NAND2_X1   g19133(.A1(new_n19389_), .A2(new_n19288_), .ZN(new_n19390_));
  AOI22_X1   g19134(.A1(new_n12922_), .A2(\b[35] ), .B1(\b[34] ), .B2(new_n12923_), .ZN(new_n19391_));
  INV_X1     g19135(.I(new_n19391_), .ZN(new_n19392_));
  NOR2_X1    g19136(.A1(new_n19392_), .A2(new_n19286_), .ZN(new_n19393_));
  NAND2_X1   g19137(.A1(new_n19392_), .A2(new_n19286_), .ZN(new_n19394_));
  INV_X1     g19138(.I(new_n19394_), .ZN(new_n19395_));
  NOR2_X1    g19139(.A1(new_n19395_), .A2(new_n19393_), .ZN(new_n19396_));
  XNOR2_X1   g19140(.A1(new_n19390_), .A2(new_n19396_), .ZN(new_n19397_));
  INV_X1     g19141(.I(new_n19397_), .ZN(new_n19398_));
  OAI22_X1   g19142(.A1(new_n12306_), .A2(new_n6285_), .B1(new_n12305_), .B2(new_n6284_), .ZN(new_n19399_));
  AOI21_X1   g19143(.A1(\b[39] ), .A2(new_n12304_), .B(new_n19399_), .ZN(new_n19400_));
  OAI21_X1   g19144(.A1(new_n6299_), .A2(new_n10985_), .B(new_n19400_), .ZN(new_n19401_));
  XOR2_X1    g19145(.A1(new_n19401_), .A2(\a[59] ), .Z(new_n19402_));
  AOI22_X1   g19146(.A1(new_n11926_), .A2(\b[38] ), .B1(new_n11924_), .B2(\b[37] ), .ZN(new_n19403_));
  OAI21_X1   g19147(.A1(new_n4886_), .A2(new_n12317_), .B(new_n19403_), .ZN(new_n19404_));
  AOI21_X1   g19148(.A1(new_n5351_), .A2(new_n11929_), .B(new_n19404_), .ZN(new_n19405_));
  XOR2_X1    g19149(.A1(new_n19405_), .A2(new_n12312_), .Z(new_n19406_));
  NOR2_X1    g19150(.A1(new_n19402_), .A2(new_n19406_), .ZN(new_n19407_));
  INV_X1     g19151(.I(new_n19407_), .ZN(new_n19408_));
  NAND2_X1   g19152(.A1(new_n19402_), .A2(new_n19406_), .ZN(new_n19409_));
  NAND2_X1   g19153(.A1(new_n19408_), .A2(new_n19409_), .ZN(new_n19410_));
  XOR2_X1    g19154(.A1(new_n19410_), .A2(new_n19398_), .Z(new_n19411_));
  NOR2_X1    g19155(.A1(new_n19411_), .A2(new_n19388_), .ZN(new_n19412_));
  INV_X1     g19156(.I(new_n19412_), .ZN(new_n19413_));
  NAND2_X1   g19157(.A1(new_n19411_), .A2(new_n19388_), .ZN(new_n19414_));
  NAND2_X1   g19158(.A1(new_n19413_), .A2(new_n19414_), .ZN(new_n19415_));
  XOR2_X1    g19159(.A1(new_n19415_), .A2(new_n19386_), .Z(new_n19416_));
  AOI22_X1   g19160(.A1(new_n9125_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n9123_), .ZN(new_n19417_));
  OAI21_X1   g19161(.A1(new_n7096_), .A2(new_n9470_), .B(new_n19417_), .ZN(new_n19418_));
  AOI21_X1   g19162(.A1(new_n7649_), .A2(new_n9129_), .B(new_n19418_), .ZN(new_n19419_));
  XOR2_X1    g19163(.A1(new_n19419_), .A2(new_n9133_), .Z(new_n19420_));
  AOI21_X1   g19164(.A1(new_n19271_), .A2(new_n19303_), .B(new_n19301_), .ZN(new_n19421_));
  NOR2_X1    g19165(.A1(new_n19420_), .A2(new_n19421_), .ZN(new_n19422_));
  AND2_X2    g19166(.A1(new_n19420_), .A2(new_n19421_), .Z(new_n19423_));
  NOR2_X1    g19167(.A1(new_n19423_), .A2(new_n19422_), .ZN(new_n19424_));
  XOR2_X1    g19168(.A1(new_n19416_), .A2(new_n19424_), .Z(new_n19425_));
  AOI21_X1   g19169(.A1(new_n19268_), .A2(new_n19309_), .B(new_n19307_), .ZN(new_n19426_));
  NOR2_X1    g19170(.A1(new_n19425_), .A2(new_n19426_), .ZN(new_n19427_));
  INV_X1     g19171(.I(new_n19427_), .ZN(new_n19428_));
  NAND2_X1   g19172(.A1(new_n19425_), .A2(new_n19426_), .ZN(new_n19429_));
  NAND2_X1   g19173(.A1(new_n19428_), .A2(new_n19429_), .ZN(new_n19430_));
  XOR2_X1    g19174(.A1(new_n19430_), .A2(new_n19381_), .Z(new_n19431_));
  INV_X1     g19175(.I(new_n19431_), .ZN(new_n19432_));
  INV_X1     g19176(.I(new_n19311_), .ZN(new_n19433_));
  AOI21_X1   g19177(.A1(new_n19433_), .A2(new_n19319_), .B(new_n19318_), .ZN(new_n19434_));
  NOR2_X1    g19178(.A1(new_n19432_), .A2(new_n19434_), .ZN(new_n19435_));
  INV_X1     g19179(.I(new_n19435_), .ZN(new_n19436_));
  NAND2_X1   g19180(.A1(new_n19432_), .A2(new_n19434_), .ZN(new_n19437_));
  NAND2_X1   g19181(.A1(new_n19436_), .A2(new_n19437_), .ZN(new_n19438_));
  XNOR2_X1   g19182(.A1(new_n19438_), .A2(new_n19377_), .ZN(new_n19439_));
  NOR2_X1    g19183(.A1(new_n19439_), .A2(new_n19373_), .ZN(new_n19440_));
  INV_X1     g19184(.I(new_n19440_), .ZN(new_n19441_));
  NAND2_X1   g19185(.A1(new_n19439_), .A2(new_n19373_), .ZN(new_n19442_));
  NAND2_X1   g19186(.A1(new_n19441_), .A2(new_n19442_), .ZN(new_n19443_));
  XNOR2_X1   g19187(.A1(new_n19443_), .A2(new_n19368_), .ZN(new_n19444_));
  OAI22_X1   g19188(.A1(new_n5852_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n5857_), .ZN(new_n19445_));
  AOI21_X1   g19189(.A1(\b[57] ), .A2(new_n6115_), .B(new_n19445_), .ZN(new_n19446_));
  OAI21_X1   g19190(.A1(new_n12203_), .A2(new_n5861_), .B(new_n19446_), .ZN(new_n19447_));
  XOR2_X1    g19191(.A1(new_n19447_), .A2(\a[41] ), .Z(new_n19448_));
  AOI21_X1   g19192(.A1(new_n19259_), .A2(new_n19332_), .B(new_n19331_), .ZN(new_n19449_));
  NOR2_X1    g19193(.A1(new_n19449_), .A2(new_n19448_), .ZN(new_n19450_));
  AND2_X2    g19194(.A1(new_n19449_), .A2(new_n19448_), .Z(new_n19451_));
  NOR2_X1    g19195(.A1(new_n19451_), .A2(new_n19450_), .ZN(new_n19452_));
  XOR2_X1    g19196(.A1(new_n19444_), .A2(new_n19452_), .Z(new_n19453_));
  OAI21_X1   g19197(.A1(new_n19254_), .A2(new_n19336_), .B(new_n19338_), .ZN(new_n19454_));
  INV_X1     g19198(.I(new_n19454_), .ZN(new_n19455_));
  NOR2_X1    g19199(.A1(new_n19453_), .A2(new_n19455_), .ZN(new_n19456_));
  INV_X1     g19200(.I(new_n19456_), .ZN(new_n19457_));
  NAND2_X1   g19201(.A1(new_n19453_), .A2(new_n19455_), .ZN(new_n19458_));
  NAND2_X1   g19202(.A1(new_n19457_), .A2(new_n19458_), .ZN(new_n19459_));
  XOR2_X1    g19203(.A1(new_n19459_), .A2(new_n19364_), .Z(new_n19460_));
  XOR2_X1    g19204(.A1(new_n19460_), .A2(new_n19359_), .Z(new_n19461_));
  INV_X1     g19205(.I(new_n19340_), .ZN(new_n19462_));
  NAND2_X1   g19206(.A1(new_n19462_), .A2(new_n19249_), .ZN(new_n19463_));
  NAND2_X1   g19207(.A1(new_n19463_), .A2(new_n19248_), .ZN(new_n19464_));
  XOR2_X1    g19208(.A1(new_n19464_), .A2(\a[35] ), .Z(new_n19465_));
  XOR2_X1    g19209(.A1(new_n19461_), .A2(new_n19465_), .Z(new_n19466_));
  NOR2_X1    g19210(.A1(new_n19466_), .A2(new_n19358_), .ZN(new_n19467_));
  NAND2_X1   g19211(.A1(new_n19466_), .A2(new_n19358_), .ZN(new_n19468_));
  INV_X1     g19212(.I(new_n19468_), .ZN(new_n19469_));
  NOR2_X1    g19213(.A1(new_n19469_), .A2(new_n19467_), .ZN(new_n19470_));
  XOR2_X1    g19214(.A1(new_n19356_), .A2(new_n19470_), .Z(\f[98] ));
  INV_X1     g19215(.I(new_n19467_), .ZN(new_n19472_));
  OAI21_X1   g19216(.A1(new_n19356_), .A2(new_n19469_), .B(new_n19472_), .ZN(new_n19473_));
  AOI22_X1   g19217(.A1(new_n5155_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n5160_), .ZN(new_n19474_));
  OAI21_X1   g19218(.A1(new_n12148_), .A2(new_n6877_), .B(new_n19474_), .ZN(new_n19475_));
  AOI21_X1   g19219(.A1(new_n12811_), .A2(new_n5166_), .B(new_n19475_), .ZN(new_n19476_));
  XOR2_X1    g19220(.A1(new_n19476_), .A2(new_n5162_), .Z(new_n19477_));
  AOI21_X1   g19221(.A1(new_n19364_), .A2(new_n19458_), .B(new_n19456_), .ZN(new_n19478_));
  OAI21_X1   g19222(.A1(new_n19368_), .A2(new_n19440_), .B(new_n19442_), .ZN(new_n19479_));
  AOI21_X1   g19223(.A1(new_n19377_), .A2(new_n19437_), .B(new_n19435_), .ZN(new_n19480_));
  AOI22_X1   g19224(.A1(new_n7403_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n7408_), .ZN(new_n19481_));
  OAI21_X1   g19225(.A1(new_n9032_), .A2(new_n9488_), .B(new_n19481_), .ZN(new_n19482_));
  AOI21_X1   g19226(.A1(new_n10884_), .A2(new_n7414_), .B(new_n19482_), .ZN(new_n19483_));
  XOR2_X1    g19227(.A1(new_n19483_), .A2(new_n7410_), .Z(new_n19484_));
  INV_X1     g19228(.I(new_n19484_), .ZN(new_n19485_));
  INV_X1     g19229(.I(new_n19381_), .ZN(new_n19486_));
  AOI21_X1   g19230(.A1(new_n19486_), .A2(new_n19429_), .B(new_n19427_), .ZN(new_n19487_));
  AOI21_X1   g19231(.A1(new_n19386_), .A2(new_n19414_), .B(new_n19412_), .ZN(new_n19488_));
  INV_X1     g19232(.I(new_n19488_), .ZN(new_n19489_));
  INV_X1     g19233(.I(new_n19393_), .ZN(new_n19490_));
  AOI21_X1   g19234(.A1(new_n19390_), .A2(new_n19490_), .B(new_n19395_), .ZN(new_n19491_));
  AOI22_X1   g19235(.A1(new_n11926_), .A2(\b[39] ), .B1(new_n11924_), .B2(\b[38] ), .ZN(new_n19492_));
  OAI21_X1   g19236(.A1(new_n5312_), .A2(new_n12317_), .B(new_n19492_), .ZN(new_n19493_));
  AOI21_X1   g19237(.A1(new_n6310_), .A2(new_n11929_), .B(new_n19493_), .ZN(new_n19494_));
  XOR2_X1    g19238(.A1(new_n19494_), .A2(new_n12312_), .Z(new_n19495_));
  INV_X1     g19239(.I(new_n19495_), .ZN(new_n19496_));
  AOI22_X1   g19240(.A1(new_n12922_), .A2(\b[36] ), .B1(\b[35] ), .B2(new_n12923_), .ZN(new_n19497_));
  NAND2_X1   g19241(.A1(new_n19497_), .A2(\a[35] ), .ZN(new_n19498_));
  OR2_X2     g19242(.A1(new_n19497_), .A2(\a[35] ), .Z(new_n19499_));
  NAND2_X1   g19243(.A1(new_n19499_), .A2(new_n19498_), .ZN(new_n19500_));
  XOR2_X1    g19244(.A1(new_n19500_), .A2(new_n19392_), .Z(new_n19501_));
  NOR2_X1    g19245(.A1(new_n19496_), .A2(new_n19501_), .ZN(new_n19502_));
  INV_X1     g19246(.I(new_n19502_), .ZN(new_n19503_));
  NAND2_X1   g19247(.A1(new_n19496_), .A2(new_n19501_), .ZN(new_n19504_));
  NAND2_X1   g19248(.A1(new_n19503_), .A2(new_n19504_), .ZN(new_n19505_));
  XOR2_X1    g19249(.A1(new_n19505_), .A2(new_n19491_), .Z(new_n19506_));
  AOI22_X1   g19250(.A1(new_n10981_), .A2(\b[42] ), .B1(new_n10979_), .B2(\b[41] ), .ZN(new_n19507_));
  OAI21_X1   g19251(.A1(new_n6284_), .A2(new_n11306_), .B(new_n19507_), .ZN(new_n19508_));
  AOI21_X1   g19252(.A1(new_n7106_), .A2(new_n10984_), .B(new_n19508_), .ZN(new_n19509_));
  XOR2_X1    g19253(.A1(new_n19509_), .A2(new_n10989_), .Z(new_n19510_));
  INV_X1     g19254(.I(new_n19510_), .ZN(new_n19511_));
  NAND2_X1   g19255(.A1(new_n19409_), .A2(new_n19398_), .ZN(new_n19512_));
  NAND2_X1   g19256(.A1(new_n19512_), .A2(new_n19408_), .ZN(new_n19513_));
  NAND2_X1   g19257(.A1(new_n19513_), .A2(new_n19511_), .ZN(new_n19514_));
  NAND3_X1   g19258(.A1(new_n19512_), .A2(new_n19408_), .A3(new_n19510_), .ZN(new_n19515_));
  NAND2_X1   g19259(.A1(new_n19514_), .A2(new_n19515_), .ZN(new_n19516_));
  XOR2_X1    g19260(.A1(new_n19516_), .A2(new_n19506_), .Z(new_n19517_));
  AOI22_X1   g19261(.A1(new_n10064_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n10062_), .ZN(new_n19518_));
  OAI21_X1   g19262(.A1(new_n6775_), .A2(new_n10399_), .B(new_n19518_), .ZN(new_n19519_));
  AOI21_X1   g19263(.A1(new_n7926_), .A2(new_n10068_), .B(new_n19519_), .ZN(new_n19520_));
  XOR2_X1    g19264(.A1(new_n19520_), .A2(new_n10057_), .Z(new_n19521_));
  NOR2_X1    g19265(.A1(new_n19517_), .A2(new_n19521_), .ZN(new_n19522_));
  NAND2_X1   g19266(.A1(new_n19517_), .A2(new_n19521_), .ZN(new_n19523_));
  INV_X1     g19267(.I(new_n19523_), .ZN(new_n19524_));
  NOR2_X1    g19268(.A1(new_n19524_), .A2(new_n19522_), .ZN(new_n19525_));
  XOR2_X1    g19269(.A1(new_n19525_), .A2(new_n19489_), .Z(new_n19526_));
  AOI22_X1   g19270(.A1(new_n9125_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n9123_), .ZN(new_n19527_));
  OAI21_X1   g19271(.A1(new_n7617_), .A2(new_n9470_), .B(new_n19527_), .ZN(new_n19528_));
  AOI21_X1   g19272(.A1(new_n8792_), .A2(new_n9129_), .B(new_n19528_), .ZN(new_n19529_));
  XOR2_X1    g19273(.A1(new_n19529_), .A2(\a[53] ), .Z(new_n19530_));
  INV_X1     g19274(.I(new_n19422_), .ZN(new_n19531_));
  OAI21_X1   g19275(.A1(new_n19416_), .A2(new_n19423_), .B(new_n19531_), .ZN(new_n19532_));
  NAND2_X1   g19276(.A1(new_n19532_), .A2(new_n19530_), .ZN(new_n19533_));
  OR2_X2     g19277(.A1(new_n19532_), .A2(new_n19530_), .Z(new_n19534_));
  NAND2_X1   g19278(.A1(new_n19534_), .A2(new_n19533_), .ZN(new_n19535_));
  XNOR2_X1   g19279(.A1(new_n19535_), .A2(new_n19526_), .ZN(new_n19536_));
  INV_X1     g19280(.I(new_n19536_), .ZN(new_n19537_));
  AOI22_X1   g19281(.A1(new_n8241_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n8246_), .ZN(new_n19538_));
  OAI21_X1   g19282(.A1(new_n8168_), .A2(new_n9114_), .B(new_n19538_), .ZN(new_n19539_));
  AOI21_X1   g19283(.A1(new_n8783_), .A2(new_n8252_), .B(new_n19539_), .ZN(new_n19540_));
  XOR2_X1    g19284(.A1(new_n19540_), .A2(new_n8248_), .Z(new_n19541_));
  NOR2_X1    g19285(.A1(new_n19537_), .A2(new_n19541_), .ZN(new_n19542_));
  INV_X1     g19286(.I(new_n19542_), .ZN(new_n19543_));
  NAND2_X1   g19287(.A1(new_n19537_), .A2(new_n19541_), .ZN(new_n19544_));
  NAND2_X1   g19288(.A1(new_n19543_), .A2(new_n19544_), .ZN(new_n19545_));
  XOR2_X1    g19289(.A1(new_n19545_), .A2(new_n19487_), .Z(new_n19546_));
  NOR2_X1    g19290(.A1(new_n19546_), .A2(new_n19485_), .ZN(new_n19547_));
  INV_X1     g19291(.I(new_n19547_), .ZN(new_n19548_));
  NAND2_X1   g19292(.A1(new_n19546_), .A2(new_n19485_), .ZN(new_n19549_));
  NAND2_X1   g19293(.A1(new_n19548_), .A2(new_n19549_), .ZN(new_n19550_));
  XOR2_X1    g19294(.A1(new_n19550_), .A2(new_n19480_), .Z(new_n19551_));
  AOI22_X1   g19295(.A1(new_n6569_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n6574_), .ZN(new_n19552_));
  OAI21_X1   g19296(.A1(new_n9972_), .A2(new_n8565_), .B(new_n19552_), .ZN(new_n19553_));
  AOI21_X1   g19297(.A1(new_n10631_), .A2(new_n6579_), .B(new_n19553_), .ZN(new_n19554_));
  XOR2_X1    g19298(.A1(new_n19554_), .A2(\a[44] ), .Z(new_n19555_));
  NAND2_X1   g19299(.A1(new_n19551_), .A2(new_n19555_), .ZN(new_n19556_));
  OR2_X2     g19300(.A1(new_n19551_), .A2(new_n19555_), .Z(new_n19557_));
  NAND2_X1   g19301(.A1(new_n19557_), .A2(new_n19556_), .ZN(new_n19558_));
  XNOR2_X1   g19302(.A1(new_n19558_), .A2(new_n19479_), .ZN(new_n19559_));
  AOI22_X1   g19303(.A1(new_n6108_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n6111_), .ZN(new_n19560_));
  OAI21_X1   g19304(.A1(new_n11195_), .A2(new_n7708_), .B(new_n19560_), .ZN(new_n19561_));
  AOI21_X1   g19305(.A1(new_n11836_), .A2(new_n6105_), .B(new_n19561_), .ZN(new_n19562_));
  XOR2_X1    g19306(.A1(new_n19562_), .A2(\a[41] ), .Z(new_n19563_));
  INV_X1     g19307(.I(new_n19450_), .ZN(new_n19564_));
  OAI21_X1   g19308(.A1(new_n19444_), .A2(new_n19451_), .B(new_n19564_), .ZN(new_n19565_));
  NAND2_X1   g19309(.A1(new_n19565_), .A2(new_n19563_), .ZN(new_n19566_));
  OR2_X2     g19310(.A1(new_n19565_), .A2(new_n19563_), .Z(new_n19567_));
  NAND2_X1   g19311(.A1(new_n19567_), .A2(new_n19566_), .ZN(new_n19568_));
  XOR2_X1    g19312(.A1(new_n19568_), .A2(new_n19559_), .Z(new_n19569_));
  NAND2_X1   g19313(.A1(new_n19569_), .A2(new_n19478_), .ZN(new_n19570_));
  NOR2_X1    g19314(.A1(new_n19569_), .A2(new_n19478_), .ZN(new_n19571_));
  INV_X1     g19315(.I(new_n19571_), .ZN(new_n19572_));
  NAND2_X1   g19316(.A1(new_n19572_), .A2(new_n19570_), .ZN(new_n19573_));
  XOR2_X1    g19317(.A1(new_n19573_), .A2(new_n19477_), .Z(new_n19574_));
  INV_X1     g19318(.I(new_n19460_), .ZN(new_n19575_));
  INV_X1     g19319(.I(new_n19464_), .ZN(new_n19576_));
  XOR2_X1    g19320(.A1(new_n19359_), .A2(new_n4446_), .Z(new_n19577_));
  AOI21_X1   g19321(.A1(new_n19460_), .A2(new_n19576_), .B(new_n19577_), .ZN(new_n19578_));
  AOI21_X1   g19322(.A1(new_n19575_), .A2(new_n19464_), .B(new_n19578_), .ZN(new_n19579_));
  INV_X1     g19323(.I(new_n19579_), .ZN(new_n19580_));
  NOR2_X1    g19324(.A1(new_n19574_), .A2(new_n19580_), .ZN(new_n19581_));
  INV_X1     g19325(.I(new_n19581_), .ZN(new_n19582_));
  NAND2_X1   g19326(.A1(new_n19574_), .A2(new_n19580_), .ZN(new_n19583_));
  AND2_X2    g19327(.A1(new_n19582_), .A2(new_n19583_), .Z(new_n19584_));
  INV_X1     g19328(.I(new_n19584_), .ZN(new_n19585_));
  XOR2_X1    g19329(.A1(new_n19473_), .A2(new_n19585_), .Z(\f[99] ));
  OAI22_X1   g19330(.A1(new_n6877_), .A2(new_n12796_), .B1(new_n12800_), .B2(new_n6129_), .ZN(new_n19587_));
  AOI21_X1   g19331(.A1(new_n13973_), .A2(new_n5166_), .B(new_n19587_), .ZN(new_n19588_));
  XOR2_X1    g19332(.A1(new_n19588_), .A2(new_n5162_), .Z(new_n19589_));
  INV_X1     g19333(.I(new_n19589_), .ZN(new_n19590_));
  INV_X1     g19334(.I(new_n19566_), .ZN(new_n19591_));
  AOI21_X1   g19335(.A1(new_n19559_), .A2(new_n19567_), .B(new_n19591_), .ZN(new_n19592_));
  INV_X1     g19336(.I(new_n19592_), .ZN(new_n19593_));
  AOI22_X1   g19337(.A1(new_n6569_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n6574_), .ZN(new_n19594_));
  OAI21_X1   g19338(.A1(new_n10308_), .A2(new_n8565_), .B(new_n19594_), .ZN(new_n19595_));
  AOI21_X1   g19339(.A1(new_n12164_), .A2(new_n6579_), .B(new_n19595_), .ZN(new_n19596_));
  XOR2_X1    g19340(.A1(new_n19596_), .A2(new_n6567_), .Z(new_n19597_));
  INV_X1     g19341(.I(new_n19597_), .ZN(new_n19598_));
  AOI22_X1   g19342(.A1(new_n8241_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n8246_), .ZN(new_n19599_));
  OAI21_X1   g19343(.A1(new_n8500_), .A2(new_n9114_), .B(new_n19599_), .ZN(new_n19600_));
  AOI21_X1   g19344(.A1(new_n9987_), .A2(new_n8252_), .B(new_n19600_), .ZN(new_n19601_));
  XOR2_X1    g19345(.A1(new_n19601_), .A2(new_n8248_), .Z(new_n19602_));
  AOI22_X1   g19346(.A1(new_n10064_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n10062_), .ZN(new_n19603_));
  OAI21_X1   g19347(.A1(new_n7074_), .A2(new_n10399_), .B(new_n19603_), .ZN(new_n19604_));
  AOI21_X1   g19348(.A1(new_n9337_), .A2(new_n10068_), .B(new_n19604_), .ZN(new_n19605_));
  XOR2_X1    g19349(.A1(new_n19605_), .A2(new_n10057_), .Z(new_n19606_));
  INV_X1     g19350(.I(new_n19606_), .ZN(new_n19607_));
  AOI22_X1   g19351(.A1(new_n11926_), .A2(\b[40] ), .B1(new_n11924_), .B2(\b[39] ), .ZN(new_n19608_));
  OAI21_X1   g19352(.A1(new_n5341_), .A2(new_n12317_), .B(new_n19608_), .ZN(new_n19609_));
  AOI21_X1   g19353(.A1(new_n5793_), .A2(new_n11929_), .B(new_n19609_), .ZN(new_n19610_));
  XOR2_X1    g19354(.A1(new_n19610_), .A2(new_n12312_), .Z(new_n19611_));
  NAND2_X1   g19355(.A1(new_n19499_), .A2(new_n19391_), .ZN(new_n19612_));
  NAND2_X1   g19356(.A1(new_n19612_), .A2(new_n19498_), .ZN(new_n19613_));
  AOI22_X1   g19357(.A1(new_n12922_), .A2(\b[37] ), .B1(\b[36] ), .B2(new_n12923_), .ZN(new_n19614_));
  INV_X1     g19358(.I(new_n19614_), .ZN(new_n19615_));
  XOR2_X1    g19359(.A1(new_n19613_), .A2(new_n19615_), .Z(new_n19616_));
  XOR2_X1    g19360(.A1(new_n19611_), .A2(new_n19616_), .Z(new_n19617_));
  INV_X1     g19361(.I(new_n19617_), .ZN(new_n19618_));
  OAI21_X1   g19362(.A1(new_n19491_), .A2(new_n19502_), .B(new_n19504_), .ZN(new_n19619_));
  INV_X1     g19363(.I(new_n19619_), .ZN(new_n19620_));
  OAI22_X1   g19364(.A1(new_n12306_), .A2(new_n6775_), .B1(new_n12305_), .B2(new_n6490_), .ZN(new_n19621_));
  AOI21_X1   g19365(.A1(\b[41] ), .A2(new_n12304_), .B(new_n19621_), .ZN(new_n19622_));
  OAI21_X1   g19366(.A1(new_n6785_), .A2(new_n10985_), .B(new_n19622_), .ZN(new_n19623_));
  XOR2_X1    g19367(.A1(new_n19623_), .A2(\a[59] ), .Z(new_n19624_));
  NOR2_X1    g19368(.A1(new_n19624_), .A2(new_n19620_), .ZN(new_n19625_));
  INV_X1     g19369(.I(new_n19625_), .ZN(new_n19626_));
  NAND2_X1   g19370(.A1(new_n19624_), .A2(new_n19620_), .ZN(new_n19627_));
  NAND2_X1   g19371(.A1(new_n19626_), .A2(new_n19627_), .ZN(new_n19628_));
  XOR2_X1    g19372(.A1(new_n19628_), .A2(new_n19618_), .Z(new_n19629_));
  NAND2_X1   g19373(.A1(new_n19515_), .A2(new_n19506_), .ZN(new_n19630_));
  NAND2_X1   g19374(.A1(new_n19630_), .A2(new_n19514_), .ZN(new_n19631_));
  INV_X1     g19375(.I(new_n19631_), .ZN(new_n19632_));
  NOR2_X1    g19376(.A1(new_n19629_), .A2(new_n19632_), .ZN(new_n19633_));
  INV_X1     g19377(.I(new_n19633_), .ZN(new_n19634_));
  NAND2_X1   g19378(.A1(new_n19629_), .A2(new_n19632_), .ZN(new_n19635_));
  NAND2_X1   g19379(.A1(new_n19634_), .A2(new_n19635_), .ZN(new_n19636_));
  XOR2_X1    g19380(.A1(new_n19636_), .A2(new_n19607_), .Z(new_n19637_));
  AOI21_X1   g19381(.A1(new_n19489_), .A2(new_n19523_), .B(new_n19522_), .ZN(new_n19638_));
  OAI22_X1   g19382(.A1(new_n10390_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n10389_), .ZN(new_n19639_));
  AOI21_X1   g19383(.A1(\b[47] ), .A2(new_n9471_), .B(new_n19639_), .ZN(new_n19640_));
  OAI21_X1   g19384(.A1(new_n9050_), .A2(new_n10388_), .B(new_n19640_), .ZN(new_n19641_));
  XOR2_X1    g19385(.A1(new_n19641_), .A2(\a[53] ), .Z(new_n19642_));
  NOR2_X1    g19386(.A1(new_n19642_), .A2(new_n19638_), .ZN(new_n19643_));
  NAND2_X1   g19387(.A1(new_n19642_), .A2(new_n19638_), .ZN(new_n19644_));
  INV_X1     g19388(.I(new_n19644_), .ZN(new_n19645_));
  NOR2_X1    g19389(.A1(new_n19645_), .A2(new_n19643_), .ZN(new_n19646_));
  XOR2_X1    g19390(.A1(new_n19637_), .A2(new_n19646_), .Z(new_n19647_));
  INV_X1     g19391(.I(new_n19533_), .ZN(new_n19648_));
  AOI21_X1   g19392(.A1(new_n19526_), .A2(new_n19534_), .B(new_n19648_), .ZN(new_n19649_));
  XOR2_X1    g19393(.A1(new_n19647_), .A2(new_n19649_), .Z(new_n19650_));
  XOR2_X1    g19394(.A1(new_n19650_), .A2(new_n19602_), .Z(new_n19651_));
  INV_X1     g19395(.I(new_n19651_), .ZN(new_n19652_));
  INV_X1     g19396(.I(new_n19487_), .ZN(new_n19653_));
  AOI21_X1   g19397(.A1(new_n19653_), .A2(new_n19544_), .B(new_n19542_), .ZN(new_n19654_));
  AOI22_X1   g19398(.A1(new_n7403_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n7408_), .ZN(new_n19655_));
  OAI21_X1   g19399(.A1(new_n9376_), .A2(new_n9488_), .B(new_n19655_), .ZN(new_n19656_));
  AOI21_X1   g19400(.A1(new_n9979_), .A2(new_n7414_), .B(new_n19656_), .ZN(new_n19657_));
  XOR2_X1    g19401(.A1(new_n19657_), .A2(new_n7410_), .Z(new_n19658_));
  NOR2_X1    g19402(.A1(new_n19654_), .A2(new_n19658_), .ZN(new_n19659_));
  INV_X1     g19403(.I(new_n19659_), .ZN(new_n19660_));
  NAND2_X1   g19404(.A1(new_n19654_), .A2(new_n19658_), .ZN(new_n19661_));
  NAND2_X1   g19405(.A1(new_n19660_), .A2(new_n19661_), .ZN(new_n19662_));
  XOR2_X1    g19406(.A1(new_n19662_), .A2(new_n19652_), .Z(new_n19663_));
  OAI21_X1   g19407(.A1(new_n19480_), .A2(new_n19547_), .B(new_n19549_), .ZN(new_n19664_));
  INV_X1     g19408(.I(new_n19664_), .ZN(new_n19665_));
  NOR2_X1    g19409(.A1(new_n19665_), .A2(new_n19663_), .ZN(new_n19666_));
  INV_X1     g19410(.I(new_n19666_), .ZN(new_n19667_));
  NAND2_X1   g19411(.A1(new_n19665_), .A2(new_n19663_), .ZN(new_n19668_));
  NAND2_X1   g19412(.A1(new_n19667_), .A2(new_n19668_), .ZN(new_n19669_));
  XOR2_X1    g19413(.A1(new_n19669_), .A2(new_n19598_), .Z(new_n19670_));
  INV_X1     g19414(.I(new_n19556_), .ZN(new_n19671_));
  AOI21_X1   g19415(.A1(new_n19479_), .A2(new_n19557_), .B(new_n19671_), .ZN(new_n19672_));
  OAI22_X1   g19416(.A1(new_n5852_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n5857_), .ZN(new_n19673_));
  AOI21_X1   g19417(.A1(\b[59] ), .A2(new_n6115_), .B(new_n19673_), .ZN(new_n19674_));
  OAI21_X1   g19418(.A1(new_n13110_), .A2(new_n5861_), .B(new_n19674_), .ZN(new_n19675_));
  XOR2_X1    g19419(.A1(new_n19675_), .A2(\a[41] ), .Z(new_n19676_));
  NOR2_X1    g19420(.A1(new_n19672_), .A2(new_n19676_), .ZN(new_n19677_));
  INV_X1     g19421(.I(new_n19677_), .ZN(new_n19678_));
  NAND2_X1   g19422(.A1(new_n19672_), .A2(new_n19676_), .ZN(new_n19679_));
  NAND2_X1   g19423(.A1(new_n19678_), .A2(new_n19679_), .ZN(new_n19680_));
  XOR2_X1    g19424(.A1(new_n19680_), .A2(new_n19670_), .Z(new_n19681_));
  NOR2_X1    g19425(.A1(new_n19681_), .A2(new_n19593_), .ZN(new_n19682_));
  INV_X1     g19426(.I(new_n19682_), .ZN(new_n19683_));
  NAND2_X1   g19427(.A1(new_n19681_), .A2(new_n19593_), .ZN(new_n19684_));
  NAND2_X1   g19428(.A1(new_n19683_), .A2(new_n19684_), .ZN(new_n19685_));
  XOR2_X1    g19429(.A1(new_n19685_), .A2(new_n19590_), .Z(new_n19686_));
  INV_X1     g19430(.I(new_n19477_), .ZN(new_n19687_));
  AOI21_X1   g19431(.A1(new_n19687_), .A2(new_n19570_), .B(new_n19571_), .ZN(new_n19688_));
  INV_X1     g19432(.I(new_n19688_), .ZN(new_n19689_));
  AOI21_X1   g19433(.A1(new_n19351_), .A2(new_n19226_), .B(new_n19348_), .ZN(new_n19690_));
  OAI21_X1   g19434(.A1(new_n19346_), .A2(new_n19690_), .B(new_n19352_), .ZN(new_n19691_));
  AOI21_X1   g19435(.A1(new_n19691_), .A2(new_n19468_), .B(new_n19467_), .ZN(new_n19692_));
  AOI21_X1   g19436(.A1(new_n19692_), .A2(new_n19584_), .B(new_n19581_), .ZN(new_n19693_));
  NOR2_X1    g19437(.A1(new_n19693_), .A2(new_n19689_), .ZN(new_n19694_));
  OAI21_X1   g19438(.A1(new_n19473_), .A2(new_n19585_), .B(new_n19582_), .ZN(new_n19695_));
  NOR2_X1    g19439(.A1(new_n19695_), .A2(new_n19688_), .ZN(new_n19696_));
  NOR2_X1    g19440(.A1(new_n19694_), .A2(new_n19696_), .ZN(new_n19697_));
  XOR2_X1    g19441(.A1(new_n19697_), .A2(new_n19686_), .Z(\f[100] ));
  AOI21_X1   g19442(.A1(new_n19695_), .A2(new_n19688_), .B(new_n19686_), .ZN(new_n19699_));
  NOR2_X1    g19443(.A1(new_n19699_), .A2(new_n19696_), .ZN(new_n19700_));
  OAI21_X1   g19444(.A1(new_n19589_), .A2(new_n19682_), .B(new_n19684_), .ZN(new_n19701_));
  INV_X1     g19445(.I(new_n19701_), .ZN(new_n19702_));
  AOI22_X1   g19446(.A1(new_n13460_), .A2(new_n5166_), .B1(\b[63] ), .B2(new_n5420_), .ZN(new_n19703_));
  AOI22_X1   g19447(.A1(new_n6108_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n6111_), .ZN(new_n19704_));
  OAI21_X1   g19448(.A1(new_n12147_), .A2(new_n7708_), .B(new_n19704_), .ZN(new_n19705_));
  AOI21_X1   g19449(.A1(new_n13444_), .A2(new_n6105_), .B(new_n19705_), .ZN(new_n19706_));
  XOR2_X1    g19450(.A1(new_n19706_), .A2(new_n5849_), .Z(new_n19707_));
  INV_X1     g19451(.I(new_n19707_), .ZN(new_n19708_));
  AOI22_X1   g19452(.A1(new_n7403_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n7408_), .ZN(new_n19709_));
  OAI21_X1   g19453(.A1(new_n9942_), .A2(new_n9488_), .B(new_n19709_), .ZN(new_n19710_));
  AOI21_X1   g19454(.A1(new_n10318_), .A2(new_n7414_), .B(new_n19710_), .ZN(new_n19711_));
  XOR2_X1    g19455(.A1(new_n19711_), .A2(new_n7410_), .Z(new_n19712_));
  INV_X1     g19456(.I(new_n19602_), .ZN(new_n19713_));
  NOR2_X1    g19457(.A1(new_n19647_), .A2(new_n19649_), .ZN(new_n19714_));
  NAND2_X1   g19458(.A1(new_n19647_), .A2(new_n19649_), .ZN(new_n19715_));
  AOI21_X1   g19459(.A1(new_n19713_), .A2(new_n19715_), .B(new_n19714_), .ZN(new_n19716_));
  INV_X1     g19460(.I(new_n19716_), .ZN(new_n19717_));
  OAI22_X1   g19461(.A1(new_n9461_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n9462_), .ZN(new_n19718_));
  AOI21_X1   g19462(.A1(\b[51] ), .A2(new_n8575_), .B(new_n19718_), .ZN(new_n19719_));
  OAI21_X1   g19463(.A1(new_n9385_), .A2(new_n9460_), .B(new_n19719_), .ZN(new_n19720_));
  XOR2_X1    g19464(.A1(new_n19720_), .A2(new_n8248_), .Z(new_n19721_));
  AOI22_X1   g19465(.A1(new_n9125_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n9123_), .ZN(new_n19722_));
  OAI21_X1   g19466(.A1(new_n8127_), .A2(new_n9470_), .B(new_n19722_), .ZN(new_n19723_));
  AOI21_X1   g19467(.A1(new_n9684_), .A2(new_n9129_), .B(new_n19723_), .ZN(new_n19724_));
  XOR2_X1    g19468(.A1(new_n19724_), .A2(new_n9133_), .Z(new_n19725_));
  NAND2_X1   g19469(.A1(new_n19613_), .A2(new_n19615_), .ZN(new_n19726_));
  NOR2_X1    g19470(.A1(new_n19613_), .A2(new_n19615_), .ZN(new_n19727_));
  OAI21_X1   g19471(.A1(new_n19611_), .A2(new_n19727_), .B(new_n19726_), .ZN(new_n19728_));
  AOI22_X1   g19472(.A1(new_n12922_), .A2(\b[38] ), .B1(\b[37] ), .B2(new_n12923_), .ZN(new_n19729_));
  INV_X1     g19473(.I(new_n19729_), .ZN(new_n19730_));
  NOR2_X1    g19474(.A1(new_n19730_), .A2(new_n19614_), .ZN(new_n19731_));
  INV_X1     g19475(.I(new_n19731_), .ZN(new_n19732_));
  NAND2_X1   g19476(.A1(new_n19730_), .A2(new_n19614_), .ZN(new_n19733_));
  NAND2_X1   g19477(.A1(new_n19732_), .A2(new_n19733_), .ZN(new_n19734_));
  XOR2_X1    g19478(.A1(new_n19728_), .A2(new_n19734_), .Z(new_n19735_));
  INV_X1     g19479(.I(new_n19735_), .ZN(new_n19736_));
  AOI22_X1   g19480(.A1(new_n10981_), .A2(\b[44] ), .B1(new_n10979_), .B2(\b[43] ), .ZN(new_n19737_));
  OAI21_X1   g19481(.A1(new_n6490_), .A2(new_n11306_), .B(new_n19737_), .ZN(new_n19738_));
  AOI21_X1   g19482(.A1(new_n7906_), .A2(new_n10984_), .B(new_n19738_), .ZN(new_n19739_));
  XOR2_X1    g19483(.A1(new_n19739_), .A2(new_n10989_), .Z(new_n19740_));
  OAI22_X1   g19484(.A1(new_n13224_), .A2(new_n6285_), .B1(new_n6284_), .B2(new_n11923_), .ZN(new_n19741_));
  AOI21_X1   g19485(.A1(\b[39] ), .A2(new_n13223_), .B(new_n19741_), .ZN(new_n19742_));
  OAI21_X1   g19486(.A1(new_n6299_), .A2(new_n11930_), .B(new_n19742_), .ZN(new_n19743_));
  XOR2_X1    g19487(.A1(new_n19743_), .A2(\a[62] ), .Z(new_n19744_));
  NOR2_X1    g19488(.A1(new_n19740_), .A2(new_n19744_), .ZN(new_n19745_));
  INV_X1     g19489(.I(new_n19745_), .ZN(new_n19746_));
  NAND2_X1   g19490(.A1(new_n19740_), .A2(new_n19744_), .ZN(new_n19747_));
  NAND2_X1   g19491(.A1(new_n19746_), .A2(new_n19747_), .ZN(new_n19748_));
  XOR2_X1    g19492(.A1(new_n19748_), .A2(new_n19736_), .Z(new_n19749_));
  AOI22_X1   g19493(.A1(new_n10064_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n10062_), .ZN(new_n19750_));
  OAI21_X1   g19494(.A1(new_n7096_), .A2(new_n10399_), .B(new_n19750_), .ZN(new_n19751_));
  AOI21_X1   g19495(.A1(new_n7649_), .A2(new_n10068_), .B(new_n19751_), .ZN(new_n19752_));
  XOR2_X1    g19496(.A1(new_n19752_), .A2(new_n10057_), .Z(new_n19753_));
  AOI21_X1   g19497(.A1(new_n19618_), .A2(new_n19627_), .B(new_n19625_), .ZN(new_n19754_));
  NOR2_X1    g19498(.A1(new_n19753_), .A2(new_n19754_), .ZN(new_n19755_));
  NAND2_X1   g19499(.A1(new_n19753_), .A2(new_n19754_), .ZN(new_n19756_));
  INV_X1     g19500(.I(new_n19756_), .ZN(new_n19757_));
  NOR2_X1    g19501(.A1(new_n19757_), .A2(new_n19755_), .ZN(new_n19758_));
  XOR2_X1    g19502(.A1(new_n19758_), .A2(new_n19749_), .Z(new_n19759_));
  AOI21_X1   g19503(.A1(new_n19607_), .A2(new_n19635_), .B(new_n19633_), .ZN(new_n19760_));
  NOR2_X1    g19504(.A1(new_n19759_), .A2(new_n19760_), .ZN(new_n19761_));
  INV_X1     g19505(.I(new_n19761_), .ZN(new_n19762_));
  NAND2_X1   g19506(.A1(new_n19759_), .A2(new_n19760_), .ZN(new_n19763_));
  NAND2_X1   g19507(.A1(new_n19762_), .A2(new_n19763_), .ZN(new_n19764_));
  XOR2_X1    g19508(.A1(new_n19764_), .A2(new_n19725_), .Z(new_n19765_));
  INV_X1     g19509(.I(new_n19765_), .ZN(new_n19766_));
  INV_X1     g19510(.I(new_n19637_), .ZN(new_n19767_));
  AOI21_X1   g19511(.A1(new_n19767_), .A2(new_n19644_), .B(new_n19643_), .ZN(new_n19768_));
  NOR2_X1    g19512(.A1(new_n19766_), .A2(new_n19768_), .ZN(new_n19769_));
  INV_X1     g19513(.I(new_n19769_), .ZN(new_n19770_));
  NAND2_X1   g19514(.A1(new_n19766_), .A2(new_n19768_), .ZN(new_n19771_));
  NAND2_X1   g19515(.A1(new_n19770_), .A2(new_n19771_), .ZN(new_n19772_));
  XNOR2_X1   g19516(.A1(new_n19772_), .A2(new_n19721_), .ZN(new_n19773_));
  NOR2_X1    g19517(.A1(new_n19773_), .A2(new_n19717_), .ZN(new_n19774_));
  INV_X1     g19518(.I(new_n19774_), .ZN(new_n19775_));
  NAND2_X1   g19519(.A1(new_n19773_), .A2(new_n19717_), .ZN(new_n19776_));
  NAND2_X1   g19520(.A1(new_n19775_), .A2(new_n19776_), .ZN(new_n19777_));
  XNOR2_X1   g19521(.A1(new_n19777_), .A2(new_n19712_), .ZN(new_n19778_));
  OAI22_X1   g19522(.A1(new_n7730_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n7731_), .ZN(new_n19779_));
  AOI21_X1   g19523(.A1(\b[57] ), .A2(new_n6887_), .B(new_n19779_), .ZN(new_n19780_));
  OAI21_X1   g19524(.A1(new_n12203_), .A2(new_n7728_), .B(new_n19780_), .ZN(new_n19781_));
  XOR2_X1    g19525(.A1(new_n19781_), .A2(\a[44] ), .Z(new_n19782_));
  AOI21_X1   g19526(.A1(new_n19652_), .A2(new_n19661_), .B(new_n19659_), .ZN(new_n19783_));
  NOR2_X1    g19527(.A1(new_n19783_), .A2(new_n19782_), .ZN(new_n19784_));
  AND2_X2    g19528(.A1(new_n19783_), .A2(new_n19782_), .Z(new_n19785_));
  NOR2_X1    g19529(.A1(new_n19785_), .A2(new_n19784_), .ZN(new_n19786_));
  XOR2_X1    g19530(.A1(new_n19778_), .A2(new_n19786_), .Z(new_n19787_));
  AOI21_X1   g19531(.A1(new_n19598_), .A2(new_n19668_), .B(new_n19666_), .ZN(new_n19788_));
  NOR2_X1    g19532(.A1(new_n19787_), .A2(new_n19788_), .ZN(new_n19789_));
  INV_X1     g19533(.I(new_n19789_), .ZN(new_n19790_));
  NAND2_X1   g19534(.A1(new_n19787_), .A2(new_n19788_), .ZN(new_n19791_));
  NAND2_X1   g19535(.A1(new_n19790_), .A2(new_n19791_), .ZN(new_n19792_));
  XOR2_X1    g19536(.A1(new_n19792_), .A2(new_n19708_), .Z(new_n19793_));
  XOR2_X1    g19537(.A1(new_n19793_), .A2(new_n19703_), .Z(new_n19794_));
  INV_X1     g19538(.I(new_n19670_), .ZN(new_n19795_));
  NAND2_X1   g19539(.A1(new_n19679_), .A2(new_n19795_), .ZN(new_n19796_));
  NAND2_X1   g19540(.A1(new_n19796_), .A2(new_n19678_), .ZN(new_n19797_));
  XOR2_X1    g19541(.A1(new_n19797_), .A2(\a[38] ), .Z(new_n19798_));
  XOR2_X1    g19542(.A1(new_n19794_), .A2(new_n19798_), .Z(new_n19799_));
  NOR2_X1    g19543(.A1(new_n19799_), .A2(new_n19702_), .ZN(new_n19800_));
  NAND2_X1   g19544(.A1(new_n19799_), .A2(new_n19702_), .ZN(new_n19801_));
  INV_X1     g19545(.I(new_n19801_), .ZN(new_n19802_));
  NOR2_X1    g19546(.A1(new_n19802_), .A2(new_n19800_), .ZN(new_n19803_));
  XOR2_X1    g19547(.A1(new_n19700_), .A2(new_n19803_), .Z(\f[101] ));
  NAND2_X1   g19548(.A1(new_n19693_), .A2(new_n19689_), .ZN(new_n19805_));
  INV_X1     g19549(.I(new_n19686_), .ZN(new_n19806_));
  OAI21_X1   g19550(.A1(new_n19693_), .A2(new_n19689_), .B(new_n19806_), .ZN(new_n19807_));
  AOI21_X1   g19551(.A1(new_n19807_), .A2(new_n19805_), .B(new_n19802_), .ZN(new_n19808_));
  AOI22_X1   g19552(.A1(new_n6108_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n6111_), .ZN(new_n19809_));
  OAI21_X1   g19553(.A1(new_n12148_), .A2(new_n7708_), .B(new_n19809_), .ZN(new_n19810_));
  AOI21_X1   g19554(.A1(new_n12811_), .A2(new_n6105_), .B(new_n19810_), .ZN(new_n19811_));
  XOR2_X1    g19555(.A1(new_n19811_), .A2(new_n5849_), .Z(new_n19812_));
  AOI21_X1   g19556(.A1(new_n19708_), .A2(new_n19791_), .B(new_n19789_), .ZN(new_n19813_));
  OAI21_X1   g19557(.A1(new_n19712_), .A2(new_n19774_), .B(new_n19776_), .ZN(new_n19814_));
  AOI21_X1   g19558(.A1(new_n19721_), .A2(new_n19771_), .B(new_n19769_), .ZN(new_n19815_));
  AOI22_X1   g19559(.A1(new_n8241_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n8246_), .ZN(new_n19816_));
  OAI21_X1   g19560(.A1(new_n9032_), .A2(new_n9114_), .B(new_n19816_), .ZN(new_n19817_));
  AOI21_X1   g19561(.A1(new_n10884_), .A2(new_n8252_), .B(new_n19817_), .ZN(new_n19818_));
  XOR2_X1    g19562(.A1(new_n19818_), .A2(new_n8248_), .Z(new_n19819_));
  INV_X1     g19563(.I(new_n19819_), .ZN(new_n19820_));
  INV_X1     g19564(.I(new_n19725_), .ZN(new_n19821_));
  AOI21_X1   g19565(.A1(new_n19821_), .A2(new_n19763_), .B(new_n19761_), .ZN(new_n19822_));
  AOI21_X1   g19566(.A1(new_n19728_), .A2(new_n19733_), .B(new_n19731_), .ZN(new_n19823_));
  AOI22_X1   g19567(.A1(new_n11926_), .A2(\b[42] ), .B1(new_n11924_), .B2(\b[41] ), .ZN(new_n19824_));
  OAI21_X1   g19568(.A1(new_n6284_), .A2(new_n12317_), .B(new_n19824_), .ZN(new_n19825_));
  AOI21_X1   g19569(.A1(new_n7106_), .A2(new_n11929_), .B(new_n19825_), .ZN(new_n19826_));
  XOR2_X1    g19570(.A1(new_n19826_), .A2(new_n12312_), .Z(new_n19827_));
  INV_X1     g19571(.I(new_n19827_), .ZN(new_n19828_));
  AOI22_X1   g19572(.A1(new_n12922_), .A2(\b[39] ), .B1(\b[38] ), .B2(new_n12923_), .ZN(new_n19829_));
  INV_X1     g19573(.I(new_n19829_), .ZN(new_n19830_));
  NOR2_X1    g19574(.A1(new_n19830_), .A2(new_n5162_), .ZN(new_n19831_));
  NOR2_X1    g19575(.A1(new_n19829_), .A2(\a[38] ), .ZN(new_n19832_));
  NOR2_X1    g19576(.A1(new_n19831_), .A2(new_n19832_), .ZN(new_n19833_));
  XOR2_X1    g19577(.A1(new_n19833_), .A2(new_n19614_), .Z(new_n19834_));
  NOR2_X1    g19578(.A1(new_n19828_), .A2(new_n19834_), .ZN(new_n19835_));
  NAND2_X1   g19579(.A1(new_n19828_), .A2(new_n19834_), .ZN(new_n19836_));
  INV_X1     g19580(.I(new_n19836_), .ZN(new_n19837_));
  NOR2_X1    g19581(.A1(new_n19837_), .A2(new_n19835_), .ZN(new_n19838_));
  XOR2_X1    g19582(.A1(new_n19838_), .A2(new_n19823_), .Z(new_n19839_));
  NAND2_X1   g19583(.A1(new_n19747_), .A2(new_n19736_), .ZN(new_n19840_));
  NAND2_X1   g19584(.A1(new_n19840_), .A2(new_n19746_), .ZN(new_n19841_));
  INV_X1     g19585(.I(new_n19841_), .ZN(new_n19842_));
  AOI22_X1   g19586(.A1(new_n10981_), .A2(\b[45] ), .B1(new_n10979_), .B2(\b[44] ), .ZN(new_n19843_));
  OAI21_X1   g19587(.A1(new_n6775_), .A2(new_n11306_), .B(new_n19843_), .ZN(new_n19844_));
  AOI21_X1   g19588(.A1(new_n7926_), .A2(new_n10984_), .B(new_n19844_), .ZN(new_n19845_));
  XOR2_X1    g19589(.A1(new_n19845_), .A2(new_n10989_), .Z(new_n19846_));
  NOR2_X1    g19590(.A1(new_n19842_), .A2(new_n19846_), .ZN(new_n19847_));
  INV_X1     g19591(.I(new_n19847_), .ZN(new_n19848_));
  NAND2_X1   g19592(.A1(new_n19842_), .A2(new_n19846_), .ZN(new_n19849_));
  NAND2_X1   g19593(.A1(new_n19848_), .A2(new_n19849_), .ZN(new_n19850_));
  XOR2_X1    g19594(.A1(new_n19850_), .A2(new_n19839_), .Z(new_n19851_));
  AOI22_X1   g19595(.A1(new_n10064_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n10062_), .ZN(new_n19852_));
  OAI21_X1   g19596(.A1(new_n7617_), .A2(new_n10399_), .B(new_n19852_), .ZN(new_n19853_));
  AOI21_X1   g19597(.A1(new_n8792_), .A2(new_n10068_), .B(new_n19853_), .ZN(new_n19854_));
  XOR2_X1    g19598(.A1(new_n19854_), .A2(\a[56] ), .Z(new_n19855_));
  INV_X1     g19599(.I(new_n19755_), .ZN(new_n19856_));
  OAI21_X1   g19600(.A1(new_n19749_), .A2(new_n19757_), .B(new_n19856_), .ZN(new_n19857_));
  NAND2_X1   g19601(.A1(new_n19857_), .A2(new_n19855_), .ZN(new_n19858_));
  OR2_X2     g19602(.A1(new_n19857_), .A2(new_n19855_), .Z(new_n19859_));
  NAND2_X1   g19603(.A1(new_n19859_), .A2(new_n19858_), .ZN(new_n19860_));
  XNOR2_X1   g19604(.A1(new_n19860_), .A2(new_n19851_), .ZN(new_n19861_));
  INV_X1     g19605(.I(new_n19861_), .ZN(new_n19862_));
  AOI22_X1   g19606(.A1(new_n9125_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n9123_), .ZN(new_n19863_));
  OAI21_X1   g19607(.A1(new_n8168_), .A2(new_n9470_), .B(new_n19863_), .ZN(new_n19864_));
  AOI21_X1   g19608(.A1(new_n8783_), .A2(new_n9129_), .B(new_n19864_), .ZN(new_n19865_));
  XOR2_X1    g19609(.A1(new_n19865_), .A2(new_n9133_), .Z(new_n19866_));
  NOR2_X1    g19610(.A1(new_n19862_), .A2(new_n19866_), .ZN(new_n19867_));
  INV_X1     g19611(.I(new_n19867_), .ZN(new_n19868_));
  NAND2_X1   g19612(.A1(new_n19862_), .A2(new_n19866_), .ZN(new_n19869_));
  NAND2_X1   g19613(.A1(new_n19868_), .A2(new_n19869_), .ZN(new_n19870_));
  XOR2_X1    g19614(.A1(new_n19870_), .A2(new_n19822_), .Z(new_n19871_));
  NOR2_X1    g19615(.A1(new_n19871_), .A2(new_n19820_), .ZN(new_n19872_));
  INV_X1     g19616(.I(new_n19872_), .ZN(new_n19873_));
  NAND2_X1   g19617(.A1(new_n19871_), .A2(new_n19820_), .ZN(new_n19874_));
  NAND2_X1   g19618(.A1(new_n19873_), .A2(new_n19874_), .ZN(new_n19875_));
  XOR2_X1    g19619(.A1(new_n19875_), .A2(new_n19815_), .Z(new_n19876_));
  AOI22_X1   g19620(.A1(new_n7403_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n7408_), .ZN(new_n19877_));
  OAI21_X1   g19621(.A1(new_n9972_), .A2(new_n9488_), .B(new_n19877_), .ZN(new_n19878_));
  AOI21_X1   g19622(.A1(new_n10631_), .A2(new_n7414_), .B(new_n19878_), .ZN(new_n19879_));
  XOR2_X1    g19623(.A1(new_n19879_), .A2(\a[47] ), .Z(new_n19880_));
  NAND2_X1   g19624(.A1(new_n19876_), .A2(new_n19880_), .ZN(new_n19881_));
  OR2_X2     g19625(.A1(new_n19876_), .A2(new_n19880_), .Z(new_n19882_));
  NAND2_X1   g19626(.A1(new_n19882_), .A2(new_n19881_), .ZN(new_n19883_));
  XNOR2_X1   g19627(.A1(new_n19883_), .A2(new_n19814_), .ZN(new_n19884_));
  AOI22_X1   g19628(.A1(new_n6569_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n6574_), .ZN(new_n19885_));
  OAI21_X1   g19629(.A1(new_n11195_), .A2(new_n8565_), .B(new_n19885_), .ZN(new_n19886_));
  AOI21_X1   g19630(.A1(new_n11836_), .A2(new_n6579_), .B(new_n19886_), .ZN(new_n19887_));
  XOR2_X1    g19631(.A1(new_n19887_), .A2(\a[44] ), .Z(new_n19888_));
  INV_X1     g19632(.I(new_n19784_), .ZN(new_n19889_));
  OAI21_X1   g19633(.A1(new_n19778_), .A2(new_n19785_), .B(new_n19889_), .ZN(new_n19890_));
  NAND2_X1   g19634(.A1(new_n19890_), .A2(new_n19888_), .ZN(new_n19891_));
  OR2_X2     g19635(.A1(new_n19890_), .A2(new_n19888_), .Z(new_n19892_));
  NAND2_X1   g19636(.A1(new_n19892_), .A2(new_n19891_), .ZN(new_n19893_));
  XOR2_X1    g19637(.A1(new_n19893_), .A2(new_n19884_), .Z(new_n19894_));
  NAND2_X1   g19638(.A1(new_n19894_), .A2(new_n19813_), .ZN(new_n19895_));
  NOR2_X1    g19639(.A1(new_n19894_), .A2(new_n19813_), .ZN(new_n19896_));
  INV_X1     g19640(.I(new_n19896_), .ZN(new_n19897_));
  NAND2_X1   g19641(.A1(new_n19897_), .A2(new_n19895_), .ZN(new_n19898_));
  XOR2_X1    g19642(.A1(new_n19898_), .A2(new_n19812_), .Z(new_n19899_));
  INV_X1     g19643(.I(new_n19793_), .ZN(new_n19900_));
  INV_X1     g19644(.I(new_n19797_), .ZN(new_n19901_));
  XOR2_X1    g19645(.A1(new_n19703_), .A2(new_n5162_), .Z(new_n19902_));
  AOI21_X1   g19646(.A1(new_n19793_), .A2(new_n19901_), .B(new_n19902_), .ZN(new_n19903_));
  AOI21_X1   g19647(.A1(new_n19900_), .A2(new_n19797_), .B(new_n19903_), .ZN(new_n19904_));
  INV_X1     g19648(.I(new_n19904_), .ZN(new_n19905_));
  NOR2_X1    g19649(.A1(new_n19899_), .A2(new_n19905_), .ZN(new_n19906_));
  INV_X1     g19650(.I(new_n19906_), .ZN(new_n19907_));
  NAND2_X1   g19651(.A1(new_n19899_), .A2(new_n19905_), .ZN(new_n19908_));
  AND2_X2    g19652(.A1(new_n19907_), .A2(new_n19908_), .Z(new_n19909_));
  INV_X1     g19653(.I(new_n19909_), .ZN(new_n19910_));
  NOR3_X1    g19654(.A1(new_n19808_), .A2(new_n19800_), .A3(new_n19910_), .ZN(new_n19911_));
  INV_X1     g19655(.I(new_n19800_), .ZN(new_n19912_));
  OAI21_X1   g19656(.A1(new_n19699_), .A2(new_n19696_), .B(new_n19801_), .ZN(new_n19913_));
  AOI21_X1   g19657(.A1(new_n19913_), .A2(new_n19912_), .B(new_n19909_), .ZN(new_n19914_));
  NOR2_X1    g19658(.A1(new_n19911_), .A2(new_n19914_), .ZN(\f[102] ));
  OAI22_X1   g19659(.A1(new_n7708_), .A2(new_n12796_), .B1(new_n12800_), .B2(new_n5857_), .ZN(new_n19916_));
  AOI21_X1   g19660(.A1(new_n13973_), .A2(new_n6105_), .B(new_n19916_), .ZN(new_n19917_));
  XOR2_X1    g19661(.A1(new_n19917_), .A2(new_n5849_), .Z(new_n19918_));
  INV_X1     g19662(.I(new_n19918_), .ZN(new_n19919_));
  INV_X1     g19663(.I(new_n19891_), .ZN(new_n19920_));
  AOI21_X1   g19664(.A1(new_n19884_), .A2(new_n19892_), .B(new_n19920_), .ZN(new_n19921_));
  INV_X1     g19665(.I(new_n19921_), .ZN(new_n19922_));
  AOI22_X1   g19666(.A1(new_n7403_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n7408_), .ZN(new_n19923_));
  OAI21_X1   g19667(.A1(new_n10308_), .A2(new_n9488_), .B(new_n19923_), .ZN(new_n19924_));
  AOI21_X1   g19668(.A1(new_n12164_), .A2(new_n7414_), .B(new_n19924_), .ZN(new_n19925_));
  XOR2_X1    g19669(.A1(new_n19925_), .A2(new_n7410_), .Z(new_n19926_));
  INV_X1     g19670(.I(new_n19926_), .ZN(new_n19927_));
  AOI22_X1   g19671(.A1(new_n9125_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n9123_), .ZN(new_n19928_));
  OAI21_X1   g19672(.A1(new_n8500_), .A2(new_n9470_), .B(new_n19928_), .ZN(new_n19929_));
  AOI21_X1   g19673(.A1(new_n9987_), .A2(new_n9129_), .B(new_n19929_), .ZN(new_n19930_));
  XOR2_X1    g19674(.A1(new_n19930_), .A2(new_n9133_), .Z(new_n19931_));
  OAI21_X1   g19675(.A1(new_n19823_), .A2(new_n19835_), .B(new_n19836_), .ZN(new_n19932_));
  INV_X1     g19676(.I(new_n19932_), .ZN(new_n19933_));
  AOI22_X1   g19677(.A1(new_n10981_), .A2(\b[46] ), .B1(new_n10979_), .B2(\b[45] ), .ZN(new_n19934_));
  OAI21_X1   g19678(.A1(new_n7074_), .A2(new_n11306_), .B(new_n19934_), .ZN(new_n19935_));
  AOI21_X1   g19679(.A1(new_n9337_), .A2(new_n10984_), .B(new_n19935_), .ZN(new_n19936_));
  XOR2_X1    g19680(.A1(new_n19936_), .A2(new_n10989_), .Z(new_n19937_));
  INV_X1     g19681(.I(new_n19937_), .ZN(new_n19938_));
  OAI22_X1   g19682(.A1(new_n13224_), .A2(new_n6775_), .B1(new_n6490_), .B2(new_n11923_), .ZN(new_n19939_));
  AOI21_X1   g19683(.A1(\b[41] ), .A2(new_n13223_), .B(new_n19939_), .ZN(new_n19940_));
  OAI21_X1   g19684(.A1(new_n6785_), .A2(new_n11930_), .B(new_n19940_), .ZN(new_n19941_));
  XOR2_X1    g19685(.A1(new_n19941_), .A2(\a[62] ), .Z(new_n19942_));
  INV_X1     g19686(.I(new_n19832_), .ZN(new_n19943_));
  AOI21_X1   g19687(.A1(new_n19614_), .A2(new_n19943_), .B(new_n19831_), .ZN(new_n19944_));
  AOI22_X1   g19688(.A1(new_n12922_), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n12923_), .ZN(new_n19945_));
  AND2_X2    g19689(.A1(new_n19944_), .A2(new_n19945_), .Z(new_n19946_));
  NOR2_X1    g19690(.A1(new_n19944_), .A2(new_n19945_), .ZN(new_n19947_));
  NOR2_X1    g19691(.A1(new_n19946_), .A2(new_n19947_), .ZN(new_n19948_));
  XNOR2_X1   g19692(.A1(new_n19942_), .A2(new_n19948_), .ZN(new_n19949_));
  NOR2_X1    g19693(.A1(new_n19938_), .A2(new_n19949_), .ZN(new_n19950_));
  NAND2_X1   g19694(.A1(new_n19938_), .A2(new_n19949_), .ZN(new_n19951_));
  INV_X1     g19695(.I(new_n19951_), .ZN(new_n19952_));
  NOR2_X1    g19696(.A1(new_n19952_), .A2(new_n19950_), .ZN(new_n19953_));
  XOR2_X1    g19697(.A1(new_n19953_), .A2(new_n19933_), .Z(new_n19954_));
  INV_X1     g19698(.I(new_n19839_), .ZN(new_n19955_));
  AOI21_X1   g19699(.A1(new_n19955_), .A2(new_n19849_), .B(new_n19847_), .ZN(new_n19956_));
  OAI22_X1   g19700(.A1(new_n11298_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n11297_), .ZN(new_n19957_));
  AOI21_X1   g19701(.A1(\b[47] ), .A2(new_n11296_), .B(new_n19957_), .ZN(new_n19958_));
  OAI21_X1   g19702(.A1(new_n9050_), .A2(new_n10069_), .B(new_n19958_), .ZN(new_n19959_));
  XOR2_X1    g19703(.A1(new_n19959_), .A2(\a[56] ), .Z(new_n19960_));
  NOR2_X1    g19704(.A1(new_n19960_), .A2(new_n19956_), .ZN(new_n19961_));
  NAND2_X1   g19705(.A1(new_n19960_), .A2(new_n19956_), .ZN(new_n19962_));
  INV_X1     g19706(.I(new_n19962_), .ZN(new_n19963_));
  NOR2_X1    g19707(.A1(new_n19963_), .A2(new_n19961_), .ZN(new_n19964_));
  XOR2_X1    g19708(.A1(new_n19964_), .A2(new_n19954_), .Z(new_n19965_));
  INV_X1     g19709(.I(new_n19858_), .ZN(new_n19966_));
  AOI21_X1   g19710(.A1(new_n19851_), .A2(new_n19859_), .B(new_n19966_), .ZN(new_n19967_));
  XOR2_X1    g19711(.A1(new_n19965_), .A2(new_n19967_), .Z(new_n19968_));
  XOR2_X1    g19712(.A1(new_n19968_), .A2(new_n19931_), .Z(new_n19969_));
  INV_X1     g19713(.I(new_n19969_), .ZN(new_n19970_));
  INV_X1     g19714(.I(new_n19822_), .ZN(new_n19971_));
  AOI21_X1   g19715(.A1(new_n19971_), .A2(new_n19869_), .B(new_n19867_), .ZN(new_n19972_));
  AOI22_X1   g19716(.A1(new_n8241_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n8246_), .ZN(new_n19973_));
  OAI21_X1   g19717(.A1(new_n9376_), .A2(new_n9114_), .B(new_n19973_), .ZN(new_n19974_));
  AOI21_X1   g19718(.A1(new_n9979_), .A2(new_n8252_), .B(new_n19974_), .ZN(new_n19975_));
  XOR2_X1    g19719(.A1(new_n19975_), .A2(new_n8248_), .Z(new_n19976_));
  NOR2_X1    g19720(.A1(new_n19972_), .A2(new_n19976_), .ZN(new_n19977_));
  INV_X1     g19721(.I(new_n19977_), .ZN(new_n19978_));
  NAND2_X1   g19722(.A1(new_n19972_), .A2(new_n19976_), .ZN(new_n19979_));
  NAND2_X1   g19723(.A1(new_n19978_), .A2(new_n19979_), .ZN(new_n19980_));
  XOR2_X1    g19724(.A1(new_n19980_), .A2(new_n19970_), .Z(new_n19981_));
  OAI21_X1   g19725(.A1(new_n19815_), .A2(new_n19872_), .B(new_n19874_), .ZN(new_n19982_));
  INV_X1     g19726(.I(new_n19982_), .ZN(new_n19983_));
  NOR2_X1    g19727(.A1(new_n19983_), .A2(new_n19981_), .ZN(new_n19984_));
  INV_X1     g19728(.I(new_n19984_), .ZN(new_n19985_));
  NAND2_X1   g19729(.A1(new_n19983_), .A2(new_n19981_), .ZN(new_n19986_));
  NAND2_X1   g19730(.A1(new_n19985_), .A2(new_n19986_), .ZN(new_n19987_));
  XOR2_X1    g19731(.A1(new_n19987_), .A2(new_n19927_), .Z(new_n19988_));
  INV_X1     g19732(.I(new_n19881_), .ZN(new_n19989_));
  AOI21_X1   g19733(.A1(new_n19814_), .A2(new_n19882_), .B(new_n19989_), .ZN(new_n19990_));
  OAI22_X1   g19734(.A1(new_n7730_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n7731_), .ZN(new_n19991_));
  AOI21_X1   g19735(.A1(\b[59] ), .A2(new_n6887_), .B(new_n19991_), .ZN(new_n19992_));
  OAI21_X1   g19736(.A1(new_n13110_), .A2(new_n7728_), .B(new_n19992_), .ZN(new_n19993_));
  XOR2_X1    g19737(.A1(new_n19993_), .A2(\a[44] ), .Z(new_n19994_));
  NOR2_X1    g19738(.A1(new_n19990_), .A2(new_n19994_), .ZN(new_n19995_));
  INV_X1     g19739(.I(new_n19995_), .ZN(new_n19996_));
  NAND2_X1   g19740(.A1(new_n19990_), .A2(new_n19994_), .ZN(new_n19997_));
  NAND2_X1   g19741(.A1(new_n19996_), .A2(new_n19997_), .ZN(new_n19998_));
  XOR2_X1    g19742(.A1(new_n19998_), .A2(new_n19988_), .Z(new_n19999_));
  NOR2_X1    g19743(.A1(new_n19999_), .A2(new_n19922_), .ZN(new_n20000_));
  INV_X1     g19744(.I(new_n20000_), .ZN(new_n20001_));
  NAND2_X1   g19745(.A1(new_n19999_), .A2(new_n19922_), .ZN(new_n20002_));
  NAND2_X1   g19746(.A1(new_n20001_), .A2(new_n20002_), .ZN(new_n20003_));
  XOR2_X1    g19747(.A1(new_n20003_), .A2(new_n19919_), .Z(new_n20004_));
  INV_X1     g19748(.I(new_n20004_), .ZN(new_n20005_));
  INV_X1     g19749(.I(new_n19812_), .ZN(new_n20006_));
  AOI21_X1   g19750(.A1(new_n20006_), .A2(new_n19895_), .B(new_n19896_), .ZN(new_n20007_));
  OAI21_X1   g19751(.A1(new_n19911_), .A2(new_n19906_), .B(new_n20007_), .ZN(new_n20008_));
  NAND3_X1   g19752(.A1(new_n19913_), .A2(new_n19912_), .A3(new_n19909_), .ZN(new_n20009_));
  INV_X1     g19753(.I(new_n20007_), .ZN(new_n20010_));
  NAND3_X1   g19754(.A1(new_n20009_), .A2(new_n19907_), .A3(new_n20010_), .ZN(new_n20011_));
  NAND2_X1   g19755(.A1(new_n20008_), .A2(new_n20011_), .ZN(new_n20012_));
  XOR2_X1    g19756(.A1(new_n20012_), .A2(new_n20005_), .Z(\f[103] ));
  AOI21_X1   g19757(.A1(new_n20009_), .A2(new_n19907_), .B(new_n20010_), .ZN(new_n20014_));
  OAI21_X1   g19758(.A1(new_n20004_), .A2(new_n20014_), .B(new_n20011_), .ZN(new_n20015_));
  OAI21_X1   g19759(.A1(new_n19918_), .A2(new_n20000_), .B(new_n20002_), .ZN(new_n20016_));
  INV_X1     g19760(.I(new_n20016_), .ZN(new_n20017_));
  AOI22_X1   g19761(.A1(new_n13460_), .A2(new_n6105_), .B1(\b[63] ), .B2(new_n6115_), .ZN(new_n20018_));
  AOI22_X1   g19762(.A1(new_n6569_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n6574_), .ZN(new_n20019_));
  OAI21_X1   g19763(.A1(new_n12147_), .A2(new_n8565_), .B(new_n20019_), .ZN(new_n20020_));
  AOI21_X1   g19764(.A1(new_n13444_), .A2(new_n6579_), .B(new_n20020_), .ZN(new_n20021_));
  XOR2_X1    g19765(.A1(new_n20021_), .A2(new_n6567_), .Z(new_n20022_));
  INV_X1     g19766(.I(new_n20022_), .ZN(new_n20023_));
  AOI22_X1   g19767(.A1(new_n8241_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n8246_), .ZN(new_n20024_));
  OAI21_X1   g19768(.A1(new_n9942_), .A2(new_n9114_), .B(new_n20024_), .ZN(new_n20025_));
  AOI21_X1   g19769(.A1(new_n10318_), .A2(new_n8252_), .B(new_n20025_), .ZN(new_n20026_));
  XOR2_X1    g19770(.A1(new_n20026_), .A2(new_n8248_), .Z(new_n20027_));
  INV_X1     g19771(.I(new_n19931_), .ZN(new_n20028_));
  NOR2_X1    g19772(.A1(new_n19965_), .A2(new_n19967_), .ZN(new_n20029_));
  NAND2_X1   g19773(.A1(new_n19965_), .A2(new_n19967_), .ZN(new_n20030_));
  AOI21_X1   g19774(.A1(new_n20028_), .A2(new_n20030_), .B(new_n20029_), .ZN(new_n20031_));
  INV_X1     g19775(.I(new_n20031_), .ZN(new_n20032_));
  OAI22_X1   g19776(.A1(new_n10390_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n10389_), .ZN(new_n20033_));
  AOI21_X1   g19777(.A1(\b[51] ), .A2(new_n9471_), .B(new_n20033_), .ZN(new_n20034_));
  OAI21_X1   g19778(.A1(new_n9385_), .A2(new_n10388_), .B(new_n20034_), .ZN(new_n20035_));
  XOR2_X1    g19779(.A1(new_n20035_), .A2(new_n9133_), .Z(new_n20036_));
  AOI22_X1   g19780(.A1(new_n10064_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n10062_), .ZN(new_n20037_));
  OAI21_X1   g19781(.A1(new_n8127_), .A2(new_n10399_), .B(new_n20037_), .ZN(new_n20038_));
  AOI21_X1   g19782(.A1(new_n9684_), .A2(new_n10068_), .B(new_n20038_), .ZN(new_n20039_));
  XOR2_X1    g19783(.A1(new_n20039_), .A2(new_n10057_), .Z(new_n20040_));
  OAI21_X1   g19784(.A1(new_n19933_), .A2(new_n19950_), .B(new_n19951_), .ZN(new_n20041_));
  AOI22_X1   g19785(.A1(new_n10981_), .A2(\b[47] ), .B1(new_n10979_), .B2(\b[46] ), .ZN(new_n20042_));
  OAI21_X1   g19786(.A1(new_n7096_), .A2(new_n11306_), .B(new_n20042_), .ZN(new_n20043_));
  AOI21_X1   g19787(.A1(new_n7649_), .A2(new_n10984_), .B(new_n20043_), .ZN(new_n20044_));
  XOR2_X1    g19788(.A1(new_n20044_), .A2(new_n10989_), .Z(new_n20045_));
  AOI22_X1   g19789(.A1(new_n11926_), .A2(\b[44] ), .B1(new_n11924_), .B2(\b[43] ), .ZN(new_n20046_));
  OAI21_X1   g19790(.A1(new_n6490_), .A2(new_n12317_), .B(new_n20046_), .ZN(new_n20047_));
  AOI21_X1   g19791(.A1(new_n7906_), .A2(new_n11929_), .B(new_n20047_), .ZN(new_n20048_));
  XOR2_X1    g19792(.A1(new_n20048_), .A2(new_n12312_), .Z(new_n20049_));
  NOR2_X1    g19793(.A1(new_n20045_), .A2(new_n20049_), .ZN(new_n20050_));
  INV_X1     g19794(.I(new_n20050_), .ZN(new_n20051_));
  NAND2_X1   g19795(.A1(new_n20045_), .A2(new_n20049_), .ZN(new_n20052_));
  NAND2_X1   g19796(.A1(new_n20051_), .A2(new_n20052_), .ZN(new_n20053_));
  INV_X1     g19797(.I(new_n19947_), .ZN(new_n20054_));
  OAI21_X1   g19798(.A1(new_n19942_), .A2(new_n19946_), .B(new_n20054_), .ZN(new_n20055_));
  AOI22_X1   g19799(.A1(new_n12922_), .A2(\b[41] ), .B1(\b[40] ), .B2(new_n12923_), .ZN(new_n20056_));
  INV_X1     g19800(.I(new_n20056_), .ZN(new_n20057_));
  NOR2_X1    g19801(.A1(new_n20057_), .A2(new_n19945_), .ZN(new_n20058_));
  INV_X1     g19802(.I(new_n20058_), .ZN(new_n20059_));
  NAND2_X1   g19803(.A1(new_n20057_), .A2(new_n19945_), .ZN(new_n20060_));
  NAND2_X1   g19804(.A1(new_n20059_), .A2(new_n20060_), .ZN(new_n20061_));
  XOR2_X1    g19805(.A1(new_n20055_), .A2(new_n20061_), .Z(new_n20062_));
  XOR2_X1    g19806(.A1(new_n20053_), .A2(new_n20062_), .Z(new_n20063_));
  NOR2_X1    g19807(.A1(new_n20063_), .A2(new_n20041_), .ZN(new_n20064_));
  INV_X1     g19808(.I(new_n20064_), .ZN(new_n20065_));
  NAND2_X1   g19809(.A1(new_n20063_), .A2(new_n20041_), .ZN(new_n20066_));
  NAND2_X1   g19810(.A1(new_n20065_), .A2(new_n20066_), .ZN(new_n20067_));
  XOR2_X1    g19811(.A1(new_n20067_), .A2(new_n20040_), .Z(new_n20068_));
  INV_X1     g19812(.I(new_n20068_), .ZN(new_n20069_));
  INV_X1     g19813(.I(new_n19954_), .ZN(new_n20070_));
  AOI21_X1   g19814(.A1(new_n20070_), .A2(new_n19962_), .B(new_n19961_), .ZN(new_n20071_));
  NOR2_X1    g19815(.A1(new_n20069_), .A2(new_n20071_), .ZN(new_n20072_));
  INV_X1     g19816(.I(new_n20072_), .ZN(new_n20073_));
  NAND2_X1   g19817(.A1(new_n20069_), .A2(new_n20071_), .ZN(new_n20074_));
  NAND2_X1   g19818(.A1(new_n20073_), .A2(new_n20074_), .ZN(new_n20075_));
  XNOR2_X1   g19819(.A1(new_n20075_), .A2(new_n20036_), .ZN(new_n20076_));
  NOR2_X1    g19820(.A1(new_n20076_), .A2(new_n20032_), .ZN(new_n20077_));
  INV_X1     g19821(.I(new_n20077_), .ZN(new_n20078_));
  NAND2_X1   g19822(.A1(new_n20076_), .A2(new_n20032_), .ZN(new_n20079_));
  NAND2_X1   g19823(.A1(new_n20078_), .A2(new_n20079_), .ZN(new_n20080_));
  XOR2_X1    g19824(.A1(new_n20080_), .A2(new_n20027_), .Z(new_n20081_));
  OAI22_X1   g19825(.A1(new_n11195_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n12151_), .ZN(new_n20082_));
  AOI21_X1   g19826(.A1(\b[57] ), .A2(new_n7719_), .B(new_n20082_), .ZN(new_n20083_));
  OAI21_X1   g19827(.A1(new_n12203_), .A2(new_n8585_), .B(new_n20083_), .ZN(new_n20084_));
  XOR2_X1    g19828(.A1(new_n20084_), .A2(\a[47] ), .Z(new_n20085_));
  AOI21_X1   g19829(.A1(new_n19970_), .A2(new_n19979_), .B(new_n19977_), .ZN(new_n20086_));
  NOR2_X1    g19830(.A1(new_n20086_), .A2(new_n20085_), .ZN(new_n20087_));
  INV_X1     g19831(.I(new_n20087_), .ZN(new_n20088_));
  NAND2_X1   g19832(.A1(new_n20086_), .A2(new_n20085_), .ZN(new_n20089_));
  NAND2_X1   g19833(.A1(new_n20088_), .A2(new_n20089_), .ZN(new_n20090_));
  XOR2_X1    g19834(.A1(new_n20081_), .A2(new_n20090_), .Z(new_n20091_));
  AOI21_X1   g19835(.A1(new_n19927_), .A2(new_n19986_), .B(new_n19984_), .ZN(new_n20092_));
  NOR2_X1    g19836(.A1(new_n20091_), .A2(new_n20092_), .ZN(new_n20093_));
  INV_X1     g19837(.I(new_n20093_), .ZN(new_n20094_));
  NAND2_X1   g19838(.A1(new_n20091_), .A2(new_n20092_), .ZN(new_n20095_));
  NAND2_X1   g19839(.A1(new_n20094_), .A2(new_n20095_), .ZN(new_n20096_));
  XOR2_X1    g19840(.A1(new_n20096_), .A2(new_n20023_), .Z(new_n20097_));
  XOR2_X1    g19841(.A1(new_n20097_), .A2(new_n20018_), .Z(new_n20098_));
  INV_X1     g19842(.I(new_n19988_), .ZN(new_n20099_));
  NAND2_X1   g19843(.A1(new_n19997_), .A2(new_n20099_), .ZN(new_n20100_));
  NAND2_X1   g19844(.A1(new_n20100_), .A2(new_n19996_), .ZN(new_n20101_));
  XOR2_X1    g19845(.A1(new_n20101_), .A2(\a[41] ), .Z(new_n20102_));
  XOR2_X1    g19846(.A1(new_n20098_), .A2(new_n20102_), .Z(new_n20103_));
  NOR2_X1    g19847(.A1(new_n20103_), .A2(new_n20017_), .ZN(new_n20104_));
  INV_X1     g19848(.I(new_n20104_), .ZN(new_n20105_));
  NAND2_X1   g19849(.A1(new_n20103_), .A2(new_n20017_), .ZN(new_n20106_));
  NAND2_X1   g19850(.A1(new_n20105_), .A2(new_n20106_), .ZN(new_n20107_));
  XOR2_X1    g19851(.A1(new_n20015_), .A2(new_n20107_), .Z(\f[104] ));
  AOI21_X1   g19852(.A1(new_n20015_), .A2(new_n20106_), .B(new_n20104_), .ZN(new_n20109_));
  AOI22_X1   g19853(.A1(new_n6569_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n6574_), .ZN(new_n20110_));
  OAI21_X1   g19854(.A1(new_n12148_), .A2(new_n8565_), .B(new_n20110_), .ZN(new_n20111_));
  AOI21_X1   g19855(.A1(new_n12811_), .A2(new_n6579_), .B(new_n20111_), .ZN(new_n20112_));
  XOR2_X1    g19856(.A1(new_n20112_), .A2(new_n6567_), .Z(new_n20113_));
  AOI21_X1   g19857(.A1(new_n20023_), .A2(new_n20095_), .B(new_n20093_), .ZN(new_n20114_));
  OAI21_X1   g19858(.A1(new_n20027_), .A2(new_n20077_), .B(new_n20079_), .ZN(new_n20115_));
  AOI22_X1   g19859(.A1(new_n8241_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n8246_), .ZN(new_n20116_));
  OAI21_X1   g19860(.A1(new_n9972_), .A2(new_n9114_), .B(new_n20116_), .ZN(new_n20117_));
  AOI21_X1   g19861(.A1(new_n10631_), .A2(new_n8252_), .B(new_n20117_), .ZN(new_n20118_));
  XOR2_X1    g19862(.A1(new_n20118_), .A2(new_n8248_), .Z(new_n20119_));
  INV_X1     g19863(.I(new_n20119_), .ZN(new_n20120_));
  AOI21_X1   g19864(.A1(new_n20036_), .A2(new_n20074_), .B(new_n20072_), .ZN(new_n20121_));
  INV_X1     g19865(.I(new_n20121_), .ZN(new_n20122_));
  AOI22_X1   g19866(.A1(new_n9125_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n9123_), .ZN(new_n20123_));
  OAI21_X1   g19867(.A1(new_n9032_), .A2(new_n9470_), .B(new_n20123_), .ZN(new_n20124_));
  AOI21_X1   g19868(.A1(new_n10884_), .A2(new_n9129_), .B(new_n20124_), .ZN(new_n20125_));
  XOR2_X1    g19869(.A1(new_n20125_), .A2(new_n9133_), .Z(new_n20126_));
  OAI21_X1   g19870(.A1(new_n20040_), .A2(new_n20064_), .B(new_n20066_), .ZN(new_n20127_));
  AOI22_X1   g19871(.A1(new_n10064_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n10062_), .ZN(new_n20128_));
  OAI21_X1   g19872(.A1(new_n8168_), .A2(new_n10399_), .B(new_n20128_), .ZN(new_n20129_));
  AOI21_X1   g19873(.A1(new_n8783_), .A2(new_n10068_), .B(new_n20129_), .ZN(new_n20130_));
  XOR2_X1    g19874(.A1(new_n20130_), .A2(new_n10057_), .Z(new_n20131_));
  INV_X1     g19875(.I(new_n20131_), .ZN(new_n20132_));
  AOI21_X1   g19876(.A1(new_n20055_), .A2(new_n20060_), .B(new_n20058_), .ZN(new_n20133_));
  AOI22_X1   g19877(.A1(new_n11926_), .A2(\b[45] ), .B1(new_n11924_), .B2(\b[44] ), .ZN(new_n20134_));
  OAI21_X1   g19878(.A1(new_n6775_), .A2(new_n12317_), .B(new_n20134_), .ZN(new_n20135_));
  AOI21_X1   g19879(.A1(new_n7926_), .A2(new_n11929_), .B(new_n20135_), .ZN(new_n20136_));
  XOR2_X1    g19880(.A1(new_n20136_), .A2(new_n12312_), .Z(new_n20137_));
  INV_X1     g19881(.I(new_n20137_), .ZN(new_n20138_));
  AOI22_X1   g19882(.A1(new_n12922_), .A2(\b[42] ), .B1(\b[41] ), .B2(new_n12923_), .ZN(new_n20139_));
  INV_X1     g19883(.I(new_n20139_), .ZN(new_n20140_));
  NOR2_X1    g19884(.A1(new_n20140_), .A2(new_n5849_), .ZN(new_n20141_));
  NOR2_X1    g19885(.A1(new_n20139_), .A2(\a[41] ), .ZN(new_n20142_));
  NOR2_X1    g19886(.A1(new_n20141_), .A2(new_n20142_), .ZN(new_n20143_));
  XOR2_X1    g19887(.A1(new_n20143_), .A2(new_n19945_), .Z(new_n20144_));
  NOR2_X1    g19888(.A1(new_n20138_), .A2(new_n20144_), .ZN(new_n20145_));
  INV_X1     g19889(.I(new_n20145_), .ZN(new_n20146_));
  NAND2_X1   g19890(.A1(new_n20138_), .A2(new_n20144_), .ZN(new_n20147_));
  NAND2_X1   g19891(.A1(new_n20146_), .A2(new_n20147_), .ZN(new_n20148_));
  XOR2_X1    g19892(.A1(new_n20148_), .A2(new_n20133_), .Z(new_n20149_));
  AOI22_X1   g19893(.A1(new_n10981_), .A2(\b[48] ), .B1(new_n10979_), .B2(\b[47] ), .ZN(new_n20150_));
  OAI21_X1   g19894(.A1(new_n7617_), .A2(new_n11306_), .B(new_n20150_), .ZN(new_n20151_));
  AOI21_X1   g19895(.A1(new_n8792_), .A2(new_n10984_), .B(new_n20151_), .ZN(new_n20152_));
  XOR2_X1    g19896(.A1(new_n20152_), .A2(\a[59] ), .Z(new_n20153_));
  INV_X1     g19897(.I(new_n20052_), .ZN(new_n20154_));
  OAI21_X1   g19898(.A1(new_n20154_), .A2(new_n20062_), .B(new_n20051_), .ZN(new_n20155_));
  NAND2_X1   g19899(.A1(new_n20155_), .A2(new_n20153_), .ZN(new_n20156_));
  OR2_X2     g19900(.A1(new_n20155_), .A2(new_n20153_), .Z(new_n20157_));
  NAND2_X1   g19901(.A1(new_n20157_), .A2(new_n20156_), .ZN(new_n20158_));
  XNOR2_X1   g19902(.A1(new_n20158_), .A2(new_n20149_), .ZN(new_n20159_));
  NOR2_X1    g19903(.A1(new_n20159_), .A2(new_n20132_), .ZN(new_n20160_));
  INV_X1     g19904(.I(new_n20160_), .ZN(new_n20161_));
  NAND2_X1   g19905(.A1(new_n20159_), .A2(new_n20132_), .ZN(new_n20162_));
  NAND2_X1   g19906(.A1(new_n20161_), .A2(new_n20162_), .ZN(new_n20163_));
  XOR2_X1    g19907(.A1(new_n20163_), .A2(new_n20127_), .Z(new_n20164_));
  NOR2_X1    g19908(.A1(new_n20164_), .A2(new_n20126_), .ZN(new_n20165_));
  NAND2_X1   g19909(.A1(new_n20164_), .A2(new_n20126_), .ZN(new_n20166_));
  INV_X1     g19910(.I(new_n20166_), .ZN(new_n20167_));
  NOR2_X1    g19911(.A1(new_n20167_), .A2(new_n20165_), .ZN(new_n20168_));
  XOR2_X1    g19912(.A1(new_n20168_), .A2(new_n20122_), .Z(new_n20169_));
  NOR2_X1    g19913(.A1(new_n20169_), .A2(new_n20120_), .ZN(new_n20170_));
  NAND2_X1   g19914(.A1(new_n20169_), .A2(new_n20120_), .ZN(new_n20171_));
  INV_X1     g19915(.I(new_n20171_), .ZN(new_n20172_));
  NOR2_X1    g19916(.A1(new_n20172_), .A2(new_n20170_), .ZN(new_n20173_));
  XOR2_X1    g19917(.A1(new_n20173_), .A2(new_n20115_), .Z(new_n20174_));
  AOI22_X1   g19918(.A1(new_n7403_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n7408_), .ZN(new_n20175_));
  OAI21_X1   g19919(.A1(new_n11195_), .A2(new_n9488_), .B(new_n20175_), .ZN(new_n20176_));
  AOI21_X1   g19920(.A1(new_n11836_), .A2(new_n7414_), .B(new_n20176_), .ZN(new_n20177_));
  XOR2_X1    g19921(.A1(new_n20177_), .A2(new_n7410_), .Z(new_n20178_));
  NAND2_X1   g19922(.A1(new_n20081_), .A2(new_n20089_), .ZN(new_n20179_));
  NAND2_X1   g19923(.A1(new_n20179_), .A2(new_n20088_), .ZN(new_n20180_));
  INV_X1     g19924(.I(new_n20180_), .ZN(new_n20181_));
  NOR2_X1    g19925(.A1(new_n20181_), .A2(new_n20178_), .ZN(new_n20182_));
  INV_X1     g19926(.I(new_n20182_), .ZN(new_n20183_));
  NAND2_X1   g19927(.A1(new_n20181_), .A2(new_n20178_), .ZN(new_n20184_));
  NAND2_X1   g19928(.A1(new_n20183_), .A2(new_n20184_), .ZN(new_n20185_));
  XOR2_X1    g19929(.A1(new_n20185_), .A2(new_n20174_), .Z(new_n20186_));
  NAND2_X1   g19930(.A1(new_n20186_), .A2(new_n20114_), .ZN(new_n20187_));
  NOR2_X1    g19931(.A1(new_n20186_), .A2(new_n20114_), .ZN(new_n20188_));
  INV_X1     g19932(.I(new_n20188_), .ZN(new_n20189_));
  NAND2_X1   g19933(.A1(new_n20189_), .A2(new_n20187_), .ZN(new_n20190_));
  XOR2_X1    g19934(.A1(new_n20190_), .A2(new_n20113_), .Z(new_n20191_));
  INV_X1     g19935(.I(new_n20097_), .ZN(new_n20192_));
  INV_X1     g19936(.I(new_n20101_), .ZN(new_n20193_));
  XOR2_X1    g19937(.A1(new_n20018_), .A2(new_n5849_), .Z(new_n20194_));
  AOI21_X1   g19938(.A1(new_n20097_), .A2(new_n20193_), .B(new_n20194_), .ZN(new_n20195_));
  AOI21_X1   g19939(.A1(new_n20192_), .A2(new_n20101_), .B(new_n20195_), .ZN(new_n20196_));
  INV_X1     g19940(.I(new_n20196_), .ZN(new_n20197_));
  NOR2_X1    g19941(.A1(new_n20191_), .A2(new_n20197_), .ZN(new_n20198_));
  INV_X1     g19942(.I(new_n20198_), .ZN(new_n20199_));
  NAND2_X1   g19943(.A1(new_n20191_), .A2(new_n20197_), .ZN(new_n20200_));
  AND2_X2    g19944(.A1(new_n20199_), .A2(new_n20200_), .Z(new_n20201_));
  XOR2_X1    g19945(.A1(new_n20109_), .A2(new_n20201_), .Z(\f[105] ));
  OAI22_X1   g19946(.A1(new_n8565_), .A2(new_n12796_), .B1(new_n12800_), .B2(new_n7731_), .ZN(new_n20203_));
  AOI21_X1   g19947(.A1(new_n13973_), .A2(new_n6579_), .B(new_n20203_), .ZN(new_n20204_));
  XOR2_X1    g19948(.A1(new_n20204_), .A2(new_n6567_), .Z(new_n20205_));
  INV_X1     g19949(.I(new_n20205_), .ZN(new_n20206_));
  NAND2_X1   g19950(.A1(new_n20184_), .A2(new_n20174_), .ZN(new_n20207_));
  NAND2_X1   g19951(.A1(new_n20207_), .A2(new_n20183_), .ZN(new_n20208_));
  INV_X1     g19952(.I(new_n20208_), .ZN(new_n20209_));
  OAI22_X1   g19953(.A1(new_n12147_), .A2(new_n8588_), .B1(new_n8587_), .B2(new_n12148_), .ZN(new_n20210_));
  AOI21_X1   g19954(.A1(\b[59] ), .A2(new_n7719_), .B(new_n20210_), .ZN(new_n20211_));
  OAI21_X1   g19955(.A1(new_n13110_), .A2(new_n8585_), .B(new_n20211_), .ZN(new_n20212_));
  XOR2_X1    g19956(.A1(new_n20212_), .A2(new_n7410_), .Z(new_n20213_));
  INV_X1     g19957(.I(new_n20170_), .ZN(new_n20214_));
  AOI21_X1   g19958(.A1(new_n20115_), .A2(new_n20214_), .B(new_n20172_), .ZN(new_n20215_));
  AOI22_X1   g19959(.A1(new_n8241_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n8246_), .ZN(new_n20216_));
  OAI21_X1   g19960(.A1(new_n10308_), .A2(new_n9114_), .B(new_n20216_), .ZN(new_n20217_));
  AOI21_X1   g19961(.A1(new_n12164_), .A2(new_n8252_), .B(new_n20217_), .ZN(new_n20218_));
  XOR2_X1    g19962(.A1(new_n20218_), .A2(new_n8248_), .Z(new_n20219_));
  AOI21_X1   g19963(.A1(new_n20122_), .A2(new_n20166_), .B(new_n20165_), .ZN(new_n20220_));
  AOI22_X1   g19964(.A1(new_n10064_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n10062_), .ZN(new_n20221_));
  OAI21_X1   g19965(.A1(new_n8500_), .A2(new_n10399_), .B(new_n20221_), .ZN(new_n20222_));
  AOI21_X1   g19966(.A1(new_n9987_), .A2(new_n10068_), .B(new_n20222_), .ZN(new_n20223_));
  XOR2_X1    g19967(.A1(new_n20223_), .A2(new_n10057_), .Z(new_n20224_));
  INV_X1     g19968(.I(new_n20224_), .ZN(new_n20225_));
  OAI21_X1   g19969(.A1(new_n20133_), .A2(new_n20145_), .B(new_n20147_), .ZN(new_n20226_));
  AOI22_X1   g19970(.A1(new_n11926_), .A2(\b[46] ), .B1(new_n11924_), .B2(\b[45] ), .ZN(new_n20227_));
  OAI21_X1   g19971(.A1(new_n7074_), .A2(new_n12317_), .B(new_n20227_), .ZN(new_n20228_));
  AOI21_X1   g19972(.A1(new_n9337_), .A2(new_n11929_), .B(new_n20228_), .ZN(new_n20229_));
  XOR2_X1    g19973(.A1(new_n20229_), .A2(\a[62] ), .Z(new_n20230_));
  INV_X1     g19974(.I(new_n20142_), .ZN(new_n20231_));
  AOI21_X1   g19975(.A1(new_n19945_), .A2(new_n20231_), .B(new_n20141_), .ZN(new_n20232_));
  AOI22_X1   g19976(.A1(new_n12922_), .A2(\b[43] ), .B1(\b[42] ), .B2(new_n12923_), .ZN(new_n20233_));
  NAND2_X1   g19977(.A1(new_n20232_), .A2(new_n20233_), .ZN(new_n20234_));
  NOR2_X1    g19978(.A1(new_n20232_), .A2(new_n20233_), .ZN(new_n20235_));
  INV_X1     g19979(.I(new_n20235_), .ZN(new_n20236_));
  NAND2_X1   g19980(.A1(new_n20236_), .A2(new_n20234_), .ZN(new_n20237_));
  XNOR2_X1   g19981(.A1(new_n20230_), .A2(new_n20237_), .ZN(new_n20238_));
  INV_X1     g19982(.I(new_n20238_), .ZN(new_n20239_));
  OAI22_X1   g19983(.A1(new_n12306_), .A2(new_n8168_), .B1(new_n12305_), .B2(new_n8127_), .ZN(new_n20240_));
  AOI21_X1   g19984(.A1(\b[47] ), .A2(new_n12304_), .B(new_n20240_), .ZN(new_n20241_));
  OAI21_X1   g19985(.A1(new_n9050_), .A2(new_n10985_), .B(new_n20241_), .ZN(new_n20242_));
  XOR2_X1    g19986(.A1(new_n20242_), .A2(\a[59] ), .Z(new_n20243_));
  NOR2_X1    g19987(.A1(new_n20243_), .A2(new_n20239_), .ZN(new_n20244_));
  NAND2_X1   g19988(.A1(new_n20243_), .A2(new_n20239_), .ZN(new_n20245_));
  INV_X1     g19989(.I(new_n20245_), .ZN(new_n20246_));
  NOR2_X1    g19990(.A1(new_n20246_), .A2(new_n20244_), .ZN(new_n20247_));
  XNOR2_X1   g19991(.A1(new_n20247_), .A2(new_n20226_), .ZN(new_n20248_));
  INV_X1     g19992(.I(new_n20156_), .ZN(new_n20249_));
  AOI21_X1   g19993(.A1(new_n20149_), .A2(new_n20157_), .B(new_n20249_), .ZN(new_n20250_));
  NOR2_X1    g19994(.A1(new_n20248_), .A2(new_n20250_), .ZN(new_n20251_));
  INV_X1     g19995(.I(new_n20251_), .ZN(new_n20252_));
  NAND2_X1   g19996(.A1(new_n20248_), .A2(new_n20250_), .ZN(new_n20253_));
  NAND2_X1   g19997(.A1(new_n20252_), .A2(new_n20253_), .ZN(new_n20254_));
  XOR2_X1    g19998(.A1(new_n20254_), .A2(new_n20225_), .Z(new_n20255_));
  INV_X1     g19999(.I(new_n20162_), .ZN(new_n20256_));
  AOI21_X1   g20000(.A1(new_n20127_), .A2(new_n20161_), .B(new_n20256_), .ZN(new_n20257_));
  AOI22_X1   g20001(.A1(new_n9125_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n9123_), .ZN(new_n20258_));
  OAI21_X1   g20002(.A1(new_n9376_), .A2(new_n9470_), .B(new_n20258_), .ZN(new_n20259_));
  AOI21_X1   g20003(.A1(new_n9979_), .A2(new_n9129_), .B(new_n20259_), .ZN(new_n20260_));
  XOR2_X1    g20004(.A1(new_n20260_), .A2(new_n9133_), .Z(new_n20261_));
  NOR2_X1    g20005(.A1(new_n20257_), .A2(new_n20261_), .ZN(new_n20262_));
  NAND2_X1   g20006(.A1(new_n20257_), .A2(new_n20261_), .ZN(new_n20263_));
  INV_X1     g20007(.I(new_n20263_), .ZN(new_n20264_));
  NOR2_X1    g20008(.A1(new_n20264_), .A2(new_n20262_), .ZN(new_n20265_));
  XOR2_X1    g20009(.A1(new_n20265_), .A2(new_n20255_), .Z(new_n20266_));
  NOR2_X1    g20010(.A1(new_n20266_), .A2(new_n20220_), .ZN(new_n20267_));
  INV_X1     g20011(.I(new_n20267_), .ZN(new_n20268_));
  NAND2_X1   g20012(.A1(new_n20266_), .A2(new_n20220_), .ZN(new_n20269_));
  NAND2_X1   g20013(.A1(new_n20268_), .A2(new_n20269_), .ZN(new_n20270_));
  XOR2_X1    g20014(.A1(new_n20270_), .A2(new_n20219_), .Z(new_n20271_));
  INV_X1     g20015(.I(new_n20271_), .ZN(new_n20272_));
  NAND2_X1   g20016(.A1(new_n20272_), .A2(new_n20215_), .ZN(new_n20273_));
  INV_X1     g20017(.I(new_n20215_), .ZN(new_n20274_));
  NAND2_X1   g20018(.A1(new_n20274_), .A2(new_n20271_), .ZN(new_n20275_));
  NAND2_X1   g20019(.A1(new_n20273_), .A2(new_n20275_), .ZN(new_n20276_));
  XOR2_X1    g20020(.A1(new_n20276_), .A2(new_n20213_), .Z(new_n20277_));
  NOR2_X1    g20021(.A1(new_n20209_), .A2(new_n20277_), .ZN(new_n20278_));
  INV_X1     g20022(.I(new_n20278_), .ZN(new_n20279_));
  NAND2_X1   g20023(.A1(new_n20209_), .A2(new_n20277_), .ZN(new_n20280_));
  NAND2_X1   g20024(.A1(new_n20279_), .A2(new_n20280_), .ZN(new_n20281_));
  XOR2_X1    g20025(.A1(new_n20281_), .A2(new_n20206_), .Z(new_n20282_));
  INV_X1     g20026(.I(new_n20113_), .ZN(new_n20283_));
  AOI21_X1   g20027(.A1(new_n20283_), .A2(new_n20187_), .B(new_n20188_), .ZN(new_n20284_));
  INV_X1     g20028(.I(new_n20284_), .ZN(new_n20285_));
  AOI21_X1   g20029(.A1(new_n20109_), .A2(new_n20201_), .B(new_n20198_), .ZN(new_n20286_));
  NOR2_X1    g20030(.A1(new_n20286_), .A2(new_n20285_), .ZN(new_n20287_));
  NOR3_X1    g20031(.A1(new_n19911_), .A2(new_n19906_), .A3(new_n20007_), .ZN(new_n20288_));
  AOI21_X1   g20032(.A1(new_n20005_), .A2(new_n20008_), .B(new_n20288_), .ZN(new_n20289_));
  INV_X1     g20033(.I(new_n20106_), .ZN(new_n20290_));
  OAI21_X1   g20034(.A1(new_n20289_), .A2(new_n20290_), .B(new_n20105_), .ZN(new_n20291_));
  INV_X1     g20035(.I(new_n20201_), .ZN(new_n20292_));
  OAI21_X1   g20036(.A1(new_n20291_), .A2(new_n20292_), .B(new_n20199_), .ZN(new_n20293_));
  NOR2_X1    g20037(.A1(new_n20293_), .A2(new_n20284_), .ZN(new_n20294_));
  NOR2_X1    g20038(.A1(new_n20294_), .A2(new_n20287_), .ZN(new_n20295_));
  XOR2_X1    g20039(.A1(new_n20295_), .A2(new_n20282_), .Z(\f[106] ));
  NAND2_X1   g20040(.A1(new_n20286_), .A2(new_n20285_), .ZN(new_n20297_));
  INV_X1     g20041(.I(new_n20282_), .ZN(new_n20298_));
  OAI21_X1   g20042(.A1(new_n20286_), .A2(new_n20285_), .B(new_n20298_), .ZN(new_n20299_));
  NAND2_X1   g20043(.A1(new_n20299_), .A2(new_n20297_), .ZN(new_n20300_));
  AOI21_X1   g20044(.A1(new_n20206_), .A2(new_n20280_), .B(new_n20278_), .ZN(new_n20301_));
  AOI22_X1   g20045(.A1(new_n13460_), .A2(new_n6579_), .B1(\b[63] ), .B2(new_n6887_), .ZN(new_n20302_));
  AOI22_X1   g20046(.A1(new_n7403_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n7408_), .ZN(new_n20303_));
  OAI21_X1   g20047(.A1(new_n12147_), .A2(new_n9488_), .B(new_n20303_), .ZN(new_n20304_));
  AOI21_X1   g20048(.A1(new_n13444_), .A2(new_n7414_), .B(new_n20304_), .ZN(new_n20305_));
  XOR2_X1    g20049(.A1(new_n20305_), .A2(\a[47] ), .Z(new_n20306_));
  AOI22_X1   g20050(.A1(new_n9125_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n9123_), .ZN(new_n20307_));
  OAI21_X1   g20051(.A1(new_n9942_), .A2(new_n9470_), .B(new_n20307_), .ZN(new_n20308_));
  AOI21_X1   g20052(.A1(new_n10318_), .A2(new_n9129_), .B(new_n20308_), .ZN(new_n20309_));
  XOR2_X1    g20053(.A1(new_n20309_), .A2(new_n9133_), .Z(new_n20310_));
  AOI21_X1   g20054(.A1(new_n20225_), .A2(new_n20253_), .B(new_n20251_), .ZN(new_n20311_));
  INV_X1     g20055(.I(new_n20311_), .ZN(new_n20312_));
  OAI22_X1   g20056(.A1(new_n11298_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n11297_), .ZN(new_n20313_));
  AOI21_X1   g20057(.A1(\b[51] ), .A2(new_n11296_), .B(new_n20313_), .ZN(new_n20314_));
  OAI21_X1   g20058(.A1(new_n9385_), .A2(new_n10069_), .B(new_n20314_), .ZN(new_n20315_));
  XOR2_X1    g20059(.A1(new_n20315_), .A2(new_n10057_), .Z(new_n20316_));
  AOI22_X1   g20060(.A1(new_n10981_), .A2(\b[50] ), .B1(new_n10979_), .B2(\b[49] ), .ZN(new_n20317_));
  OAI21_X1   g20061(.A1(new_n8127_), .A2(new_n11306_), .B(new_n20317_), .ZN(new_n20318_));
  AOI21_X1   g20062(.A1(new_n9684_), .A2(new_n10984_), .B(new_n20318_), .ZN(new_n20319_));
  XOR2_X1    g20063(.A1(new_n20319_), .A2(new_n10989_), .Z(new_n20320_));
  AOI21_X1   g20064(.A1(new_n20230_), .A2(new_n20234_), .B(new_n20235_), .ZN(new_n20321_));
  INV_X1     g20065(.I(new_n20321_), .ZN(new_n20322_));
  AOI22_X1   g20066(.A1(new_n11926_), .A2(\b[47] ), .B1(new_n11924_), .B2(\b[46] ), .ZN(new_n20323_));
  OAI21_X1   g20067(.A1(new_n7096_), .A2(new_n12317_), .B(new_n20323_), .ZN(new_n20324_));
  AOI21_X1   g20068(.A1(new_n7649_), .A2(new_n11929_), .B(new_n20324_), .ZN(new_n20325_));
  XOR2_X1    g20069(.A1(new_n20325_), .A2(\a[62] ), .Z(new_n20326_));
  INV_X1     g20070(.I(new_n20233_), .ZN(new_n20327_));
  AOI22_X1   g20071(.A1(new_n12922_), .A2(\b[44] ), .B1(\b[43] ), .B2(new_n12923_), .ZN(new_n20328_));
  NAND2_X1   g20072(.A1(new_n20327_), .A2(new_n20328_), .ZN(new_n20329_));
  INV_X1     g20073(.I(new_n20328_), .ZN(new_n20330_));
  NAND2_X1   g20074(.A1(new_n20330_), .A2(new_n20233_), .ZN(new_n20331_));
  NAND2_X1   g20075(.A1(new_n20329_), .A2(new_n20331_), .ZN(new_n20332_));
  XNOR2_X1   g20076(.A1(new_n20326_), .A2(new_n20332_), .ZN(new_n20333_));
  NOR2_X1    g20077(.A1(new_n20333_), .A2(new_n20322_), .ZN(new_n20334_));
  INV_X1     g20078(.I(new_n20334_), .ZN(new_n20335_));
  NAND2_X1   g20079(.A1(new_n20333_), .A2(new_n20322_), .ZN(new_n20336_));
  NAND2_X1   g20080(.A1(new_n20335_), .A2(new_n20336_), .ZN(new_n20337_));
  XOR2_X1    g20081(.A1(new_n20337_), .A2(new_n20320_), .Z(new_n20338_));
  INV_X1     g20082(.I(new_n20338_), .ZN(new_n20339_));
  AOI21_X1   g20083(.A1(new_n20226_), .A2(new_n20245_), .B(new_n20244_), .ZN(new_n20340_));
  NOR2_X1    g20084(.A1(new_n20339_), .A2(new_n20340_), .ZN(new_n20341_));
  INV_X1     g20085(.I(new_n20341_), .ZN(new_n20342_));
  NAND2_X1   g20086(.A1(new_n20339_), .A2(new_n20340_), .ZN(new_n20343_));
  NAND2_X1   g20087(.A1(new_n20342_), .A2(new_n20343_), .ZN(new_n20344_));
  XNOR2_X1   g20088(.A1(new_n20344_), .A2(new_n20316_), .ZN(new_n20345_));
  NOR2_X1    g20089(.A1(new_n20345_), .A2(new_n20312_), .ZN(new_n20346_));
  NAND2_X1   g20090(.A1(new_n20345_), .A2(new_n20312_), .ZN(new_n20347_));
  INV_X1     g20091(.I(new_n20347_), .ZN(new_n20348_));
  NOR2_X1    g20092(.A1(new_n20348_), .A2(new_n20346_), .ZN(new_n20349_));
  XOR2_X1    g20093(.A1(new_n20349_), .A2(new_n20310_), .Z(new_n20350_));
  OAI22_X1   g20094(.A1(new_n9461_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n9462_), .ZN(new_n20351_));
  AOI21_X1   g20095(.A1(\b[57] ), .A2(new_n8575_), .B(new_n20351_), .ZN(new_n20352_));
  OAI21_X1   g20096(.A1(new_n12203_), .A2(new_n9460_), .B(new_n20352_), .ZN(new_n20353_));
  XOR2_X1    g20097(.A1(new_n20353_), .A2(\a[50] ), .Z(new_n20354_));
  INV_X1     g20098(.I(new_n20255_), .ZN(new_n20355_));
  AOI21_X1   g20099(.A1(new_n20355_), .A2(new_n20263_), .B(new_n20262_), .ZN(new_n20356_));
  NOR2_X1    g20100(.A1(new_n20356_), .A2(new_n20354_), .ZN(new_n20357_));
  AND2_X2    g20101(.A1(new_n20356_), .A2(new_n20354_), .Z(new_n20358_));
  NOR2_X1    g20102(.A1(new_n20358_), .A2(new_n20357_), .ZN(new_n20359_));
  XOR2_X1    g20103(.A1(new_n20350_), .A2(new_n20359_), .Z(new_n20360_));
  INV_X1     g20104(.I(new_n20219_), .ZN(new_n20361_));
  AOI21_X1   g20105(.A1(new_n20361_), .A2(new_n20269_), .B(new_n20267_), .ZN(new_n20362_));
  OR2_X2     g20106(.A1(new_n20360_), .A2(new_n20362_), .Z(new_n20363_));
  NAND2_X1   g20107(.A1(new_n20360_), .A2(new_n20362_), .ZN(new_n20364_));
  NAND2_X1   g20108(.A1(new_n20363_), .A2(new_n20364_), .ZN(new_n20365_));
  XOR2_X1    g20109(.A1(new_n20365_), .A2(new_n20306_), .Z(new_n20366_));
  XOR2_X1    g20110(.A1(new_n20366_), .A2(new_n20302_), .Z(new_n20367_));
  NAND2_X1   g20111(.A1(new_n20273_), .A2(new_n20213_), .ZN(new_n20368_));
  NAND2_X1   g20112(.A1(new_n20368_), .A2(new_n20275_), .ZN(new_n20369_));
  XOR2_X1    g20113(.A1(new_n20369_), .A2(\a[44] ), .Z(new_n20370_));
  XOR2_X1    g20114(.A1(new_n20367_), .A2(new_n20370_), .Z(new_n20371_));
  NOR2_X1    g20115(.A1(new_n20371_), .A2(new_n20301_), .ZN(new_n20372_));
  INV_X1     g20116(.I(new_n20372_), .ZN(new_n20373_));
  NAND2_X1   g20117(.A1(new_n20371_), .A2(new_n20301_), .ZN(new_n20374_));
  NAND2_X1   g20118(.A1(new_n20373_), .A2(new_n20374_), .ZN(new_n20375_));
  XOR2_X1    g20119(.A1(new_n20300_), .A2(new_n20375_), .Z(\f[107] ));
  INV_X1     g20120(.I(new_n20374_), .ZN(new_n20377_));
  AOI21_X1   g20121(.A1(new_n20299_), .A2(new_n20297_), .B(new_n20377_), .ZN(new_n20378_));
  AOI22_X1   g20122(.A1(new_n7403_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n7408_), .ZN(new_n20379_));
  OAI21_X1   g20123(.A1(new_n12148_), .A2(new_n9488_), .B(new_n20379_), .ZN(new_n20380_));
  AOI21_X1   g20124(.A1(new_n12811_), .A2(new_n7414_), .B(new_n20380_), .ZN(new_n20381_));
  XOR2_X1    g20125(.A1(new_n20381_), .A2(new_n7410_), .Z(new_n20382_));
  NAND2_X1   g20126(.A1(new_n20364_), .A2(new_n20306_), .ZN(new_n20383_));
  NAND2_X1   g20127(.A1(new_n20383_), .A2(new_n20363_), .ZN(new_n20384_));
  NOR2_X1    g20128(.A1(new_n20350_), .A2(new_n20358_), .ZN(new_n20385_));
  NOR2_X1    g20129(.A1(new_n20385_), .A2(new_n20357_), .ZN(new_n20386_));
  AOI22_X1   g20130(.A1(new_n8241_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n8246_), .ZN(new_n20387_));
  OAI21_X1   g20131(.A1(new_n11195_), .A2(new_n9114_), .B(new_n20387_), .ZN(new_n20388_));
  AOI21_X1   g20132(.A1(new_n11836_), .A2(new_n8252_), .B(new_n20388_), .ZN(new_n20389_));
  XOR2_X1    g20133(.A1(new_n20389_), .A2(\a[50] ), .Z(new_n20390_));
  OAI21_X1   g20134(.A1(new_n20310_), .A2(new_n20346_), .B(new_n20347_), .ZN(new_n20391_));
  INV_X1     g20135(.I(new_n20391_), .ZN(new_n20392_));
  AOI22_X1   g20136(.A1(new_n9125_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n9123_), .ZN(new_n20393_));
  OAI21_X1   g20137(.A1(new_n9972_), .A2(new_n9470_), .B(new_n20393_), .ZN(new_n20394_));
  AOI21_X1   g20138(.A1(new_n10631_), .A2(new_n9129_), .B(new_n20394_), .ZN(new_n20395_));
  XOR2_X1    g20139(.A1(new_n20395_), .A2(new_n9133_), .Z(new_n20396_));
  INV_X1     g20140(.I(new_n20396_), .ZN(new_n20397_));
  AOI21_X1   g20141(.A1(new_n20316_), .A2(new_n20343_), .B(new_n20341_), .ZN(new_n20398_));
  AOI22_X1   g20142(.A1(new_n10064_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n10062_), .ZN(new_n20399_));
  OAI21_X1   g20143(.A1(new_n9032_), .A2(new_n10399_), .B(new_n20399_), .ZN(new_n20400_));
  AOI21_X1   g20144(.A1(new_n10884_), .A2(new_n10068_), .B(new_n20400_), .ZN(new_n20401_));
  XOR2_X1    g20145(.A1(new_n20401_), .A2(new_n10057_), .Z(new_n20402_));
  INV_X1     g20146(.I(new_n20402_), .ZN(new_n20403_));
  OAI21_X1   g20147(.A1(new_n20320_), .A2(new_n20334_), .B(new_n20336_), .ZN(new_n20404_));
  NAND2_X1   g20148(.A1(new_n20326_), .A2(new_n20331_), .ZN(new_n20405_));
  NAND2_X1   g20149(.A1(new_n20405_), .A2(new_n20329_), .ZN(new_n20406_));
  AOI22_X1   g20150(.A1(new_n11926_), .A2(\b[48] ), .B1(new_n11924_), .B2(\b[47] ), .ZN(new_n20407_));
  OAI21_X1   g20151(.A1(new_n7617_), .A2(new_n12317_), .B(new_n20407_), .ZN(new_n20408_));
  AOI21_X1   g20152(.A1(new_n8792_), .A2(new_n11929_), .B(new_n20408_), .ZN(new_n20409_));
  XOR2_X1    g20153(.A1(new_n20409_), .A2(new_n12312_), .Z(new_n20410_));
  AOI22_X1   g20154(.A1(new_n12922_), .A2(\b[45] ), .B1(\b[44] ), .B2(new_n12923_), .ZN(new_n20411_));
  XOR2_X1    g20155(.A1(new_n20411_), .A2(new_n6567_), .Z(new_n20412_));
  XOR2_X1    g20156(.A1(new_n20412_), .A2(new_n20233_), .Z(new_n20413_));
  NOR2_X1    g20157(.A1(new_n20410_), .A2(new_n20413_), .ZN(new_n20414_));
  NAND2_X1   g20158(.A1(new_n20410_), .A2(new_n20413_), .ZN(new_n20415_));
  INV_X1     g20159(.I(new_n20415_), .ZN(new_n20416_));
  NOR2_X1    g20160(.A1(new_n20416_), .A2(new_n20414_), .ZN(new_n20417_));
  XNOR2_X1   g20161(.A1(new_n20417_), .A2(new_n20406_), .ZN(new_n20418_));
  AOI22_X1   g20162(.A1(new_n10981_), .A2(\b[51] ), .B1(new_n10979_), .B2(\b[50] ), .ZN(new_n20419_));
  OAI21_X1   g20163(.A1(new_n8168_), .A2(new_n11306_), .B(new_n20419_), .ZN(new_n20420_));
  AOI21_X1   g20164(.A1(new_n8783_), .A2(new_n10984_), .B(new_n20420_), .ZN(new_n20421_));
  XOR2_X1    g20165(.A1(new_n20421_), .A2(new_n10989_), .Z(new_n20422_));
  NOR2_X1    g20166(.A1(new_n20418_), .A2(new_n20422_), .ZN(new_n20423_));
  NAND2_X1   g20167(.A1(new_n20418_), .A2(new_n20422_), .ZN(new_n20424_));
  INV_X1     g20168(.I(new_n20424_), .ZN(new_n20425_));
  NOR2_X1    g20169(.A1(new_n20425_), .A2(new_n20423_), .ZN(new_n20426_));
  XOR2_X1    g20170(.A1(new_n20426_), .A2(new_n20404_), .Z(new_n20427_));
  NOR2_X1    g20171(.A1(new_n20427_), .A2(new_n20403_), .ZN(new_n20428_));
  NAND2_X1   g20172(.A1(new_n20427_), .A2(new_n20403_), .ZN(new_n20429_));
  INV_X1     g20173(.I(new_n20429_), .ZN(new_n20430_));
  NOR2_X1    g20174(.A1(new_n20430_), .A2(new_n20428_), .ZN(new_n20431_));
  XNOR2_X1   g20175(.A1(new_n20431_), .A2(new_n20398_), .ZN(new_n20432_));
  NOR2_X1    g20176(.A1(new_n20432_), .A2(new_n20397_), .ZN(new_n20433_));
  INV_X1     g20177(.I(new_n20433_), .ZN(new_n20434_));
  NAND2_X1   g20178(.A1(new_n20432_), .A2(new_n20397_), .ZN(new_n20435_));
  NAND2_X1   g20179(.A1(new_n20434_), .A2(new_n20435_), .ZN(new_n20436_));
  XOR2_X1    g20180(.A1(new_n20436_), .A2(new_n20392_), .Z(new_n20437_));
  NOR2_X1    g20181(.A1(new_n20437_), .A2(new_n20390_), .ZN(new_n20438_));
  INV_X1     g20182(.I(new_n20438_), .ZN(new_n20439_));
  NAND2_X1   g20183(.A1(new_n20437_), .A2(new_n20390_), .ZN(new_n20440_));
  NAND2_X1   g20184(.A1(new_n20439_), .A2(new_n20440_), .ZN(new_n20441_));
  XOR2_X1    g20185(.A1(new_n20441_), .A2(new_n20386_), .Z(new_n20442_));
  NOR2_X1    g20186(.A1(new_n20442_), .A2(new_n20384_), .ZN(new_n20443_));
  INV_X1     g20187(.I(new_n20443_), .ZN(new_n20444_));
  NAND2_X1   g20188(.A1(new_n20442_), .A2(new_n20384_), .ZN(new_n20445_));
  NAND2_X1   g20189(.A1(new_n20444_), .A2(new_n20445_), .ZN(new_n20446_));
  XOR2_X1    g20190(.A1(new_n20446_), .A2(new_n20382_), .Z(new_n20447_));
  INV_X1     g20191(.I(new_n20366_), .ZN(new_n20448_));
  INV_X1     g20192(.I(new_n20369_), .ZN(new_n20449_));
  XOR2_X1    g20193(.A1(new_n20302_), .A2(new_n6567_), .Z(new_n20450_));
  AOI21_X1   g20194(.A1(new_n20366_), .A2(new_n20449_), .B(new_n20450_), .ZN(new_n20451_));
  AOI21_X1   g20195(.A1(new_n20448_), .A2(new_n20369_), .B(new_n20451_), .ZN(new_n20452_));
  INV_X1     g20196(.I(new_n20452_), .ZN(new_n20453_));
  NOR2_X1    g20197(.A1(new_n20447_), .A2(new_n20453_), .ZN(new_n20454_));
  INV_X1     g20198(.I(new_n20454_), .ZN(new_n20455_));
  NAND2_X1   g20199(.A1(new_n20447_), .A2(new_n20453_), .ZN(new_n20456_));
  AND2_X2    g20200(.A1(new_n20455_), .A2(new_n20456_), .Z(new_n20457_));
  INV_X1     g20201(.I(new_n20457_), .ZN(new_n20458_));
  NOR3_X1    g20202(.A1(new_n20378_), .A2(new_n20372_), .A3(new_n20458_), .ZN(new_n20459_));
  AOI21_X1   g20203(.A1(new_n20293_), .A2(new_n20284_), .B(new_n20282_), .ZN(new_n20460_));
  OAI21_X1   g20204(.A1(new_n20460_), .A2(new_n20294_), .B(new_n20374_), .ZN(new_n20461_));
  AOI21_X1   g20205(.A1(new_n20461_), .A2(new_n20373_), .B(new_n20457_), .ZN(new_n20462_));
  NOR2_X1    g20206(.A1(new_n20462_), .A2(new_n20459_), .ZN(\f[108] ));
  OAI22_X1   g20207(.A1(new_n9488_), .A2(new_n12796_), .B1(new_n12800_), .B2(new_n8588_), .ZN(new_n20464_));
  AOI21_X1   g20208(.A1(new_n13973_), .A2(new_n7414_), .B(new_n20464_), .ZN(new_n20465_));
  XOR2_X1    g20209(.A1(new_n20465_), .A2(new_n7410_), .Z(new_n20466_));
  INV_X1     g20210(.I(new_n20466_), .ZN(new_n20467_));
  OAI21_X1   g20211(.A1(new_n20386_), .A2(new_n20438_), .B(new_n20440_), .ZN(new_n20468_));
  OAI22_X1   g20212(.A1(new_n9461_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n9462_), .ZN(new_n20469_));
  AOI21_X1   g20213(.A1(\b[59] ), .A2(new_n8575_), .B(new_n20469_), .ZN(new_n20470_));
  OAI21_X1   g20214(.A1(new_n13110_), .A2(new_n9460_), .B(new_n20470_), .ZN(new_n20471_));
  XOR2_X1    g20215(.A1(new_n20471_), .A2(new_n8248_), .Z(new_n20472_));
  OAI21_X1   g20216(.A1(new_n20392_), .A2(new_n20433_), .B(new_n20435_), .ZN(new_n20473_));
  AOI22_X1   g20217(.A1(new_n9125_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n9123_), .ZN(new_n20474_));
  OAI21_X1   g20218(.A1(new_n10308_), .A2(new_n9470_), .B(new_n20474_), .ZN(new_n20475_));
  AOI21_X1   g20219(.A1(new_n12164_), .A2(new_n9129_), .B(new_n20475_), .ZN(new_n20476_));
  XOR2_X1    g20220(.A1(new_n20476_), .A2(new_n9133_), .Z(new_n20477_));
  OAI21_X1   g20221(.A1(new_n20398_), .A2(new_n20428_), .B(new_n20429_), .ZN(new_n20478_));
  INV_X1     g20222(.I(new_n20478_), .ZN(new_n20479_));
  AOI21_X1   g20223(.A1(new_n20404_), .A2(new_n20424_), .B(new_n20423_), .ZN(new_n20480_));
  AOI22_X1   g20224(.A1(new_n10981_), .A2(\b[52] ), .B1(new_n10979_), .B2(\b[51] ), .ZN(new_n20481_));
  OAI21_X1   g20225(.A1(new_n8500_), .A2(new_n11306_), .B(new_n20481_), .ZN(new_n20482_));
  AOI21_X1   g20226(.A1(new_n9987_), .A2(new_n10984_), .B(new_n20482_), .ZN(new_n20483_));
  XOR2_X1    g20227(.A1(new_n20483_), .A2(new_n10989_), .Z(new_n20484_));
  AOI21_X1   g20228(.A1(new_n20406_), .A2(new_n20415_), .B(new_n20414_), .ZN(new_n20485_));
  INV_X1     g20229(.I(new_n20485_), .ZN(new_n20486_));
  OAI22_X1   g20230(.A1(new_n13224_), .A2(new_n8168_), .B1(new_n8127_), .B2(new_n11923_), .ZN(new_n20487_));
  AOI21_X1   g20231(.A1(\b[47] ), .A2(new_n13223_), .B(new_n20487_), .ZN(new_n20488_));
  OAI21_X1   g20232(.A1(new_n9050_), .A2(new_n11930_), .B(new_n20488_), .ZN(new_n20489_));
  XOR2_X1    g20233(.A1(new_n20489_), .A2(new_n12312_), .Z(new_n20490_));
  NOR2_X1    g20234(.A1(new_n20411_), .A2(\a[44] ), .ZN(new_n20491_));
  NOR2_X1    g20235(.A1(new_n20491_), .A2(new_n20327_), .ZN(new_n20492_));
  AOI21_X1   g20236(.A1(\a[44] ), .A2(new_n20411_), .B(new_n20492_), .ZN(new_n20493_));
  AOI22_X1   g20237(.A1(new_n12922_), .A2(\b[46] ), .B1(\b[45] ), .B2(new_n12923_), .ZN(new_n20494_));
  NAND2_X1   g20238(.A1(new_n20493_), .A2(new_n20494_), .ZN(new_n20495_));
  OR2_X2     g20239(.A1(new_n20493_), .A2(new_n20494_), .Z(new_n20496_));
  NAND2_X1   g20240(.A1(new_n20496_), .A2(new_n20495_), .ZN(new_n20497_));
  XNOR2_X1   g20241(.A1(new_n20490_), .A2(new_n20497_), .ZN(new_n20498_));
  NOR2_X1    g20242(.A1(new_n20498_), .A2(new_n20486_), .ZN(new_n20499_));
  INV_X1     g20243(.I(new_n20499_), .ZN(new_n20500_));
  NAND2_X1   g20244(.A1(new_n20498_), .A2(new_n20486_), .ZN(new_n20501_));
  NAND2_X1   g20245(.A1(new_n20500_), .A2(new_n20501_), .ZN(new_n20502_));
  XOR2_X1    g20246(.A1(new_n20502_), .A2(new_n20484_), .Z(new_n20503_));
  INV_X1     g20247(.I(new_n20503_), .ZN(new_n20504_));
  AOI22_X1   g20248(.A1(new_n10064_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n10062_), .ZN(new_n20505_));
  OAI21_X1   g20249(.A1(new_n9376_), .A2(new_n10399_), .B(new_n20505_), .ZN(new_n20506_));
  AOI21_X1   g20250(.A1(new_n9979_), .A2(new_n10068_), .B(new_n20506_), .ZN(new_n20507_));
  XOR2_X1    g20251(.A1(new_n20507_), .A2(new_n10057_), .Z(new_n20508_));
  NOR2_X1    g20252(.A1(new_n20504_), .A2(new_n20508_), .ZN(new_n20509_));
  NAND2_X1   g20253(.A1(new_n20504_), .A2(new_n20508_), .ZN(new_n20510_));
  INV_X1     g20254(.I(new_n20510_), .ZN(new_n20511_));
  NOR2_X1    g20255(.A1(new_n20511_), .A2(new_n20509_), .ZN(new_n20512_));
  XOR2_X1    g20256(.A1(new_n20512_), .A2(new_n20480_), .Z(new_n20513_));
  NOR2_X1    g20257(.A1(new_n20513_), .A2(new_n20479_), .ZN(new_n20514_));
  INV_X1     g20258(.I(new_n20514_), .ZN(new_n20515_));
  NAND2_X1   g20259(.A1(new_n20513_), .A2(new_n20479_), .ZN(new_n20516_));
  NAND2_X1   g20260(.A1(new_n20515_), .A2(new_n20516_), .ZN(new_n20517_));
  XOR2_X1    g20261(.A1(new_n20517_), .A2(new_n20477_), .Z(new_n20518_));
  OR2_X2     g20262(.A1(new_n20518_), .A2(new_n20473_), .Z(new_n20519_));
  NAND2_X1   g20263(.A1(new_n20518_), .A2(new_n20473_), .ZN(new_n20520_));
  NAND2_X1   g20264(.A1(new_n20519_), .A2(new_n20520_), .ZN(new_n20521_));
  XNOR2_X1   g20265(.A1(new_n20521_), .A2(new_n20472_), .ZN(new_n20522_));
  NAND2_X1   g20266(.A1(new_n20522_), .A2(new_n20468_), .ZN(new_n20523_));
  NOR2_X1    g20267(.A1(new_n20522_), .A2(new_n20468_), .ZN(new_n20524_));
  INV_X1     g20268(.I(new_n20524_), .ZN(new_n20525_));
  NAND2_X1   g20269(.A1(new_n20525_), .A2(new_n20523_), .ZN(new_n20526_));
  XOR2_X1    g20270(.A1(new_n20526_), .A2(new_n20467_), .Z(new_n20527_));
  INV_X1     g20271(.I(new_n20527_), .ZN(new_n20528_));
  OAI21_X1   g20272(.A1(new_n20382_), .A2(new_n20443_), .B(new_n20445_), .ZN(new_n20529_));
  INV_X1     g20273(.I(new_n20529_), .ZN(new_n20530_));
  OAI21_X1   g20274(.A1(new_n20459_), .A2(new_n20454_), .B(new_n20530_), .ZN(new_n20531_));
  NAND3_X1   g20275(.A1(new_n20461_), .A2(new_n20373_), .A3(new_n20457_), .ZN(new_n20532_));
  NAND3_X1   g20276(.A1(new_n20532_), .A2(new_n20455_), .A3(new_n20529_), .ZN(new_n20533_));
  NAND2_X1   g20277(.A1(new_n20533_), .A2(new_n20531_), .ZN(new_n20534_));
  XOR2_X1    g20278(.A1(new_n20534_), .A2(new_n20528_), .Z(\f[109] ));
  NOR3_X1    g20279(.A1(new_n20459_), .A2(new_n20454_), .A3(new_n20530_), .ZN(new_n20536_));
  AOI21_X1   g20280(.A1(new_n20528_), .A2(new_n20531_), .B(new_n20536_), .ZN(new_n20537_));
  AOI22_X1   g20281(.A1(new_n8241_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n8246_), .ZN(new_n20538_));
  OAI21_X1   g20282(.A1(new_n12147_), .A2(new_n9114_), .B(new_n20538_), .ZN(new_n20539_));
  AOI21_X1   g20283(.A1(new_n13444_), .A2(new_n8252_), .B(new_n20539_), .ZN(new_n20540_));
  XOR2_X1    g20284(.A1(new_n20540_), .A2(\a[50] ), .Z(new_n20541_));
  AOI22_X1   g20285(.A1(new_n10064_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n10062_), .ZN(new_n20542_));
  OAI21_X1   g20286(.A1(new_n9942_), .A2(new_n10399_), .B(new_n20542_), .ZN(new_n20543_));
  AOI21_X1   g20287(.A1(new_n10318_), .A2(new_n10068_), .B(new_n20543_), .ZN(new_n20544_));
  XOR2_X1    g20288(.A1(new_n20544_), .A2(new_n10057_), .Z(new_n20545_));
  OAI21_X1   g20289(.A1(new_n20484_), .A2(new_n20499_), .B(new_n20501_), .ZN(new_n20546_));
  OAI22_X1   g20290(.A1(new_n12306_), .A2(new_n9376_), .B1(new_n12305_), .B2(new_n9032_), .ZN(new_n20547_));
  AOI21_X1   g20291(.A1(\b[51] ), .A2(new_n12304_), .B(new_n20547_), .ZN(new_n20548_));
  OAI21_X1   g20292(.A1(new_n9385_), .A2(new_n10985_), .B(new_n20548_), .ZN(new_n20549_));
  XOR2_X1    g20293(.A1(new_n20549_), .A2(new_n10989_), .Z(new_n20550_));
  AOI22_X1   g20294(.A1(new_n11926_), .A2(\b[50] ), .B1(new_n11924_), .B2(\b[49] ), .ZN(new_n20551_));
  OAI21_X1   g20295(.A1(new_n8127_), .A2(new_n12317_), .B(new_n20551_), .ZN(new_n20552_));
  AOI21_X1   g20296(.A1(new_n9684_), .A2(new_n11929_), .B(new_n20552_), .ZN(new_n20553_));
  XOR2_X1    g20297(.A1(new_n20553_), .A2(new_n12312_), .Z(new_n20554_));
  NAND2_X1   g20298(.A1(new_n20490_), .A2(new_n20495_), .ZN(new_n20555_));
  NAND2_X1   g20299(.A1(new_n20555_), .A2(new_n20496_), .ZN(new_n20556_));
  AOI22_X1   g20300(.A1(new_n12922_), .A2(\b[47] ), .B1(\b[46] ), .B2(new_n12923_), .ZN(new_n20557_));
  INV_X1     g20301(.I(new_n20557_), .ZN(new_n20558_));
  NOR2_X1    g20302(.A1(new_n20558_), .A2(new_n20494_), .ZN(new_n20559_));
  NAND2_X1   g20303(.A1(new_n20558_), .A2(new_n20494_), .ZN(new_n20560_));
  INV_X1     g20304(.I(new_n20560_), .ZN(new_n20561_));
  NOR2_X1    g20305(.A1(new_n20561_), .A2(new_n20559_), .ZN(new_n20562_));
  XNOR2_X1   g20306(.A1(new_n20556_), .A2(new_n20562_), .ZN(new_n20563_));
  NOR2_X1    g20307(.A1(new_n20563_), .A2(new_n20554_), .ZN(new_n20564_));
  INV_X1     g20308(.I(new_n20564_), .ZN(new_n20565_));
  NAND2_X1   g20309(.A1(new_n20563_), .A2(new_n20554_), .ZN(new_n20566_));
  NAND2_X1   g20310(.A1(new_n20565_), .A2(new_n20566_), .ZN(new_n20567_));
  XNOR2_X1   g20311(.A1(new_n20567_), .A2(new_n20550_), .ZN(new_n20568_));
  NOR2_X1    g20312(.A1(new_n20568_), .A2(new_n20546_), .ZN(new_n20569_));
  INV_X1     g20313(.I(new_n20569_), .ZN(new_n20570_));
  NAND2_X1   g20314(.A1(new_n20568_), .A2(new_n20546_), .ZN(new_n20571_));
  NAND2_X1   g20315(.A1(new_n20570_), .A2(new_n20571_), .ZN(new_n20572_));
  XOR2_X1    g20316(.A1(new_n20572_), .A2(new_n20545_), .Z(new_n20573_));
  OAI22_X1   g20317(.A1(new_n10390_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n10389_), .ZN(new_n20574_));
  AOI21_X1   g20318(.A1(\b[57] ), .A2(new_n9471_), .B(new_n20574_), .ZN(new_n20575_));
  OAI21_X1   g20319(.A1(new_n12203_), .A2(new_n10388_), .B(new_n20575_), .ZN(new_n20576_));
  XOR2_X1    g20320(.A1(new_n20576_), .A2(\a[53] ), .Z(new_n20577_));
  NOR2_X1    g20321(.A1(new_n20511_), .A2(new_n20480_), .ZN(new_n20578_));
  NOR2_X1    g20322(.A1(new_n20578_), .A2(new_n20509_), .ZN(new_n20579_));
  NOR2_X1    g20323(.A1(new_n20579_), .A2(new_n20577_), .ZN(new_n20580_));
  INV_X1     g20324(.I(new_n20580_), .ZN(new_n20581_));
  NAND2_X1   g20325(.A1(new_n20579_), .A2(new_n20577_), .ZN(new_n20582_));
  NAND2_X1   g20326(.A1(new_n20581_), .A2(new_n20582_), .ZN(new_n20583_));
  XOR2_X1    g20327(.A1(new_n20573_), .A2(new_n20583_), .Z(new_n20584_));
  INV_X1     g20328(.I(new_n20477_), .ZN(new_n20585_));
  AOI21_X1   g20329(.A1(new_n20585_), .A2(new_n20516_), .B(new_n20514_), .ZN(new_n20586_));
  OR2_X2     g20330(.A1(new_n20584_), .A2(new_n20586_), .Z(new_n20587_));
  NAND2_X1   g20331(.A1(new_n20584_), .A2(new_n20586_), .ZN(new_n20588_));
  NAND2_X1   g20332(.A1(new_n20587_), .A2(new_n20588_), .ZN(new_n20589_));
  XOR2_X1    g20333(.A1(new_n20589_), .A2(new_n20541_), .Z(new_n20590_));
  AOI22_X1   g20334(.A1(new_n13460_), .A2(new_n7414_), .B1(\b[63] ), .B2(new_n7719_), .ZN(new_n20591_));
  XOR2_X1    g20335(.A1(new_n20590_), .A2(new_n20591_), .Z(new_n20592_));
  NAND2_X1   g20336(.A1(new_n20519_), .A2(new_n20472_), .ZN(new_n20593_));
  NAND2_X1   g20337(.A1(new_n20593_), .A2(new_n20520_), .ZN(new_n20594_));
  XOR2_X1    g20338(.A1(new_n20594_), .A2(new_n7410_), .Z(new_n20595_));
  XNOR2_X1   g20339(.A1(new_n20592_), .A2(new_n20595_), .ZN(new_n20596_));
  OAI21_X1   g20340(.A1(new_n20466_), .A2(new_n20524_), .B(new_n20523_), .ZN(new_n20597_));
  INV_X1     g20341(.I(new_n20597_), .ZN(new_n20598_));
  NOR2_X1    g20342(.A1(new_n20596_), .A2(new_n20598_), .ZN(new_n20599_));
  NAND2_X1   g20343(.A1(new_n20596_), .A2(new_n20598_), .ZN(new_n20600_));
  INV_X1     g20344(.I(new_n20600_), .ZN(new_n20601_));
  NOR2_X1    g20345(.A1(new_n20601_), .A2(new_n20599_), .ZN(new_n20602_));
  XOR2_X1    g20346(.A1(new_n20537_), .A2(new_n20602_), .Z(\f[110] ));
  INV_X1     g20347(.I(new_n20599_), .ZN(new_n20604_));
  OAI21_X1   g20348(.A1(new_n20537_), .A2(new_n20601_), .B(new_n20604_), .ZN(new_n20605_));
  AOI22_X1   g20349(.A1(new_n8241_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n8246_), .ZN(new_n20606_));
  OAI21_X1   g20350(.A1(new_n12148_), .A2(new_n9114_), .B(new_n20606_), .ZN(new_n20607_));
  AOI21_X1   g20351(.A1(new_n12811_), .A2(new_n8252_), .B(new_n20607_), .ZN(new_n20608_));
  XOR2_X1    g20352(.A1(new_n20608_), .A2(new_n8248_), .Z(new_n20609_));
  NAND2_X1   g20353(.A1(new_n20588_), .A2(new_n20541_), .ZN(new_n20610_));
  NAND2_X1   g20354(.A1(new_n20610_), .A2(new_n20587_), .ZN(new_n20611_));
  AOI21_X1   g20355(.A1(new_n20573_), .A2(new_n20582_), .B(new_n20580_), .ZN(new_n20612_));
  AOI22_X1   g20356(.A1(new_n9125_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n9123_), .ZN(new_n20613_));
  OAI21_X1   g20357(.A1(new_n11195_), .A2(new_n9470_), .B(new_n20613_), .ZN(new_n20614_));
  AOI21_X1   g20358(.A1(new_n11836_), .A2(new_n9129_), .B(new_n20614_), .ZN(new_n20615_));
  XOR2_X1    g20359(.A1(new_n20615_), .A2(new_n9133_), .Z(new_n20616_));
  OAI21_X1   g20360(.A1(new_n20545_), .A2(new_n20569_), .B(new_n20571_), .ZN(new_n20617_));
  INV_X1     g20361(.I(new_n20617_), .ZN(new_n20618_));
  AOI22_X1   g20362(.A1(new_n10064_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n10062_), .ZN(new_n20619_));
  OAI21_X1   g20363(.A1(new_n9972_), .A2(new_n10399_), .B(new_n20619_), .ZN(new_n20620_));
  AOI21_X1   g20364(.A1(new_n10631_), .A2(new_n10068_), .B(new_n20620_), .ZN(new_n20621_));
  XOR2_X1    g20365(.A1(new_n20621_), .A2(new_n10057_), .Z(new_n20622_));
  INV_X1     g20366(.I(new_n20622_), .ZN(new_n20623_));
  AOI21_X1   g20367(.A1(new_n20550_), .A2(new_n20566_), .B(new_n20564_), .ZN(new_n20624_));
  INV_X1     g20368(.I(new_n20624_), .ZN(new_n20625_));
  AOI22_X1   g20369(.A1(new_n10981_), .A2(\b[54] ), .B1(new_n10979_), .B2(\b[53] ), .ZN(new_n20626_));
  OAI21_X1   g20370(.A1(new_n9032_), .A2(new_n11306_), .B(new_n20626_), .ZN(new_n20627_));
  AOI21_X1   g20371(.A1(new_n10884_), .A2(new_n10984_), .B(new_n20627_), .ZN(new_n20628_));
  XOR2_X1    g20372(.A1(new_n20628_), .A2(new_n10989_), .Z(new_n20629_));
  INV_X1     g20373(.I(new_n20559_), .ZN(new_n20630_));
  AOI21_X1   g20374(.A1(new_n20556_), .A2(new_n20630_), .B(new_n20561_), .ZN(new_n20631_));
  AOI22_X1   g20375(.A1(new_n11926_), .A2(\b[51] ), .B1(new_n11924_), .B2(\b[50] ), .ZN(new_n20632_));
  OAI21_X1   g20376(.A1(new_n8168_), .A2(new_n12317_), .B(new_n20632_), .ZN(new_n20633_));
  AOI21_X1   g20377(.A1(new_n8783_), .A2(new_n11929_), .B(new_n20633_), .ZN(new_n20634_));
  XOR2_X1    g20378(.A1(new_n20634_), .A2(new_n12312_), .Z(new_n20635_));
  INV_X1     g20379(.I(new_n20635_), .ZN(new_n20636_));
  AOI22_X1   g20380(.A1(new_n12922_), .A2(\b[48] ), .B1(\b[47] ), .B2(new_n12923_), .ZN(new_n20637_));
  INV_X1     g20381(.I(new_n20637_), .ZN(new_n20638_));
  NOR2_X1    g20382(.A1(new_n20638_), .A2(new_n7410_), .ZN(new_n20639_));
  NOR2_X1    g20383(.A1(new_n20637_), .A2(\a[47] ), .ZN(new_n20640_));
  NOR2_X1    g20384(.A1(new_n20639_), .A2(new_n20640_), .ZN(new_n20641_));
  XOR2_X1    g20385(.A1(new_n20641_), .A2(new_n20557_), .Z(new_n20642_));
  NOR2_X1    g20386(.A1(new_n20636_), .A2(new_n20642_), .ZN(new_n20643_));
  NAND2_X1   g20387(.A1(new_n20636_), .A2(new_n20642_), .ZN(new_n20644_));
  INV_X1     g20388(.I(new_n20644_), .ZN(new_n20645_));
  NOR2_X1    g20389(.A1(new_n20645_), .A2(new_n20643_), .ZN(new_n20646_));
  XOR2_X1    g20390(.A1(new_n20646_), .A2(new_n20631_), .Z(new_n20647_));
  NOR2_X1    g20391(.A1(new_n20647_), .A2(new_n20629_), .ZN(new_n20648_));
  NAND2_X1   g20392(.A1(new_n20647_), .A2(new_n20629_), .ZN(new_n20649_));
  INV_X1     g20393(.I(new_n20649_), .ZN(new_n20650_));
  NOR2_X1    g20394(.A1(new_n20650_), .A2(new_n20648_), .ZN(new_n20651_));
  XOR2_X1    g20395(.A1(new_n20651_), .A2(new_n20625_), .Z(new_n20652_));
  NOR2_X1    g20396(.A1(new_n20652_), .A2(new_n20623_), .ZN(new_n20653_));
  NAND2_X1   g20397(.A1(new_n20652_), .A2(new_n20623_), .ZN(new_n20654_));
  INV_X1     g20398(.I(new_n20654_), .ZN(new_n20655_));
  NOR2_X1    g20399(.A1(new_n20655_), .A2(new_n20653_), .ZN(new_n20656_));
  XOR2_X1    g20400(.A1(new_n20656_), .A2(new_n20618_), .Z(new_n20657_));
  NAND2_X1   g20401(.A1(new_n20657_), .A2(new_n20616_), .ZN(new_n20658_));
  NOR2_X1    g20402(.A1(new_n20657_), .A2(new_n20616_), .ZN(new_n20659_));
  INV_X1     g20403(.I(new_n20659_), .ZN(new_n20660_));
  NAND2_X1   g20404(.A1(new_n20660_), .A2(new_n20658_), .ZN(new_n20661_));
  XOR2_X1    g20405(.A1(new_n20661_), .A2(new_n20612_), .Z(new_n20662_));
  NOR2_X1    g20406(.A1(new_n20662_), .A2(new_n20611_), .ZN(new_n20663_));
  INV_X1     g20407(.I(new_n20663_), .ZN(new_n20664_));
  NAND2_X1   g20408(.A1(new_n20662_), .A2(new_n20611_), .ZN(new_n20665_));
  NAND2_X1   g20409(.A1(new_n20664_), .A2(new_n20665_), .ZN(new_n20666_));
  XOR2_X1    g20410(.A1(new_n20666_), .A2(new_n20609_), .Z(new_n20667_));
  INV_X1     g20411(.I(new_n20590_), .ZN(new_n20668_));
  INV_X1     g20412(.I(new_n20594_), .ZN(new_n20669_));
  XOR2_X1    g20413(.A1(new_n20591_), .A2(new_n7410_), .Z(new_n20670_));
  AOI21_X1   g20414(.A1(new_n20669_), .A2(new_n20590_), .B(new_n20670_), .ZN(new_n20671_));
  AOI21_X1   g20415(.A1(new_n20668_), .A2(new_n20594_), .B(new_n20671_), .ZN(new_n20672_));
  INV_X1     g20416(.I(new_n20672_), .ZN(new_n20673_));
  NOR2_X1    g20417(.A1(new_n20667_), .A2(new_n20673_), .ZN(new_n20674_));
  INV_X1     g20418(.I(new_n20674_), .ZN(new_n20675_));
  NAND2_X1   g20419(.A1(new_n20667_), .A2(new_n20673_), .ZN(new_n20676_));
  AND2_X2    g20420(.A1(new_n20675_), .A2(new_n20676_), .Z(new_n20677_));
  INV_X1     g20421(.I(new_n20677_), .ZN(new_n20678_));
  XOR2_X1    g20422(.A1(new_n20605_), .A2(new_n20678_), .Z(\f[111] ));
  OAI22_X1   g20423(.A1(new_n9114_), .A2(new_n12796_), .B1(new_n12800_), .B2(new_n9462_), .ZN(new_n20680_));
  AOI21_X1   g20424(.A1(new_n13973_), .A2(new_n8252_), .B(new_n20680_), .ZN(new_n20681_));
  XOR2_X1    g20425(.A1(new_n20681_), .A2(new_n8248_), .Z(new_n20682_));
  INV_X1     g20426(.I(new_n20682_), .ZN(new_n20683_));
  INV_X1     g20427(.I(new_n20612_), .ZN(new_n20684_));
  AOI21_X1   g20428(.A1(new_n20684_), .A2(new_n20658_), .B(new_n20659_), .ZN(new_n20685_));
  INV_X1     g20429(.I(new_n20685_), .ZN(new_n20686_));
  OAI22_X1   g20430(.A1(new_n10390_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n10389_), .ZN(new_n20687_));
  AOI21_X1   g20431(.A1(\b[59] ), .A2(new_n9471_), .B(new_n20687_), .ZN(new_n20688_));
  OAI21_X1   g20432(.A1(new_n13110_), .A2(new_n10388_), .B(new_n20688_), .ZN(new_n20689_));
  XOR2_X1    g20433(.A1(new_n20689_), .A2(new_n9133_), .Z(new_n20690_));
  OAI21_X1   g20434(.A1(new_n20618_), .A2(new_n20653_), .B(new_n20654_), .ZN(new_n20691_));
  AOI22_X1   g20435(.A1(new_n10064_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n10062_), .ZN(new_n20692_));
  OAI21_X1   g20436(.A1(new_n10308_), .A2(new_n10399_), .B(new_n20692_), .ZN(new_n20693_));
  AOI21_X1   g20437(.A1(new_n12164_), .A2(new_n10068_), .B(new_n20693_), .ZN(new_n20694_));
  XOR2_X1    g20438(.A1(new_n20694_), .A2(new_n10057_), .Z(new_n20695_));
  AOI21_X1   g20439(.A1(new_n20625_), .A2(new_n20649_), .B(new_n20648_), .ZN(new_n20696_));
  INV_X1     g20440(.I(new_n20696_), .ZN(new_n20697_));
  AOI22_X1   g20441(.A1(new_n10981_), .A2(\b[55] ), .B1(new_n10979_), .B2(\b[54] ), .ZN(new_n20698_));
  OAI21_X1   g20442(.A1(new_n9376_), .A2(new_n11306_), .B(new_n20698_), .ZN(new_n20699_));
  AOI21_X1   g20443(.A1(new_n9979_), .A2(new_n10984_), .B(new_n20699_), .ZN(new_n20700_));
  XOR2_X1    g20444(.A1(new_n20700_), .A2(\a[59] ), .Z(new_n20701_));
  OAI21_X1   g20445(.A1(new_n20631_), .A2(new_n20643_), .B(new_n20644_), .ZN(new_n20702_));
  INV_X1     g20446(.I(new_n20702_), .ZN(new_n20703_));
  AOI22_X1   g20447(.A1(new_n11926_), .A2(\b[52] ), .B1(new_n11924_), .B2(\b[51] ), .ZN(new_n20704_));
  OAI21_X1   g20448(.A1(new_n8500_), .A2(new_n12317_), .B(new_n20704_), .ZN(new_n20705_));
  AOI21_X1   g20449(.A1(new_n9987_), .A2(new_n11929_), .B(new_n20705_), .ZN(new_n20706_));
  XOR2_X1    g20450(.A1(new_n20706_), .A2(\a[62] ), .Z(new_n20707_));
  NOR2_X1    g20451(.A1(new_n20640_), .A2(new_n20558_), .ZN(new_n20708_));
  NOR2_X1    g20452(.A1(new_n20708_), .A2(new_n20639_), .ZN(new_n20709_));
  AOI22_X1   g20453(.A1(new_n12922_), .A2(\b[49] ), .B1(\b[48] ), .B2(new_n12923_), .ZN(new_n20710_));
  NAND2_X1   g20454(.A1(new_n20709_), .A2(new_n20710_), .ZN(new_n20711_));
  NOR2_X1    g20455(.A1(new_n20709_), .A2(new_n20710_), .ZN(new_n20712_));
  INV_X1     g20456(.I(new_n20712_), .ZN(new_n20713_));
  NAND2_X1   g20457(.A1(new_n20713_), .A2(new_n20711_), .ZN(new_n20714_));
  XNOR2_X1   g20458(.A1(new_n20707_), .A2(new_n20714_), .ZN(new_n20715_));
  INV_X1     g20459(.I(new_n20715_), .ZN(new_n20716_));
  NAND2_X1   g20460(.A1(new_n20703_), .A2(new_n20716_), .ZN(new_n20717_));
  NOR2_X1    g20461(.A1(new_n20703_), .A2(new_n20716_), .ZN(new_n20718_));
  INV_X1     g20462(.I(new_n20718_), .ZN(new_n20719_));
  NAND2_X1   g20463(.A1(new_n20719_), .A2(new_n20717_), .ZN(new_n20720_));
  XNOR2_X1   g20464(.A1(new_n20720_), .A2(new_n20701_), .ZN(new_n20721_));
  NOR2_X1    g20465(.A1(new_n20721_), .A2(new_n20697_), .ZN(new_n20722_));
  INV_X1     g20466(.I(new_n20722_), .ZN(new_n20723_));
  NAND2_X1   g20467(.A1(new_n20721_), .A2(new_n20697_), .ZN(new_n20724_));
  NAND2_X1   g20468(.A1(new_n20723_), .A2(new_n20724_), .ZN(new_n20725_));
  XOR2_X1    g20469(.A1(new_n20725_), .A2(new_n20695_), .Z(new_n20726_));
  OR2_X2     g20470(.A1(new_n20726_), .A2(new_n20691_), .Z(new_n20727_));
  NAND2_X1   g20471(.A1(new_n20726_), .A2(new_n20691_), .ZN(new_n20728_));
  NAND2_X1   g20472(.A1(new_n20727_), .A2(new_n20728_), .ZN(new_n20729_));
  XNOR2_X1   g20473(.A1(new_n20729_), .A2(new_n20690_), .ZN(new_n20730_));
  NOR2_X1    g20474(.A1(new_n20730_), .A2(new_n20686_), .ZN(new_n20731_));
  INV_X1     g20475(.I(new_n20731_), .ZN(new_n20732_));
  NAND2_X1   g20476(.A1(new_n20730_), .A2(new_n20686_), .ZN(new_n20733_));
  NAND2_X1   g20477(.A1(new_n20732_), .A2(new_n20733_), .ZN(new_n20734_));
  XOR2_X1    g20478(.A1(new_n20734_), .A2(new_n20683_), .Z(new_n20735_));
  OAI21_X1   g20479(.A1(new_n20609_), .A2(new_n20663_), .B(new_n20665_), .ZN(new_n20736_));
  AOI21_X1   g20480(.A1(new_n20532_), .A2(new_n20455_), .B(new_n20529_), .ZN(new_n20737_));
  OAI21_X1   g20481(.A1(new_n20527_), .A2(new_n20737_), .B(new_n20533_), .ZN(new_n20738_));
  AOI21_X1   g20482(.A1(new_n20738_), .A2(new_n20600_), .B(new_n20599_), .ZN(new_n20739_));
  AOI21_X1   g20483(.A1(new_n20739_), .A2(new_n20677_), .B(new_n20674_), .ZN(new_n20740_));
  NOR2_X1    g20484(.A1(new_n20740_), .A2(new_n20736_), .ZN(new_n20741_));
  INV_X1     g20485(.I(new_n20736_), .ZN(new_n20742_));
  OAI21_X1   g20486(.A1(new_n20605_), .A2(new_n20678_), .B(new_n20675_), .ZN(new_n20743_));
  NOR2_X1    g20487(.A1(new_n20743_), .A2(new_n20742_), .ZN(new_n20744_));
  NOR2_X1    g20488(.A1(new_n20741_), .A2(new_n20744_), .ZN(new_n20745_));
  XOR2_X1    g20489(.A1(new_n20745_), .A2(new_n20735_), .Z(\f[112] ));
  AOI21_X1   g20490(.A1(new_n20743_), .A2(new_n20742_), .B(new_n20735_), .ZN(new_n20747_));
  NOR2_X1    g20491(.A1(new_n20747_), .A2(new_n20744_), .ZN(new_n20748_));
  AOI22_X1   g20492(.A1(new_n9125_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n9123_), .ZN(new_n20749_));
  OAI21_X1   g20493(.A1(new_n12147_), .A2(new_n9470_), .B(new_n20749_), .ZN(new_n20750_));
  AOI21_X1   g20494(.A1(new_n13444_), .A2(new_n9129_), .B(new_n20750_), .ZN(new_n20751_));
  XOR2_X1    g20495(.A1(new_n20751_), .A2(\a[53] ), .Z(new_n20752_));
  AOI22_X1   g20496(.A1(new_n10981_), .A2(\b[56] ), .B1(new_n10979_), .B2(\b[55] ), .ZN(new_n20753_));
  OAI21_X1   g20497(.A1(new_n9942_), .A2(new_n11306_), .B(new_n20753_), .ZN(new_n20754_));
  AOI21_X1   g20498(.A1(new_n10318_), .A2(new_n10984_), .B(new_n20754_), .ZN(new_n20755_));
  XOR2_X1    g20499(.A1(new_n20755_), .A2(new_n10989_), .Z(new_n20756_));
  AOI21_X1   g20500(.A1(new_n20707_), .A2(new_n20711_), .B(new_n20712_), .ZN(new_n20757_));
  OAI22_X1   g20501(.A1(new_n13224_), .A2(new_n9376_), .B1(new_n9032_), .B2(new_n11923_), .ZN(new_n20758_));
  AOI21_X1   g20502(.A1(\b[51] ), .A2(new_n13223_), .B(new_n20758_), .ZN(new_n20759_));
  OAI21_X1   g20503(.A1(new_n9385_), .A2(new_n11930_), .B(new_n20759_), .ZN(new_n20760_));
  XOR2_X1    g20504(.A1(new_n20760_), .A2(\a[62] ), .Z(new_n20761_));
  AOI22_X1   g20505(.A1(new_n12922_), .A2(\b[50] ), .B1(\b[49] ), .B2(new_n12923_), .ZN(new_n20762_));
  INV_X1     g20506(.I(new_n20762_), .ZN(new_n20763_));
  NOR2_X1    g20507(.A1(new_n20763_), .A2(new_n20710_), .ZN(new_n20764_));
  INV_X1     g20508(.I(new_n20710_), .ZN(new_n20765_));
  NOR2_X1    g20509(.A1(new_n20765_), .A2(new_n20762_), .ZN(new_n20766_));
  NOR2_X1    g20510(.A1(new_n20764_), .A2(new_n20766_), .ZN(new_n20767_));
  XOR2_X1    g20511(.A1(new_n20761_), .A2(new_n20767_), .Z(new_n20768_));
  NOR2_X1    g20512(.A1(new_n20768_), .A2(new_n20757_), .ZN(new_n20769_));
  INV_X1     g20513(.I(new_n20769_), .ZN(new_n20770_));
  NAND2_X1   g20514(.A1(new_n20768_), .A2(new_n20757_), .ZN(new_n20771_));
  NAND2_X1   g20515(.A1(new_n20770_), .A2(new_n20771_), .ZN(new_n20772_));
  XOR2_X1    g20516(.A1(new_n20772_), .A2(new_n20756_), .Z(new_n20773_));
  OAI22_X1   g20517(.A1(new_n11298_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n11297_), .ZN(new_n20774_));
  AOI21_X1   g20518(.A1(\b[57] ), .A2(new_n11296_), .B(new_n20774_), .ZN(new_n20775_));
  OAI21_X1   g20519(.A1(new_n12203_), .A2(new_n10069_), .B(new_n20775_), .ZN(new_n20776_));
  XOR2_X1    g20520(.A1(new_n20776_), .A2(\a[56] ), .Z(new_n20777_));
  AOI21_X1   g20521(.A1(new_n20701_), .A2(new_n20717_), .B(new_n20718_), .ZN(new_n20778_));
  NOR2_X1    g20522(.A1(new_n20777_), .A2(new_n20778_), .ZN(new_n20779_));
  INV_X1     g20523(.I(new_n20779_), .ZN(new_n20780_));
  NAND2_X1   g20524(.A1(new_n20777_), .A2(new_n20778_), .ZN(new_n20781_));
  NAND2_X1   g20525(.A1(new_n20780_), .A2(new_n20781_), .ZN(new_n20782_));
  XOR2_X1    g20526(.A1(new_n20782_), .A2(new_n20773_), .Z(new_n20783_));
  OAI21_X1   g20527(.A1(new_n20695_), .A2(new_n20722_), .B(new_n20724_), .ZN(new_n20784_));
  INV_X1     g20528(.I(new_n20784_), .ZN(new_n20785_));
  OR2_X2     g20529(.A1(new_n20783_), .A2(new_n20785_), .Z(new_n20786_));
  NAND2_X1   g20530(.A1(new_n20783_), .A2(new_n20785_), .ZN(new_n20787_));
  NAND2_X1   g20531(.A1(new_n20786_), .A2(new_n20787_), .ZN(new_n20788_));
  XOR2_X1    g20532(.A1(new_n20788_), .A2(new_n20752_), .Z(new_n20789_));
  AOI22_X1   g20533(.A1(new_n13460_), .A2(new_n8252_), .B1(\b[63] ), .B2(new_n8575_), .ZN(new_n20790_));
  XOR2_X1    g20534(.A1(new_n20789_), .A2(new_n20790_), .Z(new_n20791_));
  NAND2_X1   g20535(.A1(new_n20727_), .A2(new_n20690_), .ZN(new_n20792_));
  NAND2_X1   g20536(.A1(new_n20792_), .A2(new_n20728_), .ZN(new_n20793_));
  XOR2_X1    g20537(.A1(new_n20793_), .A2(new_n8248_), .Z(new_n20794_));
  XNOR2_X1   g20538(.A1(new_n20791_), .A2(new_n20794_), .ZN(new_n20795_));
  OAI21_X1   g20539(.A1(new_n20682_), .A2(new_n20731_), .B(new_n20733_), .ZN(new_n20796_));
  INV_X1     g20540(.I(new_n20796_), .ZN(new_n20797_));
  NOR2_X1    g20541(.A1(new_n20795_), .A2(new_n20797_), .ZN(new_n20798_));
  NAND2_X1   g20542(.A1(new_n20795_), .A2(new_n20797_), .ZN(new_n20799_));
  INV_X1     g20543(.I(new_n20799_), .ZN(new_n20800_));
  NOR2_X1    g20544(.A1(new_n20800_), .A2(new_n20798_), .ZN(new_n20801_));
  XOR2_X1    g20545(.A1(new_n20748_), .A2(new_n20801_), .Z(\f[113] ));
  NAND2_X1   g20546(.A1(new_n20740_), .A2(new_n20736_), .ZN(new_n20803_));
  INV_X1     g20547(.I(new_n20735_), .ZN(new_n20804_));
  OAI21_X1   g20548(.A1(new_n20740_), .A2(new_n20736_), .B(new_n20804_), .ZN(new_n20805_));
  AOI21_X1   g20549(.A1(new_n20805_), .A2(new_n20803_), .B(new_n20800_), .ZN(new_n20806_));
  AOI22_X1   g20550(.A1(new_n9125_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n9123_), .ZN(new_n20807_));
  OAI21_X1   g20551(.A1(new_n12148_), .A2(new_n9470_), .B(new_n20807_), .ZN(new_n20808_));
  AOI21_X1   g20552(.A1(new_n12811_), .A2(new_n9129_), .B(new_n20808_), .ZN(new_n20809_));
  XOR2_X1    g20553(.A1(new_n20809_), .A2(new_n9133_), .Z(new_n20810_));
  NAND2_X1   g20554(.A1(new_n20787_), .A2(new_n20752_), .ZN(new_n20811_));
  NAND2_X1   g20555(.A1(new_n20811_), .A2(new_n20786_), .ZN(new_n20812_));
  AOI21_X1   g20556(.A1(new_n20773_), .A2(new_n20781_), .B(new_n20779_), .ZN(new_n20813_));
  AOI22_X1   g20557(.A1(new_n10064_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n10062_), .ZN(new_n20814_));
  OAI21_X1   g20558(.A1(new_n11195_), .A2(new_n10399_), .B(new_n20814_), .ZN(new_n20815_));
  AOI21_X1   g20559(.A1(new_n11836_), .A2(new_n10068_), .B(new_n20815_), .ZN(new_n20816_));
  XOR2_X1    g20560(.A1(new_n20816_), .A2(new_n10057_), .Z(new_n20817_));
  INV_X1     g20561(.I(new_n20817_), .ZN(new_n20818_));
  INV_X1     g20562(.I(new_n20756_), .ZN(new_n20819_));
  AOI21_X1   g20563(.A1(new_n20819_), .A2(new_n20771_), .B(new_n20769_), .ZN(new_n20820_));
  AOI22_X1   g20564(.A1(new_n10981_), .A2(\b[57] ), .B1(new_n10979_), .B2(\b[56] ), .ZN(new_n20821_));
  OAI21_X1   g20565(.A1(new_n9972_), .A2(new_n11306_), .B(new_n20821_), .ZN(new_n20822_));
  AOI21_X1   g20566(.A1(new_n10631_), .A2(new_n10984_), .B(new_n20822_), .ZN(new_n20823_));
  XOR2_X1    g20567(.A1(new_n20823_), .A2(new_n10989_), .Z(new_n20824_));
  INV_X1     g20568(.I(new_n20824_), .ZN(new_n20825_));
  AOI22_X1   g20569(.A1(new_n11926_), .A2(\b[54] ), .B1(new_n11924_), .B2(\b[53] ), .ZN(new_n20826_));
  OAI21_X1   g20570(.A1(new_n9032_), .A2(new_n12317_), .B(new_n20826_), .ZN(new_n20827_));
  AOI21_X1   g20571(.A1(new_n10884_), .A2(new_n11929_), .B(new_n20827_), .ZN(new_n20828_));
  XOR2_X1    g20572(.A1(new_n20828_), .A2(new_n12312_), .Z(new_n20829_));
  NOR2_X1    g20573(.A1(new_n20761_), .A2(new_n20766_), .ZN(new_n20830_));
  NOR2_X1    g20574(.A1(new_n20830_), .A2(new_n20764_), .ZN(new_n20831_));
  INV_X1     g20575(.I(new_n20831_), .ZN(new_n20832_));
  AOI22_X1   g20576(.A1(new_n12922_), .A2(\b[51] ), .B1(\b[50] ), .B2(new_n12923_), .ZN(new_n20833_));
  INV_X1     g20577(.I(new_n20833_), .ZN(new_n20834_));
  NOR2_X1    g20578(.A1(new_n20834_), .A2(new_n8248_), .ZN(new_n20835_));
  NOR2_X1    g20579(.A1(new_n20833_), .A2(\a[50] ), .ZN(new_n20836_));
  NOR2_X1    g20580(.A1(new_n20835_), .A2(new_n20836_), .ZN(new_n20837_));
  XOR2_X1    g20581(.A1(new_n20837_), .A2(new_n20710_), .Z(new_n20838_));
  NOR2_X1    g20582(.A1(new_n20832_), .A2(new_n20838_), .ZN(new_n20839_));
  INV_X1     g20583(.I(new_n20839_), .ZN(new_n20840_));
  NAND2_X1   g20584(.A1(new_n20832_), .A2(new_n20838_), .ZN(new_n20841_));
  NAND2_X1   g20585(.A1(new_n20840_), .A2(new_n20841_), .ZN(new_n20842_));
  XOR2_X1    g20586(.A1(new_n20842_), .A2(new_n20829_), .Z(new_n20843_));
  NOR2_X1    g20587(.A1(new_n20843_), .A2(new_n20825_), .ZN(new_n20844_));
  NAND2_X1   g20588(.A1(new_n20843_), .A2(new_n20825_), .ZN(new_n20845_));
  INV_X1     g20589(.I(new_n20845_), .ZN(new_n20846_));
  NOR2_X1    g20590(.A1(new_n20846_), .A2(new_n20844_), .ZN(new_n20847_));
  XNOR2_X1   g20591(.A1(new_n20847_), .A2(new_n20820_), .ZN(new_n20848_));
  NOR2_X1    g20592(.A1(new_n20848_), .A2(new_n20818_), .ZN(new_n20849_));
  INV_X1     g20593(.I(new_n20849_), .ZN(new_n20850_));
  NAND2_X1   g20594(.A1(new_n20848_), .A2(new_n20818_), .ZN(new_n20851_));
  NAND2_X1   g20595(.A1(new_n20850_), .A2(new_n20851_), .ZN(new_n20852_));
  XOR2_X1    g20596(.A1(new_n20852_), .A2(new_n20813_), .Z(new_n20853_));
  NOR2_X1    g20597(.A1(new_n20853_), .A2(new_n20812_), .ZN(new_n20854_));
  INV_X1     g20598(.I(new_n20854_), .ZN(new_n20855_));
  NAND2_X1   g20599(.A1(new_n20853_), .A2(new_n20812_), .ZN(new_n20856_));
  NAND2_X1   g20600(.A1(new_n20855_), .A2(new_n20856_), .ZN(new_n20857_));
  XOR2_X1    g20601(.A1(new_n20857_), .A2(new_n20810_), .Z(new_n20858_));
  INV_X1     g20602(.I(new_n20789_), .ZN(new_n20859_));
  INV_X1     g20603(.I(new_n20793_), .ZN(new_n20860_));
  XOR2_X1    g20604(.A1(new_n20790_), .A2(new_n8248_), .Z(new_n20861_));
  AOI21_X1   g20605(.A1(new_n20860_), .A2(new_n20789_), .B(new_n20861_), .ZN(new_n20862_));
  AOI21_X1   g20606(.A1(new_n20859_), .A2(new_n20793_), .B(new_n20862_), .ZN(new_n20863_));
  INV_X1     g20607(.I(new_n20863_), .ZN(new_n20864_));
  NOR2_X1    g20608(.A1(new_n20858_), .A2(new_n20864_), .ZN(new_n20865_));
  INV_X1     g20609(.I(new_n20865_), .ZN(new_n20866_));
  NAND2_X1   g20610(.A1(new_n20858_), .A2(new_n20864_), .ZN(new_n20867_));
  AND2_X2    g20611(.A1(new_n20866_), .A2(new_n20867_), .Z(new_n20868_));
  INV_X1     g20612(.I(new_n20868_), .ZN(new_n20869_));
  NOR3_X1    g20613(.A1(new_n20806_), .A2(new_n20798_), .A3(new_n20869_), .ZN(new_n20870_));
  INV_X1     g20614(.I(new_n20798_), .ZN(new_n20871_));
  OAI21_X1   g20615(.A1(new_n20747_), .A2(new_n20744_), .B(new_n20799_), .ZN(new_n20872_));
  AOI21_X1   g20616(.A1(new_n20872_), .A2(new_n20871_), .B(new_n20868_), .ZN(new_n20873_));
  NOR2_X1    g20617(.A1(new_n20870_), .A2(new_n20873_), .ZN(\f[114] ));
  OAI22_X1   g20618(.A1(new_n10389_), .A2(new_n12800_), .B1(new_n9470_), .B2(new_n12796_), .ZN(new_n20875_));
  AOI21_X1   g20619(.A1(new_n13973_), .A2(new_n9129_), .B(new_n20875_), .ZN(new_n20876_));
  XOR2_X1    g20620(.A1(new_n20876_), .A2(new_n9133_), .Z(new_n20877_));
  INV_X1     g20621(.I(new_n20877_), .ZN(new_n20878_));
  OAI21_X1   g20622(.A1(new_n20813_), .A2(new_n20849_), .B(new_n20851_), .ZN(new_n20879_));
  OAI22_X1   g20623(.A1(new_n11298_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n11297_), .ZN(new_n20880_));
  AOI21_X1   g20624(.A1(\b[59] ), .A2(new_n11296_), .B(new_n20880_), .ZN(new_n20881_));
  OAI21_X1   g20625(.A1(new_n13110_), .A2(new_n10069_), .B(new_n20881_), .ZN(new_n20882_));
  XOR2_X1    g20626(.A1(new_n20882_), .A2(new_n10057_), .Z(new_n20883_));
  OAI21_X1   g20627(.A1(new_n20820_), .A2(new_n20844_), .B(new_n20845_), .ZN(new_n20884_));
  AOI22_X1   g20628(.A1(new_n10981_), .A2(\b[58] ), .B1(new_n10979_), .B2(\b[57] ), .ZN(new_n20885_));
  OAI21_X1   g20629(.A1(new_n10308_), .A2(new_n11306_), .B(new_n20885_), .ZN(new_n20886_));
  AOI21_X1   g20630(.A1(new_n12164_), .A2(new_n10984_), .B(new_n20886_), .ZN(new_n20887_));
  XOR2_X1    g20631(.A1(new_n20887_), .A2(new_n10989_), .Z(new_n20888_));
  OAI21_X1   g20632(.A1(new_n20829_), .A2(new_n20839_), .B(new_n20841_), .ZN(new_n20889_));
  AOI22_X1   g20633(.A1(new_n11926_), .A2(\b[55] ), .B1(new_n11924_), .B2(\b[54] ), .ZN(new_n20890_));
  OAI21_X1   g20634(.A1(new_n9376_), .A2(new_n12317_), .B(new_n20890_), .ZN(new_n20891_));
  AOI21_X1   g20635(.A1(new_n9979_), .A2(new_n11929_), .B(new_n20891_), .ZN(new_n20892_));
  XOR2_X1    g20636(.A1(new_n20892_), .A2(new_n12312_), .Z(new_n20893_));
  INV_X1     g20637(.I(new_n20836_), .ZN(new_n20894_));
  AOI21_X1   g20638(.A1(new_n20710_), .A2(new_n20894_), .B(new_n20835_), .ZN(new_n20895_));
  AOI22_X1   g20639(.A1(new_n12922_), .A2(\b[52] ), .B1(\b[51] ), .B2(new_n12923_), .ZN(new_n20896_));
  AND2_X2    g20640(.A1(new_n20895_), .A2(new_n20896_), .Z(new_n20897_));
  NOR2_X1    g20641(.A1(new_n20895_), .A2(new_n20896_), .ZN(new_n20898_));
  NOR2_X1    g20642(.A1(new_n20897_), .A2(new_n20898_), .ZN(new_n20899_));
  XNOR2_X1   g20643(.A1(new_n20893_), .A2(new_n20899_), .ZN(new_n20900_));
  NOR2_X1    g20644(.A1(new_n20900_), .A2(new_n20889_), .ZN(new_n20901_));
  INV_X1     g20645(.I(new_n20901_), .ZN(new_n20902_));
  NAND2_X1   g20646(.A1(new_n20900_), .A2(new_n20889_), .ZN(new_n20903_));
  NAND2_X1   g20647(.A1(new_n20902_), .A2(new_n20903_), .ZN(new_n20904_));
  XOR2_X1    g20648(.A1(new_n20904_), .A2(new_n20888_), .Z(new_n20905_));
  OR2_X2     g20649(.A1(new_n20905_), .A2(new_n20884_), .Z(new_n20906_));
  NAND2_X1   g20650(.A1(new_n20905_), .A2(new_n20884_), .ZN(new_n20907_));
  NAND2_X1   g20651(.A1(new_n20906_), .A2(new_n20907_), .ZN(new_n20908_));
  XNOR2_X1   g20652(.A1(new_n20908_), .A2(new_n20883_), .ZN(new_n20909_));
  NOR2_X1    g20653(.A1(new_n20909_), .A2(new_n20879_), .ZN(new_n20910_));
  INV_X1     g20654(.I(new_n20910_), .ZN(new_n20911_));
  NAND2_X1   g20655(.A1(new_n20909_), .A2(new_n20879_), .ZN(new_n20912_));
  NAND2_X1   g20656(.A1(new_n20911_), .A2(new_n20912_), .ZN(new_n20913_));
  XOR2_X1    g20657(.A1(new_n20913_), .A2(new_n20878_), .Z(new_n20914_));
  INV_X1     g20658(.I(new_n20914_), .ZN(new_n20915_));
  OAI21_X1   g20659(.A1(new_n20810_), .A2(new_n20854_), .B(new_n20856_), .ZN(new_n20916_));
  INV_X1     g20660(.I(new_n20916_), .ZN(new_n20917_));
  OAI21_X1   g20661(.A1(new_n20870_), .A2(new_n20865_), .B(new_n20917_), .ZN(new_n20918_));
  NAND3_X1   g20662(.A1(new_n20872_), .A2(new_n20871_), .A3(new_n20868_), .ZN(new_n20919_));
  NAND3_X1   g20663(.A1(new_n20919_), .A2(new_n20866_), .A3(new_n20916_), .ZN(new_n20920_));
  NAND2_X1   g20664(.A1(new_n20918_), .A2(new_n20920_), .ZN(new_n20921_));
  XOR2_X1    g20665(.A1(new_n20921_), .A2(new_n20915_), .Z(\f[115] ));
  AOI21_X1   g20666(.A1(new_n20919_), .A2(new_n20866_), .B(new_n20916_), .ZN(new_n20923_));
  OAI21_X1   g20667(.A1(new_n20914_), .A2(new_n20923_), .B(new_n20920_), .ZN(new_n20924_));
  AOI22_X1   g20668(.A1(new_n13460_), .A2(new_n9129_), .B1(\b[63] ), .B2(new_n9471_), .ZN(new_n20925_));
  AOI22_X1   g20669(.A1(new_n10064_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n10062_), .ZN(new_n20926_));
  OAI21_X1   g20670(.A1(new_n12147_), .A2(new_n10399_), .B(new_n20926_), .ZN(new_n20927_));
  AOI21_X1   g20671(.A1(new_n13444_), .A2(new_n10068_), .B(new_n20927_), .ZN(new_n20928_));
  XOR2_X1    g20672(.A1(new_n20928_), .A2(new_n10057_), .Z(new_n20929_));
  OAI21_X1   g20673(.A1(new_n20888_), .A2(new_n20901_), .B(new_n20903_), .ZN(new_n20930_));
  OAI22_X1   g20674(.A1(new_n12306_), .A2(new_n12151_), .B1(new_n12305_), .B2(new_n11195_), .ZN(new_n20931_));
  AOI21_X1   g20675(.A1(\b[57] ), .A2(new_n12304_), .B(new_n20931_), .ZN(new_n20932_));
  OAI21_X1   g20676(.A1(new_n12203_), .A2(new_n10985_), .B(new_n20932_), .ZN(new_n20933_));
  XOR2_X1    g20677(.A1(new_n20933_), .A2(\a[59] ), .Z(new_n20934_));
  AOI22_X1   g20678(.A1(new_n11926_), .A2(\b[56] ), .B1(new_n11924_), .B2(\b[55] ), .ZN(new_n20935_));
  OAI21_X1   g20679(.A1(new_n9942_), .A2(new_n12317_), .B(new_n20935_), .ZN(new_n20936_));
  AOI21_X1   g20680(.A1(new_n10318_), .A2(new_n11929_), .B(new_n20936_), .ZN(new_n20937_));
  XOR2_X1    g20681(.A1(new_n20937_), .A2(new_n12312_), .Z(new_n20938_));
  NOR2_X1    g20682(.A1(new_n20934_), .A2(new_n20938_), .ZN(new_n20939_));
  INV_X1     g20683(.I(new_n20939_), .ZN(new_n20940_));
  NAND2_X1   g20684(.A1(new_n20934_), .A2(new_n20938_), .ZN(new_n20941_));
  NAND2_X1   g20685(.A1(new_n20940_), .A2(new_n20941_), .ZN(new_n20942_));
  NOR2_X1    g20686(.A1(new_n20893_), .A2(new_n20897_), .ZN(new_n20943_));
  NOR2_X1    g20687(.A1(new_n20943_), .A2(new_n20898_), .ZN(new_n20944_));
  AOI22_X1   g20688(.A1(new_n12922_), .A2(\b[53] ), .B1(\b[52] ), .B2(new_n12923_), .ZN(new_n20945_));
  INV_X1     g20689(.I(new_n20945_), .ZN(new_n20946_));
  NOR2_X1    g20690(.A1(new_n20946_), .A2(new_n20896_), .ZN(new_n20947_));
  INV_X1     g20691(.I(new_n20896_), .ZN(new_n20948_));
  NOR2_X1    g20692(.A1(new_n20948_), .A2(new_n20945_), .ZN(new_n20949_));
  OR2_X2     g20693(.A1(new_n20947_), .A2(new_n20949_), .Z(new_n20950_));
  XNOR2_X1   g20694(.A1(new_n20944_), .A2(new_n20950_), .ZN(new_n20951_));
  XOR2_X1    g20695(.A1(new_n20942_), .A2(new_n20951_), .Z(new_n20952_));
  NOR2_X1    g20696(.A1(new_n20952_), .A2(new_n20930_), .ZN(new_n20953_));
  NAND2_X1   g20697(.A1(new_n20952_), .A2(new_n20930_), .ZN(new_n20954_));
  INV_X1     g20698(.I(new_n20954_), .ZN(new_n20955_));
  NOR2_X1    g20699(.A1(new_n20955_), .A2(new_n20953_), .ZN(new_n20956_));
  XOR2_X1    g20700(.A1(new_n20956_), .A2(new_n20929_), .Z(new_n20957_));
  XOR2_X1    g20701(.A1(new_n20957_), .A2(new_n20925_), .Z(new_n20958_));
  NAND2_X1   g20702(.A1(new_n20906_), .A2(new_n20883_), .ZN(new_n20959_));
  NAND2_X1   g20703(.A1(new_n20959_), .A2(new_n20907_), .ZN(new_n20960_));
  XOR2_X1    g20704(.A1(new_n20960_), .A2(\a[53] ), .Z(new_n20961_));
  XOR2_X1    g20705(.A1(new_n20958_), .A2(new_n20961_), .Z(new_n20962_));
  OAI21_X1   g20706(.A1(new_n20877_), .A2(new_n20910_), .B(new_n20912_), .ZN(new_n20963_));
  INV_X1     g20707(.I(new_n20963_), .ZN(new_n20964_));
  NOR2_X1    g20708(.A1(new_n20962_), .A2(new_n20964_), .ZN(new_n20965_));
  INV_X1     g20709(.I(new_n20965_), .ZN(new_n20966_));
  NAND2_X1   g20710(.A1(new_n20962_), .A2(new_n20964_), .ZN(new_n20967_));
  NAND2_X1   g20711(.A1(new_n20966_), .A2(new_n20967_), .ZN(new_n20968_));
  XOR2_X1    g20712(.A1(new_n20924_), .A2(new_n20968_), .Z(\f[116] ));
  INV_X1     g20713(.I(new_n20960_), .ZN(new_n20970_));
  NAND2_X1   g20714(.A1(new_n20957_), .A2(new_n20970_), .ZN(new_n20971_));
  XOR2_X1    g20715(.A1(new_n20925_), .A2(\a[53] ), .Z(new_n20972_));
  NAND2_X1   g20716(.A1(new_n20971_), .A2(new_n20972_), .ZN(new_n20973_));
  OAI21_X1   g20717(.A1(new_n20957_), .A2(new_n20970_), .B(new_n20973_), .ZN(new_n20974_));
  OAI21_X1   g20718(.A1(new_n20929_), .A2(new_n20953_), .B(new_n20954_), .ZN(new_n20975_));
  AOI22_X1   g20719(.A1(new_n10064_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n10062_), .ZN(new_n20976_));
  OAI21_X1   g20720(.A1(new_n12148_), .A2(new_n10399_), .B(new_n20976_), .ZN(new_n20977_));
  AOI21_X1   g20721(.A1(new_n12811_), .A2(new_n10068_), .B(new_n20977_), .ZN(new_n20978_));
  XOR2_X1    g20722(.A1(new_n20978_), .A2(new_n10057_), .Z(new_n20979_));
  INV_X1     g20723(.I(new_n20951_), .ZN(new_n20980_));
  AOI21_X1   g20724(.A1(new_n20980_), .A2(new_n20941_), .B(new_n20939_), .ZN(new_n20981_));
  AOI22_X1   g20725(.A1(new_n10981_), .A2(\b[60] ), .B1(new_n10979_), .B2(\b[59] ), .ZN(new_n20982_));
  OAI21_X1   g20726(.A1(new_n11195_), .A2(new_n11306_), .B(new_n20982_), .ZN(new_n20983_));
  AOI21_X1   g20727(.A1(new_n11836_), .A2(new_n10984_), .B(new_n20983_), .ZN(new_n20984_));
  XOR2_X1    g20728(.A1(new_n20984_), .A2(new_n10989_), .Z(new_n20985_));
  INV_X1     g20729(.I(new_n20985_), .ZN(new_n20986_));
  INV_X1     g20730(.I(new_n20949_), .ZN(new_n20987_));
  OAI21_X1   g20731(.A1(new_n20944_), .A2(new_n20947_), .B(new_n20987_), .ZN(new_n20988_));
  INV_X1     g20732(.I(new_n20988_), .ZN(new_n20989_));
  AOI22_X1   g20733(.A1(new_n11926_), .A2(\b[57] ), .B1(new_n11924_), .B2(\b[56] ), .ZN(new_n20990_));
  OAI21_X1   g20734(.A1(new_n9972_), .A2(new_n12317_), .B(new_n20990_), .ZN(new_n20991_));
  AOI21_X1   g20735(.A1(new_n10631_), .A2(new_n11929_), .B(new_n20991_), .ZN(new_n20992_));
  XOR2_X1    g20736(.A1(new_n20992_), .A2(new_n12312_), .Z(new_n20993_));
  INV_X1     g20737(.I(new_n20993_), .ZN(new_n20994_));
  AOI22_X1   g20738(.A1(new_n12922_), .A2(\b[54] ), .B1(\b[53] ), .B2(new_n12923_), .ZN(new_n20995_));
  INV_X1     g20739(.I(new_n20995_), .ZN(new_n20996_));
  NOR2_X1    g20740(.A1(new_n20996_), .A2(new_n9133_), .ZN(new_n20997_));
  NOR2_X1    g20741(.A1(new_n20995_), .A2(\a[53] ), .ZN(new_n20998_));
  NOR2_X1    g20742(.A1(new_n20997_), .A2(new_n20998_), .ZN(new_n20999_));
  XOR2_X1    g20743(.A1(new_n20999_), .A2(new_n20945_), .Z(new_n21000_));
  NOR2_X1    g20744(.A1(new_n20994_), .A2(new_n21000_), .ZN(new_n21001_));
  INV_X1     g20745(.I(new_n21001_), .ZN(new_n21002_));
  NAND2_X1   g20746(.A1(new_n20994_), .A2(new_n21000_), .ZN(new_n21003_));
  NAND2_X1   g20747(.A1(new_n21002_), .A2(new_n21003_), .ZN(new_n21004_));
  XOR2_X1    g20748(.A1(new_n21004_), .A2(new_n20989_), .Z(new_n21005_));
  NOR2_X1    g20749(.A1(new_n21005_), .A2(new_n20986_), .ZN(new_n21006_));
  NAND2_X1   g20750(.A1(new_n21005_), .A2(new_n20986_), .ZN(new_n21007_));
  INV_X1     g20751(.I(new_n21007_), .ZN(new_n21008_));
  NOR2_X1    g20752(.A1(new_n21008_), .A2(new_n21006_), .ZN(new_n21009_));
  XOR2_X1    g20753(.A1(new_n21009_), .A2(new_n20981_), .Z(new_n21010_));
  NOR2_X1    g20754(.A1(new_n21010_), .A2(new_n20979_), .ZN(new_n21011_));
  NAND2_X1   g20755(.A1(new_n21010_), .A2(new_n20979_), .ZN(new_n21012_));
  INV_X1     g20756(.I(new_n21012_), .ZN(new_n21013_));
  NOR2_X1    g20757(.A1(new_n21013_), .A2(new_n21011_), .ZN(new_n21014_));
  XOR2_X1    g20758(.A1(new_n21014_), .A2(new_n20975_), .Z(new_n21015_));
  XNOR2_X1   g20759(.A1(new_n21015_), .A2(new_n20974_), .ZN(new_n21016_));
  INV_X1     g20760(.I(new_n21016_), .ZN(new_n21017_));
  AOI21_X1   g20761(.A1(new_n20924_), .A2(new_n20967_), .B(new_n20965_), .ZN(new_n21018_));
  XOR2_X1    g20762(.A1(new_n21018_), .A2(new_n21017_), .Z(\f[117] ));
  OAI22_X1   g20763(.A1(new_n11297_), .A2(new_n12800_), .B1(new_n12796_), .B2(new_n10399_), .ZN(new_n21020_));
  AOI21_X1   g20764(.A1(new_n13973_), .A2(new_n10068_), .B(new_n21020_), .ZN(new_n21021_));
  XOR2_X1    g20765(.A1(new_n21021_), .A2(new_n10057_), .Z(new_n21022_));
  INV_X1     g20766(.I(new_n21022_), .ZN(new_n21023_));
  OAI21_X1   g20767(.A1(new_n20981_), .A2(new_n21006_), .B(new_n21007_), .ZN(new_n21024_));
  OAI22_X1   g20768(.A1(new_n12306_), .A2(new_n12148_), .B1(new_n12305_), .B2(new_n12147_), .ZN(new_n21025_));
  AOI21_X1   g20769(.A1(\b[59] ), .A2(new_n12304_), .B(new_n21025_), .ZN(new_n21026_));
  OAI21_X1   g20770(.A1(new_n13110_), .A2(new_n10985_), .B(new_n21026_), .ZN(new_n21027_));
  XOR2_X1    g20771(.A1(new_n21027_), .A2(new_n10989_), .Z(new_n21028_));
  OAI21_X1   g20772(.A1(new_n20989_), .A2(new_n21001_), .B(new_n21003_), .ZN(new_n21029_));
  AOI22_X1   g20773(.A1(new_n11926_), .A2(\b[58] ), .B1(new_n11924_), .B2(\b[57] ), .ZN(new_n21030_));
  OAI21_X1   g20774(.A1(new_n10308_), .A2(new_n12317_), .B(new_n21030_), .ZN(new_n21031_));
  AOI21_X1   g20775(.A1(new_n12164_), .A2(new_n11929_), .B(new_n21031_), .ZN(new_n21032_));
  XOR2_X1    g20776(.A1(new_n21032_), .A2(\a[62] ), .Z(new_n21033_));
  NOR2_X1    g20777(.A1(new_n20998_), .A2(new_n20946_), .ZN(new_n21034_));
  NOR2_X1    g20778(.A1(new_n21034_), .A2(new_n20997_), .ZN(new_n21035_));
  AOI22_X1   g20779(.A1(new_n12922_), .A2(\b[55] ), .B1(\b[54] ), .B2(new_n12923_), .ZN(new_n21036_));
  NAND2_X1   g20780(.A1(new_n21035_), .A2(new_n21036_), .ZN(new_n21037_));
  NOR2_X1    g20781(.A1(new_n21035_), .A2(new_n21036_), .ZN(new_n21038_));
  INV_X1     g20782(.I(new_n21038_), .ZN(new_n21039_));
  NAND2_X1   g20783(.A1(new_n21039_), .A2(new_n21037_), .ZN(new_n21040_));
  XNOR2_X1   g20784(.A1(new_n21033_), .A2(new_n21040_), .ZN(new_n21041_));
  OR2_X2     g20785(.A1(new_n21029_), .A2(new_n21041_), .Z(new_n21042_));
  NAND2_X1   g20786(.A1(new_n21029_), .A2(new_n21041_), .ZN(new_n21043_));
  NAND2_X1   g20787(.A1(new_n21042_), .A2(new_n21043_), .ZN(new_n21044_));
  XNOR2_X1   g20788(.A1(new_n21028_), .A2(new_n21044_), .ZN(new_n21045_));
  NOR2_X1    g20789(.A1(new_n21045_), .A2(new_n21024_), .ZN(new_n21046_));
  INV_X1     g20790(.I(new_n21046_), .ZN(new_n21047_));
  NAND2_X1   g20791(.A1(new_n21045_), .A2(new_n21024_), .ZN(new_n21048_));
  NAND2_X1   g20792(.A1(new_n21047_), .A2(new_n21048_), .ZN(new_n21049_));
  XOR2_X1    g20793(.A1(new_n21049_), .A2(new_n21023_), .Z(new_n21050_));
  AOI21_X1   g20794(.A1(new_n20975_), .A2(new_n21012_), .B(new_n21011_), .ZN(new_n21051_));
  INV_X1     g20795(.I(new_n21051_), .ZN(new_n21052_));
  NOR2_X1    g20796(.A1(new_n21015_), .A2(new_n20974_), .ZN(new_n21053_));
  AOI21_X1   g20797(.A1(new_n21018_), .A2(new_n21017_), .B(new_n21053_), .ZN(new_n21054_));
  NOR2_X1    g20798(.A1(new_n21054_), .A2(new_n21052_), .ZN(new_n21055_));
  NOR3_X1    g20799(.A1(new_n20870_), .A2(new_n20865_), .A3(new_n20917_), .ZN(new_n21056_));
  AOI21_X1   g20800(.A1(new_n20915_), .A2(new_n20918_), .B(new_n21056_), .ZN(new_n21057_));
  INV_X1     g20801(.I(new_n20967_), .ZN(new_n21058_));
  OAI21_X1   g20802(.A1(new_n21057_), .A2(new_n21058_), .B(new_n20966_), .ZN(new_n21059_));
  INV_X1     g20803(.I(new_n21053_), .ZN(new_n21060_));
  OAI21_X1   g20804(.A1(new_n21059_), .A2(new_n21016_), .B(new_n21060_), .ZN(new_n21061_));
  NOR2_X1    g20805(.A1(new_n21061_), .A2(new_n21051_), .ZN(new_n21062_));
  NOR2_X1    g20806(.A1(new_n21062_), .A2(new_n21055_), .ZN(new_n21063_));
  XOR2_X1    g20807(.A1(new_n21063_), .A2(new_n21050_), .Z(\f[118] ));
  NAND2_X1   g20808(.A1(new_n21054_), .A2(new_n21052_), .ZN(new_n21065_));
  INV_X1     g20809(.I(new_n21050_), .ZN(new_n21066_));
  OAI21_X1   g20810(.A1(new_n21054_), .A2(new_n21052_), .B(new_n21066_), .ZN(new_n21067_));
  NAND2_X1   g20811(.A1(new_n21067_), .A2(new_n21065_), .ZN(new_n21068_));
  AOI22_X1   g20812(.A1(new_n10981_), .A2(\b[62] ), .B1(new_n10979_), .B2(\b[61] ), .ZN(new_n21069_));
  OAI21_X1   g20813(.A1(new_n12147_), .A2(new_n11306_), .B(new_n21069_), .ZN(new_n21070_));
  AOI21_X1   g20814(.A1(new_n13444_), .A2(new_n10984_), .B(new_n21070_), .ZN(new_n21071_));
  XOR2_X1    g20815(.A1(new_n21071_), .A2(new_n10989_), .Z(new_n21072_));
  AOI21_X1   g20816(.A1(new_n21033_), .A2(new_n21037_), .B(new_n21038_), .ZN(new_n21073_));
  OAI22_X1   g20817(.A1(new_n13224_), .A2(new_n12151_), .B1(new_n11195_), .B2(new_n11923_), .ZN(new_n21074_));
  AOI21_X1   g20818(.A1(\b[57] ), .A2(new_n13223_), .B(new_n21074_), .ZN(new_n21075_));
  OAI21_X1   g20819(.A1(new_n12203_), .A2(new_n11930_), .B(new_n21075_), .ZN(new_n21076_));
  XOR2_X1    g20820(.A1(new_n21076_), .A2(new_n12312_), .Z(new_n21077_));
  AOI22_X1   g20821(.A1(new_n12922_), .A2(\b[56] ), .B1(\b[55] ), .B2(new_n12923_), .ZN(new_n21078_));
  INV_X1     g20822(.I(new_n21078_), .ZN(new_n21079_));
  NOR2_X1    g20823(.A1(new_n21079_), .A2(new_n21036_), .ZN(new_n21080_));
  INV_X1     g20824(.I(new_n21080_), .ZN(new_n21081_));
  NAND2_X1   g20825(.A1(new_n21079_), .A2(new_n21036_), .ZN(new_n21082_));
  NAND2_X1   g20826(.A1(new_n21081_), .A2(new_n21082_), .ZN(new_n21083_));
  XOR2_X1    g20827(.A1(new_n21077_), .A2(new_n21083_), .Z(new_n21084_));
  NOR2_X1    g20828(.A1(new_n21084_), .A2(new_n21073_), .ZN(new_n21085_));
  NAND2_X1   g20829(.A1(new_n21084_), .A2(new_n21073_), .ZN(new_n21086_));
  INV_X1     g20830(.I(new_n21086_), .ZN(new_n21087_));
  NOR2_X1    g20831(.A1(new_n21087_), .A2(new_n21085_), .ZN(new_n21088_));
  XOR2_X1    g20832(.A1(new_n21088_), .A2(new_n21072_), .Z(new_n21089_));
  AOI22_X1   g20833(.A1(new_n13460_), .A2(new_n10068_), .B1(\b[63] ), .B2(new_n11296_), .ZN(new_n21090_));
  XNOR2_X1   g20834(.A1(new_n21089_), .A2(new_n21090_), .ZN(new_n21091_));
  NAND2_X1   g20835(.A1(new_n21028_), .A2(new_n21042_), .ZN(new_n21092_));
  NAND2_X1   g20836(.A1(new_n21092_), .A2(new_n21043_), .ZN(new_n21093_));
  XOR2_X1    g20837(.A1(new_n21093_), .A2(new_n10057_), .Z(new_n21094_));
  XOR2_X1    g20838(.A1(new_n21091_), .A2(new_n21094_), .Z(new_n21095_));
  OAI21_X1   g20839(.A1(new_n21022_), .A2(new_n21046_), .B(new_n21048_), .ZN(new_n21096_));
  INV_X1     g20840(.I(new_n21096_), .ZN(new_n21097_));
  NOR2_X1    g20841(.A1(new_n21095_), .A2(new_n21097_), .ZN(new_n21098_));
  INV_X1     g20842(.I(new_n21098_), .ZN(new_n21099_));
  NAND2_X1   g20843(.A1(new_n21095_), .A2(new_n21097_), .ZN(new_n21100_));
  NAND2_X1   g20844(.A1(new_n21099_), .A2(new_n21100_), .ZN(new_n21101_));
  XOR2_X1    g20845(.A1(new_n21068_), .A2(new_n21101_), .Z(\f[119] ));
  INV_X1     g20846(.I(new_n21100_), .ZN(new_n21103_));
  AOI21_X1   g20847(.A1(new_n21067_), .A2(new_n21065_), .B(new_n21103_), .ZN(new_n21104_));
  NOR2_X1    g20848(.A1(new_n21104_), .A2(new_n21098_), .ZN(new_n21105_));
  NOR2_X1    g20849(.A1(new_n21072_), .A2(new_n21087_), .ZN(new_n21106_));
  NOR2_X1    g20850(.A1(new_n21106_), .A2(new_n21085_), .ZN(new_n21107_));
  AOI22_X1   g20851(.A1(new_n10981_), .A2(\b[63] ), .B1(new_n10979_), .B2(\b[62] ), .ZN(new_n21108_));
  OAI21_X1   g20852(.A1(new_n12148_), .A2(new_n11306_), .B(new_n21108_), .ZN(new_n21109_));
  AOI21_X1   g20853(.A1(new_n12811_), .A2(new_n10984_), .B(new_n21109_), .ZN(new_n21110_));
  XOR2_X1    g20854(.A1(new_n21110_), .A2(new_n10989_), .Z(new_n21111_));
  INV_X1     g20855(.I(new_n21111_), .ZN(new_n21112_));
  AOI21_X1   g20856(.A1(new_n21077_), .A2(new_n21082_), .B(new_n21080_), .ZN(new_n21113_));
  AOI22_X1   g20857(.A1(new_n11926_), .A2(\b[60] ), .B1(new_n11924_), .B2(\b[59] ), .ZN(new_n21114_));
  OAI21_X1   g20858(.A1(new_n11195_), .A2(new_n12317_), .B(new_n21114_), .ZN(new_n21115_));
  AOI21_X1   g20859(.A1(new_n11836_), .A2(new_n11929_), .B(new_n21115_), .ZN(new_n21116_));
  XOR2_X1    g20860(.A1(new_n21116_), .A2(new_n12312_), .Z(new_n21117_));
  AOI22_X1   g20861(.A1(new_n12922_), .A2(\b[57] ), .B1(\b[56] ), .B2(new_n12923_), .ZN(new_n21118_));
  XOR2_X1    g20862(.A1(new_n21118_), .A2(new_n10057_), .Z(new_n21119_));
  XOR2_X1    g20863(.A1(new_n21119_), .A2(new_n21036_), .Z(new_n21120_));
  NOR2_X1    g20864(.A1(new_n21117_), .A2(new_n21120_), .ZN(new_n21121_));
  INV_X1     g20865(.I(new_n21121_), .ZN(new_n21122_));
  NAND2_X1   g20866(.A1(new_n21117_), .A2(new_n21120_), .ZN(new_n21123_));
  NAND2_X1   g20867(.A1(new_n21122_), .A2(new_n21123_), .ZN(new_n21124_));
  XOR2_X1    g20868(.A1(new_n21124_), .A2(new_n21113_), .Z(new_n21125_));
  NOR2_X1    g20869(.A1(new_n21125_), .A2(new_n21112_), .ZN(new_n21126_));
  NAND2_X1   g20870(.A1(new_n21125_), .A2(new_n21112_), .ZN(new_n21127_));
  INV_X1     g20871(.I(new_n21127_), .ZN(new_n21128_));
  NOR2_X1    g20872(.A1(new_n21128_), .A2(new_n21126_), .ZN(new_n21129_));
  XOR2_X1    g20873(.A1(new_n21129_), .A2(new_n21107_), .Z(new_n21130_));
  INV_X1     g20874(.I(new_n21130_), .ZN(new_n21131_));
  INV_X1     g20875(.I(new_n21093_), .ZN(new_n21132_));
  NOR2_X1    g20876(.A1(new_n21132_), .A2(new_n21089_), .ZN(new_n21133_));
  XOR2_X1    g20877(.A1(new_n21090_), .A2(new_n10057_), .Z(new_n21134_));
  AOI21_X1   g20878(.A1(new_n21132_), .A2(new_n21089_), .B(new_n21134_), .ZN(new_n21135_));
  NOR2_X1    g20879(.A1(new_n21135_), .A2(new_n21133_), .ZN(new_n21136_));
  INV_X1     g20880(.I(new_n21136_), .ZN(new_n21137_));
  NOR2_X1    g20881(.A1(new_n21131_), .A2(new_n21137_), .ZN(new_n21138_));
  INV_X1     g20882(.I(new_n21138_), .ZN(new_n21139_));
  NAND2_X1   g20883(.A1(new_n21131_), .A2(new_n21137_), .ZN(new_n21140_));
  AND2_X2    g20884(.A1(new_n21139_), .A2(new_n21140_), .Z(new_n21141_));
  XOR2_X1    g20885(.A1(new_n21105_), .A2(new_n21141_), .Z(\f[120] ));
  OAI22_X1   g20886(.A1(new_n12305_), .A2(new_n12800_), .B1(new_n11306_), .B2(new_n12796_), .ZN(new_n21143_));
  AOI21_X1   g20887(.A1(new_n13973_), .A2(new_n10984_), .B(new_n21143_), .ZN(new_n21144_));
  XOR2_X1    g20888(.A1(new_n21144_), .A2(new_n10989_), .Z(new_n21145_));
  INV_X1     g20889(.I(new_n21145_), .ZN(new_n21146_));
  INV_X1     g20890(.I(new_n21113_), .ZN(new_n21147_));
  AOI21_X1   g20891(.A1(new_n21147_), .A2(new_n21123_), .B(new_n21121_), .ZN(new_n21148_));
  INV_X1     g20892(.I(new_n21148_), .ZN(new_n21149_));
  OAI22_X1   g20893(.A1(new_n13224_), .A2(new_n12148_), .B1(new_n12147_), .B2(new_n11923_), .ZN(new_n21150_));
  AOI21_X1   g20894(.A1(\b[59] ), .A2(new_n13223_), .B(new_n21150_), .ZN(new_n21151_));
  OAI21_X1   g20895(.A1(new_n13110_), .A2(new_n11930_), .B(new_n21151_), .ZN(new_n21152_));
  XOR2_X1    g20896(.A1(new_n21152_), .A2(new_n12312_), .Z(new_n21153_));
  OAI21_X1   g20897(.A1(\a[56] ), .A2(new_n21118_), .B(new_n21036_), .ZN(new_n21154_));
  INV_X1     g20898(.I(new_n21154_), .ZN(new_n21155_));
  AOI21_X1   g20899(.A1(\a[56] ), .A2(new_n21118_), .B(new_n21155_), .ZN(new_n21156_));
  AOI22_X1   g20900(.A1(new_n12922_), .A2(\b[58] ), .B1(\b[57] ), .B2(new_n12923_), .ZN(new_n21157_));
  NAND2_X1   g20901(.A1(new_n21156_), .A2(new_n21157_), .ZN(new_n21158_));
  OR2_X2     g20902(.A1(new_n21156_), .A2(new_n21157_), .Z(new_n21159_));
  NAND2_X1   g20903(.A1(new_n21159_), .A2(new_n21158_), .ZN(new_n21160_));
  XNOR2_X1   g20904(.A1(new_n21153_), .A2(new_n21160_), .ZN(new_n21161_));
  NOR2_X1    g20905(.A1(new_n21161_), .A2(new_n21149_), .ZN(new_n21162_));
  INV_X1     g20906(.I(new_n21162_), .ZN(new_n21163_));
  NAND2_X1   g20907(.A1(new_n21161_), .A2(new_n21149_), .ZN(new_n21164_));
  NAND2_X1   g20908(.A1(new_n21163_), .A2(new_n21164_), .ZN(new_n21165_));
  XOR2_X1    g20909(.A1(new_n21165_), .A2(new_n21146_), .Z(new_n21166_));
  INV_X1     g20910(.I(new_n21166_), .ZN(new_n21167_));
  OAI21_X1   g20911(.A1(new_n21107_), .A2(new_n21126_), .B(new_n21127_), .ZN(new_n21168_));
  INV_X1     g20912(.I(new_n21168_), .ZN(new_n21169_));
  INV_X1     g20913(.I(new_n21141_), .ZN(new_n21170_));
  NOR3_X1    g20914(.A1(new_n21104_), .A2(new_n21098_), .A3(new_n21170_), .ZN(new_n21171_));
  OAI21_X1   g20915(.A1(new_n21171_), .A2(new_n21138_), .B(new_n21169_), .ZN(new_n21172_));
  AOI21_X1   g20916(.A1(new_n21061_), .A2(new_n21051_), .B(new_n21050_), .ZN(new_n21173_));
  OAI21_X1   g20917(.A1(new_n21173_), .A2(new_n21062_), .B(new_n21100_), .ZN(new_n21174_));
  NAND3_X1   g20918(.A1(new_n21174_), .A2(new_n21099_), .A3(new_n21141_), .ZN(new_n21175_));
  NAND3_X1   g20919(.A1(new_n21175_), .A2(new_n21139_), .A3(new_n21168_), .ZN(new_n21176_));
  NAND2_X1   g20920(.A1(new_n21176_), .A2(new_n21172_), .ZN(new_n21177_));
  XOR2_X1    g20921(.A1(new_n21177_), .A2(new_n21167_), .Z(\f[121] ));
  NOR3_X1    g20922(.A1(new_n21171_), .A2(new_n21138_), .A3(new_n21169_), .ZN(new_n21179_));
  AOI21_X1   g20923(.A1(new_n21167_), .A2(new_n21172_), .B(new_n21179_), .ZN(new_n21180_));
  OAI21_X1   g20924(.A1(new_n21145_), .A2(new_n21162_), .B(new_n21164_), .ZN(new_n21181_));
  AOI22_X1   g20925(.A1(new_n13460_), .A2(new_n10984_), .B1(\b[63] ), .B2(new_n12304_), .ZN(new_n21182_));
  NAND2_X1   g20926(.A1(new_n21153_), .A2(new_n21158_), .ZN(new_n21183_));
  NAND2_X1   g20927(.A1(new_n21183_), .A2(new_n21159_), .ZN(new_n21184_));
  AOI22_X1   g20928(.A1(new_n12922_), .A2(\b[59] ), .B1(\b[58] ), .B2(new_n12923_), .ZN(new_n21185_));
  INV_X1     g20929(.I(new_n21185_), .ZN(new_n21186_));
  NOR2_X1    g20930(.A1(new_n21186_), .A2(new_n21157_), .ZN(new_n21187_));
  NAND2_X1   g20931(.A1(new_n21186_), .A2(new_n21157_), .ZN(new_n21188_));
  INV_X1     g20932(.I(new_n21188_), .ZN(new_n21189_));
  NOR2_X1    g20933(.A1(new_n21189_), .A2(new_n21187_), .ZN(new_n21190_));
  XNOR2_X1   g20934(.A1(new_n21184_), .A2(new_n21190_), .ZN(new_n21191_));
  XOR2_X1    g20935(.A1(new_n21191_), .A2(new_n21182_), .Z(new_n21192_));
  AOI22_X1   g20936(.A1(new_n11926_), .A2(\b[62] ), .B1(new_n11924_), .B2(\b[61] ), .ZN(new_n21193_));
  OAI21_X1   g20937(.A1(new_n12147_), .A2(new_n12317_), .B(new_n21193_), .ZN(new_n21194_));
  AOI21_X1   g20938(.A1(new_n13444_), .A2(new_n11929_), .B(new_n21194_), .ZN(new_n21195_));
  XOR2_X1    g20939(.A1(new_n21195_), .A2(new_n12312_), .Z(new_n21196_));
  XOR2_X1    g20940(.A1(new_n21196_), .A2(new_n10989_), .Z(new_n21197_));
  XOR2_X1    g20941(.A1(new_n21192_), .A2(new_n21197_), .Z(new_n21198_));
  INV_X1     g20942(.I(new_n21198_), .ZN(new_n21199_));
  NAND2_X1   g20943(.A1(new_n21199_), .A2(new_n21181_), .ZN(new_n21200_));
  NOR2_X1    g20944(.A1(new_n21199_), .A2(new_n21181_), .ZN(new_n21201_));
  INV_X1     g20945(.I(new_n21201_), .ZN(new_n21202_));
  AND2_X2    g20946(.A1(new_n21202_), .A2(new_n21200_), .Z(new_n21203_));
  XOR2_X1    g20947(.A1(new_n21180_), .A2(new_n21203_), .Z(\f[122] ));
  NOR2_X1    g20948(.A1(new_n21191_), .A2(new_n21196_), .ZN(new_n21205_));
  NAND2_X1   g20949(.A1(new_n21191_), .A2(new_n21196_), .ZN(new_n21206_));
  XOR2_X1    g20950(.A1(new_n21182_), .A2(new_n10989_), .Z(new_n21207_));
  INV_X1     g20951(.I(new_n21207_), .ZN(new_n21208_));
  AOI21_X1   g20952(.A1(new_n21206_), .A2(new_n21208_), .B(new_n21205_), .ZN(new_n21209_));
  INV_X1     g20953(.I(new_n21187_), .ZN(new_n21210_));
  AOI21_X1   g20954(.A1(new_n21184_), .A2(new_n21210_), .B(new_n21189_), .ZN(new_n21211_));
  AOI22_X1   g20955(.A1(new_n11926_), .A2(\b[63] ), .B1(new_n11924_), .B2(\b[62] ), .ZN(new_n21212_));
  OAI21_X1   g20956(.A1(new_n12148_), .A2(new_n12317_), .B(new_n21212_), .ZN(new_n21213_));
  AOI21_X1   g20957(.A1(new_n12811_), .A2(new_n11929_), .B(new_n21213_), .ZN(new_n21214_));
  XOR2_X1    g20958(.A1(new_n21214_), .A2(new_n12312_), .Z(new_n21215_));
  INV_X1     g20959(.I(new_n21215_), .ZN(new_n21216_));
  AOI22_X1   g20960(.A1(new_n12922_), .A2(\b[60] ), .B1(\b[59] ), .B2(new_n12923_), .ZN(new_n21217_));
  INV_X1     g20961(.I(new_n21217_), .ZN(new_n21218_));
  NOR2_X1    g20962(.A1(new_n21218_), .A2(new_n10989_), .ZN(new_n21219_));
  NOR2_X1    g20963(.A1(new_n21217_), .A2(\a[59] ), .ZN(new_n21220_));
  NOR2_X1    g20964(.A1(new_n21219_), .A2(new_n21220_), .ZN(new_n21221_));
  XOR2_X1    g20965(.A1(new_n21221_), .A2(new_n21185_), .Z(new_n21222_));
  NOR2_X1    g20966(.A1(new_n21216_), .A2(new_n21222_), .ZN(new_n21223_));
  NAND2_X1   g20967(.A1(new_n21216_), .A2(new_n21222_), .ZN(new_n21224_));
  INV_X1     g20968(.I(new_n21224_), .ZN(new_n21225_));
  NOR2_X1    g20969(.A1(new_n21225_), .A2(new_n21223_), .ZN(new_n21226_));
  XOR2_X1    g20970(.A1(new_n21226_), .A2(new_n21211_), .Z(new_n21227_));
  NAND2_X1   g20971(.A1(new_n21209_), .A2(new_n21227_), .ZN(new_n21228_));
  INV_X1     g20972(.I(new_n21228_), .ZN(new_n21229_));
  NOR2_X1    g20973(.A1(new_n21209_), .A2(new_n21227_), .ZN(new_n21230_));
  NOR2_X1    g20974(.A1(new_n21229_), .A2(new_n21230_), .ZN(new_n21231_));
  INV_X1     g20975(.I(new_n21231_), .ZN(new_n21232_));
  AOI21_X1   g20976(.A1(new_n21180_), .A2(new_n21203_), .B(new_n21201_), .ZN(new_n21233_));
  XOR2_X1    g20977(.A1(new_n21233_), .A2(new_n21232_), .Z(\f[123] ));
  OAI21_X1   g20978(.A1(new_n21211_), .A2(new_n21223_), .B(new_n21224_), .ZN(new_n21235_));
  OAI22_X1   g20979(.A1(new_n12317_), .A2(new_n12796_), .B1(new_n11923_), .B2(new_n12800_), .ZN(new_n21236_));
  AOI21_X1   g20980(.A1(new_n13973_), .A2(new_n11929_), .B(new_n21236_), .ZN(new_n21237_));
  XOR2_X1    g20981(.A1(new_n21237_), .A2(\a[62] ), .Z(new_n21238_));
  NOR2_X1    g20982(.A1(new_n21220_), .A2(new_n21186_), .ZN(new_n21239_));
  NOR2_X1    g20983(.A1(new_n21239_), .A2(new_n21219_), .ZN(new_n21240_));
  AOI22_X1   g20984(.A1(new_n12922_), .A2(\b[61] ), .B1(\b[60] ), .B2(new_n12923_), .ZN(new_n21241_));
  NAND2_X1   g20985(.A1(new_n21240_), .A2(new_n21241_), .ZN(new_n21242_));
  NOR2_X1    g20986(.A1(new_n21240_), .A2(new_n21241_), .ZN(new_n21243_));
  INV_X1     g20987(.I(new_n21243_), .ZN(new_n21244_));
  NAND2_X1   g20988(.A1(new_n21244_), .A2(new_n21242_), .ZN(new_n21245_));
  XNOR2_X1   g20989(.A1(new_n21238_), .A2(new_n21245_), .ZN(new_n21246_));
  INV_X1     g20990(.I(new_n21246_), .ZN(new_n21247_));
  OAI21_X1   g20991(.A1(new_n21233_), .A2(new_n21232_), .B(new_n21228_), .ZN(new_n21248_));
  NAND2_X1   g20992(.A1(new_n21248_), .A2(new_n21247_), .ZN(new_n21249_));
  AOI21_X1   g20993(.A1(new_n21175_), .A2(new_n21139_), .B(new_n21168_), .ZN(new_n21250_));
  OAI21_X1   g20994(.A1(new_n21166_), .A2(new_n21250_), .B(new_n21176_), .ZN(new_n21251_));
  INV_X1     g20995(.I(new_n21203_), .ZN(new_n21252_));
  OAI21_X1   g20996(.A1(new_n21251_), .A2(new_n21252_), .B(new_n21202_), .ZN(new_n21253_));
  AOI21_X1   g20997(.A1(new_n21253_), .A2(new_n21231_), .B(new_n21229_), .ZN(new_n21254_));
  NAND2_X1   g20998(.A1(new_n21254_), .A2(new_n21246_), .ZN(new_n21255_));
  NAND2_X1   g20999(.A1(new_n21255_), .A2(new_n21249_), .ZN(new_n21256_));
  XOR2_X1    g21000(.A1(new_n21256_), .A2(new_n21235_), .Z(\f[124] ));
  NOR2_X1    g21001(.A1(new_n21248_), .A2(new_n21247_), .ZN(new_n21258_));
  INV_X1     g21002(.I(new_n21235_), .ZN(new_n21259_));
  AOI21_X1   g21003(.A1(new_n21248_), .A2(new_n21247_), .B(new_n21259_), .ZN(new_n21260_));
  NOR2_X1    g21004(.A1(new_n21260_), .A2(new_n21258_), .ZN(new_n21261_));
  AOI21_X1   g21005(.A1(new_n21238_), .A2(new_n21242_), .B(new_n21243_), .ZN(new_n21262_));
  INV_X1     g21006(.I(new_n21262_), .ZN(new_n21263_));
  INV_X1     g21007(.I(new_n21241_), .ZN(new_n21264_));
  AOI22_X1   g21008(.A1(new_n13460_), .A2(new_n11929_), .B1(\b[63] ), .B2(new_n13223_), .ZN(new_n21265_));
  XOR2_X1    g21009(.A1(new_n21265_), .A2(new_n21264_), .Z(new_n21266_));
  AOI22_X1   g21010(.A1(new_n12922_), .A2(\b[62] ), .B1(\b[61] ), .B2(new_n12923_), .ZN(new_n21267_));
  XOR2_X1    g21011(.A1(new_n21267_), .A2(new_n12312_), .Z(new_n21268_));
  XOR2_X1    g21012(.A1(new_n21265_), .A2(new_n21241_), .Z(new_n21269_));
  MUX2_X1    g21013(.I0(new_n21269_), .I1(new_n21266_), .S(new_n21268_), .Z(new_n21270_));
  NOR2_X1    g21014(.A1(new_n21263_), .A2(new_n21270_), .ZN(new_n21271_));
  NAND2_X1   g21015(.A1(new_n21263_), .A2(new_n21270_), .ZN(new_n21272_));
  INV_X1     g21016(.I(new_n21272_), .ZN(new_n21273_));
  NOR2_X1    g21017(.A1(new_n21273_), .A2(new_n21271_), .ZN(new_n21274_));
  XOR2_X1    g21018(.A1(new_n21261_), .A2(new_n21274_), .Z(\f[125] ));
  INV_X1     g21019(.I(new_n21271_), .ZN(new_n21276_));
  OAI21_X1   g21020(.A1(new_n21260_), .A2(new_n21258_), .B(new_n21276_), .ZN(new_n21277_));
  NAND2_X1   g21021(.A1(new_n21277_), .A2(new_n21272_), .ZN(new_n21278_));
  INV_X1     g21022(.I(new_n21267_), .ZN(new_n21279_));
  NOR2_X1    g21023(.A1(new_n21265_), .A2(new_n12312_), .ZN(new_n21280_));
  INV_X1     g21024(.I(new_n21280_), .ZN(new_n21281_));
  NAND2_X1   g21025(.A1(new_n21265_), .A2(new_n12312_), .ZN(new_n21282_));
  AOI22_X1   g21026(.A1(new_n21281_), .A2(new_n21282_), .B1(new_n21241_), .B2(new_n21279_), .ZN(new_n21283_));
  AOI21_X1   g21027(.A1(new_n21264_), .A2(new_n21267_), .B(new_n21283_), .ZN(new_n21284_));
  INV_X1     g21028(.I(new_n21284_), .ZN(new_n21285_));
  AOI22_X1   g21029(.A1(new_n12922_), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n12923_), .ZN(new_n21286_));
  NAND2_X1   g21030(.A1(new_n21286_), .A2(\a[62] ), .ZN(new_n21287_));
  NOR2_X1    g21031(.A1(new_n21286_), .A2(\a[62] ), .ZN(new_n21288_));
  INV_X1     g21032(.I(new_n21288_), .ZN(new_n21289_));
  NAND2_X1   g21033(.A1(new_n21289_), .A2(new_n21287_), .ZN(new_n21290_));
  XOR2_X1    g21034(.A1(new_n21290_), .A2(new_n21264_), .Z(new_n21291_));
  NOR2_X1    g21035(.A1(new_n21285_), .A2(new_n21291_), .ZN(new_n21292_));
  NAND2_X1   g21036(.A1(new_n21285_), .A2(new_n21291_), .ZN(new_n21293_));
  INV_X1     g21037(.I(new_n21293_), .ZN(new_n21294_));
  NOR2_X1    g21038(.A1(new_n21294_), .A2(new_n21292_), .ZN(new_n21295_));
  INV_X1     g21039(.I(new_n21295_), .ZN(new_n21296_));
  XOR2_X1    g21040(.A1(new_n21278_), .A2(new_n21296_), .Z(\f[126] ));
  INV_X1     g21041(.I(new_n21292_), .ZN(new_n21298_));
  NAND3_X1   g21042(.A1(new_n21277_), .A2(new_n21272_), .A3(new_n21293_), .ZN(new_n21299_));
  NAND2_X1   g21043(.A1(new_n12923_), .A2(\b[63] ), .ZN(new_n21300_));
  OAI21_X1   g21044(.A1(new_n21264_), .A2(new_n21288_), .B(new_n21287_), .ZN(new_n21301_));
  XNOR2_X1   g21045(.A1(new_n21301_), .A2(new_n21300_), .ZN(new_n21302_));
  NAND3_X1   g21046(.A1(new_n21299_), .A2(new_n21298_), .A3(new_n21302_), .ZN(new_n21303_));
  OAI21_X1   g21047(.A1(new_n21254_), .A2(new_n21246_), .B(new_n21235_), .ZN(new_n21304_));
  AOI21_X1   g21048(.A1(new_n21304_), .A2(new_n21255_), .B(new_n21271_), .ZN(new_n21305_));
  NOR3_X1    g21049(.A1(new_n21305_), .A2(new_n21273_), .A3(new_n21294_), .ZN(new_n21306_));
  INV_X1     g21050(.I(new_n21302_), .ZN(new_n21307_));
  OAI21_X1   g21051(.A1(new_n21306_), .A2(new_n21292_), .B(new_n21307_), .ZN(new_n21308_));
  NAND2_X1   g21052(.A1(new_n21308_), .A2(new_n21303_), .ZN(\f[127] ));
endmodule


