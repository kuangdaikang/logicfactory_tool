// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:43 2022

module x6dn  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
    v30, v31, v32, v33, v34, v35, v36, v37, v38,
    \v39.0 , \v39.1 , \v39.2 , \v39.3 , \v39.4   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28,
    v29, v30, v31, v32, v33, v34, v35, v36, v37, v38;
  output \v39.0 , \v39.1 , \v39.2 , \v39.3 , \v39.4 ;
  wire new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_;
  assign new_n45_ = ~v9 & ~v10;
  assign new_n46_ = ~v11 & v12;
  assign new_n47_ = new_n45_ & new_n46_;
  assign new_n48_ = ~v9 & ~new_n47_;
  assign new_n49_ = ~v8 & ~new_n48_;
  assign new_n50_ = ~v8 & v9;
  assign new_n51_ = ~v13 & ~new_n50_;
  assign new_n52_ = ~v11 & new_n51_;
  assign new_n53_ = v10 & new_n52_;
  assign new_n54_ = ~new_n49_ & ~new_n53_;
  assign new_n55_ = v7 & ~new_n54_;
  assign new_n56_ = v7 & ~new_n55_;
  assign new_n57_ = v6 & ~new_n56_;
  assign new_n58_ = ~v2 & new_n57_;
  assign new_n59_ = v17 & v19;
  assign new_n60_ = v16 & ~new_n59_;
  assign new_n61_ = ~v17 & ~v19;
  assign new_n62_ = ~v16 & ~new_n61_;
  assign new_n63_ = ~v17 & v19;
  assign new_n64_ = v17 & ~v19;
  assign new_n65_ = v25 & ~new_n64_;
  assign new_n66_ = ~new_n63_ & new_n65_;
  assign new_n67_ = ~new_n62_ & new_n66_;
  assign new_n68_ = ~new_n60_ & new_n67_;
  assign new_n69_ = v14 & ~new_n68_;
  assign new_n70_ = v2 & new_n69_;
  assign new_n71_ = ~new_n58_ & ~new_n70_;
  assign new_n72_ = ~v4 & ~new_n71_;
  assign new_n73_ = v22 & v23;
  assign new_n74_ = v19 & ~v20;
  assign new_n75_ = v18 & new_n74_;
  assign new_n76_ = v21 & ~new_n75_;
  assign new_n77_ = ~new_n73_ & ~new_n76_;
  assign new_n78_ = ~v17 & new_n77_;
  assign new_n79_ = ~v13 & v17;
  assign new_n80_ = ~new_n78_ & ~new_n79_;
  assign new_n81_ = v2 & ~new_n80_;
  assign new_n82_ = ~v2 & v16;
  assign new_n83_ = ~new_n81_ & ~new_n82_;
  assign new_n84_ = ~v14 & ~new_n83_;
  assign new_n85_ = v4 & new_n84_;
  assign new_n86_ = ~new_n72_ & ~new_n85_;
  assign new_n87_ = ~v3 & ~new_n86_;
  assign new_n88_ = v27 & v28;
  assign new_n89_ = ~new_n73_ & ~new_n88_;
  assign new_n90_ = v26 & new_n89_;
  assign new_n91_ = v19 & new_n90_;
  assign new_n92_ = v14 & new_n91_;
  assign new_n93_ = ~v2 & new_n92_;
  assign new_n94_ = v2 & ~v14;
  assign new_n95_ = ~new_n93_ & ~new_n94_;
  assign new_n96_ = v4 & ~new_n95_;
  assign new_n97_ = v3 & new_n96_;
  assign new_n98_ = ~new_n87_ & ~new_n97_;
  assign new_n99_ = ~v0 & ~new_n98_;
  assign new_n100_ = ~v3 & v4;
  assign new_n101_ = v3 & ~v4;
  assign new_n102_ = ~new_n100_ & ~new_n101_;
  assign new_n103_ = ~v2 & ~new_n102_;
  assign new_n104_ = ~v22 & ~v23;
  assign new_n105_ = ~v23 & ~new_n104_;
  assign new_n106_ = ~v22 & new_n105_;
  assign new_n107_ = v3 & ~new_n106_;
  assign new_n108_ = v3 & ~new_n107_;
  assign new_n109_ = v2 & ~new_n108_;
  assign new_n110_ = ~new_n103_ & ~new_n109_;
  assign new_n111_ = v0 & ~new_n110_;
  assign new_n112_ = v17 & ~v20;
  assign new_n113_ = v21 & ~new_n112_;
  assign new_n114_ = v4 & ~new_n113_;
  assign new_n115_ = v3 & new_n114_;
  assign new_n116_ = ~v2 & new_n115_;
  assign new_n117_ = ~new_n111_ & ~new_n116_;
  assign new_n118_ = ~v14 & ~new_n117_;
  assign new_n119_ = v0 & ~v2;
  assign new_n120_ = v3 & v14;
  assign new_n121_ = new_n119_ & new_n120_;
  assign new_n122_ = ~new_n118_ & ~new_n121_;
  assign new_n123_ = ~new_n99_ & new_n122_;
  assign new_n124_ = ~v5 & ~new_n123_;
  assign new_n125_ = ~v4 & v14;
  assign new_n126_ = v0 & new_n125_;
  assign new_n127_ = v4 & v5;
  assign new_n128_ = ~v0 & new_n127_;
  assign new_n129_ = v23 & ~v24;
  assign new_n130_ = ~v14 & new_n129_;
  assign new_n131_ = new_n128_ & new_n130_;
  assign new_n132_ = ~new_n126_ & ~new_n131_;
  assign new_n133_ = ~v3 & ~new_n132_;
  assign new_n134_ = v5 & ~v14;
  assign new_n135_ = v4 & new_n134_;
  assign new_n136_ = ~new_n125_ & ~new_n135_;
  assign new_n137_ = v0 & ~new_n136_;
  assign new_n138_ = ~v14 & v17;
  assign new_n139_ = ~v13 & new_n138_;
  assign new_n140_ = new_n128_ & new_n139_;
  assign new_n141_ = ~new_n137_ & ~new_n140_;
  assign new_n142_ = ~new_n104_ & ~new_n141_;
  assign new_n143_ = ~v14 & new_n104_;
  assign new_n144_ = ~v14 & ~new_n143_;
  assign new_n145_ = v5 & ~new_n144_;
  assign new_n146_ = v4 & new_n145_;
  assign new_n147_ = new_n104_ & new_n125_;
  assign new_n148_ = ~new_n146_ & ~new_n147_;
  assign new_n149_ = v0 & ~new_n148_;
  assign new_n150_ = ~v4 & new_n134_;
  assign new_n151_ = v18 & ~v20;
  assign new_n152_ = ~v17 & new_n151_;
  assign new_n153_ = new_n150_ & new_n152_;
  assign new_n154_ = ~new_n149_ & ~new_n153_;
  assign new_n155_ = ~new_n142_ & new_n154_;
  assign new_n156_ = v3 & ~new_n155_;
  assign new_n157_ = ~new_n133_ & ~new_n156_;
  assign new_n158_ = v2 & ~new_n157_;
  assign new_n159_ = ~v2 & v4;
  assign new_n160_ = ~v4 & v5;
  assign new_n161_ = ~new_n159_ & ~new_n160_;
  assign new_n162_ = v3 & ~new_n161_;
  assign new_n163_ = ~v3 & new_n127_;
  assign new_n164_ = ~new_n162_ & ~new_n163_;
  assign new_n165_ = ~v14 & ~new_n164_;
  assign new_n166_ = v4 & v14;
  assign new_n167_ = v4 & ~new_n166_;
  assign new_n168_ = ~v3 & ~new_n167_;
  assign new_n169_ = ~v2 & new_n168_;
  assign new_n170_ = ~new_n165_ & ~new_n169_;
  assign new_n171_ = v0 & ~new_n170_;
  assign new_n172_ = ~new_n158_ & ~new_n171_;
  assign new_n173_ = ~new_n124_ & new_n172_;
  assign \v39.0  = v1 & ~new_n173_;
  assign new_n175_ = ~v11 & v13;
  assign new_n176_ = ~v9 & new_n175_;
  assign new_n177_ = ~v11 & ~new_n176_;
  assign new_n178_ = v8 & ~new_n177_;
  assign new_n179_ = ~v9 & v11;
  assign new_n180_ = ~new_n178_ & ~new_n179_;
  assign new_n181_ = v10 & ~new_n180_;
  assign new_n182_ = v10 & ~new_n175_;
  assign new_n183_ = v8 & ~new_n182_;
  assign new_n184_ = v8 & ~new_n183_;
  assign new_n185_ = v9 & ~new_n184_;
  assign new_n186_ = ~new_n181_ & ~new_n185_;
  assign new_n187_ = v7 & ~new_n186_;
  assign new_n188_ = v7 & ~new_n187_;
  assign new_n189_ = v6 & ~new_n188_;
  assign new_n190_ = ~v4 & new_n189_;
  assign new_n191_ = ~v14 & v16;
  assign new_n192_ = v4 & new_n191_;
  assign new_n193_ = ~new_n190_ & ~new_n192_;
  assign new_n194_ = ~v3 & ~new_n193_;
  assign new_n195_ = v19 & v34;
  assign new_n196_ = v34 & ~new_n195_;
  assign new_n197_ = ~new_n112_ & ~new_n196_;
  assign new_n198_ = v21 & new_n197_;
  assign new_n199_ = ~v14 & new_n198_;
  assign new_n200_ = v26 & ~new_n73_;
  assign new_n201_ = v19 & new_n200_;
  assign new_n202_ = ~new_n73_ & ~new_n201_;
  assign new_n203_ = ~new_n88_ & ~new_n202_;
  assign new_n204_ = v14 & new_n203_;
  assign new_n205_ = ~new_n199_ & ~new_n204_;
  assign new_n206_ = v4 & ~new_n205_;
  assign new_n207_ = v14 & v19;
  assign new_n208_ = new_n88_ & new_n207_;
  assign new_n209_ = ~new_n206_ & ~new_n208_;
  assign new_n210_ = v3 & ~new_n209_;
  assign new_n211_ = ~new_n194_ & ~new_n210_;
  assign new_n212_ = ~v2 & ~new_n211_;
  assign new_n213_ = ~v4 & new_n69_;
  assign new_n214_ = ~v14 & new_n78_;
  assign new_n215_ = v4 & new_n214_;
  assign new_n216_ = ~new_n213_ & ~new_n215_;
  assign new_n217_ = ~v3 & ~new_n216_;
  assign new_n218_ = v2 & new_n217_;
  assign new_n219_ = ~new_n212_ & ~new_n218_;
  assign new_n220_ = ~v0 & ~new_n219_;
  assign new_n221_ = v0 & ~new_n102_;
  assign new_n222_ = ~v4 & v29;
  assign new_n223_ = ~v3 & new_n222_;
  assign new_n224_ = v30 & v31;
  assign new_n225_ = ~v32 & v33;
  assign new_n226_ = new_n224_ & new_n225_;
  assign new_n227_ = new_n223_ & new_n226_;
  assign new_n228_ = ~new_n115_ & ~new_n227_;
  assign new_n229_ = ~new_n221_ & new_n228_;
  assign new_n230_ = ~v2 & ~new_n229_;
  assign new_n231_ = v0 & new_n109_;
  assign new_n232_ = ~new_n230_ & ~new_n231_;
  assign new_n233_ = ~v14 & ~new_n232_;
  assign new_n234_ = ~new_n121_ & ~new_n233_;
  assign new_n235_ = ~new_n220_ & new_n234_;
  assign new_n236_ = ~v5 & ~new_n235_;
  assign new_n237_ = ~new_n106_ & ~new_n136_;
  assign new_n238_ = v5 & v14;
  assign new_n239_ = v4 & new_n238_;
  assign new_n240_ = ~new_n237_ & ~new_n239_;
  assign new_n241_ = v2 & ~new_n240_;
  assign new_n242_ = ~v14 & ~new_n161_;
  assign new_n243_ = ~new_n241_ & ~new_n242_;
  assign new_n244_ = v3 & ~new_n243_;
  assign new_n245_ = ~v2 & ~new_n167_;
  assign new_n246_ = v2 & new_n125_;
  assign new_n247_ = ~new_n135_ & ~new_n246_;
  assign new_n248_ = ~new_n245_ & new_n247_;
  assign new_n249_ = ~v3 & ~new_n248_;
  assign new_n250_ = ~new_n244_ & ~new_n249_;
  assign new_n251_ = v0 & ~new_n250_;
  assign new_n252_ = v2 & ~v3;
  assign new_n253_ = new_n129_ & new_n252_;
  assign new_n254_ = ~v2 & v3;
  assign new_n255_ = v19 & v35;
  assign new_n256_ = new_n254_ & new_n255_;
  assign new_n257_ = ~new_n253_ & ~new_n256_;
  assign new_n258_ = v4 & ~new_n257_;
  assign new_n259_ = ~v0 & new_n258_;
  assign new_n260_ = v2 & new_n101_;
  assign new_n261_ = new_n152_ & new_n260_;
  assign new_n262_ = ~new_n259_ & ~new_n261_;
  assign new_n263_ = ~v14 & ~new_n262_;
  assign new_n264_ = ~v2 & ~v3;
  assign new_n265_ = ~v0 & new_n264_;
  assign new_n266_ = v14 & v16;
  assign new_n267_ = v4 & new_n266_;
  assign new_n268_ = new_n265_ & new_n267_;
  assign new_n269_ = ~new_n263_ & ~new_n268_;
  assign new_n270_ = v5 & ~new_n269_;
  assign new_n271_ = ~new_n251_ & ~new_n270_;
  assign new_n272_ = ~new_n236_ & new_n271_;
  assign \v39.1  = v1 & ~new_n272_;
  assign new_n274_ = v10 & ~v13;
  assign new_n275_ = ~v11 & ~new_n274_;
  assign new_n276_ = v8 & new_n275_;
  assign new_n277_ = v8 & ~new_n276_;
  assign new_n278_ = v9 & ~new_n277_;
  assign new_n279_ = v7 & new_n278_;
  assign new_n280_ = v6 & new_n279_;
  assign new_n281_ = ~v14 & v32;
  assign new_n282_ = ~new_n280_ & ~new_n281_;
  assign new_n283_ = ~v2 & ~new_n282_;
  assign new_n284_ = ~new_n70_ & ~new_n283_;
  assign new_n285_ = ~v4 & ~new_n284_;
  assign new_n286_ = ~v14 & ~new_n191_;
  assign new_n287_ = ~v2 & ~new_n286_;
  assign new_n288_ = v21 & v34;
  assign new_n289_ = v21 & ~new_n288_;
  assign new_n290_ = v23 & ~new_n289_;
  assign new_n291_ = v22 & new_n290_;
  assign new_n292_ = v34 & ~new_n75_;
  assign new_n293_ = v21 & new_n292_;
  assign new_n294_ = ~new_n291_ & ~new_n293_;
  assign new_n295_ = ~new_n77_ & new_n294_;
  assign new_n296_ = ~v17 & ~new_n295_;
  assign new_n297_ = v13 & v16;
  assign new_n298_ = new_n59_ & new_n297_;
  assign new_n299_ = ~new_n296_ & ~new_n298_;
  assign new_n300_ = ~v14 & ~new_n299_;
  assign new_n301_ = v2 & new_n300_;
  assign new_n302_ = ~new_n287_ & ~new_n301_;
  assign new_n303_ = v4 & ~new_n302_;
  assign new_n304_ = ~new_n285_ & ~new_n303_;
  assign new_n305_ = ~v3 & ~new_n304_;
  assign new_n306_ = v4 & new_n90_;
  assign new_n307_ = ~new_n88_ & ~new_n306_;
  assign new_n308_ = v19 & ~new_n307_;
  assign new_n309_ = v14 & new_n308_;
  assign new_n310_ = v3 & new_n309_;
  assign new_n311_ = ~v2 & new_n310_;
  assign new_n312_ = ~new_n305_ & ~new_n311_;
  assign new_n313_ = ~v0 & ~new_n312_;
  assign new_n314_ = v29 & new_n224_;
  assign new_n315_ = v33 & ~new_n314_;
  assign new_n316_ = ~v32 & new_n315_;
  assign new_n317_ = ~v4 & new_n316_;
  assign new_n318_ = ~v3 & new_n317_;
  assign new_n319_ = ~new_n115_ & ~new_n318_;
  assign new_n320_ = ~new_n221_ & new_n319_;
  assign new_n321_ = ~v2 & ~new_n320_;
  assign new_n322_ = ~new_n231_ & ~new_n321_;
  assign new_n323_ = ~v14 & ~new_n322_;
  assign new_n324_ = ~new_n121_ & ~new_n323_;
  assign new_n325_ = ~new_n313_ & new_n324_;
  assign new_n326_ = ~v5 & ~new_n325_;
  assign new_n327_ = v3 & ~v14;
  assign new_n328_ = new_n152_ & new_n327_;
  assign new_n329_ = ~v3 & v13;
  assign new_n330_ = ~v0 & new_n329_;
  assign new_n331_ = v17 & ~v37;
  assign new_n332_ = v14 & new_n331_;
  assign new_n333_ = new_n330_ & new_n332_;
  assign new_n334_ = ~new_n328_ & ~new_n333_;
  assign new_n335_ = ~v4 & ~new_n334_;
  assign new_n336_ = v35 & ~new_n129_;
  assign new_n337_ = v19 & new_n336_;
  assign new_n338_ = ~new_n129_ & ~new_n337_;
  assign new_n339_ = ~v3 & ~new_n338_;
  assign new_n340_ = ~v0 & new_n339_;
  assign new_n341_ = v0 & new_n107_;
  assign new_n342_ = ~new_n340_ & ~new_n341_;
  assign new_n343_ = ~v14 & ~new_n342_;
  assign new_n344_ = v0 & new_n120_;
  assign new_n345_ = ~new_n343_ & ~new_n344_;
  assign new_n346_ = v4 & ~new_n345_;
  assign new_n347_ = ~new_n335_ & ~new_n346_;
  assign new_n348_ = v5 & ~new_n347_;
  assign new_n349_ = v14 & ~new_n108_;
  assign new_n350_ = ~v4 & new_n349_;
  assign new_n351_ = v0 & new_n350_;
  assign new_n352_ = ~new_n348_ & ~new_n351_;
  assign new_n353_ = v2 & ~new_n352_;
  assign new_n354_ = ~v14 & v38;
  assign new_n355_ = new_n160_ & new_n354_;
  assign new_n356_ = new_n265_ & new_n355_;
  assign new_n357_ = ~new_n171_ & ~new_n356_;
  assign new_n358_ = ~new_n353_ & new_n357_;
  assign new_n359_ = ~new_n326_ & new_n358_;
  assign \v39.2  = v1 & ~new_n359_;
  assign new_n361_ = ~v10 & v11;
  assign new_n362_ = ~v11 & ~v13;
  assign new_n363_ = v10 & new_n362_;
  assign new_n364_ = ~new_n361_ & ~new_n363_;
  assign new_n365_ = ~new_n50_ & ~new_n364_;
  assign new_n366_ = ~v9 & ~v11;
  assign new_n367_ = v8 & new_n366_;
  assign new_n368_ = ~new_n50_ & ~new_n367_;
  assign new_n369_ = ~new_n365_ & new_n368_;
  assign new_n370_ = v7 & ~new_n369_;
  assign new_n371_ = v6 & new_n370_;
  assign new_n372_ = ~new_n281_ & ~new_n371_;
  assign new_n373_ = ~v2 & ~new_n372_;
  assign new_n374_ = ~new_n70_ & ~new_n373_;
  assign new_n375_ = ~v4 & ~new_n374_;
  assign new_n376_ = ~new_n85_ & ~new_n375_;
  assign new_n377_ = ~v3 & ~new_n376_;
  assign new_n378_ = v4 & new_n201_;
  assign new_n379_ = v4 & ~new_n378_;
  assign new_n380_ = ~new_n88_ & ~new_n379_;
  assign new_n381_ = ~v4 & new_n88_;
  assign new_n382_ = ~new_n380_ & ~new_n381_;
  assign new_n383_ = v14 & ~new_n382_;
  assign new_n384_ = v3 & new_n383_;
  assign new_n385_ = ~v2 & new_n384_;
  assign new_n386_ = ~new_n377_ & ~new_n385_;
  assign new_n387_ = ~v0 & ~new_n386_;
  assign new_n388_ = v0 & v3;
  assign new_n389_ = v29 & v30;
  assign new_n390_ = ~v3 & new_n389_;
  assign new_n391_ = v31 & new_n225_;
  assign new_n392_ = new_n390_ & new_n391_;
  assign new_n393_ = ~new_n388_ & ~new_n392_;
  assign new_n394_ = ~v2 & ~new_n393_;
  assign new_n395_ = ~new_n252_ & ~new_n394_;
  assign new_n396_ = ~v4 & ~new_n395_;
  assign new_n397_ = ~v2 & new_n114_;
  assign new_n398_ = v2 & ~new_n106_;
  assign new_n399_ = v0 & new_n398_;
  assign new_n400_ = ~new_n397_ & ~new_n399_;
  assign new_n401_ = v3 & ~new_n400_;
  assign new_n402_ = ~new_n396_ & ~new_n401_;
  assign new_n403_ = ~v14 & ~new_n402_;
  assign new_n404_ = ~new_n121_ & ~new_n403_;
  assign new_n405_ = ~new_n387_ & new_n404_;
  assign new_n406_ = ~v5 & ~new_n405_;
  assign new_n407_ = v4 & ~v14;
  assign new_n408_ = new_n129_ & new_n407_;
  assign new_n409_ = new_n125_ & new_n331_;
  assign new_n410_ = ~new_n408_ & ~new_n409_;
  assign new_n411_ = ~v3 & ~new_n410_;
  assign new_n412_ = ~v14 & ~new_n152_;
  assign new_n413_ = ~v4 & new_n412_;
  assign new_n414_ = v3 & new_n413_;
  assign new_n415_ = ~new_n411_ & ~new_n414_;
  assign new_n416_ = ~v0 & ~new_n415_;
  assign new_n417_ = ~v14 & ~new_n106_;
  assign new_n418_ = ~v14 & ~new_n417_;
  assign new_n419_ = v4 & ~new_n418_;
  assign new_n420_ = v0 & new_n419_;
  assign new_n421_ = ~v4 & ~v14;
  assign new_n422_ = new_n152_ & new_n421_;
  assign new_n423_ = ~new_n420_ & ~new_n422_;
  assign new_n424_ = v3 & ~new_n423_;
  assign new_n425_ = ~new_n416_ & ~new_n424_;
  assign new_n426_ = v5 & ~new_n425_;
  assign new_n427_ = ~new_n125_ & ~new_n407_;
  assign new_n428_ = ~v3 & ~new_n427_;
  assign new_n429_ = v14 & ~new_n106_;
  assign new_n430_ = ~v4 & new_n429_;
  assign new_n431_ = v3 & new_n430_;
  assign new_n432_ = ~new_n428_ & ~new_n431_;
  assign new_n433_ = v0 & ~new_n432_;
  assign new_n434_ = ~new_n426_ & ~new_n433_;
  assign new_n435_ = v2 & ~new_n434_;
  assign new_n436_ = ~new_n168_ & ~new_n407_;
  assign new_n437_ = ~v2 & ~new_n436_;
  assign new_n438_ = new_n101_ & new_n134_;
  assign new_n439_ = ~new_n437_ & ~new_n438_;
  assign new_n440_ = v0 & ~new_n439_;
  assign new_n441_ = ~new_n356_ & ~new_n440_;
  assign new_n442_ = ~new_n435_ & new_n441_;
  assign new_n443_ = ~new_n406_ & new_n442_;
  assign \v39.3  = v1 & ~new_n443_;
  assign new_n445_ = ~v9 & v10;
  assign new_n446_ = ~v9 & ~new_n445_;
  assign new_n447_ = v13 & ~new_n446_;
  assign new_n448_ = v10 & ~new_n447_;
  assign new_n449_ = ~v11 & ~new_n448_;
  assign new_n450_ = v8 & new_n449_;
  assign new_n451_ = ~new_n49_ & ~new_n450_;
  assign new_n452_ = v7 & ~new_n451_;
  assign new_n453_ = v6 & new_n452_;
  assign new_n454_ = ~v2 & new_n453_;
  assign new_n455_ = v16 & new_n59_;
  assign new_n456_ = ~v16 & new_n61_;
  assign new_n457_ = ~new_n455_ & ~new_n456_;
  assign new_n458_ = v25 & ~new_n457_;
  assign new_n459_ = new_n68_ & ~new_n458_;
  assign new_n460_ = v14 & ~new_n459_;
  assign new_n461_ = v2 & new_n460_;
  assign new_n462_ = ~new_n454_ & ~new_n461_;
  assign new_n463_ = ~v4 & ~new_n462_;
  assign new_n464_ = ~v16 & v36;
  assign new_n465_ = ~v16 & ~new_n464_;
  assign new_n466_ = v17 & ~new_n465_;
  assign new_n467_ = v13 & new_n466_;
  assign new_n468_ = v18 & v19;
  assign new_n469_ = ~v20 & ~new_n73_;
  assign new_n470_ = new_n468_ & new_n469_;
  assign new_n471_ = v34 & ~new_n470_;
  assign new_n472_ = v21 & new_n471_;
  assign new_n473_ = ~new_n77_ & ~new_n472_;
  assign new_n474_ = ~v17 & ~new_n473_;
  assign new_n475_ = ~new_n467_ & ~new_n474_;
  assign new_n476_ = v2 & ~new_n475_;
  assign new_n477_ = ~new_n82_ & ~new_n476_;
  assign new_n478_ = ~v14 & ~new_n477_;
  assign new_n479_ = v4 & new_n478_;
  assign new_n480_ = ~new_n463_ & ~new_n479_;
  assign new_n481_ = ~v3 & ~new_n480_;
  assign new_n482_ = v34 & ~new_n112_;
  assign new_n483_ = v21 & new_n482_;
  assign new_n484_ = ~v14 & new_n483_;
  assign new_n485_ = v19 & v26;
  assign new_n486_ = v26 & ~new_n485_;
  assign new_n487_ = v19 & new_n486_;
  assign new_n488_ = ~new_n73_ & ~new_n487_;
  assign new_n489_ = ~new_n88_ & new_n488_;
  assign new_n490_ = ~new_n88_ & ~new_n489_;
  assign new_n491_ = v14 & ~new_n490_;
  assign new_n492_ = ~new_n484_ & ~new_n491_;
  assign new_n493_ = v4 & ~new_n492_;
  assign new_n494_ = ~v2 & new_n493_;
  assign new_n495_ = v14 & ~new_n88_;
  assign new_n496_ = v14 & ~new_n495_;
  assign new_n497_ = v36 & ~new_n496_;
  assign new_n498_ = v2 & new_n497_;
  assign new_n499_ = v14 & new_n88_;
  assign new_n500_ = ~new_n498_ & ~new_n499_;
  assign new_n501_ = ~v4 & ~new_n500_;
  assign new_n502_ = ~new_n494_ & ~new_n501_;
  assign new_n503_ = v3 & ~new_n502_;
  assign new_n504_ = ~new_n481_ & ~new_n503_;
  assign new_n505_ = ~v0 & ~new_n504_;
  assign new_n506_ = ~v3 & new_n407_;
  assign new_n507_ = ~new_n120_ & ~new_n506_;
  assign new_n508_ = ~v2 & ~new_n507_;
  assign new_n509_ = v3 & ~new_n104_;
  assign new_n510_ = v3 & ~new_n509_;
  assign new_n511_ = ~v14 & ~new_n510_;
  assign new_n512_ = v2 & new_n511_;
  assign new_n513_ = ~new_n508_ & ~new_n512_;
  assign new_n514_ = v0 & ~new_n513_;
  assign new_n515_ = new_n254_ & new_n421_;
  assign new_n516_ = ~new_n514_ & ~new_n515_;
  assign new_n517_ = ~new_n505_ & new_n516_;
  assign new_n518_ = ~v5 & ~new_n517_;
  assign new_n519_ = ~new_n104_ & ~new_n136_;
  assign new_n520_ = ~new_n166_ & ~new_n421_;
  assign new_n521_ = v5 & ~new_n520_;
  assign new_n522_ = ~new_n519_ & ~new_n521_;
  assign new_n523_ = v3 & ~new_n522_;
  assign new_n524_ = ~v3 & new_n125_;
  assign new_n525_ = ~new_n523_ & ~new_n524_;
  assign new_n526_ = v0 & ~new_n525_;
  assign new_n527_ = v36 & v37;
  assign new_n528_ = v13 & new_n331_;
  assign new_n529_ = ~new_n527_ & ~new_n528_;
  assign new_n530_ = v14 & ~new_n529_;
  assign new_n531_ = ~v4 & new_n530_;
  assign new_n532_ = ~new_n408_ & ~new_n531_;
  assign new_n533_ = ~v3 & ~new_n532_;
  assign new_n534_ = ~v0 & new_n533_;
  assign new_n535_ = v3 & new_n421_;
  assign new_n536_ = new_n152_ & new_n535_;
  assign new_n537_ = ~new_n534_ & ~new_n536_;
  assign new_n538_ = v5 & ~new_n537_;
  assign new_n539_ = ~new_n526_ & ~new_n538_;
  assign new_n540_ = v2 & ~new_n539_;
  assign new_n541_ = ~v2 & v14;
  assign new_n542_ = ~new_n134_ & ~new_n541_;
  assign new_n543_ = v0 & ~new_n542_;
  assign new_n544_ = ~v2 & v5;
  assign new_n545_ = ~v0 & new_n544_;
  assign new_n546_ = v14 & new_n464_;
  assign new_n547_ = new_n545_ & new_n546_;
  assign new_n548_ = ~new_n543_ & ~new_n547_;
  assign new_n549_ = v4 & ~new_n548_;
  assign new_n550_ = ~v2 & ~v4;
  assign new_n551_ = v0 & new_n550_;
  assign new_n552_ = ~new_n549_ & ~new_n551_;
  assign new_n553_ = ~v3 & ~new_n552_;
  assign new_n554_ = ~new_n540_ & ~new_n553_;
  assign new_n555_ = ~new_n518_ & new_n554_;
  assign \v39.4  = v1 & ~new_n555_;
endmodule


