// Benchmark "source.pla" written by ABC on Fri Feb 25 15:13:04 2022

module xparc  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
    v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40,
    \v41.0 , \v41.1 , \v41.2 , \v41.3 , \v41.4 , \v41.5 , \v41.6 , \v41.7 ,
    \v41.8 , \v41.9 , \v41.10 , \v41.11 , \v41.12 , \v41.13 , \v41.14 ,
    \v41.15 , \v41.16 , \v41.17 , \v41.18 , \v41.19 , \v41.20 , \v41.21 ,
    \v41.22 , \v41.23 , \v41.24 , \v41.25 , \v41.26 , \v41.27 , \v41.28 ,
    \v41.29 , \v41.30 , \v41.31 , \v41.32 , \v41.33 , \v41.34 , \v41.35 ,
    \v41.36 , \v41.37 , \v41.38 , \v41.39 , \v41.40 , \v41.41 , \v41.42 ,
    \v41.43 , \v41.44 , \v41.45 , \v41.46 , \v41.47 , \v41.48 , \v41.49 ,
    \v41.50 , \v41.51 , \v41.52 , \v41.53 , \v41.54 , \v41.55 , \v41.56 ,
    \v41.57 , \v41.58 , \v41.59 , \v41.60 , \v41.61 , \v41.62 , \v41.63 ,
    \v41.64 , \v41.65 , \v41.66 , \v41.67 , \v41.68 , \v41.69 , \v41.70 ,
    \v41.71 , \v41.72   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28,
    v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40;
  output \v41.0 , \v41.1 , \v41.2 , \v41.3 , \v41.4 , \v41.5 , \v41.6 ,
    \v41.7 , \v41.8 , \v41.9 , \v41.10 , \v41.11 , \v41.12 , \v41.13 ,
    \v41.14 , \v41.15 , \v41.16 , \v41.17 , \v41.18 , \v41.19 , \v41.20 ,
    \v41.21 , \v41.22 , \v41.23 , \v41.24 , \v41.25 , \v41.26 , \v41.27 ,
    \v41.28 , \v41.29 , \v41.30 , \v41.31 , \v41.32 , \v41.33 , \v41.34 ,
    \v41.35 , \v41.36 , \v41.37 , \v41.38 , \v41.39 , \v41.40 , \v41.41 ,
    \v41.42 , \v41.43 , \v41.44 , \v41.45 , \v41.46 , \v41.47 , \v41.48 ,
    \v41.49 , \v41.50 , \v41.51 , \v41.52 , \v41.53 , \v41.54 , \v41.55 ,
    \v41.56 , \v41.57 , \v41.58 , \v41.59 , \v41.60 , \v41.61 , \v41.62 ,
    \v41.63 , \v41.64 , \v41.65 , \v41.66 , \v41.67 , \v41.68 , \v41.69 ,
    \v41.70 , \v41.71 , \v41.72 ;
  wire new_n116_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_,
    new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_,
    new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_,
    new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_,
    new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_,
    new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_,
    new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_,
    new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_,
    new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_,
    new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_,
    new_n1845_, new_n1846_, new_n1848_, new_n1849_, new_n1850_, new_n1851_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_,
    new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_,
    new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_,
    new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_,
    new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_,
    new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_,
    new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_,
    new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_,
    new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_,
    new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_,
    new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_,
    new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_,
    new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_,
    new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_,
    new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_,
    new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_,
    new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_,
    new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_,
    new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_,
    new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_,
    new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_,
    new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_,
    new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_,
    new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_,
    new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_,
    new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_,
    new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_,
    new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_,
    new_n2630_, new_n2631_, new_n2632_, new_n2634_, new_n2635_, new_n2636_,
    new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_,
    new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_,
    new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_,
    new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_,
    new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_,
    new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_,
    new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_,
    new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_,
    new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_,
    new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_,
    new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_,
    new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_,
    new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_,
    new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_,
    new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_,
    new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_,
    new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_,
    new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_,
    new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_,
    new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_,
    new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_,
    new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_,
    new_n2769_, new_n2770_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_,
    new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_,
    new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_,
    new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_,
    new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_,
    new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_,
    new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_,
    new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_,
    new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_,
    new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_,
    new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_,
    new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_,
    new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_,
    new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_,
    new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_,
    new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_,
    new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_,
    new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_,
    new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_,
    new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_,
    new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_,
    new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_,
    new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_,
    new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_,
    new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_,
    new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_,
    new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_,
    new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_,
    new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_,
    new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_,
    new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_,
    new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_,
    new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_,
    new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_,
    new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_,
    new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_,
    new_n3191_, new_n3192_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3215_, new_n3216_,
    new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_,
    new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_,
    new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_,
    new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_,
    new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_,
    new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_,
    new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_,
    new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_,
    new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_,
    new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_,
    new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_,
    new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_,
    new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_,
    new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_,
    new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_,
    new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_,
    new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_,
    new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_,
    new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_,
    new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3355_, new_n3356_,
    new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3399_, new_n3400_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3424_, new_n3425_, new_n3426_,
    new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_,
    new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_,
    new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_,
    new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_,
    new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_,
    new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_,
    new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_,
    new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_,
    new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_,
    new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_,
    new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_,
    new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_,
    new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_,
    new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3530_,
    new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_,
    new_n3549_, new_n3550_, new_n3551_, new_n3553_, new_n3554_, new_n3555_,
    new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_,
    new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_,
    new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_,
    new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_,
    new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_,
    new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_,
    new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_,
    new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_,
    new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_,
    new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_,
    new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_,
    new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_,
    new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_,
    new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_,
    new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_,
    new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_,
    new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_,
    new_n3719_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3809_, new_n3810_,
    new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_,
    new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_,
    new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_,
    new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_,
    new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_,
    new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_,
    new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_,
    new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_,
    new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_,
    new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_,
    new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_,
    new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_,
    new_n3883_, new_n3884_, new_n3886_, new_n3887_, new_n3888_, new_n3889_,
    new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_,
    new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_,
    new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_,
    new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_,
    new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_,
    new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_,
    new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_,
    new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_,
    new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_,
    new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_,
    new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_,
    new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3968_,
    new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_,
    new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_,
    new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_,
    new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_,
    new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_,
    new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_,
    new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_,
    new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_,
    new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_,
    new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_,
    new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_,
    new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_,
    new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_,
    new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_,
    new_n4053_, new_n4054_, new_n4056_, new_n4057_, new_n4058_, new_n4059_,
    new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_,
    new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_,
    new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_,
    new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_,
    new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_,
    new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_,
    new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_,
    new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_,
    new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_,
    new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_,
    new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_,
    new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_,
    new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_,
    new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_,
    new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_,
    new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_,
    new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_,
    new_n4259_, new_n4260_, new_n4261_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4307_, new_n4308_,
    new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_,
    new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_,
    new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_,
    new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_,
    new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_,
    new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_,
    new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_,
    new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_,
    new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_,
    new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_,
    new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_,
    new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_,
    new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_,
    new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_,
    new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4502_,
    new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_,
    new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_,
    new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_,
    new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_,
    new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_,
    new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4580_, new_n4581_,
    new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_,
    new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_,
    new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_,
    new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_,
    new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_,
    new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_,
    new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_,
    new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_,
    new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_,
    new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_,
    new_n4679_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_,
    new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_,
    new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_,
    new_n4698_, new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_,
    new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_,
    new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_,
    new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_,
    new_n4754_, new_n4755_, new_n4757_, new_n4758_, new_n4759_, new_n4760_,
    new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_,
    new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_,
    new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4778_, new_n4779_,
    new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_,
    new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_,
    new_n4792_, new_n4793_, new_n4795_, new_n4796_, new_n4797_, new_n4798_,
    new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_,
    new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_,
    new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_,
    new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_,
    new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_,
    new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_,
    new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_,
    new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_,
    new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_,
    new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_,
    new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_,
    new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_,
    new_n4885_, new_n4886_, new_n4887_, new_n4889_, new_n4890_, new_n4891_,
    new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_,
    new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_,
    new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_,
    new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_,
    new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_,
    new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4935_,
    new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_,
    new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_,
    new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_,
    new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_,
    new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_,
    new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_,
    new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_,
    new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_,
    new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_,
    new_n5039_, new_n5040_, new_n5041_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5093_, new_n5094_,
    new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_,
    new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_,
    new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_,
    new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_,
    new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_,
    new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_,
    new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_,
    new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5162_,
    new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_,
    new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_,
    new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_,
    new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_,
    new_n5187_, new_n5188_, new_n5189_, new_n5191_, new_n5192_, new_n5193_,
    new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_,
    new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_,
    new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_,
    new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_,
    new_n5218_, new_n5219_;
  assign new_n116_ = ~v15 & v16;
  assign new_n117_ = v15 & ~v16;
  assign new_n118_ = ~new_n116_ & ~new_n117_;
  assign new_n119_ = ~v17 & ~v18;
  assign new_n120_ = v18 & v19;
  assign new_n121_ = v17 & new_n120_;
  assign new_n122_ = ~new_n119_ & ~new_n121_;
  assign new_n123_ = ~new_n118_ & ~new_n122_;
  assign new_n124_ = v16 & new_n119_;
  assign new_n125_ = v15 & new_n124_;
  assign new_n126_ = ~new_n123_ & ~new_n125_;
  assign new_n127_ = ~v12 & ~new_n126_;
  assign new_n128_ = v25 & v28;
  assign new_n129_ = v24 & new_n128_;
  assign new_n130_ = ~v28 & ~v31;
  assign new_n131_ = ~new_n129_ & ~new_n130_;
  assign new_n132_ = ~v15 & ~new_n131_;
  assign new_n133_ = ~v15 & ~new_n132_;
  assign new_n134_ = v12 & ~new_n133_;
  assign new_n135_ = ~new_n127_ & ~new_n134_;
  assign new_n136_ = v40 & ~new_n135_;
  assign new_n137_ = ~v5 & new_n136_;
  assign new_n138_ = v15 & new_n119_;
  assign new_n139_ = new_n116_ & new_n121_;
  assign new_n140_ = ~new_n138_ & ~new_n139_;
  assign new_n141_ = ~v12 & ~new_n140_;
  assign new_n142_ = v5 & new_n141_;
  assign new_n143_ = ~new_n137_ & ~new_n142_;
  assign new_n144_ = ~v4 & ~new_n143_;
  assign new_n145_ = v4 & new_n141_;
  assign new_n146_ = ~new_n144_ & ~new_n145_;
  assign new_n147_ = ~v3 & ~new_n146_;
  assign new_n148_ = v3 & new_n141_;
  assign new_n149_ = ~new_n147_ & ~new_n148_;
  assign new_n150_ = ~v2 & ~new_n149_;
  assign new_n151_ = v2 & new_n141_;
  assign new_n152_ = ~new_n150_ & ~new_n151_;
  assign new_n153_ = ~v1 & ~new_n152_;
  assign new_n154_ = ~v16 & v19;
  assign new_n155_ = v16 & ~v19;
  assign new_n156_ = ~new_n154_ & ~new_n155_;
  assign new_n157_ = ~v18 & ~new_n156_;
  assign new_n158_ = ~v17 & new_n157_;
  assign new_n159_ = v15 & new_n158_;
  assign new_n160_ = ~new_n139_ & ~new_n159_;
  assign new_n161_ = ~v2 & ~v3;
  assign new_n162_ = ~v4 & v15;
  assign new_n163_ = new_n161_ & new_n162_;
  assign new_n164_ = v16 & ~v17;
  assign new_n165_ = ~v18 & v19;
  assign new_n166_ = new_n164_ & new_n165_;
  assign new_n167_ = new_n163_ & new_n166_;
  assign new_n168_ = new_n160_ & ~new_n167_;
  assign new_n169_ = ~v4 & ~v5;
  assign new_n170_ = new_n161_ & new_n169_;
  assign new_n171_ = ~v18 & ~v19;
  assign new_n172_ = ~v17 & new_n171_;
  assign new_n173_ = new_n117_ & new_n172_;
  assign new_n174_ = new_n170_ & new_n173_;
  assign new_n175_ = new_n168_ & ~new_n174_;
  assign new_n176_ = ~v12 & ~new_n175_;
  assign new_n177_ = v1 & new_n176_;
  assign new_n178_ = ~new_n153_ & ~new_n177_;
  assign new_n179_ = v13 & ~new_n178_;
  assign new_n180_ = v15 & v19;
  assign new_n181_ = ~v15 & ~v19;
  assign new_n182_ = ~new_n180_ & ~new_n181_;
  assign new_n183_ = v17 & ~v19;
  assign new_n184_ = v15 & new_n183_;
  assign new_n185_ = new_n182_ & ~new_n184_;
  assign new_n186_ = ~v18 & ~new_n185_;
  assign new_n187_ = ~v15 & v19;
  assign new_n188_ = v15 & ~v19;
  assign new_n189_ = ~new_n187_ & ~new_n188_;
  assign new_n190_ = v18 & ~new_n189_;
  assign new_n191_ = v17 & new_n190_;
  assign new_n192_ = ~new_n186_ & ~new_n191_;
  assign new_n193_ = ~v16 & ~new_n192_;
  assign new_n194_ = ~v18 & ~new_n165_;
  assign new_n195_ = v17 & ~new_n194_;
  assign new_n196_ = v16 & new_n195_;
  assign new_n197_ = ~v15 & new_n196_;
  assign new_n198_ = ~new_n193_ & ~new_n197_;
  assign new_n199_ = v40 & ~new_n198_;
  assign new_n200_ = ~v5 & new_n199_;
  assign new_n201_ = ~v15 & ~v16;
  assign new_n202_ = v5 & new_n201_;
  assign new_n203_ = v17 & new_n171_;
  assign new_n204_ = new_n202_ & new_n203_;
  assign new_n205_ = ~new_n200_ & ~new_n204_;
  assign new_n206_ = ~v3 & ~new_n205_;
  assign new_n207_ = ~v5 & ~v15;
  assign new_n208_ = v3 & new_n207_;
  assign new_n209_ = ~v16 & v17;
  assign new_n210_ = new_n171_ & new_n209_;
  assign new_n211_ = new_n208_ & new_n210_;
  assign new_n212_ = ~new_n206_ & ~new_n211_;
  assign new_n213_ = ~v13 & ~new_n212_;
  assign new_n214_ = v12 & new_n213_;
  assign new_n215_ = ~v4 & new_n214_;
  assign new_n216_ = ~v2 & new_n215_;
  assign new_n217_ = ~v1 & new_n216_;
  assign new_n218_ = ~new_n179_ & ~new_n217_;
  assign new_n219_ = ~v14 & ~new_n218_;
  assign new_n220_ = v13 & v16;
  assign new_n221_ = new_n172_ & new_n220_;
  assign new_n222_ = v13 & ~new_n221_;
  assign new_n223_ = ~v15 & new_n171_;
  assign new_n224_ = ~new_n180_ & ~new_n223_;
  assign new_n225_ = ~v17 & ~new_n224_;
  assign new_n226_ = ~v15 & v17;
  assign new_n227_ = new_n120_ & new_n226_;
  assign new_n228_ = ~new_n225_ & ~new_n227_;
  assign new_n229_ = ~v16 & ~new_n228_;
  assign new_n230_ = ~v17 & ~new_n194_;
  assign new_n231_ = v16 & new_n230_;
  assign new_n232_ = v15 & new_n231_;
  assign new_n233_ = ~new_n229_ & ~new_n232_;
  assign new_n234_ = v13 & ~new_n233_;
  assign new_n235_ = new_n222_ & ~new_n234_;
  assign new_n236_ = v40 & ~new_n235_;
  assign new_n237_ = v14 & new_n236_;
  assign new_n238_ = v12 & new_n237_;
  assign new_n239_ = ~v5 & new_n238_;
  assign new_n240_ = ~v4 & new_n239_;
  assign new_n241_ = ~v3 & new_n240_;
  assign new_n242_ = ~v2 & new_n241_;
  assign new_n243_ = ~v1 & new_n242_;
  assign new_n244_ = ~new_n219_ & ~new_n243_;
  assign new_n245_ = ~v0 & ~new_n244_;
  assign new_n246_ = v15 & ~v17;
  assign new_n247_ = new_n171_ & new_n246_;
  assign new_n248_ = ~new_n227_ & ~new_n247_;
  assign new_n249_ = v4 & ~v5;
  assign new_n250_ = v4 & ~new_n249_;
  assign new_n251_ = ~v3 & ~new_n250_;
  assign new_n252_ = v3 & new_n169_;
  assign new_n253_ = ~new_n251_ & ~new_n252_;
  assign new_n254_ = ~new_n248_ & ~new_n253_;
  assign new_n255_ = v16 & new_n254_;
  assign new_n256_ = ~v3 & ~v4;
  assign new_n257_ = ~v5 & v15;
  assign new_n258_ = new_n256_ & new_n257_;
  assign new_n259_ = ~v16 & ~v17;
  assign new_n260_ = new_n165_ & new_n259_;
  assign new_n261_ = new_n258_ & new_n260_;
  assign new_n262_ = ~new_n255_ & ~new_n261_;
  assign new_n263_ = v13 & ~new_n262_;
  assign new_n264_ = ~v12 & new_n263_;
  assign new_n265_ = v12 & ~v13;
  assign new_n266_ = ~v5 & new_n265_;
  assign new_n267_ = new_n256_ & new_n266_;
  assign new_n268_ = new_n201_ & new_n203_;
  assign new_n269_ = new_n267_ & new_n268_;
  assign new_n270_ = ~new_n264_ & ~new_n269_;
  assign new_n271_ = ~v14 & ~new_n270_;
  assign new_n272_ = ~v2 & new_n271_;
  assign new_n273_ = ~v1 & new_n272_;
  assign new_n274_ = v0 & new_n273_;
  assign new_n275_ = ~new_n245_ & ~new_n274_;
  assign new_n276_ = ~v36 & ~new_n275_;
  assign new_n277_ = ~v11 & new_n276_;
  assign new_n278_ = ~v10 & new_n277_;
  assign new_n279_ = ~v9 & new_n278_;
  assign \v41.0  = ~v8 & new_n279_;
  assign new_n281_ = new_n165_ & new_n226_;
  assign new_n282_ = ~new_n246_ & ~new_n281_;
  assign new_n283_ = ~v16 & ~new_n282_;
  assign new_n284_ = v13 & new_n283_;
  assign new_n285_ = v13 & ~new_n284_;
  assign new_n286_ = v14 & ~new_n285_;
  assign new_n287_ = ~v15 & ~v28;
  assign new_n288_ = ~v14 & new_n287_;
  assign new_n289_ = v13 & new_n288_;
  assign new_n290_ = ~new_n286_ & ~new_n289_;
  assign new_n291_ = v40 & ~new_n290_;
  assign new_n292_ = ~v36 & new_n291_;
  assign new_n293_ = v12 & new_n292_;
  assign new_n294_ = ~v11 & new_n293_;
  assign new_n295_ = ~v10 & new_n294_;
  assign new_n296_ = ~v9 & new_n295_;
  assign new_n297_ = ~v8 & new_n296_;
  assign new_n298_ = ~v5 & new_n297_;
  assign new_n299_ = ~v4 & new_n298_;
  assign new_n300_ = ~v3 & new_n299_;
  assign new_n301_ = ~v2 & new_n300_;
  assign new_n302_ = ~v1 & new_n301_;
  assign \v41.2  = ~v0 & new_n302_;
  assign new_n304_ = v15 & new_n259_;
  assign new_n305_ = v13 & new_n304_;
  assign new_n306_ = v13 & ~new_n305_;
  assign new_n307_ = v14 & ~new_n306_;
  assign new_n308_ = v24 & ~v25;
  assign new_n309_ = v24 & ~new_n308_;
  assign new_n310_ = v28 & ~new_n309_;
  assign new_n311_ = v28 & ~new_n310_;
  assign new_n312_ = ~v15 & ~new_n311_;
  assign new_n313_ = ~v14 & new_n312_;
  assign new_n314_ = v13 & new_n313_;
  assign new_n315_ = ~new_n307_ & ~new_n314_;
  assign new_n316_ = v40 & ~new_n315_;
  assign new_n317_ = ~v36 & new_n316_;
  assign new_n318_ = v12 & new_n317_;
  assign new_n319_ = ~v11 & new_n318_;
  assign new_n320_ = ~v10 & new_n319_;
  assign new_n321_ = ~v9 & new_n320_;
  assign new_n322_ = ~v8 & new_n321_;
  assign new_n323_ = ~v5 & new_n322_;
  assign new_n324_ = ~v4 & new_n323_;
  assign new_n325_ = ~v3 & new_n324_;
  assign new_n326_ = ~v2 & new_n325_;
  assign new_n327_ = ~v1 & new_n326_;
  assign \v41.3  = ~v0 & new_n327_;
  assign new_n329_ = ~v2 & v3;
  assign new_n330_ = ~v2 & ~new_n329_;
  assign new_n331_ = ~v14 & ~new_n330_;
  assign new_n332_ = ~v12 & new_n331_;
  assign new_n333_ = v14 & v40;
  assign new_n334_ = v12 & new_n333_;
  assign new_n335_ = new_n161_ & new_n334_;
  assign new_n336_ = ~new_n332_ & ~new_n335_;
  assign new_n337_ = ~v18 & ~new_n336_;
  assign new_n338_ = ~v3 & v12;
  assign new_n339_ = ~v2 & new_n338_;
  assign new_n340_ = v18 & v40;
  assign new_n341_ = v14 & new_n340_;
  assign new_n342_ = new_n339_ & new_n341_;
  assign new_n343_ = ~new_n337_ & ~new_n342_;
  assign new_n344_ = ~v5 & ~new_n343_;
  assign new_n345_ = ~v18 & ~new_n330_;
  assign new_n346_ = ~v14 & new_n345_;
  assign new_n347_ = ~v12 & new_n346_;
  assign new_n348_ = v5 & new_n347_;
  assign new_n349_ = ~new_n344_ & ~new_n348_;
  assign new_n350_ = ~v4 & ~new_n349_;
  assign new_n351_ = ~v3 & v5;
  assign new_n352_ = ~v2 & new_n351_;
  assign new_n353_ = new_n330_ & ~new_n352_;
  assign new_n354_ = ~v18 & ~new_n353_;
  assign new_n355_ = ~v14 & new_n354_;
  assign new_n356_ = ~v12 & new_n355_;
  assign new_n357_ = v4 & new_n356_;
  assign new_n358_ = ~new_n350_ & ~new_n357_;
  assign new_n359_ = ~v16 & ~new_n358_;
  assign new_n360_ = v4 & v5;
  assign new_n361_ = new_n161_ & new_n360_;
  assign new_n362_ = new_n330_ & ~new_n361_;
  assign new_n363_ = ~v18 & ~new_n362_;
  assign new_n364_ = v16 & new_n363_;
  assign new_n365_ = ~v14 & new_n364_;
  assign new_n366_ = ~v12 & new_n365_;
  assign new_n367_ = ~new_n359_ & ~new_n366_;
  assign new_n368_ = ~v1 & ~new_n367_;
  assign new_n369_ = v5 & v16;
  assign new_n370_ = v5 & ~new_n369_;
  assign new_n371_ = ~v18 & ~new_n370_;
  assign new_n372_ = ~v14 & new_n371_;
  assign new_n373_ = ~v12 & new_n372_;
  assign new_n374_ = ~v4 & new_n373_;
  assign new_n375_ = ~v3 & new_n374_;
  assign new_n376_ = ~v2 & new_n375_;
  assign new_n377_ = v1 & new_n376_;
  assign new_n378_ = ~new_n368_ & ~new_n377_;
  assign new_n379_ = v15 & ~new_n378_;
  assign new_n380_ = ~v1 & ~v2;
  assign new_n381_ = ~v3 & new_n169_;
  assign new_n382_ = new_n380_ & new_n381_;
  assign new_n383_ = ~v14 & ~v15;
  assign new_n384_ = ~v12 & new_n383_;
  assign new_n385_ = ~v18 & v40;
  assign new_n386_ = v16 & new_n385_;
  assign new_n387_ = new_n384_ & new_n386_;
  assign new_n388_ = new_n382_ & new_n387_;
  assign new_n389_ = ~new_n379_ & ~new_n388_;
  assign new_n390_ = ~v3 & v4;
  assign new_n391_ = ~v2 & new_n390_;
  assign new_n392_ = new_n330_ & ~new_n391_;
  assign new_n393_ = v1 & ~new_n392_;
  assign new_n394_ = ~v1 & new_n161_;
  assign new_n395_ = ~v5 & v40;
  assign new_n396_ = ~v4 & new_n395_;
  assign new_n397_ = new_n394_ & new_n396_;
  assign new_n398_ = ~new_n393_ & ~new_n397_;
  assign new_n399_ = ~new_n156_ & ~new_n398_;
  assign new_n400_ = v16 & v19;
  assign new_n401_ = ~v16 & ~v19;
  assign new_n402_ = ~new_n400_ & ~new_n401_;
  assign new_n403_ = ~v4 & v5;
  assign new_n404_ = ~new_n249_ & ~new_n403_;
  assign new_n405_ = ~new_n402_ & ~new_n404_;
  assign new_n406_ = ~v1 & new_n405_;
  assign new_n407_ = v1 & ~v4;
  assign new_n408_ = v5 & new_n154_;
  assign new_n409_ = new_n407_ & new_n408_;
  assign new_n410_ = ~new_n406_ & ~new_n409_;
  assign new_n411_ = ~v3 & ~new_n410_;
  assign new_n412_ = ~v2 & new_n411_;
  assign new_n413_ = ~new_n399_ & ~new_n412_;
  assign new_n414_ = ~v18 & ~new_n413_;
  assign new_n415_ = v15 & new_n414_;
  assign new_n416_ = ~v14 & new_n415_;
  assign new_n417_ = ~v12 & new_n416_;
  assign new_n418_ = new_n389_ & ~new_n417_;
  assign new_n419_ = ~v17 & ~new_n418_;
  assign new_n420_ = ~v3 & v40;
  assign new_n421_ = ~v3 & ~new_n420_;
  assign new_n422_ = ~v2 & ~new_n421_;
  assign new_n423_ = ~v2 & ~new_n422_;
  assign new_n424_ = v16 & ~new_n423_;
  assign new_n425_ = ~v15 & new_n424_;
  assign new_n426_ = ~v16 & v40;
  assign new_n427_ = v15 & new_n426_;
  assign new_n428_ = new_n161_ & new_n427_;
  assign new_n429_ = ~new_n425_ & ~new_n428_;
  assign new_n430_ = v19 & ~new_n429_;
  assign new_n431_ = v18 & new_n430_;
  assign new_n432_ = v17 & new_n431_;
  assign new_n433_ = ~v12 & new_n432_;
  assign new_n434_ = ~v15 & v24;
  assign new_n435_ = v27 & v28;
  assign new_n436_ = v25 & new_n435_;
  assign new_n437_ = new_n434_ & new_n436_;
  assign new_n438_ = v15 & v29;
  assign new_n439_ = ~new_n437_ & ~new_n438_;
  assign new_n440_ = v40 & ~new_n439_;
  assign new_n441_ = v12 & new_n440_;
  assign new_n442_ = ~v3 & new_n441_;
  assign new_n443_ = ~v2 & new_n442_;
  assign new_n444_ = ~new_n433_ & ~new_n443_;
  assign new_n445_ = ~v1 & ~new_n444_;
  assign new_n446_ = v16 & new_n121_;
  assign new_n447_ = ~v15 & new_n446_;
  assign new_n448_ = ~v12 & new_n447_;
  assign new_n449_ = v1 & new_n448_;
  assign new_n450_ = ~new_n445_ & ~new_n449_;
  assign new_n451_ = ~v5 & ~new_n450_;
  assign new_n452_ = ~v1 & v2;
  assign new_n453_ = ~v1 & ~new_n452_;
  assign new_n454_ = ~v1 & new_n329_;
  assign new_n455_ = new_n453_ & ~new_n454_;
  assign new_n456_ = v19 & ~new_n455_;
  assign new_n457_ = v18 & new_n456_;
  assign new_n458_ = v17 & new_n457_;
  assign new_n459_ = v16 & new_n458_;
  assign new_n460_ = ~v15 & new_n459_;
  assign new_n461_ = ~v12 & new_n460_;
  assign new_n462_ = v5 & new_n461_;
  assign new_n463_ = ~new_n451_ & ~new_n462_;
  assign new_n464_ = ~v4 & ~new_n463_;
  assign new_n465_ = new_n351_ & new_n380_;
  assign new_n466_ = new_n455_ & ~new_n465_;
  assign new_n467_ = v19 & ~new_n466_;
  assign new_n468_ = v18 & new_n467_;
  assign new_n469_ = v17 & new_n468_;
  assign new_n470_ = v16 & new_n469_;
  assign new_n471_ = ~v15 & new_n470_;
  assign new_n472_ = ~v12 & new_n471_;
  assign new_n473_ = v4 & new_n472_;
  assign new_n474_ = ~new_n464_ & ~new_n473_;
  assign new_n475_ = ~v14 & ~new_n474_;
  assign new_n476_ = ~new_n419_ & ~new_n475_;
  assign new_n477_ = ~v0 & ~new_n476_;
  assign new_n478_ = ~v14 & ~new_n262_;
  assign new_n479_ = ~v12 & new_n478_;
  assign new_n480_ = ~v2 & new_n479_;
  assign new_n481_ = ~v1 & new_n480_;
  assign new_n482_ = v0 & new_n481_;
  assign new_n483_ = ~new_n477_ & ~new_n482_;
  assign new_n484_ = v13 & ~new_n483_;
  assign new_n485_ = v16 & v18;
  assign new_n486_ = ~v16 & ~v18;
  assign new_n487_ = ~new_n485_ & ~new_n486_;
  assign new_n488_ = ~v15 & ~new_n487_;
  assign new_n489_ = ~v16 & v18;
  assign new_n490_ = v15 & new_n489_;
  assign new_n491_ = ~new_n488_ & ~new_n490_;
  assign new_n492_ = v40 & ~new_n491_;
  assign new_n493_ = ~v3 & new_n492_;
  assign new_n494_ = v3 & ~v15;
  assign new_n495_ = new_n486_ & new_n494_;
  assign new_n496_ = ~new_n493_ & ~new_n495_;
  assign new_n497_ = ~v0 & ~new_n496_;
  assign new_n498_ = v0 & ~v3;
  assign new_n499_ = ~v15 & new_n486_;
  assign new_n500_ = new_n498_ & new_n499_;
  assign new_n501_ = ~new_n497_ & ~new_n500_;
  assign new_n502_ = ~v19 & ~new_n501_;
  assign new_n503_ = v17 & new_n502_;
  assign new_n504_ = ~v14 & new_n503_;
  assign new_n505_ = ~v13 & new_n504_;
  assign new_n506_ = v12 & new_n505_;
  assign new_n507_ = ~v5 & new_n506_;
  assign new_n508_ = ~v4 & new_n507_;
  assign new_n509_ = ~v2 & new_n508_;
  assign new_n510_ = ~v1 & new_n509_;
  assign new_n511_ = ~new_n484_ & ~new_n510_;
  assign new_n512_ = ~v36 & ~new_n511_;
  assign new_n513_ = ~v11 & new_n512_;
  assign new_n514_ = ~v10 & new_n513_;
  assign new_n515_ = ~v9 & new_n514_;
  assign \v41.4  = ~v8 & new_n515_;
  assign new_n517_ = v17 & v18;
  assign new_n518_ = ~new_n119_ & ~new_n517_;
  assign new_n519_ = ~new_n118_ & ~new_n518_;
  assign new_n520_ = v19 & new_n519_;
  assign new_n521_ = v16 & new_n172_;
  assign new_n522_ = ~new_n520_ & ~new_n521_;
  assign new_n523_ = ~v12 & ~new_n522_;
  assign new_n524_ = v25 & v27;
  assign new_n525_ = v25 & ~new_n524_;
  assign new_n526_ = v24 & ~new_n525_;
  assign new_n527_ = v24 & ~new_n526_;
  assign new_n528_ = v28 & ~new_n527_;
  assign new_n529_ = v28 & ~new_n528_;
  assign new_n530_ = ~v15 & ~new_n529_;
  assign new_n531_ = ~new_n438_ & ~new_n530_;
  assign new_n532_ = v12 & ~new_n531_;
  assign new_n533_ = ~new_n523_ & ~new_n532_;
  assign new_n534_ = v40 & ~new_n533_;
  assign new_n535_ = ~v3 & new_n534_;
  assign new_n536_ = ~new_n148_ & ~new_n535_;
  assign new_n537_ = ~v2 & ~new_n536_;
  assign new_n538_ = ~new_n151_ & ~new_n537_;
  assign new_n539_ = ~v5 & ~new_n538_;
  assign new_n540_ = v2 & ~new_n156_;
  assign new_n541_ = new_n402_ & ~new_n540_;
  assign new_n542_ = ~v18 & ~new_n541_;
  assign new_n543_ = ~v17 & new_n542_;
  assign new_n544_ = v15 & new_n543_;
  assign new_n545_ = v2 & new_n116_;
  assign new_n546_ = new_n121_ & new_n545_;
  assign new_n547_ = ~new_n544_ & ~new_n546_;
  assign new_n548_ = v3 & ~new_n160_;
  assign new_n549_ = ~v2 & new_n548_;
  assign new_n550_ = new_n547_ & ~new_n549_;
  assign new_n551_ = ~v12 & ~new_n550_;
  assign new_n552_ = v5 & new_n551_;
  assign new_n553_ = ~new_n539_ & ~new_n552_;
  assign new_n554_ = ~v4 & ~new_n553_;
  assign new_n555_ = v5 & ~new_n160_;
  assign new_n556_ = ~v3 & new_n555_;
  assign new_n557_ = ~v2 & new_n556_;
  assign new_n558_ = new_n550_ & ~new_n557_;
  assign new_n559_ = ~v12 & ~new_n558_;
  assign new_n560_ = v4 & new_n559_;
  assign new_n561_ = ~new_n554_ & ~new_n560_;
  assign new_n562_ = ~v1 & ~new_n561_;
  assign new_n563_ = ~new_n177_ & ~new_n562_;
  assign new_n564_ = ~v0 & ~new_n563_;
  assign new_n565_ = ~v12 & ~new_n262_;
  assign new_n566_ = ~v2 & new_n565_;
  assign new_n567_ = ~v1 & new_n566_;
  assign new_n568_ = v0 & new_n567_;
  assign new_n569_ = ~new_n564_ & ~new_n568_;
  assign new_n570_ = v13 & ~new_n569_;
  assign new_n571_ = ~v13 & new_n503_;
  assign new_n572_ = v12 & new_n571_;
  assign new_n573_ = ~v5 & new_n572_;
  assign new_n574_ = ~v4 & new_n573_;
  assign new_n575_ = ~v2 & new_n574_;
  assign new_n576_ = ~v1 & new_n575_;
  assign new_n577_ = ~new_n570_ & ~new_n576_;
  assign new_n578_ = ~v14 & ~new_n577_;
  assign new_n579_ = ~v17 & v40;
  assign new_n580_ = ~v16 & new_n579_;
  assign new_n581_ = v15 & new_n580_;
  assign new_n582_ = v14 & new_n581_;
  assign new_n583_ = v13 & new_n582_;
  assign new_n584_ = v12 & new_n583_;
  assign new_n585_ = ~v5 & new_n584_;
  assign new_n586_ = ~v4 & new_n585_;
  assign new_n587_ = ~v3 & new_n586_;
  assign new_n588_ = ~v2 & new_n587_;
  assign new_n589_ = ~v1 & new_n588_;
  assign new_n590_ = ~v0 & new_n589_;
  assign new_n591_ = ~new_n578_ & ~new_n590_;
  assign new_n592_ = ~v36 & ~new_n591_;
  assign new_n593_ = ~v11 & new_n592_;
  assign new_n594_ = ~v10 & new_n593_;
  assign new_n595_ = ~v9 & new_n594_;
  assign \v41.5  = ~v8 & new_n595_;
  assign new_n597_ = new_n117_ & new_n517_;
  assign new_n598_ = new_n116_ & new_n119_;
  assign new_n599_ = ~new_n597_ & ~new_n598_;
  assign new_n600_ = v40 & ~new_n599_;
  assign new_n601_ = ~v5 & new_n600_;
  assign new_n602_ = new_n116_ & new_n517_;
  assign new_n603_ = ~new_n138_ & ~new_n602_;
  assign new_n604_ = v5 & ~new_n603_;
  assign new_n605_ = ~new_n601_ & ~new_n604_;
  assign new_n606_ = v19 & ~new_n605_;
  assign new_n607_ = v5 & v15;
  assign new_n608_ = v16 & v40;
  assign new_n609_ = new_n207_ & new_n608_;
  assign new_n610_ = ~new_n607_ & ~new_n609_;
  assign new_n611_ = ~v19 & ~new_n610_;
  assign new_n612_ = ~v18 & new_n611_;
  assign new_n613_ = ~v17 & new_n612_;
  assign new_n614_ = ~new_n606_ & ~new_n613_;
  assign new_n615_ = ~v12 & ~new_n614_;
  assign new_n616_ = v40 & ~new_n531_;
  assign new_n617_ = v12 & new_n616_;
  assign new_n618_ = ~v5 & new_n617_;
  assign new_n619_ = ~new_n615_ & ~new_n618_;
  assign new_n620_ = ~v4 & ~new_n619_;
  assign new_n621_ = ~new_n145_ & ~new_n620_;
  assign new_n622_ = ~v3 & ~new_n621_;
  assign new_n623_ = ~new_n148_ & ~new_n622_;
  assign new_n624_ = ~v2 & ~new_n623_;
  assign new_n625_ = ~new_n151_ & ~new_n624_;
  assign new_n626_ = ~v1 & ~new_n625_;
  assign new_n627_ = ~new_n177_ & ~new_n626_;
  assign new_n628_ = ~v0 & ~new_n627_;
  assign new_n629_ = ~new_n248_ & ~new_n250_;
  assign new_n630_ = v16 & new_n629_;
  assign new_n631_ = ~v4 & new_n257_;
  assign new_n632_ = new_n260_ & new_n631_;
  assign new_n633_ = ~new_n630_ & ~new_n632_;
  assign new_n634_ = ~v12 & ~new_n633_;
  assign new_n635_ = ~v3 & new_n634_;
  assign new_n636_ = ~v2 & new_n635_;
  assign new_n637_ = ~v1 & new_n636_;
  assign new_n638_ = v0 & new_n637_;
  assign new_n639_ = ~new_n628_ & ~new_n638_;
  assign new_n640_ = ~v14 & ~new_n639_;
  assign new_n641_ = v12 & new_n582_;
  assign new_n642_ = ~v5 & new_n641_;
  assign new_n643_ = ~v4 & new_n642_;
  assign new_n644_ = ~v3 & new_n643_;
  assign new_n645_ = ~v2 & new_n644_;
  assign new_n646_ = ~v1 & new_n645_;
  assign new_n647_ = ~v0 & new_n646_;
  assign new_n648_ = ~new_n640_ & ~new_n647_;
  assign new_n649_ = v13 & ~new_n648_;
  assign new_n650_ = v40 & ~new_n118_;
  assign new_n651_ = v18 & new_n650_;
  assign new_n652_ = ~v5 & new_n651_;
  assign new_n653_ = v5 & ~v15;
  assign new_n654_ = new_n486_ & new_n653_;
  assign new_n655_ = ~new_n652_ & ~new_n654_;
  assign new_n656_ = ~v19 & ~new_n655_;
  assign new_n657_ = v17 & new_n656_;
  assign new_n658_ = ~v14 & new_n657_;
  assign new_n659_ = ~v13 & new_n658_;
  assign new_n660_ = v12 & new_n659_;
  assign new_n661_ = ~v4 & new_n660_;
  assign new_n662_ = ~v3 & new_n661_;
  assign new_n663_ = ~v2 & new_n662_;
  assign new_n664_ = ~v1 & new_n663_;
  assign new_n665_ = ~v0 & new_n664_;
  assign new_n666_ = ~new_n649_ & ~new_n665_;
  assign new_n667_ = ~v36 & ~new_n666_;
  assign new_n668_ = ~v11 & new_n667_;
  assign new_n669_ = ~v10 & new_n668_;
  assign new_n670_ = ~v9 & new_n669_;
  assign \v41.6  = ~v8 & new_n670_;
  assign new_n672_ = ~v5 & ~new_n395_;
  assign new_n673_ = v16 & v17;
  assign new_n674_ = ~v15 & new_n673_;
  assign new_n675_ = ~new_n246_ & ~new_n674_;
  assign new_n676_ = ~v18 & ~new_n675_;
  assign new_n677_ = v13 & new_n676_;
  assign new_n678_ = ~v12 & new_n677_;
  assign new_n679_ = v20 & ~v21;
  assign new_n680_ = v22 & ~v23;
  assign new_n681_ = v22 & ~new_n680_;
  assign new_n682_ = ~v24 & ~new_n681_;
  assign new_n683_ = v21 & new_n682_;
  assign new_n684_ = ~v20 & new_n683_;
  assign new_n685_ = ~new_n679_ & ~new_n684_;
  assign new_n686_ = v24 & ~v26;
  assign new_n687_ = v24 & ~new_n686_;
  assign new_n688_ = v23 & ~new_n687_;
  assign new_n689_ = ~v23 & v24;
  assign new_n690_ = ~new_n688_ & ~new_n689_;
  assign new_n691_ = v22 & ~new_n690_;
  assign new_n692_ = ~v22 & v24;
  assign new_n693_ = ~new_n691_ & ~new_n692_;
  assign new_n694_ = v27 & ~new_n693_;
  assign new_n695_ = v21 & new_n694_;
  assign new_n696_ = ~v20 & new_n695_;
  assign new_n697_ = new_n685_ & ~new_n696_;
  assign new_n698_ = v18 & ~new_n697_;
  assign new_n699_ = v17 & new_n698_;
  assign new_n700_ = ~v16 & new_n699_;
  assign new_n701_ = ~v15 & new_n700_;
  assign new_n702_ = ~v13 & new_n701_;
  assign new_n703_ = v12 & new_n702_;
  assign new_n704_ = ~new_n678_ & ~new_n703_;
  assign new_n705_ = ~v19 & ~new_n704_;
  assign new_n706_ = v19 & ~new_n603_;
  assign new_n707_ = v13 & new_n706_;
  assign new_n708_ = ~v12 & new_n707_;
  assign new_n709_ = ~new_n705_ & ~new_n708_;
  assign new_n710_ = ~new_n672_ & ~new_n709_;
  assign new_n711_ = v32 & v33;
  assign new_n712_ = v30 & new_n711_;
  assign new_n713_ = ~v30 & ~v31;
  assign new_n714_ = ~new_n712_ & ~new_n713_;
  assign new_n715_ = v13 & ~new_n714_;
  assign new_n716_ = v26 & v27;
  assign new_n717_ = v27 & ~new_n716_;
  assign new_n718_ = v24 & ~new_n717_;
  assign new_n719_ = ~v24 & ~v27;
  assign new_n720_ = ~new_n718_ & ~new_n719_;
  assign new_n721_ = v23 & ~new_n720_;
  assign new_n722_ = v24 & ~v27;
  assign new_n723_ = ~v23 & new_n722_;
  assign new_n724_ = ~new_n721_ & ~new_n723_;
  assign new_n725_ = v22 & ~new_n724_;
  assign new_n726_ = ~v22 & new_n722_;
  assign new_n727_ = ~new_n725_ & ~new_n726_;
  assign new_n728_ = v21 & ~new_n727_;
  assign new_n729_ = ~v20 & new_n728_;
  assign new_n730_ = v17 & new_n729_;
  assign new_n731_ = ~v16 & new_n730_;
  assign new_n732_ = ~v15 & new_n731_;
  assign new_n733_ = new_n118_ & ~new_n732_;
  assign new_n734_ = ~v19 & ~new_n733_;
  assign new_n735_ = ~v17 & v19;
  assign new_n736_ = new_n117_ & new_n735_;
  assign new_n737_ = ~new_n734_ & ~new_n736_;
  assign new_n738_ = v18 & ~new_n737_;
  assign new_n739_ = v19 & ~new_n118_;
  assign new_n740_ = v38 & v39;
  assign new_n741_ = ~v19 & ~new_n740_;
  assign new_n742_ = v16 & new_n741_;
  assign new_n743_ = ~v15 & new_n742_;
  assign new_n744_ = ~new_n739_ & ~new_n743_;
  assign new_n745_ = ~v18 & ~new_n744_;
  assign new_n746_ = v17 & new_n745_;
  assign new_n747_ = ~new_n738_ & ~new_n746_;
  assign new_n748_ = ~v13 & ~new_n747_;
  assign new_n749_ = ~new_n715_ & ~new_n748_;
  assign new_n750_ = v12 & ~new_n749_;
  assign new_n751_ = v15 & new_n209_;
  assign new_n752_ = ~new_n598_ & ~new_n751_;
  assign new_n753_ = ~v17 & v18;
  assign new_n754_ = v17 & ~v18;
  assign new_n755_ = ~new_n753_ & ~new_n754_;
  assign new_n756_ = v19 & ~new_n755_;
  assign new_n757_ = v16 & new_n756_;
  assign new_n758_ = ~v15 & new_n757_;
  assign new_n759_ = new_n752_ & ~new_n758_;
  assign new_n760_ = v13 & ~new_n759_;
  assign new_n761_ = ~v12 & new_n760_;
  assign new_n762_ = ~new_n750_ & ~new_n761_;
  assign new_n763_ = v40 & ~new_n762_;
  assign new_n764_ = ~v5 & new_n763_;
  assign new_n765_ = v5 & v12;
  assign new_n766_ = ~v13 & ~v15;
  assign new_n767_ = new_n765_ & new_n766_;
  assign new_n768_ = new_n210_ & new_n767_;
  assign new_n769_ = ~new_n764_ & ~new_n768_;
  assign new_n770_ = ~new_n710_ & new_n769_;
  assign new_n771_ = ~v4 & ~new_n770_;
  assign new_n772_ = v13 & new_n138_;
  assign new_n773_ = ~v12 & new_n772_;
  assign new_n774_ = v27 & ~new_n685_;
  assign new_n775_ = ~v19 & new_n774_;
  assign new_n776_ = v18 & new_n775_;
  assign new_n777_ = v17 & new_n776_;
  assign new_n778_ = ~v15 & new_n777_;
  assign new_n779_ = ~v13 & new_n778_;
  assign new_n780_ = v12 & new_n779_;
  assign new_n781_ = ~new_n773_ & ~new_n780_;
  assign new_n782_ = ~v16 & ~new_n781_;
  assign new_n783_ = ~new_n138_ & ~new_n227_;
  assign new_n784_ = v16 & ~new_n783_;
  assign new_n785_ = v13 & new_n784_;
  assign new_n786_ = ~v12 & new_n785_;
  assign new_n787_ = ~new_n782_ & ~new_n786_;
  assign new_n788_ = v4 & ~new_n787_;
  assign new_n789_ = ~new_n771_ & ~new_n788_;
  assign new_n790_ = ~v3 & ~new_n789_;
  assign new_n791_ = v13 & ~new_n140_;
  assign new_n792_ = ~v12 & new_n791_;
  assign new_n793_ = v3 & new_n792_;
  assign new_n794_ = ~new_n790_ & ~new_n793_;
  assign new_n795_ = ~v2 & ~new_n794_;
  assign new_n796_ = v2 & new_n792_;
  assign new_n797_ = ~new_n795_ & ~new_n796_;
  assign new_n798_ = ~v1 & ~new_n797_;
  assign new_n799_ = v13 & ~new_n175_;
  assign new_n800_ = ~v12 & new_n799_;
  assign new_n801_ = v1 & new_n800_;
  assign new_n802_ = ~new_n798_ & ~new_n801_;
  assign new_n803_ = ~v0 & ~new_n802_;
  assign new_n804_ = v13 & ~new_n633_;
  assign new_n805_ = ~v12 & new_n804_;
  assign new_n806_ = new_n169_ & new_n265_;
  assign new_n807_ = new_n268_ & new_n806_;
  assign new_n808_ = ~new_n805_ & ~new_n807_;
  assign new_n809_ = ~v3 & ~new_n808_;
  assign new_n810_ = ~v2 & new_n809_;
  assign new_n811_ = ~v1 & new_n810_;
  assign new_n812_ = v0 & new_n811_;
  assign new_n813_ = ~new_n803_ & ~new_n812_;
  assign new_n814_ = ~v14 & ~new_n813_;
  assign new_n815_ = new_n116_ & new_n171_;
  assign new_n816_ = ~new_n490_ & ~new_n815_;
  assign new_n817_ = ~v17 & ~new_n816_;
  assign new_n818_ = v12 & new_n817_;
  assign new_n819_ = v12 & ~new_n818_;
  assign new_n820_ = v13 & ~new_n819_;
  assign new_n821_ = ~v13 & v15;
  assign new_n822_ = v12 & new_n821_;
  assign new_n823_ = ~new_n820_ & ~new_n822_;
  assign new_n824_ = v40 & ~new_n823_;
  assign new_n825_ = v14 & new_n824_;
  assign new_n826_ = ~v5 & new_n825_;
  assign new_n827_ = ~v4 & new_n826_;
  assign new_n828_ = ~v3 & new_n827_;
  assign new_n829_ = ~v2 & new_n828_;
  assign new_n830_ = ~v1 & new_n829_;
  assign new_n831_ = ~v0 & new_n830_;
  assign new_n832_ = ~new_n814_ & ~new_n831_;
  assign new_n833_ = ~v36 & ~new_n832_;
  assign new_n834_ = ~v11 & new_n833_;
  assign new_n835_ = ~v10 & new_n834_;
  assign new_n836_ = ~v9 & new_n835_;
  assign \v41.7  = ~v8 & new_n836_;
  assign new_n838_ = v10 & v11;
  assign new_n839_ = v10 & ~new_n838_;
  assign new_n840_ = v9 & ~new_n839_;
  assign new_n841_ = ~v15 & new_n485_;
  assign new_n842_ = v15 & new_n486_;
  assign new_n843_ = ~v38 & ~v39;
  assign new_n844_ = ~v37 & new_n843_;
  assign new_n845_ = new_n842_ & new_n844_;
  assign new_n846_ = ~new_n841_ & ~new_n845_;
  assign new_n847_ = ~v13 & ~new_n846_;
  assign new_n848_ = v12 & new_n847_;
  assign new_n849_ = ~v12 & v13;
  assign new_n850_ = new_n117_ & new_n849_;
  assign new_n851_ = v18 & ~v37;
  assign new_n852_ = new_n843_ & new_n851_;
  assign new_n853_ = new_n850_ & new_n852_;
  assign new_n854_ = ~new_n848_ & ~new_n853_;
  assign new_n855_ = ~v19 & ~new_n854_;
  assign new_n856_ = new_n120_ & new_n844_;
  assign new_n857_ = new_n850_ & new_n856_;
  assign new_n858_ = ~new_n855_ & ~new_n857_;
  assign new_n859_ = ~v17 & ~new_n858_;
  assign new_n860_ = ~v18 & new_n741_;
  assign new_n861_ = v17 & new_n860_;
  assign new_n862_ = v16 & new_n861_;
  assign new_n863_ = ~v15 & new_n862_;
  assign new_n864_ = ~v13 & new_n863_;
  assign new_n865_ = v12 & new_n864_;
  assign new_n866_ = ~new_n859_ & ~new_n865_;
  assign new_n867_ = v40 & ~new_n866_;
  assign new_n868_ = ~v36 & new_n867_;
  assign new_n869_ = ~v14 & new_n868_;
  assign new_n870_ = ~v11 & new_n869_;
  assign new_n871_ = ~v10 & new_n870_;
  assign new_n872_ = ~v9 & new_n871_;
  assign new_n873_ = ~v5 & new_n872_;
  assign new_n874_ = ~v4 & new_n873_;
  assign new_n875_ = ~v3 & new_n874_;
  assign new_n876_ = ~v2 & new_n875_;
  assign new_n877_ = ~v1 & new_n876_;
  assign new_n878_ = ~v0 & new_n877_;
  assign new_n879_ = ~new_n840_ & ~new_n878_;
  assign \v41.8  = ~v8 & ~new_n879_;
  assign new_n881_ = ~v15 & ~v30;
  assign new_n882_ = ~v14 & new_n881_;
  assign new_n883_ = ~v16 & new_n753_;
  assign new_n884_ = v14 & new_n883_;
  assign new_n885_ = ~v14 & ~v30;
  assign new_n886_ = ~new_n884_ & ~new_n885_;
  assign new_n887_ = v15 & ~new_n886_;
  assign new_n888_ = ~new_n882_ & ~new_n887_;
  assign new_n889_ = v13 & ~new_n888_;
  assign new_n890_ = ~v18 & ~new_n740_;
  assign new_n891_ = v17 & new_n890_;
  assign new_n892_ = ~new_n753_ & ~new_n891_;
  assign new_n893_ = ~v19 & ~new_n892_;
  assign new_n894_ = v16 & new_n893_;
  assign new_n895_ = ~v15 & new_n894_;
  assign new_n896_ = ~v14 & new_n895_;
  assign new_n897_ = ~v13 & new_n896_;
  assign new_n898_ = ~new_n889_ & ~new_n897_;
  assign new_n899_ = v12 & ~new_n898_;
  assign new_n900_ = v14 & ~v15;
  assign new_n901_ = new_n849_ & new_n900_;
  assign new_n902_ = ~new_n899_ & ~new_n901_;
  assign new_n903_ = v40 & ~new_n902_;
  assign new_n904_ = ~v36 & new_n903_;
  assign new_n905_ = ~v11 & new_n904_;
  assign new_n906_ = ~v10 & new_n905_;
  assign new_n907_ = ~v9 & new_n906_;
  assign new_n908_ = ~v8 & new_n907_;
  assign new_n909_ = ~v5 & new_n908_;
  assign new_n910_ = ~v4 & new_n909_;
  assign new_n911_ = ~v3 & new_n910_;
  assign new_n912_ = ~v2 & new_n911_;
  assign new_n913_ = ~v1 & new_n912_;
  assign \v41.9  = ~v0 & new_n913_;
  assign new_n915_ = ~v14 & ~v16;
  assign new_n916_ = ~v14 & ~new_n915_;
  assign new_n917_ = ~v12 & ~new_n916_;
  assign new_n918_ = v32 & ~v33;
  assign new_n919_ = v32 & ~new_n918_;
  assign new_n920_ = v30 & ~new_n919_;
  assign new_n921_ = v30 & ~new_n920_;
  assign new_n922_ = ~v14 & ~new_n921_;
  assign new_n923_ = v12 & new_n922_;
  assign new_n924_ = ~new_n917_ & ~new_n923_;
  assign new_n925_ = ~v15 & ~new_n924_;
  assign new_n926_ = ~new_n884_ & ~new_n922_;
  assign new_n927_ = v15 & ~new_n926_;
  assign new_n928_ = v12 & new_n927_;
  assign new_n929_ = ~new_n925_ & ~new_n928_;
  assign new_n930_ = v13 & ~new_n929_;
  assign new_n931_ = v12 & new_n897_;
  assign new_n932_ = ~new_n930_ & ~new_n931_;
  assign new_n933_ = v40 & ~new_n932_;
  assign new_n934_ = ~v36 & new_n933_;
  assign new_n935_ = ~v11 & new_n934_;
  assign new_n936_ = ~v10 & new_n935_;
  assign new_n937_ = ~v9 & new_n936_;
  assign new_n938_ = ~v8 & new_n937_;
  assign new_n939_ = ~v5 & new_n938_;
  assign new_n940_ = ~v4 & new_n939_;
  assign new_n941_ = ~v3 & new_n940_;
  assign new_n942_ = ~v2 & new_n941_;
  assign new_n943_ = ~v1 & new_n942_;
  assign \v41.10  = ~v0 & new_n943_;
  assign new_n945_ = v18 & ~new_n852_;
  assign new_n946_ = ~v14 & ~new_n945_;
  assign new_n947_ = ~v12 & new_n946_;
  assign new_n948_ = v14 & v18;
  assign new_n949_ = v12 & new_n948_;
  assign new_n950_ = ~new_n947_ & ~new_n949_;
  assign new_n951_ = ~v16 & ~new_n950_;
  assign new_n952_ = ~v12 & ~v14;
  assign new_n953_ = v16 & ~v18;
  assign new_n954_ = new_n952_ & new_n953_;
  assign new_n955_ = ~new_n951_ & ~new_n954_;
  assign new_n956_ = ~v17 & ~new_n955_;
  assign new_n957_ = v33 & v35;
  assign new_n958_ = v33 & ~new_n957_;
  assign new_n959_ = v32 & ~new_n958_;
  assign new_n960_ = v32 & ~new_n959_;
  assign new_n961_ = v30 & ~new_n960_;
  assign new_n962_ = v30 & ~new_n961_;
  assign new_n963_ = ~v14 & ~new_n962_;
  assign new_n964_ = v12 & new_n963_;
  assign new_n965_ = ~new_n956_ & ~new_n964_;
  assign new_n966_ = v15 & ~new_n965_;
  assign new_n967_ = v12 & ~new_n962_;
  assign new_n968_ = ~v12 & v16;
  assign new_n969_ = new_n121_ & new_n968_;
  assign new_n970_ = ~new_n967_ & ~new_n969_;
  assign new_n971_ = ~v15 & ~new_n970_;
  assign new_n972_ = ~v14 & new_n971_;
  assign new_n973_ = ~new_n966_ & ~new_n972_;
  assign new_n974_ = v13 & ~new_n973_;
  assign new_n975_ = v17 & v19;
  assign new_n976_ = ~v17 & ~v19;
  assign new_n977_ = new_n844_ & new_n976_;
  assign new_n978_ = ~new_n975_ & ~new_n977_;
  assign new_n979_ = ~v16 & ~new_n978_;
  assign new_n980_ = v15 & new_n979_;
  assign new_n981_ = new_n116_ & new_n975_;
  assign new_n982_ = ~new_n980_ & ~new_n981_;
  assign new_n983_ = ~v18 & ~new_n982_;
  assign new_n984_ = ~v14 & new_n983_;
  assign new_n985_ = ~v13 & new_n984_;
  assign new_n986_ = v12 & new_n985_;
  assign new_n987_ = ~new_n974_ & ~new_n986_;
  assign new_n988_ = v40 & ~new_n987_;
  assign new_n989_ = ~v5 & new_n988_;
  assign new_n990_ = ~v16 & new_n698_;
  assign new_n991_ = ~v13 & new_n990_;
  assign new_n992_ = v12 & new_n991_;
  assign new_n993_ = new_n849_ & new_n953_;
  assign new_n994_ = ~new_n992_ & ~new_n993_;
  assign new_n995_ = ~v19 & ~new_n994_;
  assign new_n996_ = v17 & new_n995_;
  assign new_n997_ = ~v15 & new_n996_;
  assign new_n998_ = ~v14 & new_n997_;
  assign new_n999_ = v5 & new_n998_;
  assign new_n1000_ = ~new_n989_ & ~new_n999_;
  assign new_n1001_ = ~v4 & ~new_n1000_;
  assign new_n1002_ = ~v16 & new_n777_;
  assign new_n1003_ = ~v15 & new_n1002_;
  assign new_n1004_ = ~v14 & new_n1003_;
  assign new_n1005_ = ~v13 & new_n1004_;
  assign new_n1006_ = v12 & new_n1005_;
  assign new_n1007_ = v4 & new_n1006_;
  assign new_n1008_ = ~new_n1001_ & ~new_n1007_;
  assign new_n1009_ = ~v0 & ~new_n1008_;
  assign new_n1010_ = v0 & ~v4;
  assign new_n1011_ = new_n266_ & new_n1010_;
  assign new_n1012_ = ~v14 & new_n201_;
  assign new_n1013_ = new_n203_ & new_n1012_;
  assign new_n1014_ = new_n1011_ & new_n1013_;
  assign new_n1015_ = ~new_n1009_ & ~new_n1014_;
  assign new_n1016_ = ~v36 & ~new_n1015_;
  assign new_n1017_ = ~v11 & new_n1016_;
  assign new_n1018_ = ~v10 & new_n1017_;
  assign new_n1019_ = ~v9 & new_n1018_;
  assign new_n1020_ = ~v3 & new_n1019_;
  assign new_n1021_ = ~v2 & new_n1020_;
  assign new_n1022_ = ~v1 & new_n1021_;
  assign new_n1023_ = ~new_n840_ & ~new_n1022_;
  assign \v41.11  = ~v8 & ~new_n1023_;
  assign new_n1025_ = ~v5 & new_n1006_;
  assign new_n1026_ = v4 & new_n1025_;
  assign new_n1027_ = ~new_n1001_ & ~new_n1026_;
  assign new_n1028_ = ~v0 & ~new_n1027_;
  assign new_n1029_ = ~new_n1014_ & ~new_n1028_;
  assign new_n1030_ = ~v36 & ~new_n1029_;
  assign new_n1031_ = ~v11 & new_n1030_;
  assign new_n1032_ = ~v10 & new_n1031_;
  assign new_n1033_ = ~v9 & new_n1032_;
  assign new_n1034_ = ~v8 & new_n1033_;
  assign new_n1035_ = ~v3 & new_n1034_;
  assign new_n1036_ = ~v2 & new_n1035_;
  assign \v41.12  = ~v1 & new_n1036_;
  assign new_n1038_ = v18 & ~v19;
  assign new_n1039_ = ~v17 & new_n1038_;
  assign new_n1040_ = new_n116_ & new_n1039_;
  assign new_n1041_ = ~new_n746_ & ~new_n1040_;
  assign new_n1042_ = ~v13 & ~new_n1041_;
  assign new_n1043_ = v13 & ~new_n962_;
  assign new_n1044_ = ~new_n1042_ & ~new_n1043_;
  assign new_n1045_ = v40 & ~new_n1044_;
  assign new_n1046_ = ~v5 & new_n1045_;
  assign new_n1047_ = ~v19 & ~new_n697_;
  assign new_n1048_ = v18 & new_n1047_;
  assign new_n1049_ = v17 & new_n1048_;
  assign new_n1050_ = ~v16 & new_n1049_;
  assign new_n1051_ = ~v15 & new_n1050_;
  assign new_n1052_ = ~v13 & new_n1051_;
  assign new_n1053_ = v5 & new_n1052_;
  assign new_n1054_ = ~new_n1046_ & ~new_n1053_;
  assign new_n1055_ = v12 & ~new_n1054_;
  assign new_n1056_ = v40 & ~new_n783_;
  assign new_n1057_ = ~v5 & new_n1056_;
  assign new_n1058_ = new_n203_ & new_n653_;
  assign new_n1059_ = ~new_n1057_ & ~new_n1058_;
  assign new_n1060_ = v16 & ~new_n1059_;
  assign new_n1061_ = ~v17 & new_n385_;
  assign new_n1062_ = ~v16 & new_n1061_;
  assign new_n1063_ = v15 & new_n1062_;
  assign new_n1064_ = ~v5 & new_n1063_;
  assign new_n1065_ = ~new_n1060_ & ~new_n1064_;
  assign new_n1066_ = v13 & ~new_n1065_;
  assign new_n1067_ = ~v12 & new_n1066_;
  assign new_n1068_ = ~new_n1055_ & ~new_n1067_;
  assign new_n1069_ = ~v4 & ~new_n1068_;
  assign new_n1070_ = ~v13 & new_n1003_;
  assign new_n1071_ = v12 & new_n1070_;
  assign new_n1072_ = v5 & new_n1071_;
  assign new_n1073_ = v4 & new_n1072_;
  assign new_n1074_ = ~new_n1069_ & ~new_n1073_;
  assign new_n1075_ = ~v0 & ~new_n1074_;
  assign new_n1076_ = new_n268_ & new_n1011_;
  assign new_n1077_ = ~new_n1075_ & ~new_n1076_;
  assign new_n1078_ = ~v36 & ~new_n1077_;
  assign new_n1079_ = ~v14 & new_n1078_;
  assign new_n1080_ = ~v11 & new_n1079_;
  assign new_n1081_ = ~v10 & new_n1080_;
  assign new_n1082_ = ~v9 & new_n1081_;
  assign new_n1083_ = ~v3 & new_n1082_;
  assign new_n1084_ = ~v2 & new_n1083_;
  assign new_n1085_ = ~v1 & new_n1084_;
  assign new_n1086_ = ~new_n840_ & ~new_n1085_;
  assign \v41.13  = ~v8 & ~new_n1086_;
  assign new_n1088_ = new_n249_ & new_n400_;
  assign new_n1089_ = new_n401_ & new_n403_;
  assign new_n1090_ = ~new_n1088_ & ~new_n1089_;
  assign new_n1091_ = v15 & ~new_n1090_;
  assign new_n1092_ = v1 & new_n1091_;
  assign new_n1093_ = ~v15 & new_n608_;
  assign new_n1094_ = ~v5 & new_n1093_;
  assign new_n1095_ = ~v4 & new_n1094_;
  assign new_n1096_ = ~v1 & new_n1095_;
  assign new_n1097_ = ~new_n1092_ & ~new_n1096_;
  assign new_n1098_ = ~v18 & ~new_n1097_;
  assign new_n1099_ = v16 & new_n340_;
  assign new_n1100_ = ~v15 & new_n1099_;
  assign new_n1101_ = ~v5 & new_n1100_;
  assign new_n1102_ = ~v4 & new_n1101_;
  assign new_n1103_ = ~v1 & new_n1102_;
  assign new_n1104_ = ~new_n1098_ & ~new_n1103_;
  assign new_n1105_ = ~v17 & ~new_n1104_;
  assign new_n1106_ = ~new_n165_ & ~new_n1038_;
  assign new_n1107_ = v17 & ~new_n1106_;
  assign new_n1108_ = v16 & new_n1107_;
  assign new_n1109_ = v16 & ~new_n1108_;
  assign new_n1110_ = ~v15 & ~new_n1109_;
  assign new_n1111_ = new_n117_ & new_n121_;
  assign new_n1112_ = ~new_n1110_ & ~new_n1111_;
  assign new_n1113_ = v40 & ~new_n1112_;
  assign new_n1114_ = ~v5 & new_n1113_;
  assign new_n1115_ = v5 & new_n116_;
  assign new_n1116_ = new_n203_ & new_n1115_;
  assign new_n1117_ = ~new_n1114_ & ~new_n1116_;
  assign new_n1118_ = ~v4 & ~new_n1117_;
  assign new_n1119_ = ~v1 & new_n1118_;
  assign new_n1120_ = ~new_n1105_ & ~new_n1119_;
  assign new_n1121_ = ~v12 & ~new_n1120_;
  assign new_n1122_ = v15 & ~new_n117_;
  assign new_n1123_ = v40 & ~new_n1122_;
  assign new_n1124_ = v12 & new_n1123_;
  assign new_n1125_ = ~v5 & new_n1124_;
  assign new_n1126_ = ~v4 & new_n1125_;
  assign new_n1127_ = ~v1 & new_n1126_;
  assign new_n1128_ = ~new_n1121_ & ~new_n1127_;
  assign new_n1129_ = v13 & ~new_n1128_;
  assign new_n1130_ = v4 & v15;
  assign new_n1131_ = new_n735_ & new_n1130_;
  assign new_n1132_ = ~v4 & new_n226_;
  assign new_n1133_ = v20 & v21;
  assign new_n1134_ = ~v19 & new_n1133_;
  assign new_n1135_ = new_n1132_ & new_n1134_;
  assign new_n1136_ = ~new_n1131_ & ~new_n1135_;
  assign new_n1137_ = v5 & ~new_n1136_;
  assign new_n1138_ = ~v15 & new_n976_;
  assign new_n1139_ = new_n189_ & ~new_n1138_;
  assign new_n1140_ = v40 & ~new_n1139_;
  assign new_n1141_ = ~v5 & new_n1140_;
  assign new_n1142_ = ~v4 & new_n1141_;
  assign new_n1143_ = ~new_n1137_ & ~new_n1142_;
  assign new_n1144_ = v18 & ~new_n1143_;
  assign new_n1145_ = v15 & v17;
  assign new_n1146_ = ~v15 & ~v17;
  assign new_n1147_ = ~new_n1145_ & ~new_n1146_;
  assign new_n1148_ = ~v38 & v39;
  assign new_n1149_ = v37 & new_n1148_;
  assign new_n1150_ = v17 & ~new_n1149_;
  assign new_n1151_ = ~v15 & new_n1150_;
  assign new_n1152_ = ~new_n246_ & ~new_n1151_;
  assign new_n1153_ = v19 & ~new_n1152_;
  assign new_n1154_ = new_n1147_ & ~new_n1153_;
  assign new_n1155_ = v40 & ~new_n1154_;
  assign new_n1156_ = ~v18 & new_n1155_;
  assign new_n1157_ = ~v5 & new_n1156_;
  assign new_n1158_ = ~v4 & new_n1157_;
  assign new_n1159_ = ~new_n1144_ & ~new_n1158_;
  assign new_n1160_ = ~v16 & ~new_n1159_;
  assign new_n1161_ = ~v19 & ~new_n741_;
  assign new_n1162_ = v17 & ~new_n1161_;
  assign new_n1163_ = ~new_n976_ & ~new_n1162_;
  assign new_n1164_ = ~v18 & ~new_n1163_;
  assign new_n1165_ = ~v18 & ~new_n1164_;
  assign new_n1166_ = v40 & ~new_n1165_;
  assign new_n1167_ = v16 & new_n1166_;
  assign new_n1168_ = ~v15 & new_n1167_;
  assign new_n1169_ = ~v5 & new_n1168_;
  assign new_n1170_ = ~v4 & new_n1169_;
  assign new_n1171_ = ~new_n1160_ & ~new_n1170_;
  assign new_n1172_ = ~v13 & ~new_n1171_;
  assign new_n1173_ = v12 & new_n1172_;
  assign new_n1174_ = ~v1 & new_n1173_;
  assign new_n1175_ = ~new_n1129_ & ~new_n1174_;
  assign new_n1176_ = ~v14 & ~new_n1175_;
  assign new_n1177_ = v18 & ~new_n1038_;
  assign new_n1178_ = ~v16 & ~new_n1177_;
  assign new_n1179_ = v16 & new_n171_;
  assign new_n1180_ = ~new_n1178_ & ~new_n1179_;
  assign new_n1181_ = ~v17 & ~new_n1180_;
  assign new_n1182_ = v13 & new_n1181_;
  assign new_n1183_ = v13 & ~new_n1182_;
  assign new_n1184_ = ~v17 & ~new_n156_;
  assign new_n1185_ = v15 & new_n1184_;
  assign new_n1186_ = ~v15 & new_n209_;
  assign new_n1187_ = ~new_n1185_ & ~new_n1186_;
  assign new_n1188_ = v18 & ~new_n1187_;
  assign new_n1189_ = v17 & new_n165_;
  assign new_n1190_ = new_n201_ & new_n1189_;
  assign new_n1191_ = ~new_n1188_ & ~new_n1190_;
  assign new_n1192_ = v13 & ~new_n1191_;
  assign new_n1193_ = new_n1183_ & ~new_n1192_;
  assign new_n1194_ = v12 & ~new_n1193_;
  assign new_n1195_ = ~v15 & new_n883_;
  assign new_n1196_ = ~v13 & new_n1195_;
  assign new_n1197_ = ~v13 & ~new_n1196_;
  assign new_n1198_ = ~v12 & ~new_n1197_;
  assign new_n1199_ = ~new_n1194_ & ~new_n1198_;
  assign new_n1200_ = v40 & ~new_n1199_;
  assign new_n1201_ = v14 & new_n1200_;
  assign new_n1202_ = ~v5 & new_n1201_;
  assign new_n1203_ = ~v4 & new_n1202_;
  assign new_n1204_ = ~v1 & new_n1203_;
  assign new_n1205_ = ~new_n1176_ & ~new_n1204_;
  assign new_n1206_ = ~v3 & ~new_n1205_;
  assign new_n1207_ = v23 & ~v24;
  assign new_n1208_ = v22 & new_n1207_;
  assign new_n1209_ = ~new_n692_ & ~new_n1208_;
  assign new_n1210_ = v4 & v27;
  assign new_n1211_ = ~v4 & ~v27;
  assign new_n1212_ = ~new_n1210_ & ~new_n1211_;
  assign new_n1213_ = ~new_n1209_ & ~new_n1212_;
  assign new_n1214_ = v23 & ~v25;
  assign new_n1215_ = v23 & ~new_n1214_;
  assign new_n1216_ = ~v27 & ~new_n1215_;
  assign new_n1217_ = v24 & new_n1216_;
  assign new_n1218_ = v22 & new_n1217_;
  assign new_n1219_ = ~v4 & new_n1218_;
  assign new_n1220_ = ~new_n1213_ & ~new_n1219_;
  assign new_n1221_ = ~v5 & ~new_n1220_;
  assign new_n1222_ = v24 & v27;
  assign new_n1223_ = ~new_n719_ & ~new_n1222_;
  assign new_n1224_ = ~v23 & ~new_n1223_;
  assign new_n1225_ = v25 & ~v27;
  assign new_n1226_ = ~v27 & ~new_n1225_;
  assign new_n1227_ = v24 & ~new_n1226_;
  assign new_n1228_ = v23 & new_n1227_;
  assign new_n1229_ = ~new_n1224_ & ~new_n1228_;
  assign new_n1230_ = v22 & ~new_n1229_;
  assign new_n1231_ = ~v22 & new_n719_;
  assign new_n1232_ = ~new_n1230_ & ~new_n1231_;
  assign new_n1233_ = v5 & ~new_n1232_;
  assign new_n1234_ = ~v4 & new_n1233_;
  assign new_n1235_ = ~new_n1221_ & ~new_n1234_;
  assign new_n1236_ = v21 & ~new_n1235_;
  assign new_n1237_ = ~v20 & new_n1236_;
  assign new_n1238_ = ~v21 & ~v27;
  assign new_n1239_ = v20 & new_n1238_;
  assign new_n1240_ = new_n403_ & new_n1239_;
  assign new_n1241_ = ~new_n1237_ & ~new_n1240_;
  assign new_n1242_ = v18 & ~new_n1241_;
  assign new_n1243_ = ~v5 & ~v18;
  assign new_n1244_ = ~v4 & new_n1243_;
  assign new_n1245_ = ~new_n1242_ & ~new_n1244_;
  assign new_n1246_ = ~v19 & ~new_n1245_;
  assign new_n1247_ = v17 & new_n1246_;
  assign new_n1248_ = ~v16 & new_n1247_;
  assign new_n1249_ = ~v15 & new_n1248_;
  assign new_n1250_ = ~v14 & new_n1249_;
  assign new_n1251_ = ~v13 & new_n1250_;
  assign new_n1252_ = v12 & new_n1251_;
  assign new_n1253_ = v3 & new_n1252_;
  assign new_n1254_ = ~v1 & new_n1253_;
  assign new_n1255_ = ~new_n1206_ & ~new_n1254_;
  assign new_n1256_ = ~v0 & ~new_n1255_;
  assign new_n1257_ = v3 & ~new_n248_;
  assign new_n1258_ = ~v3 & v15;
  assign new_n1259_ = ~v17 & new_n165_;
  assign new_n1260_ = new_n1258_ & new_n1259_;
  assign new_n1261_ = ~new_n1257_ & ~new_n1260_;
  assign new_n1262_ = v16 & ~new_n1261_;
  assign new_n1263_ = ~v3 & new_n117_;
  assign new_n1264_ = new_n172_ & new_n1263_;
  assign new_n1265_ = ~new_n1262_ & ~new_n1264_;
  assign new_n1266_ = v13 & ~new_n1265_;
  assign new_n1267_ = ~v12 & new_n1266_;
  assign new_n1268_ = new_n338_ & new_n766_;
  assign new_n1269_ = new_n210_ & new_n1268_;
  assign new_n1270_ = ~new_n1267_ & ~new_n1269_;
  assign new_n1271_ = ~v14 & ~new_n1270_;
  assign new_n1272_ = ~v5 & new_n1271_;
  assign new_n1273_ = ~v4 & new_n1272_;
  assign new_n1274_ = ~v1 & new_n1273_;
  assign new_n1275_ = v0 & new_n1274_;
  assign new_n1276_ = ~new_n1256_ & ~new_n1275_;
  assign new_n1277_ = ~v2 & ~new_n1276_;
  assign new_n1278_ = ~v5 & new_n684_;
  assign new_n1279_ = v5 & new_n679_;
  assign new_n1280_ = ~new_n1278_ & ~new_n1279_;
  assign new_n1281_ = v27 & ~new_n1280_;
  assign new_n1282_ = ~v19 & new_n1281_;
  assign new_n1283_ = v18 & new_n1282_;
  assign new_n1284_ = v17 & new_n1283_;
  assign new_n1285_ = ~v16 & new_n1284_;
  assign new_n1286_ = ~v15 & new_n1285_;
  assign new_n1287_ = ~v14 & new_n1286_;
  assign new_n1288_ = ~v13 & new_n1287_;
  assign new_n1289_ = v12 & new_n1288_;
  assign new_n1290_ = ~v4 & new_n1289_;
  assign new_n1291_ = ~v3 & new_n1290_;
  assign new_n1292_ = v2 & new_n1291_;
  assign new_n1293_ = ~v1 & new_n1292_;
  assign new_n1294_ = ~v0 & new_n1293_;
  assign new_n1295_ = ~new_n1277_ & ~new_n1294_;
  assign new_n1296_ = ~v36 & ~new_n1295_;
  assign new_n1297_ = ~v11 & new_n1296_;
  assign new_n1298_ = ~v10 & new_n1297_;
  assign new_n1299_ = ~v9 & new_n1298_;
  assign \v41.14  = ~v8 & new_n1299_;
  assign new_n1301_ = v8 & ~v36;
  assign new_n1302_ = ~v5 & new_n1301_;
  assign new_n1303_ = ~v4 & new_n1302_;
  assign new_n1304_ = ~v3 & new_n1303_;
  assign new_n1305_ = ~v2 & new_n1304_;
  assign new_n1306_ = ~v1 & new_n1305_;
  assign new_n1307_ = ~v0 & new_n1306_;
  assign new_n1308_ = ~v8 & v10;
  assign new_n1309_ = ~new_n1307_ & ~new_n1308_;
  assign new_n1310_ = ~v9 & ~new_n1309_;
  assign new_n1311_ = v9 & ~v10;
  assign \v41.71  = ~v8 & new_n1311_;
  assign new_n1313_ = ~new_n1310_ & ~\v41.71 ;
  assign new_n1314_ = ~v16 & new_n843_;
  assign new_n1315_ = ~v16 & ~new_n1314_;
  assign new_n1316_ = v13 & ~new_n1315_;
  assign new_n1317_ = v13 & ~new_n1316_;
  assign new_n1318_ = ~v17 & ~new_n1317_;
  assign new_n1319_ = v13 & ~new_n220_;
  assign new_n1320_ = v17 & ~new_n1319_;
  assign new_n1321_ = ~new_n1318_ & ~new_n1320_;
  assign new_n1322_ = v18 & ~new_n1321_;
  assign new_n1323_ = v13 & new_n673_;
  assign new_n1324_ = v13 & ~new_n1323_;
  assign new_n1325_ = ~v18 & ~new_n1324_;
  assign new_n1326_ = ~new_n1322_ & ~new_n1325_;
  assign new_n1327_ = v15 & ~new_n1326_;
  assign new_n1328_ = ~new_n766_ & ~new_n1327_;
  assign new_n1329_ = ~v14 & ~new_n1328_;
  assign new_n1330_ = ~v5 & new_n1329_;
  assign new_n1331_ = ~v15 & ~new_n116_;
  assign new_n1332_ = ~new_n1186_ & new_n1331_;
  assign new_n1333_ = v14 & ~new_n1332_;
  assign new_n1334_ = ~v13 & new_n1333_;
  assign new_n1335_ = v5 & new_n1334_;
  assign new_n1336_ = ~new_n1330_ & ~new_n1335_;
  assign new_n1337_ = ~v12 & ~new_n1336_;
  assign new_n1338_ = v13 & v14;
  assign new_n1339_ = ~v14 & v16;
  assign new_n1340_ = ~v13 & new_n1339_;
  assign new_n1341_ = ~new_n1338_ & ~new_n1340_;
  assign new_n1342_ = v17 & ~new_n1341_;
  assign new_n1343_ = ~v13 & ~v14;
  assign new_n1344_ = new_n164_ & new_n1343_;
  assign new_n1345_ = ~new_n1342_ & ~new_n1344_;
  assign new_n1346_ = v15 & ~new_n1345_;
  assign new_n1347_ = new_n674_ & new_n1338_;
  assign new_n1348_ = ~new_n1346_ & ~new_n1347_;
  assign new_n1349_ = v13 & new_n900_;
  assign new_n1350_ = v16 & new_n753_;
  assign new_n1351_ = new_n1349_ & new_n1350_;
  assign new_n1352_ = new_n1348_ & ~new_n1351_;
  assign new_n1353_ = v12 & ~new_n1352_;
  assign new_n1354_ = v5 & new_n1353_;
  assign new_n1355_ = ~new_n1337_ & ~new_n1354_;
  assign new_n1356_ = ~v14 & v15;
  assign new_n1357_ = ~v13 & new_n1356_;
  assign new_n1358_ = ~v16 & new_n517_;
  assign new_n1359_ = new_n1357_ & new_n1358_;
  assign new_n1360_ = new_n124_ & new_n1349_;
  assign new_n1361_ = ~new_n1359_ & ~new_n1360_;
  assign new_n1362_ = v5 & ~new_n1361_;
  assign new_n1363_ = ~v5 & ~v13;
  assign new_n1364_ = new_n383_ & new_n1363_;
  assign new_n1365_ = v37 & ~v38;
  assign new_n1366_ = ~v18 & new_n1365_;
  assign new_n1367_ = new_n209_ & new_n1366_;
  assign new_n1368_ = new_n1364_ & new_n1367_;
  assign new_n1369_ = ~new_n1362_ & ~new_n1368_;
  assign new_n1370_ = v19 & ~new_n1369_;
  assign new_n1371_ = ~v19 & new_n843_;
  assign new_n1372_ = ~v18 & new_n1371_;
  assign new_n1373_ = ~v17 & new_n1372_;
  assign new_n1374_ = ~v16 & new_n1373_;
  assign new_n1375_ = v15 & new_n1374_;
  assign new_n1376_ = ~v14 & new_n1375_;
  assign new_n1377_ = ~v13 & new_n1376_;
  assign new_n1378_ = ~v5 & new_n1377_;
  assign new_n1379_ = ~new_n1370_ & ~new_n1378_;
  assign new_n1380_ = v12 & ~new_n1379_;
  assign new_n1381_ = new_n1355_ & ~new_n1380_;
  assign new_n1382_ = v40 & ~new_n1381_;
  assign new_n1383_ = ~v36 & new_n1382_;
  assign new_n1384_ = ~v11 & new_n1383_;
  assign new_n1385_ = ~v10 & new_n1384_;
  assign new_n1386_ = ~v9 & new_n1385_;
  assign new_n1387_ = ~v4 & new_n1386_;
  assign new_n1388_ = ~v3 & new_n1387_;
  assign new_n1389_ = ~v2 & new_n1388_;
  assign new_n1390_ = ~v1 & new_n1389_;
  assign new_n1391_ = ~v0 & new_n1390_;
  assign new_n1392_ = v9 & new_n838_;
  assign new_n1393_ = ~new_n1391_ & ~new_n1392_;
  assign new_n1394_ = ~v8 & ~new_n1393_;
  assign \v41.15  = ~new_n1313_ | new_n1394_;
  assign new_n1396_ = v9 & v10;
  assign new_n1397_ = ~v4 & ~new_n672_;
  assign new_n1398_ = ~v4 & ~new_n1397_;
  assign new_n1399_ = ~v14 & ~new_n1398_;
  assign new_n1400_ = v13 & new_n1399_;
  assign new_n1401_ = ~v13 & new_n333_;
  assign new_n1402_ = new_n169_ & new_n1401_;
  assign new_n1403_ = ~new_n1400_ & ~new_n1402_;
  assign new_n1404_ = ~v18 & ~new_n1403_;
  assign new_n1405_ = ~v4 & new_n1363_;
  assign new_n1406_ = new_n341_ & new_n1405_;
  assign new_n1407_ = ~new_n1404_ & ~new_n1406_;
  assign new_n1408_ = ~v17 & ~new_n1407_;
  assign new_n1409_ = v17 & v40;
  assign new_n1410_ = v14 & new_n1409_;
  assign new_n1411_ = ~v13 & new_n1410_;
  assign new_n1412_ = ~v5 & new_n1411_;
  assign new_n1413_ = ~v4 & new_n1412_;
  assign new_n1414_ = ~new_n1408_ & ~new_n1413_;
  assign new_n1415_ = v15 & ~new_n1414_;
  assign new_n1416_ = ~v17 & ~new_n119_;
  assign new_n1417_ = v40 & ~new_n1416_;
  assign new_n1418_ = ~v15 & new_n1417_;
  assign new_n1419_ = v14 & new_n1418_;
  assign new_n1420_ = ~v13 & new_n1419_;
  assign new_n1421_ = ~v5 & new_n1420_;
  assign new_n1422_ = ~v4 & new_n1421_;
  assign new_n1423_ = ~new_n1415_ & ~new_n1422_;
  assign new_n1424_ = ~v12 & ~new_n1423_;
  assign new_n1425_ = v15 & new_n1409_;
  assign new_n1426_ = v14 & new_n1425_;
  assign new_n1427_ = v13 & new_n1426_;
  assign new_n1428_ = v12 & new_n1427_;
  assign new_n1429_ = ~v5 & new_n1428_;
  assign new_n1430_ = ~v4 & new_n1429_;
  assign new_n1431_ = ~new_n1424_ & ~new_n1430_;
  assign new_n1432_ = ~v3 & ~new_n1431_;
  assign new_n1433_ = ~v14 & new_n138_;
  assign new_n1434_ = v13 & new_n1433_;
  assign new_n1435_ = ~v12 & new_n1434_;
  assign new_n1436_ = v3 & new_n1435_;
  assign new_n1437_ = ~new_n1432_ & ~new_n1436_;
  assign new_n1438_ = ~v2 & ~new_n1437_;
  assign new_n1439_ = v2 & new_n1435_;
  assign new_n1440_ = ~new_n1438_ & ~new_n1439_;
  assign new_n1441_ = ~v1 & ~new_n1440_;
  assign new_n1442_ = v1 & ~v2;
  assign new_n1443_ = new_n381_ & new_n1442_;
  assign new_n1444_ = v13 & ~v14;
  assign new_n1445_ = ~v12 & new_n1444_;
  assign new_n1446_ = new_n138_ & new_n1445_;
  assign new_n1447_ = new_n1443_ & new_n1446_;
  assign new_n1448_ = ~new_n1441_ & ~new_n1447_;
  assign new_n1449_ = ~v18 & ~new_n1398_;
  assign new_n1450_ = v17 & new_n1449_;
  assign new_n1451_ = ~v39 & ~new_n844_;
  assign new_n1452_ = ~v38 & new_n1451_;
  assign new_n1453_ = v40 & ~new_n1452_;
  assign new_n1454_ = v18 & new_n1453_;
  assign new_n1455_ = ~v17 & new_n1454_;
  assign new_n1456_ = ~v5 & new_n1455_;
  assign new_n1457_ = ~v4 & new_n1456_;
  assign new_n1458_ = ~new_n1450_ & ~new_n1457_;
  assign new_n1459_ = ~v16 & ~new_n1458_;
  assign new_n1460_ = v13 & new_n1459_;
  assign new_n1461_ = ~v12 & new_n1460_;
  assign new_n1462_ = ~v13 & new_n608_;
  assign new_n1463_ = v12 & new_n1462_;
  assign new_n1464_ = ~v5 & new_n1463_;
  assign new_n1465_ = ~v4 & new_n1464_;
  assign new_n1466_ = ~new_n1461_ & ~new_n1465_;
  assign new_n1467_ = v15 & ~new_n1466_;
  assign new_n1468_ = ~v14 & new_n1467_;
  assign new_n1469_ = ~v17 & ~new_n753_;
  assign new_n1470_ = v13 & ~new_n1469_;
  assign new_n1471_ = v12 & new_n1470_;
  assign new_n1472_ = ~v12 & ~v13;
  assign new_n1473_ = new_n753_ & new_n1472_;
  assign new_n1474_ = ~new_n1471_ & ~new_n1473_;
  assign new_n1475_ = v40 & ~new_n1474_;
  assign new_n1476_ = v16 & new_n1475_;
  assign new_n1477_ = ~v15 & new_n1476_;
  assign new_n1478_ = v14 & new_n1477_;
  assign new_n1479_ = ~v5 & new_n1478_;
  assign new_n1480_ = ~v4 & new_n1479_;
  assign new_n1481_ = ~new_n1468_ & ~new_n1480_;
  assign new_n1482_ = ~v3 & ~new_n1481_;
  assign new_n1483_ = v3 & ~v4;
  assign new_n1484_ = ~v5 & new_n849_;
  assign new_n1485_ = new_n1483_ & new_n1484_;
  assign new_n1486_ = ~v16 & new_n754_;
  assign new_n1487_ = new_n1356_ & new_n1486_;
  assign new_n1488_ = new_n1485_ & new_n1487_;
  assign new_n1489_ = ~new_n1482_ & ~new_n1488_;
  assign new_n1490_ = ~v1 & ~new_n1489_;
  assign new_n1491_ = v1 & ~v3;
  assign new_n1492_ = v5 & ~v12;
  assign new_n1493_ = ~v4 & new_n1492_;
  assign new_n1494_ = new_n1491_ & new_n1493_;
  assign new_n1495_ = v13 & new_n1356_;
  assign new_n1496_ = new_n124_ & new_n1495_;
  assign new_n1497_ = new_n1494_ & new_n1496_;
  assign new_n1498_ = ~new_n1490_ & ~new_n1497_;
  assign new_n1499_ = ~v2 & ~new_n1498_;
  assign new_n1500_ = new_n1448_ & ~new_n1499_;
  assign new_n1501_ = ~new_n304_ & ~new_n674_;
  assign new_n1502_ = ~new_n843_ & ~new_n1501_;
  assign new_n1503_ = new_n246_ & new_n844_;
  assign new_n1504_ = ~new_n226_ & ~new_n1503_;
  assign new_n1505_ = ~v16 & ~new_n1504_;
  assign new_n1506_ = ~new_n1502_ & ~new_n1505_;
  assign new_n1507_ = ~v18 & ~new_n1506_;
  assign new_n1508_ = new_n681_ & ~new_n1208_;
  assign new_n1509_ = v21 & ~new_n1508_;
  assign new_n1510_ = ~v20 & new_n1509_;
  assign new_n1511_ = ~new_n679_ & ~new_n1510_;
  assign new_n1512_ = v23 & v24;
  assign new_n1513_ = v22 & new_n1512_;
  assign new_n1514_ = ~v20 & new_n1513_;
  assign new_n1515_ = ~v20 & ~new_n1514_;
  assign new_n1516_ = v21 & ~new_n1515_;
  assign new_n1517_ = new_n1511_ & ~new_n1516_;
  assign new_n1518_ = v18 & ~new_n1517_;
  assign new_n1519_ = v17 & new_n1518_;
  assign new_n1520_ = ~v16 & new_n1519_;
  assign new_n1521_ = ~v15 & new_n1520_;
  assign new_n1522_ = ~new_n1507_ & ~new_n1521_;
  assign new_n1523_ = v40 & ~new_n1522_;
  assign new_n1524_ = ~v5 & new_n1523_;
  assign new_n1525_ = v21 & new_n1513_;
  assign new_n1526_ = ~v20 & new_n1525_;
  assign new_n1527_ = new_n1511_ & ~new_n1526_;
  assign new_n1528_ = v18 & ~new_n1527_;
  assign new_n1529_ = v18 & ~new_n1528_;
  assign new_n1530_ = v17 & ~new_n1529_;
  assign new_n1531_ = ~v16 & new_n1530_;
  assign new_n1532_ = ~v15 & new_n1531_;
  assign new_n1533_ = v5 & new_n1532_;
  assign new_n1534_ = ~new_n1524_ & ~new_n1533_;
  assign new_n1535_ = ~v4 & ~new_n1534_;
  assign new_n1536_ = v4 & new_n1532_;
  assign new_n1537_ = ~new_n1535_ & ~new_n1536_;
  assign new_n1538_ = ~v3 & ~new_n1537_;
  assign new_n1539_ = v24 & ~new_n1222_;
  assign new_n1540_ = ~new_n681_ & ~new_n1539_;
  assign new_n1541_ = ~v24 & v27;
  assign new_n1542_ = ~new_n1227_ & ~new_n1541_;
  assign new_n1543_ = v23 & ~new_n1542_;
  assign new_n1544_ = v22 & new_n1543_;
  assign new_n1545_ = ~new_n1540_ & ~new_n1544_;
  assign new_n1546_ = ~v5 & ~new_n1545_;
  assign new_n1547_ = v24 & ~new_n692_;
  assign new_n1548_ = v27 & ~new_n1547_;
  assign new_n1549_ = v5 & new_n1548_;
  assign new_n1550_ = ~new_n1546_ & ~new_n1549_;
  assign new_n1551_ = ~v4 & ~new_n1550_;
  assign new_n1552_ = v27 & ~new_n681_;
  assign new_n1553_ = ~v24 & new_n1552_;
  assign new_n1554_ = v4 & new_n1553_;
  assign new_n1555_ = ~new_n1551_ & ~new_n1554_;
  assign new_n1556_ = v21 & ~new_n1555_;
  assign new_n1557_ = ~v20 & new_n1556_;
  assign new_n1558_ = ~v5 & ~v27;
  assign new_n1559_ = ~v4 & new_n1558_;
  assign new_n1560_ = ~v27 & ~new_n1559_;
  assign new_n1561_ = ~v21 & ~new_n1560_;
  assign new_n1562_ = v20 & new_n1561_;
  assign new_n1563_ = ~new_n1557_ & ~new_n1562_;
  assign new_n1564_ = v18 & ~new_n1563_;
  assign new_n1565_ = v17 & new_n1564_;
  assign new_n1566_ = ~v16 & new_n1565_;
  assign new_n1567_ = ~v15 & new_n1566_;
  assign new_n1568_ = v3 & new_n1567_;
  assign new_n1569_ = ~new_n1538_ & ~new_n1568_;
  assign new_n1570_ = ~v19 & ~new_n1569_;
  assign new_n1571_ = v15 & v18;
  assign new_n1572_ = ~v18 & v39;
  assign new_n1573_ = new_n226_ & new_n1572_;
  assign new_n1574_ = ~new_n1571_ & ~new_n1573_;
  assign new_n1575_ = v40 & ~new_n1574_;
  assign new_n1576_ = ~v5 & new_n1575_;
  assign new_n1577_ = new_n607_ & new_n753_;
  assign new_n1578_ = ~new_n1576_ & ~new_n1577_;
  assign new_n1579_ = ~v4 & ~new_n1578_;
  assign new_n1580_ = v15 & new_n753_;
  assign new_n1581_ = new_n249_ & new_n1580_;
  assign new_n1582_ = ~new_n1579_ & ~new_n1581_;
  assign new_n1583_ = v19 & ~new_n1582_;
  assign new_n1584_ = ~v16 & new_n1583_;
  assign new_n1585_ = ~v3 & new_n1584_;
  assign new_n1586_ = ~new_n1570_ & ~new_n1585_;
  assign new_n1587_ = ~v13 & ~new_n1586_;
  assign new_n1588_ = v12 & new_n1587_;
  assign new_n1589_ = ~v15 & new_n400_;
  assign new_n1590_ = v15 & new_n401_;
  assign new_n1591_ = ~new_n1589_ & ~new_n1590_;
  assign new_n1592_ = ~new_n672_ & ~new_n1591_;
  assign new_n1593_ = v18 & new_n1592_;
  assign new_n1594_ = ~v5 & new_n116_;
  assign new_n1595_ = ~v19 & v40;
  assign new_n1596_ = ~v18 & new_n1595_;
  assign new_n1597_ = new_n1594_ & new_n1596_;
  assign new_n1598_ = ~new_n1593_ & ~new_n1597_;
  assign new_n1599_ = ~v4 & ~new_n1598_;
  assign new_n1600_ = v18 & ~new_n1591_;
  assign new_n1601_ = v4 & new_n1600_;
  assign new_n1602_ = ~new_n1599_ & ~new_n1601_;
  assign new_n1603_ = ~v3 & ~new_n1602_;
  assign new_n1604_ = v16 & new_n120_;
  assign new_n1605_ = ~v15 & new_n1604_;
  assign new_n1606_ = v3 & new_n1605_;
  assign new_n1607_ = ~new_n1603_ & ~new_n1606_;
  assign new_n1608_ = v17 & ~new_n1607_;
  assign new_n1609_ = v13 & new_n1608_;
  assign new_n1610_ = ~v12 & new_n1609_;
  assign new_n1611_ = ~new_n1588_ & ~new_n1610_;
  assign new_n1612_ = ~v1 & ~new_n1611_;
  assign new_n1613_ = ~v3 & new_n116_;
  assign new_n1614_ = new_n121_ & new_n1613_;
  assign new_n1615_ = ~new_n548_ & ~new_n1614_;
  assign new_n1616_ = v4 & new_n159_;
  assign new_n1617_ = ~v3 & new_n1616_;
  assign new_n1618_ = new_n1615_ & ~new_n1617_;
  assign new_n1619_ = new_n256_ & new_n607_;
  assign new_n1620_ = new_n260_ & new_n1619_;
  assign new_n1621_ = new_n1618_ & ~new_n1620_;
  assign new_n1622_ = v13 & ~new_n1621_;
  assign new_n1623_ = ~v12 & new_n1622_;
  assign new_n1624_ = v1 & new_n1623_;
  assign new_n1625_ = ~new_n1612_ & ~new_n1624_;
  assign new_n1626_ = ~v2 & ~new_n1625_;
  assign new_n1627_ = v1 & ~new_n160_;
  assign new_n1628_ = ~v1 & new_n116_;
  assign new_n1629_ = new_n121_ & new_n1628_;
  assign new_n1630_ = ~new_n1627_ & ~new_n1629_;
  assign new_n1631_ = v13 & ~new_n1630_;
  assign new_n1632_ = ~v12 & new_n1631_;
  assign new_n1633_ = ~v1 & new_n256_;
  assign new_n1634_ = ~v5 & v12;
  assign new_n1635_ = new_n766_ & new_n1634_;
  assign new_n1636_ = new_n1633_ & new_n1635_;
  assign new_n1637_ = ~v19 & v20;
  assign new_n1638_ = ~v21 & v27;
  assign new_n1639_ = new_n1637_ & new_n1638_;
  assign new_n1640_ = new_n1358_ & new_n1639_;
  assign new_n1641_ = new_n1636_ & new_n1640_;
  assign new_n1642_ = ~new_n1632_ & ~new_n1641_;
  assign new_n1643_ = v2 & ~new_n1642_;
  assign new_n1644_ = ~new_n1626_ & ~new_n1643_;
  assign new_n1645_ = ~v14 & ~new_n1644_;
  assign new_n1646_ = v12 & v13;
  assign new_n1647_ = new_n900_ & new_n1646_;
  assign new_n1648_ = v19 & v40;
  assign new_n1649_ = ~v18 & new_n1648_;
  assign new_n1650_ = new_n164_ & new_n1649_;
  assign new_n1651_ = new_n1647_ & new_n1650_;
  assign new_n1652_ = v40 & ~new_n1651_;
  assign new_n1653_ = ~v5 & ~new_n1652_;
  assign new_n1654_ = ~v4 & new_n1653_;
  assign new_n1655_ = ~v3 & new_n1654_;
  assign new_n1656_ = ~v2 & new_n1655_;
  assign new_n1657_ = ~v1 & new_n1656_;
  assign new_n1658_ = ~new_n1645_ & ~new_n1657_;
  assign new_n1659_ = new_n1500_ & new_n1658_;
  assign new_n1660_ = ~v0 & ~new_n1659_;
  assign new_n1661_ = v16 & ~new_n248_;
  assign new_n1662_ = ~new_n632_ & ~new_n1661_;
  assign new_n1663_ = ~v14 & ~new_n1662_;
  assign new_n1664_ = v13 & new_n1663_;
  assign new_n1665_ = ~v12 & new_n1664_;
  assign new_n1666_ = ~v3 & new_n1665_;
  assign new_n1667_ = ~v2 & new_n1666_;
  assign new_n1668_ = ~v1 & new_n1667_;
  assign new_n1669_ = v0 & new_n1668_;
  assign new_n1670_ = ~new_n1660_ & ~new_n1669_;
  assign new_n1671_ = ~v36 & ~new_n1670_;
  assign new_n1672_ = ~v36 & ~new_n1671_;
  assign new_n1673_ = ~v11 & ~new_n1672_;
  assign new_n1674_ = ~v10 & new_n1673_;
  assign new_n1675_ = ~v9 & new_n1674_;
  assign new_n1676_ = ~new_n1396_ & ~new_n1675_;
  assign \v41.16  = ~v8 & ~new_n1676_;
  assign new_n1678_ = ~v13 & ~v18;
  assign new_n1679_ = ~v12 & new_n1678_;
  assign new_n1680_ = new_n120_ & new_n1646_;
  assign new_n1681_ = ~new_n1679_ & ~new_n1680_;
  assign new_n1682_ = ~v16 & ~new_n1681_;
  assign new_n1683_ = ~v15 & new_n1682_;
  assign new_n1684_ = v15 & new_n400_;
  assign new_n1685_ = v13 & new_n1684_;
  assign new_n1686_ = v12 & new_n1685_;
  assign new_n1687_ = ~new_n1683_ & ~new_n1686_;
  assign new_n1688_ = ~v17 & ~new_n1687_;
  assign new_n1689_ = v13 & ~v15;
  assign new_n1690_ = v12 & new_n1689_;
  assign new_n1691_ = new_n210_ & new_n1690_;
  assign new_n1692_ = ~new_n1688_ & ~new_n1691_;
  assign new_n1693_ = v14 & ~new_n1692_;
  assign new_n1694_ = v13 & v15;
  assign new_n1695_ = new_n766_ & new_n1259_;
  assign new_n1696_ = ~new_n1694_ & ~new_n1695_;
  assign new_n1697_ = v16 & ~new_n1696_;
  assign new_n1698_ = ~v14 & new_n1697_;
  assign new_n1699_ = v12 & new_n1698_;
  assign new_n1700_ = ~new_n1693_ & ~new_n1699_;
  assign new_n1701_ = v40 & ~new_n1700_;
  assign new_n1702_ = ~v36 & new_n1701_;
  assign new_n1703_ = ~v11 & new_n1702_;
  assign new_n1704_ = ~v10 & new_n1703_;
  assign new_n1705_ = ~v9 & new_n1704_;
  assign new_n1706_ = ~v8 & new_n1705_;
  assign new_n1707_ = ~v5 & new_n1706_;
  assign new_n1708_ = ~v4 & new_n1707_;
  assign new_n1709_ = ~v3 & new_n1708_;
  assign new_n1710_ = ~v2 & new_n1709_;
  assign new_n1711_ = ~v1 & new_n1710_;
  assign \v41.17  = ~v0 & new_n1711_;
  assign new_n1713_ = ~v17 & new_n120_;
  assign new_n1714_ = ~new_n203_ & ~new_n1713_;
  assign new_n1715_ = v13 & ~new_n1714_;
  assign new_n1716_ = v12 & new_n1715_;
  assign new_n1717_ = ~v13 & new_n119_;
  assign new_n1718_ = ~v12 & new_n1717_;
  assign new_n1719_ = ~new_n1716_ & ~new_n1718_;
  assign new_n1720_ = v14 & ~new_n1719_;
  assign new_n1721_ = ~v14 & v17;
  assign new_n1722_ = new_n265_ & new_n1721_;
  assign new_n1723_ = new_n165_ & new_n1365_;
  assign new_n1724_ = new_n1722_ & new_n1723_;
  assign new_n1725_ = ~new_n1720_ & ~new_n1724_;
  assign new_n1726_ = ~v15 & ~new_n1725_;
  assign new_n1727_ = v13 & v18;
  assign new_n1728_ = ~v12 & new_n1727_;
  assign new_n1729_ = new_n171_ & new_n265_;
  assign new_n1730_ = ~new_n1728_ & ~new_n1729_;
  assign new_n1731_ = ~v39 & ~new_n1730_;
  assign new_n1732_ = ~v38 & new_n1731_;
  assign new_n1733_ = v37 & new_n1732_;
  assign new_n1734_ = ~v17 & new_n1733_;
  assign new_n1735_ = v15 & new_n1734_;
  assign new_n1736_ = ~v14 & new_n1735_;
  assign new_n1737_ = ~new_n1726_ & ~new_n1736_;
  assign new_n1738_ = v40 & ~new_n1737_;
  assign new_n1739_ = ~v16 & new_n1738_;
  assign new_n1740_ = ~v11 & new_n1739_;
  assign new_n1741_ = ~v10 & new_n1740_;
  assign new_n1742_ = ~v8 & new_n1741_;
  assign new_n1743_ = ~v8 & ~new_n1742_;
  assign new_n1744_ = ~v3 & ~new_n1743_;
  assign new_n1745_ = v17 & ~new_n1177_;
  assign new_n1746_ = ~v16 & new_n1745_;
  assign new_n1747_ = v15 & new_n1746_;
  assign new_n1748_ = ~v14 & new_n1747_;
  assign new_n1749_ = v13 & new_n1748_;
  assign new_n1750_ = ~v12 & new_n1749_;
  assign new_n1751_ = ~v11 & new_n1750_;
  assign new_n1752_ = ~v10 & new_n1751_;
  assign new_n1753_ = ~v8 & new_n1752_;
  assign new_n1754_ = v3 & new_n1753_;
  assign new_n1755_ = ~new_n1744_ & ~new_n1754_;
  assign new_n1756_ = ~v36 & ~new_n1755_;
  assign new_n1757_ = ~v5 & new_n1756_;
  assign new_n1758_ = ~v4 & new_n1757_;
  assign new_n1759_ = ~v2 & new_n1758_;
  assign new_n1760_ = ~v1 & new_n1759_;
  assign new_n1761_ = ~v0 & new_n1760_;
  assign new_n1762_ = ~new_n1308_ & ~new_n1761_;
  assign new_n1763_ = ~v9 & ~new_n1762_;
  assign new_n1764_ = ~v8 & new_n840_;
  assign \v41.18  = new_n1763_ | new_n1764_;
  assign new_n1766_ = ~v13 & new_n900_;
  assign new_n1767_ = ~v16 & new_n119_;
  assign new_n1768_ = new_n1766_ & new_n1767_;
  assign new_n1769_ = ~new_n1329_ & ~new_n1768_;
  assign new_n1770_ = ~v12 & ~new_n1769_;
  assign new_n1771_ = v15 & v16;
  assign new_n1772_ = new_n735_ & new_n1771_;
  assign new_n1773_ = new_n183_ & new_n201_;
  assign new_n1774_ = ~new_n1772_ & ~new_n1773_;
  assign new_n1775_ = v14 & ~new_n1774_;
  assign new_n1776_ = v13 & new_n1775_;
  assign new_n1777_ = ~v19 & ~v39;
  assign new_n1778_ = ~v17 & new_n1777_;
  assign new_n1779_ = v15 & new_n1778_;
  assign new_n1780_ = v19 & v37;
  assign new_n1781_ = new_n226_ & new_n1780_;
  assign new_n1782_ = ~new_n1779_ & ~new_n1781_;
  assign new_n1783_ = ~v38 & ~new_n1782_;
  assign new_n1784_ = ~v16 & new_n1783_;
  assign new_n1785_ = new_n116_ & new_n735_;
  assign new_n1786_ = ~new_n1784_ & ~new_n1785_;
  assign new_n1787_ = ~v14 & ~new_n1786_;
  assign new_n1788_ = ~v13 & new_n1787_;
  assign new_n1789_ = ~new_n1776_ & ~new_n1788_;
  assign new_n1790_ = ~v18 & ~new_n1789_;
  assign new_n1791_ = ~new_n201_ & ~new_n1771_;
  assign new_n1792_ = v19 & ~new_n1791_;
  assign new_n1793_ = v18 & new_n1792_;
  assign new_n1794_ = ~v17 & new_n1793_;
  assign new_n1795_ = v14 & new_n1794_;
  assign new_n1796_ = ~v14 & new_n1771_;
  assign new_n1797_ = ~new_n1795_ & ~new_n1796_;
  assign new_n1798_ = v13 & ~new_n1797_;
  assign new_n1799_ = ~new_n1790_ & ~new_n1798_;
  assign new_n1800_ = v12 & ~new_n1799_;
  assign new_n1801_ = ~new_n1770_ & ~new_n1800_;
  assign new_n1802_ = v40 & ~new_n1801_;
  assign new_n1803_ = ~v11 & new_n1802_;
  assign new_n1804_ = ~v10 & new_n1803_;
  assign new_n1805_ = ~v8 & new_n1804_;
  assign new_n1806_ = ~v8 & ~new_n1805_;
  assign new_n1807_ = ~v5 & ~new_n1806_;
  assign new_n1808_ = v14 & ~new_n1331_;
  assign new_n1809_ = ~v12 & new_n1808_;
  assign new_n1810_ = v12 & ~v14;
  assign new_n1811_ = new_n1771_ & new_n1810_;
  assign new_n1812_ = ~new_n1809_ & ~new_n1811_;
  assign new_n1813_ = ~v12 & v14;
  assign new_n1814_ = new_n1186_ & new_n1813_;
  assign new_n1815_ = new_n1812_ & ~new_n1814_;
  assign new_n1816_ = ~v13 & ~new_n1815_;
  assign new_n1817_ = v17 & ~new_n1331_;
  assign new_n1818_ = v14 & new_n1817_;
  assign new_n1819_ = v13 & new_n1818_;
  assign new_n1820_ = v12 & new_n1819_;
  assign new_n1821_ = ~new_n1816_ & ~new_n1820_;
  assign new_n1822_ = v12 & new_n1338_;
  assign new_n1823_ = new_n116_ & new_n753_;
  assign new_n1824_ = new_n1822_ & new_n1823_;
  assign new_n1825_ = new_n1821_ & ~new_n1824_;
  assign new_n1826_ = v19 & ~new_n1361_;
  assign new_n1827_ = v12 & new_n1826_;
  assign new_n1828_ = new_n1825_ & ~new_n1827_;
  assign new_n1829_ = v40 & ~new_n1828_;
  assign new_n1830_ = ~v11 & new_n1829_;
  assign new_n1831_ = ~v10 & new_n1830_;
  assign new_n1832_ = ~v8 & new_n1831_;
  assign new_n1833_ = v5 & new_n1832_;
  assign new_n1834_ = ~new_n1807_ & ~new_n1833_;
  assign new_n1835_ = ~v3 & ~new_n1834_;
  assign new_n1836_ = ~v5 & new_n1753_;
  assign new_n1837_ = v3 & new_n1836_;
  assign new_n1838_ = ~new_n1835_ & ~new_n1837_;
  assign new_n1839_ = ~v36 & ~new_n1838_;
  assign new_n1840_ = ~v4 & new_n1839_;
  assign new_n1841_ = ~v2 & new_n1840_;
  assign new_n1842_ = ~v1 & new_n1841_;
  assign new_n1843_ = ~v0 & new_n1842_;
  assign new_n1844_ = ~v8 & new_n838_;
  assign new_n1845_ = ~new_n1843_ & ~new_n1844_;
  assign new_n1846_ = ~v9 & ~new_n1845_;
  assign \v41.19  = new_n1764_ | new_n1846_;
  assign new_n1848_ = ~v29 & ~v31;
  assign new_n1849_ = v21 & v29;
  assign new_n1850_ = v20 & new_n1849_;
  assign new_n1851_ = ~new_n1848_ & ~new_n1850_;
  assign new_n1852_ = ~v14 & ~new_n1851_;
  assign new_n1853_ = ~v16 & ~new_n1358_;
  assign new_n1854_ = ~new_n975_ & ~new_n976_;
  assign new_n1855_ = ~v18 & ~new_n1854_;
  assign new_n1856_ = ~v16 & new_n1855_;
  assign new_n1857_ = new_n1853_ & ~new_n1856_;
  assign new_n1858_ = v14 & ~new_n1857_;
  assign new_n1859_ = ~new_n1852_ & ~new_n1858_;
  assign new_n1860_ = ~v15 & ~new_n1859_;
  assign new_n1861_ = ~v17 & ~new_n1767_;
  assign new_n1862_ = v15 & ~new_n1861_;
  assign new_n1863_ = v14 & new_n1862_;
  assign new_n1864_ = ~new_n1860_ & ~new_n1863_;
  assign new_n1865_ = v13 & ~new_n1864_;
  assign new_n1866_ = ~new_n120_ & ~new_n171_;
  assign new_n1867_ = ~v16 & ~new_n209_;
  assign new_n1868_ = v15 & ~new_n1867_;
  assign new_n1869_ = ~new_n1186_ & ~new_n1868_;
  assign new_n1870_ = ~new_n1866_ & ~new_n1869_;
  assign new_n1871_ = v15 & new_n155_;
  assign new_n1872_ = new_n118_ & ~new_n1871_;
  assign new_n1873_ = v18 & ~new_n1872_;
  assign new_n1874_ = ~v15 & new_n401_;
  assign new_n1875_ = ~new_n180_ & ~new_n1874_;
  assign new_n1876_ = ~v18 & ~new_n1875_;
  assign new_n1877_ = ~new_n1873_ & ~new_n1876_;
  assign new_n1878_ = ~v17 & ~new_n1877_;
  assign new_n1879_ = v15 & ~new_n1106_;
  assign new_n1880_ = ~new_n120_ & ~new_n860_;
  assign new_n1881_ = ~v15 & ~new_n1880_;
  assign new_n1882_ = ~new_n1879_ & ~new_n1881_;
  assign new_n1883_ = v17 & ~new_n1882_;
  assign new_n1884_ = v16 & new_n1883_;
  assign new_n1885_ = ~new_n1878_ & ~new_n1884_;
  assign new_n1886_ = ~new_n1870_ & new_n1885_;
  assign new_n1887_ = ~v14 & ~new_n1886_;
  assign new_n1888_ = ~new_n900_ & ~new_n1887_;
  assign new_n1889_ = ~v13 & ~new_n1888_;
  assign new_n1890_ = ~new_n1865_ & ~new_n1889_;
  assign new_n1891_ = v12 & ~new_n1890_;
  assign new_n1892_ = ~v13 & new_n1808_;
  assign new_n1893_ = new_n116_ & new_n1444_;
  assign new_n1894_ = ~new_n1892_ & ~new_n1893_;
  assign new_n1895_ = ~new_n1866_ & ~new_n1894_;
  assign new_n1896_ = ~new_n1106_ & ~new_n1331_;
  assign new_n1897_ = new_n120_ & new_n201_;
  assign new_n1898_ = ~new_n1896_ & ~new_n1897_;
  assign new_n1899_ = v14 & ~new_n1898_;
  assign new_n1900_ = ~v13 & new_n1899_;
  assign new_n1901_ = ~new_n1895_ & ~new_n1900_;
  assign new_n1902_ = ~v13 & v14;
  assign new_n1903_ = new_n226_ & new_n1902_;
  assign new_n1904_ = new_n246_ & new_n1444_;
  assign new_n1905_ = ~new_n1903_ & ~new_n1904_;
  assign new_n1906_ = ~v18 & ~new_n1905_;
  assign new_n1907_ = new_n120_ & new_n1145_;
  assign new_n1908_ = v15 & ~new_n1907_;
  assign new_n1909_ = ~v14 & ~new_n1908_;
  assign new_n1910_ = v13 & new_n1909_;
  assign new_n1911_ = v17 & new_n1038_;
  assign new_n1912_ = new_n1766_ & new_n1911_;
  assign new_n1913_ = ~new_n1910_ & ~new_n1912_;
  assign new_n1914_ = ~new_n1906_ & new_n1913_;
  assign new_n1915_ = ~v16 & ~new_n1914_;
  assign new_n1916_ = ~v15 & new_n975_;
  assign new_n1917_ = ~new_n246_ & ~new_n1916_;
  assign new_n1918_ = ~v18 & ~new_n1917_;
  assign new_n1919_ = v16 & new_n1918_;
  assign new_n1920_ = ~v14 & new_n1919_;
  assign new_n1921_ = ~v14 & ~new_n1920_;
  assign new_n1922_ = v13 & ~new_n1921_;
  assign new_n1923_ = ~new_n1915_ & ~new_n1922_;
  assign new_n1924_ = new_n1901_ & new_n1923_;
  assign new_n1925_ = ~v12 & ~new_n1924_;
  assign new_n1926_ = ~new_n1891_ & ~new_n1925_;
  assign new_n1927_ = v40 & ~new_n1926_;
  assign new_n1928_ = ~v3 & new_n1927_;
  assign new_n1929_ = v22 & new_n721_;
  assign new_n1930_ = ~new_n726_ & ~new_n1929_;
  assign new_n1931_ = v21 & ~new_n1930_;
  assign new_n1932_ = ~v20 & new_n1931_;
  assign new_n1933_ = ~v19 & new_n1932_;
  assign new_n1934_ = v18 & new_n1933_;
  assign new_n1935_ = v17 & new_n1934_;
  assign new_n1936_ = ~v16 & new_n1935_;
  assign new_n1937_ = ~v15 & new_n1936_;
  assign new_n1938_ = ~v13 & new_n1937_;
  assign new_n1939_ = v12 & new_n1938_;
  assign new_n1940_ = ~new_n792_ & ~new_n1939_;
  assign new_n1941_ = ~v14 & ~new_n1940_;
  assign new_n1942_ = v3 & new_n1941_;
  assign new_n1943_ = ~new_n1928_ & ~new_n1942_;
  assign new_n1944_ = ~v5 & ~new_n1943_;
  assign new_n1945_ = ~v22 & ~new_n1223_;
  assign new_n1946_ = ~new_n1544_ & ~new_n1945_;
  assign new_n1947_ = v21 & ~new_n1946_;
  assign new_n1948_ = ~v20 & new_n1947_;
  assign new_n1949_ = ~new_n1239_ & ~new_n1948_;
  assign new_n1950_ = ~v19 & ~new_n1949_;
  assign new_n1951_ = v18 & new_n1950_;
  assign new_n1952_ = v17 & new_n1951_;
  assign new_n1953_ = ~v15 & new_n1952_;
  assign new_n1954_ = ~v13 & new_n1953_;
  assign new_n1955_ = v12 & new_n1954_;
  assign new_n1956_ = ~new_n773_ & ~new_n1955_;
  assign new_n1957_ = ~v16 & ~new_n1956_;
  assign new_n1958_ = ~new_n786_ & ~new_n1957_;
  assign new_n1959_ = v3 & ~new_n1958_;
  assign new_n1960_ = ~v15 & new_n183_;
  assign new_n1961_ = ~new_n246_ & ~new_n1960_;
  assign new_n1962_ = ~v18 & ~new_n1961_;
  assign new_n1963_ = ~new_n227_ & ~new_n1962_;
  assign new_n1964_ = v16 & ~new_n1963_;
  assign new_n1965_ = v15 & new_n1767_;
  assign new_n1966_ = ~new_n1964_ & ~new_n1965_;
  assign new_n1967_ = v13 & ~new_n1966_;
  assign new_n1968_ = ~v12 & new_n1967_;
  assign new_n1969_ = ~v3 & new_n1968_;
  assign new_n1970_ = ~new_n1959_ & ~new_n1969_;
  assign new_n1971_ = ~v14 & ~new_n1970_;
  assign new_n1972_ = v5 & new_n1971_;
  assign new_n1973_ = ~new_n1944_ & ~new_n1972_;
  assign new_n1974_ = ~v4 & ~new_n1973_;
  assign new_n1975_ = ~v5 & ~new_n1209_;
  assign new_n1976_ = ~v22 & ~v24;
  assign new_n1977_ = v5 & new_n1976_;
  assign new_n1978_ = ~new_n1975_ & ~new_n1977_;
  assign new_n1979_ = v27 & ~new_n1978_;
  assign new_n1980_ = v21 & new_n1979_;
  assign new_n1981_ = ~v20 & new_n1980_;
  assign new_n1982_ = ~v19 & new_n1981_;
  assign new_n1983_ = v18 & new_n1982_;
  assign new_n1984_ = v17 & new_n1983_;
  assign new_n1985_ = ~v15 & new_n1984_;
  assign new_n1986_ = ~v13 & new_n1985_;
  assign new_n1987_ = v12 & new_n1986_;
  assign new_n1988_ = ~new_n773_ & ~new_n1987_;
  assign new_n1989_ = ~v16 & ~new_n1988_;
  assign new_n1990_ = ~new_n786_ & ~new_n1989_;
  assign new_n1991_ = v3 & ~new_n1990_;
  assign new_n1992_ = ~v3 & new_n792_;
  assign new_n1993_ = ~new_n1991_ & ~new_n1992_;
  assign new_n1994_ = ~v14 & ~new_n1993_;
  assign new_n1995_ = v4 & new_n1994_;
  assign new_n1996_ = ~new_n1974_ & ~new_n1995_;
  assign new_n1997_ = ~v2 & ~new_n1996_;
  assign new_n1998_ = ~v4 & v12;
  assign new_n1999_ = ~v3 & new_n1998_;
  assign new_n2000_ = ~v13 & new_n201_;
  assign new_n2001_ = new_n1999_ & new_n2000_;
  assign new_n2002_ = v20 & new_n1638_;
  assign new_n2003_ = new_n1911_ & new_n2002_;
  assign new_n2004_ = new_n2001_ & new_n2003_;
  assign new_n2005_ = ~new_n792_ & ~new_n2004_;
  assign new_n2006_ = new_n201_ & new_n265_;
  assign new_n2007_ = new_n381_ & new_n2006_;
  assign new_n2008_ = ~v19 & ~v20;
  assign new_n2009_ = new_n517_ & new_n2008_;
  assign new_n2010_ = v21 & ~v22;
  assign new_n2011_ = new_n1541_ & new_n2010_;
  assign new_n2012_ = new_n2009_ & new_n2011_;
  assign new_n2013_ = new_n2007_ & new_n2012_;
  assign new_n2014_ = new_n2005_ & ~new_n2013_;
  assign new_n2015_ = ~v14 & ~new_n2014_;
  assign new_n2016_ = v2 & new_n2015_;
  assign new_n2017_ = ~new_n1997_ & ~new_n2016_;
  assign new_n2018_ = ~v1 & ~new_n2017_;
  assign new_n2019_ = ~v18 & ~new_n402_;
  assign new_n2020_ = ~v17 & new_n2019_;
  assign new_n2021_ = v15 & new_n2020_;
  assign new_n2022_ = ~v4 & new_n2021_;
  assign new_n2023_ = ~v3 & new_n2022_;
  assign new_n2024_ = ~v2 & new_n2023_;
  assign new_n2025_ = new_n160_ & ~new_n2024_;
  assign new_n2026_ = new_n161_ & new_n249_;
  assign new_n2027_ = new_n1259_ & new_n1771_;
  assign new_n2028_ = new_n2026_ & new_n2027_;
  assign new_n2029_ = new_n2025_ & ~new_n2028_;
  assign new_n2030_ = ~v14 & ~new_n2029_;
  assign new_n2031_ = v13 & new_n2030_;
  assign new_n2032_ = ~v12 & new_n2031_;
  assign new_n2033_ = v1 & new_n2032_;
  assign new_n2034_ = ~new_n2018_ & ~new_n2033_;
  assign new_n2035_ = ~v0 & ~new_n2034_;
  assign new_n2036_ = v3 & ~new_n252_;
  assign new_n2037_ = ~new_n248_ & ~new_n2036_;
  assign new_n2038_ = new_n165_ & new_n246_;
  assign new_n2039_ = new_n381_ & new_n2038_;
  assign new_n2040_ = ~new_n2037_ & ~new_n2039_;
  assign new_n2041_ = v16 & ~new_n2040_;
  assign new_n2042_ = ~v5 & new_n1965_;
  assign new_n2043_ = ~v4 & new_n2042_;
  assign new_n2044_ = ~v3 & new_n2043_;
  assign new_n2045_ = ~new_n2041_ & ~new_n2044_;
  assign new_n2046_ = ~v14 & ~new_n2045_;
  assign new_n2047_ = v13 & new_n2046_;
  assign new_n2048_ = ~v12 & new_n2047_;
  assign new_n2049_ = ~v2 & new_n2048_;
  assign new_n2050_ = ~v1 & new_n2049_;
  assign new_n2051_ = v0 & new_n2050_;
  assign new_n2052_ = ~new_n2035_ & ~new_n2051_;
  assign new_n2053_ = ~v36 & ~new_n2052_;
  assign new_n2054_ = ~v11 & new_n2053_;
  assign new_n2055_ = ~v10 & new_n2054_;
  assign new_n2056_ = ~v9 & new_n2055_;
  assign \v41.20  = ~v8 & new_n2056_;
  assign new_n2058_ = new_n265_ & new_n753_;
  assign new_n2059_ = new_n754_ & new_n849_;
  assign new_n2060_ = ~new_n2058_ & ~new_n2059_;
  assign new_n2061_ = new_n849_ & new_n1911_;
  assign new_n2062_ = new_n2060_ & ~new_n2061_;
  assign new_n2063_ = v40 & ~new_n2062_;
  assign new_n2064_ = ~v36 & new_n2063_;
  assign new_n2065_ = ~v16 & new_n2064_;
  assign new_n2066_ = v15 & new_n2065_;
  assign new_n2067_ = ~v14 & new_n2066_;
  assign new_n2068_ = ~v11 & new_n2067_;
  assign new_n2069_ = ~v10 & new_n2068_;
  assign new_n2070_ = ~v9 & new_n2069_;
  assign new_n2071_ = ~v8 & new_n2070_;
  assign new_n2072_ = ~v5 & new_n2071_;
  assign new_n2073_ = ~v4 & new_n2072_;
  assign new_n2074_ = ~v3 & new_n2073_;
  assign new_n2075_ = ~v2 & new_n2074_;
  assign new_n2076_ = ~v1 & new_n2075_;
  assign \v41.21  = ~v0 & new_n2076_;
  assign new_n2078_ = ~v19 & ~new_n1517_;
  assign new_n2079_ = v17 & new_n2078_;
  assign new_n2080_ = ~v15 & new_n2079_;
  assign new_n2081_ = v15 & new_n735_;
  assign new_n2082_ = ~new_n2080_ & ~new_n2081_;
  assign new_n2083_ = ~new_n672_ & ~new_n2082_;
  assign new_n2084_ = ~v15 & ~new_n1146_;
  assign new_n2085_ = ~v19 & ~new_n2084_;
  assign new_n2086_ = ~v15 & new_n735_;
  assign new_n2087_ = ~new_n2085_ & ~new_n2086_;
  assign new_n2088_ = ~v5 & ~new_n2087_;
  assign new_n2089_ = new_n607_ & new_n975_;
  assign new_n2090_ = ~new_n2088_ & ~new_n2089_;
  assign new_n2091_ = v40 & ~new_n2090_;
  assign new_n2092_ = ~new_n2083_ & ~new_n2091_;
  assign new_n2093_ = v18 & ~new_n2092_;
  assign new_n2094_ = v15 & new_n976_;
  assign new_n2095_ = ~new_n1916_ & ~new_n2094_;
  assign new_n2096_ = ~new_n843_ & ~new_n2095_;
  assign new_n2097_ = v37 & v39;
  assign new_n2098_ = v17 & ~new_n2097_;
  assign new_n2099_ = v17 & ~new_n2098_;
  assign new_n2100_ = ~v15 & ~new_n2099_;
  assign new_n2101_ = ~new_n1145_ & ~new_n2100_;
  assign new_n2102_ = v19 & ~new_n2101_;
  assign new_n2103_ = ~new_n2096_ & ~new_n2102_;
  assign new_n2104_ = ~new_n1783_ & new_n2103_;
  assign new_n2105_ = v40 & ~new_n2104_;
  assign new_n2106_ = ~v5 & new_n2105_;
  assign new_n2107_ = new_n183_ & new_n653_;
  assign new_n2108_ = ~new_n2106_ & ~new_n2107_;
  assign new_n2109_ = ~v18 & ~new_n2108_;
  assign new_n2110_ = ~new_n2093_ & ~new_n2109_;
  assign new_n2111_ = v12 & ~new_n2110_;
  assign new_n2112_ = ~v12 & v40;
  assign new_n2113_ = ~v5 & new_n2112_;
  assign new_n2114_ = ~new_n2111_ & ~new_n2113_;
  assign new_n2115_ = ~v16 & ~new_n2114_;
  assign new_n2116_ = ~v5 & ~v12;
  assign new_n2117_ = v12 & v15;
  assign new_n2118_ = v5 & new_n2117_;
  assign new_n2119_ = ~new_n2116_ & ~new_n2118_;
  assign new_n2120_ = ~v15 & new_n119_;
  assign new_n2121_ = new_n1634_ & new_n2120_;
  assign new_n2122_ = new_n2119_ & ~new_n2121_;
  assign new_n2123_ = ~v19 & ~new_n843_;
  assign new_n2124_ = ~v19 & ~new_n2123_;
  assign new_n2125_ = ~v18 & ~new_n2124_;
  assign new_n2126_ = ~new_n1038_ & ~new_n2125_;
  assign new_n2127_ = v17 & ~new_n2126_;
  assign new_n2128_ = ~v15 & new_n2127_;
  assign new_n2129_ = v12 & new_n2128_;
  assign new_n2130_ = ~v5 & new_n2129_;
  assign new_n2131_ = new_n2122_ & ~new_n2130_;
  assign new_n2132_ = v40 & ~new_n2131_;
  assign new_n2133_ = v16 & new_n2132_;
  assign new_n2134_ = ~new_n2115_ & ~new_n2133_;
  assign new_n2135_ = ~v14 & ~new_n2134_;
  assign new_n2136_ = v5 & ~new_n1332_;
  assign new_n2137_ = new_n207_ & new_n1767_;
  assign new_n2138_ = ~new_n2136_ & ~new_n2137_;
  assign new_n2139_ = ~v5 & new_n201_;
  assign new_n2140_ = new_n1039_ & new_n2139_;
  assign new_n2141_ = new_n2138_ & ~new_n2140_;
  assign new_n2142_ = ~v12 & ~new_n2141_;
  assign new_n2143_ = ~v5 & new_n2117_;
  assign new_n2144_ = ~new_n2142_ & ~new_n2143_;
  assign new_n2145_ = v40 & ~new_n2144_;
  assign new_n2146_ = v14 & new_n2145_;
  assign new_n2147_ = ~new_n2135_ & ~new_n2146_;
  assign new_n2148_ = ~v13 & ~new_n2147_;
  assign new_n2149_ = v12 & ~v29;
  assign new_n2150_ = ~v17 & ~new_n1106_;
  assign new_n2151_ = ~new_n1911_ & ~new_n2150_;
  assign new_n2152_ = v16 & ~new_n2151_;
  assign new_n2153_ = ~v12 & new_n2152_;
  assign new_n2154_ = ~new_n2149_ & ~new_n2153_;
  assign new_n2155_ = ~v15 & ~new_n2154_;
  assign new_n2156_ = v16 & ~new_n1469_;
  assign new_n2157_ = ~new_n883_ & ~new_n2156_;
  assign new_n2158_ = ~v12 & ~new_n2157_;
  assign new_n2159_ = ~v12 & ~new_n2158_;
  assign new_n2160_ = v15 & ~new_n2159_;
  assign new_n2161_ = ~new_n2155_ & ~new_n2160_;
  assign new_n2162_ = ~v14 & ~new_n2161_;
  assign new_n2163_ = ~v15 & new_n489_;
  assign new_n2164_ = ~v15 & ~new_n2163_;
  assign new_n2165_ = new_n165_ & new_n201_;
  assign new_n2166_ = new_n2164_ & ~new_n2165_;
  assign new_n2167_ = ~v17 & ~new_n2166_;
  assign new_n2168_ = ~new_n268_ & ~new_n2167_;
  assign new_n2169_ = v12 & ~new_n2168_;
  assign new_n2170_ = ~v12 & v15;
  assign new_n2171_ = ~new_n2169_ & ~new_n2170_;
  assign new_n2172_ = v14 & ~new_n2171_;
  assign new_n2173_ = ~new_n2162_ & ~new_n2172_;
  assign new_n2174_ = ~v5 & ~new_n2173_;
  assign new_n2175_ = ~new_n1817_ & ~new_n1823_;
  assign new_n2176_ = new_n116_ & new_n1259_;
  assign new_n2177_ = new_n2175_ & ~new_n2176_;
  assign new_n2178_ = v14 & ~new_n2177_;
  assign new_n2179_ = v12 & new_n2178_;
  assign new_n2180_ = v5 & new_n2179_;
  assign new_n2181_ = ~new_n2174_ & ~new_n2180_;
  assign new_n2182_ = v40 & ~new_n2181_;
  assign new_n2183_ = ~v12 & new_n1748_;
  assign new_n2184_ = v5 & new_n2183_;
  assign new_n2185_ = ~new_n2182_ & ~new_n2184_;
  assign new_n2186_ = v13 & ~new_n2185_;
  assign new_n2187_ = ~v5 & ~v40;
  assign new_n2188_ = ~new_n2186_ & ~new_n2187_;
  assign new_n2189_ = ~new_n2148_ & new_n2188_;
  assign new_n2190_ = ~v4 & ~new_n2189_;
  assign new_n2191_ = new_n265_ & new_n735_;
  assign new_n2192_ = new_n183_ & new_n849_;
  assign new_n2193_ = ~new_n2191_ & ~new_n2192_;
  assign new_n2194_ = v18 & ~new_n2193_;
  assign new_n2195_ = v13 & new_n754_;
  assign new_n2196_ = ~v12 & new_n2195_;
  assign new_n2197_ = ~new_n2194_ & ~new_n2196_;
  assign new_n2198_ = v15 & ~new_n2197_;
  assign new_n2199_ = ~v19 & ~new_n1529_;
  assign new_n2200_ = v17 & new_n2199_;
  assign new_n2201_ = ~v15 & new_n2200_;
  assign new_n2202_ = ~v13 & new_n2201_;
  assign new_n2203_ = v12 & new_n2202_;
  assign new_n2204_ = ~new_n2198_ & ~new_n2203_;
  assign new_n2205_ = ~v16 & ~new_n2204_;
  assign new_n2206_ = ~v14 & new_n2205_;
  assign new_n2207_ = v4 & new_n2206_;
  assign new_n2208_ = ~new_n2190_ & ~new_n2207_;
  assign new_n2209_ = ~v3 & ~new_n2208_;
  assign new_n2210_ = ~v12 & new_n1694_;
  assign new_n2211_ = ~new_n680_ & ~new_n1976_;
  assign new_n2212_ = v21 & ~new_n2211_;
  assign new_n2213_ = ~v20 & new_n2212_;
  assign new_n2214_ = ~new_n679_ & ~new_n2213_;
  assign new_n2215_ = v22 & new_n688_;
  assign new_n2216_ = ~new_n692_ & ~new_n2215_;
  assign new_n2217_ = v27 & ~new_n2216_;
  assign new_n2218_ = v21 & new_n2217_;
  assign new_n2219_ = ~v20 & new_n2218_;
  assign new_n2220_ = new_n2214_ & ~new_n2219_;
  assign new_n2221_ = v18 & ~new_n2220_;
  assign new_n2222_ = v18 & ~new_n2221_;
  assign new_n2223_ = ~v15 & ~new_n2222_;
  assign new_n2224_ = ~v13 & new_n2223_;
  assign new_n2225_ = v12 & new_n2224_;
  assign new_n2226_ = ~new_n2210_ & ~new_n2225_;
  assign new_n2227_ = ~v5 & ~new_n2226_;
  assign new_n2228_ = ~v23 & ~new_n1539_;
  assign new_n2229_ = v22 & new_n2228_;
  assign new_n2230_ = ~v22 & new_n1541_;
  assign new_n2231_ = ~new_n2229_ & ~new_n2230_;
  assign new_n2232_ = v21 & ~new_n2231_;
  assign new_n2233_ = ~v20 & new_n2232_;
  assign new_n2234_ = ~new_n2002_ & ~new_n2233_;
  assign new_n2235_ = v18 & ~new_n2234_;
  assign new_n2236_ = ~v15 & new_n2235_;
  assign new_n2237_ = ~v13 & new_n2236_;
  assign new_n2238_ = v12 & new_n2237_;
  assign new_n2239_ = v5 & new_n2238_;
  assign new_n2240_ = ~new_n2227_ & ~new_n2239_;
  assign new_n2241_ = ~v4 & ~new_n2240_;
  assign new_n2242_ = ~v20 & v21;
  assign new_n2243_ = ~v23 & ~v24;
  assign new_n2244_ = v22 & new_n2243_;
  assign new_n2245_ = new_n2242_ & new_n2244_;
  assign new_n2246_ = ~new_n679_ & ~new_n2245_;
  assign new_n2247_ = ~v5 & ~v20;
  assign new_n2248_ = v21 & new_n1976_;
  assign new_n2249_ = new_n2247_ & new_n2248_;
  assign new_n2250_ = new_n2246_ & ~new_n2249_;
  assign new_n2251_ = v27 & ~new_n2250_;
  assign new_n2252_ = v18 & new_n2251_;
  assign new_n2253_ = ~v15 & new_n2252_;
  assign new_n2254_ = ~v13 & new_n2253_;
  assign new_n2255_ = v12 & new_n2254_;
  assign new_n2256_ = v4 & new_n2255_;
  assign new_n2257_ = ~new_n2241_ & ~new_n2256_;
  assign new_n2258_ = ~v19 & ~new_n2257_;
  assign new_n2259_ = ~v4 & new_n2116_;
  assign new_n2260_ = new_n165_ & new_n1694_;
  assign new_n2261_ = new_n2259_ & new_n2260_;
  assign new_n2262_ = ~new_n2258_ & ~new_n2261_;
  assign new_n2263_ = v17 & ~new_n2262_;
  assign new_n2264_ = ~v16 & new_n2263_;
  assign new_n2265_ = ~v14 & new_n2264_;
  assign new_n2266_ = v3 & new_n2265_;
  assign new_n2267_ = ~new_n2209_ & ~new_n2266_;
  assign new_n2268_ = ~v2 & ~new_n2267_;
  assign new_n2269_ = v2 & ~v3;
  assign new_n2270_ = new_n169_ & new_n2269_;
  assign new_n2271_ = new_n265_ & new_n1012_;
  assign new_n2272_ = new_n2270_ & new_n2271_;
  assign new_n2273_ = v21 & v22;
  assign new_n2274_ = ~v23 & new_n1541_;
  assign new_n2275_ = new_n2273_ & new_n2274_;
  assign new_n2276_ = new_n2009_ & new_n2275_;
  assign new_n2277_ = new_n2272_ & new_n2276_;
  assign new_n2278_ = ~new_n2268_ & ~new_n2277_;
  assign new_n2279_ = ~v0 & ~new_n2278_;
  assign new_n2280_ = v0 & new_n161_;
  assign new_n2281_ = ~v4 & new_n1634_;
  assign new_n2282_ = new_n2280_ & new_n2281_;
  assign new_n2283_ = ~v13 & new_n383_;
  assign new_n2284_ = new_n210_ & new_n2283_;
  assign new_n2285_ = new_n2282_ & new_n2284_;
  assign new_n2286_ = ~new_n2279_ & ~new_n2285_;
  assign new_n2287_ = ~v36 & ~new_n2286_;
  assign new_n2288_ = ~v1 & new_n2287_;
  assign new_n2289_ = ~v36 & ~new_n2288_;
  assign new_n2290_ = ~v10 & ~new_n2289_;
  assign new_n2291_ = ~v10 & ~new_n2290_;
  assign new_n2292_ = ~v9 & ~new_n2291_;
  assign new_n2293_ = ~v9 & ~new_n2292_;
  assign new_n2294_ = ~v11 & ~new_n2293_;
  assign new_n2295_ = ~v9 & v10;
  assign new_n2296_ = ~v9 & ~new_n2295_;
  assign new_n2297_ = v11 & ~new_n2296_;
  assign new_n2298_ = ~new_n2294_ & ~new_n2297_;
  assign new_n2299_ = ~v8 & ~new_n2298_;
  assign new_n2300_ = ~v9 & ~v36;
  assign new_n2301_ = v8 & new_n2300_;
  assign new_n2302_ = ~v5 & new_n2301_;
  assign new_n2303_ = ~v4 & new_n2302_;
  assign new_n2304_ = ~v3 & new_n2303_;
  assign new_n2305_ = ~v2 & new_n2304_;
  assign new_n2306_ = ~v1 & new_n2305_;
  assign new_n2307_ = ~v0 & new_n2306_;
  assign \v41.22  = new_n2299_ | new_n2307_;
  assign new_n2309_ = v20 & ~new_n679_;
  assign new_n2310_ = v29 & ~new_n2309_;
  assign new_n2311_ = v29 & ~new_n2310_;
  assign new_n2312_ = ~v15 & ~new_n2311_;
  assign new_n2313_ = ~v14 & new_n2312_;
  assign new_n2314_ = v13 & new_n2313_;
  assign new_n2315_ = ~v14 & v18;
  assign new_n2316_ = ~v13 & new_n2315_;
  assign new_n2317_ = v14 & ~v18;
  assign new_n2318_ = v13 & new_n2317_;
  assign new_n2319_ = ~new_n2316_ & ~new_n2318_;
  assign new_n2320_ = ~v17 & ~new_n2319_;
  assign new_n2321_ = ~v16 & new_n2320_;
  assign new_n2322_ = v15 & new_n2321_;
  assign new_n2323_ = ~new_n2314_ & ~new_n2322_;
  assign new_n2324_ = v12 & ~new_n2323_;
  assign new_n2325_ = v14 & v15;
  assign new_n2326_ = new_n849_ & new_n2325_;
  assign new_n2327_ = ~new_n2324_ & ~new_n2326_;
  assign new_n2328_ = v40 & ~new_n2327_;
  assign new_n2329_ = ~v36 & new_n2328_;
  assign new_n2330_ = ~v11 & new_n2329_;
  assign new_n2331_ = ~v10 & new_n2330_;
  assign new_n2332_ = ~v9 & new_n2331_;
  assign new_n2333_ = ~v8 & new_n2332_;
  assign new_n2334_ = ~v5 & new_n2333_;
  assign new_n2335_ = ~v4 & new_n2334_;
  assign new_n2336_ = ~v3 & new_n2335_;
  assign new_n2337_ = ~v2 & new_n2336_;
  assign new_n2338_ = ~v1 & new_n2337_;
  assign \v41.23  = ~v0 & new_n2338_;
  assign new_n2340_ = ~v8 & v9;
  assign new_n2341_ = ~v0 & ~v1;
  assign new_n2342_ = new_n161_ & new_n2341_;
  assign new_n2343_ = new_n169_ & new_n2301_;
  assign new_n2344_ = new_n2342_ & new_n2343_;
  assign new_n2345_ = ~new_n2340_ & ~new_n2344_;
  assign new_n2346_ = ~v8 & new_n2295_;
  assign new_n2347_ = new_n2345_ & ~new_n2346_;
  assign new_n2348_ = ~new_n390_ & ~new_n1483_;
  assign new_n2349_ = ~v15 & new_n1049_;
  assign new_n2350_ = ~v13 & new_n2349_;
  assign new_n2351_ = v12 & new_n2350_;
  assign new_n2352_ = ~new_n773_ & ~new_n2351_;
  assign new_n2353_ = ~v16 & ~new_n2352_;
  assign new_n2354_ = ~new_n786_ & ~new_n2353_;
  assign new_n2355_ = ~v2 & ~new_n2354_;
  assign new_n2356_ = ~new_n796_ & ~new_n2355_;
  assign new_n2357_ = ~v1 & ~new_n2356_;
  assign new_n2358_ = v13 & ~new_n160_;
  assign new_n2359_ = ~v12 & new_n2358_;
  assign new_n2360_ = v1 & new_n2359_;
  assign new_n2361_ = ~new_n2357_ & ~new_n2360_;
  assign new_n2362_ = ~new_n2348_ & ~new_n2361_;
  assign new_n2363_ = v3 & v4;
  assign new_n2364_ = ~v2 & new_n2363_;
  assign new_n2365_ = v2 & new_n256_;
  assign new_n2366_ = ~new_n2364_ & ~new_n2365_;
  assign new_n2367_ = ~v1 & new_n2021_;
  assign new_n2368_ = new_n160_ & ~new_n2367_;
  assign new_n2369_ = v13 & ~new_n2368_;
  assign new_n2370_ = ~v12 & new_n2369_;
  assign new_n2371_ = ~v1 & v12;
  assign new_n2372_ = new_n2000_ & new_n2371_;
  assign new_n2373_ = new_n2003_ & new_n2372_;
  assign new_n2374_ = ~new_n2370_ & ~new_n2373_;
  assign new_n2375_ = ~new_n2366_ & ~new_n2374_;
  assign new_n2376_ = ~v3 & v17;
  assign new_n2377_ = ~v2 & new_n2376_;
  assign new_n2378_ = v3 & ~v17;
  assign new_n2379_ = v2 & new_n2378_;
  assign new_n2380_ = ~new_n2377_ & ~new_n2379_;
  assign new_n2381_ = ~v18 & ~new_n2380_;
  assign new_n2382_ = new_n161_ & new_n1911_;
  assign new_n2383_ = ~new_n2381_ & ~new_n2382_;
  assign new_n2384_ = v13 & ~new_n2383_;
  assign new_n2385_ = ~v12 & new_n2384_;
  assign new_n2386_ = ~v13 & ~v17;
  assign new_n2387_ = new_n120_ & new_n2386_;
  assign new_n2388_ = new_n339_ & new_n2387_;
  assign new_n2389_ = ~new_n2385_ & ~new_n2388_;
  assign new_n2390_ = v15 & ~new_n2389_;
  assign new_n2391_ = v3 & new_n1541_;
  assign new_n2392_ = ~v3 & new_n722_;
  assign new_n2393_ = ~new_n2391_ & ~new_n2392_;
  assign new_n2394_ = ~new_n681_ & ~new_n2393_;
  assign new_n2395_ = ~v3 & new_n1929_;
  assign new_n2396_ = ~new_n2394_ & ~new_n2395_;
  assign new_n2397_ = v21 & ~new_n2396_;
  assign new_n2398_ = ~v20 & new_n2397_;
  assign new_n2399_ = v18 & new_n2398_;
  assign new_n2400_ = ~v3 & ~v18;
  assign new_n2401_ = ~new_n2399_ & ~new_n2400_;
  assign new_n2402_ = ~v19 & ~new_n2401_;
  assign new_n2403_ = v17 & new_n2402_;
  assign new_n2404_ = ~v15 & new_n2403_;
  assign new_n2405_ = ~v13 & new_n2404_;
  assign new_n2406_ = v12 & new_n2405_;
  assign new_n2407_ = ~v2 & new_n2406_;
  assign new_n2408_ = ~new_n2390_ & ~new_n2407_;
  assign new_n2409_ = ~v16 & ~new_n2408_;
  assign new_n2410_ = v3 & new_n786_;
  assign new_n2411_ = v2 & new_n2410_;
  assign new_n2412_ = ~new_n2409_ & ~new_n2411_;
  assign new_n2413_ = ~v1 & ~new_n2412_;
  assign new_n2414_ = v3 & new_n2359_;
  assign new_n2415_ = v2 & new_n2414_;
  assign new_n2416_ = v1 & new_n2415_;
  assign new_n2417_ = ~new_n2413_ & ~new_n2416_;
  assign new_n2418_ = v4 & ~new_n2417_;
  assign new_n2419_ = ~v16 & ~new_n154_;
  assign new_n2420_ = ~v18 & ~new_n2419_;
  assign new_n2421_ = ~v17 & new_n2420_;
  assign new_n2422_ = v15 & new_n2421_;
  assign new_n2423_ = ~new_n139_ & ~new_n2422_;
  assign new_n2424_ = v13 & ~new_n2423_;
  assign new_n2425_ = ~v12 & new_n2424_;
  assign new_n2426_ = ~v4 & new_n2425_;
  assign new_n2427_ = ~v3 & new_n2426_;
  assign new_n2428_ = ~v2 & new_n2427_;
  assign new_n2429_ = v1 & new_n2428_;
  assign new_n2430_ = ~new_n2418_ & ~new_n2429_;
  assign new_n2431_ = ~new_n2375_ & new_n2430_;
  assign new_n2432_ = ~new_n2362_ & new_n2431_;
  assign new_n2433_ = ~v0 & ~new_n2432_;
  assign new_n2434_ = v13 & new_n1661_;
  assign new_n2435_ = ~v12 & new_n2434_;
  assign new_n2436_ = ~v3 & new_n2435_;
  assign new_n2437_ = ~v2 & new_n2436_;
  assign new_n2438_ = ~v1 & new_n2437_;
  assign new_n2439_ = v0 & new_n2438_;
  assign new_n2440_ = ~new_n2433_ & ~new_n2439_;
  assign new_n2441_ = ~v2 & ~new_n672_;
  assign new_n2442_ = v2 & ~v5;
  assign new_n2443_ = new_n1541_ & new_n2442_;
  assign new_n2444_ = ~new_n2441_ & ~new_n2443_;
  assign new_n2445_ = ~new_n681_ & ~new_n2444_;
  assign new_n2446_ = v23 & ~new_n672_;
  assign new_n2447_ = v22 & new_n2446_;
  assign new_n2448_ = ~v2 & new_n2447_;
  assign new_n2449_ = ~new_n2445_ & ~new_n2448_;
  assign new_n2450_ = ~v20 & ~new_n2449_;
  assign new_n2451_ = v20 & ~new_n672_;
  assign new_n2452_ = ~v2 & new_n2451_;
  assign new_n2453_ = ~new_n2450_ & ~new_n2452_;
  assign new_n2454_ = v21 & ~new_n2453_;
  assign new_n2455_ = ~v21 & ~new_n672_;
  assign new_n2456_ = v20 & new_n2455_;
  assign new_n2457_ = ~v2 & new_n2456_;
  assign new_n2458_ = ~new_n2454_ & ~new_n2457_;
  assign new_n2459_ = v18 & ~new_n2458_;
  assign new_n2460_ = v5 & ~v18;
  assign new_n2461_ = ~v2 & new_n2460_;
  assign new_n2462_ = ~new_n2459_ & ~new_n2461_;
  assign new_n2463_ = ~v19 & ~new_n2462_;
  assign new_n2464_ = ~v5 & new_n1649_;
  assign new_n2465_ = ~v2 & new_n2464_;
  assign new_n2466_ = ~new_n2463_ & ~new_n2465_;
  assign new_n2467_ = v17 & ~new_n2466_;
  assign new_n2468_ = v40 & ~new_n194_;
  assign new_n2469_ = ~v17 & new_n2468_;
  assign new_n2470_ = ~v5 & new_n2469_;
  assign new_n2471_ = ~v2 & new_n2470_;
  assign new_n2472_ = ~new_n2467_ & ~new_n2471_;
  assign new_n2473_ = ~v15 & ~new_n2472_;
  assign new_n2474_ = v17 & ~new_n1409_;
  assign new_n2475_ = v19 & ~new_n2474_;
  assign new_n2476_ = v5 & new_n2475_;
  assign new_n2477_ = ~v5 & v17;
  assign new_n2478_ = new_n1595_ & new_n2477_;
  assign new_n2479_ = ~new_n2476_ & ~new_n2478_;
  assign new_n2480_ = v18 & ~new_n2479_;
  assign new_n2481_ = v40 & ~new_n1854_;
  assign new_n2482_ = ~v18 & new_n2481_;
  assign new_n2483_ = ~v5 & new_n2482_;
  assign new_n2484_ = ~new_n2480_ & ~new_n2483_;
  assign new_n2485_ = v15 & ~new_n2484_;
  assign new_n2486_ = ~v2 & new_n2485_;
  assign new_n2487_ = ~new_n2473_ & ~new_n2486_;
  assign new_n2488_ = v12 & ~new_n2487_;
  assign new_n2489_ = ~v2 & new_n2113_;
  assign new_n2490_ = ~new_n2488_ & ~new_n2489_;
  assign new_n2491_ = ~v16 & ~new_n2490_;
  assign new_n2492_ = ~v2 & new_n2133_;
  assign new_n2493_ = ~new_n2491_ & ~new_n2492_;
  assign new_n2494_ = ~v13 & ~new_n2493_;
  assign new_n2495_ = ~v15 & ~v18;
  assign new_n2496_ = ~new_n1571_ & ~new_n2495_;
  assign new_n2497_ = v15 & new_n754_;
  assign new_n2498_ = new_n2496_ & ~new_n2497_;
  assign new_n2499_ = v16 & ~new_n2498_;
  assign new_n2500_ = ~v16 & ~new_n1469_;
  assign new_n2501_ = v15 & new_n2500_;
  assign new_n2502_ = ~new_n2499_ & ~new_n2501_;
  assign new_n2503_ = v40 & ~new_n2502_;
  assign new_n2504_ = ~v5 & new_n2503_;
  assign new_n2505_ = new_n607_ & new_n1486_;
  assign new_n2506_ = ~new_n2504_ & ~new_n2505_;
  assign new_n2507_ = v5 & ~new_n518_;
  assign new_n2508_ = ~v5 & ~v17;
  assign new_n2509_ = new_n385_ & new_n2508_;
  assign new_n2510_ = ~new_n2507_ & ~new_n2509_;
  assign new_n2511_ = ~v16 & ~new_n2510_;
  assign new_n2512_ = v15 & new_n2511_;
  assign new_n2513_ = ~new_n1101_ & ~new_n2512_;
  assign new_n2514_ = ~v19 & ~new_n2513_;
  assign new_n2515_ = v19 & ~new_n672_;
  assign new_n2516_ = ~v18 & new_n2515_;
  assign new_n2517_ = ~v17 & new_n2516_;
  assign new_n2518_ = v16 & new_n2517_;
  assign new_n2519_ = v15 & new_n2518_;
  assign new_n2520_ = ~new_n2514_ & ~new_n2519_;
  assign new_n2521_ = new_n2506_ & new_n2520_;
  assign new_n2522_ = ~v12 & ~new_n2521_;
  assign new_n2523_ = ~v15 & new_n1133_;
  assign new_n2524_ = v23 & v29;
  assign new_n2525_ = ~v22 & new_n2524_;
  assign new_n2526_ = new_n2523_ & new_n2525_;
  assign new_n2527_ = ~v15 & ~new_n2526_;
  assign new_n2528_ = v40 & ~new_n2527_;
  assign new_n2529_ = v12 & new_n2528_;
  assign new_n2530_ = ~v5 & new_n2529_;
  assign new_n2531_ = ~new_n2522_ & ~new_n2530_;
  assign new_n2532_ = v13 & ~new_n2531_;
  assign new_n2533_ = ~v2 & new_n2532_;
  assign new_n2534_ = ~new_n2494_ & ~new_n2533_;
  assign new_n2535_ = ~v3 & ~new_n2534_;
  assign new_n2536_ = v18 & new_n2242_;
  assign new_n2537_ = new_n680_ & new_n722_;
  assign new_n2538_ = new_n2536_ & new_n2537_;
  assign new_n2539_ = v18 & ~new_n2538_;
  assign new_n2540_ = ~v15 & ~new_n2539_;
  assign new_n2541_ = ~v13 & new_n2540_;
  assign new_n2542_ = v12 & new_n2541_;
  assign new_n2543_ = ~new_n2210_ & ~new_n2542_;
  assign new_n2544_ = ~v19 & ~new_n2543_;
  assign new_n2545_ = v15 & new_n165_;
  assign new_n2546_ = new_n849_ & new_n2545_;
  assign new_n2547_ = ~new_n2544_ & ~new_n2546_;
  assign new_n2548_ = v17 & ~new_n2547_;
  assign new_n2549_ = ~v16 & new_n2548_;
  assign new_n2550_ = ~v5 & new_n2549_;
  assign new_n2551_ = v3 & new_n2550_;
  assign new_n2552_ = ~v2 & new_n2551_;
  assign new_n2553_ = ~new_n2535_ & ~new_n2552_;
  assign new_n2554_ = ~v0 & ~new_n2553_;
  assign new_n2555_ = ~v3 & new_n1965_;
  assign new_n2556_ = ~new_n1262_ & ~new_n2555_;
  assign new_n2557_ = v13 & ~new_n2556_;
  assign new_n2558_ = ~v12 & new_n2557_;
  assign new_n2559_ = ~new_n1269_ & ~new_n2558_;
  assign new_n2560_ = ~v5 & ~new_n2559_;
  assign new_n2561_ = ~v2 & new_n2560_;
  assign new_n2562_ = v0 & new_n2561_;
  assign new_n2563_ = ~new_n2554_ & ~new_n2562_;
  assign new_n2564_ = ~v1 & ~new_n2563_;
  assign new_n2565_ = ~v0 & new_n1442_;
  assign new_n2566_ = ~v3 & new_n2116_;
  assign new_n2567_ = new_n2565_ & new_n2566_;
  assign new_n2568_ = v13 & new_n117_;
  assign new_n2569_ = new_n172_ & new_n2568_;
  assign new_n2570_ = new_n2567_ & new_n2569_;
  assign new_n2571_ = ~new_n2564_ & ~new_n2570_;
  assign new_n2572_ = ~v4 & ~new_n2571_;
  assign new_n2573_ = new_n2440_ & ~new_n2572_;
  assign new_n2574_ = ~v14 & ~new_n2573_;
  assign new_n2575_ = v12 & new_n1727_;
  assign new_n2576_ = ~new_n1679_ & ~new_n2575_;
  assign new_n2577_ = ~v15 & new_n164_;
  assign new_n2578_ = ~new_n1817_ & ~new_n2577_;
  assign new_n2579_ = v5 & ~new_n2578_;
  assign new_n2580_ = new_n207_ & new_n259_;
  assign new_n2581_ = ~new_n2579_ & ~new_n2580_;
  assign new_n2582_ = ~new_n2576_ & ~new_n2581_;
  assign new_n2583_ = ~v5 & new_n1646_;
  assign new_n2584_ = v5 & new_n1472_;
  assign new_n2585_ = ~new_n2583_ & ~new_n2584_;
  assign new_n2586_ = ~v17 & ~new_n2585_;
  assign new_n2587_ = v15 & new_n2586_;
  assign new_n2588_ = new_n1186_ & new_n2584_;
  assign new_n2589_ = ~new_n2587_ & ~new_n2588_;
  assign new_n2590_ = ~v13 & v18;
  assign new_n2591_ = ~v12 & new_n2590_;
  assign new_n2592_ = v13 & ~v18;
  assign new_n2593_ = v12 & new_n2592_;
  assign new_n2594_ = ~new_n2591_ & ~new_n2593_;
  assign new_n2595_ = ~new_n1331_ & ~new_n2594_;
  assign new_n2596_ = v17 & new_n2595_;
  assign new_n2597_ = ~v12 & new_n766_;
  assign new_n2598_ = new_n1350_ & new_n2597_;
  assign new_n2599_ = ~new_n2596_ & ~new_n2598_;
  assign new_n2600_ = v5 & ~new_n2599_;
  assign new_n2601_ = new_n2589_ & ~new_n2600_;
  assign new_n2602_ = ~new_n2582_ & new_n2601_;
  assign new_n2603_ = ~new_n183_ & ~new_n735_;
  assign new_n2604_ = ~v18 & ~new_n2603_;
  assign new_n2605_ = ~v16 & new_n2604_;
  assign new_n2606_ = ~v15 & new_n2605_;
  assign new_n2607_ = v13 & new_n2606_;
  assign new_n2608_ = ~new_n821_ & ~new_n2607_;
  assign new_n2609_ = v12 & ~new_n2608_;
  assign new_n2610_ = new_n259_ & new_n1038_;
  assign new_n2611_ = new_n2597_ & new_n2610_;
  assign new_n2612_ = ~new_n2609_ & ~new_n2611_;
  assign new_n2613_ = ~v5 & ~new_n2612_;
  assign new_n2614_ = new_n765_ & new_n1689_;
  assign new_n2615_ = new_n166_ & new_n2614_;
  assign new_n2616_ = ~new_n2613_ & ~new_n2615_;
  assign new_n2617_ = new_n2602_ & new_n2616_;
  assign new_n2618_ = v40 & ~new_n2617_;
  assign new_n2619_ = v14 & new_n2618_;
  assign new_n2620_ = ~new_n2187_ & ~new_n2619_;
  assign new_n2621_ = ~v4 & ~new_n2620_;
  assign new_n2622_ = ~v3 & new_n2621_;
  assign new_n2623_ = ~v2 & new_n2622_;
  assign new_n2624_ = ~v1 & new_n2623_;
  assign new_n2625_ = ~v0 & new_n2624_;
  assign new_n2626_ = ~new_n2574_ & ~new_n2625_;
  assign new_n2627_ = ~v36 & ~new_n2626_;
  assign new_n2628_ = ~v36 & ~new_n2627_;
  assign new_n2629_ = ~v11 & ~new_n2628_;
  assign new_n2630_ = ~v10 & new_n2629_;
  assign new_n2631_ = ~v9 & new_n2630_;
  assign new_n2632_ = ~v8 & new_n2631_;
  assign \v41.24  = ~new_n2347_ | new_n2632_;
  assign new_n2634_ = v29 & v40;
  assign new_n2635_ = v13 & new_n2634_;
  assign new_n2636_ = ~v5 & new_n2635_;
  assign new_n2637_ = ~v3 & new_n2636_;
  assign new_n2638_ = ~new_n1231_ & ~new_n2217_;
  assign new_n2639_ = v21 & ~new_n2638_;
  assign new_n2640_ = ~v19 & new_n2639_;
  assign new_n2641_ = v18 & new_n2640_;
  assign new_n2642_ = v17 & new_n2641_;
  assign new_n2643_ = ~v16 & new_n2642_;
  assign new_n2644_ = ~v13 & new_n2643_;
  assign new_n2645_ = v5 & new_n2644_;
  assign new_n2646_ = v3 & new_n2645_;
  assign new_n2647_ = ~new_n2637_ & ~new_n2646_;
  assign new_n2648_ = ~v20 & ~new_n2647_;
  assign new_n2649_ = ~v22 & v23;
  assign new_n2650_ = v21 & new_n2649_;
  assign new_n2651_ = v21 & ~new_n2650_;
  assign new_n2652_ = v40 & ~new_n2651_;
  assign new_n2653_ = v29 & new_n2652_;
  assign new_n2654_ = v13 & new_n2653_;
  assign new_n2655_ = ~v5 & new_n2654_;
  assign new_n2656_ = ~v3 & new_n2655_;
  assign new_n2657_ = v3 & v5;
  assign new_n2658_ = ~v13 & ~v16;
  assign new_n2659_ = new_n2657_ & new_n2658_;
  assign new_n2660_ = ~v19 & new_n1238_;
  assign new_n2661_ = new_n517_ & new_n2660_;
  assign new_n2662_ = new_n2659_ & new_n2661_;
  assign new_n2663_ = ~new_n2656_ & ~new_n2662_;
  assign new_n2664_ = v20 & ~new_n2663_;
  assign new_n2665_ = ~v29 & v40;
  assign new_n2666_ = v13 & new_n2665_;
  assign new_n2667_ = ~v5 & new_n2666_;
  assign new_n2668_ = ~v3 & new_n2667_;
  assign new_n2669_ = ~new_n2664_ & ~new_n2668_;
  assign new_n2670_ = ~new_n2648_ & new_n2669_;
  assign new_n2671_ = v12 & ~new_n2670_;
  assign new_n2672_ = v3 & v18;
  assign new_n2673_ = ~v3 & ~v5;
  assign new_n2674_ = new_n385_ & new_n2673_;
  assign new_n2675_ = ~new_n2672_ & ~new_n2674_;
  assign new_n2676_ = v19 & ~new_n2675_;
  assign new_n2677_ = new_n1596_ & new_n2673_;
  assign new_n2678_ = ~new_n2676_ & ~new_n2677_;
  assign new_n2679_ = v17 & ~new_n2678_;
  assign new_n2680_ = ~v3 & new_n2508_;
  assign new_n2681_ = new_n1596_ & new_n2680_;
  assign new_n2682_ = ~new_n2679_ & ~new_n2681_;
  assign new_n2683_ = v16 & ~new_n2682_;
  assign new_n2684_ = v13 & new_n2683_;
  assign new_n2685_ = ~v12 & new_n2684_;
  assign new_n2686_ = ~new_n2671_ & ~new_n2685_;
  assign new_n2687_ = ~v15 & ~new_n2686_;
  assign new_n2688_ = ~v3 & new_n1595_;
  assign new_n2689_ = ~v3 & ~new_n2688_;
  assign new_n2690_ = ~v18 & ~new_n2689_;
  assign new_n2691_ = ~v17 & new_n2690_;
  assign new_n2692_ = v18 & new_n1648_;
  assign new_n2693_ = new_n2376_ & new_n2692_;
  assign new_n2694_ = ~new_n2691_ & ~new_n2693_;
  assign new_n2695_ = ~v16 & ~new_n2694_;
  assign new_n2696_ = ~v3 & new_n1648_;
  assign new_n2697_ = ~v3 & ~new_n2696_;
  assign new_n2698_ = ~v18 & ~new_n2697_;
  assign new_n2699_ = ~v17 & new_n2698_;
  assign new_n2700_ = v16 & new_n2699_;
  assign new_n2701_ = ~new_n2695_ & ~new_n2700_;
  assign new_n2702_ = ~v5 & ~new_n2701_;
  assign new_n2703_ = v3 & ~new_n156_;
  assign new_n2704_ = new_n402_ & ~new_n2703_;
  assign new_n2705_ = ~v18 & ~new_n2704_;
  assign new_n2706_ = ~v17 & new_n2705_;
  assign new_n2707_ = v5 & new_n2706_;
  assign new_n2708_ = ~new_n2702_ & ~new_n2707_;
  assign new_n2709_ = v15 & ~new_n2708_;
  assign new_n2710_ = v13 & new_n2709_;
  assign new_n2711_ = ~v12 & new_n2710_;
  assign new_n2712_ = ~new_n2687_ & ~new_n2711_;
  assign new_n2713_ = ~v2 & ~new_n2712_;
  assign new_n2714_ = new_n138_ & new_n849_;
  assign new_n2715_ = new_n226_ & new_n265_;
  assign new_n2716_ = v18 & v20;
  assign new_n2717_ = new_n1638_ & new_n2716_;
  assign new_n2718_ = new_n2715_ & new_n2717_;
  assign new_n2719_ = ~new_n2714_ & ~new_n2718_;
  assign new_n2720_ = v5 & ~new_n2719_;
  assign new_n2721_ = ~v15 & new_n517_;
  assign new_n2722_ = new_n265_ & new_n2721_;
  assign new_n2723_ = new_n2230_ & new_n2242_;
  assign new_n2724_ = new_n2722_ & new_n2723_;
  assign new_n2725_ = ~new_n2714_ & ~new_n2724_;
  assign new_n2726_ = ~v5 & ~new_n2725_;
  assign new_n2727_ = ~new_n2720_ & ~new_n2726_;
  assign new_n2728_ = ~v19 & ~new_n2727_;
  assign new_n2729_ = v15 & new_n1259_;
  assign new_n2730_ = v13 & new_n2729_;
  assign new_n2731_ = ~v12 & new_n2730_;
  assign new_n2732_ = ~new_n2728_ & ~new_n2731_;
  assign new_n2733_ = ~v16 & ~new_n2732_;
  assign new_n2734_ = ~new_n786_ & ~new_n2733_;
  assign new_n2735_ = ~v3 & ~new_n2734_;
  assign new_n2736_ = ~new_n793_ & ~new_n2735_;
  assign new_n2737_ = v2 & ~new_n2736_;
  assign new_n2738_ = ~new_n2713_ & ~new_n2737_;
  assign new_n2739_ = ~v4 & ~new_n2738_;
  assign new_n2740_ = v4 & new_n792_;
  assign new_n2741_ = ~new_n2739_ & ~new_n2740_;
  assign new_n2742_ = ~v1 & ~new_n2741_;
  assign new_n2743_ = ~new_n801_ & ~new_n2742_;
  assign new_n2744_ = ~v0 & ~new_n2743_;
  assign new_n2745_ = v13 & ~new_n2045_;
  assign new_n2746_ = ~v12 & new_n2745_;
  assign new_n2747_ = ~v2 & new_n2746_;
  assign new_n2748_ = ~v1 & new_n2747_;
  assign new_n2749_ = v0 & new_n2748_;
  assign new_n2750_ = ~new_n2744_ & ~new_n2749_;
  assign new_n2751_ = ~v14 & ~new_n2750_;
  assign new_n2752_ = ~v15 & ~new_n187_;
  assign new_n2753_ = v40 & ~new_n2752_;
  assign new_n2754_ = ~v18 & new_n2753_;
  assign new_n2755_ = ~v17 & new_n2754_;
  assign new_n2756_ = ~v16 & new_n2755_;
  assign new_n2757_ = v14 & new_n2756_;
  assign new_n2758_ = v13 & new_n2757_;
  assign new_n2759_ = v12 & new_n2758_;
  assign new_n2760_ = ~v5 & new_n2759_;
  assign new_n2761_ = ~v4 & new_n2760_;
  assign new_n2762_ = ~v3 & new_n2761_;
  assign new_n2763_ = ~v2 & new_n2762_;
  assign new_n2764_ = ~v1 & new_n2763_;
  assign new_n2765_ = ~v0 & new_n2764_;
  assign new_n2766_ = ~new_n2751_ & ~new_n2765_;
  assign new_n2767_ = ~v36 & ~new_n2766_;
  assign new_n2768_ = ~v11 & new_n2767_;
  assign new_n2769_ = ~v10 & new_n2768_;
  assign new_n2770_ = ~v9 & new_n2769_;
  assign \v41.25  = ~v8 & new_n2770_;
  assign new_n2772_ = v2 & v18;
  assign new_n2773_ = new_n2002_ & new_n2772_;
  assign new_n2774_ = ~v2 & new_n385_;
  assign new_n2775_ = ~new_n2773_ & ~new_n2774_;
  assign new_n2776_ = ~v5 & ~new_n2775_;
  assign new_n2777_ = ~v3 & new_n2776_;
  assign new_n2778_ = v18 & ~new_n1949_;
  assign new_n2779_ = v5 & new_n2778_;
  assign new_n2780_ = v3 & new_n2779_;
  assign new_n2781_ = ~v2 & new_n2780_;
  assign new_n2782_ = ~new_n2777_ & ~new_n2781_;
  assign new_n2783_ = v17 & ~new_n2782_;
  assign new_n2784_ = ~v15 & new_n2783_;
  assign new_n2785_ = ~v2 & new_n2673_;
  assign new_n2786_ = new_n246_ & new_n340_;
  assign new_n2787_ = new_n2785_ & new_n2786_;
  assign new_n2788_ = ~new_n2784_ & ~new_n2787_;
  assign new_n2789_ = ~v13 & ~new_n2788_;
  assign new_n2790_ = v12 & new_n2789_;
  assign new_n2791_ = ~v3 & ~new_n672_;
  assign new_n2792_ = ~v2 & new_n2791_;
  assign new_n2793_ = new_n330_ & ~new_n2792_;
  assign new_n2794_ = ~v18 & ~new_n2793_;
  assign new_n2795_ = ~v17 & new_n2794_;
  assign new_n2796_ = v15 & new_n2795_;
  assign new_n2797_ = v13 & new_n2796_;
  assign new_n2798_ = ~v12 & new_n2797_;
  assign new_n2799_ = ~new_n2790_ & ~new_n2798_;
  assign new_n2800_ = ~v16 & ~new_n2799_;
  assign new_n2801_ = ~v3 & ~new_n2791_;
  assign new_n2802_ = v15 & ~new_n2801_;
  assign new_n2803_ = ~v15 & v40;
  assign new_n2804_ = new_n2673_ & new_n2803_;
  assign new_n2805_ = ~new_n2802_ & ~new_n2804_;
  assign new_n2806_ = ~v17 & ~new_n2805_;
  assign new_n2807_ = ~v15 & new_n1409_;
  assign new_n2808_ = new_n2673_ & new_n2807_;
  assign new_n2809_ = ~new_n2806_ & ~new_n2808_;
  assign new_n2810_ = v13 & ~new_n2809_;
  assign new_n2811_ = ~v12 & new_n2810_;
  assign new_n2812_ = v17 & ~new_n740_;
  assign new_n2813_ = ~v15 & new_n2812_;
  assign new_n2814_ = ~v15 & ~new_n2813_;
  assign new_n2815_ = v40 & ~new_n2814_;
  assign new_n2816_ = ~v13 & new_n2815_;
  assign new_n2817_ = v12 & new_n2816_;
  assign new_n2818_ = ~v5 & new_n2817_;
  assign new_n2819_ = ~v3 & new_n2818_;
  assign new_n2820_ = ~new_n2811_ & ~new_n2819_;
  assign new_n2821_ = ~v18 & ~new_n2820_;
  assign new_n2822_ = v40 & ~new_n2084_;
  assign new_n2823_ = v18 & new_n2822_;
  assign new_n2824_ = ~v13 & new_n2823_;
  assign new_n2825_ = v12 & new_n2824_;
  assign new_n2826_ = ~v5 & new_n2825_;
  assign new_n2827_ = ~v3 & new_n2826_;
  assign new_n2828_ = ~new_n2821_ & ~new_n2827_;
  assign new_n2829_ = ~v2 & ~new_n2828_;
  assign new_n2830_ = v2 & new_n773_;
  assign new_n2831_ = ~new_n2829_ & ~new_n2830_;
  assign new_n2832_ = v16 & ~new_n2831_;
  assign new_n2833_ = ~new_n2800_ & ~new_n2832_;
  assign new_n2834_ = ~v19 & ~new_n2833_;
  assign new_n2835_ = v19 & ~new_n1469_;
  assign new_n2836_ = v16 & new_n2835_;
  assign new_n2837_ = v16 & ~new_n2836_;
  assign new_n2838_ = ~v12 & ~new_n2837_;
  assign new_n2839_ = ~v22 & ~new_n2649_;
  assign new_n2840_ = v29 & ~new_n2839_;
  assign new_n2841_ = v21 & new_n2840_;
  assign new_n2842_ = v20 & new_n2841_;
  assign new_n2843_ = v12 & new_n2842_;
  assign new_n2844_ = ~new_n2838_ & ~new_n2843_;
  assign new_n2845_ = ~v15 & ~new_n2844_;
  assign new_n2846_ = ~v16 & ~new_n518_;
  assign new_n2847_ = ~new_n124_ & ~new_n2846_;
  assign new_n2848_ = v19 & ~new_n2847_;
  assign new_n2849_ = v15 & new_n2848_;
  assign new_n2850_ = ~v12 & new_n2849_;
  assign new_n2851_ = ~new_n2845_ & ~new_n2850_;
  assign new_n2852_ = v40 & ~new_n2851_;
  assign new_n2853_ = ~v5 & new_n2852_;
  assign new_n2854_ = ~v12 & new_n706_;
  assign new_n2855_ = v5 & new_n2854_;
  assign new_n2856_ = ~new_n2853_ & ~new_n2855_;
  assign new_n2857_ = ~v3 & ~new_n2856_;
  assign new_n2858_ = v3 & new_n2854_;
  assign new_n2859_ = ~new_n2857_ & ~new_n2858_;
  assign new_n2860_ = ~v2 & ~new_n2859_;
  assign new_n2861_ = v2 & new_n2854_;
  assign new_n2862_ = ~new_n2860_ & ~new_n2861_;
  assign new_n2863_ = v13 & ~new_n2862_;
  assign new_n2864_ = ~v16 & ~new_n259_;
  assign new_n2865_ = ~new_n1358_ & new_n2864_;
  assign new_n2866_ = v15 & ~new_n2865_;
  assign new_n2867_ = ~new_n1823_ & ~new_n2866_;
  assign new_n2868_ = v40 & ~new_n2867_;
  assign new_n2869_ = v19 & new_n2868_;
  assign new_n2870_ = ~v13 & new_n2869_;
  assign new_n2871_ = v12 & new_n2870_;
  assign new_n2872_ = ~v5 & new_n2871_;
  assign new_n2873_ = ~v3 & new_n2872_;
  assign new_n2874_ = ~v2 & new_n2873_;
  assign new_n2875_ = ~new_n2863_ & ~new_n2874_;
  assign new_n2876_ = ~new_n2834_ & new_n2875_;
  assign new_n2877_ = ~v4 & ~new_n2876_;
  assign new_n2878_ = ~v2 & new_n2657_;
  assign new_n2879_ = new_n2006_ & new_n2878_;
  assign new_n2880_ = new_n2012_ & new_n2879_;
  assign new_n2881_ = ~new_n792_ & ~new_n2880_;
  assign new_n2882_ = v4 & ~new_n2881_;
  assign new_n2883_ = ~new_n2877_ & ~new_n2882_;
  assign new_n2884_ = ~v1 & ~new_n2883_;
  assign new_n2885_ = ~new_n801_ & ~new_n2884_;
  assign new_n2886_ = ~v14 & ~new_n2885_;
  assign new_n2887_ = ~v15 & ~new_n226_;
  assign new_n2888_ = ~v13 & ~new_n2887_;
  assign new_n2889_ = ~v12 & new_n2888_;
  assign new_n2890_ = new_n1145_ & new_n1646_;
  assign new_n2891_ = ~new_n2889_ & ~new_n2890_;
  assign new_n2892_ = v13 & v17;
  assign new_n2893_ = v12 & new_n2892_;
  assign new_n2894_ = ~v12 & new_n2386_;
  assign new_n2895_ = ~new_n2893_ & ~new_n2894_;
  assign new_n2896_ = v16 & ~new_n2895_;
  assign new_n2897_ = ~v15 & new_n2896_;
  assign new_n2898_ = new_n2891_ & ~new_n2897_;
  assign new_n2899_ = new_n1350_ & new_n1690_;
  assign new_n2900_ = new_n2898_ & ~new_n2899_;
  assign new_n2901_ = new_n1713_ & new_n2658_;
  assign new_n2902_ = ~v13 & ~new_n2901_;
  assign new_n2903_ = ~v12 & ~new_n2902_;
  assign new_n2904_ = ~new_n1107_ & ~new_n1259_;
  assign new_n2905_ = ~v16 & ~new_n2904_;
  assign new_n2906_ = ~new_n166_ & ~new_n2905_;
  assign new_n2907_ = v13 & ~new_n2906_;
  assign new_n2908_ = v13 & ~new_n2907_;
  assign new_n2909_ = v12 & ~new_n2908_;
  assign new_n2910_ = ~new_n2903_ & ~new_n2909_;
  assign new_n2911_ = ~v15 & ~new_n2910_;
  assign new_n2912_ = new_n2900_ & ~new_n2911_;
  assign new_n2913_ = v40 & ~new_n2912_;
  assign new_n2914_ = v14 & new_n2913_;
  assign new_n2915_ = ~v5 & new_n2914_;
  assign new_n2916_ = ~v4 & new_n2915_;
  assign new_n2917_ = ~v3 & new_n2916_;
  assign new_n2918_ = ~v2 & new_n2917_;
  assign new_n2919_ = ~v1 & new_n2918_;
  assign new_n2920_ = ~new_n2886_ & ~new_n2919_;
  assign new_n2921_ = ~v0 & ~new_n2920_;
  assign new_n2922_ = new_n631_ & new_n1259_;
  assign new_n2923_ = ~new_n629_ & ~new_n2922_;
  assign new_n2924_ = v16 & ~new_n2923_;
  assign new_n2925_ = ~new_n2043_ & ~new_n2924_;
  assign new_n2926_ = ~v14 & ~new_n2925_;
  assign new_n2927_ = v13 & new_n2926_;
  assign new_n2928_ = ~v12 & new_n2927_;
  assign new_n2929_ = ~v3 & new_n2928_;
  assign new_n2930_ = ~v2 & new_n2929_;
  assign new_n2931_ = ~v1 & new_n2930_;
  assign new_n2932_ = v0 & new_n2931_;
  assign new_n2933_ = ~new_n2921_ & ~new_n2932_;
  assign new_n2934_ = ~v36 & ~new_n2933_;
  assign new_n2935_ = ~v11 & new_n2934_;
  assign new_n2936_ = ~v10 & new_n2935_;
  assign new_n2937_ = ~v9 & new_n2936_;
  assign \v41.26  = ~v8 & new_n2937_;
  assign new_n2939_ = ~v19 & ~new_n1511_;
  assign new_n2940_ = v18 & new_n2939_;
  assign new_n2941_ = v17 & new_n2940_;
  assign new_n2942_ = ~v16 & new_n2941_;
  assign new_n2943_ = ~v13 & new_n2942_;
  assign new_n2944_ = v13 & v24;
  assign new_n2945_ = new_n128_ & new_n2944_;
  assign new_n2946_ = ~new_n2943_ & ~new_n2945_;
  assign new_n2947_ = new_n1911_ & new_n2658_;
  assign new_n2948_ = ~v20 & new_n2273_;
  assign new_n2949_ = v23 & new_n722_;
  assign new_n2950_ = new_n2948_ & new_n2949_;
  assign new_n2951_ = new_n2947_ & new_n2950_;
  assign new_n2952_ = ~v24 & v28;
  assign new_n2953_ = v13 & new_n2952_;
  assign new_n2954_ = ~new_n2951_ & ~new_n2953_;
  assign new_n2955_ = v23 & new_n1222_;
  assign new_n2956_ = v22 & new_n2955_;
  assign new_n2957_ = ~v20 & new_n2956_;
  assign new_n2958_ = ~v20 & ~new_n2957_;
  assign new_n2959_ = v21 & ~new_n2958_;
  assign new_n2960_ = ~v19 & new_n2959_;
  assign new_n2961_ = ~v19 & ~new_n2960_;
  assign new_n2962_ = v18 & ~new_n2961_;
  assign new_n2963_ = v18 & ~new_n2962_;
  assign new_n2964_ = ~v16 & ~new_n2963_;
  assign new_n2965_ = ~v16 & ~new_n2964_;
  assign new_n2966_ = v17 & ~new_n2965_;
  assign new_n2967_ = v17 & ~new_n2966_;
  assign new_n2968_ = ~v13 & ~new_n2967_;
  assign new_n2969_ = ~v25 & v28;
  assign new_n2970_ = v24 & new_n2969_;
  assign new_n2971_ = v28 & ~new_n2970_;
  assign new_n2972_ = v13 & ~new_n2971_;
  assign new_n2973_ = ~new_n2968_ & ~new_n2972_;
  assign new_n2974_ = new_n2954_ & new_n2973_;
  assign new_n2975_ = new_n2946_ & new_n2974_;
  assign new_n2976_ = v12 & ~new_n2975_;
  assign new_n2977_ = v13 & ~v16;
  assign new_n2978_ = new_n1319_ & ~new_n2977_;
  assign new_n2979_ = ~v12 & ~new_n2978_;
  assign new_n2980_ = ~new_n2976_ & ~new_n2979_;
  assign new_n2981_ = ~v15 & ~new_n2980_;
  assign new_n2982_ = ~v12 & ~new_n1319_;
  assign new_n2983_ = ~v13 & v16;
  assign new_n2984_ = v12 & new_n2983_;
  assign new_n2985_ = ~new_n2982_ & ~new_n2984_;
  assign new_n2986_ = ~new_n265_ & ~new_n849_;
  assign new_n2987_ = v17 & ~new_n2986_;
  assign new_n2988_ = ~v16 & new_n2987_;
  assign new_n2989_ = new_n2985_ & ~new_n2988_;
  assign new_n2990_ = v37 & new_n843_;
  assign new_n2991_ = ~v39 & ~new_n2990_;
  assign new_n2992_ = ~v38 & new_n2991_;
  assign new_n2993_ = v18 & ~new_n2992_;
  assign new_n2994_ = v18 & ~new_n2993_;
  assign new_n2995_ = v13 & ~new_n2994_;
  assign new_n2996_ = ~v12 & new_n2995_;
  assign new_n2997_ = v12 & new_n2590_;
  assign new_n2998_ = ~new_n2996_ & ~new_n2997_;
  assign new_n2999_ = ~v17 & ~new_n2998_;
  assign new_n3000_ = ~v16 & new_n2999_;
  assign new_n3001_ = new_n2989_ & ~new_n3000_;
  assign new_n3002_ = ~v19 & ~new_n2992_;
  assign new_n3003_ = ~v19 & ~new_n3002_;
  assign new_n3004_ = ~v18 & ~new_n3003_;
  assign new_n3005_ = ~v17 & new_n3004_;
  assign new_n3006_ = ~v16 & new_n3005_;
  assign new_n3007_ = ~v13 & new_n3006_;
  assign new_n3008_ = ~v13 & ~new_n3007_;
  assign new_n3009_ = v12 & ~new_n3008_;
  assign new_n3010_ = new_n3001_ & ~new_n3009_;
  assign new_n3011_ = v15 & ~new_n3010_;
  assign new_n3012_ = ~new_n2981_ & ~new_n3011_;
  assign new_n3013_ = ~v14 & ~new_n3012_;
  assign new_n3014_ = ~new_n1472_ & ~new_n1646_;
  assign new_n3015_ = new_n2986_ & new_n3014_;
  assign new_n3016_ = v14 & ~new_n3015_;
  assign new_n3017_ = ~new_n3013_ & ~new_n3016_;
  assign new_n3018_ = v40 & ~new_n3017_;
  assign new_n3019_ = v40 & ~new_n3018_;
  assign new_n3020_ = ~v10 & ~new_n3019_;
  assign new_n3021_ = ~v8 & new_n3020_;
  assign new_n3022_ = ~v8 & ~new_n3021_;
  assign new_n3023_ = ~v5 & ~new_n3022_;
  assign new_n3024_ = ~v12 & new_n333_;
  assign new_n3025_ = ~v14 & new_n2078_;
  assign new_n3026_ = v12 & new_n3025_;
  assign new_n3027_ = ~new_n3024_ & ~new_n3026_;
  assign new_n3028_ = ~v15 & ~new_n3027_;
  assign new_n3029_ = ~v14 & v19;
  assign new_n3030_ = v12 & new_n3029_;
  assign new_n3031_ = ~new_n1813_ & ~new_n3030_;
  assign new_n3032_ = v40 & ~new_n3031_;
  assign new_n3033_ = v15 & new_n3032_;
  assign new_n3034_ = ~new_n3028_ & ~new_n3033_;
  assign new_n3035_ = ~v16 & ~new_n3034_;
  assign new_n3036_ = v12 & new_n1356_;
  assign new_n3037_ = ~new_n1813_ & ~new_n3036_;
  assign new_n3038_ = v40 & ~new_n3037_;
  assign new_n3039_ = v16 & new_n3038_;
  assign new_n3040_ = ~new_n3035_ & ~new_n3039_;
  assign new_n3041_ = v18 & ~new_n3040_;
  assign new_n3042_ = ~new_n1811_ & ~new_n1813_;
  assign new_n3043_ = v40 & ~new_n3042_;
  assign new_n3044_ = new_n1810_ & new_n1874_;
  assign new_n3045_ = ~new_n3043_ & ~new_n3044_;
  assign new_n3046_ = ~v18 & ~new_n3045_;
  assign new_n3047_ = ~new_n3041_ & ~new_n3046_;
  assign new_n3048_ = v17 & ~new_n3047_;
  assign new_n3049_ = v40 & ~new_n1812_;
  assign new_n3050_ = ~v16 & new_n120_;
  assign new_n3051_ = new_n3036_ & new_n3050_;
  assign new_n3052_ = ~new_n3049_ & ~new_n3051_;
  assign new_n3053_ = ~v17 & ~new_n3052_;
  assign new_n3054_ = ~new_n3048_ & ~new_n3053_;
  assign new_n3055_ = ~v13 & ~new_n3054_;
  assign new_n3056_ = new_n842_ & new_n952_;
  assign new_n3057_ = v12 & new_n900_;
  assign new_n3058_ = new_n1099_ & new_n3057_;
  assign new_n3059_ = ~new_n3056_ & ~new_n3058_;
  assign new_n3060_ = ~v15 & new_n953_;
  assign new_n3061_ = ~v15 & ~new_n3060_;
  assign new_n3062_ = v40 & ~new_n3061_;
  assign new_n3063_ = v17 & new_n3062_;
  assign new_n3064_ = v14 & new_n3063_;
  assign new_n3065_ = v12 & new_n3064_;
  assign new_n3066_ = ~v12 & new_n1356_;
  assign new_n3067_ = new_n124_ & new_n3066_;
  assign new_n3068_ = ~new_n3065_ & ~new_n3067_;
  assign new_n3069_ = new_n3059_ & new_n3068_;
  assign new_n3070_ = v16 & ~new_n1866_;
  assign new_n3071_ = ~v15 & new_n3070_;
  assign new_n3072_ = new_n117_ & new_n1038_;
  assign new_n3073_ = ~new_n3071_ & ~new_n3072_;
  assign new_n3074_ = v17 & ~new_n3073_;
  assign new_n3075_ = ~v14 & new_n3074_;
  assign new_n3076_ = ~v12 & new_n3075_;
  assign new_n3077_ = v12 & v14;
  assign new_n3078_ = new_n116_ & new_n3077_;
  assign new_n3079_ = new_n119_ & new_n1648_;
  assign new_n3080_ = new_n3078_ & new_n3079_;
  assign new_n3081_ = ~new_n3076_ & ~new_n3080_;
  assign new_n3082_ = new_n3069_ & new_n3081_;
  assign new_n3083_ = v13 & ~new_n3082_;
  assign new_n3084_ = ~new_n3055_ & ~new_n3083_;
  assign new_n3085_ = ~v10 & ~new_n3084_;
  assign new_n3086_ = ~v8 & new_n3085_;
  assign new_n3087_ = v5 & new_n3086_;
  assign new_n3088_ = ~new_n3023_ & ~new_n3087_;
  assign new_n3089_ = ~v4 & ~new_n3088_;
  assign new_n3090_ = ~v15 & ~new_n1529_;
  assign new_n3091_ = ~v13 & new_n3090_;
  assign new_n3092_ = v12 & new_n3091_;
  assign new_n3093_ = ~new_n2210_ & ~new_n3092_;
  assign new_n3094_ = ~v19 & ~new_n3093_;
  assign new_n3095_ = ~new_n2546_ & ~new_n3094_;
  assign new_n3096_ = v17 & ~new_n3095_;
  assign new_n3097_ = ~v12 & new_n2592_;
  assign new_n3098_ = new_n120_ & new_n265_;
  assign new_n3099_ = ~new_n3097_ & ~new_n3098_;
  assign new_n3100_ = ~v17 & ~new_n3099_;
  assign new_n3101_ = v15 & new_n3100_;
  assign new_n3102_ = ~new_n3096_ & ~new_n3101_;
  assign new_n3103_ = ~v16 & ~new_n3102_;
  assign new_n3104_ = ~new_n786_ & ~new_n3103_;
  assign new_n3105_ = ~v14 & ~new_n3104_;
  assign new_n3106_ = ~v10 & new_n3105_;
  assign new_n3107_ = ~v8 & new_n3106_;
  assign new_n3108_ = v4 & new_n3107_;
  assign new_n3109_ = ~new_n3089_ & ~new_n3108_;
  assign new_n3110_ = ~v3 & ~new_n3109_;
  assign new_n3111_ = ~new_n681_ & ~new_n1223_;
  assign new_n3112_ = ~new_n1544_ & ~new_n3111_;
  assign new_n3113_ = v21 & ~new_n3112_;
  assign new_n3114_ = ~v20 & new_n3113_;
  assign new_n3115_ = ~new_n1239_ & ~new_n3114_;
  assign new_n3116_ = ~v19 & ~new_n3115_;
  assign new_n3117_ = v18 & new_n3116_;
  assign new_n3118_ = v17 & new_n3117_;
  assign new_n3119_ = ~v15 & new_n3118_;
  assign new_n3120_ = ~v13 & new_n3119_;
  assign new_n3121_ = v12 & new_n3120_;
  assign new_n3122_ = ~v4 & new_n3121_;
  assign new_n3123_ = new_n781_ & ~new_n3122_;
  assign new_n3124_ = ~v16 & ~new_n3123_;
  assign new_n3125_ = ~new_n786_ & ~new_n3124_;
  assign new_n3126_ = v21 & ~new_n1220_;
  assign new_n3127_ = ~v20 & new_n3126_;
  assign new_n3128_ = v18 & new_n3127_;
  assign new_n3129_ = ~v4 & ~v18;
  assign new_n3130_ = ~new_n3128_ & ~new_n3129_;
  assign new_n3131_ = ~v15 & ~new_n3130_;
  assign new_n3132_ = ~v13 & new_n3131_;
  assign new_n3133_ = v12 & new_n3132_;
  assign new_n3134_ = ~v4 & new_n2210_;
  assign new_n3135_ = ~new_n3133_ & ~new_n3134_;
  assign new_n3136_ = ~v19 & ~new_n3135_;
  assign new_n3137_ = ~v4 & new_n849_;
  assign new_n3138_ = new_n2545_ & new_n3137_;
  assign new_n3139_ = ~new_n3136_ & ~new_n3138_;
  assign new_n3140_ = v17 & ~new_n3139_;
  assign new_n3141_ = ~v16 & new_n3140_;
  assign new_n3142_ = ~v5 & new_n3141_;
  assign new_n3143_ = new_n3125_ & ~new_n3142_;
  assign new_n3144_ = ~v14 & ~new_n3143_;
  assign new_n3145_ = ~v10 & new_n3144_;
  assign new_n3146_ = ~v8 & new_n3145_;
  assign new_n3147_ = v3 & new_n3146_;
  assign new_n3148_ = ~new_n3110_ & ~new_n3147_;
  assign new_n3149_ = ~v2 & ~new_n3148_;
  assign new_n3150_ = v21 & new_n1553_;
  assign new_n3151_ = ~v20 & new_n3150_;
  assign new_n3152_ = ~v19 & new_n3151_;
  assign new_n3153_ = v18 & new_n3152_;
  assign new_n3154_ = v17 & new_n3153_;
  assign new_n3155_ = ~v16 & new_n3154_;
  assign new_n3156_ = ~v15 & new_n3155_;
  assign new_n3157_ = ~v13 & new_n3156_;
  assign new_n3158_ = v12 & new_n3157_;
  assign new_n3159_ = ~v5 & new_n3158_;
  assign new_n3160_ = ~v4 & new_n3159_;
  assign new_n3161_ = ~v3 & new_n3160_;
  assign new_n3162_ = new_n2005_ & ~new_n3161_;
  assign new_n3163_ = ~v14 & ~new_n3162_;
  assign new_n3164_ = ~v10 & new_n3163_;
  assign new_n3165_ = ~v8 & new_n3164_;
  assign new_n3166_ = v2 & new_n3165_;
  assign new_n3167_ = ~new_n3149_ & ~new_n3166_;
  assign new_n3168_ = ~v1 & ~new_n3167_;
  assign new_n3169_ = ~v10 & new_n2032_;
  assign new_n3170_ = ~v8 & new_n3169_;
  assign new_n3171_ = v1 & new_n3170_;
  assign new_n3172_ = ~new_n3168_ & ~new_n3171_;
  assign new_n3173_ = ~v0 & ~new_n3172_;
  assign new_n3174_ = ~new_n269_ & ~new_n2746_;
  assign new_n3175_ = ~v14 & ~new_n3174_;
  assign new_n3176_ = ~v10 & new_n3175_;
  assign new_n3177_ = ~v8 & new_n3176_;
  assign new_n3178_ = ~v2 & new_n3177_;
  assign new_n3179_ = ~v1 & new_n3178_;
  assign new_n3180_ = v0 & new_n3179_;
  assign new_n3181_ = ~new_n3173_ & ~new_n3180_;
  assign new_n3182_ = ~v36 & ~new_n3181_;
  assign new_n3183_ = ~v10 & v36;
  assign new_n3184_ = ~v10 & ~new_n3183_;
  assign new_n3185_ = ~v8 & ~new_n3184_;
  assign new_n3186_ = ~new_n3182_ & ~new_n3185_;
  assign new_n3187_ = ~v11 & ~new_n3186_;
  assign new_n3188_ = v11 & ~new_n1309_;
  assign new_n3189_ = ~new_n3187_ & ~new_n3188_;
  assign new_n3190_ = ~v9 & ~new_n3189_;
  assign new_n3191_ = v10 & ~v11;
  assign new_n3192_ = new_n2340_ & new_n3191_;
  assign \v41.27  = new_n3190_ | new_n3192_;
  assign new_n3194_ = v40 & ~new_n1730_;
  assign new_n3195_ = ~v39 & new_n3194_;
  assign new_n3196_ = ~v38 & new_n3195_;
  assign new_n3197_ = ~v37 & new_n3196_;
  assign new_n3198_ = ~v36 & new_n3197_;
  assign new_n3199_ = ~v17 & new_n3198_;
  assign new_n3200_ = ~v16 & new_n3199_;
  assign new_n3201_ = v15 & new_n3200_;
  assign new_n3202_ = ~v14 & new_n3201_;
  assign new_n3203_ = ~v11 & new_n3202_;
  assign new_n3204_ = ~v10 & new_n3203_;
  assign new_n3205_ = ~v5 & new_n3204_;
  assign new_n3206_ = ~v4 & new_n3205_;
  assign new_n3207_ = ~v3 & new_n3206_;
  assign new_n3208_ = ~v2 & new_n3207_;
  assign new_n3209_ = ~v1 & new_n3208_;
  assign new_n3210_ = ~v0 & new_n3209_;
  assign new_n3211_ = ~v10 & ~new_n3210_;
  assign new_n3212_ = ~v9 & ~new_n3211_;
  assign new_n3213_ = ~new_n840_ & ~new_n3212_;
  assign \v41.28  = ~v8 & ~new_n3213_;
  assign new_n3215_ = v18 & ~new_n1518_;
  assign new_n3216_ = ~v15 & ~new_n3215_;
  assign new_n3217_ = ~v13 & new_n3216_;
  assign new_n3218_ = v12 & new_n3217_;
  assign new_n3219_ = ~new_n2210_ & ~new_n3218_;
  assign new_n3220_ = ~v19 & ~new_n3219_;
  assign new_n3221_ = ~new_n2546_ & ~new_n3220_;
  assign new_n3222_ = v17 & ~new_n3221_;
  assign new_n3223_ = ~new_n3101_ & ~new_n3222_;
  assign new_n3224_ = ~v16 & ~new_n3223_;
  assign new_n3225_ = v13 & new_n1964_;
  assign new_n3226_ = ~v12 & new_n3225_;
  assign new_n3227_ = ~new_n3224_ & ~new_n3226_;
  assign new_n3228_ = ~new_n672_ & ~new_n3227_;
  assign new_n3229_ = ~v18 & ~new_n1572_;
  assign new_n3230_ = v17 & ~new_n3229_;
  assign new_n3231_ = v17 & ~new_n3230_;
  assign new_n3232_ = ~new_n156_ & ~new_n3231_;
  assign new_n3233_ = ~v16 & new_n976_;
  assign new_n3234_ = ~new_n400_ & ~new_n3233_;
  assign new_n3235_ = ~v38 & new_n740_;
  assign new_n3236_ = ~v19 & ~new_n3235_;
  assign new_n3237_ = ~v18 & new_n3236_;
  assign new_n3238_ = v17 & new_n3237_;
  assign new_n3239_ = v16 & new_n3238_;
  assign new_n3240_ = new_n3234_ & ~new_n3239_;
  assign new_n3241_ = ~new_n3232_ & new_n3240_;
  assign new_n3242_ = ~v13 & ~new_n3241_;
  assign new_n3243_ = ~v13 & ~new_n3242_;
  assign new_n3244_ = v12 & ~new_n3243_;
  assign new_n3245_ = ~new_n1106_ & ~new_n1319_;
  assign new_n3246_ = v13 & new_n164_;
  assign new_n3247_ = v13 & ~new_n3246_;
  assign new_n3248_ = ~new_n1866_ & ~new_n3247_;
  assign new_n3249_ = ~new_n2977_ & ~new_n3248_;
  assign new_n3250_ = ~new_n3245_ & new_n3249_;
  assign new_n3251_ = ~v12 & ~new_n3250_;
  assign new_n3252_ = ~new_n3244_ & ~new_n3251_;
  assign new_n3253_ = ~v15 & ~new_n3252_;
  assign new_n3254_ = v17 & ~new_n1320_;
  assign new_n3255_ = v18 & ~new_n3254_;
  assign new_n3256_ = ~new_n1325_ & ~new_n3255_;
  assign new_n3257_ = ~v12 & ~new_n3256_;
  assign new_n3258_ = ~v13 & ~new_n1867_;
  assign new_n3259_ = v12 & new_n3258_;
  assign new_n3260_ = ~new_n3257_ & ~new_n3259_;
  assign new_n3261_ = ~v12 & v17;
  assign new_n3262_ = new_n120_ & new_n3261_;
  assign new_n3263_ = ~v12 & ~new_n3262_;
  assign new_n3264_ = v13 & ~new_n3263_;
  assign new_n3265_ = ~v17 & ~new_n1177_;
  assign new_n3266_ = ~v13 & new_n3265_;
  assign new_n3267_ = v12 & new_n3266_;
  assign new_n3268_ = ~new_n3264_ & ~new_n3267_;
  assign new_n3269_ = ~v16 & ~new_n3268_;
  assign new_n3270_ = v12 & new_n220_;
  assign new_n3271_ = ~new_n3269_ & ~new_n3270_;
  assign new_n3272_ = new_n3260_ & new_n3271_;
  assign new_n3273_ = v15 & ~new_n3272_;
  assign new_n3274_ = ~new_n3253_ & ~new_n3273_;
  assign new_n3275_ = ~v5 & ~new_n3274_;
  assign new_n3276_ = new_n120_ & new_n209_;
  assign new_n3277_ = ~v16 & ~new_n3276_;
  assign new_n3278_ = v15 & ~new_n3277_;
  assign new_n3279_ = ~v13 & new_n3278_;
  assign new_n3280_ = v12 & new_n3279_;
  assign new_n3281_ = v5 & new_n3280_;
  assign new_n3282_ = ~new_n3275_ & ~new_n3281_;
  assign new_n3283_ = v40 & ~new_n3282_;
  assign new_n3284_ = ~new_n3228_ & ~new_n3283_;
  assign new_n3285_ = ~v14 & ~new_n3284_;
  assign new_n3286_ = ~v5 & ~new_n3014_;
  assign new_n3287_ = new_n821_ & new_n1492_;
  assign new_n3288_ = ~new_n3286_ & ~new_n3287_;
  assign new_n3289_ = v12 & new_n1694_;
  assign new_n3290_ = ~new_n2597_ & ~new_n3289_;
  assign new_n3291_ = v17 & ~new_n3290_;
  assign new_n3292_ = v5 & new_n3291_;
  assign new_n3293_ = new_n3288_ & ~new_n3292_;
  assign new_n3294_ = v5 & new_n2897_;
  assign new_n3295_ = new_n3293_ & ~new_n3294_;
  assign new_n3296_ = v5 & new_n1646_;
  assign new_n3297_ = new_n1823_ & new_n3296_;
  assign new_n3298_ = new_n3295_ & ~new_n3297_;
  assign new_n3299_ = ~v5 & ~new_n2986_;
  assign new_n3300_ = ~new_n2615_ & ~new_n3299_;
  assign new_n3301_ = new_n3298_ & new_n3300_;
  assign new_n3302_ = v40 & ~new_n3301_;
  assign new_n3303_ = v14 & new_n3302_;
  assign new_n3304_ = ~new_n2187_ & ~new_n3303_;
  assign new_n3305_ = ~new_n3285_ & new_n3304_;
  assign new_n3306_ = ~v4 & ~new_n3305_;
  assign new_n3307_ = v4 & new_n3105_;
  assign new_n3308_ = ~new_n3306_ & ~new_n3307_;
  assign new_n3309_ = ~v3 & ~new_n3308_;
  assign new_n3310_ = v3 & new_n3144_;
  assign new_n3311_ = ~new_n3309_ & ~new_n3310_;
  assign new_n3312_ = ~v2 & ~new_n3311_;
  assign new_n3313_ = v2 & new_n3163_;
  assign new_n3314_ = ~new_n3312_ & ~new_n3313_;
  assign new_n3315_ = ~v1 & ~new_n3314_;
  assign new_n3316_ = ~new_n2033_ & ~new_n3315_;
  assign new_n3317_ = ~v0 & ~new_n3316_;
  assign new_n3318_ = ~v2 & new_n3175_;
  assign new_n3319_ = ~v1 & new_n3318_;
  assign new_n3320_ = v0 & new_n3319_;
  assign new_n3321_ = ~new_n3317_ & ~new_n3320_;
  assign new_n3322_ = ~v36 & ~new_n3321_;
  assign new_n3323_ = ~v36 & ~new_n3322_;
  assign new_n3324_ = ~v10 & ~new_n3323_;
  assign new_n3325_ = ~v10 & ~new_n3324_;
  assign new_n3326_ = ~v9 & ~new_n3325_;
  assign new_n3327_ = ~v9 & ~new_n3326_;
  assign new_n3328_ = ~v11 & ~new_n3327_;
  assign new_n3329_ = ~new_n2297_ & ~new_n3328_;
  assign new_n3330_ = ~v8 & ~new_n3329_;
  assign \v41.29  = new_n2307_ | new_n3330_;
  assign new_n3332_ = v39 & ~new_n1365_;
  assign new_n3333_ = new_n1365_ & new_n3332_;
  assign new_n3334_ = v17 & ~new_n3333_;
  assign new_n3335_ = v17 & ~new_n3334_;
  assign new_n3336_ = v40 & ~new_n3335_;
  assign new_n3337_ = ~v36 & new_n3336_;
  assign new_n3338_ = v19 & new_n3337_;
  assign new_n3339_ = ~v18 & new_n3338_;
  assign new_n3340_ = ~v16 & new_n3339_;
  assign new_n3341_ = ~v15 & new_n3340_;
  assign new_n3342_ = ~v14 & new_n3341_;
  assign new_n3343_ = ~v13 & new_n3342_;
  assign new_n3344_ = v12 & new_n3343_;
  assign new_n3345_ = ~v11 & new_n3344_;
  assign new_n3346_ = ~v10 & new_n3345_;
  assign new_n3347_ = ~v9 & new_n3346_;
  assign new_n3348_ = ~v8 & new_n3347_;
  assign new_n3349_ = ~v5 & new_n3348_;
  assign new_n3350_ = ~v4 & new_n3349_;
  assign new_n3351_ = ~v3 & new_n3350_;
  assign new_n3352_ = ~v2 & new_n3351_;
  assign new_n3353_ = ~v1 & new_n3352_;
  assign \v41.30  = ~v0 & new_n3353_;
  assign new_n3355_ = ~v5 & new_n3346_;
  assign new_n3356_ = ~v4 & new_n3355_;
  assign new_n3357_ = ~v3 & new_n3356_;
  assign new_n3358_ = ~v2 & new_n3357_;
  assign new_n3359_ = ~v1 & new_n3358_;
  assign new_n3360_ = ~v0 & new_n3359_;
  assign new_n3361_ = ~v10 & ~new_n3360_;
  assign new_n3362_ = ~v9 & ~new_n3361_;
  assign \v41.33  = ~v8 & new_n3362_;
  assign new_n3364_ = ~new_n883_ & new_n1867_;
  assign new_n3365_ = ~v13 & ~new_n3364_;
  assign new_n3366_ = v12 & new_n3365_;
  assign new_n3367_ = v12 & ~new_n3366_;
  assign new_n3368_ = ~v13 & new_n1767_;
  assign new_n3369_ = ~v13 & ~new_n3368_;
  assign new_n3370_ = v12 & ~new_n3369_;
  assign new_n3371_ = new_n3367_ & ~new_n3370_;
  assign new_n3372_ = v15 & ~new_n3371_;
  assign new_n3373_ = ~new_n2981_ & ~new_n3372_;
  assign new_n3374_ = ~v14 & ~new_n3373_;
  assign new_n3375_ = ~new_n3016_ & ~new_n3374_;
  assign new_n3376_ = v40 & ~new_n3375_;
  assign new_n3377_ = v40 & ~new_n3376_;
  assign new_n3378_ = ~v10 & ~new_n3377_;
  assign new_n3379_ = ~v8 & new_n3378_;
  assign new_n3380_ = ~v8 & ~new_n3379_;
  assign new_n3381_ = ~v5 & ~new_n3380_;
  assign new_n3382_ = ~new_n3087_ & ~new_n3381_;
  assign new_n3383_ = ~v4 & ~new_n3382_;
  assign new_n3384_ = ~new_n3108_ & ~new_n3383_;
  assign new_n3385_ = ~v3 & ~new_n3384_;
  assign new_n3386_ = ~new_n3147_ & ~new_n3385_;
  assign new_n3387_ = ~v2 & ~new_n3386_;
  assign new_n3388_ = ~new_n3166_ & ~new_n3387_;
  assign new_n3389_ = ~v1 & ~new_n3388_;
  assign new_n3390_ = ~new_n3171_ & ~new_n3389_;
  assign new_n3391_ = ~v0 & ~new_n3390_;
  assign new_n3392_ = ~new_n3180_ & ~new_n3391_;
  assign new_n3393_ = ~v36 & ~new_n3392_;
  assign new_n3394_ = ~new_n3185_ & ~new_n3393_;
  assign new_n3395_ = ~v11 & ~new_n3394_;
  assign new_n3396_ = ~new_n3188_ & ~new_n3395_;
  assign new_n3397_ = ~v9 & ~new_n3396_;
  assign \v41.34  = new_n3192_ | new_n3397_;
  assign new_n3399_ = ~new_n1311_ & ~new_n2295_;
  assign new_n3400_ = ~new_n1392_ & new_n3399_;
  assign \v41.35  = ~v8 & ~new_n3400_;
  assign new_n3402_ = v15 & new_n1372_;
  assign new_n3403_ = ~v15 & new_n120_;
  assign new_n3404_ = ~new_n3402_ & ~new_n3403_;
  assign new_n3405_ = v40 & ~new_n3404_;
  assign new_n3406_ = ~v36 & new_n3405_;
  assign new_n3407_ = ~v17 & new_n3406_;
  assign new_n3408_ = ~v16 & new_n3407_;
  assign new_n3409_ = ~v14 & new_n3408_;
  assign new_n3410_ = ~v13 & new_n3409_;
  assign new_n3411_ = v12 & new_n3410_;
  assign new_n3412_ = ~v11 & new_n3411_;
  assign new_n3413_ = ~v10 & new_n3412_;
  assign new_n3414_ = ~v5 & new_n3413_;
  assign new_n3415_ = ~v4 & new_n3414_;
  assign new_n3416_ = ~v3 & new_n3415_;
  assign new_n3417_ = ~v2 & new_n3416_;
  assign new_n3418_ = ~v1 & new_n3417_;
  assign new_n3419_ = ~v0 & new_n3418_;
  assign new_n3420_ = ~v10 & ~new_n3419_;
  assign new_n3421_ = ~v9 & ~new_n3420_;
  assign new_n3422_ = ~new_n840_ & ~new_n3421_;
  assign \v41.36  = ~v8 & ~new_n3422_;
  assign new_n3424_ = v18 & ~new_n1452_;
  assign new_n3425_ = v18 & ~new_n3424_;
  assign new_n3426_ = v13 & ~new_n3425_;
  assign new_n3427_ = ~v12 & new_n3426_;
  assign new_n3428_ = ~new_n2997_ & ~new_n3427_;
  assign new_n3429_ = ~v17 & ~new_n3428_;
  assign new_n3430_ = ~v16 & new_n3429_;
  assign new_n3431_ = new_n2989_ & ~new_n3430_;
  assign new_n3432_ = ~new_n3370_ & new_n3431_;
  assign new_n3433_ = v15 & ~new_n3432_;
  assign new_n3434_ = ~new_n2981_ & ~new_n3433_;
  assign new_n3435_ = ~v14 & ~new_n3434_;
  assign new_n3436_ = ~new_n3016_ & ~new_n3435_;
  assign new_n3437_ = v40 & ~new_n3436_;
  assign new_n3438_ = v40 & ~new_n3437_;
  assign new_n3439_ = ~v11 & ~new_n3438_;
  assign new_n3440_ = ~v10 & new_n3439_;
  assign new_n3441_ = ~v8 & new_n3440_;
  assign new_n3442_ = ~v8 & ~new_n3441_;
  assign new_n3443_ = ~v5 & ~new_n3442_;
  assign new_n3444_ = ~v11 & ~new_n3084_;
  assign new_n3445_ = ~v10 & new_n3444_;
  assign new_n3446_ = ~v8 & new_n3445_;
  assign new_n3447_ = v5 & new_n3446_;
  assign new_n3448_ = ~new_n3443_ & ~new_n3447_;
  assign new_n3449_ = ~v4 & ~new_n3448_;
  assign new_n3450_ = ~v11 & new_n3105_;
  assign new_n3451_ = ~v10 & new_n3450_;
  assign new_n3452_ = ~v8 & new_n3451_;
  assign new_n3453_ = v4 & new_n3452_;
  assign new_n3454_ = ~new_n3449_ & ~new_n3453_;
  assign new_n3455_ = ~v3 & ~new_n3454_;
  assign new_n3456_ = ~v11 & new_n3144_;
  assign new_n3457_ = ~v10 & new_n3456_;
  assign new_n3458_ = ~v8 & new_n3457_;
  assign new_n3459_ = v3 & new_n3458_;
  assign new_n3460_ = ~new_n3455_ & ~new_n3459_;
  assign new_n3461_ = ~v2 & ~new_n3460_;
  assign new_n3462_ = ~v11 & new_n3163_;
  assign new_n3463_ = ~v10 & new_n3462_;
  assign new_n3464_ = ~v8 & new_n3463_;
  assign new_n3465_ = v2 & new_n3464_;
  assign new_n3466_ = ~new_n3461_ & ~new_n3465_;
  assign new_n3467_ = ~v1 & ~new_n3466_;
  assign new_n3468_ = ~v11 & new_n2032_;
  assign new_n3469_ = ~v10 & new_n3468_;
  assign new_n3470_ = ~v8 & new_n3469_;
  assign new_n3471_ = v1 & new_n3470_;
  assign new_n3472_ = ~new_n3467_ & ~new_n3471_;
  assign new_n3473_ = ~v0 & ~new_n3472_;
  assign new_n3474_ = ~v11 & new_n3175_;
  assign new_n3475_ = ~v10 & new_n3474_;
  assign new_n3476_ = ~v8 & new_n3475_;
  assign new_n3477_ = ~v2 & new_n3476_;
  assign new_n3478_ = ~v1 & new_n3477_;
  assign new_n3479_ = v0 & new_n3478_;
  assign new_n3480_ = ~new_n3473_ & ~new_n3479_;
  assign new_n3481_ = ~v36 & ~new_n3480_;
  assign new_n3482_ = ~v8 & ~v10;
  assign new_n3483_ = ~v11 & v36;
  assign new_n3484_ = new_n3482_ & new_n3483_;
  assign new_n3485_ = ~new_n3481_ & ~new_n3484_;
  assign new_n3486_ = ~v9 & ~new_n3485_;
  assign \v41.37  = new_n3192_ | new_n3486_;
  assign new_n3488_ = ~v16 & ~new_n486_;
  assign new_n3489_ = ~v17 & ~new_n3488_;
  assign new_n3490_ = ~new_n2966_ & ~new_n3489_;
  assign new_n3491_ = ~v13 & ~new_n3490_;
  assign new_n3492_ = ~new_n2972_ & ~new_n3491_;
  assign new_n3493_ = new_n2954_ & new_n3492_;
  assign new_n3494_ = new_n2946_ & new_n3493_;
  assign new_n3495_ = v12 & ~new_n3494_;
  assign new_n3496_ = ~new_n2979_ & ~new_n3495_;
  assign new_n3497_ = ~v15 & ~new_n3496_;
  assign new_n3498_ = ~v17 & new_n2125_;
  assign new_n3499_ = ~v16 & new_n3498_;
  assign new_n3500_ = ~v13 & new_n3499_;
  assign new_n3501_ = ~v13 & ~new_n3500_;
  assign new_n3502_ = v12 & ~new_n3501_;
  assign new_n3503_ = new_n3431_ & ~new_n3502_;
  assign new_n3504_ = v15 & ~new_n3503_;
  assign new_n3505_ = ~new_n3497_ & ~new_n3504_;
  assign new_n3506_ = ~v14 & ~new_n3505_;
  assign new_n3507_ = ~new_n3016_ & ~new_n3506_;
  assign new_n3508_ = v40 & ~new_n3507_;
  assign new_n3509_ = v40 & ~new_n3508_;
  assign new_n3510_ = ~v11 & ~new_n3509_;
  assign new_n3511_ = ~v10 & new_n3510_;
  assign new_n3512_ = ~v8 & new_n3511_;
  assign new_n3513_ = ~v8 & ~new_n3512_;
  assign new_n3514_ = ~v5 & ~new_n3513_;
  assign new_n3515_ = ~new_n3447_ & ~new_n3514_;
  assign new_n3516_ = ~v4 & ~new_n3515_;
  assign new_n3517_ = ~new_n3453_ & ~new_n3516_;
  assign new_n3518_ = ~v3 & ~new_n3517_;
  assign new_n3519_ = ~new_n3459_ & ~new_n3518_;
  assign new_n3520_ = ~v2 & ~new_n3519_;
  assign new_n3521_ = ~new_n3465_ & ~new_n3520_;
  assign new_n3522_ = ~v1 & ~new_n3521_;
  assign new_n3523_ = ~new_n3471_ & ~new_n3522_;
  assign new_n3524_ = ~v0 & ~new_n3523_;
  assign new_n3525_ = ~new_n3479_ & ~new_n3524_;
  assign new_n3526_ = ~v36 & ~new_n3525_;
  assign new_n3527_ = ~new_n3484_ & ~new_n3526_;
  assign new_n3528_ = ~v9 & ~new_n3527_;
  assign \v41.38  = new_n3192_ | new_n3528_;
  assign new_n3530_ = ~v18 & new_n843_;
  assign new_n3531_ = v15 & new_n3530_;
  assign new_n3532_ = ~v15 & v18;
  assign new_n3533_ = ~new_n3531_ & ~new_n3532_;
  assign new_n3534_ = ~v19 & ~new_n3533_;
  assign new_n3535_ = ~new_n3403_ & ~new_n3534_;
  assign new_n3536_ = v40 & ~new_n3535_;
  assign new_n3537_ = ~v36 & new_n3536_;
  assign new_n3538_ = ~v17 & new_n3537_;
  assign new_n3539_ = ~v16 & new_n3538_;
  assign new_n3540_ = ~v14 & new_n3539_;
  assign new_n3541_ = ~v13 & new_n3540_;
  assign new_n3542_ = v12 & new_n3541_;
  assign new_n3543_ = ~v11 & new_n3542_;
  assign new_n3544_ = ~v10 & new_n3543_;
  assign new_n3545_ = ~v9 & new_n3544_;
  assign new_n3546_ = ~v8 & new_n3545_;
  assign new_n3547_ = ~v5 & new_n3546_;
  assign new_n3548_ = ~v4 & new_n3547_;
  assign new_n3549_ = ~v3 & new_n3548_;
  assign new_n3550_ = ~v2 & new_n3549_;
  assign new_n3551_ = ~v1 & new_n3550_;
  assign \v41.40  = ~v0 & new_n3551_;
  assign new_n3553_ = v0 & new_n1257_;
  assign new_n3554_ = v17 & ~new_n975_;
  assign new_n3555_ = ~v18 & ~new_n3554_;
  assign new_n3556_ = ~new_n1039_ & ~new_n3555_;
  assign new_n3557_ = v40 & ~new_n3556_;
  assign new_n3558_ = ~v15 & new_n3557_;
  assign new_n3559_ = ~v3 & new_n3558_;
  assign new_n3560_ = ~v0 & new_n3559_;
  assign new_n3561_ = ~new_n3553_ & ~new_n3560_;
  assign new_n3562_ = v16 & ~new_n3561_;
  assign new_n3563_ = v3 & ~v19;
  assign new_n3564_ = ~v3 & v18;
  assign new_n3565_ = new_n1648_ & new_n3564_;
  assign new_n3566_ = ~new_n3563_ & ~new_n3565_;
  assign new_n3567_ = v17 & ~new_n3566_;
  assign new_n3568_ = ~v16 & new_n3567_;
  assign new_n3569_ = v15 & new_n3568_;
  assign new_n3570_ = ~v0 & new_n3569_;
  assign new_n3571_ = ~new_n3562_ & ~new_n3570_;
  assign new_n3572_ = ~v12 & ~new_n3571_;
  assign new_n3573_ = v25 & v26;
  assign new_n3574_ = new_n434_ & new_n3573_;
  assign new_n3575_ = ~v15 & ~new_n3574_;
  assign new_n3576_ = v40 & ~new_n3575_;
  assign new_n3577_ = v28 & new_n3576_;
  assign new_n3578_ = v12 & new_n3577_;
  assign new_n3579_ = ~v3 & new_n3578_;
  assign new_n3580_ = ~v0 & new_n3579_;
  assign new_n3581_ = ~new_n3572_ & ~new_n3580_;
  assign new_n3582_ = v13 & ~new_n3581_;
  assign new_n3583_ = ~new_n118_ & ~new_n1106_;
  assign new_n3584_ = v40 & new_n3583_;
  assign new_n3585_ = ~v3 & new_n3584_;
  assign new_n3586_ = ~v16 & new_n1038_;
  assign new_n3587_ = new_n494_ & new_n3586_;
  assign new_n3588_ = new_n723_ & new_n2948_;
  assign new_n3589_ = new_n3587_ & new_n3588_;
  assign new_n3590_ = ~new_n3585_ & ~new_n3589_;
  assign new_n3591_ = v17 & ~new_n3590_;
  assign new_n3592_ = ~v13 & new_n3591_;
  assign new_n3593_ = v12 & new_n3592_;
  assign new_n3594_ = ~v0 & new_n3593_;
  assign new_n3595_ = ~new_n3582_ & ~new_n3594_;
  assign new_n3596_ = ~v5 & ~new_n3595_;
  assign new_n3597_ = ~v26 & v27;
  assign new_n3598_ = new_n1512_ & new_n3597_;
  assign new_n3599_ = ~new_n1224_ & ~new_n3598_;
  assign new_n3600_ = v22 & ~new_n3599_;
  assign new_n3601_ = ~new_n1231_ & ~new_n3600_;
  assign new_n3602_ = v21 & ~new_n3601_;
  assign new_n3603_ = ~v20 & new_n3602_;
  assign new_n3604_ = ~new_n1239_ & ~new_n3603_;
  assign new_n3605_ = ~v19 & ~new_n3604_;
  assign new_n3606_ = v18 & new_n3605_;
  assign new_n3607_ = v17 & new_n3606_;
  assign new_n3608_ = ~v16 & new_n3607_;
  assign new_n3609_ = ~v15 & new_n3608_;
  assign new_n3610_ = ~v13 & new_n3609_;
  assign new_n3611_ = v12 & new_n3610_;
  assign new_n3612_ = v5 & new_n3611_;
  assign new_n3613_ = v3 & new_n3612_;
  assign new_n3614_ = ~v0 & new_n3613_;
  assign new_n3615_ = ~new_n3596_ & ~new_n3614_;
  assign new_n3616_ = ~v14 & ~new_n3615_;
  assign new_n3617_ = v16 & new_n579_;
  assign new_n3618_ = v15 & new_n3617_;
  assign new_n3619_ = v14 & new_n3618_;
  assign new_n3620_ = v13 & new_n3619_;
  assign new_n3621_ = v12 & new_n3620_;
  assign new_n3622_ = ~v5 & new_n3621_;
  assign new_n3623_ = ~v3 & new_n3622_;
  assign new_n3624_ = ~v0 & new_n3623_;
  assign new_n3625_ = ~new_n3616_ & ~new_n3624_;
  assign new_n3626_ = ~v2 & ~new_n3625_;
  assign new_n3627_ = ~v3 & new_n1289_;
  assign new_n3628_ = v2 & new_n3627_;
  assign new_n3629_ = ~v0 & new_n3628_;
  assign new_n3630_ = ~new_n3626_ & ~new_n3629_;
  assign new_n3631_ = ~v4 & ~new_n3630_;
  assign new_n3632_ = new_n735_ & new_n1258_;
  assign new_n3633_ = v17 & new_n2008_;
  assign new_n3634_ = new_n494_ & new_n3633_;
  assign new_n3635_ = new_n2275_ & new_n3634_;
  assign new_n3636_ = ~new_n3632_ & ~new_n3635_;
  assign new_n3637_ = v18 & ~new_n3636_;
  assign new_n3638_ = ~v16 & new_n3637_;
  assign new_n3639_ = ~v14 & new_n3638_;
  assign new_n3640_ = ~v13 & new_n3639_;
  assign new_n3641_ = v12 & new_n3640_;
  assign new_n3642_ = v5 & new_n3641_;
  assign new_n3643_ = v4 & new_n3642_;
  assign new_n3644_ = ~v2 & new_n3643_;
  assign new_n3645_ = ~v0 & new_n3644_;
  assign new_n3646_ = ~new_n3631_ & ~new_n3645_;
  assign new_n3647_ = ~v36 & ~new_n3646_;
  assign new_n3648_ = ~v11 & new_n3647_;
  assign new_n3649_ = ~v10 & new_n3648_;
  assign new_n3650_ = ~v9 & new_n3649_;
  assign new_n3651_ = ~v8 & new_n3650_;
  assign \v41.41  = ~v1 & new_n3651_;
  assign new_n3653_ = ~v5 & new_n1552_;
  assign new_n3654_ = ~v3 & new_n3653_;
  assign new_n3655_ = v2 & new_n3654_;
  assign new_n3656_ = ~v23 & ~v27;
  assign new_n3657_ = v22 & new_n3656_;
  assign new_n3658_ = new_n2878_ & new_n3657_;
  assign new_n3659_ = ~new_n3655_ & ~new_n3658_;
  assign new_n3660_ = ~v24 & ~new_n3659_;
  assign new_n3661_ = new_n680_ & new_n1222_;
  assign new_n3662_ = new_n2878_ & new_n3661_;
  assign new_n3663_ = ~new_n3660_ & ~new_n3662_;
  assign new_n3664_ = v21 & ~new_n3663_;
  assign new_n3665_ = ~v20 & new_n3664_;
  assign new_n3666_ = v2 & new_n351_;
  assign new_n3667_ = new_n2002_ & new_n3666_;
  assign new_n3668_ = ~new_n3665_ & ~new_n3667_;
  assign new_n3669_ = ~v15 & ~new_n3668_;
  assign new_n3670_ = v15 & v40;
  assign new_n3671_ = ~v5 & new_n3670_;
  assign new_n3672_ = new_n161_ & new_n3671_;
  assign new_n3673_ = ~new_n3669_ & ~new_n3672_;
  assign new_n3674_ = ~v19 & ~new_n3673_;
  assign new_n3675_ = v18 & new_n3674_;
  assign new_n3676_ = v15 & ~v18;
  assign new_n3677_ = new_n1648_ & new_n3676_;
  assign new_n3678_ = new_n2785_ & new_n3677_;
  assign new_n3679_ = ~new_n3675_ & ~new_n3678_;
  assign new_n3680_ = v17 & ~new_n3679_;
  assign new_n3681_ = new_n161_ & new_n257_;
  assign new_n3682_ = new_n753_ & new_n1595_;
  assign new_n3683_ = new_n3681_ & new_n3682_;
  assign new_n3684_ = ~new_n3680_ & ~new_n3683_;
  assign new_n3685_ = ~v16 & ~new_n3684_;
  assign new_n3686_ = new_n161_ & new_n207_;
  assign new_n3687_ = new_n673_ & new_n1649_;
  assign new_n3688_ = new_n3686_ & new_n3687_;
  assign new_n3689_ = ~new_n3685_ & ~new_n3688_;
  assign new_n3690_ = ~v13 & ~new_n3689_;
  assign new_n3691_ = v34 & v40;
  assign new_n3692_ = v33 & new_n3691_;
  assign new_n3693_ = v32 & new_n3692_;
  assign new_n3694_ = v30 & new_n3693_;
  assign new_n3695_ = v13 & new_n3694_;
  assign new_n3696_ = ~v5 & new_n3695_;
  assign new_n3697_ = ~v3 & new_n3696_;
  assign new_n3698_ = ~v2 & new_n3697_;
  assign new_n3699_ = ~new_n3690_ & ~new_n3698_;
  assign new_n3700_ = ~v14 & ~new_n3699_;
  assign new_n3701_ = new_n1902_ & new_n3670_;
  assign new_n3702_ = new_n2785_ & new_n3701_;
  assign new_n3703_ = ~new_n3700_ & ~new_n3702_;
  assign new_n3704_ = v12 & ~new_n3703_;
  assign new_n3705_ = new_n161_ & new_n2116_;
  assign new_n3706_ = new_n1338_ & new_n3670_;
  assign new_n3707_ = new_n3705_ & new_n3706_;
  assign new_n3708_ = ~new_n3704_ & ~new_n3707_;
  assign new_n3709_ = ~v4 & ~new_n3708_;
  assign new_n3710_ = new_n329_ & new_n360_;
  assign new_n3711_ = new_n2271_ & new_n3710_;
  assign new_n3712_ = new_n2276_ & new_n3711_;
  assign new_n3713_ = ~new_n3709_ & ~new_n3712_;
  assign new_n3714_ = ~v36 & ~new_n3713_;
  assign new_n3715_ = ~v11 & new_n3714_;
  assign new_n3716_ = ~v10 & new_n3715_;
  assign new_n3717_ = ~v9 & new_n3716_;
  assign new_n3718_ = ~v8 & new_n3717_;
  assign new_n3719_ = ~v1 & new_n3718_;
  assign \v41.42  = ~v0 & new_n3719_;
  assign new_n3721_ = ~new_n716_ & ~new_n1225_;
  assign new_n3722_ = v24 & ~new_n3721_;
  assign new_n3723_ = v23 & new_n3722_;
  assign new_n3724_ = v22 & new_n3723_;
  assign new_n3725_ = v21 & new_n3724_;
  assign new_n3726_ = ~v20 & new_n3725_;
  assign new_n3727_ = ~v14 & new_n3726_;
  assign new_n3728_ = v12 & new_n3727_;
  assign new_n3729_ = v3 & new_n3728_;
  assign new_n3730_ = ~v3 & ~v12;
  assign new_n3731_ = new_n333_ & new_n3730_;
  assign new_n3732_ = ~new_n3729_ & ~new_n3731_;
  assign new_n3733_ = ~v19 & ~new_n3732_;
  assign new_n3734_ = v14 & new_n1648_;
  assign new_n3735_ = new_n3730_ & new_n3734_;
  assign new_n3736_ = ~new_n3733_ & ~new_n3735_;
  assign new_n3737_ = ~v15 & ~new_n3736_;
  assign new_n3738_ = ~v3 & new_n3033_;
  assign new_n3739_ = ~new_n3737_ & ~new_n3738_;
  assign new_n3740_ = ~v16 & ~new_n3739_;
  assign new_n3741_ = ~v3 & new_n3039_;
  assign new_n3742_ = ~new_n3740_ & ~new_n3741_;
  assign new_n3743_ = v18 & ~new_n3742_;
  assign new_n3744_ = ~v18 & new_n3043_;
  assign new_n3745_ = ~v3 & new_n3744_;
  assign new_n3746_ = ~new_n3743_ & ~new_n3745_;
  assign new_n3747_ = v17 & ~new_n3746_;
  assign new_n3748_ = ~v17 & new_n3049_;
  assign new_n3749_ = ~v3 & new_n3748_;
  assign new_n3750_ = ~new_n3747_ & ~new_n3749_;
  assign new_n3751_ = ~v13 & ~new_n3750_;
  assign new_n3752_ = v40 & ~new_n2177_;
  assign new_n3753_ = v14 & new_n3752_;
  assign new_n3754_ = v13 & new_n3753_;
  assign new_n3755_ = v12 & new_n3754_;
  assign new_n3756_ = ~v3 & new_n3755_;
  assign new_n3757_ = ~new_n3751_ & ~new_n3756_;
  assign new_n3758_ = v5 & ~new_n3757_;
  assign new_n3759_ = ~v16 & ~new_n1106_;
  assign new_n3760_ = v14 & new_n3759_;
  assign new_n3761_ = v13 & new_n3760_;
  assign new_n3762_ = v16 & new_n860_;
  assign new_n3763_ = ~v14 & new_n3762_;
  assign new_n3764_ = ~v13 & new_n3763_;
  assign new_n3765_ = ~new_n3761_ & ~new_n3764_;
  assign new_n3766_ = v17 & ~new_n3765_;
  assign new_n3767_ = ~v14 & new_n1350_;
  assign new_n3768_ = ~v14 & ~new_n3767_;
  assign new_n3769_ = ~v13 & ~new_n3768_;
  assign new_n3770_ = ~v14 & v20;
  assign new_n3771_ = v13 & new_n3770_;
  assign new_n3772_ = new_n2273_ & new_n2524_;
  assign new_n3773_ = new_n3771_ & new_n3772_;
  assign new_n3774_ = ~new_n3769_ & ~new_n3773_;
  assign new_n3775_ = ~new_n3766_ & new_n3774_;
  assign new_n3776_ = v12 & ~new_n3775_;
  assign new_n3777_ = v14 & ~new_n2902_;
  assign new_n3778_ = new_n120_ & new_n164_;
  assign new_n3779_ = v16 & ~new_n3778_;
  assign new_n3780_ = ~v14 & ~new_n3779_;
  assign new_n3781_ = v13 & new_n3780_;
  assign new_n3782_ = ~new_n3777_ & ~new_n3781_;
  assign new_n3783_ = ~v12 & ~new_n3782_;
  assign new_n3784_ = ~new_n3776_ & ~new_n3783_;
  assign new_n3785_ = ~v15 & ~new_n3784_;
  assign new_n3786_ = new_n265_ & new_n1356_;
  assign new_n3787_ = new_n260_ & new_n3786_;
  assign new_n3788_ = ~new_n3785_ & ~new_n3787_;
  assign new_n3789_ = v40 & ~new_n3788_;
  assign new_n3790_ = ~v3 & new_n3789_;
  assign new_n3791_ = v3 & v12;
  assign new_n3792_ = new_n1343_ & new_n3791_;
  assign new_n3793_ = new_n268_ & new_n3792_;
  assign new_n3794_ = ~new_n3790_ & ~new_n3793_;
  assign new_n3795_ = ~v5 & ~new_n3794_;
  assign new_n3796_ = ~new_n3758_ & ~new_n3795_;
  assign new_n3797_ = ~v0 & ~new_n3796_;
  assign new_n3798_ = new_n266_ & new_n498_;
  assign new_n3799_ = new_n1013_ & new_n3798_;
  assign new_n3800_ = ~new_n3797_ & ~new_n3799_;
  assign new_n3801_ = ~v36 & ~new_n3800_;
  assign new_n3802_ = ~v11 & new_n3801_;
  assign new_n3803_ = ~v10 & new_n3802_;
  assign new_n3804_ = ~v9 & new_n3803_;
  assign new_n3805_ = ~v8 & new_n3804_;
  assign new_n3806_ = ~v4 & new_n3805_;
  assign new_n3807_ = ~v2 & new_n3806_;
  assign \v41.43  = ~v1 & new_n3807_;
  assign new_n3809_ = ~new_n421_ & ~new_n727_;
  assign new_n3810_ = new_n681_ & ~new_n2215_;
  assign new_n3811_ = v27 & ~new_n3810_;
  assign new_n3812_ = ~v27 & ~new_n681_;
  assign new_n3813_ = ~v24 & new_n3812_;
  assign new_n3814_ = ~new_n3811_ & ~new_n3813_;
  assign new_n3815_ = v40 & ~new_n3814_;
  assign new_n3816_ = ~v3 & new_n3815_;
  assign new_n3817_ = ~new_n3809_ & ~new_n3816_;
  assign new_n3818_ = ~v5 & ~new_n3817_;
  assign new_n3819_ = v27 & ~new_n687_;
  assign new_n3820_ = v23 & new_n3819_;
  assign new_n3821_ = v22 & new_n3820_;
  assign new_n3822_ = ~new_n3111_ & ~new_n3821_;
  assign new_n3823_ = v3 & new_n3723_;
  assign new_n3824_ = ~v3 & ~v23;
  assign new_n3825_ = new_n1541_ & new_n3824_;
  assign new_n3826_ = ~new_n3823_ & ~new_n3825_;
  assign new_n3827_ = v22 & ~new_n3826_;
  assign new_n3828_ = ~v3 & ~v22;
  assign new_n3829_ = new_n1541_ & new_n3828_;
  assign new_n3830_ = ~new_n3827_ & ~new_n3829_;
  assign new_n3831_ = new_n3822_ & new_n3830_;
  assign new_n3832_ = v5 & ~new_n3831_;
  assign new_n3833_ = ~new_n3818_ & ~new_n3832_;
  assign new_n3834_ = ~v4 & ~new_n3833_;
  assign new_n3835_ = v3 & ~new_n2657_;
  assign new_n3836_ = ~new_n681_ & ~new_n3835_;
  assign new_n3837_ = v22 & v23;
  assign new_n3838_ = v3 & ~v5;
  assign new_n3839_ = new_n3837_ & new_n3838_;
  assign new_n3840_ = ~new_n3836_ & ~new_n3839_;
  assign new_n3841_ = ~v24 & ~new_n3840_;
  assign new_n3842_ = new_n692_ & new_n3838_;
  assign new_n3843_ = ~new_n3841_ & ~new_n3842_;
  assign new_n3844_ = v27 & ~new_n3843_;
  assign new_n3845_ = v4 & new_n3844_;
  assign new_n3846_ = ~new_n3834_ & ~new_n3845_;
  assign new_n3847_ = ~v20 & ~new_n3846_;
  assign new_n3848_ = v20 & v40;
  assign new_n3849_ = ~v5 & new_n3848_;
  assign new_n3850_ = new_n256_ & new_n3849_;
  assign new_n3851_ = ~new_n3847_ & ~new_n3850_;
  assign new_n3852_ = v21 & ~new_n3851_;
  assign new_n3853_ = v27 & ~new_n1398_;
  assign new_n3854_ = ~v27 & ~new_n672_;
  assign new_n3855_ = ~v4 & new_n3854_;
  assign new_n3856_ = ~new_n3853_ & ~new_n3855_;
  assign new_n3857_ = ~v3 & ~new_n3856_;
  assign new_n3858_ = v5 & ~v27;
  assign new_n3859_ = new_n1483_ & new_n3858_;
  assign new_n3860_ = ~new_n3857_ & ~new_n3859_;
  assign new_n3861_ = ~v21 & ~new_n3860_;
  assign new_n3862_ = v20 & new_n3861_;
  assign new_n3863_ = ~new_n3852_ & ~new_n3862_;
  assign new_n3864_ = ~v2 & ~new_n3863_;
  assign new_n3865_ = ~new_n679_ & ~new_n1278_;
  assign new_n3866_ = v27 & ~new_n3865_;
  assign new_n3867_ = ~v4 & new_n3866_;
  assign new_n3868_ = ~v3 & new_n3867_;
  assign new_n3869_ = v2 & new_n3868_;
  assign new_n3870_ = ~new_n3864_ & ~new_n3869_;
  assign new_n3871_ = ~v36 & ~new_n3870_;
  assign new_n3872_ = ~v19 & new_n3871_;
  assign new_n3873_ = v18 & new_n3872_;
  assign new_n3874_ = v17 & new_n3873_;
  assign new_n3875_ = ~v16 & new_n3874_;
  assign new_n3876_ = ~v15 & new_n3875_;
  assign new_n3877_ = ~v14 & new_n3876_;
  assign new_n3878_ = ~v13 & new_n3877_;
  assign new_n3879_ = v12 & new_n3878_;
  assign new_n3880_ = ~v11 & new_n3879_;
  assign new_n3881_ = ~v10 & new_n3880_;
  assign new_n3882_ = ~v9 & new_n3881_;
  assign new_n3883_ = ~v8 & new_n3882_;
  assign new_n3884_ = ~v1 & new_n3883_;
  assign \v41.44  = ~v0 & new_n3884_;
  assign new_n3886_ = new_n685_ & ~new_n1133_;
  assign new_n3887_ = ~v19 & ~new_n3886_;
  assign new_n3888_ = ~v19 & ~new_n3887_;
  assign new_n3889_ = ~v16 & ~new_n3888_;
  assign new_n3890_ = ~v16 & ~new_n3889_;
  assign new_n3891_ = v40 & ~new_n3890_;
  assign new_n3892_ = ~v5 & new_n3891_;
  assign new_n3893_ = ~v16 & new_n775_;
  assign new_n3894_ = v5 & new_n3893_;
  assign new_n3895_ = ~new_n3892_ & ~new_n3894_;
  assign new_n3896_ = ~v15 & ~new_n3895_;
  assign new_n3897_ = ~new_n3671_ & ~new_n3896_;
  assign new_n3898_ = ~v14 & ~new_n3897_;
  assign new_n3899_ = ~v13 & new_n3898_;
  assign new_n3900_ = v13 & new_n333_;
  assign new_n3901_ = ~v5 & new_n3900_;
  assign new_n3902_ = ~new_n3899_ & ~new_n3901_;
  assign new_n3903_ = v18 & ~new_n3902_;
  assign new_n3904_ = v13 & new_n2325_;
  assign new_n3905_ = ~new_n1343_ & ~new_n3904_;
  assign new_n3906_ = ~new_n402_ & ~new_n3905_;
  assign new_n3907_ = ~new_n1338_ & ~new_n1357_;
  assign new_n3908_ = ~new_n156_ & ~new_n3907_;
  assign new_n3909_ = new_n1338_ & new_n1589_;
  assign new_n3910_ = ~new_n3908_ & ~new_n3909_;
  assign new_n3911_ = ~new_n3906_ & new_n3910_;
  assign new_n3912_ = v40 & ~new_n3911_;
  assign new_n3913_ = ~v18 & new_n3912_;
  assign new_n3914_ = ~v5 & new_n3913_;
  assign new_n3915_ = ~new_n3903_ & ~new_n3914_;
  assign new_n3916_ = v17 & ~new_n3915_;
  assign new_n3917_ = ~v16 & new_n171_;
  assign new_n3918_ = ~new_n1604_ & ~new_n3917_;
  assign new_n3919_ = ~new_n1338_ & ~new_n2283_;
  assign new_n3920_ = ~new_n3918_ & ~new_n3919_;
  assign new_n3921_ = ~v15 & new_n165_;
  assign new_n3922_ = ~new_n1879_ & ~new_n3921_;
  assign new_n3923_ = v14 & ~new_n3922_;
  assign new_n3924_ = v13 & new_n3923_;
  assign new_n3925_ = new_n1343_ & new_n2545_;
  assign new_n3926_ = ~new_n3924_ & ~new_n3925_;
  assign new_n3927_ = ~new_n1349_ & ~new_n1357_;
  assign new_n3928_ = new_n1338_ & new_n3676_;
  assign new_n3929_ = new_n3927_ & ~new_n3928_;
  assign new_n3930_ = ~v19 & ~new_n3929_;
  assign new_n3931_ = v15 & new_n120_;
  assign new_n3932_ = new_n1343_ & new_n3931_;
  assign new_n3933_ = ~new_n3930_ & ~new_n3932_;
  assign new_n3934_ = v16 & ~new_n3933_;
  assign new_n3935_ = new_n3050_ & new_n3904_;
  assign new_n3936_ = ~new_n3934_ & ~new_n3935_;
  assign new_n3937_ = new_n3926_ & new_n3936_;
  assign new_n3938_ = ~new_n3920_ & new_n3937_;
  assign new_n3939_ = ~v17 & ~new_n3938_;
  assign new_n3940_ = ~new_n1902_ & ~new_n3939_;
  assign new_n3941_ = v40 & ~new_n3940_;
  assign new_n3942_ = ~v5 & new_n3941_;
  assign new_n3943_ = ~new_n3916_ & ~new_n3942_;
  assign new_n3944_ = v12 & ~new_n3943_;
  assign new_n3945_ = new_n201_ & new_n1713_;
  assign new_n3946_ = new_n1332_ & ~new_n3945_;
  assign new_n3947_ = v40 & ~new_n3946_;
  assign new_n3948_ = v14 & new_n3947_;
  assign new_n3949_ = ~v13 & new_n3948_;
  assign new_n3950_ = ~v12 & new_n3949_;
  assign new_n3951_ = ~v5 & new_n3950_;
  assign new_n3952_ = ~new_n3944_ & ~new_n3951_;
  assign new_n3953_ = ~v3 & ~new_n3952_;
  assign new_n3954_ = v12 & new_n1343_;
  assign new_n3955_ = new_n3838_ & new_n3954_;
  assign new_n3956_ = new_n268_ & new_n3955_;
  assign new_n3957_ = ~new_n3953_ & ~new_n3956_;
  assign new_n3958_ = ~v0 & ~new_n3957_;
  assign new_n3959_ = ~new_n3799_ & ~new_n3958_;
  assign new_n3960_ = ~v36 & ~new_n3959_;
  assign new_n3961_ = ~v11 & new_n3960_;
  assign new_n3962_ = ~v10 & new_n3961_;
  assign new_n3963_ = ~v9 & new_n3962_;
  assign new_n3964_ = ~v8 & new_n3963_;
  assign new_n3965_ = ~v4 & new_n3964_;
  assign new_n3966_ = ~v2 & new_n3965_;
  assign \v41.45  = ~v1 & new_n3966_;
  assign new_n3968_ = new_n1134_ & new_n1810_;
  assign new_n3969_ = ~new_n1813_ & ~new_n3968_;
  assign new_n3970_ = v40 & ~new_n3969_;
  assign new_n3971_ = ~v3 & new_n3970_;
  assign new_n3972_ = ~v19 & new_n729_;
  assign new_n3973_ = ~v14 & new_n3972_;
  assign new_n3974_ = v12 & new_n3973_;
  assign new_n3975_ = v3 & new_n3974_;
  assign new_n3976_ = ~new_n3971_ & ~new_n3975_;
  assign new_n3977_ = ~v5 & ~new_n3976_;
  assign new_n3978_ = ~v14 & new_n3116_;
  assign new_n3979_ = v12 & new_n3978_;
  assign new_n3980_ = v5 & new_n3979_;
  assign new_n3981_ = v3 & new_n3980_;
  assign new_n3982_ = ~new_n3977_ & ~new_n3981_;
  assign new_n3983_ = ~v2 & ~new_n3982_;
  assign new_n3984_ = ~v19 & new_n3866_;
  assign new_n3985_ = ~v14 & new_n3984_;
  assign new_n3986_ = v12 & new_n3985_;
  assign new_n3987_ = ~v3 & new_n3986_;
  assign new_n3988_ = v2 & new_n3987_;
  assign new_n3989_ = ~new_n3983_ & ~new_n3988_;
  assign new_n3990_ = ~v15 & ~new_n3989_;
  assign new_n3991_ = ~v5 & new_n3033_;
  assign new_n3992_ = ~v3 & new_n3991_;
  assign new_n3993_ = ~v2 & new_n3992_;
  assign new_n3994_ = ~new_n3990_ & ~new_n3993_;
  assign new_n3995_ = ~v16 & ~new_n3994_;
  assign new_n3996_ = ~v5 & new_n3039_;
  assign new_n3997_ = ~v3 & new_n3996_;
  assign new_n3998_ = ~v2 & new_n3997_;
  assign new_n3999_ = ~new_n3995_ & ~new_n3998_;
  assign new_n4000_ = v18 & ~new_n3999_;
  assign new_n4001_ = ~v5 & new_n3744_;
  assign new_n4002_ = ~v3 & new_n4001_;
  assign new_n4003_ = ~v2 & new_n4002_;
  assign new_n4004_ = ~new_n4000_ & ~new_n4003_;
  assign new_n4005_ = v17 & ~new_n4004_;
  assign new_n4006_ = ~v12 & new_n900_;
  assign new_n4007_ = new_n3050_ & new_n4006_;
  assign new_n4008_ = new_n1812_ & ~new_n4007_;
  assign new_n4009_ = v40 & ~new_n4008_;
  assign new_n4010_ = ~v17 & new_n4009_;
  assign new_n4011_ = ~v5 & new_n4010_;
  assign new_n4012_ = ~v3 & new_n4011_;
  assign new_n4013_ = ~v2 & new_n4012_;
  assign new_n4014_ = ~new_n4005_ & ~new_n4013_;
  assign new_n4015_ = ~v13 & ~new_n4014_;
  assign new_n4016_ = ~v15 & new_n2846_;
  assign new_n4017_ = new_n2578_ & ~new_n4016_;
  assign new_n4018_ = ~new_n1190_ & new_n4017_;
  assign new_n4019_ = v40 & ~new_n4018_;
  assign new_n4020_ = v14 & new_n4019_;
  assign new_n4021_ = v13 & new_n4020_;
  assign new_n4022_ = v12 & new_n4021_;
  assign new_n4023_ = ~v5 & new_n4022_;
  assign new_n4024_ = ~v3 & new_n4023_;
  assign new_n4025_ = ~v2 & new_n4024_;
  assign new_n4026_ = ~new_n4015_ & ~new_n4025_;
  assign new_n4027_ = ~v4 & ~new_n4026_;
  assign new_n4028_ = v5 & ~new_n681_;
  assign new_n4029_ = ~v5 & new_n3837_;
  assign new_n4030_ = ~new_n4028_ & ~new_n4029_;
  assign new_n4031_ = ~v24 & ~new_n4030_;
  assign new_n4032_ = ~v5 & new_n692_;
  assign new_n4033_ = ~new_n4031_ & ~new_n4032_;
  assign new_n4034_ = v27 & ~new_n4033_;
  assign new_n4035_ = v21 & new_n4034_;
  assign new_n4036_ = ~v20 & new_n4035_;
  assign new_n4037_ = ~v19 & new_n4036_;
  assign new_n4038_ = v18 & new_n4037_;
  assign new_n4039_ = v17 & new_n4038_;
  assign new_n4040_ = ~v16 & new_n4039_;
  assign new_n4041_ = ~v15 & new_n4040_;
  assign new_n4042_ = ~v14 & new_n4041_;
  assign new_n4043_ = ~v13 & new_n4042_;
  assign new_n4044_ = v12 & new_n4043_;
  assign new_n4045_ = v4 & new_n4044_;
  assign new_n4046_ = v3 & new_n4045_;
  assign new_n4047_ = ~v2 & new_n4046_;
  assign new_n4048_ = ~new_n4027_ & ~new_n4047_;
  assign new_n4049_ = ~v36 & ~new_n4048_;
  assign new_n4050_ = ~v11 & new_n4049_;
  assign new_n4051_ = ~v10 & new_n4050_;
  assign new_n4052_ = ~v9 & new_n4051_;
  assign new_n4053_ = ~v8 & new_n4052_;
  assign new_n4054_ = ~v1 & new_n4053_;
  assign \v41.46  = ~v0 & new_n4054_;
  assign new_n4056_ = ~new_n1279_ & ~new_n2249_;
  assign new_n4057_ = v2 & ~new_n4056_;
  assign new_n4058_ = v21 & ~new_n3810_;
  assign new_n4059_ = ~v20 & new_n4058_;
  assign new_n4060_ = ~new_n679_ & ~new_n4059_;
  assign new_n4061_ = v40 & ~new_n4060_;
  assign new_n4062_ = ~v5 & new_n4061_;
  assign new_n4063_ = ~v2 & new_n4062_;
  assign new_n4064_ = ~new_n4057_ & ~new_n4063_;
  assign new_n4065_ = v27 & ~new_n4064_;
  assign new_n4066_ = ~v2 & ~v5;
  assign new_n4067_ = v21 & v40;
  assign new_n4068_ = v20 & new_n4067_;
  assign new_n4069_ = new_n4066_ & new_n4068_;
  assign new_n4070_ = ~new_n4065_ & ~new_n4069_;
  assign new_n4071_ = v18 & ~new_n4070_;
  assign new_n4072_ = ~v16 & new_n4071_;
  assign new_n4073_ = v40 & ~new_n740_;
  assign new_n4074_ = ~v18 & new_n4073_;
  assign new_n4075_ = v16 & new_n4074_;
  assign new_n4076_ = ~v5 & new_n4075_;
  assign new_n4077_ = ~v2 & new_n4076_;
  assign new_n4078_ = ~new_n4072_ & ~new_n4077_;
  assign new_n4079_ = ~v14 & ~new_n4078_;
  assign new_n4080_ = v12 & new_n4079_;
  assign new_n4081_ = ~v5 & new_n3024_;
  assign new_n4082_ = ~v2 & new_n4081_;
  assign new_n4083_ = ~new_n4080_ & ~new_n4082_;
  assign new_n4084_ = ~v15 & ~new_n4083_;
  assign new_n4085_ = v12 & new_n1339_;
  assign new_n4086_ = ~new_n1813_ & ~new_n4085_;
  assign new_n4087_ = v40 & ~new_n4086_;
  assign new_n4088_ = v15 & new_n4087_;
  assign new_n4089_ = ~v5 & new_n4088_;
  assign new_n4090_ = ~v2 & new_n4089_;
  assign new_n4091_ = ~new_n4084_ & ~new_n4090_;
  assign new_n4092_ = ~v19 & ~new_n4091_;
  assign new_n4093_ = new_n490_ & new_n1810_;
  assign new_n4094_ = new_n3042_ & ~new_n4093_;
  assign new_n4095_ = v40 & ~new_n4094_;
  assign new_n4096_ = v19 & new_n4095_;
  assign new_n4097_ = ~v5 & new_n4096_;
  assign new_n4098_ = ~v2 & new_n4097_;
  assign new_n4099_ = ~new_n4092_ & ~new_n4098_;
  assign new_n4100_ = v17 & ~new_n4099_;
  assign new_n4101_ = new_n1813_ & new_n3403_;
  assign new_n4102_ = new_n1810_ & new_n3676_;
  assign new_n4103_ = ~v19 & ~v37;
  assign new_n4104_ = new_n843_ & new_n4103_;
  assign new_n4105_ = new_n4102_ & new_n4104_;
  assign new_n4106_ = ~new_n4101_ & ~new_n4105_;
  assign new_n4107_ = ~v16 & ~new_n4106_;
  assign new_n4108_ = new_n1812_ & ~new_n4107_;
  assign new_n4109_ = v40 & ~new_n4108_;
  assign new_n4110_ = ~v17 & new_n4109_;
  assign new_n4111_ = ~v5 & new_n4110_;
  assign new_n4112_ = ~v2 & new_n4111_;
  assign new_n4113_ = ~new_n4100_ & ~new_n4112_;
  assign new_n4114_ = ~v13 & ~new_n4113_;
  assign new_n4115_ = ~new_n674_ & ~new_n1868_;
  assign new_n4116_ = ~new_n1823_ & new_n4115_;
  assign new_n4117_ = v14 & ~new_n4116_;
  assign new_n4118_ = v12 & new_n4117_;
  assign new_n4119_ = new_n117_ & new_n952_;
  assign new_n4120_ = new_n753_ & new_n844_;
  assign new_n4121_ = new_n4119_ & new_n4120_;
  assign new_n4122_ = ~new_n4118_ & ~new_n4121_;
  assign new_n4123_ = new_n166_ & new_n3057_;
  assign new_n4124_ = new_n4122_ & ~new_n4123_;
  assign new_n4125_ = v40 & ~new_n4124_;
  assign new_n4126_ = v13 & new_n4125_;
  assign new_n4127_ = ~v5 & new_n4126_;
  assign new_n4128_ = ~v2 & new_n4127_;
  assign new_n4129_ = ~new_n4114_ & ~new_n4128_;
  assign new_n4130_ = ~v4 & ~new_n4129_;
  assign new_n4131_ = ~v2 & new_n1026_;
  assign new_n4132_ = ~new_n4130_ & ~new_n4131_;
  assign new_n4133_ = ~v3 & ~new_n4132_;
  assign new_n4134_ = v4 & new_n1975_;
  assign new_n4135_ = v5 & v22;
  assign new_n4136_ = ~v4 & new_n4135_;
  assign new_n4137_ = v24 & v26;
  assign new_n4138_ = v23 & new_n4137_;
  assign new_n4139_ = new_n4136_ & new_n4138_;
  assign new_n4140_ = ~new_n4134_ & ~new_n4139_;
  assign new_n4141_ = v27 & ~new_n4140_;
  assign new_n4142_ = new_n1225_ & new_n1512_;
  assign new_n4143_ = new_n4136_ & new_n4142_;
  assign new_n4144_ = ~new_n4141_ & ~new_n4143_;
  assign new_n4145_ = v21 & ~new_n4144_;
  assign new_n4146_ = ~v20 & new_n4145_;
  assign new_n4147_ = ~v19 & new_n4146_;
  assign new_n4148_ = v18 & new_n4147_;
  assign new_n4149_ = v17 & new_n4148_;
  assign new_n4150_ = ~v16 & new_n4149_;
  assign new_n4151_ = ~v15 & new_n4150_;
  assign new_n4152_ = ~v14 & new_n4151_;
  assign new_n4153_ = ~v13 & new_n4152_;
  assign new_n4154_ = v12 & new_n4153_;
  assign new_n4155_ = v3 & new_n4154_;
  assign new_n4156_ = ~v2 & new_n4155_;
  assign new_n4157_ = ~new_n4133_ & ~new_n4156_;
  assign new_n4158_ = ~v36 & ~new_n4157_;
  assign new_n4159_ = ~v9 & new_n4158_;
  assign new_n4160_ = ~v1 & new_n4159_;
  assign new_n4161_ = ~v0 & new_n4160_;
  assign new_n4162_ = ~v9 & ~new_n4161_;
  assign new_n4163_ = ~v11 & ~new_n4162_;
  assign new_n4164_ = v9 & v11;
  assign new_n4165_ = ~new_n4163_ & ~new_n4164_;
  assign new_n4166_ = ~v10 & ~new_n4165_;
  assign new_n4167_ = ~new_n1392_ & ~new_n4166_;
  assign \v41.47  = ~v8 & ~new_n4167_;
  assign new_n4169_ = ~new_n2283_ & ~new_n3904_;
  assign new_n4170_ = v12 & ~new_n4169_;
  assign new_n4171_ = new_n1472_ & new_n2325_;
  assign new_n4172_ = ~new_n4170_ & ~new_n4171_;
  assign new_n4173_ = new_n1145_ & new_n1343_;
  assign new_n4174_ = new_n1146_ & new_n1338_;
  assign new_n4175_ = ~new_n4173_ & ~new_n4174_;
  assign new_n4176_ = v12 & ~new_n4175_;
  assign new_n4177_ = v14 & new_n226_;
  assign new_n4178_ = new_n1472_ & new_n4177_;
  assign new_n4179_ = ~new_n4176_ & ~new_n4178_;
  assign new_n4180_ = new_n4172_ & new_n4179_;
  assign new_n4181_ = ~new_n3918_ & ~new_n4180_;
  assign new_n4182_ = v12 & ~new_n2319_;
  assign new_n4183_ = ~v12 & new_n1902_;
  assign new_n4184_ = ~new_n4182_ & ~new_n4183_;
  assign new_n4185_ = v17 & ~new_n4184_;
  assign new_n4186_ = v14 & new_n753_;
  assign new_n4187_ = new_n1472_ & new_n4186_;
  assign new_n4188_ = ~new_n4185_ & ~new_n4187_;
  assign new_n4189_ = v13 & new_n948_;
  assign new_n4190_ = ~v14 & ~v18;
  assign new_n4191_ = ~v13 & new_n4190_;
  assign new_n4192_ = ~new_n4189_ & ~new_n4191_;
  assign new_n4193_ = new_n119_ & new_n1338_;
  assign new_n4194_ = new_n4192_ & ~new_n4193_;
  assign new_n4195_ = v12 & ~new_n4194_;
  assign new_n4196_ = v14 & new_n119_;
  assign new_n4197_ = new_n1472_ & new_n4196_;
  assign new_n4198_ = ~new_n4195_ & ~new_n4197_;
  assign new_n4199_ = v15 & ~new_n4198_;
  assign new_n4200_ = new_n4188_ & ~new_n4199_;
  assign new_n4201_ = ~new_n156_ & ~new_n4200_;
  assign new_n4202_ = v16 & new_n165_;
  assign new_n4203_ = new_n209_ & new_n1038_;
  assign new_n4204_ = ~new_n4202_ & ~new_n4203_;
  assign new_n4205_ = v13 & ~new_n4204_;
  assign new_n4206_ = v13 & ~new_n4205_;
  assign new_n4207_ = ~v16 & new_n165_;
  assign new_n4208_ = v16 & new_n1038_;
  assign new_n4209_ = ~new_n4207_ & ~new_n4208_;
  assign new_n4210_ = ~v15 & ~new_n4209_;
  assign new_n4211_ = ~new_n3072_ & ~new_n4210_;
  assign new_n4212_ = ~v17 & ~new_n4211_;
  assign new_n4213_ = v16 & new_n517_;
  assign new_n4214_ = ~v15 & new_n4213_;
  assign new_n4215_ = ~new_n4212_ & ~new_n4214_;
  assign new_n4216_ = v13 & ~new_n4215_;
  assign new_n4217_ = new_n4206_ & ~new_n4216_;
  assign new_n4218_ = v14 & ~new_n4217_;
  assign new_n4219_ = ~new_n230_ & ~new_n1189_;
  assign new_n4220_ = v15 & ~new_n4219_;
  assign new_n4221_ = ~v18 & ~new_n1161_;
  assign new_n4222_ = v17 & new_n4221_;
  assign new_n4223_ = ~v15 & new_n4222_;
  assign new_n4224_ = ~new_n4220_ & ~new_n4223_;
  assign new_n4225_ = v16 & ~new_n4224_;
  assign new_n4226_ = new_n117_ & new_n1911_;
  assign new_n4227_ = ~new_n4225_ & ~new_n4226_;
  assign new_n4228_ = ~v14 & ~new_n4227_;
  assign new_n4229_ = ~v13 & new_n4228_;
  assign new_n4230_ = ~new_n4218_ & ~new_n4229_;
  assign new_n4231_ = v12 & ~new_n4230_;
  assign new_n4232_ = ~new_n3586_ & ~new_n4202_;
  assign new_n4233_ = v15 & ~new_n4232_;
  assign new_n4234_ = new_n116_ & new_n165_;
  assign new_n4235_ = ~new_n4233_ & ~new_n4234_;
  assign new_n4236_ = ~v17 & ~new_n1866_;
  assign new_n4237_ = v16 & new_n4236_;
  assign new_n4238_ = ~new_n4203_ & ~new_n4237_;
  assign new_n4239_ = ~v15 & ~new_n4238_;
  assign new_n4240_ = new_n4235_ & ~new_n4239_;
  assign new_n4241_ = v14 & ~new_n4240_;
  assign new_n4242_ = ~v13 & new_n4241_;
  assign new_n4243_ = ~v12 & new_n4242_;
  assign new_n4244_ = ~new_n4231_ & ~new_n4243_;
  assign new_n4245_ = ~new_n4201_ & new_n4244_;
  assign new_n4246_ = ~new_n4181_ & new_n4245_;
  assign new_n4247_ = v40 & ~new_n4246_;
  assign new_n4248_ = ~v3 & new_n4247_;
  assign new_n4249_ = ~new_n3793_ & ~new_n4248_;
  assign new_n4250_ = ~v0 & ~new_n4249_;
  assign new_n4251_ = new_n498_ & new_n3954_;
  assign new_n4252_ = new_n268_ & new_n4251_;
  assign new_n4253_ = ~new_n4250_ & ~new_n4252_;
  assign new_n4254_ = ~v36 & ~new_n4253_;
  assign new_n4255_ = ~v11 & new_n4254_;
  assign new_n4256_ = ~v10 & new_n4255_;
  assign new_n4257_ = ~v9 & new_n4256_;
  assign new_n4258_ = ~v8 & new_n4257_;
  assign new_n4259_ = ~v5 & new_n4258_;
  assign new_n4260_ = ~v4 & new_n4259_;
  assign new_n4261_ = ~v2 & new_n4260_;
  assign \v41.48  = ~v1 & new_n4261_;
  assign new_n4263_ = ~v1 & ~new_n392_;
  assign new_n4264_ = new_n256_ & new_n1442_;
  assign new_n4265_ = ~new_n4263_ & ~new_n4264_;
  assign new_n4266_ = ~v3 & new_n1397_;
  assign new_n4267_ = ~v2 & new_n4266_;
  assign new_n4268_ = ~v1 & new_n4267_;
  assign new_n4269_ = new_n4265_ & ~new_n4268_;
  assign new_n4270_ = v1 & new_n161_;
  assign new_n4271_ = ~v5 & v16;
  assign new_n4272_ = v4 & new_n4271_;
  assign new_n4273_ = new_n4270_ & new_n4272_;
  assign new_n4274_ = new_n4269_ & ~new_n4273_;
  assign new_n4275_ = ~new_n156_ & ~new_n362_;
  assign new_n4276_ = ~v5 & new_n154_;
  assign new_n4277_ = new_n391_ & new_n4276_;
  assign new_n4278_ = ~new_n4275_ & ~new_n4277_;
  assign new_n4279_ = v1 & ~new_n4278_;
  assign new_n4280_ = new_n4274_ & ~new_n4279_;
  assign new_n4281_ = ~v18 & ~new_n4280_;
  assign new_n4282_ = ~v17 & new_n4281_;
  assign new_n4283_ = v15 & new_n4282_;
  assign new_n4284_ = new_n380_ & new_n390_;
  assign new_n4285_ = new_n455_ & ~new_n4284_;
  assign new_n4286_ = ~new_n4268_ & new_n4285_;
  assign new_n4287_ = v19 & ~new_n4286_;
  assign new_n4288_ = v18 & new_n4287_;
  assign new_n4289_ = v17 & new_n4288_;
  assign new_n4290_ = v16 & new_n4289_;
  assign new_n4291_ = ~v15 & new_n4290_;
  assign new_n4292_ = ~new_n4283_ & ~new_n4291_;
  assign new_n4293_ = ~v0 & ~new_n4292_;
  assign new_n4294_ = ~v3 & ~new_n1662_;
  assign new_n4295_ = ~v2 & new_n4294_;
  assign new_n4296_ = ~v1 & new_n4295_;
  assign new_n4297_ = v0 & new_n4296_;
  assign new_n4298_ = ~new_n4293_ & ~new_n4297_;
  assign new_n4299_ = ~v36 & ~new_n4298_;
  assign new_n4300_ = ~v14 & new_n4299_;
  assign new_n4301_ = v13 & new_n4300_;
  assign new_n4302_ = ~v12 & new_n4301_;
  assign new_n4303_ = ~v11 & new_n4302_;
  assign new_n4304_ = ~v10 & new_n4303_;
  assign new_n4305_ = ~v9 & new_n4304_;
  assign \v41.49  = ~v8 & new_n4305_;
  assign new_n4307_ = ~v12 & new_n158_;
  assign new_n4308_ = v4 & new_n4307_;
  assign new_n4309_ = v12 & v40;
  assign new_n4310_ = ~v4 & new_n4309_;
  assign new_n4311_ = ~new_n4308_ & ~new_n4310_;
  assign new_n4312_ = ~v3 & ~new_n4311_;
  assign new_n4313_ = v3 & new_n4307_;
  assign new_n4314_ = ~new_n4312_ & ~new_n4313_;
  assign new_n4315_ = ~v2 & ~new_n4314_;
  assign new_n4316_ = v2 & new_n4307_;
  assign new_n4317_ = ~new_n4315_ & ~new_n4316_;
  assign new_n4318_ = ~v1 & ~new_n4317_;
  assign new_n4319_ = v1 & new_n4307_;
  assign new_n4320_ = ~new_n4318_ & ~new_n4319_;
  assign new_n4321_ = ~v5 & ~new_n4320_;
  assign new_n4322_ = ~new_n156_ & ~new_n4285_;
  assign new_n4323_ = ~v18 & new_n4322_;
  assign new_n4324_ = ~v17 & new_n4323_;
  assign new_n4325_ = ~v12 & new_n4324_;
  assign new_n4326_ = v5 & new_n4325_;
  assign new_n4327_ = ~new_n4321_ & ~new_n4326_;
  assign new_n4328_ = v15 & ~new_n4327_;
  assign new_n4329_ = ~v3 & ~new_n390_;
  assign new_n4330_ = v18 & ~new_n4329_;
  assign new_n4331_ = v17 & new_n4330_;
  assign new_n4332_ = new_n256_ & new_n1061_;
  assign new_n4333_ = ~new_n4331_ & ~new_n4332_;
  assign new_n4334_ = v19 & ~new_n4333_;
  assign new_n4335_ = v16 & new_n4334_;
  assign new_n4336_ = ~v12 & new_n4335_;
  assign new_n4337_ = new_n256_ & new_n4309_;
  assign new_n4338_ = ~new_n4336_ & ~new_n4337_;
  assign new_n4339_ = ~v2 & ~new_n4338_;
  assign new_n4340_ = ~v12 & new_n446_;
  assign new_n4341_ = v2 & new_n4340_;
  assign new_n4342_ = ~new_n4339_ & ~new_n4341_;
  assign new_n4343_ = ~v1 & ~new_n4342_;
  assign new_n4344_ = v1 & new_n4340_;
  assign new_n4345_ = ~new_n4343_ & ~new_n4344_;
  assign new_n4346_ = ~v5 & ~new_n4345_;
  assign new_n4347_ = v19 & ~new_n4285_;
  assign new_n4348_ = v18 & new_n4347_;
  assign new_n4349_ = v17 & new_n4348_;
  assign new_n4350_ = v16 & new_n4349_;
  assign new_n4351_ = ~v12 & new_n4350_;
  assign new_n4352_ = v5 & new_n4351_;
  assign new_n4353_ = ~new_n4346_ & ~new_n4352_;
  assign new_n4354_ = ~v15 & ~new_n4353_;
  assign new_n4355_ = ~new_n4328_ & ~new_n4354_;
  assign new_n4356_ = ~v0 & ~new_n4355_;
  assign new_n4357_ = ~new_n638_ & ~new_n4356_;
  assign new_n4358_ = v13 & ~new_n4357_;
  assign new_n4359_ = ~v16 & ~new_n1866_;
  assign new_n4360_ = ~new_n1604_ & ~new_n4359_;
  assign new_n4361_ = ~v15 & ~new_n4360_;
  assign new_n4362_ = ~new_n3583_ & ~new_n4361_;
  assign new_n4363_ = v17 & ~new_n4362_;
  assign new_n4364_ = new_n117_ & new_n1259_;
  assign new_n4365_ = ~new_n4363_ & ~new_n4364_;
  assign new_n4366_ = v40 & ~new_n4365_;
  assign new_n4367_ = ~v5 & new_n4366_;
  assign new_n4368_ = ~new_n204_ & ~new_n4367_;
  assign new_n4369_ = ~v3 & ~new_n4368_;
  assign new_n4370_ = ~new_n211_ & ~new_n4369_;
  assign new_n4371_ = ~v0 & ~new_n4370_;
  assign new_n4372_ = new_n207_ & new_n498_;
  assign new_n4373_ = new_n210_ & new_n4372_;
  assign new_n4374_ = ~new_n4371_ & ~new_n4373_;
  assign new_n4375_ = ~v13 & ~new_n4374_;
  assign new_n4376_ = v12 & new_n4375_;
  assign new_n4377_ = ~v4 & new_n4376_;
  assign new_n4378_ = ~v2 & new_n4377_;
  assign new_n4379_ = ~v1 & new_n4378_;
  assign new_n4380_ = ~new_n4358_ & ~new_n4379_;
  assign new_n4381_ = ~v14 & ~new_n4380_;
  assign new_n4382_ = ~new_n246_ & ~new_n1190_;
  assign new_n4383_ = v13 & ~new_n4382_;
  assign new_n4384_ = v13 & ~new_n4383_;
  assign new_n4385_ = v40 & ~new_n4384_;
  assign new_n4386_ = v14 & new_n4385_;
  assign new_n4387_ = v12 & new_n4386_;
  assign new_n4388_ = ~v5 & new_n4387_;
  assign new_n4389_ = ~v4 & new_n4388_;
  assign new_n4390_ = ~v3 & new_n4389_;
  assign new_n4391_ = ~v2 & new_n4390_;
  assign new_n4392_ = ~v1 & new_n4391_;
  assign new_n4393_ = ~v0 & new_n4392_;
  assign new_n4394_ = ~new_n4381_ & ~new_n4393_;
  assign new_n4395_ = ~v36 & ~new_n4394_;
  assign new_n4396_ = ~v11 & new_n4395_;
  assign new_n4397_ = ~v10 & new_n4396_;
  assign new_n4398_ = ~v9 & new_n4397_;
  assign \v41.50  = ~v8 & new_n4398_;
  assign new_n4400_ = v1 & ~new_n1090_;
  assign new_n4401_ = ~new_n156_ & ~new_n672_;
  assign new_n4402_ = ~v4 & new_n4401_;
  assign new_n4403_ = ~v1 & new_n4402_;
  assign new_n4404_ = ~new_n4400_ & ~new_n4403_;
  assign new_n4405_ = ~v14 & ~new_n4404_;
  assign new_n4406_ = ~v12 & new_n4405_;
  assign new_n4407_ = ~v5 & new_n334_;
  assign new_n4408_ = ~v4 & new_n4407_;
  assign new_n4409_ = ~v1 & new_n4408_;
  assign new_n4410_ = ~new_n4406_ & ~new_n4409_;
  assign new_n4411_ = v15 & ~new_n4410_;
  assign new_n4412_ = ~v12 & ~new_n952_;
  assign new_n4413_ = ~v19 & ~new_n4412_;
  assign new_n4414_ = ~v12 & new_n3029_;
  assign new_n4415_ = ~new_n4413_ & ~new_n4414_;
  assign new_n4416_ = v16 & ~new_n4415_;
  assign new_n4417_ = new_n401_ & new_n3077_;
  assign new_n4418_ = ~new_n4416_ & ~new_n4417_;
  assign new_n4419_ = v40 & ~new_n4418_;
  assign new_n4420_ = ~v15 & new_n4419_;
  assign new_n4421_ = ~v5 & new_n4420_;
  assign new_n4422_ = ~v4 & new_n4421_;
  assign new_n4423_ = ~v1 & new_n4422_;
  assign new_n4424_ = ~new_n4411_ & ~new_n4423_;
  assign new_n4425_ = ~v18 & ~new_n4424_;
  assign new_n4426_ = v15 & new_n340_;
  assign new_n4427_ = v14 & new_n4426_;
  assign new_n4428_ = v12 & new_n4427_;
  assign new_n4429_ = ~v5 & new_n4428_;
  assign new_n4430_ = ~v4 & new_n4429_;
  assign new_n4431_ = ~v1 & new_n4430_;
  assign new_n4432_ = ~new_n4425_ & ~new_n4431_;
  assign new_n4433_ = ~v17 & ~new_n4432_;
  assign new_n4434_ = ~v12 & ~v16;
  assign new_n4435_ = new_n121_ & new_n4434_;
  assign new_n4436_ = ~v12 & ~new_n4435_;
  assign new_n4437_ = v15 & ~new_n4436_;
  assign new_n4438_ = ~v12 & new_n116_;
  assign new_n4439_ = new_n121_ & new_n4438_;
  assign new_n4440_ = ~new_n4437_ & ~new_n4439_;
  assign new_n4441_ = ~v14 & ~new_n4440_;
  assign new_n4442_ = ~v16 & new_n975_;
  assign new_n4443_ = ~v15 & new_n4442_;
  assign new_n4444_ = v14 & new_n4443_;
  assign new_n4445_ = v12 & new_n4444_;
  assign new_n4446_ = ~new_n4441_ & ~new_n4445_;
  assign new_n4447_ = v40 & ~new_n4446_;
  assign new_n4448_ = ~v5 & new_n4447_;
  assign new_n4449_ = new_n383_ & new_n1492_;
  assign new_n4450_ = new_n120_ & new_n673_;
  assign new_n4451_ = new_n4449_ & new_n4450_;
  assign new_n4452_ = ~new_n4448_ & ~new_n4451_;
  assign new_n4453_ = ~v4 & ~new_n4452_;
  assign new_n4454_ = ~v1 & new_n4453_;
  assign new_n4455_ = ~new_n4433_ & ~new_n4454_;
  assign new_n4456_ = v13 & ~new_n4455_;
  assign new_n4457_ = new_n203_ & new_n915_;
  assign new_n4458_ = ~v14 & ~new_n4457_;
  assign new_n4459_ = ~new_n121_ & ~new_n172_;
  assign new_n4460_ = ~v15 & ~new_n4459_;
  assign new_n4461_ = v15 & ~new_n2904_;
  assign new_n4462_ = ~new_n4460_ & ~new_n4461_;
  assign new_n4463_ = ~v16 & ~new_n4462_;
  assign new_n4464_ = ~new_n197_ & ~new_n4463_;
  assign new_n4465_ = ~v14 & ~new_n4464_;
  assign new_n4466_ = new_n4458_ & ~new_n4465_;
  assign new_n4467_ = v40 & ~new_n4466_;
  assign new_n4468_ = ~v5 & new_n4467_;
  assign new_n4469_ = v5 & new_n383_;
  assign new_n4470_ = new_n210_ & new_n4469_;
  assign new_n4471_ = ~new_n4468_ & ~new_n4470_;
  assign new_n4472_ = ~v13 & ~new_n4471_;
  assign new_n4473_ = v12 & new_n4472_;
  assign new_n4474_ = ~v4 & new_n4473_;
  assign new_n4475_ = ~v1 & new_n4474_;
  assign new_n4476_ = ~new_n4456_ & ~new_n4475_;
  assign new_n4477_ = ~v0 & ~new_n4476_;
  assign new_n4478_ = v4 & new_n2435_;
  assign new_n4479_ = ~new_n807_ & ~new_n4478_;
  assign new_n4480_ = ~v14 & ~new_n4479_;
  assign new_n4481_ = ~v1 & new_n4480_;
  assign new_n4482_ = v0 & new_n4481_;
  assign new_n4483_ = ~new_n4477_ & ~new_n4482_;
  assign new_n4484_ = ~v3 & ~new_n4483_;
  assign new_n4485_ = v0 & new_n2435_;
  assign new_n4486_ = ~v0 & v12;
  assign new_n4487_ = new_n766_ & new_n4486_;
  assign new_n4488_ = new_n210_ & new_n4487_;
  assign new_n4489_ = ~new_n4485_ & ~new_n4488_;
  assign new_n4490_ = ~v14 & ~new_n4489_;
  assign new_n4491_ = ~v5 & new_n4490_;
  assign new_n4492_ = ~v4 & new_n4491_;
  assign new_n4493_ = v3 & new_n4492_;
  assign new_n4494_ = ~v1 & new_n4493_;
  assign new_n4495_ = ~new_n4484_ & ~new_n4494_;
  assign new_n4496_ = ~v36 & ~new_n4495_;
  assign new_n4497_ = ~v11 & new_n4496_;
  assign new_n4498_ = ~v10 & new_n4497_;
  assign new_n4499_ = ~v9 & new_n4498_;
  assign new_n4500_ = ~v8 & new_n4499_;
  assign \v41.51  = ~v2 & new_n4500_;
  assign new_n4502_ = v13 & ~new_n610_;
  assign new_n4503_ = ~v12 & new_n4502_;
  assign new_n4504_ = ~v15 & new_n426_;
  assign new_n4505_ = new_n266_ & new_n4504_;
  assign new_n4506_ = ~new_n4503_ & ~new_n4505_;
  assign new_n4507_ = ~v17 & ~new_n4506_;
  assign new_n4508_ = new_n117_ & new_n1409_;
  assign new_n4509_ = new_n266_ & new_n4508_;
  assign new_n4510_ = ~new_n4507_ & ~new_n4509_;
  assign new_n4511_ = ~v19 & ~new_n4510_;
  assign new_n4512_ = v13 & new_n2081_;
  assign new_n4513_ = ~v12 & new_n4512_;
  assign new_n4514_ = v5 & new_n4513_;
  assign new_n4515_ = ~new_n4511_ & ~new_n4514_;
  assign new_n4516_ = ~v4 & ~new_n4515_;
  assign new_n4517_ = ~v17 & ~new_n402_;
  assign new_n4518_ = v15 & new_n4517_;
  assign new_n4519_ = v13 & new_n4518_;
  assign new_n4520_ = ~v12 & new_n4519_;
  assign new_n4521_ = v4 & new_n4520_;
  assign new_n4522_ = ~new_n4516_ & ~new_n4521_;
  assign new_n4523_ = ~v3 & ~new_n4522_;
  assign new_n4524_ = v3 & new_n4520_;
  assign new_n4525_ = ~new_n4523_ & ~new_n4524_;
  assign new_n4526_ = ~v2 & ~new_n4525_;
  assign new_n4527_ = v2 & new_n4520_;
  assign new_n4528_ = ~new_n4526_ & ~new_n4527_;
  assign new_n4529_ = ~v18 & ~new_n4528_;
  assign new_n4530_ = new_n257_ & new_n426_;
  assign new_n4531_ = ~new_n1115_ & ~new_n4530_;
  assign new_n4532_ = v19 & ~new_n4531_;
  assign new_n4533_ = v18 & new_n4532_;
  assign new_n4534_ = v17 & new_n4533_;
  assign new_n4535_ = v13 & new_n4534_;
  assign new_n4536_ = ~v12 & new_n4535_;
  assign new_n4537_ = ~v4 & new_n4536_;
  assign new_n4538_ = ~v3 & new_n4537_;
  assign new_n4539_ = ~v2 & new_n4538_;
  assign new_n4540_ = ~new_n4529_ & ~new_n4539_;
  assign new_n4541_ = ~v0 & ~new_n4540_;
  assign new_n4542_ = ~new_n351_ & ~new_n3838_;
  assign new_n4543_ = ~new_n248_ & ~new_n4542_;
  assign new_n4544_ = v16 & new_n4543_;
  assign new_n4545_ = v13 & new_n4544_;
  assign new_n4546_ = ~v12 & new_n4545_;
  assign new_n4547_ = ~v4 & new_n4546_;
  assign new_n4548_ = ~v2 & new_n4547_;
  assign new_n4549_ = v0 & new_n4548_;
  assign new_n4550_ = ~new_n4541_ & ~new_n4549_;
  assign new_n4551_ = ~v1 & ~new_n4550_;
  assign new_n4552_ = ~v5 & ~new_n402_;
  assign new_n4553_ = v5 & new_n400_;
  assign new_n4554_ = ~new_n4552_ & ~new_n4553_;
  assign new_n4555_ = ~v18 & ~new_n4554_;
  assign new_n4556_ = ~v17 & new_n4555_;
  assign new_n4557_ = v15 & new_n4556_;
  assign new_n4558_ = v13 & new_n4557_;
  assign new_n4559_ = ~v12 & new_n4558_;
  assign new_n4560_ = ~v4 & new_n4559_;
  assign new_n4561_ = ~v3 & new_n4560_;
  assign new_n4562_ = ~v2 & new_n4561_;
  assign new_n4563_ = v1 & new_n4562_;
  assign new_n4564_ = ~v0 & new_n4563_;
  assign new_n4565_ = ~new_n4551_ & ~new_n4564_;
  assign new_n4566_ = ~v14 & ~new_n4565_;
  assign new_n4567_ = ~v0 & new_n380_;
  assign new_n4568_ = new_n256_ & new_n1634_;
  assign new_n4569_ = new_n4567_ & new_n4568_;
  assign new_n4570_ = new_n201_ & new_n1338_;
  assign new_n4571_ = new_n119_ & new_n1595_;
  assign new_n4572_ = new_n4570_ & new_n4571_;
  assign new_n4573_ = new_n4569_ & new_n4572_;
  assign new_n4574_ = ~new_n4566_ & ~new_n4573_;
  assign new_n4575_ = ~v36 & ~new_n4574_;
  assign new_n4576_ = ~v11 & new_n4575_;
  assign new_n4577_ = ~v10 & new_n4576_;
  assign new_n4578_ = ~v9 & new_n4577_;
  assign \v41.52  = ~v8 & new_n4578_;
  assign new_n4580_ = new_n265_ & new_n1186_;
  assign new_n4581_ = v15 & new_n164_;
  assign new_n4582_ = new_n849_ & new_n4581_;
  assign new_n4583_ = ~new_n4580_ & ~new_n4582_;
  assign new_n4584_ = v5 & ~new_n4583_;
  assign new_n4585_ = new_n209_ & new_n265_;
  assign new_n4586_ = new_n164_ & new_n849_;
  assign new_n4587_ = ~new_n4585_ & ~new_n4586_;
  assign new_n4588_ = v40 & ~new_n4587_;
  assign new_n4589_ = v15 & new_n4588_;
  assign new_n4590_ = ~v5 & new_n4589_;
  assign new_n4591_ = ~new_n4584_ & ~new_n4590_;
  assign new_n4592_ = ~v19 & ~new_n4591_;
  assign new_n4593_ = v40 & ~new_n1331_;
  assign new_n4594_ = v19 & new_n4593_;
  assign new_n4595_ = ~v17 & new_n4594_;
  assign new_n4596_ = v13 & new_n4595_;
  assign new_n4597_ = ~v12 & new_n4596_;
  assign new_n4598_ = ~v5 & new_n4597_;
  assign new_n4599_ = ~new_n4592_ & ~new_n4598_;
  assign new_n4600_ = ~v18 & ~new_n4599_;
  assign new_n4601_ = v40 & ~new_n4440_;
  assign new_n4602_ = v13 & new_n4601_;
  assign new_n4603_ = ~v5 & new_n4602_;
  assign new_n4604_ = ~new_n4600_ & ~new_n4603_;
  assign new_n4605_ = ~v14 & ~new_n4604_;
  assign new_n4606_ = new_n164_ & new_n171_;
  assign new_n4607_ = ~new_n3276_ & ~new_n4606_;
  assign new_n4608_ = ~v15 & ~new_n4607_;
  assign new_n4609_ = ~new_n4581_ & ~new_n4608_;
  assign new_n4610_ = v40 & ~new_n4609_;
  assign new_n4611_ = v14 & new_n4610_;
  assign new_n4612_ = v13 & new_n4611_;
  assign new_n4613_ = v12 & new_n4612_;
  assign new_n4614_ = ~v5 & new_n4613_;
  assign new_n4615_ = ~new_n4605_ & ~new_n4614_;
  assign new_n4616_ = ~v1 & ~new_n4615_;
  assign new_n4617_ = v1 & v5;
  assign new_n4618_ = new_n1445_ & new_n4617_;
  assign new_n4619_ = new_n2027_ & new_n4618_;
  assign new_n4620_ = ~new_n4616_ & ~new_n4619_;
  assign new_n4621_ = ~v0 & ~new_n4620_;
  assign new_n4622_ = v0 & ~v1;
  assign new_n4623_ = v5 & new_n849_;
  assign new_n4624_ = new_n4622_ & new_n4623_;
  assign new_n4625_ = ~v14 & new_n116_;
  assign new_n4626_ = new_n121_ & new_n4625_;
  assign new_n4627_ = new_n4624_ & new_n4626_;
  assign new_n4628_ = ~new_n4621_ & ~new_n4627_;
  assign new_n4629_ = ~v36 & ~new_n4628_;
  assign new_n4630_ = ~v11 & new_n4629_;
  assign new_n4631_ = ~v10 & new_n4630_;
  assign new_n4632_ = ~v9 & new_n4631_;
  assign new_n4633_ = ~v8 & new_n4632_;
  assign new_n4634_ = ~v4 & new_n4633_;
  assign new_n4635_ = ~v3 & new_n4634_;
  assign \v41.53  = ~v2 & new_n4635_;
  assign new_n4637_ = new_n117_ & new_n119_;
  assign new_n4638_ = ~new_n602_ & ~new_n4637_;
  assign new_n4639_ = v4 & ~new_n4638_;
  assign new_n4640_ = ~v4 & new_n600_;
  assign new_n4641_ = ~new_n4639_ & ~new_n4640_;
  assign new_n4642_ = v19 & ~new_n4641_;
  assign new_n4643_ = ~v4 & new_n116_;
  assign new_n4644_ = new_n4571_ & new_n4643_;
  assign new_n4645_ = ~new_n4642_ & ~new_n4644_;
  assign new_n4646_ = ~v12 & ~new_n4645_;
  assign new_n4647_ = ~v15 & ~new_n2721_;
  assign new_n4648_ = ~new_n2176_ & new_n4647_;
  assign new_n4649_ = v40 & ~new_n4648_;
  assign new_n4650_ = v12 & new_n4649_;
  assign new_n4651_ = ~v4 & new_n4650_;
  assign new_n4652_ = ~new_n4646_ & ~new_n4651_;
  assign new_n4653_ = v13 & ~new_n4652_;
  assign new_n4654_ = v40 & ~new_n1147_;
  assign new_n4655_ = ~v19 & new_n4654_;
  assign new_n4656_ = ~v18 & new_n4655_;
  assign new_n4657_ = ~v16 & new_n4656_;
  assign new_n4658_ = ~v13 & new_n4657_;
  assign new_n4659_ = v12 & new_n4658_;
  assign new_n4660_ = ~v4 & new_n4659_;
  assign new_n4661_ = ~new_n4653_ & ~new_n4660_;
  assign new_n4662_ = ~v14 & ~new_n4661_;
  assign new_n4663_ = new_n1349_ & new_n1998_;
  assign new_n4664_ = new_n259_ & new_n1596_;
  assign new_n4665_ = new_n4663_ & new_n4664_;
  assign new_n4666_ = ~new_n4662_ & ~new_n4665_;
  assign new_n4667_ = ~v5 & ~new_n4666_;
  assign new_n4668_ = new_n403_ & new_n1445_;
  assign new_n4669_ = new_n172_ & new_n1771_;
  assign new_n4670_ = new_n4668_ & new_n4669_;
  assign new_n4671_ = ~new_n4667_ & ~new_n4670_;
  assign new_n4672_ = ~v36 & ~new_n4671_;
  assign new_n4673_ = ~v11 & new_n4672_;
  assign new_n4674_ = ~v10 & new_n4673_;
  assign new_n4675_ = ~v9 & new_n4674_;
  assign new_n4676_ = ~v8 & new_n4675_;
  assign new_n4677_ = ~v3 & new_n4676_;
  assign new_n4678_ = ~v2 & new_n4677_;
  assign new_n4679_ = ~v1 & new_n4678_;
  assign \v41.54  = ~v0 & new_n4679_;
  assign new_n4681_ = v14 & new_n2150_;
  assign new_n4682_ = v14 & ~new_n4681_;
  assign new_n4683_ = v16 & ~new_n4682_;
  assign new_n4684_ = ~new_n915_ & ~new_n4683_;
  assign new_n4685_ = v40 & ~new_n4684_;
  assign new_n4686_ = ~v36 & new_n4685_;
  assign new_n4687_ = v15 & new_n4686_;
  assign new_n4688_ = v13 & new_n4687_;
  assign new_n4689_ = v12 & new_n4688_;
  assign new_n4690_ = ~v11 & new_n4689_;
  assign new_n4691_ = ~v10 & new_n4690_;
  assign new_n4692_ = ~v9 & new_n4691_;
  assign new_n4693_ = ~v8 & new_n4692_;
  assign new_n4694_ = ~v5 & new_n4693_;
  assign new_n4695_ = ~v4 & new_n4694_;
  assign new_n4696_ = ~v3 & new_n4695_;
  assign new_n4697_ = ~v2 & new_n4696_;
  assign new_n4698_ = ~v1 & new_n4697_;
  assign \v41.55  = ~v0 & new_n4698_;
  assign new_n4700_ = v19 & ~new_n4638_;
  assign new_n4701_ = ~v12 & new_n4700_;
  assign new_n4702_ = v4 & new_n4701_;
  assign new_n4703_ = ~v15 & ~new_n602_;
  assign new_n4704_ = v40 & ~new_n4703_;
  assign new_n4705_ = v12 & new_n4704_;
  assign new_n4706_ = ~v4 & new_n4705_;
  assign new_n4707_ = ~new_n4702_ & ~new_n4706_;
  assign new_n4708_ = ~v5 & ~new_n4707_;
  assign new_n4709_ = new_n403_ & new_n2170_;
  assign new_n4710_ = new_n4606_ & new_n4709_;
  assign new_n4711_ = ~new_n4708_ & ~new_n4710_;
  assign new_n4712_ = ~v36 & ~new_n4711_;
  assign new_n4713_ = ~v14 & new_n4712_;
  assign new_n4714_ = v13 & new_n4713_;
  assign new_n4715_ = ~v11 & new_n4714_;
  assign new_n4716_ = ~v10 & new_n4715_;
  assign new_n4717_ = ~v9 & new_n4716_;
  assign new_n4718_ = ~v8 & new_n4717_;
  assign new_n4719_ = ~v3 & new_n4718_;
  assign new_n4720_ = ~v2 & new_n4719_;
  assign new_n4721_ = ~v1 & new_n4720_;
  assign \v41.56  = ~v0 & new_n4721_;
  assign new_n4723_ = v16 & new_n1061_;
  assign new_n4724_ = ~v4 & new_n4723_;
  assign new_n4725_ = ~new_n4639_ & ~new_n4724_;
  assign new_n4726_ = v19 & ~new_n4725_;
  assign new_n4727_ = ~v4 & new_n117_;
  assign new_n4728_ = new_n4571_ & new_n4727_;
  assign new_n4729_ = ~new_n4726_ & ~new_n4728_;
  assign new_n4730_ = ~v12 & ~new_n4729_;
  assign new_n4731_ = ~v15 & ~new_n2176_;
  assign new_n4732_ = v40 & ~new_n4731_;
  assign new_n4733_ = v12 & new_n4732_;
  assign new_n4734_ = ~v4 & new_n4733_;
  assign new_n4735_ = ~new_n4730_ & ~new_n4734_;
  assign new_n4736_ = ~v14 & ~new_n4735_;
  assign new_n4737_ = v12 & new_n3619_;
  assign new_n4738_ = ~v4 & new_n4737_;
  assign new_n4739_ = ~new_n4736_ & ~new_n4738_;
  assign new_n4740_ = ~v5 & ~new_n4739_;
  assign new_n4741_ = new_n403_ & new_n952_;
  assign new_n4742_ = new_n4669_ & new_n4741_;
  assign new_n4743_ = ~new_n4740_ & ~new_n4742_;
  assign new_n4744_ = v13 & ~new_n4743_;
  assign new_n4745_ = new_n403_ & new_n3954_;
  assign new_n4746_ = new_n268_ & new_n4745_;
  assign new_n4747_ = ~new_n4744_ & ~new_n4746_;
  assign new_n4748_ = ~v36 & ~new_n4747_;
  assign new_n4749_ = ~v11 & new_n4748_;
  assign new_n4750_ = ~v10 & new_n4749_;
  assign new_n4751_ = ~v9 & new_n4750_;
  assign new_n4752_ = ~v8 & new_n4751_;
  assign new_n4753_ = ~v3 & new_n4752_;
  assign new_n4754_ = ~v2 & new_n4753_;
  assign new_n4755_ = ~v1 & new_n4754_;
  assign \v41.57  = ~v0 & new_n4755_;
  assign new_n4757_ = v40 & ~new_n402_;
  assign new_n4758_ = ~v17 & new_n4757_;
  assign new_n4759_ = v15 & new_n4758_;
  assign new_n4760_ = v13 & new_n4759_;
  assign new_n4761_ = ~v12 & new_n4760_;
  assign new_n4762_ = ~v5 & new_n4761_;
  assign new_n4763_ = v5 & new_n265_;
  assign new_n4764_ = new_n1773_ & new_n4763_;
  assign new_n4765_ = ~new_n4762_ & ~new_n4764_;
  assign new_n4766_ = ~v36 & ~new_n4765_;
  assign new_n4767_ = ~v18 & new_n4766_;
  assign new_n4768_ = ~v14 & new_n4767_;
  assign new_n4769_ = ~v11 & new_n4768_;
  assign new_n4770_ = ~v10 & new_n4769_;
  assign new_n4771_ = ~v9 & new_n4770_;
  assign new_n4772_ = ~v8 & new_n4771_;
  assign new_n4773_ = ~v4 & new_n4772_;
  assign new_n4774_ = ~v3 & new_n4773_;
  assign new_n4775_ = ~v2 & new_n4774_;
  assign new_n4776_ = ~v1 & new_n4775_;
  assign \v41.58  = ~v0 & new_n4776_;
  assign new_n4778_ = v14 & new_n164_;
  assign new_n4779_ = v14 & ~new_n4778_;
  assign new_n4780_ = v40 & ~new_n4779_;
  assign new_n4781_ = ~v36 & new_n4780_;
  assign new_n4782_ = v15 & new_n4781_;
  assign new_n4783_ = v13 & new_n4782_;
  assign new_n4784_ = v12 & new_n4783_;
  assign new_n4785_ = ~v11 & new_n4784_;
  assign new_n4786_ = ~v10 & new_n4785_;
  assign new_n4787_ = ~v9 & new_n4786_;
  assign new_n4788_ = ~v8 & new_n4787_;
  assign new_n4789_ = ~v5 & new_n4788_;
  assign new_n4790_ = ~v4 & new_n4789_;
  assign new_n4791_ = ~v3 & new_n4790_;
  assign new_n4792_ = ~v2 & new_n4791_;
  assign new_n4793_ = ~v1 & new_n4792_;
  assign \v41.59  = ~v0 & new_n4793_;
  assign new_n4795_ = ~v2 & new_n2341_;
  assign new_n4796_ = ~v3 & new_n4795_;
  assign new_n4797_ = ~v4 & new_n4796_;
  assign new_n4798_ = v5 & new_n4797_;
  assign new_n4799_ = ~v8 & new_n4798_;
  assign new_n4800_ = ~v9 & new_n4799_;
  assign new_n4801_ = ~v10 & new_n4800_;
  assign new_n4802_ = ~v11 & new_n4801_;
  assign new_n4803_ = ~v12 & new_n4802_;
  assign new_n4804_ = v13 & new_n4803_;
  assign new_n4805_ = ~v14 & new_n4804_;
  assign new_n4806_ = ~v15 & new_n4805_;
  assign new_n4807_ = v16 & new_n4806_;
  assign new_n4808_ = v17 & new_n4807_;
  assign new_n4809_ = ~v18 & new_n4808_;
  assign new_n4810_ = ~v19 & new_n4809_;
  assign \v41.60  = ~v36 & new_n4810_;
  assign new_n4812_ = ~v9 & new_n3204_;
  assign new_n4813_ = ~v8 & new_n4812_;
  assign new_n4814_ = ~v5 & new_n4813_;
  assign new_n4815_ = ~v4 & new_n4814_;
  assign new_n4816_ = ~v3 & new_n4815_;
  assign new_n4817_ = ~v2 & new_n4816_;
  assign new_n4818_ = ~v1 & new_n4817_;
  assign \v41.61  = ~v0 & new_n4818_;
  assign new_n4820_ = ~v5 & ~v14;
  assign new_n4821_ = v5 & new_n2325_;
  assign new_n4822_ = ~new_n4820_ & ~new_n4821_;
  assign new_n4823_ = v5 & v14;
  assign new_n4824_ = new_n226_ & new_n4823_;
  assign new_n4825_ = new_n4822_ & ~new_n4824_;
  assign new_n4826_ = ~v13 & ~new_n4825_;
  assign new_n4827_ = ~v12 & new_n4826_;
  assign new_n4828_ = v14 & new_n1145_;
  assign new_n4829_ = new_n3296_ & new_n4828_;
  assign new_n4830_ = ~new_n4827_ & ~new_n4829_;
  assign new_n4831_ = ~v5 & v13;
  assign new_n4832_ = ~v14 & new_n1145_;
  assign new_n4833_ = new_n4831_ & new_n4832_;
  assign new_n4834_ = v5 & ~v13;
  assign new_n4835_ = v14 & new_n1146_;
  assign new_n4836_ = new_n4834_ & new_n4835_;
  assign new_n4837_ = ~new_n4833_ & ~new_n4836_;
  assign new_n4838_ = ~v12 & ~new_n4837_;
  assign new_n4839_ = new_n226_ & new_n1338_;
  assign new_n4840_ = ~new_n1357_ & ~new_n4839_;
  assign new_n4841_ = v12 & ~new_n4840_;
  assign new_n4842_ = v5 & new_n4841_;
  assign new_n4843_ = ~new_n4838_ & ~new_n4842_;
  assign new_n4844_ = v16 & ~new_n4843_;
  assign new_n4845_ = new_n4830_ & ~new_n4844_;
  assign new_n4846_ = new_n1356_ & new_n2116_;
  assign new_n4847_ = new_n765_ & new_n900_;
  assign new_n4848_ = ~new_n4846_ & ~new_n4847_;
  assign new_n4849_ = v18 & ~new_n4848_;
  assign new_n4850_ = ~v17 & new_n4849_;
  assign new_n4851_ = v16 & new_n4850_;
  assign new_n4852_ = v13 & new_n4851_;
  assign new_n4853_ = new_n4845_ & ~new_n4852_;
  assign new_n4854_ = v40 & ~new_n4853_;
  assign new_n4855_ = ~v3 & new_n4854_;
  assign new_n4856_ = new_n849_ & new_n3838_;
  assign new_n4857_ = new_n1487_ & new_n4856_;
  assign new_n4858_ = ~new_n4855_ & ~new_n4857_;
  assign new_n4859_ = new_n900_ & new_n4831_;
  assign new_n4860_ = new_n210_ & new_n4859_;
  assign new_n4861_ = ~new_n1370_ & ~new_n4860_;
  assign new_n4862_ = v12 & ~new_n4861_;
  assign new_n4863_ = new_n1902_ & new_n2116_;
  assign new_n4864_ = new_n172_ & new_n201_;
  assign new_n4865_ = new_n4863_ & new_n4864_;
  assign new_n4866_ = ~new_n4862_ & ~new_n4865_;
  assign new_n4867_ = v40 & ~new_n4866_;
  assign new_n4868_ = ~v3 & new_n4867_;
  assign new_n4869_ = new_n4858_ & ~new_n4868_;
  assign new_n4870_ = ~v8 & ~new_n4869_;
  assign new_n4871_ = ~v5 & v8;
  assign new_n4872_ = ~v3 & new_n4871_;
  assign new_n4873_ = ~new_n4870_ & ~new_n4872_;
  assign new_n4874_ = ~v11 & ~new_n4873_;
  assign new_n4875_ = v8 & v11;
  assign new_n4876_ = new_n2673_ & new_n4875_;
  assign new_n4877_ = ~new_n4874_ & ~new_n4876_;
  assign new_n4878_ = ~v10 & ~new_n4877_;
  assign new_n4879_ = v8 & v10;
  assign new_n4880_ = ~v5 & new_n4879_;
  assign new_n4881_ = ~v3 & new_n4880_;
  assign new_n4882_ = ~new_n4878_ & ~new_n4881_;
  assign new_n4883_ = ~v36 & ~new_n4882_;
  assign new_n4884_ = ~v9 & new_n4883_;
  assign new_n4885_ = ~v4 & new_n4884_;
  assign new_n4886_ = ~v2 & new_n4885_;
  assign new_n4887_ = ~v1 & new_n4886_;
  assign \v41.62  = ~v0 & new_n4887_;
  assign new_n4889_ = new_n246_ & new_n1777_;
  assign new_n4890_ = ~new_n1916_ & ~new_n4889_;
  assign new_n4891_ = ~v18 & ~new_n4890_;
  assign new_n4892_ = ~v13 & new_n4891_;
  assign new_n4893_ = v12 & new_n4892_;
  assign new_n4894_ = v18 & ~v39;
  assign new_n4895_ = ~v17 & new_n4894_;
  assign new_n4896_ = v15 & new_n4895_;
  assign new_n4897_ = v13 & new_n4896_;
  assign new_n4898_ = ~v12 & new_n4897_;
  assign new_n4899_ = ~new_n4893_ & ~new_n4898_;
  assign new_n4900_ = v40 & ~new_n4899_;
  assign new_n4901_ = ~v38 & new_n4900_;
  assign new_n4902_ = v37 & new_n4901_;
  assign new_n4903_ = ~v16 & new_n4902_;
  assign new_n4904_ = ~v14 & new_n4903_;
  assign new_n4905_ = ~v11 & new_n4904_;
  assign new_n4906_ = ~v10 & new_n4905_;
  assign new_n4907_ = ~v8 & new_n4906_;
  assign new_n4908_ = ~v8 & ~new_n4907_;
  assign new_n4909_ = ~v36 & ~new_n4908_;
  assign new_n4910_ = ~v9 & new_n4909_;
  assign new_n4911_ = ~v5 & new_n4910_;
  assign new_n4912_ = ~v4 & new_n4911_;
  assign new_n4913_ = ~v3 & new_n4912_;
  assign new_n4914_ = ~v2 & new_n4913_;
  assign new_n4915_ = ~v1 & new_n4914_;
  assign \v41.63  = ~v0 & new_n4915_;
  assign new_n4917_ = ~v5 & new_n4797_;
  assign new_n4918_ = ~v8 & new_n4917_;
  assign new_n4919_ = ~v9 & new_n4918_;
  assign new_n4920_ = ~v10 & new_n4919_;
  assign new_n4921_ = ~v11 & new_n4920_;
  assign new_n4922_ = ~v12 & new_n4921_;
  assign new_n4923_ = v13 & new_n4922_;
  assign new_n4924_ = ~v14 & new_n4923_;
  assign new_n4925_ = v15 & new_n4924_;
  assign new_n4926_ = ~v16 & new_n4925_;
  assign new_n4927_ = ~v17 & new_n4926_;
  assign new_n4928_ = v18 & new_n4927_;
  assign new_n4929_ = v19 & new_n4928_;
  assign new_n4930_ = ~v36 & new_n4929_;
  assign new_n4931_ = ~v37 & new_n4930_;
  assign new_n4932_ = ~v38 & new_n4931_;
  assign new_n4933_ = ~v39 & new_n4932_;
  assign \v41.64  = v40 & new_n4933_;
  assign new_n4935_ = v14 & new_n304_;
  assign new_n4936_ = v13 & new_n4935_;
  assign new_n4937_ = new_n2283_ & new_n4213_;
  assign new_n4938_ = ~new_n4936_ & ~new_n4937_;
  assign new_n4939_ = v14 & ~v16;
  assign new_n4940_ = new_n975_ & new_n4939_;
  assign new_n4941_ = new_n976_ & new_n1339_;
  assign new_n4942_ = ~new_n4940_ & ~new_n4941_;
  assign new_n4943_ = v13 & ~new_n4942_;
  assign new_n4944_ = v17 & ~new_n402_;
  assign new_n4945_ = ~v14 & new_n4944_;
  assign new_n4946_ = ~v13 & new_n4945_;
  assign new_n4947_ = ~new_n4943_ & ~new_n4946_;
  assign new_n4948_ = ~v18 & ~new_n4947_;
  assign new_n4949_ = new_n121_ & new_n915_;
  assign new_n4950_ = ~v14 & ~new_n4949_;
  assign new_n4951_ = ~v13 & ~new_n4950_;
  assign new_n4952_ = ~new_n4948_ & ~new_n4951_;
  assign new_n4953_ = ~v15 & ~new_n4952_;
  assign new_n4954_ = ~v14 & new_n2905_;
  assign new_n4955_ = ~v14 & ~new_n4954_;
  assign new_n4956_ = v15 & ~new_n4955_;
  assign new_n4957_ = ~v13 & new_n4956_;
  assign new_n4958_ = ~new_n4953_ & ~new_n4957_;
  assign new_n4959_ = new_n4938_ & new_n4958_;
  assign new_n4960_ = v12 & ~new_n4959_;
  assign new_n4961_ = new_n849_ & new_n1356_;
  assign new_n4962_ = new_n165_ & new_n209_;
  assign new_n4963_ = new_n4961_ & new_n4962_;
  assign new_n4964_ = ~new_n4960_ & ~new_n4963_;
  assign new_n4965_ = v40 & ~new_n4964_;
  assign new_n4966_ = ~v3 & new_n4965_;
  assign new_n4967_ = ~new_n3793_ & ~new_n4966_;
  assign new_n4968_ = ~v0 & ~new_n4967_;
  assign new_n4969_ = ~new_n4252_ & ~new_n4968_;
  assign new_n4970_ = ~v36 & ~new_n4969_;
  assign new_n4971_ = ~v11 & new_n4970_;
  assign new_n4972_ = ~v10 & new_n4971_;
  assign new_n4973_ = ~v9 & new_n4972_;
  assign new_n4974_ = ~v8 & new_n4973_;
  assign new_n4975_ = ~v5 & new_n4974_;
  assign new_n4976_ = ~v4 & new_n4975_;
  assign new_n4977_ = ~v2 & new_n4976_;
  assign \v41.65  = ~v1 & new_n4977_;
  assign new_n4979_ = ~v2 & v4;
  assign new_n4980_ = v2 & ~v4;
  assign new_n4981_ = ~new_n4979_ & ~new_n4980_;
  assign new_n4982_ = ~v21 & ~new_n4981_;
  assign new_n4983_ = v20 & new_n4982_;
  assign new_n4984_ = v4 & new_n684_;
  assign new_n4985_ = ~v2 & new_n4984_;
  assign new_n4986_ = ~new_n4983_ & ~new_n4985_;
  assign new_n4987_ = ~new_n672_ & ~new_n4060_;
  assign new_n4988_ = new_n2247_ & new_n2273_;
  assign new_n4989_ = v26 & v40;
  assign new_n4990_ = new_n1512_ & new_n4989_;
  assign new_n4991_ = new_n4988_ & new_n4990_;
  assign new_n4992_ = ~new_n4987_ & ~new_n4991_;
  assign new_n4993_ = ~v4 & ~new_n4992_;
  assign new_n4994_ = ~v2 & new_n4993_;
  assign new_n4995_ = new_n4986_ & ~new_n4994_;
  assign new_n4996_ = v27 & ~new_n4995_;
  assign new_n4997_ = ~new_n672_ & ~new_n685_;
  assign new_n4998_ = ~v23 & ~new_n689_;
  assign new_n4999_ = v22 & ~new_n4998_;
  assign new_n5000_ = ~new_n692_ & ~new_n4999_;
  assign new_n5001_ = v40 & ~new_n5000_;
  assign new_n5002_ = v21 & new_n5001_;
  assign new_n5003_ = ~v20 & new_n5002_;
  assign new_n5004_ = ~v5 & new_n5003_;
  assign new_n5005_ = ~new_n4997_ & ~new_n5004_;
  assign new_n5006_ = ~v27 & ~new_n5005_;
  assign new_n5007_ = ~v5 & v20;
  assign new_n5008_ = new_n4067_ & new_n5007_;
  assign new_n5009_ = ~new_n5006_ & ~new_n5008_;
  assign new_n5010_ = ~v4 & ~new_n5009_;
  assign new_n5011_ = ~v2 & new_n5010_;
  assign new_n5012_ = ~new_n4996_ & ~new_n5011_;
  assign new_n5013_ = ~v19 & ~new_n5012_;
  assign new_n5014_ = ~v2 & ~v4;
  assign new_n5015_ = ~v5 & new_n1648_;
  assign new_n5016_ = new_n5014_ & new_n5015_;
  assign new_n5017_ = ~new_n5013_ & ~new_n5016_;
  assign new_n5018_ = v18 & ~new_n5017_;
  assign new_n5019_ = ~v16 & new_n5018_;
  assign new_n5020_ = ~v2 & new_n169_;
  assign new_n5021_ = new_n953_ & new_n1648_;
  assign new_n5022_ = new_n5020_ & new_n5021_;
  assign new_n5023_ = ~new_n5019_ & ~new_n5022_;
  assign new_n5024_ = ~v3 & ~new_n5023_;
  assign new_n5025_ = v5 & ~v16;
  assign new_n5026_ = ~v4 & new_n5025_;
  assign new_n5027_ = new_n329_ & new_n5026_;
  assign new_n5028_ = new_n1038_ & new_n1239_;
  assign new_n5029_ = new_n5027_ & new_n5028_;
  assign new_n5030_ = ~new_n5024_ & ~new_n5029_;
  assign new_n5031_ = ~v36 & ~new_n5030_;
  assign new_n5032_ = v17 & new_n5031_;
  assign new_n5033_ = ~v15 & new_n5032_;
  assign new_n5034_ = ~v14 & new_n5033_;
  assign new_n5035_ = ~v13 & new_n5034_;
  assign new_n5036_ = v12 & new_n5035_;
  assign new_n5037_ = ~v11 & new_n5036_;
  assign new_n5038_ = ~v10 & new_n5037_;
  assign new_n5039_ = ~v9 & new_n5038_;
  assign new_n5040_ = ~v8 & new_n5039_;
  assign new_n5041_ = ~v1 & new_n5040_;
  assign \v41.66  = ~v0 & new_n5041_;
  assign new_n5043_ = v5 & ~new_n1223_;
  assign new_n5044_ = ~v5 & new_n722_;
  assign new_n5045_ = ~new_n5043_ & ~new_n5044_;
  assign new_n5046_ = v3 & ~new_n5045_;
  assign new_n5047_ = ~v2 & new_n5046_;
  assign new_n5048_ = ~v5 & new_n1541_;
  assign new_n5049_ = new_n2269_ & new_n5048_;
  assign new_n5050_ = ~new_n5047_ & ~new_n5049_;
  assign new_n5051_ = ~v4 & ~new_n5050_;
  assign new_n5052_ = v5 & new_n1541_;
  assign new_n5053_ = new_n2364_ & new_n5052_;
  assign new_n5054_ = ~new_n5051_ & ~new_n5053_;
  assign new_n5055_ = ~new_n681_ & ~new_n5054_;
  assign new_n5056_ = v4 & ~new_n1209_;
  assign new_n5057_ = ~v4 & v22;
  assign new_n5058_ = new_n4138_ & new_n5057_;
  assign new_n5059_ = ~new_n5056_ & ~new_n5058_;
  assign new_n5060_ = v27 & ~new_n5059_;
  assign new_n5061_ = v23 & ~v27;
  assign new_n5062_ = v22 & new_n5061_;
  assign new_n5063_ = ~v4 & new_n5062_;
  assign new_n5064_ = ~new_n5060_ & ~new_n5063_;
  assign new_n5065_ = ~v5 & ~new_n5064_;
  assign new_n5066_ = v5 & new_n1544_;
  assign new_n5067_ = ~v4 & new_n5066_;
  assign new_n5068_ = ~new_n5065_ & ~new_n5067_;
  assign new_n5069_ = v3 & ~new_n5068_;
  assign new_n5070_ = ~v2 & new_n5069_;
  assign new_n5071_ = ~new_n5055_ & ~new_n5070_;
  assign new_n5072_ = v21 & ~new_n5071_;
  assign new_n5073_ = ~v20 & new_n5072_;
  assign new_n5074_ = v18 & new_n5073_;
  assign new_n5075_ = ~v2 & new_n256_;
  assign new_n5076_ = ~v5 & new_n385_;
  assign new_n5077_ = new_n5075_ & new_n5076_;
  assign new_n5078_ = ~new_n5074_ & ~new_n5077_;
  assign new_n5079_ = ~v36 & ~new_n5078_;
  assign new_n5080_ = ~v19 & new_n5079_;
  assign new_n5081_ = v17 & new_n5080_;
  assign new_n5082_ = ~v16 & new_n5081_;
  assign new_n5083_ = ~v15 & new_n5082_;
  assign new_n5084_ = ~v14 & new_n5083_;
  assign new_n5085_ = ~v13 & new_n5084_;
  assign new_n5086_ = v12 & new_n5085_;
  assign new_n5087_ = ~v11 & new_n5086_;
  assign new_n5088_ = ~v10 & new_n5087_;
  assign new_n5089_ = ~v9 & new_n5088_;
  assign new_n5090_ = ~v8 & new_n5089_;
  assign new_n5091_ = ~v1 & new_n5090_;
  assign \v41.67  = ~v0 & new_n5091_;
  assign new_n5093_ = v14 & ~v17;
  assign new_n5094_ = v13 & new_n5093_;
  assign new_n5095_ = new_n183_ & new_n1343_;
  assign new_n5096_ = ~new_n5094_ & ~new_n5095_;
  assign new_n5097_ = v15 & ~new_n5096_;
  assign new_n5098_ = ~v14 & new_n2080_;
  assign new_n5099_ = ~v13 & new_n5098_;
  assign new_n5100_ = ~new_n5097_ & ~new_n5099_;
  assign new_n5101_ = v40 & ~new_n5100_;
  assign new_n5102_ = ~v5 & new_n5101_;
  assign new_n5103_ = v17 & new_n1047_;
  assign new_n5104_ = ~v15 & new_n5103_;
  assign new_n5105_ = ~v14 & new_n5104_;
  assign new_n5106_ = ~v13 & new_n5105_;
  assign new_n5107_ = v5 & new_n5106_;
  assign new_n5108_ = ~new_n5102_ & ~new_n5107_;
  assign new_n5109_ = ~v4 & ~new_n5108_;
  assign new_n5110_ = v17 & new_n775_;
  assign new_n5111_ = ~v15 & new_n5110_;
  assign new_n5112_ = ~v14 & new_n5111_;
  assign new_n5113_ = ~v13 & new_n5112_;
  assign new_n5114_ = v4 & new_n5113_;
  assign new_n5115_ = ~new_n5109_ & ~new_n5114_;
  assign new_n5116_ = v18 & ~new_n5115_;
  assign new_n5117_ = new_n169_ & new_n1343_;
  assign new_n5118_ = new_n1145_ & new_n1649_;
  assign new_n5119_ = new_n5117_ & new_n5118_;
  assign new_n5120_ = ~new_n5116_ & ~new_n5119_;
  assign new_n5121_ = ~v16 & ~new_n5120_;
  assign new_n5122_ = ~v15 & new_n1108_;
  assign new_n5123_ = ~v14 & new_n5122_;
  assign new_n5124_ = ~new_n2325_ & ~new_n5123_;
  assign new_n5125_ = v40 & ~new_n5124_;
  assign new_n5126_ = ~v13 & new_n5125_;
  assign new_n5127_ = ~v5 & new_n5126_;
  assign new_n5128_ = ~v4 & new_n5127_;
  assign new_n5129_ = ~new_n5121_ & ~new_n5128_;
  assign new_n5130_ = ~v0 & ~new_n5129_;
  assign new_n5131_ = ~v5 & new_n1343_;
  assign new_n5132_ = new_n1010_ & new_n5131_;
  assign new_n5133_ = new_n268_ & new_n5132_;
  assign new_n5134_ = ~new_n5130_ & ~new_n5133_;
  assign new_n5135_ = ~v36 & ~new_n5134_;
  assign new_n5136_ = v12 & new_n5135_;
  assign new_n5137_ = ~v11 & new_n5136_;
  assign new_n5138_ = ~v10 & new_n5137_;
  assign new_n5139_ = ~v9 & new_n5138_;
  assign new_n5140_ = ~v8 & new_n5139_;
  assign new_n5141_ = ~v3 & new_n5140_;
  assign new_n5142_ = ~v2 & new_n5141_;
  assign \v41.68  = ~v1 & new_n5142_;
  assign new_n5144_ = v16 & new_n976_;
  assign new_n5145_ = v14 & new_n5144_;
  assign new_n5146_ = ~new_n915_ & ~new_n5145_;
  assign new_n5147_ = v40 & ~new_n5146_;
  assign new_n5148_ = ~v36 & new_n5147_;
  assign new_n5149_ = v15 & new_n5148_;
  assign new_n5150_ = v13 & new_n5149_;
  assign new_n5151_ = v12 & new_n5150_;
  assign new_n5152_ = ~v11 & new_n5151_;
  assign new_n5153_ = ~v10 & new_n5152_;
  assign new_n5154_ = ~v9 & new_n5153_;
  assign new_n5155_ = ~v8 & new_n5154_;
  assign new_n5156_ = ~v5 & new_n5155_;
  assign new_n5157_ = ~v4 & new_n5156_;
  assign new_n5158_ = ~v3 & new_n5157_;
  assign new_n5159_ = ~v2 & new_n5158_;
  assign new_n5160_ = ~v1 & new_n5159_;
  assign \v41.69  = ~v0 & new_n5160_;
  assign new_n5162_ = v14 & new_n4581_;
  assign new_n5163_ = v13 & new_n5162_;
  assign new_n5164_ = new_n201_ & new_n1343_;
  assign new_n5165_ = new_n754_ & new_n1365_;
  assign new_n5166_ = new_n5164_ & new_n5165_;
  assign new_n5167_ = ~new_n5163_ & ~new_n5166_;
  assign new_n5168_ = ~v5 & ~new_n5167_;
  assign new_n5169_ = ~new_n1362_ & ~new_n5168_;
  assign new_n5170_ = v19 & ~new_n5169_;
  assign new_n5171_ = v14 & new_n201_;
  assign new_n5172_ = new_n203_ & new_n5171_;
  assign new_n5173_ = ~new_n1796_ & ~new_n5172_;
  assign new_n5174_ = v13 & ~new_n5173_;
  assign new_n5175_ = ~v5 & new_n5174_;
  assign new_n5176_ = ~new_n5170_ & ~new_n5175_;
  assign new_n5177_ = v12 & ~new_n5176_;
  assign new_n5178_ = ~new_n4865_ & ~new_n5177_;
  assign new_n5179_ = v40 & ~new_n5178_;
  assign new_n5180_ = ~v3 & new_n5179_;
  assign new_n5181_ = new_n4858_ & ~new_n5180_;
  assign new_n5182_ = ~v36 & ~new_n5181_;
  assign new_n5183_ = ~v11 & new_n5182_;
  assign new_n5184_ = ~v10 & new_n5183_;
  assign new_n5185_ = ~v9 & new_n5184_;
  assign new_n5186_ = ~v8 & new_n5185_;
  assign new_n5187_ = ~v4 & new_n5186_;
  assign new_n5188_ = ~v2 & new_n5187_;
  assign new_n5189_ = ~v1 & new_n5188_;
  assign \v41.70  = ~v0 & new_n5189_;
  assign new_n5191_ = ~v18 & ~new_n1501_;
  assign new_n5192_ = ~v13 & new_n5191_;
  assign new_n5193_ = v12 & new_n5192_;
  assign new_n5194_ = new_n883_ & new_n2210_;
  assign new_n5195_ = ~new_n5193_ & ~new_n5194_;
  assign new_n5196_ = ~v19 & ~new_n5195_;
  assign new_n5197_ = new_n120_ & new_n259_;
  assign new_n5198_ = new_n2210_ & new_n5197_;
  assign new_n5199_ = ~new_n5196_ & ~new_n5198_;
  assign new_n5200_ = ~new_n843_ & ~new_n5199_;
  assign new_n5201_ = v19 & v39;
  assign new_n5202_ = new_n754_ & new_n5201_;
  assign new_n5203_ = new_n2006_ & new_n5202_;
  assign new_n5204_ = ~new_n5200_ & ~new_n5203_;
  assign new_n5205_ = v40 & ~new_n5204_;
  assign new_n5206_ = ~v14 & new_n5205_;
  assign new_n5207_ = v40 & ~new_n5206_;
  assign new_n5208_ = ~v36 & ~new_n5207_;
  assign new_n5209_ = ~v5 & new_n5208_;
  assign new_n5210_ = ~v4 & new_n5209_;
  assign new_n5211_ = ~v3 & new_n5210_;
  assign new_n5212_ = ~v2 & new_n5211_;
  assign new_n5213_ = ~v1 & new_n5212_;
  assign new_n5214_ = ~v0 & new_n5213_;
  assign new_n5215_ = ~v36 & ~new_n5214_;
  assign new_n5216_ = ~v10 & ~new_n5215_;
  assign new_n5217_ = ~v9 & new_n5216_;
  assign new_n5218_ = ~new_n1396_ & ~new_n5217_;
  assign new_n5219_ = ~v11 & ~new_n5218_;
  assign \v41.72  = ~v8 & new_n5219_;
  assign \v41.1  = 1'b0;
  assign \v41.31  = 1'b0;
  assign \v41.32  = 1'b0;
  assign \v41.39  = 1'b0;
endmodule


