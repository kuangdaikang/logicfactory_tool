// Benchmark "i10" written by ABC on Fri Feb 25 15:12:52 2022

module i10 ( 
    \V32(0) , \V32(1) , \V32(2) , \V32(3) , \V56(0) , \V289(0) , \V10(0) ,
    \V13(0) , \V35(0) , \V203(0) , \V288(6) , \V288(7) , \V248(0) ,
    \V249(0) , \V62(0) , \V59(0) , \V174(0) , \V215(0) , \V66(0) ,
    \V70(0) , \V43(0) , \V214(0) , \V37(0) , \V271(0) , \V40(0) , \V45(0) ,
    \V149(7) , \V149(6) , \V149(5) , \V149(4) , \V1(0) , \V7(0) , \V34(0) ,
    \V243(0) , \V244(0) , \V245(0) , \V246(0) , \V247(0) , \V293(0) ,
    \V302(0) , \V270(0) , \V269(0) , \V274(0) , \V202(0) , \V275(0) ,
    \V257(7) , \V257(5) , \V257(3) , \V257(1) , \V257(2) , \V257(4) ,
    \V257(6) , \V9(0) , \V149(0) , \V149(1) , \V149(2) , \V149(3) ,
    \V169(1) , \V165(0) , \V165(2) , \V165(4) , \V165(5) , \V165(6) ,
    \V165(7) , \V165(1) , \V88(2) , \V88(3) , \V55(0) , \V169(0) ,
    \V52(0) , \V5(0) , \V6(0) , \V12(0) , \V11(0) , \V4(0) , \V165(3) ,
    \V51(0) , \V65(0) , \V290(0) , \V279(0) , \V280(0) , \V288(4) ,
    \V288(2) , \V288(0) , \V258(0) , \V229(5) , \V229(4) , \V229(3) ,
    \V229(2) , \V229(1) , \V229(0) , \V223(5) , \V223(4) , \V223(3) ,
    \V223(2) , \V223(1) , \V223(0) , \V189(5) , \V189(4) , \V189(3) ,
    \V189(2) , \V189(1) , \V189(0) , \V183(5) , \V183(4) , \V183(3) ,
    \V183(2) , \V183(1) , \V183(0) , \V239(4) , \V239(3) , \V239(2) ,
    \V239(1) , \V239(0) , \V234(4) , \V234(3) , \V234(2) , \V234(1) ,
    \V234(0) , \V199(4) , \V199(3) , \V199(2) , \V199(1) , \V199(0) ,
    \V194(4) , \V194(3) , \V194(2) , \V194(1) , \V194(0) , \V257(0) ,
    \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(11) , \V32(10) ,
    \V32(9) , \V88(1) , \V88(0) , \V84(5) , \V84(4) , \V84(3) , \V84(2) ,
    \V84(1) , \V84(0) , \V78(5) , \V78(4) , \V2(0) , \V3(0) , \V14(0) ,
    \V213(0) , \V213(5) , \V213(4) , \V213(3) , \V213(2) , \V213(1) ,
    \V268(5) , \V268(3) , \V268(1) , \V268(2) , \V268(4) , \V8(0) ,
    \V60(0) , \V53(0) , \V57(0) , \V109(0) , \V277(0) , \V278(0) ,
    \V259(0) , \V260(0) , \V67(0) , \V68(0) , \V69(0) , \V216(0) ,
    \V175(0) , \V177(0) , \V172(0) , \V171(0) , \V50(0) , \V63(0) ,
    \V71(0) , \V292(0) , \V291(0) , \V91(0) , \V91(1) , \V294(0) ,
    \V207(0) , \V295(0) , \V204(0) , \V205(0) , \V261(0) , \V262(0) ,
    \V100(0) , \V100(5) , \V100(4) , \V100(3) , \V100(2) , \V100(1) ,
    \V240(0) , \V242(0) , \V241(0) , \V33(0) , \V16(0) , \V15(0) ,
    \V101(0) , \V268(0) , \V288(1) , \V288(3) , \V288(5) , \V301(0) ,
    \V108(0) , \V108(1) , \V108(2) , \V108(3) , \V108(4) , \V108(5) ,
    \V124(5) , \V124(4) , \V124(3) , \V124(2) , \V124(1) , \V124(0) ,
    \V132(7) , \V132(6) , \V132(5) , \V132(4) , \V132(3) , \V132(2) ,
    \V132(1) , \V132(0) , \V118(5) , \V118(4) , \V118(3) , \V118(2) ,
    \V118(1) , \V118(0) , \V118(7) , \V118(6) , \V46(0) , \V48(0) ,
    \V102(0) , \V110(0) , \V134(1) , \V134(0) , \V272(0) , \V78(2) ,
    \V78(3) , \V39(0) , \V38(0) , \V42(0) , \V44(0) , \V41(0) , \V78(1) ,
    \V78(0) , \V94(0) , \V94(1) ,
    \V321(2) , V356, V357, V373, \V375(0) , V377, \V393(0) , \V398(0) ,
    \V410(0) , \V423(0) , V432, \V435(0) , \V500(0) , \V508(0) , \V511(0) ,
    V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546,
    V547, V548, \V572(9) , \V572(8) , \V572(7) , \V572(6) , \V572(5) ,
    \V572(4) , \V572(3) , \V572(2) , \V572(1) , \V572(0) , \V585(0) , V587,
    \V591(0) , \V597(0) , \V603(0) , \V609(0) , V620, V621, V630,
    \V634(0) , \V640(0) , V657, V707, V763, V775, V778, V779, V780, V781,
    V782, V783, V784, V787, V789, \V798(0) , V801, \V802(0) , \V821(0) ,
    \V826(0) , V966, V986, \V1213(11) , \V1213(10) , \V1213(9) ,
    \V1213(8) , \V1213(7) , \V1213(6) , \V1213(5) , \V1213(4) , \V1213(3) ,
    \V1213(2) , \V1213(1) , \V1213(0) , \V1243(9) , \V1243(8) , \V1243(7) ,
    \V1243(6) , \V1243(5) , \V1243(4) , \V1243(3) , \V1243(2) , \V1243(1) ,
    \V1243(0) , V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263,
    V1264, V1265, V1266, V1267, \V1274(0) , \V1281(0) , \V1297(4) ,
    \V1297(3) , \V1297(2) , \V1297(1) , \V1297(0) , V1365, V1375, V1378,
    V1380, V1382, V1384, V1386, V1387, \V1392(0) , V1423, V1426, V1428,
    V1429, V1431, V1432, \V1439(0) , \V1440(0) , \V1451(0) , \V1459(0) ,
    \V1467(0) , V1470, \V1480(0) , \V1481(0) , \V1492(0) , \V1495(0) ,
    \V1512(3) , \V1512(2) , \V1512(1) , \V1536(0) , V1537, V1539,
    \V1552(1) , \V1552(0) , \V1613(0) , \V1613(1) , \V1620(0) , \V1629(0) ,
    \V1645(0) , \V1652(0) , V1669, \V1671(0) , \V1679(0) , \V1693(0) ,
    \V1709(4) , \V1709(3) , \V1709(2) , \V1709(1) , \V1709(0) , \V1717(0) ,
    V1719, \V1726(0) , V1736, \V1741(0) , \V1745(0) , \V1757(0) ,
    \V1758(0) , \V1759(0) , \V1760(0) , \V1771(1) , \V1771(0) , \V1781(1) ,
    \V1781(0) , \V1829(9) , \V1829(8) , \V1829(7) , \V1829(6) , \V1829(5) ,
    \V1829(4) , \V1829(3) , \V1829(2) , \V1829(1) , \V1829(0) , V1832,
    \V1833(0) , \V1863(0) , \V1864(0) , \V1896(0) , \V1897(0) , \V1898(0) ,
    \V1899(0) , \V1900(0) , \V1901(0) , \V1921(5) , \V1921(4) , \V1921(3) ,
    \V1921(2) , \V1921(1) , \V1921(0) , \V1953(1) , \V1953(7) , \V1953(6) ,
    \V1953(5) , \V1953(4) , \V1953(3) , \V1953(2) , \V1953(0) , \V1960(1) ,
    \V1960(0) , \V1968(0) , \V1992(1) , \V1992(0) , V650, V651, V652, V653,
    V654, V655, V656, V1370, V1371, V1372, V1373, V1374  );
  input  \V32(0) , \V32(1) , \V32(2) , \V32(3) , \V56(0) , \V289(0) ,
    \V10(0) , \V13(0) , \V35(0) , \V203(0) , \V288(6) , \V288(7) ,
    \V248(0) , \V249(0) , \V62(0) , \V59(0) , \V174(0) , \V215(0) ,
    \V66(0) , \V70(0) , \V43(0) , \V214(0) , \V37(0) , \V271(0) , \V40(0) ,
    \V45(0) , \V149(7) , \V149(6) , \V149(5) , \V149(4) , \V1(0) , \V7(0) ,
    \V34(0) , \V243(0) , \V244(0) , \V245(0) , \V246(0) , \V247(0) ,
    \V293(0) , \V302(0) , \V270(0) , \V269(0) , \V274(0) , \V202(0) ,
    \V275(0) , \V257(7) , \V257(5) , \V257(3) , \V257(1) , \V257(2) ,
    \V257(4) , \V257(6) , \V9(0) , \V149(0) , \V149(1) , \V149(2) ,
    \V149(3) , \V169(1) , \V165(0) , \V165(2) , \V165(4) , \V165(5) ,
    \V165(6) , \V165(7) , \V165(1) , \V88(2) , \V88(3) , \V55(0) ,
    \V169(0) , \V52(0) , \V5(0) , \V6(0) , \V12(0) , \V11(0) , \V4(0) ,
    \V165(3) , \V51(0) , \V65(0) , \V290(0) , \V279(0) , \V280(0) ,
    \V288(4) , \V288(2) , \V288(0) , \V258(0) , \V229(5) , \V229(4) ,
    \V229(3) , \V229(2) , \V229(1) , \V229(0) , \V223(5) , \V223(4) ,
    \V223(3) , \V223(2) , \V223(1) , \V223(0) , \V189(5) , \V189(4) ,
    \V189(3) , \V189(2) , \V189(1) , \V189(0) , \V183(5) , \V183(4) ,
    \V183(3) , \V183(2) , \V183(1) , \V183(0) , \V239(4) , \V239(3) ,
    \V239(2) , \V239(1) , \V239(0) , \V234(4) , \V234(3) , \V234(2) ,
    \V234(1) , \V234(0) , \V199(4) , \V199(3) , \V199(2) , \V199(1) ,
    \V199(0) , \V194(4) , \V194(3) , \V194(2) , \V194(1) , \V194(0) ,
    \V257(0) , \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(11) ,
    \V32(10) , \V32(9) , \V88(1) , \V88(0) , \V84(5) , \V84(4) , \V84(3) ,
    \V84(2) , \V84(1) , \V84(0) , \V78(5) , \V78(4) , \V2(0) , \V3(0) ,
    \V14(0) , \V213(0) , \V213(5) , \V213(4) , \V213(3) , \V213(2) ,
    \V213(1) , \V268(5) , \V268(3) , \V268(1) , \V268(2) , \V268(4) ,
    \V8(0) , \V60(0) , \V53(0) , \V57(0) , \V109(0) , \V277(0) , \V278(0) ,
    \V259(0) , \V260(0) , \V67(0) , \V68(0) , \V69(0) , \V216(0) ,
    \V175(0) , \V177(0) , \V172(0) , \V171(0) , \V50(0) , \V63(0) ,
    \V71(0) , \V292(0) , \V291(0) , \V91(0) , \V91(1) , \V294(0) ,
    \V207(0) , \V295(0) , \V204(0) , \V205(0) , \V261(0) , \V262(0) ,
    \V100(0) , \V100(5) , \V100(4) , \V100(3) , \V100(2) , \V100(1) ,
    \V240(0) , \V242(0) , \V241(0) , \V33(0) , \V16(0) , \V15(0) ,
    \V101(0) , \V268(0) , \V288(1) , \V288(3) , \V288(5) , \V301(0) ,
    \V108(0) , \V108(1) , \V108(2) , \V108(3) , \V108(4) , \V108(5) ,
    \V124(5) , \V124(4) , \V124(3) , \V124(2) , \V124(1) , \V124(0) ,
    \V132(7) , \V132(6) , \V132(5) , \V132(4) , \V132(3) , \V132(2) ,
    \V132(1) , \V132(0) , \V118(5) , \V118(4) , \V118(3) , \V118(2) ,
    \V118(1) , \V118(0) , \V118(7) , \V118(6) , \V46(0) , \V48(0) ,
    \V102(0) , \V110(0) , \V134(1) , \V134(0) , \V272(0) , \V78(2) ,
    \V78(3) , \V39(0) , \V38(0) , \V42(0) , \V44(0) , \V41(0) , \V78(1) ,
    \V78(0) , \V94(0) , \V94(1) ;
  output \V321(2) , V356, V357, V373, \V375(0) , V377, \V393(0) , \V398(0) ,
    \V410(0) , \V423(0) , V432, \V435(0) , \V500(0) , \V508(0) , \V511(0) ,
    V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546,
    V547, V548, \V572(9) , \V572(8) , \V572(7) , \V572(6) , \V572(5) ,
    \V572(4) , \V572(3) , \V572(2) , \V572(1) , \V572(0) , \V585(0) , V587,
    \V591(0) , \V597(0) , \V603(0) , \V609(0) , V620, V621, V630,
    \V634(0) , \V640(0) , V657, V707, V763, V775, V778, V779, V780, V781,
    V782, V783, V784, V787, V789, \V798(0) , V801, \V802(0) , \V821(0) ,
    \V826(0) , V966, V986, \V1213(11) , \V1213(10) , \V1213(9) ,
    \V1213(8) , \V1213(7) , \V1213(6) , \V1213(5) , \V1213(4) , \V1213(3) ,
    \V1213(2) , \V1213(1) , \V1213(0) , \V1243(9) , \V1243(8) , \V1243(7) ,
    \V1243(6) , \V1243(5) , \V1243(4) , \V1243(3) , \V1243(2) , \V1243(1) ,
    \V1243(0) , V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263,
    V1264, V1265, V1266, V1267, \V1274(0) , \V1281(0) , \V1297(4) ,
    \V1297(3) , \V1297(2) , \V1297(1) , \V1297(0) , V1365, V1375, V1378,
    V1380, V1382, V1384, V1386, V1387, \V1392(0) , V1423, V1426, V1428,
    V1429, V1431, V1432, \V1439(0) , \V1440(0) , \V1451(0) , \V1459(0) ,
    \V1467(0) , V1470, \V1480(0) , \V1481(0) , \V1492(0) , \V1495(0) ,
    \V1512(3) , \V1512(2) , \V1512(1) , \V1536(0) , V1537, V1539,
    \V1552(1) , \V1552(0) , \V1613(0) , \V1613(1) , \V1620(0) , \V1629(0) ,
    \V1645(0) , \V1652(0) , V1669, \V1671(0) , \V1679(0) , \V1693(0) ,
    \V1709(4) , \V1709(3) , \V1709(2) , \V1709(1) , \V1709(0) , \V1717(0) ,
    V1719, \V1726(0) , V1736, \V1741(0) , \V1745(0) , \V1757(0) ,
    \V1758(0) , \V1759(0) , \V1760(0) , \V1771(1) , \V1771(0) , \V1781(1) ,
    \V1781(0) , \V1829(9) , \V1829(8) , \V1829(7) , \V1829(6) , \V1829(5) ,
    \V1829(4) , \V1829(3) , \V1829(2) , \V1829(1) , \V1829(0) , V1832,
    \V1833(0) , \V1863(0) , \V1864(0) , \V1896(0) , \V1897(0) , \V1898(0) ,
    \V1899(0) , \V1900(0) , \V1901(0) , \V1921(5) , \V1921(4) , \V1921(3) ,
    \V1921(2) , \V1921(1) , \V1921(0) , \V1953(1) , \V1953(7) , \V1953(6) ,
    \V1953(5) , \V1953(4) , \V1953(3) , \V1953(2) , \V1953(0) , \V1960(1) ,
    \V1960(0) , \V1968(0) , \V1992(1) , \V1992(0) , V650, V651, V652, V653,
    V654, V655, V656, V1370, V1371, V1372, V1373, V1374;
  wire new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1279_, new_n1280_, new_n1281_, new_n1289_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1477_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1633_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_,
    new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_,
    new_n1724_, new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_,
    new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1750_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_,
    new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_,
    new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_,
    new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_,
    new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1899_, new_n1900_,
    new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_,
    new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_,
    new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_,
    new_n1919_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2044_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2139_,
    new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2161_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2195_,
    new_n2196_, new_n2197_, new_n2199_, new_n2200_, new_n2202_, new_n2203_,
    new_n2204_, new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_,
    new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_,
    new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_,
    new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_,
    new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_,
    new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_,
    new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_,
    new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2259_,
    new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2329_, new_n2330_, new_n2331_,
    new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_,
    new_n2338_, new_n2339_, new_n2342_, new_n2343_, new_n2344_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2363_, new_n2364_, new_n2365_, new_n2366_,
    new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_,
    new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_,
    new_n2387_, new_n2388_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_,
    new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_,
    new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2443_, new_n2444_,
    new_n2445_, new_n2446_, new_n2447_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2481_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_,
    new_n2494_, new_n2495_, new_n2496_, new_n2498_, new_n2499_, new_n2500_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2525_,
    new_n2527_, new_n2528_, new_n2531_, new_n2532_, new_n2533_, new_n2534_,
    new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_,
    new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_,
    new_n2548_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2558_, new_n2559_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2574_, new_n2575_, new_n2576_,
    new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_,
    new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_,
    new_n2589_, new_n2590_, new_n2592_, new_n2593_, new_n2594_, new_n2595_,
    new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2624_, new_n2626_, new_n2627_, new_n2629_, new_n2630_,
    new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2636_, new_n2637_,
    new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_,
    new_n2645_, new_n2646_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_,
    new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_,
    new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_,
    new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_,
    new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2790_, new_n2791_, new_n2792_,
    new_n2793_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2832_, new_n2833_,
    new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_,
    new_n2840_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_,
    new_n2847_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2872_, new_n2873_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2880_, new_n2881_, new_n2882_,
    new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_,
    new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_,
    new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_,
    new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_,
    new_n2921_, new_n2922_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2942_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2948_, new_n2949_,
    new_n2950_, new_n2951_, new_n2952_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2968_, new_n2969_, new_n2971_,
    new_n2972_, new_n2974_, new_n2976_, new_n2977_, new_n2978_, new_n2979_,
    new_n2980_, new_n2981_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2998_, new_n2999_, new_n3000_, new_n3001_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3008_, new_n3009_,
    new_n3010_, new_n3011_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3023_, new_n3024_,
    new_n3025_, new_n3026_, new_n3028_, new_n3029_, new_n3030_, new_n3031_,
    new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3038_, new_n3039_,
    new_n3040_, new_n3041_, new_n3043_, new_n3044_, new_n3045_, new_n3046_,
    new_n3048_, new_n3049_, new_n3051_, new_n3052_, new_n3053_, new_n3054_,
    new_n3056_, new_n3057_, new_n3058_, new_n3060_, new_n3061_, new_n3063_,
    new_n3064_, new_n3066_, new_n3067_, new_n3069_, new_n3071_, new_n3073_,
    new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_,
    new_n3080_, new_n3081_, new_n3083_, new_n3084_, new_n3085_, new_n3086_,
    new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_,
    new_n3107_, new_n3108_, new_n3109_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3127_, new_n3128_,
    new_n3129_, new_n3131_, new_n3132_, new_n3133_, new_n3135_, new_n3136_,
    new_n3138_, new_n3139_, new_n3141_, new_n3142_, new_n3143_, new_n3144_,
    new_n3146_, new_n3147_, new_n3148_, new_n3150_, new_n3151_, new_n3152_,
    new_n3154_, new_n3155_;
  assign new_n482_ = \V149(4)  & ~\V149(0) ;
  assign new_n483_ = \V149(1)  & new_n482_;
  assign new_n484_ = \V149(2)  & new_n483_;
  assign new_n485_ = ~\V149(3)  & new_n484_;
  assign new_n486_ = ~\V149(0)  & ~\V149(2) ;
  assign new_n487_ = ~\V149(1)  & new_n486_;
  assign new_n488_ = \V149(1)  & ~\V149(2) ;
  assign new_n489_ = ~\V149(0)  & new_n488_;
  assign new_n490_ = \V149(7)  & \V149(5) ;
  assign new_n491_ = ~\V149(3)  & new_n490_;
  assign new_n492_ = new_n489_ & new_n491_;
  assign new_n493_ = \V149(4)  & new_n492_;
  assign new_n494_ = \V149(6)  & new_n493_;
  assign new_n495_ = ~\V149(7)  & \V149(5) ;
  assign new_n496_ = ~\V149(3)  & new_n495_;
  assign new_n497_ = new_n489_ & new_n496_;
  assign new_n498_ = \V149(4)  & new_n497_;
  assign new_n499_ = \V149(6)  & new_n498_;
  assign new_n500_ = ~new_n494_ & ~new_n499_;
  assign \V802(0)  = \V52(0)  | \V51(0) ;
  assign new_n502_ = ~\V55(0)  & ~new_n500_;
  assign new_n503_ = ~\V802(0)  & new_n502_;
  assign new_n504_ = ~new_n485_ & ~new_n487_;
  assign new_n505_ = ~new_n503_ & new_n504_;
  assign new_n506_ = \V70(0)  & ~\V165(5) ;
  assign new_n507_ = \V165(3)  & new_n506_;
  assign new_n508_ = ~\V165(4)  & new_n507_;
  assign new_n509_ = ~\V165(6)  & new_n508_;
  assign new_n510_ = \V169(0)  & ~new_n505_;
  assign new_n511_ = ~\V291(0)  & new_n510_;
  assign new_n512_ = ~new_n509_ & new_n511_;
  assign V763 = ~\V292(0)  & new_n512_;
  assign new_n514_ = \V70(0)  & \V165(7) ;
  assign new_n515_ = \V261(0)  & new_n514_;
  assign new_n516_ = \V165(5)  & new_n515_;
  assign new_n517_ = \V165(3)  & new_n516_;
  assign new_n518_ = \V165(4)  & new_n517_;
  assign new_n519_ = \V165(6)  & new_n518_;
  assign new_n520_ = \V165(0)  & new_n519_;
  assign new_n521_ = \V165(1)  & new_n520_;
  assign new_n522_ = \V165(2)  & new_n521_;
  assign new_n523_ = V763 & new_n522_;
  assign new_n524_ = \V165(6)  & \V165(7) ;
  assign new_n525_ = \V165(5)  & new_n524_;
  assign new_n526_ = \V165(3)  & new_n525_;
  assign new_n527_ = \V165(4)  & new_n526_;
  assign new_n528_ = \V261(0)  & new_n527_;
  assign new_n529_ = ~\V204(0)  & new_n528_;
  assign new_n530_ = \V165(0)  & new_n529_;
  assign new_n531_ = \V165(1)  & new_n530_;
  assign new_n532_ = \V165(2)  & new_n531_;
  assign new_n533_ = ~new_n523_ & ~new_n532_;
  assign new_n534_ = ~\V262(0)  & new_n533_;
  assign new_n535_ = \V149(2)  & \V149(3) ;
  assign new_n536_ = \V149(1)  & new_n535_;
  assign new_n537_ = ~\V149(0)  & new_n536_;
  assign new_n538_ = ~\V174(0)  & new_n485_;
  assign new_n539_ = \V277(0)  & new_n538_;
  assign new_n540_ = \V278(0)  & ~new_n539_;
  assign new_n541_ = new_n537_ & ~new_n540_;
  assign new_n542_ = ~\V59(0)  & new_n541_;
  assign new_n543_ = ~\V149(1)  & \V149(2) ;
  assign new_n544_ = ~\V149(0)  & new_n543_;
  assign new_n545_ = ~new_n487_ & ~new_n544_;
  assign new_n546_ = ~\V149(4)  & ~\V149(0) ;
  assign new_n547_ = \V149(1)  & new_n546_;
  assign new_n548_ = \V149(2)  & new_n547_;
  assign new_n549_ = ~\V149(3)  & new_n548_;
  assign new_n550_ = ~new_n538_ & new_n545_;
  assign new_n551_ = ~new_n549_ & new_n550_;
  assign new_n552_ = ~\V174(0)  & ~new_n551_;
  assign new_n553_ = new_n537_ & new_n540_;
  assign new_n554_ = ~\V59(0)  & ~\V60(0) ;
  assign new_n555_ = new_n541_ & ~new_n554_;
  assign new_n556_ = ~new_n552_ & ~new_n553_;
  assign new_n557_ = ~new_n555_ & new_n556_;
  assign new_n558_ = \V257(7)  & ~new_n534_;
  assign new_n559_ = ~new_n542_ & new_n558_;
  assign new_n560_ = new_n557_ & new_n559_;
  assign new_n561_ = ~\V59(0)  & \V149(4) ;
  assign new_n562_ = ~new_n540_ & new_n561_;
  assign new_n563_ = new_n537_ & new_n562_;
  assign new_n564_ = new_n534_ & new_n563_;
  assign new_n565_ = new_n557_ & new_n564_;
  assign new_n566_ = ~new_n537_ & ~new_n538_;
  assign new_n567_ = ~new_n549_ & new_n566_;
  assign new_n568_ = \V234(0)  & ~new_n545_;
  assign new_n569_ = new_n567_ & new_n568_;
  assign new_n570_ = \V194(0)  & new_n545_;
  assign new_n571_ = ~new_n567_ & new_n570_;
  assign new_n572_ = ~new_n569_ & ~new_n571_;
  assign new_n573_ = new_n534_ & ~new_n572_;
  assign new_n574_ = ~new_n542_ & new_n573_;
  assign new_n575_ = ~new_n557_ & new_n574_;
  assign new_n576_ = ~new_n560_ & ~new_n565_;
  assign new_n577_ = ~new_n575_ & new_n576_;
  assign new_n578_ = V763 & new_n534_;
  assign new_n579_ = ~new_n577_ & ~new_n578_;
  assign new_n580_ = ~new_n578_ & new_n579_;
  assign new_n581_ = ~\V56(0)  & ~\V59(0) ;
  assign new_n582_ = ~\V60(0)  & new_n581_;
  assign new_n583_ = V763 & ~new_n582_;
  assign new_n584_ = \V32(2)  & new_n583_;
  assign new_n585_ = \V32(5)  & ~new_n583_;
  assign new_n586_ = ~new_n583_ & new_n585_;
  assign new_n587_ = ~new_n584_ & ~new_n586_;
  assign new_n588_ = new_n578_ & ~new_n587_;
  assign new_n589_ = new_n578_ & new_n588_;
  assign new_n590_ = ~new_n580_ & ~new_n589_;
  assign new_n591_ = \V149(3)  & new_n544_;
  assign new_n592_ = ~new_n538_ & ~new_n591_;
  assign new_n593_ = \V60(0)  & ~new_n592_;
  assign new_n594_ = \V149(7)  & ~\V149(5) ;
  assign new_n595_ = ~\V149(3)  & new_n594_;
  assign new_n596_ = new_n489_ & new_n595_;
  assign new_n597_ = \V149(4)  & new_n596_;
  assign new_n598_ = \V149(6)  & new_n597_;
  assign new_n599_ = ~\V174(0)  & new_n487_;
  assign new_n600_ = ~\V149(4)  & ~\V149(3) ;
  assign new_n601_ = new_n599_ & new_n600_;
  assign new_n602_ = \V149(5)  & new_n601_;
  assign new_n603_ = \V88(2)  & new_n602_;
  assign new_n604_ = ~\V88(3)  & new_n603_;
  assign new_n605_ = ~\V88(2)  & new_n602_;
  assign new_n606_ = ~\V88(3)  & new_n605_;
  assign V707 = ~\V149(3)  & new_n599_;
  assign new_n608_ = ~\V149(5)  & ~\V149(4) ;
  assign new_n609_ = V707 & new_n608_;
  assign new_n610_ = \V88(2)  & new_n609_;
  assign new_n611_ = ~\V88(3)  & new_n610_;
  assign new_n612_ = \V149(5)  & V707;
  assign new_n613_ = \V149(4)  & new_n612_;
  assign new_n614_ = ~\V149(5)  & V707;
  assign new_n615_ = \V149(4)  & new_n614_;
  assign new_n616_ = ~\V88(2)  & new_n609_;
  assign new_n617_ = \V88(3)  & new_n616_;
  assign new_n618_ = \V88(3)  & new_n610_;
  assign new_n619_ = \V88(3)  & new_n605_;
  assign new_n620_ = ~new_n611_ & ~new_n613_;
  assign new_n621_ = ~new_n604_ & ~new_n606_;
  assign new_n622_ = new_n620_ & new_n621_;
  assign new_n623_ = ~new_n618_ & ~new_n619_;
  assign new_n624_ = ~new_n615_ & ~new_n617_;
  assign new_n625_ = new_n623_ & new_n624_;
  assign new_n626_ = new_n622_ & new_n625_;
  assign new_n627_ = \V169(1)  & ~new_n545_;
  assign new_n628_ = ~new_n626_ & new_n627_;
  assign new_n629_ = \V60(0)  & new_n628_;
  assign new_n630_ = \V149(3)  & new_n599_;
  assign new_n631_ = new_n627_ & new_n630_;
  assign new_n632_ = \V60(0)  & new_n631_;
  assign new_n633_ = \V56(0)  & new_n631_;
  assign new_n634_ = \V56(0)  & new_n628_;
  assign new_n635_ = ~new_n633_ & ~new_n634_;
  assign new_n636_ = ~new_n629_ & ~new_n632_;
  assign new_n637_ = new_n635_ & new_n636_;
  assign new_n638_ = new_n538_ & ~new_n540_;
  assign new_n639_ = ~\V149(5)  & ~\V149(3) ;
  assign new_n640_ = new_n544_ & new_n639_;
  assign new_n641_ = \V149(4)  & new_n640_;
  assign new_n642_ = ~\V149(4)  & new_n640_;
  assign new_n643_ = \V149(5)  & ~\V149(3) ;
  assign new_n644_ = new_n544_ & new_n643_;
  assign new_n645_ = ~\V149(4)  & new_n644_;
  assign new_n646_ = ~new_n641_ & ~new_n642_;
  assign new_n647_ = ~new_n645_ & new_n646_;
  assign new_n648_ = ~new_n591_ & new_n626_;
  assign new_n649_ = ~new_n638_ & new_n647_;
  assign new_n650_ = ~new_n630_ & new_n649_;
  assign new_n651_ = new_n648_ & new_n650_;
  assign new_n652_ = ~\V56(0)  & ~\V53(0) ;
  assign new_n653_ = ~\V57(0)  & new_n652_;
  assign new_n654_ = new_n637_ & ~new_n651_;
  assign new_n655_ = ~new_n653_ & new_n654_;
  assign new_n656_ = new_n534_ & ~new_n549_;
  assign new_n657_ = ~new_n537_ & new_n656_;
  assign new_n658_ = \V53(0)  & new_n657_;
  assign new_n659_ = ~\V56(0)  & new_n658_;
  assign new_n660_ = ~new_n598_ & ~new_n655_;
  assign new_n661_ = ~new_n659_ & new_n660_;
  assign new_n662_ = ~new_n593_ & ~new_n661_;
  assign new_n663_ = ~new_n590_ & ~new_n662_;
  assign new_n664_ = new_n661_ & new_n663_;
  assign new_n665_ = \V78(4)  & new_n662_;
  assign new_n666_ = ~new_n661_ & new_n665_;
  assign \V321(2)  = ~new_n664_ & ~new_n666_;
  assign new_n668_ = ~\V149(7)  & ~\V149(5) ;
  assign new_n669_ = \V149(3)  & new_n668_;
  assign new_n670_ = new_n489_ & new_n669_;
  assign new_n671_ = ~\V149(4)  & new_n670_;
  assign new_n672_ = ~\V149(6)  & new_n671_;
  assign new_n673_ = ~\V802(0)  & new_n672_;
  assign new_n674_ = new_n534_ & ~new_n673_;
  assign new_n675_ = ~\V288(0)  & \V288(1) ;
  assign new_n676_ = ~\V288(2)  & \V288(3) ;
  assign new_n677_ = ~\V288(4)  & \V288(5) ;
  assign new_n678_ = ~\V288(6)  & \V288(7) ;
  assign new_n679_ = new_n677_ & new_n678_;
  assign new_n680_ = ~new_n677_ & ~new_n678_;
  assign new_n681_ = ~new_n679_ & ~new_n680_;
  assign new_n682_ = new_n676_ & new_n681_;
  assign new_n683_ = ~new_n676_ & ~new_n681_;
  assign new_n684_ = ~new_n682_ & ~new_n683_;
  assign new_n685_ = new_n675_ & new_n684_;
  assign new_n686_ = ~new_n675_ & ~new_n684_;
  assign new_n687_ = ~new_n685_ & ~new_n686_;
  assign new_n688_ = new_n675_ & ~new_n687_;
  assign new_n689_ = new_n675_ & new_n688_;
  assign new_n690_ = \V288(0)  & ~\V288(1) ;
  assign new_n691_ = ~new_n687_ & new_n690_;
  assign new_n692_ = new_n690_ & new_n691_;
  assign new_n693_ = ~new_n687_ & ~new_n690_;
  assign new_n694_ = ~new_n690_ & new_n693_;
  assign new_n695_ = ~new_n692_ & ~new_n694_;
  assign new_n696_ = ~new_n675_ & new_n695_;
  assign new_n697_ = ~new_n675_ & new_n696_;
  assign new_n698_ = ~new_n689_ & ~new_n697_;
  assign new_n699_ = \V223(3)  & ~new_n545_;
  assign new_n700_ = new_n567_ & new_n699_;
  assign new_n701_ = \V183(3)  & new_n545_;
  assign new_n702_ = ~new_n567_ & new_n701_;
  assign new_n703_ = ~new_n700_ & ~new_n702_;
  assign new_n704_ = ~new_n557_ & ~new_n578_;
  assign new_n705_ = ~new_n703_ & new_n704_;
  assign new_n706_ = new_n534_ & new_n705_;
  assign new_n707_ = ~new_n542_ & new_n706_;
  assign new_n708_ = ~new_n578_ & new_n707_;
  assign new_n709_ = ~new_n662_ & new_n708_;
  assign new_n710_ = new_n661_ & new_n709_;
  assign new_n711_ = \V32(3)  & new_n662_;
  assign new_n712_ = ~new_n661_ & new_n711_;
  assign \V1213(3)  = new_n710_ | new_n712_;
  assign new_n714_ = ~new_n698_ & ~\V1213(3) ;
  assign new_n715_ = new_n698_ & \V1213(3) ;
  assign new_n716_ = ~new_n714_ & ~new_n715_;
  assign new_n717_ = \V288(2)  & ~\V288(3) ;
  assign new_n718_ = \V288(4)  & ~\V288(5) ;
  assign new_n719_ = \V288(6)  & ~\V288(7) ;
  assign new_n720_ = ~new_n678_ & ~new_n719_;
  assign new_n721_ = new_n718_ & ~new_n720_;
  assign new_n722_ = ~new_n718_ & new_n720_;
  assign new_n723_ = ~new_n721_ & ~new_n722_;
  assign new_n724_ = new_n677_ & ~new_n678_;
  assign new_n725_ = ~new_n723_ & ~new_n724_;
  assign new_n726_ = new_n723_ & new_n724_;
  assign new_n727_ = ~new_n725_ & ~new_n726_;
  assign new_n728_ = new_n717_ & new_n727_;
  assign new_n729_ = ~new_n717_ & ~new_n727_;
  assign new_n730_ = ~new_n728_ & ~new_n729_;
  assign new_n731_ = new_n676_ & ~new_n681_;
  assign new_n732_ = ~new_n730_ & ~new_n731_;
  assign new_n733_ = new_n730_ & new_n731_;
  assign new_n734_ = ~new_n732_ & ~new_n733_;
  assign new_n735_ = new_n690_ & ~new_n734_;
  assign new_n736_ = new_n675_ & ~new_n684_;
  assign new_n737_ = new_n690_ & new_n736_;
  assign new_n738_ = ~new_n734_ & new_n736_;
  assign new_n739_ = ~new_n735_ & ~new_n737_;
  assign new_n740_ = ~new_n738_ & new_n739_;
  assign new_n741_ = \V288(0)  & \V288(1) ;
  assign new_n742_ = new_n717_ & ~new_n727_;
  assign new_n743_ = new_n717_ & new_n731_;
  assign new_n744_ = ~new_n727_ & new_n731_;
  assign new_n745_ = ~new_n742_ & ~new_n743_;
  assign new_n746_ = ~new_n744_ & new_n745_;
  assign new_n747_ = \V288(2)  & \V288(3) ;
  assign new_n748_ = new_n718_ & new_n720_;
  assign new_n749_ = new_n718_ & new_n724_;
  assign new_n750_ = new_n720_ & new_n724_;
  assign new_n751_ = ~new_n748_ & ~new_n749_;
  assign new_n752_ = ~new_n750_ & new_n751_;
  assign new_n753_ = \V288(4)  & \V288(5) ;
  assign new_n754_ = ~\V288(6)  & ~\V288(7) ;
  assign new_n755_ = new_n753_ & ~new_n754_;
  assign new_n756_ = ~new_n753_ & new_n754_;
  assign new_n757_ = ~new_n755_ & ~new_n756_;
  assign new_n758_ = ~new_n752_ & new_n757_;
  assign new_n759_ = new_n752_ & ~new_n757_;
  assign new_n760_ = ~new_n758_ & ~new_n759_;
  assign new_n761_ = new_n747_ & new_n760_;
  assign new_n762_ = ~new_n747_ & ~new_n760_;
  assign new_n763_ = ~new_n761_ & ~new_n762_;
  assign new_n764_ = ~new_n746_ & new_n763_;
  assign new_n765_ = new_n746_ & ~new_n763_;
  assign new_n766_ = ~new_n764_ & ~new_n765_;
  assign new_n767_ = new_n741_ & new_n766_;
  assign new_n768_ = ~new_n741_ & ~new_n766_;
  assign new_n769_ = ~new_n767_ & ~new_n768_;
  assign new_n770_ = ~new_n740_ & new_n769_;
  assign new_n771_ = new_n740_ & ~new_n769_;
  assign new_n772_ = ~new_n770_ & ~new_n771_;
  assign new_n773_ = new_n675_ & ~new_n772_;
  assign new_n774_ = new_n675_ & new_n773_;
  assign new_n775_ = new_n690_ & ~new_n772_;
  assign new_n776_ = new_n690_ & new_n775_;
  assign new_n777_ = new_n690_ & new_n734_;
  assign new_n778_ = ~new_n690_ & ~new_n734_;
  assign new_n779_ = ~new_n777_ & ~new_n778_;
  assign new_n780_ = ~new_n736_ & ~new_n779_;
  assign new_n781_ = new_n736_ & new_n779_;
  assign new_n782_ = ~new_n780_ & ~new_n781_;
  assign new_n783_ = new_n687_ & new_n782_;
  assign new_n784_ = ~new_n772_ & ~new_n783_;
  assign new_n785_ = new_n772_ & new_n783_;
  assign new_n786_ = ~new_n784_ & ~new_n785_;
  assign new_n787_ = ~new_n687_ & ~new_n782_;
  assign new_n788_ = ~new_n783_ & ~new_n787_;
  assign new_n789_ = ~new_n687_ & new_n788_;
  assign new_n790_ = ~new_n786_ & ~new_n789_;
  assign new_n791_ = new_n786_ & new_n789_;
  assign new_n792_ = ~new_n790_ & ~new_n791_;
  assign new_n793_ = ~new_n690_ & ~new_n792_;
  assign new_n794_ = ~new_n690_ & new_n793_;
  assign new_n795_ = ~new_n776_ & ~new_n794_;
  assign new_n796_ = new_n690_ & ~new_n782_;
  assign new_n797_ = new_n690_ & new_n796_;
  assign new_n798_ = new_n687_ & ~new_n788_;
  assign new_n799_ = ~new_n789_ & ~new_n798_;
  assign new_n800_ = ~new_n690_ & ~new_n799_;
  assign new_n801_ = ~new_n690_ & new_n800_;
  assign new_n802_ = ~new_n797_ & ~new_n801_;
  assign new_n803_ = new_n695_ & new_n802_;
  assign new_n804_ = ~new_n795_ & ~new_n803_;
  assign new_n805_ = new_n795_ & new_n803_;
  assign new_n806_ = ~new_n804_ & ~new_n805_;
  assign new_n807_ = ~new_n675_ & ~new_n806_;
  assign new_n808_ = ~new_n675_ & new_n807_;
  assign new_n809_ = ~new_n774_ & ~new_n808_;
  assign new_n810_ = \V223(1)  & ~new_n545_;
  assign new_n811_ = new_n567_ & new_n810_;
  assign new_n812_ = \V183(1)  & new_n545_;
  assign new_n813_ = ~new_n567_ & new_n812_;
  assign new_n814_ = ~new_n811_ & ~new_n813_;
  assign new_n815_ = new_n704_ & ~new_n814_;
  assign new_n816_ = new_n534_ & new_n815_;
  assign new_n817_ = ~new_n542_ & new_n816_;
  assign new_n818_ = ~new_n578_ & new_n817_;
  assign new_n819_ = ~new_n662_ & new_n818_;
  assign new_n820_ = new_n661_ & new_n819_;
  assign new_n821_ = \V32(1)  & new_n662_;
  assign new_n822_ = ~new_n661_ & new_n821_;
  assign \V1213(1)  = new_n820_ | new_n822_;
  assign new_n824_ = ~new_n809_ & ~\V1213(1) ;
  assign new_n825_ = new_n809_ & \V1213(1) ;
  assign new_n826_ = ~new_n824_ & ~new_n825_;
  assign new_n827_ = new_n753_ & new_n754_;
  assign new_n828_ = ~new_n752_ & new_n753_;
  assign new_n829_ = ~new_n752_ & new_n754_;
  assign new_n830_ = ~new_n827_ & ~new_n828_;
  assign new_n831_ = ~new_n829_ & new_n830_;
  assign new_n832_ = new_n754_ & new_n831_;
  assign new_n833_ = ~new_n754_ & ~new_n831_;
  assign new_n834_ = ~new_n832_ & ~new_n833_;
  assign new_n835_ = new_n747_ & ~new_n760_;
  assign new_n836_ = ~new_n746_ & new_n747_;
  assign new_n837_ = ~new_n746_ & ~new_n760_;
  assign new_n838_ = ~new_n835_ & ~new_n836_;
  assign new_n839_ = ~new_n837_ & new_n838_;
  assign new_n840_ = ~new_n834_ & new_n839_;
  assign new_n841_ = new_n834_ & ~new_n839_;
  assign new_n842_ = ~new_n840_ & ~new_n841_;
  assign new_n843_ = new_n741_ & ~new_n766_;
  assign new_n844_ = ~new_n740_ & new_n741_;
  assign new_n845_ = ~new_n740_ & ~new_n766_;
  assign new_n846_ = ~new_n843_ & ~new_n844_;
  assign new_n847_ = ~new_n845_ & new_n846_;
  assign new_n848_ = ~new_n842_ & new_n847_;
  assign new_n849_ = new_n842_ & ~new_n847_;
  assign new_n850_ = ~new_n848_ & ~new_n849_;
  assign new_n851_ = new_n675_ & ~new_n850_;
  assign new_n852_ = new_n675_ & new_n851_;
  assign new_n853_ = new_n690_ & ~new_n850_;
  assign new_n854_ = new_n690_ & new_n853_;
  assign new_n855_ = ~new_n785_ & ~new_n850_;
  assign new_n856_ = new_n785_ & new_n850_;
  assign new_n857_ = ~new_n855_ & ~new_n856_;
  assign new_n858_ = ~new_n791_ & ~new_n857_;
  assign new_n859_ = new_n791_ & new_n857_;
  assign new_n860_ = ~new_n858_ & ~new_n859_;
  assign new_n861_ = ~new_n690_ & ~new_n860_;
  assign new_n862_ = ~new_n690_ & new_n861_;
  assign new_n863_ = ~new_n854_ & ~new_n862_;
  assign new_n864_ = ~new_n805_ & ~new_n863_;
  assign new_n865_ = new_n805_ & new_n863_;
  assign new_n866_ = ~new_n864_ & ~new_n865_;
  assign new_n867_ = ~new_n675_ & ~new_n866_;
  assign new_n868_ = ~new_n675_ & new_n867_;
  assign new_n869_ = ~new_n852_ & ~new_n868_;
  assign new_n870_ = \V223(0)  & ~new_n545_;
  assign new_n871_ = new_n567_ & new_n870_;
  assign new_n872_ = \V183(0)  & new_n545_;
  assign new_n873_ = ~new_n567_ & new_n872_;
  assign new_n874_ = ~new_n871_ & ~new_n873_;
  assign new_n875_ = new_n704_ & ~new_n874_;
  assign new_n876_ = new_n534_ & new_n875_;
  assign new_n877_ = ~new_n542_ & new_n876_;
  assign new_n878_ = ~new_n578_ & new_n877_;
  assign new_n879_ = ~new_n662_ & new_n878_;
  assign new_n880_ = new_n661_ & new_n879_;
  assign new_n881_ = \V32(0)  & new_n662_;
  assign new_n882_ = ~new_n661_ & new_n881_;
  assign \V1213(0)  = new_n880_ | new_n882_;
  assign new_n884_ = ~new_n869_ & ~\V1213(0) ;
  assign new_n885_ = new_n869_ & \V1213(0) ;
  assign new_n886_ = ~new_n884_ & ~new_n885_;
  assign new_n887_ = new_n675_ & ~new_n782_;
  assign new_n888_ = new_n675_ & new_n887_;
  assign new_n889_ = ~new_n695_ & ~new_n802_;
  assign new_n890_ = ~new_n803_ & ~new_n889_;
  assign new_n891_ = ~new_n675_ & ~new_n890_;
  assign new_n892_ = ~new_n675_ & new_n891_;
  assign new_n893_ = ~new_n888_ & ~new_n892_;
  assign new_n894_ = \V223(2)  & ~new_n545_;
  assign new_n895_ = new_n567_ & new_n894_;
  assign new_n896_ = \V183(2)  & new_n545_;
  assign new_n897_ = ~new_n567_ & new_n896_;
  assign new_n898_ = ~new_n895_ & ~new_n897_;
  assign new_n899_ = new_n704_ & ~new_n898_;
  assign new_n900_ = new_n534_ & new_n899_;
  assign new_n901_ = ~new_n542_ & new_n900_;
  assign new_n902_ = ~new_n578_ & new_n901_;
  assign new_n903_ = ~new_n662_ & new_n902_;
  assign new_n904_ = new_n661_ & new_n903_;
  assign new_n905_ = \V32(2)  & new_n662_;
  assign new_n906_ = ~new_n661_ & new_n905_;
  assign \V1213(2)  = new_n904_ | new_n906_;
  assign new_n908_ = ~new_n893_ & ~\V1213(2) ;
  assign new_n909_ = new_n893_ & \V1213(2) ;
  assign new_n910_ = ~new_n908_ & ~new_n909_;
  assign new_n911_ = ~\V288(0)  & ~\V288(1) ;
  assign new_n912_ = ~new_n673_ & new_n716_;
  assign new_n913_ = new_n826_ & new_n912_;
  assign new_n914_ = new_n886_ & new_n913_;
  assign new_n915_ = new_n910_ & new_n914_;
  assign new_n916_ = ~new_n911_ & new_n915_;
  assign new_n917_ = new_n676_ & ~new_n684_;
  assign new_n918_ = new_n676_ & new_n917_;
  assign new_n919_ = ~new_n684_ & new_n717_;
  assign new_n920_ = new_n717_ & new_n919_;
  assign new_n921_ = ~new_n684_ & ~new_n717_;
  assign new_n922_ = ~new_n717_ & new_n921_;
  assign new_n923_ = ~new_n920_ & ~new_n922_;
  assign new_n924_ = ~new_n676_ & new_n923_;
  assign new_n925_ = ~new_n676_ & new_n924_;
  assign new_n926_ = ~new_n918_ & ~new_n925_;
  assign new_n927_ = ~\V1213(3)  & ~new_n926_;
  assign new_n928_ = \V1213(3)  & new_n926_;
  assign new_n929_ = ~new_n927_ & ~new_n928_;
  assign new_n930_ = new_n676_ & ~new_n766_;
  assign new_n931_ = new_n676_ & new_n930_;
  assign new_n932_ = new_n717_ & ~new_n766_;
  assign new_n933_ = new_n717_ & new_n932_;
  assign new_n934_ = new_n684_ & new_n734_;
  assign new_n935_ = ~new_n766_ & ~new_n934_;
  assign new_n936_ = new_n766_ & new_n934_;
  assign new_n937_ = ~new_n935_ & ~new_n936_;
  assign new_n938_ = ~new_n684_ & ~new_n734_;
  assign new_n939_ = ~new_n934_ & ~new_n938_;
  assign new_n940_ = ~new_n684_ & new_n939_;
  assign new_n941_ = ~new_n937_ & ~new_n940_;
  assign new_n942_ = new_n937_ & new_n940_;
  assign new_n943_ = ~new_n941_ & ~new_n942_;
  assign new_n944_ = ~new_n717_ & ~new_n943_;
  assign new_n945_ = ~new_n717_ & new_n944_;
  assign new_n946_ = ~new_n933_ & ~new_n945_;
  assign new_n947_ = new_n717_ & ~new_n734_;
  assign new_n948_ = new_n717_ & new_n947_;
  assign new_n949_ = new_n684_ & ~new_n939_;
  assign new_n950_ = ~new_n940_ & ~new_n949_;
  assign new_n951_ = ~new_n717_ & ~new_n950_;
  assign new_n952_ = ~new_n717_ & new_n951_;
  assign new_n953_ = ~new_n948_ & ~new_n952_;
  assign new_n954_ = new_n923_ & new_n953_;
  assign new_n955_ = ~new_n946_ & ~new_n954_;
  assign new_n956_ = new_n946_ & new_n954_;
  assign new_n957_ = ~new_n955_ & ~new_n956_;
  assign new_n958_ = ~new_n676_ & ~new_n957_;
  assign new_n959_ = ~new_n676_ & new_n958_;
  assign new_n960_ = ~new_n931_ & ~new_n959_;
  assign new_n961_ = ~\V1213(1)  & ~new_n960_;
  assign new_n962_ = \V1213(1)  & new_n960_;
  assign new_n963_ = ~new_n961_ & ~new_n962_;
  assign new_n964_ = new_n676_ & ~new_n842_;
  assign new_n965_ = new_n676_ & new_n964_;
  assign new_n966_ = new_n717_ & ~new_n842_;
  assign new_n967_ = new_n717_ & new_n966_;
  assign new_n968_ = ~new_n842_ & ~new_n936_;
  assign new_n969_ = new_n842_ & new_n936_;
  assign new_n970_ = ~new_n968_ & ~new_n969_;
  assign new_n971_ = ~new_n942_ & ~new_n970_;
  assign new_n972_ = new_n942_ & new_n970_;
  assign new_n973_ = ~new_n971_ & ~new_n972_;
  assign new_n974_ = ~new_n717_ & ~new_n973_;
  assign new_n975_ = ~new_n717_ & new_n974_;
  assign new_n976_ = ~new_n967_ & ~new_n975_;
  assign new_n977_ = ~new_n956_ & ~new_n976_;
  assign new_n978_ = new_n956_ & new_n976_;
  assign new_n979_ = ~new_n977_ & ~new_n978_;
  assign new_n980_ = ~new_n676_ & ~new_n979_;
  assign new_n981_ = ~new_n676_ & new_n980_;
  assign new_n982_ = ~new_n965_ & ~new_n981_;
  assign new_n983_ = ~\V1213(0)  & ~new_n982_;
  assign new_n984_ = \V1213(0)  & new_n982_;
  assign new_n985_ = ~new_n983_ & ~new_n984_;
  assign new_n986_ = new_n676_ & ~new_n734_;
  assign new_n987_ = new_n676_ & new_n986_;
  assign new_n988_ = ~new_n923_ & ~new_n953_;
  assign new_n989_ = ~new_n954_ & ~new_n988_;
  assign new_n990_ = ~new_n676_ & ~new_n989_;
  assign new_n991_ = ~new_n676_ & new_n990_;
  assign new_n992_ = ~new_n987_ & ~new_n991_;
  assign new_n993_ = ~\V1213(2)  & ~new_n992_;
  assign new_n994_ = \V1213(2)  & new_n992_;
  assign new_n995_ = ~new_n993_ & ~new_n994_;
  assign new_n996_ = ~\V288(2)  & ~\V288(3) ;
  assign new_n997_ = ~new_n673_ & new_n929_;
  assign new_n998_ = new_n963_ & new_n997_;
  assign new_n999_ = new_n985_ & new_n998_;
  assign new_n1000_ = new_n995_ & new_n999_;
  assign new_n1001_ = ~new_n996_ & new_n1000_;
  assign new_n1002_ = new_n677_ & ~new_n681_;
  assign new_n1003_ = new_n677_ & new_n1002_;
  assign new_n1004_ = ~new_n681_ & new_n718_;
  assign new_n1005_ = new_n718_ & new_n1004_;
  assign new_n1006_ = ~new_n681_ & ~new_n718_;
  assign new_n1007_ = ~new_n718_ & new_n1006_;
  assign new_n1008_ = ~new_n1005_ & ~new_n1007_;
  assign new_n1009_ = ~new_n677_ & new_n1008_;
  assign new_n1010_ = ~new_n677_ & new_n1009_;
  assign new_n1011_ = ~new_n1003_ & ~new_n1010_;
  assign new_n1012_ = ~\V1213(3)  & ~new_n1011_;
  assign new_n1013_ = \V1213(3)  & new_n1011_;
  assign new_n1014_ = ~new_n1012_ & ~new_n1013_;
  assign new_n1015_ = new_n677_ & ~new_n760_;
  assign new_n1016_ = new_n677_ & new_n1015_;
  assign new_n1017_ = new_n718_ & ~new_n760_;
  assign new_n1018_ = new_n718_ & new_n1017_;
  assign new_n1019_ = new_n681_ & new_n727_;
  assign new_n1020_ = ~new_n760_ & ~new_n1019_;
  assign new_n1021_ = new_n760_ & new_n1019_;
  assign new_n1022_ = ~new_n1020_ & ~new_n1021_;
  assign new_n1023_ = ~new_n681_ & ~new_n727_;
  assign new_n1024_ = ~new_n1019_ & ~new_n1023_;
  assign new_n1025_ = ~new_n681_ & new_n1024_;
  assign new_n1026_ = ~new_n1022_ & ~new_n1025_;
  assign new_n1027_ = new_n1022_ & new_n1025_;
  assign new_n1028_ = ~new_n1026_ & ~new_n1027_;
  assign new_n1029_ = ~new_n718_ & ~new_n1028_;
  assign new_n1030_ = ~new_n718_ & new_n1029_;
  assign new_n1031_ = ~new_n1018_ & ~new_n1030_;
  assign new_n1032_ = new_n718_ & ~new_n727_;
  assign new_n1033_ = new_n718_ & new_n1032_;
  assign new_n1034_ = new_n681_ & ~new_n1024_;
  assign new_n1035_ = ~new_n1025_ & ~new_n1034_;
  assign new_n1036_ = ~new_n718_ & ~new_n1035_;
  assign new_n1037_ = ~new_n718_ & new_n1036_;
  assign new_n1038_ = ~new_n1033_ & ~new_n1037_;
  assign new_n1039_ = new_n1008_ & new_n1038_;
  assign new_n1040_ = ~new_n1031_ & ~new_n1039_;
  assign new_n1041_ = new_n1031_ & new_n1039_;
  assign new_n1042_ = ~new_n1040_ & ~new_n1041_;
  assign new_n1043_ = ~new_n677_ & ~new_n1042_;
  assign new_n1044_ = ~new_n677_ & new_n1043_;
  assign new_n1045_ = ~new_n1016_ & ~new_n1044_;
  assign new_n1046_ = ~\V1213(1)  & ~new_n1045_;
  assign new_n1047_ = \V1213(1)  & new_n1045_;
  assign new_n1048_ = ~new_n1046_ & ~new_n1047_;
  assign new_n1049_ = new_n677_ & ~new_n834_;
  assign new_n1050_ = new_n677_ & new_n1049_;
  assign new_n1051_ = new_n718_ & ~new_n834_;
  assign new_n1052_ = new_n718_ & new_n1051_;
  assign new_n1053_ = ~new_n834_ & ~new_n1021_;
  assign new_n1054_ = new_n834_ & new_n1021_;
  assign new_n1055_ = ~new_n1053_ & ~new_n1054_;
  assign new_n1056_ = ~new_n1027_ & ~new_n1055_;
  assign new_n1057_ = new_n1027_ & new_n1055_;
  assign new_n1058_ = ~new_n1056_ & ~new_n1057_;
  assign new_n1059_ = ~new_n718_ & ~new_n1058_;
  assign new_n1060_ = ~new_n718_ & new_n1059_;
  assign new_n1061_ = ~new_n1052_ & ~new_n1060_;
  assign new_n1062_ = ~new_n1041_ & ~new_n1061_;
  assign new_n1063_ = new_n1041_ & new_n1061_;
  assign new_n1064_ = ~new_n1062_ & ~new_n1063_;
  assign new_n1065_ = ~new_n677_ & ~new_n1064_;
  assign new_n1066_ = ~new_n677_ & new_n1065_;
  assign new_n1067_ = ~new_n1050_ & ~new_n1066_;
  assign new_n1068_ = ~\V1213(0)  & ~new_n1067_;
  assign new_n1069_ = \V1213(0)  & new_n1067_;
  assign new_n1070_ = ~new_n1068_ & ~new_n1069_;
  assign new_n1071_ = new_n677_ & ~new_n727_;
  assign new_n1072_ = new_n677_ & new_n1071_;
  assign new_n1073_ = ~new_n1008_ & ~new_n1038_;
  assign new_n1074_ = ~new_n1039_ & ~new_n1073_;
  assign new_n1075_ = ~new_n677_ & ~new_n1074_;
  assign new_n1076_ = ~new_n677_ & new_n1075_;
  assign new_n1077_ = ~new_n1072_ & ~new_n1076_;
  assign new_n1078_ = ~\V1213(2)  & ~new_n1077_;
  assign new_n1079_ = \V1213(2)  & new_n1077_;
  assign new_n1080_ = ~new_n1078_ & ~new_n1079_;
  assign new_n1081_ = ~\V288(4)  & ~\V288(5) ;
  assign new_n1082_ = ~new_n673_ & new_n1014_;
  assign new_n1083_ = new_n1048_ & new_n1082_;
  assign new_n1084_ = new_n1070_ & new_n1083_;
  assign new_n1085_ = new_n1080_ & new_n1084_;
  assign new_n1086_ = ~new_n1081_ & new_n1085_;
  assign new_n1087_ = ~new_n673_ & ~\V1213(3) ;
  assign new_n1088_ = ~\V1213(1)  & new_n1087_;
  assign new_n1089_ = ~\V1213(0)  & new_n1088_;
  assign new_n1090_ = ~\V1213(2)  & new_n1089_;
  assign new_n1091_ = ~new_n754_ & new_n1090_;
  assign new_n1092_ = ~new_n673_ & \V1213(2) ;
  assign new_n1093_ = ~\V1213(1)  & new_n1092_;
  assign new_n1094_ = ~\V1213(0)  & new_n1093_;
  assign new_n1095_ = ~\V1213(3)  & new_n1094_;
  assign new_n1096_ = \V288(6)  & new_n1095_;
  assign new_n1097_ = \V288(7)  & new_n1096_;
  assign new_n1098_ = new_n681_ & ~\V1213(3) ;
  assign new_n1099_ = ~new_n681_ & \V1213(3) ;
  assign new_n1100_ = ~new_n1098_ & ~new_n1099_;
  assign new_n1101_ = ~\V1213(1)  & ~new_n1022_;
  assign new_n1102_ = \V1213(1)  & new_n1022_;
  assign new_n1103_ = ~new_n1101_ & ~new_n1102_;
  assign new_n1104_ = ~\V1213(0)  & ~new_n1055_;
  assign new_n1105_ = \V1213(0)  & new_n1055_;
  assign new_n1106_ = ~new_n1104_ & ~new_n1105_;
  assign new_n1107_ = ~\V1213(2)  & ~new_n1024_;
  assign new_n1108_ = \V1213(2)  & new_n1024_;
  assign new_n1109_ = ~new_n1107_ & ~new_n1108_;
  assign new_n1110_ = ~new_n673_ & new_n1100_;
  assign new_n1111_ = new_n1103_ & new_n1110_;
  assign new_n1112_ = new_n1106_ & new_n1111_;
  assign new_n1113_ = new_n1109_ & new_n1112_;
  assign new_n1114_ = new_n753_ & new_n1113_;
  assign new_n1115_ = new_n684_ & ~\V1213(3) ;
  assign new_n1116_ = ~new_n684_ & \V1213(3) ;
  assign new_n1117_ = ~new_n1115_ & ~new_n1116_;
  assign new_n1118_ = ~\V1213(1)  & ~new_n937_;
  assign new_n1119_ = \V1213(1)  & new_n937_;
  assign new_n1120_ = ~new_n1118_ & ~new_n1119_;
  assign new_n1121_ = ~\V1213(0)  & ~new_n970_;
  assign new_n1122_ = \V1213(0)  & new_n970_;
  assign new_n1123_ = ~new_n1121_ & ~new_n1122_;
  assign new_n1124_ = ~\V1213(2)  & ~new_n939_;
  assign new_n1125_ = \V1213(2)  & new_n939_;
  assign new_n1126_ = ~new_n1124_ & ~new_n1125_;
  assign new_n1127_ = ~new_n673_ & new_n1117_;
  assign new_n1128_ = new_n1120_ & new_n1127_;
  assign new_n1129_ = new_n1123_ & new_n1128_;
  assign new_n1130_ = new_n1126_ & new_n1129_;
  assign new_n1131_ = new_n747_ & new_n1130_;
  assign new_n1132_ = new_n687_ & ~\V1213(3) ;
  assign new_n1133_ = ~new_n687_ & \V1213(3) ;
  assign new_n1134_ = ~new_n1132_ & ~new_n1133_;
  assign new_n1135_ = ~new_n786_ & ~\V1213(1) ;
  assign new_n1136_ = new_n786_ & \V1213(1) ;
  assign new_n1137_ = ~new_n1135_ & ~new_n1136_;
  assign new_n1138_ = ~new_n857_ & ~\V1213(0) ;
  assign new_n1139_ = new_n857_ & \V1213(0) ;
  assign new_n1140_ = ~new_n1138_ & ~new_n1139_;
  assign new_n1141_ = ~new_n788_ & ~\V1213(2) ;
  assign new_n1142_ = new_n788_ & \V1213(2) ;
  assign new_n1143_ = ~new_n1141_ & ~new_n1142_;
  assign new_n1144_ = ~new_n673_ & new_n1134_;
  assign new_n1145_ = new_n1137_ & new_n1144_;
  assign new_n1146_ = new_n1140_ & new_n1145_;
  assign new_n1147_ = new_n1143_ & new_n1146_;
  assign new_n1148_ = new_n741_ & new_n1147_;
  assign new_n1149_ = new_n674_ & ~new_n916_;
  assign new_n1150_ = ~new_n1001_ & new_n1149_;
  assign new_n1151_ = ~new_n1086_ & new_n1150_;
  assign new_n1152_ = ~new_n1091_ & new_n1151_;
  assign new_n1153_ = ~new_n1097_ & new_n1152_;
  assign new_n1154_ = ~new_n1114_ & new_n1153_;
  assign new_n1155_ = ~new_n1131_ & new_n1154_;
  assign V356 = ~new_n1148_ & new_n1155_;
  assign new_n1157_ = ~new_n695_ & ~\V1213(3) ;
  assign new_n1158_ = new_n695_ & \V1213(3) ;
  assign new_n1159_ = ~new_n1157_ & ~new_n1158_;
  assign new_n1160_ = ~new_n795_ & ~\V1213(1) ;
  assign new_n1161_ = new_n795_ & \V1213(1) ;
  assign new_n1162_ = ~new_n1160_ & ~new_n1161_;
  assign new_n1163_ = ~new_n863_ & ~\V1213(0) ;
  assign new_n1164_ = new_n863_ & \V1213(0) ;
  assign new_n1165_ = ~new_n1163_ & ~new_n1164_;
  assign new_n1166_ = ~new_n802_ & ~\V1213(2) ;
  assign new_n1167_ = new_n802_ & \V1213(2) ;
  assign new_n1168_ = ~new_n1166_ & ~new_n1167_;
  assign new_n1169_ = ~new_n673_ & new_n1159_;
  assign new_n1170_ = new_n1162_ & new_n1169_;
  assign new_n1171_ = new_n1165_ & new_n1170_;
  assign new_n1172_ = new_n1168_ & new_n1171_;
  assign new_n1173_ = \V288(0)  & new_n1172_;
  assign new_n1174_ = ~\V1213(3)  & ~new_n923_;
  assign new_n1175_ = \V1213(3)  & new_n923_;
  assign new_n1176_ = ~new_n1174_ & ~new_n1175_;
  assign new_n1177_ = ~\V1213(1)  & ~new_n946_;
  assign new_n1178_ = \V1213(1)  & new_n946_;
  assign new_n1179_ = ~new_n1177_ & ~new_n1178_;
  assign new_n1180_ = ~\V1213(0)  & ~new_n976_;
  assign new_n1181_ = \V1213(0)  & new_n976_;
  assign new_n1182_ = ~new_n1180_ & ~new_n1181_;
  assign new_n1183_ = ~\V1213(2)  & ~new_n953_;
  assign new_n1184_ = \V1213(2)  & new_n953_;
  assign new_n1185_ = ~new_n1183_ & ~new_n1184_;
  assign new_n1186_ = ~new_n673_ & new_n1176_;
  assign new_n1187_ = new_n1179_ & new_n1186_;
  assign new_n1188_ = new_n1182_ & new_n1187_;
  assign new_n1189_ = new_n1185_ & new_n1188_;
  assign new_n1190_ = \V288(2)  & new_n1189_;
  assign new_n1191_ = ~\V1213(3)  & ~new_n1008_;
  assign new_n1192_ = \V1213(3)  & new_n1008_;
  assign new_n1193_ = ~new_n1191_ & ~new_n1192_;
  assign new_n1194_ = ~\V1213(1)  & ~new_n1031_;
  assign new_n1195_ = \V1213(1)  & new_n1031_;
  assign new_n1196_ = ~new_n1194_ & ~new_n1195_;
  assign new_n1197_ = ~\V1213(0)  & ~new_n1061_;
  assign new_n1198_ = \V1213(0)  & new_n1061_;
  assign new_n1199_ = ~new_n1197_ & ~new_n1198_;
  assign new_n1200_ = ~\V1213(2)  & ~new_n1038_;
  assign new_n1201_ = \V1213(2)  & new_n1038_;
  assign new_n1202_ = ~new_n1200_ & ~new_n1201_;
  assign new_n1203_ = ~new_n673_ & new_n1193_;
  assign new_n1204_ = new_n1196_ & new_n1203_;
  assign new_n1205_ = new_n1199_ & new_n1204_;
  assign new_n1206_ = new_n1202_ & new_n1205_;
  assign new_n1207_ = \V288(4)  & new_n1206_;
  assign new_n1208_ = ~new_n673_ & \V1213(3) ;
  assign new_n1209_ = ~\V1213(1)  & new_n1208_;
  assign new_n1210_ = ~\V1213(0)  & new_n1209_;
  assign new_n1211_ = ~\V1213(2)  & new_n1210_;
  assign new_n1212_ = \V288(6)  & new_n1211_;
  assign new_n1213_ = ~new_n673_ & ~\V1213(1) ;
  assign new_n1214_ = ~\V1213(0)  & new_n1213_;
  assign new_n1215_ = \V1213(2)  & new_n1214_;
  assign new_n1216_ = \V1213(3)  & new_n1215_;
  assign new_n1217_ = \V288(6)  & new_n1216_;
  assign new_n1218_ = \V288(7)  & new_n1217_;
  assign new_n1219_ = ~new_n681_ & ~\V1213(3) ;
  assign new_n1220_ = new_n681_ & \V1213(3) ;
  assign new_n1221_ = ~new_n1219_ & ~new_n1220_;
  assign new_n1222_ = ~new_n760_ & ~\V1213(1) ;
  assign new_n1223_ = new_n760_ & \V1213(1) ;
  assign new_n1224_ = ~new_n1222_ & ~new_n1223_;
  assign new_n1225_ = ~new_n834_ & ~\V1213(0) ;
  assign new_n1226_ = new_n834_ & \V1213(0) ;
  assign new_n1227_ = ~new_n1225_ & ~new_n1226_;
  assign new_n1228_ = ~new_n727_ & ~\V1213(2) ;
  assign new_n1229_ = new_n727_ & \V1213(2) ;
  assign new_n1230_ = ~new_n1228_ & ~new_n1229_;
  assign new_n1231_ = ~new_n673_ & new_n1221_;
  assign new_n1232_ = new_n1224_ & new_n1231_;
  assign new_n1233_ = new_n1227_ & new_n1232_;
  assign new_n1234_ = new_n1230_ & new_n1233_;
  assign new_n1235_ = new_n753_ & new_n1234_;
  assign new_n1236_ = ~new_n684_ & ~\V1213(3) ;
  assign new_n1237_ = new_n684_ & \V1213(3) ;
  assign new_n1238_ = ~new_n1236_ & ~new_n1237_;
  assign new_n1239_ = ~new_n766_ & ~\V1213(1) ;
  assign new_n1240_ = new_n766_ & \V1213(1) ;
  assign new_n1241_ = ~new_n1239_ & ~new_n1240_;
  assign new_n1242_ = ~new_n842_ & ~\V1213(0) ;
  assign new_n1243_ = new_n842_ & \V1213(0) ;
  assign new_n1244_ = ~new_n1242_ & ~new_n1243_;
  assign new_n1245_ = ~new_n734_ & ~\V1213(2) ;
  assign new_n1246_ = new_n734_ & \V1213(2) ;
  assign new_n1247_ = ~new_n1245_ & ~new_n1246_;
  assign new_n1248_ = ~new_n673_ & new_n1238_;
  assign new_n1249_ = new_n1241_ & new_n1248_;
  assign new_n1250_ = new_n1244_ & new_n1249_;
  assign new_n1251_ = new_n1247_ & new_n1250_;
  assign new_n1252_ = new_n747_ & new_n1251_;
  assign new_n1253_ = ~new_n687_ & ~\V1213(3) ;
  assign new_n1254_ = new_n687_ & \V1213(3) ;
  assign new_n1255_ = ~new_n1253_ & ~new_n1254_;
  assign new_n1256_ = ~new_n772_ & ~\V1213(1) ;
  assign new_n1257_ = new_n772_ & \V1213(1) ;
  assign new_n1258_ = ~new_n1256_ & ~new_n1257_;
  assign new_n1259_ = ~new_n850_ & ~\V1213(0) ;
  assign new_n1260_ = new_n850_ & \V1213(0) ;
  assign new_n1261_ = ~new_n1259_ & ~new_n1260_;
  assign new_n1262_ = ~new_n782_ & ~\V1213(2) ;
  assign new_n1263_ = new_n782_ & \V1213(2) ;
  assign new_n1264_ = ~new_n1262_ & ~new_n1263_;
  assign new_n1265_ = ~new_n673_ & new_n1255_;
  assign new_n1266_ = new_n1258_ & new_n1265_;
  assign new_n1267_ = new_n1261_ & new_n1266_;
  assign new_n1268_ = new_n1264_ & new_n1267_;
  assign new_n1269_ = new_n741_ & new_n1268_;
  assign new_n1270_ = new_n534_ & ~new_n1173_;
  assign new_n1271_ = ~new_n1190_ & new_n1270_;
  assign new_n1272_ = ~new_n1207_ & new_n1271_;
  assign new_n1273_ = ~new_n1212_ & new_n1272_;
  assign new_n1274_ = ~new_n1218_ & new_n1273_;
  assign new_n1275_ = ~new_n1235_ & new_n1274_;
  assign new_n1276_ = ~new_n1252_ & new_n1275_;
  assign V357 = ~new_n1269_ & new_n1276_;
  assign V373 = \V10(0)  & \V13(0) ;
  assign new_n1279_ = \V202(0)  & \V71(0) ;
  assign new_n1280_ = ~\V13(0)  & new_n1279_;
  assign new_n1281_ = \V9(0)  & ~new_n1280_;
  assign V789 = \V4(0)  & new_n1281_;
  assign V1263 = \V9(0)  & \V4(0) ;
  assign V1259 = \V9(0)  & \V3(0) ;
  assign V1387 = \V9(0)  & \V8(0) ;
  assign V780 = \V9(0)  & \V6(0) ;
  assign V778 = \V9(0)  & \V5(0) ;
  assign V787 = \V7(0)  & \V9(0) ;
  assign new_n1289_ = ~\V13(0)  & \V109(0) ;
  assign V1423 = \V1(0)  & \V9(0) ;
  assign V1431 = ~new_n1289_ & V1423;
  assign V1258 = \V9(0)  & \V2(0) ;
  assign new_n1293_ = ~V787 & ~V1431;
  assign new_n1294_ = ~V1258 & new_n1293_;
  assign new_n1295_ = ~V1423 & new_n1294_;
  assign new_n1296_ = ~V1387 & ~V780;
  assign new_n1297_ = ~V778 & new_n1296_;
  assign new_n1298_ = ~V789 & ~V1263;
  assign new_n1299_ = ~V1259 & new_n1298_;
  assign new_n1300_ = new_n1297_ & new_n1299_;
  assign \V375(0)  = ~new_n1295_ | ~new_n1300_;
  assign new_n1302_ = \V203(0)  & \V165(1) ;
  assign new_n1303_ = ~\V165(0)  & new_n1302_;
  assign new_n1304_ = \V165(2)  & new_n1303_;
  assign new_n1305_ = ~\V35(0)  & ~new_n1304_;
  assign V377 = \V203(0)  & ~new_n1305_;
  assign new_n1307_ = \V243(0)  & \V244(0) ;
  assign new_n1308_ = \V245(0)  & new_n1307_;
  assign new_n1309_ = \V246(0)  & new_n1308_;
  assign new_n1310_ = \V165(0)  & ~\V165(2) ;
  assign new_n1311_ = \V165(1)  & new_n1310_;
  assign new_n1312_ = \V240(0)  & ~new_n1311_;
  assign V1719 = ~\V172(0)  & new_n1312_;
  assign new_n1314_ = ~\V248(0)  & new_n1309_;
  assign new_n1315_ = V1719 & new_n1314_;
  assign new_n1316_ = \V247(0)  & new_n1315_;
  assign new_n1317_ = new_n534_ & ~new_n1091_;
  assign new_n1318_ = ~new_n1212_ & new_n1317_;
  assign new_n1319_ = new_n534_ & ~new_n1097_;
  assign new_n1320_ = ~new_n1218_ & new_n1319_;
  assign new_n1321_ = new_n1318_ & new_n1320_;
  assign new_n1322_ = \V288(6)  & ~new_n1321_;
  assign new_n1323_ = \V288(7)  & new_n1322_;
  assign new_n1324_ = new_n534_ & ~new_n1001_;
  assign new_n1325_ = ~new_n1190_ & new_n1324_;
  assign new_n1326_ = new_n534_ & ~new_n1131_;
  assign new_n1327_ = ~new_n1252_ & new_n1326_;
  assign new_n1328_ = new_n1325_ & new_n1327_;
  assign new_n1329_ = new_n747_ & ~new_n1328_;
  assign new_n1330_ = new_n534_ & ~new_n916_;
  assign new_n1331_ = ~new_n1173_ & new_n1330_;
  assign new_n1332_ = new_n534_ & ~new_n1148_;
  assign new_n1333_ = ~new_n1269_ & new_n1332_;
  assign new_n1334_ = new_n1331_ & new_n1333_;
  assign new_n1335_ = new_n741_ & ~new_n1334_;
  assign new_n1336_ = new_n534_ & ~new_n1086_;
  assign new_n1337_ = ~new_n1207_ & new_n1336_;
  assign new_n1338_ = new_n534_ & ~new_n1114_;
  assign new_n1339_ = ~new_n1235_ & new_n1338_;
  assign new_n1340_ = new_n1337_ & new_n1339_;
  assign new_n1341_ = new_n753_ & ~new_n1340_;
  assign new_n1342_ = ~new_n1335_ & ~new_n1341_;
  assign new_n1343_ = ~new_n1323_ & ~new_n1329_;
  assign new_n1344_ = new_n1342_ & new_n1343_;
  assign new_n1345_ = \V239(3)  & ~new_n545_;
  assign new_n1346_ = new_n567_ & new_n1345_;
  assign new_n1347_ = \V199(3)  & new_n545_;
  assign new_n1348_ = ~new_n567_ & new_n1347_;
  assign new_n1349_ = ~new_n1346_ & ~new_n1348_;
  assign new_n1350_ = ~new_n557_ & ~new_n1349_;
  assign new_n1351_ = new_n534_ & new_n1350_;
  assign new_n1352_ = ~new_n542_ & new_n1351_;
  assign new_n1353_ = ~new_n578_ & new_n1352_;
  assign new_n1354_ = ~new_n578_ & new_n1353_;
  assign new_n1355_ = \V32(10)  & new_n583_;
  assign new_n1356_ = new_n578_ & new_n1355_;
  assign new_n1357_ = new_n578_ & new_n1356_;
  assign new_n1358_ = ~new_n1354_ & ~new_n1357_;
  assign new_n1359_ = ~new_n662_ & ~new_n1358_;
  assign new_n1360_ = new_n661_ & new_n1359_;
  assign new_n1361_ = \V88(0)  & new_n662_;
  assign new_n1362_ = ~new_n661_ & new_n1361_;
  assign \V1243(8)  = new_n1360_ | new_n1362_;
  assign new_n1364_ = \V239(2)  & ~new_n545_;
  assign new_n1365_ = new_n567_ & new_n1364_;
  assign new_n1366_ = \V199(2)  & new_n545_;
  assign new_n1367_ = ~new_n567_ & new_n1366_;
  assign new_n1368_ = ~new_n1365_ & ~new_n1367_;
  assign new_n1369_ = ~new_n557_ & ~new_n1368_;
  assign new_n1370_ = new_n534_ & new_n1369_;
  assign new_n1371_ = ~new_n542_ & new_n1370_;
  assign new_n1372_ = ~new_n578_ & new_n1371_;
  assign new_n1373_ = ~new_n578_ & new_n1372_;
  assign new_n1374_ = \V32(9)  & new_n583_;
  assign new_n1375_ = new_n578_ & new_n1374_;
  assign new_n1376_ = new_n578_ & new_n1375_;
  assign new_n1377_ = ~new_n1373_ & ~new_n1376_;
  assign new_n1378_ = ~new_n662_ & ~new_n1377_;
  assign new_n1379_ = new_n661_ & new_n1378_;
  assign new_n1380_ = \V84(5)  & new_n662_;
  assign new_n1381_ = ~new_n661_ & new_n1380_;
  assign \V1243(7)  = new_n1379_ | new_n1381_;
  assign new_n1383_ = \V239(4)  & ~new_n545_;
  assign new_n1384_ = new_n567_ & new_n1383_;
  assign new_n1385_ = \V199(4)  & new_n545_;
  assign new_n1386_ = ~new_n567_ & new_n1385_;
  assign new_n1387_ = ~new_n1384_ & ~new_n1386_;
  assign new_n1388_ = ~new_n557_ & ~new_n1387_;
  assign new_n1389_ = new_n534_ & new_n1388_;
  assign new_n1390_ = ~new_n542_ & new_n1389_;
  assign new_n1391_ = ~new_n578_ & new_n1390_;
  assign new_n1392_ = ~new_n578_ & new_n1391_;
  assign new_n1393_ = \V32(11)  & new_n583_;
  assign new_n1394_ = new_n578_ & new_n1393_;
  assign new_n1395_ = new_n578_ & new_n1394_;
  assign new_n1396_ = ~new_n1392_ & ~new_n1395_;
  assign new_n1397_ = ~new_n662_ & ~new_n1396_;
  assign new_n1398_ = new_n661_ & new_n1397_;
  assign new_n1399_ = \V88(1)  & new_n662_;
  assign new_n1400_ = ~new_n661_ & new_n1399_;
  assign \V1243(9)  = new_n1398_ | new_n1400_;
  assign new_n1402_ = ~\V248(0)  & ~new_n1344_;
  assign new_n1403_ = \V1243(8)  & new_n1402_;
  assign new_n1404_ = \V1243(7)  & new_n1403_;
  assign new_n1405_ = \V1243(9)  & new_n1404_;
  assign new_n1406_ = V1719 & new_n1405_;
  assign new_n1407_ = \V199(4)  & \V199(2) ;
  assign new_n1408_ = \V199(0)  & new_n1407_;
  assign new_n1409_ = \V194(3)  & new_n1408_;
  assign new_n1410_ = \V194(1)  & new_n1409_;
  assign new_n1411_ = \V194(2)  & new_n1410_;
  assign new_n1412_ = \V194(4)  & new_n1411_;
  assign new_n1413_ = \V199(1)  & new_n1412_;
  assign new_n1414_ = \V199(3)  & new_n1413_;
  assign new_n1415_ = ~\V248(0)  & new_n1414_;
  assign new_n1416_ = V1719 & new_n1415_;
  assign new_n1417_ = ~new_n1316_ & ~new_n1406_;
  assign \V393(0)  = new_n1416_ | ~new_n1417_;
  assign new_n1419_ = ~V763 & ~new_n627_;
  assign new_n1420_ = \V802(0)  & ~new_n1419_;
  assign new_n1421_ = ~new_n540_ & ~new_n567_;
  assign new_n1422_ = \V802(0)  & new_n1421_;
  assign new_n1423_ = \V66(0)  & ~new_n1311_;
  assign new_n1424_ = V763 & new_n1423_;
  assign new_n1425_ = ~\V215(0)  & new_n1424_;
  assign new_n1426_ = \V149(4)  & new_n644_;
  assign new_n1427_ = \V88(3)  & new_n603_;
  assign new_n1428_ = ~\V88(3)  & new_n616_;
  assign new_n1429_ = ~new_n1427_ & ~new_n1428_;
  assign new_n1430_ = ~new_n627_ & ~new_n1429_;
  assign new_n1431_ = ~new_n1426_ & ~new_n1430_;
  assign new_n1432_ = ~\V174(0)  & ~new_n631_;
  assign new_n1433_ = ~new_n628_ & new_n1431_;
  assign new_n1434_ = new_n1432_ & new_n1433_;
  assign new_n1435_ = \V56(0)  & ~new_n1434_;
  assign new_n1436_ = new_n534_ & new_n647_;
  assign new_n1437_ = ~new_n630_ & new_n1436_;
  assign new_n1438_ = new_n648_ & new_n1437_;
  assign new_n1439_ = \V802(0)  & ~new_n1438_;
  assign new_n1440_ = new_n627_ & ~new_n1429_;
  assign new_n1441_ = ~new_n626_ & ~new_n627_;
  assign new_n1442_ = new_n647_ & ~new_n1440_;
  assign new_n1443_ = ~new_n1441_ & new_n1442_;
  assign new_n1444_ = new_n534_ & new_n1443_;
  assign new_n1445_ = \V59(0)  & ~new_n1444_;
  assign new_n1446_ = \V62(0)  & new_n628_;
  assign new_n1447_ = \V70(0)  & ~new_n534_;
  assign new_n1448_ = ~new_n1425_ & ~new_n1435_;
  assign new_n1449_ = ~V1719 & ~new_n1422_;
  assign new_n1450_ = new_n1448_ & new_n1449_;
  assign new_n1451_ = ~new_n1446_ & ~new_n1447_;
  assign new_n1452_ = ~new_n1439_ & ~new_n1445_;
  assign new_n1453_ = new_n1451_ & new_n1452_;
  assign \V423(0)  = ~new_n1450_ | ~new_n1453_;
  assign new_n1455_ = \V248(0)  & V1719;
  assign new_n1456_ = ~\V423(0)  & ~new_n1455_;
  assign new_n1457_ = ~\V165(7)  & new_n1311_;
  assign new_n1458_ = V1719 & new_n1457_;
  assign new_n1459_ = \V302(0)  & V1719;
  assign new_n1460_ = new_n1304_ & V1719;
  assign new_n1461_ = ~\V214(0)  & ~new_n1420_;
  assign new_n1462_ = ~new_n1456_ & new_n1461_;
  assign new_n1463_ = ~\V43(0)  & new_n1462_;
  assign new_n1464_ = ~new_n1458_ & new_n1463_;
  assign new_n1465_ = ~new_n1459_ & new_n1464_;
  assign new_n1466_ = ~new_n1416_ & new_n1465_;
  assign new_n1467_ = ~new_n1406_ & new_n1466_;
  assign new_n1468_ = ~new_n1460_ & new_n1467_;
  assign \V398(0)  = new_n1316_ | ~new_n1468_;
  assign new_n1470_ = \V56(0)  & ~new_n1431_;
  assign new_n1471_ = \V59(0)  & ~new_n1443_;
  assign new_n1472_ = ~new_n1446_ & ~new_n1470_;
  assign new_n1473_ = ~new_n1471_ & new_n1472_;
  assign new_n1474_ = ~\V16(0)  & \V15(0) ;
  assign new_n1475_ = \V16(0)  & \V15(0) ;
  assign \V1757(0)  = new_n1474_ | new_n1475_;
  assign new_n1477_ = ~new_n1311_ & ~new_n1473_;
  assign \V410(0)  = \V1757(0)  | ~new_n1477_;
  assign new_n1479_ = \V215(0)  & \V66(0) ;
  assign new_n1480_ = ~\V32(2)  & ~new_n782_;
  assign new_n1481_ = \V32(2)  & new_n782_;
  assign new_n1482_ = ~new_n1480_ & ~new_n1481_;
  assign new_n1483_ = ~\V32(0)  & ~new_n850_;
  assign new_n1484_ = \V32(0)  & new_n850_;
  assign new_n1485_ = ~new_n1483_ & ~new_n1484_;
  assign new_n1486_ = ~\V32(1)  & ~new_n772_;
  assign new_n1487_ = \V32(1)  & new_n772_;
  assign new_n1488_ = ~new_n1486_ & ~new_n1487_;
  assign new_n1489_ = new_n1482_ & new_n1485_;
  assign new_n1490_ = \V32(3)  & new_n1489_;
  assign new_n1491_ = new_n687_ & new_n1490_;
  assign new_n1492_ = new_n1488_ & new_n1491_;
  assign new_n1493_ = \V32(1)  & new_n1485_;
  assign new_n1494_ = new_n772_ & new_n1493_;
  assign new_n1495_ = new_n782_ & new_n1488_;
  assign new_n1496_ = \V32(2)  & new_n1495_;
  assign new_n1497_ = new_n1485_ & new_n1496_;
  assign new_n1498_ = ~new_n1484_ & ~new_n1497_;
  assign new_n1499_ = ~new_n1492_ & ~new_n1494_;
  assign new_n1500_ = new_n1498_ & new_n1499_;
  assign new_n1501_ = \V66(0)  & V763;
  assign new_n1502_ = ~\V149(4)  & new_n596_;
  assign new_n1503_ = \V149(6)  & new_n1502_;
  assign new_n1504_ = \V66(0)  & new_n1503_;
  assign new_n1505_ = ~new_n538_ & ~new_n599_;
  assign new_n1506_ = \V802(0)  & ~new_n1505_;
  assign new_n1507_ = ~V763 & new_n1506_;
  assign new_n1508_ = \V802(0)  & new_n544_;
  assign new_n1509_ = ~\V174(0)  & new_n494_;
  assign new_n1510_ = ~\V149(4)  & new_n497_;
  assign new_n1511_ = \V149(6)  & new_n1510_;
  assign new_n1512_ = ~\V149(4)  & new_n492_;
  assign new_n1513_ = \V149(6)  & new_n1512_;
  assign new_n1514_ = ~\V149(6)  & new_n1512_;
  assign new_n1515_ = ~new_n1513_ & ~new_n1514_;
  assign new_n1516_ = ~new_n1509_ & ~new_n1511_;
  assign new_n1517_ = new_n1515_ & new_n1516_;
  assign new_n1518_ = \V56(0)  & ~new_n1517_;
  assign new_n1519_ = ~new_n1508_ & ~new_n1518_;
  assign new_n1520_ = ~new_n1501_ & ~new_n1504_;
  assign new_n1521_ = ~new_n1507_ & new_n1520_;
  assign new_n1522_ = new_n1519_ & new_n1521_;
  assign new_n1523_ = ~new_n1500_ & ~new_n1522_;
  assign new_n1524_ = ~\V88(2)  & \V88(3) ;
  assign new_n1525_ = \V88(2)  & ~\V88(3) ;
  assign new_n1526_ = ~new_n1524_ & ~new_n1525_;
  assign new_n1527_ = \V88(1)  & ~\V88(0) ;
  assign new_n1528_ = ~\V88(1)  & \V88(0) ;
  assign new_n1529_ = ~new_n1527_ & ~new_n1528_;
  assign new_n1530_ = ~new_n1526_ & new_n1529_;
  assign new_n1531_ = new_n1526_ & ~new_n1529_;
  assign new_n1532_ = ~new_n1530_ & ~new_n1531_;
  assign new_n1533_ = \V84(5)  & ~\V84(4) ;
  assign new_n1534_ = ~\V84(5)  & \V84(4) ;
  assign new_n1535_ = ~new_n1533_ & ~new_n1534_;
  assign new_n1536_ = \V84(3)  & ~\V84(2) ;
  assign new_n1537_ = ~\V84(3)  & \V84(2) ;
  assign new_n1538_ = ~new_n1536_ & ~new_n1537_;
  assign new_n1539_ = ~new_n1535_ & new_n1538_;
  assign new_n1540_ = new_n1535_ & ~new_n1538_;
  assign new_n1541_ = ~new_n1539_ & ~new_n1540_;
  assign new_n1542_ = ~new_n1532_ & new_n1541_;
  assign new_n1543_ = new_n1532_ & ~new_n1541_;
  assign new_n1544_ = ~new_n1542_ & ~new_n1543_;
  assign new_n1545_ = \V94(1)  & new_n1544_;
  assign new_n1546_ = ~\V94(1)  & ~new_n1544_;
  assign new_n1547_ = ~new_n1545_ & ~new_n1546_;
  assign new_n1548_ = \V84(1)  & ~\V84(0) ;
  assign new_n1549_ = ~\V84(1)  & \V84(0) ;
  assign new_n1550_ = ~new_n1548_ & ~new_n1549_;
  assign new_n1551_ = \V78(5)  & ~\V78(4) ;
  assign new_n1552_ = ~\V78(5)  & \V78(4) ;
  assign new_n1553_ = ~new_n1551_ & ~new_n1552_;
  assign new_n1554_ = ~new_n1550_ & new_n1553_;
  assign new_n1555_ = new_n1550_ & ~new_n1553_;
  assign new_n1556_ = ~new_n1554_ & ~new_n1555_;
  assign new_n1557_ = ~\V78(2)  & \V78(3) ;
  assign new_n1558_ = \V78(2)  & ~\V78(3) ;
  assign new_n1559_ = ~new_n1557_ & ~new_n1558_;
  assign new_n1560_ = \V78(1)  & ~\V78(0) ;
  assign new_n1561_ = ~\V78(1)  & \V78(0) ;
  assign new_n1562_ = ~new_n1560_ & ~new_n1561_;
  assign new_n1563_ = ~new_n1559_ & new_n1562_;
  assign new_n1564_ = new_n1559_ & ~new_n1562_;
  assign new_n1565_ = ~new_n1563_ & ~new_n1564_;
  assign new_n1566_ = ~new_n1556_ & new_n1565_;
  assign new_n1567_ = new_n1556_ & ~new_n1565_;
  assign new_n1568_ = ~new_n1566_ & ~new_n1567_;
  assign new_n1569_ = \V94(0)  & new_n1568_;
  assign new_n1570_ = ~\V94(0)  & ~new_n1568_;
  assign new_n1571_ = ~new_n1569_ & ~new_n1570_;
  assign new_n1572_ = ~new_n1547_ & ~new_n1571_;
  assign new_n1573_ = ~\V149(3)  & new_n668_;
  assign new_n1574_ = new_n489_ & new_n1573_;
  assign new_n1575_ = \V149(4)  & new_n1574_;
  assign new_n1576_ = \V149(6)  & new_n1575_;
  assign new_n1577_ = ~new_n598_ & ~new_n1514_;
  assign new_n1578_ = ~new_n1576_ & new_n1577_;
  assign new_n1579_ = \V56(0)  & ~new_n1578_;
  assign new_n1580_ = ~new_n544_ & ~new_n599_;
  assign new_n1581_ = ~new_n538_ & new_n1580_;
  assign new_n1582_ = \V802(0)  & ~new_n1581_;
  assign new_n1583_ = ~new_n1579_ & ~new_n1582_;
  assign new_n1584_ = ~new_n1572_ & ~new_n1583_;
  assign new_n1585_ = \V56(0)  & \V172(0) ;
  assign new_n1586_ = \V207(0)  & ~new_n1585_;
  assign new_n1587_ = ~\V43(0)  & ~\V214(0) ;
  assign new_n1588_ = new_n534_ & new_n1587_;
  assign new_n1589_ = ~new_n1479_ & new_n1588_;
  assign new_n1590_ = ~new_n1523_ & new_n1589_;
  assign new_n1591_ = ~\V1757(0)  & new_n1590_;
  assign new_n1592_ = ~new_n1420_ & new_n1591_;
  assign new_n1593_ = ~new_n1584_ & new_n1592_;
  assign new_n1594_ = ~new_n1586_ & new_n1593_;
  assign new_n1595_ = \V423(0)  & new_n1594_;
  assign new_n1596_ = ~new_n1458_ & new_n1595_;
  assign new_n1597_ = ~new_n1459_ & new_n1596_;
  assign new_n1598_ = ~new_n1416_ & new_n1597_;
  assign new_n1599_ = ~new_n1406_ & new_n1598_;
  assign new_n1600_ = ~new_n1460_ & new_n1599_;
  assign V432 = ~new_n1316_ & new_n1600_;
  assign new_n1602_ = \V56(0)  & new_n598_;
  assign new_n1603_ = \V241(0)  & ~new_n566_;
  assign new_n1604_ = ~new_n549_ & ~new_n1603_;
  assign new_n1605_ = \V59(0)  & new_n540_;
  assign new_n1606_ = ~new_n1604_ & new_n1605_;
  assign new_n1607_ = ~new_n538_ & ~new_n549_;
  assign new_n1608_ = ~new_n537_ & new_n1607_;
  assign new_n1609_ = new_n540_ & ~new_n1608_;
  assign new_n1610_ = \V802(0)  & new_n1609_;
  assign new_n1611_ = ~\V270(0)  & ~new_n1610_;
  assign new_n1612_ = ~new_n1602_ & ~new_n1606_;
  assign new_n1613_ = new_n1611_ & new_n1612_;
  assign new_n1614_ = \V62(0)  & new_n598_;
  assign new_n1615_ = ~\V302(0)  & ~new_n1613_;
  assign V630 = ~new_n1614_ & new_n1615_;
  assign \V435(0)  = V432 | V630;
  assign \V500(0)  = \V271(0)  | ~\V14(0) ;
  assign new_n1619_ = \V59(0)  & new_n631_;
  assign new_n1620_ = new_n1514_ & ~new_n1584_;
  assign new_n1621_ = ~new_n627_ & new_n630_;
  assign new_n1622_ = ~new_n537_ & ~new_n591_;
  assign new_n1623_ = ~new_n538_ & ~new_n1620_;
  assign new_n1624_ = ~new_n1621_ & new_n1623_;
  assign new_n1625_ = new_n1622_ & new_n1624_;
  assign new_n1626_ = \V56(0)  & ~new_n1625_;
  assign new_n1627_ = \V62(0)  & new_n1513_;
  assign new_n1628_ = ~new_n1511_ & ~new_n1513_;
  assign new_n1629_ = \V56(0)  & ~new_n1628_;
  assign new_n1630_ = ~new_n1627_ & ~new_n1629_;
  assign new_n1631_ = ~new_n1619_ & ~new_n1626_;
  assign \V508(0)  = ~new_n1630_ | ~new_n1631_;
  assign new_n1633_ = ~\V43(0)  & \V45(0) ;
  assign \V511(0)  = \V40(0)  | new_n1633_;
  assign new_n1635_ = \V42(0)  & ~\V44(0) ;
  assign new_n1636_ = ~\V42(0)  & \V44(0) ;
  assign new_n1637_ = ~new_n1635_ & ~new_n1636_;
  assign new_n1638_ = \V39(0)  & ~\V38(0) ;
  assign new_n1639_ = ~\V39(0)  & \V38(0) ;
  assign new_n1640_ = ~new_n1638_ & ~new_n1639_;
  assign V512 = new_n1637_ & new_n1640_;
  assign new_n1642_ = \V59(0)  & ~new_n627_;
  assign new_n1643_ = ~new_n626_ & new_n1642_;
  assign new_n1644_ = \V56(0)  & new_n1426_;
  assign new_n1645_ = \V56(0)  & new_n1430_;
  assign new_n1646_ = \V59(0)  & new_n1440_;
  assign new_n1647_ = \V59(0)  & ~new_n647_;
  assign new_n1648_ = ~new_n1446_ & ~new_n1643_;
  assign new_n1649_ = ~new_n1644_ & new_n1648_;
  assign new_n1650_ = ~new_n1645_ & new_n1649_;
  assign new_n1651_ = ~new_n1646_ & new_n1650_;
  assign new_n1652_ = ~new_n1647_ & new_n1651_;
  assign new_n1653_ = ~\V214(0)  & ~new_n1586_;
  assign new_n1654_ = ~new_n1652_ & new_n1653_;
  assign new_n1655_ = ~new_n1311_ & new_n1654_;
  assign V527 = ~\V43(0)  & new_n1655_;
  assign V537 = new_n538_ & \V1213(0) ;
  assign V538 = new_n538_ & \V1213(1) ;
  assign V539 = new_n538_ & \V1213(2) ;
  assign V540 = new_n538_ & \V1213(3) ;
  assign new_n1661_ = \V257(6)  & ~new_n534_;
  assign new_n1662_ = ~new_n542_ & new_n1661_;
  assign new_n1663_ = new_n557_ & new_n1662_;
  assign new_n1664_ = \V223(4)  & ~new_n545_;
  assign new_n1665_ = new_n567_ & new_n1664_;
  assign new_n1666_ = \V183(4)  & new_n545_;
  assign new_n1667_ = ~new_n567_ & new_n1666_;
  assign new_n1668_ = ~new_n1665_ & ~new_n1667_;
  assign new_n1669_ = new_n534_ & ~new_n1668_;
  assign new_n1670_ = ~new_n542_ & new_n1669_;
  assign new_n1671_ = ~new_n557_ & new_n1670_;
  assign new_n1672_ = ~new_n1663_ & ~new_n1671_;
  assign new_n1673_ = ~new_n578_ & ~new_n1672_;
  assign new_n1674_ = ~new_n578_ & new_n1673_;
  assign new_n1675_ = ~new_n662_ & new_n1674_;
  assign new_n1676_ = new_n661_ & new_n1675_;
  assign new_n1677_ = \V32(4)  & new_n662_;
  assign new_n1678_ = ~new_n661_ & new_n1677_;
  assign \V1213(4)  = new_n1676_ | new_n1678_;
  assign V541 = new_n538_ & \V1213(4) ;
  assign new_n1681_ = \V257(0)  & ~new_n534_;
  assign new_n1682_ = ~new_n542_ & new_n1681_;
  assign new_n1683_ = new_n557_ & new_n1682_;
  assign new_n1684_ = \V223(5)  & ~new_n545_;
  assign new_n1685_ = new_n567_ & new_n1684_;
  assign new_n1686_ = \V183(5)  & new_n545_;
  assign new_n1687_ = ~new_n567_ & new_n1686_;
  assign new_n1688_ = ~new_n1685_ & ~new_n1687_;
  assign new_n1689_ = new_n534_ & ~new_n1688_;
  assign new_n1690_ = ~new_n542_ & new_n1689_;
  assign new_n1691_ = ~new_n557_ & new_n1690_;
  assign new_n1692_ = ~new_n1683_ & ~new_n1691_;
  assign new_n1693_ = ~new_n578_ & ~new_n1692_;
  assign new_n1694_ = ~new_n578_ & new_n1693_;
  assign new_n1695_ = new_n578_ & ~new_n583_;
  assign new_n1696_ = new_n578_ & new_n1695_;
  assign new_n1697_ = ~new_n1694_ & ~new_n1696_;
  assign new_n1698_ = ~new_n662_ & ~new_n1697_;
  assign new_n1699_ = new_n661_ & new_n1698_;
  assign new_n1700_ = \V32(5)  & new_n662_;
  assign new_n1701_ = ~new_n661_ & new_n1700_;
  assign \V1213(5)  = new_n1699_ | new_n1701_;
  assign V542 = new_n538_ & \V1213(5) ;
  assign new_n1704_ = \V257(1)  & ~new_n534_;
  assign new_n1705_ = ~new_n542_ & new_n1704_;
  assign new_n1706_ = new_n557_ & new_n1705_;
  assign new_n1707_ = \V229(0)  & ~new_n545_;
  assign new_n1708_ = new_n567_ & new_n1707_;
  assign new_n1709_ = \V189(0)  & new_n545_;
  assign new_n1710_ = ~new_n567_ & new_n1709_;
  assign new_n1711_ = ~new_n1708_ & ~new_n1710_;
  assign new_n1712_ = new_n534_ & ~new_n1711_;
  assign new_n1713_ = ~new_n542_ & new_n1712_;
  assign new_n1714_ = ~new_n557_ & new_n1713_;
  assign new_n1715_ = ~new_n1706_ & ~new_n1714_;
  assign new_n1716_ = ~new_n578_ & ~new_n1715_;
  assign new_n1717_ = ~new_n578_ & new_n1716_;
  assign new_n1718_ = new_n578_ & new_n583_;
  assign new_n1719_ = new_n578_ & new_n1718_;
  assign new_n1720_ = ~new_n1717_ & ~new_n1719_;
  assign new_n1721_ = ~new_n662_ & ~new_n1720_;
  assign new_n1722_ = new_n661_ & new_n1721_;
  assign new_n1723_ = \V32(6)  & new_n662_;
  assign new_n1724_ = ~new_n661_ & new_n1723_;
  assign \V1213(6)  = new_n1722_ | new_n1724_;
  assign V543 = new_n538_ & \V1213(6) ;
  assign new_n1727_ = \V257(2)  & ~new_n534_;
  assign new_n1728_ = ~new_n542_ & new_n1727_;
  assign new_n1729_ = new_n557_ & new_n1728_;
  assign new_n1730_ = \V229(1)  & ~new_n545_;
  assign new_n1731_ = new_n567_ & new_n1730_;
  assign new_n1732_ = \V189(1)  & new_n545_;
  assign new_n1733_ = ~new_n567_ & new_n1732_;
  assign new_n1734_ = ~new_n1731_ & ~new_n1733_;
  assign new_n1735_ = new_n534_ & ~new_n1734_;
  assign new_n1736_ = ~new_n542_ & new_n1735_;
  assign new_n1737_ = ~new_n557_ & new_n1736_;
  assign new_n1738_ = ~new_n1729_ & ~new_n1737_;
  assign new_n1739_ = ~new_n578_ & ~new_n1738_;
  assign new_n1740_ = ~new_n578_ & new_n1739_;
  assign new_n1741_ = \V32(0)  & ~new_n583_;
  assign new_n1742_ = ~new_n583_ & new_n1741_;
  assign new_n1743_ = ~new_n583_ & ~new_n1742_;
  assign new_n1744_ = new_n578_ & ~new_n1743_;
  assign new_n1745_ = new_n578_ & new_n1744_;
  assign new_n1746_ = ~new_n1740_ & ~new_n1745_;
  assign new_n1747_ = ~new_n662_ & ~new_n1746_;
  assign new_n1748_ = new_n661_ & new_n1747_;
  assign new_n1749_ = \V32(7)  & new_n662_;
  assign new_n1750_ = ~new_n661_ & new_n1749_;
  assign \V1213(7)  = new_n1748_ | new_n1750_;
  assign V544 = new_n538_ & \V1213(7) ;
  assign new_n1753_ = \V257(3)  & ~new_n534_;
  assign new_n1754_ = ~new_n542_ & new_n1753_;
  assign new_n1755_ = new_n557_ & new_n1754_;
  assign new_n1756_ = \V229(2)  & ~new_n545_;
  assign new_n1757_ = new_n567_ & new_n1756_;
  assign new_n1758_ = \V189(2)  & new_n545_;
  assign new_n1759_ = ~new_n567_ & new_n1758_;
  assign new_n1760_ = ~new_n1757_ & ~new_n1759_;
  assign new_n1761_ = new_n534_ & ~new_n1760_;
  assign new_n1762_ = ~new_n542_ & new_n1761_;
  assign new_n1763_ = ~new_n557_ & new_n1762_;
  assign new_n1764_ = ~new_n1755_ & ~new_n1763_;
  assign new_n1765_ = ~new_n578_ & ~new_n1764_;
  assign new_n1766_ = ~new_n578_ & new_n1765_;
  assign new_n1767_ = \V32(1)  & ~new_n583_;
  assign new_n1768_ = ~new_n583_ & new_n1767_;
  assign new_n1769_ = ~new_n583_ & ~new_n1768_;
  assign new_n1770_ = new_n578_ & ~new_n1769_;
  assign new_n1771_ = new_n578_ & new_n1770_;
  assign new_n1772_ = ~new_n1766_ & ~new_n1771_;
  assign new_n1773_ = ~new_n662_ & ~new_n1772_;
  assign new_n1774_ = new_n661_ & new_n1773_;
  assign new_n1775_ = \V32(8)  & new_n662_;
  assign new_n1776_ = ~new_n661_ & new_n1775_;
  assign \V1213(8)  = new_n1774_ | new_n1776_;
  assign V545 = new_n538_ & \V1213(8) ;
  assign new_n1779_ = \V257(4)  & ~new_n534_;
  assign new_n1780_ = ~new_n542_ & new_n1779_;
  assign new_n1781_ = new_n557_ & new_n1780_;
  assign new_n1782_ = \V229(3)  & ~new_n545_;
  assign new_n1783_ = new_n567_ & new_n1782_;
  assign new_n1784_ = \V189(3)  & new_n545_;
  assign new_n1785_ = ~new_n567_ & new_n1784_;
  assign new_n1786_ = ~new_n1783_ & ~new_n1785_;
  assign new_n1787_ = new_n534_ & ~new_n1786_;
  assign new_n1788_ = ~new_n542_ & new_n1787_;
  assign new_n1789_ = ~new_n557_ & new_n1788_;
  assign new_n1790_ = ~new_n1781_ & ~new_n1789_;
  assign new_n1791_ = ~new_n578_ & ~new_n1790_;
  assign new_n1792_ = ~new_n578_ & new_n1791_;
  assign new_n1793_ = \V32(2)  & ~new_n583_;
  assign new_n1794_ = ~new_n583_ & new_n1793_;
  assign new_n1795_ = ~new_n583_ & ~new_n1794_;
  assign new_n1796_ = new_n578_ & ~new_n1795_;
  assign new_n1797_ = new_n578_ & new_n1796_;
  assign new_n1798_ = ~new_n1792_ & ~new_n1797_;
  assign new_n1799_ = ~new_n662_ & ~new_n1798_;
  assign new_n1800_ = new_n661_ & new_n1799_;
  assign new_n1801_ = \V32(9)  & new_n662_;
  assign new_n1802_ = ~new_n661_ & new_n1801_;
  assign \V1213(9)  = new_n1800_ | new_n1802_;
  assign V546 = new_n538_ & \V1213(9) ;
  assign new_n1805_ = \V257(5)  & ~new_n534_;
  assign new_n1806_ = ~new_n542_ & new_n1805_;
  assign new_n1807_ = new_n557_ & new_n1806_;
  assign new_n1808_ = \V229(4)  & ~new_n545_;
  assign new_n1809_ = new_n567_ & new_n1808_;
  assign new_n1810_ = \V189(4)  & new_n545_;
  assign new_n1811_ = ~new_n567_ & new_n1810_;
  assign new_n1812_ = ~new_n1809_ & ~new_n1811_;
  assign new_n1813_ = new_n534_ & ~new_n1812_;
  assign new_n1814_ = ~new_n542_ & new_n1813_;
  assign new_n1815_ = ~new_n557_ & new_n1814_;
  assign new_n1816_ = ~new_n1807_ & ~new_n1815_;
  assign new_n1817_ = ~new_n578_ & ~new_n1816_;
  assign new_n1818_ = ~new_n578_ & new_n1817_;
  assign new_n1819_ = \V32(0)  & new_n583_;
  assign new_n1820_ = \V32(3)  & ~new_n583_;
  assign new_n1821_ = ~new_n583_ & new_n1820_;
  assign new_n1822_ = ~new_n1819_ & ~new_n1821_;
  assign new_n1823_ = new_n578_ & ~new_n1822_;
  assign new_n1824_ = new_n578_ & new_n1823_;
  assign new_n1825_ = ~new_n1818_ & ~new_n1824_;
  assign new_n1826_ = ~new_n662_ & ~new_n1825_;
  assign new_n1827_ = new_n661_ & new_n1826_;
  assign new_n1828_ = \V32(10)  & new_n662_;
  assign new_n1829_ = ~new_n661_ & new_n1828_;
  assign \V1213(10)  = new_n1827_ | new_n1829_;
  assign V547 = new_n538_ & \V1213(10) ;
  assign new_n1832_ = \V229(5)  & ~new_n545_;
  assign new_n1833_ = new_n567_ & new_n1832_;
  assign new_n1834_ = \V189(5)  & new_n545_;
  assign new_n1835_ = ~new_n567_ & new_n1834_;
  assign new_n1836_ = ~new_n1833_ & ~new_n1835_;
  assign new_n1837_ = new_n534_ & ~new_n1836_;
  assign new_n1838_ = ~new_n542_ & new_n1837_;
  assign new_n1839_ = ~new_n557_ & new_n1838_;
  assign new_n1840_ = ~new_n1663_ & ~new_n1839_;
  assign new_n1841_ = ~new_n578_ & ~new_n1840_;
  assign new_n1842_ = ~new_n578_ & new_n1841_;
  assign new_n1843_ = \V32(1)  & new_n583_;
  assign new_n1844_ = \V32(4)  & ~new_n583_;
  assign new_n1845_ = ~new_n583_ & new_n1844_;
  assign new_n1846_ = ~new_n1843_ & ~new_n1845_;
  assign new_n1847_ = new_n578_ & ~new_n1846_;
  assign new_n1848_ = new_n578_ & new_n1847_;
  assign new_n1849_ = ~new_n1842_ & ~new_n1848_;
  assign new_n1850_ = ~new_n662_ & ~new_n1849_;
  assign new_n1851_ = new_n661_ & new_n1850_;
  assign new_n1852_ = \V32(11)  & new_n662_;
  assign new_n1853_ = ~new_n661_ & new_n1852_;
  assign \V1213(11)  = new_n1851_ | new_n1853_;
  assign V548 = new_n538_ & \V1213(11) ;
  assign new_n1856_ = ~\V802(0)  & ~new_n540_;
  assign new_n1857_ = ~new_n567_ & new_n1856_;
  assign new_n1858_ = \V194(0)  & new_n1414_;
  assign new_n1859_ = \V271(0)  & ~new_n598_;
  assign new_n1860_ = ~\V274(0)  & new_n1859_;
  assign new_n1861_ = ~new_n1858_ & new_n1860_;
  assign new_n1862_ = new_n540_ & new_n1861_;
  assign new_n1863_ = \V134(0)  & new_n1862_;
  assign new_n1864_ = \V134(1)  & new_n1863_;
  assign new_n1865_ = ~new_n1857_ & ~new_n1864_;
  assign new_n1866_ = \V802(0)  & new_n537_;
  assign new_n1867_ = \V802(0)  & \V1243(9) ;
  assign new_n1868_ = new_n538_ & new_n1867_;
  assign new_n1869_ = new_n1865_ & new_n1868_;
  assign new_n1870_ = ~new_n1866_ & new_n1869_;
  assign new_n1871_ = \V802(0)  & new_n538_;
  assign new_n1872_ = ~\V199(4)  & ~new_n1866_;
  assign new_n1873_ = ~new_n1865_ & new_n1872_;
  assign new_n1874_ = ~new_n1871_ & new_n1873_;
  assign \V572(9)  = new_n1870_ | new_n1874_;
  assign new_n1876_ = \V802(0)  & \V1243(8) ;
  assign new_n1877_ = new_n538_ & new_n1876_;
  assign new_n1878_ = new_n1865_ & new_n1877_;
  assign new_n1879_ = ~new_n1866_ & new_n1878_;
  assign new_n1880_ = ~\V199(4)  & \V199(3) ;
  assign new_n1881_ = \V199(4)  & ~\V199(3) ;
  assign new_n1882_ = ~new_n1880_ & ~new_n1881_;
  assign new_n1883_ = ~new_n1866_ & ~new_n1882_;
  assign new_n1884_ = ~new_n1865_ & new_n1883_;
  assign new_n1885_ = ~new_n1871_ & new_n1884_;
  assign \V572(8)  = new_n1879_ | new_n1885_;
  assign new_n1887_ = \V802(0)  & \V1243(7) ;
  assign new_n1888_ = new_n538_ & new_n1887_;
  assign new_n1889_ = new_n1865_ & new_n1888_;
  assign new_n1890_ = ~new_n1866_ & new_n1889_;
  assign new_n1891_ = \V199(4)  & \V199(3) ;
  assign new_n1892_ = \V199(2)  & ~new_n1891_;
  assign new_n1893_ = ~\V199(2)  & new_n1891_;
  assign new_n1894_ = ~new_n1892_ & ~new_n1893_;
  assign new_n1895_ = ~new_n1866_ & ~new_n1894_;
  assign new_n1896_ = ~new_n1865_ & new_n1895_;
  assign new_n1897_ = ~new_n1871_ & new_n1896_;
  assign \V572(7)  = new_n1890_ | new_n1897_;
  assign new_n1899_ = \V239(1)  & ~new_n545_;
  assign new_n1900_ = new_n567_ & new_n1899_;
  assign new_n1901_ = \V199(1)  & new_n545_;
  assign new_n1902_ = ~new_n567_ & new_n1901_;
  assign new_n1903_ = ~new_n1900_ & ~new_n1902_;
  assign new_n1904_ = ~new_n557_ & ~new_n1903_;
  assign new_n1905_ = new_n534_ & new_n1904_;
  assign new_n1906_ = ~new_n542_ & new_n1905_;
  assign new_n1907_ = ~new_n578_ & new_n1906_;
  assign new_n1908_ = ~new_n578_ & new_n1907_;
  assign new_n1909_ = \V32(8)  & new_n583_;
  assign new_n1910_ = \V32(11)  & ~new_n583_;
  assign new_n1911_ = ~new_n583_ & new_n1910_;
  assign new_n1912_ = ~new_n1909_ & ~new_n1911_;
  assign new_n1913_ = new_n578_ & ~new_n1912_;
  assign new_n1914_ = new_n578_ & new_n1913_;
  assign new_n1915_ = ~new_n1908_ & ~new_n1914_;
  assign new_n1916_ = ~new_n662_ & ~new_n1915_;
  assign new_n1917_ = new_n661_ & new_n1916_;
  assign new_n1918_ = \V84(4)  & new_n662_;
  assign new_n1919_ = ~new_n661_ & new_n1918_;
  assign \V1243(6)  = new_n1917_ | new_n1919_;
  assign new_n1921_ = \V802(0)  & \V1243(6) ;
  assign new_n1922_ = new_n538_ & new_n1921_;
  assign new_n1923_ = new_n1865_ & new_n1922_;
  assign new_n1924_ = ~new_n1866_ & new_n1923_;
  assign new_n1925_ = \V199(3)  & new_n1407_;
  assign new_n1926_ = \V199(1)  & ~new_n1925_;
  assign new_n1927_ = ~\V199(1)  & new_n1925_;
  assign new_n1928_ = ~new_n1926_ & ~new_n1927_;
  assign new_n1929_ = ~new_n1866_ & ~new_n1928_;
  assign new_n1930_ = ~new_n1865_ & new_n1929_;
  assign new_n1931_ = ~new_n1871_ & new_n1930_;
  assign \V572(6)  = new_n1924_ | new_n1931_;
  assign new_n1933_ = \V239(0)  & ~new_n545_;
  assign new_n1934_ = new_n567_ & new_n1933_;
  assign new_n1935_ = \V199(0)  & new_n545_;
  assign new_n1936_ = ~new_n567_ & new_n1935_;
  assign new_n1937_ = ~new_n1934_ & ~new_n1936_;
  assign new_n1938_ = ~new_n557_ & ~new_n1937_;
  assign new_n1939_ = new_n534_ & new_n1938_;
  assign new_n1940_ = ~new_n542_ & new_n1939_;
  assign new_n1941_ = ~new_n578_ & new_n1940_;
  assign new_n1942_ = ~new_n578_ & new_n1941_;
  assign new_n1943_ = \V32(7)  & new_n583_;
  assign new_n1944_ = \V32(10)  & ~new_n583_;
  assign new_n1945_ = ~new_n583_ & new_n1944_;
  assign new_n1946_ = ~new_n1943_ & ~new_n1945_;
  assign new_n1947_ = new_n578_ & ~new_n1946_;
  assign new_n1948_ = new_n578_ & new_n1947_;
  assign new_n1949_ = ~new_n1942_ & ~new_n1948_;
  assign new_n1950_ = ~new_n662_ & ~new_n1949_;
  assign new_n1951_ = new_n661_ & new_n1950_;
  assign new_n1952_ = \V84(3)  & new_n662_;
  assign new_n1953_ = ~new_n661_ & new_n1952_;
  assign \V1243(5)  = new_n1951_ | new_n1953_;
  assign new_n1955_ = \V802(0)  & \V1243(5) ;
  assign new_n1956_ = new_n538_ & new_n1955_;
  assign new_n1957_ = new_n1865_ & new_n1956_;
  assign new_n1958_ = ~new_n1866_ & new_n1957_;
  assign new_n1959_ = \V199(1)  & new_n1407_;
  assign new_n1960_ = \V199(3)  & new_n1959_;
  assign new_n1961_ = \V199(0)  & ~new_n1960_;
  assign new_n1962_ = ~\V199(0)  & new_n1960_;
  assign new_n1963_ = ~new_n1961_ & ~new_n1962_;
  assign new_n1964_ = ~new_n1866_ & ~new_n1963_;
  assign new_n1965_ = ~new_n1865_ & new_n1964_;
  assign new_n1966_ = ~new_n1871_ & new_n1965_;
  assign \V572(5)  = new_n1958_ | new_n1966_;
  assign new_n1968_ = \V234(4)  & ~new_n545_;
  assign new_n1969_ = new_n567_ & new_n1968_;
  assign new_n1970_ = \V194(4)  & new_n545_;
  assign new_n1971_ = ~new_n567_ & new_n1970_;
  assign new_n1972_ = ~new_n1969_ & ~new_n1971_;
  assign new_n1973_ = ~new_n557_ & ~new_n1972_;
  assign new_n1974_ = new_n534_ & new_n1973_;
  assign new_n1975_ = ~new_n542_ & new_n1974_;
  assign new_n1976_ = ~new_n578_ & new_n1975_;
  assign new_n1977_ = ~new_n578_ & new_n1976_;
  assign new_n1978_ = \V32(6)  & new_n583_;
  assign new_n1979_ = \V32(9)  & ~new_n583_;
  assign new_n1980_ = ~new_n583_ & new_n1979_;
  assign new_n1981_ = ~new_n1978_ & ~new_n1980_;
  assign new_n1982_ = new_n578_ & ~new_n1981_;
  assign new_n1983_ = new_n578_ & new_n1982_;
  assign new_n1984_ = ~new_n1977_ & ~new_n1983_;
  assign new_n1985_ = ~new_n662_ & ~new_n1984_;
  assign new_n1986_ = new_n661_ & new_n1985_;
  assign new_n1987_ = \V84(2)  & new_n662_;
  assign new_n1988_ = ~new_n661_ & new_n1987_;
  assign \V1243(4)  = new_n1986_ | new_n1988_;
  assign new_n1990_ = \V802(0)  & \V1243(4) ;
  assign new_n1991_ = new_n538_ & new_n1990_;
  assign new_n1992_ = new_n1865_ & new_n1991_;
  assign new_n1993_ = ~new_n1866_ & new_n1992_;
  assign new_n1994_ = \V199(1)  & new_n1408_;
  assign new_n1995_ = \V199(3)  & new_n1994_;
  assign new_n1996_ = \V194(4)  & ~new_n1995_;
  assign new_n1997_ = ~\V194(4)  & new_n1995_;
  assign new_n1998_ = ~new_n1996_ & ~new_n1997_;
  assign new_n1999_ = ~new_n1866_ & ~new_n1998_;
  assign new_n2000_ = ~new_n1865_ & new_n1999_;
  assign new_n2001_ = ~new_n1871_ & new_n2000_;
  assign \V572(4)  = new_n1993_ | new_n2001_;
  assign new_n2003_ = \V149(7)  & \V802(0) ;
  assign new_n2004_ = new_n537_ & new_n2003_;
  assign new_n2005_ = new_n1865_ & new_n2004_;
  assign new_n2006_ = ~new_n1871_ & new_n2005_;
  assign new_n2007_ = \V194(4)  & new_n1408_;
  assign new_n2008_ = \V199(1)  & new_n2007_;
  assign new_n2009_ = \V199(3)  & new_n2008_;
  assign new_n2010_ = \V194(3)  & ~new_n2009_;
  assign new_n2011_ = ~\V194(3)  & new_n2009_;
  assign new_n2012_ = ~new_n2010_ & ~new_n2011_;
  assign new_n2013_ = ~new_n1866_ & ~new_n2012_;
  assign new_n2014_ = ~new_n1865_ & new_n2013_;
  assign new_n2015_ = ~new_n1871_ & new_n2014_;
  assign new_n2016_ = \V234(3)  & ~new_n545_;
  assign new_n2017_ = new_n567_ & new_n2016_;
  assign new_n2018_ = \V194(3)  & new_n545_;
  assign new_n2019_ = ~new_n567_ & new_n2018_;
  assign new_n2020_ = ~new_n2017_ & ~new_n2019_;
  assign new_n2021_ = new_n534_ & ~new_n2020_;
  assign new_n2022_ = ~new_n542_ & new_n2021_;
  assign new_n2023_ = ~new_n557_ & new_n2022_;
  assign new_n2024_ = ~\V59(0)  & \V149(7) ;
  assign new_n2025_ = ~new_n540_ & new_n2024_;
  assign new_n2026_ = new_n537_ & new_n2025_;
  assign new_n2027_ = new_n534_ & new_n2026_;
  assign new_n2028_ = new_n557_ & new_n2027_;
  assign new_n2029_ = ~new_n2023_ & ~new_n2028_;
  assign new_n2030_ = ~new_n578_ & ~new_n2029_;
  assign new_n2031_ = ~new_n578_ & new_n2030_;
  assign new_n2032_ = \V32(5)  & new_n583_;
  assign new_n2033_ = \V32(8)  & ~new_n583_;
  assign new_n2034_ = ~new_n583_ & new_n2033_;
  assign new_n2035_ = ~new_n2032_ & ~new_n2034_;
  assign new_n2036_ = new_n578_ & ~new_n2035_;
  assign new_n2037_ = new_n578_ & new_n2036_;
  assign new_n2038_ = ~new_n2031_ & ~new_n2037_;
  assign new_n2039_ = ~new_n662_ & ~new_n2038_;
  assign new_n2040_ = new_n661_ & new_n2039_;
  assign new_n2041_ = \V84(1)  & new_n662_;
  assign new_n2042_ = ~new_n661_ & new_n2041_;
  assign \V1243(3)  = new_n2040_ | new_n2042_;
  assign new_n2044_ = \V802(0)  & \V1243(3) ;
  assign new_n2045_ = new_n538_ & new_n2044_;
  assign new_n2046_ = new_n1865_ & new_n2045_;
  assign new_n2047_ = ~new_n1866_ & new_n2046_;
  assign new_n2048_ = ~new_n2006_ & ~new_n2015_;
  assign \V572(3)  = new_n2047_ | ~new_n2048_;
  assign new_n2050_ = \V149(6)  & \V802(0) ;
  assign new_n2051_ = new_n537_ & new_n2050_;
  assign new_n2052_ = new_n1865_ & new_n2051_;
  assign new_n2053_ = ~new_n1871_ & new_n2052_;
  assign new_n2054_ = \V194(4)  & new_n1409_;
  assign new_n2055_ = \V199(1)  & new_n2054_;
  assign new_n2056_ = \V199(3)  & new_n2055_;
  assign new_n2057_ = \V194(2)  & ~new_n2056_;
  assign new_n2058_ = ~\V194(2)  & new_n2056_;
  assign new_n2059_ = ~new_n2057_ & ~new_n2058_;
  assign new_n2060_ = ~new_n1866_ & ~new_n2059_;
  assign new_n2061_ = ~new_n1865_ & new_n2060_;
  assign new_n2062_ = ~new_n1871_ & new_n2061_;
  assign new_n2063_ = \V234(2)  & ~new_n545_;
  assign new_n2064_ = new_n567_ & new_n2063_;
  assign new_n2065_ = \V194(2)  & new_n545_;
  assign new_n2066_ = ~new_n567_ & new_n2065_;
  assign new_n2067_ = ~new_n2064_ & ~new_n2066_;
  assign new_n2068_ = new_n534_ & ~new_n2067_;
  assign new_n2069_ = ~new_n542_ & new_n2068_;
  assign new_n2070_ = ~new_n557_ & new_n2069_;
  assign new_n2071_ = ~\V59(0)  & \V149(6) ;
  assign new_n2072_ = ~new_n540_ & new_n2071_;
  assign new_n2073_ = new_n537_ & new_n2072_;
  assign new_n2074_ = new_n534_ & new_n2073_;
  assign new_n2075_ = new_n557_ & new_n2074_;
  assign new_n2076_ = ~new_n2070_ & ~new_n2075_;
  assign new_n2077_ = ~new_n578_ & ~new_n2076_;
  assign new_n2078_ = ~new_n578_ & new_n2077_;
  assign new_n2079_ = \V32(4)  & new_n583_;
  assign new_n2080_ = \V32(7)  & ~new_n583_;
  assign new_n2081_ = ~new_n583_ & new_n2080_;
  assign new_n2082_ = ~new_n2079_ & ~new_n2081_;
  assign new_n2083_ = new_n578_ & ~new_n2082_;
  assign new_n2084_ = new_n578_ & new_n2083_;
  assign new_n2085_ = ~new_n2078_ & ~new_n2084_;
  assign new_n2086_ = ~new_n662_ & ~new_n2085_;
  assign new_n2087_ = new_n661_ & new_n2086_;
  assign new_n2088_ = \V84(0)  & new_n662_;
  assign new_n2089_ = ~new_n661_ & new_n2088_;
  assign \V1243(2)  = new_n2087_ | new_n2089_;
  assign new_n2091_ = \V802(0)  & \V1243(2) ;
  assign new_n2092_ = new_n538_ & new_n2091_;
  assign new_n2093_ = new_n1865_ & new_n2092_;
  assign new_n2094_ = ~new_n1866_ & new_n2093_;
  assign new_n2095_ = ~new_n2053_ & ~new_n2062_;
  assign \V572(2)  = new_n2094_ | ~new_n2095_;
  assign new_n2097_ = \V149(5)  & \V802(0) ;
  assign new_n2098_ = new_n537_ & new_n2097_;
  assign new_n2099_ = new_n1865_ & new_n2098_;
  assign new_n2100_ = ~new_n1871_ & new_n2099_;
  assign new_n2101_ = \V194(2)  & new_n1409_;
  assign new_n2102_ = \V194(4)  & new_n2101_;
  assign new_n2103_ = \V199(1)  & new_n2102_;
  assign new_n2104_ = \V199(3)  & new_n2103_;
  assign new_n2105_ = \V194(1)  & ~new_n2104_;
  assign new_n2106_ = ~\V194(1)  & new_n2104_;
  assign new_n2107_ = ~new_n2105_ & ~new_n2106_;
  assign new_n2108_ = ~new_n1866_ & ~new_n2107_;
  assign new_n2109_ = ~new_n1865_ & new_n2108_;
  assign new_n2110_ = ~new_n1871_ & new_n2109_;
  assign new_n2111_ = \V234(1)  & ~new_n545_;
  assign new_n2112_ = new_n567_ & new_n2111_;
  assign new_n2113_ = \V194(1)  & new_n545_;
  assign new_n2114_ = ~new_n567_ & new_n2113_;
  assign new_n2115_ = ~new_n2112_ & ~new_n2114_;
  assign new_n2116_ = new_n534_ & ~new_n2115_;
  assign new_n2117_ = ~new_n542_ & new_n2116_;
  assign new_n2118_ = ~new_n557_ & new_n2117_;
  assign new_n2119_ = ~\V59(0)  & \V149(5) ;
  assign new_n2120_ = ~new_n540_ & new_n2119_;
  assign new_n2121_ = new_n537_ & new_n2120_;
  assign new_n2122_ = new_n534_ & new_n2121_;
  assign new_n2123_ = new_n557_ & new_n2122_;
  assign new_n2124_ = ~new_n2118_ & ~new_n2123_;
  assign new_n2125_ = ~new_n578_ & ~new_n2124_;
  assign new_n2126_ = ~new_n578_ & new_n2125_;
  assign new_n2127_ = \V32(3)  & new_n583_;
  assign new_n2128_ = \V32(6)  & ~new_n583_;
  assign new_n2129_ = ~new_n583_ & new_n2128_;
  assign new_n2130_ = ~new_n2127_ & ~new_n2129_;
  assign new_n2131_ = new_n578_ & ~new_n2130_;
  assign new_n2132_ = new_n578_ & new_n2131_;
  assign new_n2133_ = ~new_n2126_ & ~new_n2132_;
  assign new_n2134_ = ~new_n662_ & ~new_n2133_;
  assign new_n2135_ = new_n661_ & new_n2134_;
  assign new_n2136_ = \V78(5)  & new_n662_;
  assign new_n2137_ = ~new_n661_ & new_n2136_;
  assign \V1243(1)  = new_n2135_ | new_n2137_;
  assign new_n2139_ = \V802(0)  & \V1243(1) ;
  assign new_n2140_ = new_n538_ & new_n2139_;
  assign new_n2141_ = new_n1865_ & new_n2140_;
  assign new_n2142_ = ~new_n1866_ & new_n2141_;
  assign new_n2143_ = ~new_n2100_ & ~new_n2110_;
  assign \V572(1)  = new_n2142_ | ~new_n2143_;
  assign new_n2145_ = \V149(4)  & \V802(0) ;
  assign new_n2146_ = new_n537_ & new_n2145_;
  assign new_n2147_ = new_n1865_ & new_n2146_;
  assign new_n2148_ = ~new_n1871_ & new_n2147_;
  assign new_n2149_ = \V194(0)  & ~new_n1414_;
  assign new_n2150_ = ~\V194(0)  & new_n1414_;
  assign new_n2151_ = ~new_n2149_ & ~new_n2150_;
  assign new_n2152_ = ~new_n1866_ & ~new_n2151_;
  assign new_n2153_ = ~new_n1865_ & new_n2152_;
  assign new_n2154_ = ~new_n1871_ & new_n2153_;
  assign new_n2155_ = \V802(0)  & ~\V321(2) ;
  assign new_n2156_ = new_n538_ & new_n2155_;
  assign new_n2157_ = new_n1865_ & new_n2156_;
  assign new_n2158_ = ~new_n1866_ & new_n2157_;
  assign new_n2159_ = ~new_n2148_ & ~new_n2154_;
  assign \V572(0)  = new_n2158_ | ~new_n2159_;
  assign new_n2161_ = \V802(0)  & ~new_n567_;
  assign V587 = ~\V243(0)  & ~new_n2161_;
  assign new_n2163_ = ~\V243(0)  & \V244(0) ;
  assign new_n2164_ = ~new_n2161_ & new_n2163_;
  assign new_n2165_ = \V243(0)  & ~\V244(0) ;
  assign new_n2166_ = ~new_n2161_ & new_n2165_;
  assign \V591(0)  = new_n2164_ | new_n2166_;
  assign new_n2168_ = \V245(0)  & ~new_n1307_;
  assign new_n2169_ = ~new_n2161_ & new_n2168_;
  assign new_n2170_ = ~\V245(0)  & new_n1307_;
  assign new_n2171_ = ~new_n2161_ & new_n2170_;
  assign \V597(0)  = new_n2169_ | new_n2171_;
  assign new_n2173_ = \V246(0)  & ~new_n1308_;
  assign new_n2174_ = ~new_n2161_ & new_n2173_;
  assign new_n2175_ = ~\V246(0)  & new_n1308_;
  assign new_n2176_ = ~new_n2161_ & new_n2175_;
  assign \V603(0)  = new_n2174_ | new_n2176_;
  assign new_n2178_ = \V247(0)  & ~new_n1309_;
  assign new_n2179_ = ~new_n2161_ & new_n2178_;
  assign new_n2180_ = ~\V247(0)  & new_n1309_;
  assign new_n2181_ = ~new_n2161_ & new_n2180_;
  assign \V609(0)  = new_n2179_ | new_n2181_;
  assign new_n2183_ = \V62(0)  & ~\V214(0) ;
  assign new_n2184_ = new_n1513_ & new_n2183_;
  assign new_n2185_ = ~new_n1311_ & new_n2184_;
  assign new_n2186_ = ~new_n1311_ & ~new_n1586_;
  assign new_n2187_ = new_n1626_ & new_n2186_;
  assign new_n2188_ = ~\V214(0)  & new_n2187_;
  assign new_n2189_ = ~new_n631_ & ~new_n1620_;
  assign new_n2190_ = \V59(0)  & ~\V214(0) ;
  assign new_n2191_ = ~new_n2189_ & new_n2190_;
  assign new_n2192_ = ~new_n1311_ & new_n2191_;
  assign new_n2193_ = ~new_n2185_ & ~new_n2188_;
  assign V620 = ~new_n2192_ & new_n2193_;
  assign new_n2195_ = ~\V45(0)  & \V41(0) ;
  assign new_n2196_ = \V45(0)  & ~\V41(0) ;
  assign new_n2197_ = ~new_n2195_ & ~new_n2196_;
  assign V621 = \V293(0)  & new_n2197_;
  assign new_n2199_ = \V274(0)  & ~\V202(0) ;
  assign new_n2200_ = ~\V271(0)  & new_n2199_;
  assign \V640(0)  = \V271(0)  | new_n2200_;
  assign new_n2202_ = \V274(0)  & ~\V640(0) ;
  assign new_n2203_ = \V271(0)  & ~new_n2200_;
  assign new_n2204_ = \V269(0)  & new_n2203_;
  assign \V634(0)  = ~new_n2202_ & ~new_n2204_;
  assign new_n2206_ = ~\V290(0)  & new_n1311_;
  assign new_n2207_ = \V165(7)  & new_n2206_;
  assign new_n2208_ = \V261(0)  & ~new_n1604_;
  assign new_n2209_ = ~\V802(0)  & new_n2208_;
  assign new_n2210_ = \V272(0)  & new_n2209_;
  assign new_n2211_ = ~\V275(0)  & new_n2210_;
  assign new_n2212_ = new_n540_ & new_n2211_;
  assign new_n2213_ = ~\V149(6)  & new_n1510_;
  assign new_n2214_ = ~new_n544_ & new_n2213_;
  assign new_n2215_ = new_n1586_ & new_n2214_;
  assign new_n2216_ = \V62(0)  & new_n2215_;
  assign new_n2217_ = ~new_n544_ & new_n627_;
  assign new_n2218_ = new_n1586_ & new_n2217_;
  assign new_n2219_ = \V59(0)  & new_n2218_;
  assign new_n2220_ = \V67(0)  & \V172(0) ;
  assign new_n2221_ = \V215(0)  & new_n2220_;
  assign new_n2222_ = ~new_n544_ & new_n1586_;
  assign new_n2223_ = ~new_n1509_ & new_n2222_;
  assign new_n2224_ = ~new_n2213_ & new_n2223_;
  assign new_n2225_ = ~new_n627_ & new_n2224_;
  assign new_n2226_ = \V59(0)  & ~new_n544_;
  assign new_n2227_ = new_n1586_ & new_n2226_;
  assign new_n2228_ = new_n1509_ & new_n2227_;
  assign new_n2229_ = ~new_n2221_ & ~new_n2225_;
  assign new_n2230_ = ~new_n2228_ & new_n2229_;
  assign new_n2231_ = ~new_n2216_ & ~new_n2219_;
  assign new_n2232_ = ~\V214(0)  & new_n2231_;
  assign new_n2233_ = new_n2230_ & new_n2232_;
  assign new_n2234_ = \V56(0)  & ~new_n566_;
  assign new_n2235_ = ~new_n540_ & ~new_n2234_;
  assign new_n2236_ = \V242(0)  & new_n2235_;
  assign new_n2237_ = ~\V802(0)  & new_n2236_;
  assign new_n2238_ = ~new_n567_ & new_n2237_;
  assign new_n2239_ = \V261(0)  & ~new_n540_;
  assign new_n2240_ = ~new_n1604_ & new_n2239_;
  assign new_n2241_ = ~\V802(0)  & new_n2240_;
  assign new_n2242_ = \V134(1)  & \V134(0) ;
  assign new_n2243_ = \V242(0)  & new_n2242_;
  assign new_n2244_ = ~\V802(0)  & new_n2243_;
  assign new_n2245_ = \V272(0)  & new_n2244_;
  assign new_n2246_ = ~\V275(0)  & new_n2245_;
  assign new_n2247_ = new_n540_ & new_n2246_;
  assign new_n2248_ = ~new_n2241_ & ~new_n2247_;
  assign new_n2249_ = ~new_n2212_ & new_n2233_;
  assign new_n2250_ = ~new_n2238_ & new_n2249_;
  assign new_n2251_ = new_n2248_ & new_n2250_;
  assign new_n2252_ = ~new_n1457_ & new_n2251_;
  assign new_n2253_ = ~\V302(0)  & ~new_n2207_;
  assign new_n2254_ = new_n2252_ & new_n2253_;
  assign new_n2255_ = \V70(0)  & ~new_n533_;
  assign new_n2256_ = V763 & new_n2255_;
  assign new_n2257_ = new_n2254_ & new_n2256_;
  assign V775 = \V14(0)  & new_n2257_;
  assign new_n2259_ = \V10(0)  & ~\V13(0) ;
  assign V779 = \V6(0)  & new_n2259_;
  assign new_n2261_ = \V56(0)  & ~new_n500_;
  assign new_n2262_ = ~\V174(0)  & new_n2261_;
  assign new_n2263_ = ~\V52(0)  & ~new_n2262_;
  assign new_n2264_ = \V12(0)  & ~new_n2263_;
  assign V781 = \V6(0)  & new_n2264_;
  assign V782 = \V7(0)  & new_n2259_;
  assign V783 = \V5(0)  & \V11(0) ;
  assign V784 = \V7(0)  & \V11(0) ;
  assign new_n2269_ = ~\V149(7)  & ~\V149(3) ;
  assign new_n2270_ = \V149(4)  & new_n2269_;
  assign new_n2271_ = new_n489_ & new_n2270_;
  assign new_n2272_ = \V149(5)  & new_n2271_;
  assign new_n2273_ = ~\V149(6)  & new_n2272_;
  assign new_n2274_ = \V149(3)  & new_n594_;
  assign new_n2275_ = new_n489_ & new_n2274_;
  assign new_n2276_ = ~\V149(4)  & new_n2275_;
  assign new_n2277_ = ~\V149(6)  & new_n2276_;
  assign new_n2278_ = \V149(6)  & new_n671_;
  assign new_n2279_ = ~new_n672_ & ~new_n2277_;
  assign new_n2280_ = new_n489_ & new_n2279_;
  assign new_n2281_ = \V149(3)  & new_n2280_;
  assign new_n2282_ = ~new_n2278_ & new_n2281_;
  assign new_n2283_ = ~\V149(4)  & new_n1574_;
  assign new_n2284_ = ~\V149(6)  & new_n2283_;
  assign new_n2285_ = ~new_n2273_ & ~new_n2282_;
  assign new_n2286_ = ~new_n2284_ & new_n2285_;
  assign new_n2287_ = ~\V302(0)  & ~new_n2286_;
  assign new_n2288_ = \V149(0)  & \V149(2) ;
  assign new_n2289_ = \V149(1)  & new_n2288_;
  assign new_n2290_ = \V149(0)  & ~\V149(1) ;
  assign new_n2291_ = \V149(2)  & new_n2290_;
  assign new_n2292_ = \V149(0)  & ~\V149(2) ;
  assign new_n2293_ = \V149(1)  & new_n2292_;
  assign new_n2294_ = ~new_n2289_ & ~new_n2291_;
  assign new_n2295_ = new_n2286_ & new_n2294_;
  assign new_n2296_ = ~new_n2293_ & new_n2295_;
  assign new_n2297_ = new_n534_ & ~new_n2287_;
  assign new_n2298_ = ~new_n2296_ & new_n2297_;
  assign new_n2299_ = \V290(0)  & ~new_n1311_;
  assign new_n2300_ = ~\V149(6)  & new_n493_;
  assign new_n2301_ = ~\V149(6)  & new_n1575_;
  assign new_n2302_ = ~\V59(0)  & ~new_n534_;
  assign new_n2303_ = ~\V259(0)  & new_n2302_;
  assign new_n2304_ = ~\V260(0)  & new_n2303_;
  assign new_n2305_ = \V258(0)  & new_n2304_;
  assign new_n2306_ = \V149(6)  & new_n2283_;
  assign new_n2307_ = ~\V149(6)  & new_n597_;
  assign new_n2308_ = ~\V149(6)  & new_n1502_;
  assign new_n2309_ = ~new_n1576_ & ~new_n2300_;
  assign new_n2310_ = ~new_n2301_ & new_n2309_;
  assign new_n2311_ = ~new_n2305_ & new_n2310_;
  assign new_n2312_ = ~new_n2306_ & new_n2311_;
  assign new_n2313_ = ~new_n2307_ & new_n2312_;
  assign new_n2314_ = ~new_n2308_ & new_n2313_;
  assign new_n2315_ = \V56(0)  & ~new_n2314_;
  assign new_n2316_ = \V65(0)  & new_n1513_;
  assign new_n2317_ = ~new_n1511_ & ~new_n1514_;
  assign new_n2318_ = \V62(0)  & ~new_n2317_;
  assign new_n2319_ = ~new_n2315_ & ~new_n2316_;
  assign new_n2320_ = ~new_n2318_ & new_n2319_;
  assign new_n2321_ = ~new_n1311_ & new_n2219_;
  assign new_n2322_ = \V290(0)  & new_n1311_;
  assign new_n2323_ = ~new_n1311_ & new_n2225_;
  assign new_n2324_ = ~new_n1311_ & new_n2228_;
  assign new_n2325_ = ~new_n2323_ & ~new_n2324_;
  assign new_n2326_ = ~new_n2216_ & ~new_n2321_;
  assign new_n2327_ = ~new_n2322_ & new_n2326_;
  assign \V1741(0)  = ~new_n2325_ | ~new_n2327_;
  assign new_n2329_ = ~new_n1457_ & ~new_n2320_;
  assign new_n2330_ = ~\V1741(0)  & new_n2329_;
  assign new_n2331_ = ~new_n1304_ & new_n2254_;
  assign new_n2332_ = ~new_n1604_ & ~new_n2331_;
  assign new_n2333_ = ~\V289(0)  & ~new_n2330_;
  assign new_n2334_ = ~\V302(0)  & ~new_n2299_;
  assign new_n2335_ = new_n2333_ & new_n2334_;
  assign new_n2336_ = ~\V214(0)  & ~new_n2332_;
  assign new_n2337_ = ~new_n2207_ & new_n2336_;
  assign new_n2338_ = new_n2335_ & new_n2337_;
  assign new_n2339_ = \V14(0)  & ~new_n2298_;
  assign \V798(0)  = ~new_n2338_ | ~new_n2339_;
  assign V801 = new_n500_ & new_n509_;
  assign new_n2342_ = \V802(0)  & new_n591_;
  assign new_n2343_ = ~\V279(0)  & ~new_n2342_;
  assign new_n2344_ = \V149(5)  & new_n2342_;
  assign \V821(0)  = new_n2343_ | new_n2344_;
  assign new_n2346_ = \V280(0)  & ~new_n2342_;
  assign new_n2347_ = \V279(0)  & new_n2346_;
  assign new_n2348_ = \V149(4)  & new_n2342_;
  assign new_n2349_ = ~\V280(0)  & new_n2343_;
  assign new_n2350_ = ~new_n2347_ & ~new_n2348_;
  assign \V826(0)  = new_n2349_ | ~new_n2350_;
  assign new_n2352_ = ~new_n500_ & new_n509_;
  assign new_n2353_ = \V56(0)  & V763;
  assign new_n2354_ = ~new_n500_ & new_n2353_;
  assign new_n2355_ = ~new_n2263_ & new_n2354_;
  assign new_n2356_ = \V802(0)  & ~new_n2298_;
  assign new_n2357_ = \V56(0)  & ~new_n2286_;
  assign new_n2358_ = ~new_n2356_ & ~new_n2357_;
  assign new_n2359_ = ~new_n2352_ & ~new_n2355_;
  assign new_n2360_ = new_n2358_ & new_n2359_;
  assign new_n2361_ = new_n2254_ & ~new_n2360_;
  assign V966 = \V14(0)  & new_n2361_;
  assign new_n2363_ = \V62(0)  & ~new_n534_;
  assign new_n2364_ = \V56(0)  & new_n2286_;
  assign new_n2365_ = new_n2314_ & new_n2364_;
  assign new_n2366_ = ~new_n2355_ & new_n2365_;
  assign new_n2367_ = new_n567_ & ~new_n591_;
  assign new_n2368_ = ~new_n1621_ & new_n2367_;
  assign new_n2369_ = \V59(0)  & ~new_n2368_;
  assign new_n2370_ = ~new_n2363_ & ~new_n2366_;
  assign new_n2371_ = ~new_n2369_ & new_n2370_;
  assign new_n2372_ = new_n2254_ & ~new_n2371_;
  assign V986 = \V14(0)  & new_n2372_;
  assign V1256 = \V2(0)  & new_n2259_;
  assign new_n2375_ = ~\V57(0)  & new_n1514_;
  assign new_n2376_ = ~new_n630_ & new_n647_;
  assign new_n2377_ = ~new_n538_ & new_n2376_;
  assign new_n2378_ = ~new_n591_ & new_n1429_;
  assign new_n2379_ = new_n626_ & new_n2378_;
  assign new_n2380_ = new_n2377_ & new_n2379_;
  assign new_n2381_ = \V57(0)  & ~new_n2380_;
  assign new_n2382_ = ~\V60(0)  & ~\V63(0) ;
  assign new_n2383_ = new_n598_ & ~new_n2382_;
  assign new_n2384_ = \V12(0)  & \V2(0) ;
  assign new_n2385_ = ~\V174(0)  & new_n2384_;
  assign new_n2386_ = ~new_n2375_ & new_n2385_;
  assign new_n2387_ = ~new_n2381_ & new_n2386_;
  assign new_n2388_ = ~new_n2383_ & new_n2387_;
  assign V1257 = ~\V35(0)  & new_n2388_;
  assign V1260 = \V11(0)  & \V3(0) ;
  assign V1261 = ~\V62(0)  & V1260;
  assign V1262 = \V4(0)  & new_n2259_;
  assign V1264 = \V12(0)  & \V4(0) ;
  assign V1265 = \V52(0)  & V1264;
  assign V1266 = \V11(0)  & \V4(0) ;
  assign V1267 = \V11(0)  & \V2(0) ;
  assign new_n2397_ = \V14(0)  & new_n2254_;
  assign new_n2398_ = new_n631_ & new_n2397_;
  assign new_n2399_ = \V62(0)  & new_n2398_;
  assign new_n2400_ = ~new_n538_ & ~new_n1621_;
  assign new_n2401_ = ~new_n537_ & ~new_n1426_;
  assign new_n2402_ = new_n2400_ & new_n2401_;
  assign new_n2403_ = ~new_n549_ & ~new_n1430_;
  assign new_n2404_ = ~new_n591_ & new_n2403_;
  assign new_n2405_ = new_n2402_ & new_n2404_;
  assign new_n2406_ = ~\V174(0)  & new_n499_;
  assign new_n2407_ = \V59(0)  & ~V1719;
  assign new_n2408_ = ~new_n1509_ & new_n2407_;
  assign new_n2409_ = new_n2405_ & new_n2408_;
  assign new_n2410_ = ~new_n2406_ & new_n2409_;
  assign new_n2411_ = ~new_n672_ & new_n2410_;
  assign new_n2412_ = new_n2254_ & new_n2411_;
  assign new_n2413_ = \V14(0)  & new_n2412_;
  assign \V1274(0)  = new_n2399_ | new_n2413_;
  assign new_n2415_ = \V56(0)  & new_n2308_;
  assign new_n2416_ = ~\V302(0)  & new_n544_;
  assign new_n2417_ = new_n599_ & new_n627_;
  assign new_n2418_ = ~new_n2213_ & ~new_n2417_;
  assign new_n2419_ = ~new_n1509_ & ~new_n2416_;
  assign new_n2420_ = new_n2418_ & new_n2419_;
  assign new_n2421_ = ~\V289(0)  & \V14(0) ;
  assign new_n2422_ = ~new_n2420_ & new_n2421_;
  assign new_n2423_ = new_n1586_ & new_n2422_;
  assign new_n2424_ = ~new_n1311_ & new_n2423_;
  assign new_n2425_ = new_n485_ & ~new_n1311_;
  assign new_n2426_ = new_n1586_ & new_n2425_;
  assign new_n2427_ = ~new_n2424_ & new_n2426_;
  assign new_n2428_ = ~new_n499_ & new_n2427_;
  assign new_n2429_ = new_n485_ & new_n2322_;
  assign new_n2430_ = ~new_n2428_ & ~new_n2429_;
  assign new_n2431_ = \V14(0)  & ~new_n2415_;
  assign new_n2432_ = \V213(0)  & new_n2431_;
  assign new_n2433_ = new_n2430_ & new_n2432_;
  assign new_n2434_ = new_n2430_ & new_n2433_;
  assign new_n2435_ = ~\V165(5)  & ~\V165(7) ;
  assign new_n2436_ = ~\V165(3)  & new_n2435_;
  assign new_n2437_ = ~\V165(4)  & new_n2436_;
  assign new_n2438_ = ~\V165(6)  & new_n2437_;
  assign new_n2439_ = ~new_n1586_ & ~new_n2438_;
  assign new_n2440_ = ~new_n2430_ & ~new_n2439_;
  assign new_n2441_ = ~new_n2430_ & new_n2440_;
  assign \V1281(0)  = new_n2434_ | new_n2441_;
  assign new_n2443_ = \V213(5)  & new_n2431_;
  assign new_n2444_ = ~new_n2429_ & new_n2443_;
  assign new_n2445_ = ~new_n2429_ & new_n2444_;
  assign new_n2446_ = \V165(7)  & new_n2429_;
  assign new_n2447_ = new_n2429_ & new_n2446_;
  assign \V1297(4)  = new_n2445_ | new_n2447_;
  assign new_n2449_ = \V213(4)  & new_n2431_;
  assign new_n2450_ = ~new_n2429_ & new_n2449_;
  assign new_n2451_ = ~new_n2429_ & new_n2450_;
  assign new_n2452_ = \V165(6)  & new_n2429_;
  assign new_n2453_ = new_n2429_ & new_n2452_;
  assign \V1297(3)  = new_n2451_ | new_n2453_;
  assign new_n2455_ = \V213(3)  & new_n2431_;
  assign new_n2456_ = ~new_n2429_ & new_n2455_;
  assign new_n2457_ = ~new_n2429_ & new_n2456_;
  assign new_n2458_ = \V165(5)  & new_n2429_;
  assign new_n2459_ = new_n2429_ & new_n2458_;
  assign \V1297(2)  = new_n2457_ | new_n2459_;
  assign new_n2461_ = \V213(2)  & new_n2431_;
  assign new_n2462_ = ~new_n2429_ & new_n2461_;
  assign new_n2463_ = ~new_n2429_ & new_n2462_;
  assign new_n2464_ = \V165(4)  & new_n2429_;
  assign new_n2465_ = new_n2429_ & new_n2464_;
  assign \V1297(1)  = new_n2463_ | new_n2465_;
  assign new_n2467_ = \V213(1)  & new_n2431_;
  assign new_n2468_ = ~new_n2429_ & new_n2467_;
  assign new_n2469_ = ~new_n2429_ & new_n2468_;
  assign new_n2470_ = \V165(3)  & new_n2429_;
  assign new_n2471_ = new_n2429_ & new_n2470_;
  assign \V1297(0)  = new_n2469_ | new_n2471_;
  assign new_n2473_ = ~new_n1514_ & new_n2397_;
  assign new_n2474_ = ~new_n2213_ & new_n2473_;
  assign new_n2475_ = ~new_n1440_ & new_n2474_;
  assign new_n2476_ = new_n534_ & new_n2475_;
  assign new_n2477_ = ~new_n1441_ & new_n2476_;
  assign new_n2478_ = new_n647_ & new_n2477_;
  assign new_n2479_ = ~new_n1511_ & new_n2478_;
  assign V1365 = \V62(0)  & new_n2479_;
  assign new_n2481_ = \V802(0)  & ~new_n566_;
  assign V1378 = V782 & new_n2481_;
  assign new_n2483_ = ~\V802(0)  & new_n1858_;
  assign new_n2484_ = ~\V802(0)  & new_n540_;
  assign new_n2485_ = \V248(0)  & ~\V802(0) ;
  assign new_n2486_ = ~new_n2241_ & ~new_n2483_;
  assign new_n2487_ = ~new_n566_ & new_n2486_;
  assign new_n2488_ = ~new_n2484_ & new_n2487_;
  assign new_n2489_ = ~new_n2485_ & new_n2488_;
  assign new_n2490_ = ~new_n2241_ & ~new_n2485_;
  assign new_n2491_ = ~new_n540_ & new_n2490_;
  assign new_n2492_ = ~\V802(0)  & new_n2491_;
  assign new_n2493_ = new_n549_ & new_n2492_;
  assign new_n2494_ = ~new_n1858_ & new_n2493_;
  assign new_n2495_ = ~new_n1864_ & ~new_n2489_;
  assign new_n2496_ = ~new_n2494_ & new_n2495_;
  assign V1380 = V782 & ~new_n2496_;
  assign new_n2498_ = \V802(0)  & ~new_n1580_;
  assign new_n2499_ = ~new_n591_ & ~new_n2498_;
  assign new_n2500_ = \V7(0)  & ~new_n2499_;
  assign V1382 = new_n2259_ & new_n2500_;
  assign new_n2502_ = \V56(0)  & ~new_n1311_;
  assign new_n2503_ = new_n1576_ & new_n2502_;
  assign new_n2504_ = ~new_n1584_ & new_n2503_;
  assign new_n2505_ = \V7(0)  & new_n2504_;
  assign V1384 = new_n2259_ & new_n2505_;
  assign new_n2507_ = ~\V56(0)  & ~\V50(0) ;
  assign new_n2508_ = ~\V62(0)  & new_n2507_;
  assign new_n2509_ = ~new_n534_ & ~new_n2508_;
  assign new_n2510_ = \V7(0)  & new_n2509_;
  assign V1386 = new_n2259_ & new_n2510_;
  assign new_n2512_ = V763 & new_n2397_;
  assign new_n2513_ = ~\V165(5)  & new_n2512_;
  assign new_n2514_ = \V165(3)  & new_n2513_;
  assign new_n2515_ = ~\V165(4)  & new_n2514_;
  assign new_n2516_ = \V165(6)  & new_n2515_;
  assign new_n2517_ = \V70(0)  & new_n2516_;
  assign new_n2518_ = ~new_n1513_ & new_n2397_;
  assign new_n2519_ = \V65(0)  & new_n2518_;
  assign new_n2520_ = ~new_n628_ & new_n2519_;
  assign \V1392(0)  = new_n2517_ | new_n2520_;
  assign V1426 = \V1(0)  & new_n2259_;
  assign V1428 = \V1(0)  & \V11(0) ;
  assign V1429 = \V1(0)  & \V12(0) ;
  assign new_n2525_ = \V66(0)  & new_n2254_;
  assign V1432 = \V14(0)  & new_n2525_;
  assign new_n2527_ = \V277(0)  & ~new_n538_;
  assign new_n2528_ = \V14(0)  & new_n2527_;
  assign \V1439(0)  = new_n2300_ | new_n2528_;
  assign \V1440(0)  = ~\V14(0)  | new_n540_;
  assign new_n2531_ = \V268(5)  & \V268(3) ;
  assign new_n2532_ = \V268(1)  & new_n2531_;
  assign new_n2533_ = \V268(2)  & new_n2532_;
  assign new_n2534_ = \V268(4)  & new_n2533_;
  assign new_n2535_ = \V268(0)  & new_n2534_;
  assign new_n2536_ = ~new_n2509_ & ~new_n2535_;
  assign new_n2537_ = \V14(0)  & new_n2536_;
  assign new_n2538_ = \V258(0)  & new_n2537_;
  assign new_n2539_ = \V14(0)  & ~new_n2536_;
  assign new_n2540_ = ~\V258(0)  & new_n2539_;
  assign \V1451(0)  = new_n2538_ | new_n2540_;
  assign new_n2542_ = ~\V258(0)  & new_n2509_;
  assign new_n2543_ = \V258(0)  & new_n2535_;
  assign new_n2544_ = ~new_n2542_ & ~new_n2543_;
  assign new_n2545_ = \V259(0)  & new_n2544_;
  assign new_n2546_ = \V14(0)  & new_n2545_;
  assign new_n2547_ = ~\V259(0)  & ~new_n2544_;
  assign new_n2548_ = \V14(0)  & new_n2547_;
  assign \V1459(0)  = new_n2546_ | new_n2548_;
  assign new_n2550_ = ~\V259(0)  & new_n2542_;
  assign new_n2551_ = \V259(0)  & new_n2543_;
  assign new_n2552_ = ~new_n2550_ & ~new_n2551_;
  assign new_n2553_ = \V260(0)  & new_n2552_;
  assign new_n2554_ = \V14(0)  & new_n2553_;
  assign new_n2555_ = ~\V260(0)  & ~new_n2552_;
  assign new_n2556_ = \V14(0)  & new_n2555_;
  assign \V1467(0)  = new_n2554_ | new_n2556_;
  assign new_n2558_ = \V14(0)  & ~new_n1503_;
  assign new_n2559_ = new_n2254_ & new_n2558_;
  assign V1470 = \V67(0)  & new_n2559_;
  assign new_n2561_ = \V802(0)  & \V1757(0) ;
  assign new_n2562_ = new_n544_ & new_n2561_;
  assign new_n2563_ = ~new_n544_ & \V1757(0) ;
  assign new_n2564_ = ~new_n1584_ & ~new_n2562_;
  assign \V1480(0)  = new_n2563_ | ~new_n2564_;
  assign new_n2566_ = ~\V214(0)  & \V216(0) ;
  assign new_n2567_ = ~\V70(0)  & ~\V68(0) ;
  assign new_n2568_ = ~\V66(0)  & new_n2567_;
  assign new_n2569_ = ~\V69(0)  & new_n2568_;
  assign new_n2570_ = \V215(0)  & \V14(0) ;
  assign new_n2571_ = ~new_n2569_ & new_n2570_;
  assign new_n2572_ = new_n2233_ & new_n2571_;
  assign \V1492(0)  = new_n2566_ | new_n2572_;
  assign new_n2574_ = \V56(0)  & ~new_n545_;
  assign new_n2575_ = \V171(0)  & new_n2574_;
  assign new_n2576_ = \V278(0)  & ~new_n567_;
  assign new_n2577_ = ~new_n2575_ & ~new_n2576_;
  assign new_n2578_ = \V177(0)  & new_n2577_;
  assign new_n2579_ = ~\V248(0)  & new_n2578_;
  assign new_n2580_ = ~new_n1585_ & new_n2579_;
  assign new_n2581_ = ~\V271(0)  & ~\V274(0) ;
  assign new_n2582_ = ~\V172(0)  & new_n1470_;
  assign new_n2583_ = ~new_n1646_ & ~new_n2580_;
  assign new_n2584_ = ~new_n2581_ & new_n2583_;
  assign new_n2585_ = ~new_n2582_ & new_n2584_;
  assign new_n2586_ = new_n544_ & new_n1586_;
  assign new_n2587_ = \V56(0)  & new_n544_;
  assign new_n2588_ = \V149(7)  & new_n2587_;
  assign new_n2589_ = ~new_n2586_ & ~new_n2588_;
  assign new_n2590_ = new_n2251_ & ~new_n2585_;
  assign \V1536(0)  = ~new_n2589_ | ~new_n2590_;
  assign new_n2592_ = new_n2251_ & \V1536(0) ;
  assign new_n2593_ = ~new_n1252_ & ~new_n1269_;
  assign new_n2594_ = ~new_n1235_ & new_n2593_;
  assign new_n2595_ = ~new_n1218_ & new_n2594_;
  assign new_n2596_ = ~new_n1097_ & new_n2595_;
  assign new_n2597_ = ~new_n1114_ & new_n2596_;
  assign new_n2598_ = ~new_n1131_ & new_n2597_;
  assign new_n2599_ = ~new_n1148_ & new_n2598_;
  assign new_n2600_ = ~\V1536(0)  & ~new_n2599_;
  assign \V1512(3)  = new_n2592_ | new_n2600_;
  assign new_n2602_ = new_n2251_ & ~new_n2261_;
  assign new_n2603_ = ~new_n2589_ & new_n2602_;
  assign new_n2604_ = \V1536(0)  & ~new_n2603_;
  assign new_n2605_ = ~new_n1173_ & ~new_n1269_;
  assign new_n2606_ = ~new_n1235_ & new_n2605_;
  assign new_n2607_ = ~new_n1207_ & new_n2606_;
  assign new_n2608_ = ~new_n1086_ & new_n2607_;
  assign new_n2609_ = ~new_n1114_ & new_n2608_;
  assign new_n2610_ = ~new_n916_ & new_n2609_;
  assign new_n2611_ = ~new_n1148_ & new_n2610_;
  assign new_n2612_ = ~\V1536(0)  & ~new_n2611_;
  assign \V1512(2)  = new_n2604_ | new_n2612_;
  assign new_n2614_ = new_n2251_ & new_n2261_;
  assign new_n2615_ = \V1536(0)  & ~new_n2614_;
  assign new_n2616_ = ~new_n1252_ & new_n2605_;
  assign new_n2617_ = ~new_n1190_ & new_n2616_;
  assign new_n2618_ = ~new_n1001_ & new_n2617_;
  assign new_n2619_ = ~new_n1131_ & new_n2618_;
  assign new_n2620_ = ~new_n916_ & new_n2619_;
  assign new_n2621_ = ~new_n1148_ & new_n2620_;
  assign new_n2622_ = ~\V1536(0)  & ~new_n2621_;
  assign \V1512(1)  = new_n2615_ | new_n2622_;
  assign new_n2624_ = \V68(0)  & new_n2254_;
  assign V1537 = \V14(0)  & new_n2624_;
  assign new_n2626_ = ~\V69(0)  & ~\V50(0) ;
  assign new_n2627_ = new_n2254_ & ~new_n2626_;
  assign V1539 = \V14(0)  & new_n2627_;
  assign new_n2629_ = ~\V239(4)  & ~\V802(0) ;
  assign new_n2630_ = new_n591_ & new_n2629_;
  assign new_n2631_ = ~new_n2498_ & new_n2630_;
  assign new_n2632_ = ~\V802(0)  & new_n591_;
  assign new_n2633_ = \V1243(9)  & ~new_n2632_;
  assign new_n2634_ = new_n2498_ & new_n2633_;
  assign \V1552(1)  = new_n2631_ | new_n2634_;
  assign new_n2636_ = \V239(4)  & ~\V239(3) ;
  assign new_n2637_ = ~\V239(4)  & \V239(3) ;
  assign new_n2638_ = ~new_n2636_ & ~new_n2637_;
  assign new_n2639_ = ~\V802(0)  & ~new_n2638_;
  assign new_n2640_ = new_n591_ & new_n2639_;
  assign new_n2641_ = ~new_n2498_ & new_n2640_;
  assign new_n2642_ = \V1243(8)  & ~new_n2632_;
  assign new_n2643_ = new_n2498_ & new_n2642_;
  assign \V1552(0)  = new_n2641_ | new_n2643_;
  assign new_n2645_ = \V132(1)  & new_n2301_;
  assign new_n2646_ = ~new_n2307_ & new_n2645_;
  assign \V1953(1)  = ~new_n2278_ & new_n2646_;
  assign new_n2648_ = \V132(0)  & new_n2301_;
  assign new_n2649_ = ~new_n2307_ & new_n2648_;
  assign new_n2650_ = ~new_n2278_ & new_n2649_;
  assign new_n2651_ = \V108(5)  & ~new_n2301_;
  assign new_n2652_ = ~new_n2307_ & new_n2651_;
  assign new_n2653_ = new_n2278_ & new_n2652_;
  assign \V1953(0)  = new_n2650_ | new_n2653_;
  assign new_n2655_ = \V1953(1)  & ~\V1953(0) ;
  assign new_n2656_ = ~\V1953(1)  & \V1953(0) ;
  assign new_n2657_ = ~new_n2655_ & ~new_n2656_;
  assign new_n2658_ = \V100(5)  & new_n2306_;
  assign new_n2659_ = ~new_n2308_ & new_n2658_;
  assign new_n2660_ = ~new_n2301_ & new_n2659_;
  assign new_n2661_ = ~new_n2277_ & new_n2660_;
  assign new_n2662_ = \V213(5)  & ~new_n2306_;
  assign new_n2663_ = new_n2308_ & new_n2662_;
  assign new_n2664_ = ~new_n2301_ & new_n2663_;
  assign new_n2665_ = ~new_n2277_ & new_n2664_;
  assign new_n2666_ = \V124(5)  & ~new_n2306_;
  assign new_n2667_ = ~new_n2308_ & new_n2666_;
  assign new_n2668_ = new_n2301_ & new_n2667_;
  assign new_n2669_ = ~new_n2277_ & new_n2668_;
  assign new_n2670_ = ~new_n2661_ & ~new_n2665_;
  assign \V1921(5)  = new_n2669_ | ~new_n2670_;
  assign new_n2672_ = \V100(4)  & new_n2306_;
  assign new_n2673_ = ~new_n2308_ & new_n2672_;
  assign new_n2674_ = ~new_n2301_ & new_n2673_;
  assign new_n2675_ = ~new_n2277_ & new_n2674_;
  assign new_n2676_ = \V213(4)  & ~new_n2306_;
  assign new_n2677_ = new_n2308_ & new_n2676_;
  assign new_n2678_ = ~new_n2301_ & new_n2677_;
  assign new_n2679_ = ~new_n2277_ & new_n2678_;
  assign new_n2680_ = \V124(4)  & ~new_n2306_;
  assign new_n2681_ = ~new_n2308_ & new_n2680_;
  assign new_n2682_ = new_n2301_ & new_n2681_;
  assign new_n2683_ = ~new_n2277_ & new_n2682_;
  assign new_n2684_ = \V108(4)  & ~new_n2306_;
  assign new_n2685_ = ~new_n2308_ & new_n2684_;
  assign new_n2686_ = ~new_n2301_ & new_n2685_;
  assign new_n2687_ = new_n2277_ & new_n2686_;
  assign new_n2688_ = ~new_n2683_ & ~new_n2687_;
  assign new_n2689_ = ~new_n2675_ & ~new_n2679_;
  assign \V1921(4)  = ~new_n2688_ | ~new_n2689_;
  assign new_n2691_ = \V1921(5)  & ~\V1921(4) ;
  assign new_n2692_ = ~\V1921(5)  & \V1921(4) ;
  assign new_n2693_ = ~new_n2691_ & ~new_n2692_;
  assign new_n2694_ = ~new_n2657_ & new_n2693_;
  assign new_n2695_ = new_n2657_ & ~new_n2693_;
  assign new_n2696_ = ~new_n2694_ & ~new_n2695_;
  assign new_n2697_ = \V100(3)  & new_n2306_;
  assign new_n2698_ = ~new_n2308_ & new_n2697_;
  assign new_n2699_ = ~new_n2301_ & new_n2698_;
  assign new_n2700_ = ~new_n2277_ & new_n2699_;
  assign new_n2701_ = \V213(3)  & ~new_n2306_;
  assign new_n2702_ = new_n2308_ & new_n2701_;
  assign new_n2703_ = ~new_n2301_ & new_n2702_;
  assign new_n2704_ = ~new_n2277_ & new_n2703_;
  assign new_n2705_ = \V124(3)  & ~new_n2306_;
  assign new_n2706_ = ~new_n2308_ & new_n2705_;
  assign new_n2707_ = new_n2301_ & new_n2706_;
  assign new_n2708_ = ~new_n2277_ & new_n2707_;
  assign new_n2709_ = \V108(3)  & ~new_n2306_;
  assign new_n2710_ = ~new_n2308_ & new_n2709_;
  assign new_n2711_ = ~new_n2301_ & new_n2710_;
  assign new_n2712_ = new_n2277_ & new_n2711_;
  assign new_n2713_ = ~new_n2708_ & ~new_n2712_;
  assign new_n2714_ = ~new_n2700_ & ~new_n2704_;
  assign \V1921(3)  = ~new_n2713_ | ~new_n2714_;
  assign new_n2716_ = \V100(2)  & new_n2306_;
  assign new_n2717_ = ~new_n2308_ & new_n2716_;
  assign new_n2718_ = ~new_n2301_ & new_n2717_;
  assign new_n2719_ = ~new_n2277_ & new_n2718_;
  assign new_n2720_ = \V213(2)  & ~new_n2306_;
  assign new_n2721_ = new_n2308_ & new_n2720_;
  assign new_n2722_ = ~new_n2301_ & new_n2721_;
  assign new_n2723_ = ~new_n2277_ & new_n2722_;
  assign new_n2724_ = \V124(2)  & ~new_n2306_;
  assign new_n2725_ = ~new_n2308_ & new_n2724_;
  assign new_n2726_ = new_n2301_ & new_n2725_;
  assign new_n2727_ = ~new_n2277_ & new_n2726_;
  assign new_n2728_ = \V108(2)  & ~new_n2306_;
  assign new_n2729_ = ~new_n2308_ & new_n2728_;
  assign new_n2730_ = ~new_n2301_ & new_n2729_;
  assign new_n2731_ = new_n2277_ & new_n2730_;
  assign new_n2732_ = ~new_n2727_ & ~new_n2731_;
  assign new_n2733_ = ~new_n2719_ & ~new_n2723_;
  assign \V1921(2)  = ~new_n2732_ | ~new_n2733_;
  assign new_n2735_ = \V1921(3)  & ~\V1921(2) ;
  assign new_n2736_ = ~\V1921(3)  & \V1921(2) ;
  assign new_n2737_ = ~new_n2735_ & ~new_n2736_;
  assign new_n2738_ = \V100(1)  & new_n2306_;
  assign new_n2739_ = ~new_n2308_ & new_n2738_;
  assign new_n2740_ = ~new_n2301_ & new_n2739_;
  assign new_n2741_ = ~new_n2277_ & new_n2740_;
  assign new_n2742_ = \V213(1)  & ~new_n2306_;
  assign new_n2743_ = new_n2308_ & new_n2742_;
  assign new_n2744_ = ~new_n2301_ & new_n2743_;
  assign new_n2745_ = ~new_n2277_ & new_n2744_;
  assign new_n2746_ = \V124(1)  & ~new_n2306_;
  assign new_n2747_ = ~new_n2308_ & new_n2746_;
  assign new_n2748_ = new_n2301_ & new_n2747_;
  assign new_n2749_ = ~new_n2277_ & new_n2748_;
  assign new_n2750_ = \V108(1)  & ~new_n2306_;
  assign new_n2751_ = ~new_n2308_ & new_n2750_;
  assign new_n2752_ = ~new_n2301_ & new_n2751_;
  assign new_n2753_ = new_n2277_ & new_n2752_;
  assign new_n2754_ = ~new_n2749_ & ~new_n2753_;
  assign new_n2755_ = ~new_n2741_ & ~new_n2745_;
  assign \V1921(1)  = ~new_n2754_ | ~new_n2755_;
  assign new_n2757_ = \V100(0)  & new_n2306_;
  assign new_n2758_ = ~new_n2308_ & new_n2757_;
  assign new_n2759_ = ~new_n2301_ & new_n2758_;
  assign new_n2760_ = ~new_n2277_ & new_n2759_;
  assign new_n2761_ = \V213(0)  & ~new_n2306_;
  assign new_n2762_ = new_n2308_ & new_n2761_;
  assign new_n2763_ = ~new_n2301_ & new_n2762_;
  assign new_n2764_ = ~new_n2277_ & new_n2763_;
  assign new_n2765_ = \V124(0)  & ~new_n2306_;
  assign new_n2766_ = ~new_n2308_ & new_n2765_;
  assign new_n2767_ = new_n2301_ & new_n2766_;
  assign new_n2768_ = ~new_n2277_ & new_n2767_;
  assign new_n2769_ = \V108(0)  & ~new_n2306_;
  assign new_n2770_ = ~new_n2308_ & new_n2769_;
  assign new_n2771_ = ~new_n2301_ & new_n2770_;
  assign new_n2772_ = new_n2277_ & new_n2771_;
  assign new_n2773_ = ~new_n2768_ & ~new_n2772_;
  assign new_n2774_ = ~new_n2760_ & ~new_n2764_;
  assign \V1921(0)  = ~new_n2773_ | ~new_n2774_;
  assign new_n2776_ = \V1921(1)  & ~\V1921(0) ;
  assign new_n2777_ = ~\V1921(1)  & \V1921(0) ;
  assign new_n2778_ = ~new_n2776_ & ~new_n2777_;
  assign new_n2779_ = ~new_n2737_ & new_n2778_;
  assign new_n2780_ = new_n2737_ & ~new_n2778_;
  assign new_n2781_ = ~new_n2779_ & ~new_n2780_;
  assign new_n2782_ = ~new_n2696_ & new_n2781_;
  assign new_n2783_ = new_n2696_ & ~new_n2781_;
  assign \V1613(0)  = ~new_n2782_ & ~new_n2783_;
  assign new_n2785_ = \V118(7)  & new_n2307_;
  assign new_n2786_ = new_n1628_ & new_n2785_;
  assign new_n2787_ = \V46(0)  & ~new_n2307_;
  assign new_n2788_ = ~new_n1628_ & new_n2787_;
  assign \V1960(1)  = new_n2786_ | new_n2788_;
  assign new_n2790_ = \V118(6)  & new_n2307_;
  assign new_n2791_ = new_n1628_ & new_n2790_;
  assign new_n2792_ = \V48(0)  & ~new_n2307_;
  assign new_n2793_ = ~new_n1628_ & new_n2792_;
  assign \V1960(0)  = new_n2791_ | new_n2793_;
  assign new_n2795_ = \V1960(1)  & ~\V1960(0) ;
  assign new_n2796_ = ~\V1960(1)  & \V1960(0) ;
  assign new_n2797_ = ~new_n2795_ & ~new_n2796_;
  assign new_n2798_ = \V132(7)  & new_n2301_;
  assign new_n2799_ = ~new_n2307_ & new_n2798_;
  assign new_n2800_ = ~new_n2278_ & new_n2799_;
  assign new_n2801_ = \V118(5)  & ~new_n2301_;
  assign new_n2802_ = new_n2307_ & new_n2801_;
  assign new_n2803_ = ~new_n2278_ & new_n2802_;
  assign \V1953(7)  = new_n2800_ | new_n2803_;
  assign new_n2805_ = \V132(6)  & new_n2301_;
  assign new_n2806_ = ~new_n2307_ & new_n2805_;
  assign new_n2807_ = ~new_n2278_ & new_n2806_;
  assign new_n2808_ = \V118(4)  & ~new_n2301_;
  assign new_n2809_ = new_n2307_ & new_n2808_;
  assign new_n2810_ = ~new_n2278_ & new_n2809_;
  assign \V1953(6)  = new_n2807_ | new_n2810_;
  assign new_n2812_ = \V1953(7)  & ~\V1953(6) ;
  assign new_n2813_ = ~\V1953(7)  & \V1953(6) ;
  assign new_n2814_ = ~new_n2812_ & ~new_n2813_;
  assign new_n2815_ = ~new_n2797_ & new_n2814_;
  assign new_n2816_ = new_n2797_ & ~new_n2814_;
  assign new_n2817_ = ~new_n2815_ & ~new_n2816_;
  assign new_n2818_ = \V132(5)  & new_n2301_;
  assign new_n2819_ = ~new_n2307_ & new_n2818_;
  assign new_n2820_ = ~new_n2278_ & new_n2819_;
  assign new_n2821_ = \V118(3)  & ~new_n2301_;
  assign new_n2822_ = new_n2307_ & new_n2821_;
  assign new_n2823_ = ~new_n2278_ & new_n2822_;
  assign \V1953(5)  = new_n2820_ | new_n2823_;
  assign new_n2825_ = \V132(4)  & new_n2301_;
  assign new_n2826_ = ~new_n2307_ & new_n2825_;
  assign new_n2827_ = ~new_n2278_ & new_n2826_;
  assign new_n2828_ = \V118(2)  & ~new_n2301_;
  assign new_n2829_ = new_n2307_ & new_n2828_;
  assign new_n2830_ = ~new_n2278_ & new_n2829_;
  assign \V1953(4)  = new_n2827_ | new_n2830_;
  assign new_n2832_ = \V1953(5)  & ~\V1953(4) ;
  assign new_n2833_ = ~\V1953(5)  & \V1953(4) ;
  assign new_n2834_ = ~new_n2832_ & ~new_n2833_;
  assign new_n2835_ = \V132(3)  & new_n2301_;
  assign new_n2836_ = ~new_n2307_ & new_n2835_;
  assign new_n2837_ = ~new_n2278_ & new_n2836_;
  assign new_n2838_ = \V118(1)  & ~new_n2301_;
  assign new_n2839_ = new_n2307_ & new_n2838_;
  assign new_n2840_ = ~new_n2278_ & new_n2839_;
  assign \V1953(3)  = new_n2837_ | new_n2840_;
  assign new_n2842_ = \V132(2)  & new_n2301_;
  assign new_n2843_ = ~new_n2307_ & new_n2842_;
  assign new_n2844_ = ~new_n2278_ & new_n2843_;
  assign new_n2845_ = \V118(0)  & ~new_n2301_;
  assign new_n2846_ = new_n2307_ & new_n2845_;
  assign new_n2847_ = ~new_n2278_ & new_n2846_;
  assign \V1953(2)  = new_n2844_ | new_n2847_;
  assign new_n2849_ = \V1953(3)  & ~\V1953(2) ;
  assign new_n2850_ = ~\V1953(3)  & \V1953(2) ;
  assign new_n2851_ = ~new_n2849_ & ~new_n2850_;
  assign new_n2852_ = ~new_n2834_ & new_n2851_;
  assign new_n2853_ = new_n2834_ & ~new_n2851_;
  assign new_n2854_ = ~new_n2852_ & ~new_n2853_;
  assign new_n2855_ = ~new_n2817_ & new_n2854_;
  assign new_n2856_ = new_n2817_ & ~new_n2854_;
  assign \V1613(1)  = ~new_n2855_ & ~new_n2856_;
  assign new_n2858_ = \V174(0)  & new_n1311_;
  assign new_n2859_ = ~\V302(0)  & \V292(0) ;
  assign new_n2860_ = \V174(0)  & ~new_n2251_;
  assign new_n2861_ = ~new_n2859_ & ~new_n2860_;
  assign new_n2862_ = ~new_n509_ & ~new_n2858_;
  assign \V1620(0)  = ~new_n2861_ | ~new_n2862_;
  assign new_n2864_ = \V62(0)  & \V91(1) ;
  assign new_n2865_ = \V59(0)  & \V91(0) ;
  assign new_n2866_ = ~new_n2864_ & ~new_n2865_;
  assign new_n2867_ = new_n1514_ & ~new_n2866_;
  assign new_n2868_ = ~\V294(0)  & ~new_n1513_;
  assign new_n2869_ = ~new_n1620_ & new_n2868_;
  assign new_n2870_ = new_n2197_ & ~new_n2867_;
  assign \V1629(0)  = new_n2869_ | ~new_n2870_;
  assign new_n2872_ = \V149(7)  & new_n1508_;
  assign new_n2873_ = ~new_n2424_ & ~new_n2872_;
  assign \V1645(0)  = new_n1523_ | ~new_n2873_;
  assign new_n2875_ = ~\V289(0)  & new_n534_;
  assign new_n2876_ = ~\V249(0)  & new_n2875_;
  assign new_n2877_ = ~new_n1609_ & new_n2876_;
  assign new_n2878_ = \V295(0)  & new_n2877_;
  assign \V1652(0)  = \V290(0)  | ~new_n2878_;
  assign new_n2880_ = ~\V59(0)  & ~\V259(0) ;
  assign new_n2881_ = ~\V260(0)  & new_n2880_;
  assign new_n2882_ = \V258(0)  & new_n2881_;
  assign new_n2883_ = \V14(0)  & \V262(0) ;
  assign new_n2884_ = ~new_n2882_ & new_n2883_;
  assign new_n2885_ = \V262(0)  & new_n2884_;
  assign new_n2886_ = new_n533_ & ~new_n2885_;
  assign new_n2887_ = ~new_n2301_ & ~new_n2308_;
  assign new_n2888_ = ~new_n1576_ & new_n2886_;
  assign new_n2889_ = new_n2887_ & new_n2888_;
  assign new_n2890_ = ~new_n2306_ & ~new_n2307_;
  assign new_n2891_ = ~new_n2300_ & new_n2890_;
  assign new_n2892_ = new_n2889_ & new_n2891_;
  assign new_n2893_ = ~\V289(0)  & new_n2892_;
  assign new_n2894_ = \V1741(0)  & new_n2893_;
  assign new_n2895_ = new_n2317_ & new_n2892_;
  assign new_n2896_ = new_n2886_ & new_n2895_;
  assign new_n2897_ = ~new_n1513_ & new_n2896_;
  assign new_n2898_ = ~\V289(0)  & new_n2320_;
  assign new_n2899_ = new_n2251_ & new_n2898_;
  assign new_n2900_ = ~new_n2897_ & new_n2899_;
  assign new_n2901_ = ~new_n2207_ & new_n2900_;
  assign new_n2902_ = ~\V289(0)  & new_n1457_;
  assign new_n2903_ = ~\V802(0)  & new_n2902_;
  assign new_n2904_ = ~new_n1504_ & ~new_n2894_;
  assign new_n2905_ = ~new_n2901_ & new_n2904_;
  assign V1669 = ~new_n2903_ & new_n2905_;
  assign \V1679(0)  = ~new_n533_ | new_n2884_;
  assign new_n2908_ = \V56(0)  & new_n2306_;
  assign new_n2909_ = ~new_n487_ & ~new_n489_;
  assign new_n2910_ = new_n1311_ & ~new_n2909_;
  assign new_n2911_ = \V290(0)  & new_n2910_;
  assign new_n2912_ = ~new_n1311_ & ~new_n2909_;
  assign new_n2913_ = new_n1586_ & new_n2912_;
  assign new_n2914_ = ~new_n2424_ & new_n2913_;
  assign new_n2915_ = ~new_n499_ & new_n2914_;
  assign new_n2916_ = ~new_n2911_ & ~new_n2915_;
  assign new_n2917_ = \V14(0)  & ~new_n2908_;
  assign new_n2918_ = \V100(0)  & new_n2917_;
  assign new_n2919_ = new_n2916_ & new_n2918_;
  assign new_n2920_ = new_n2916_ & new_n2919_;
  assign new_n2921_ = ~new_n2439_ & ~new_n2916_;
  assign new_n2922_ = ~new_n2916_ & new_n2921_;
  assign \V1693(0)  = new_n2920_ | new_n2922_;
  assign new_n2924_ = \V100(5)  & new_n2917_;
  assign new_n2925_ = ~new_n2911_ & new_n2924_;
  assign new_n2926_ = ~new_n2911_ & new_n2925_;
  assign new_n2927_ = \V165(7)  & new_n2911_;
  assign new_n2928_ = new_n2911_ & new_n2927_;
  assign \V1709(4)  = new_n2926_ | new_n2928_;
  assign new_n2930_ = \V100(4)  & new_n2917_;
  assign new_n2931_ = ~new_n2911_ & new_n2930_;
  assign new_n2932_ = ~new_n2911_ & new_n2931_;
  assign new_n2933_ = \V165(6)  & new_n2911_;
  assign new_n2934_ = new_n2911_ & new_n2933_;
  assign \V1709(3)  = new_n2932_ | new_n2934_;
  assign new_n2936_ = \V100(3)  & new_n2917_;
  assign new_n2937_ = ~new_n2911_ & new_n2936_;
  assign new_n2938_ = ~new_n2911_ & new_n2937_;
  assign new_n2939_ = \V165(5)  & new_n2911_;
  assign new_n2940_ = new_n2911_ & new_n2939_;
  assign \V1709(2)  = new_n2938_ | new_n2940_;
  assign new_n2942_ = \V100(2)  & new_n2917_;
  assign new_n2943_ = ~new_n2911_ & new_n2942_;
  assign new_n2944_ = ~new_n2911_ & new_n2943_;
  assign new_n2945_ = \V165(4)  & new_n2911_;
  assign new_n2946_ = new_n2911_ & new_n2945_;
  assign \V1709(1)  = new_n2944_ | new_n2946_;
  assign new_n2948_ = \V100(1)  & new_n2917_;
  assign new_n2949_ = ~new_n2911_ & new_n2948_;
  assign new_n2950_ = ~new_n2911_ & new_n2949_;
  assign new_n2951_ = \V165(3)  & new_n2911_;
  assign new_n2952_ = new_n2911_ & new_n2951_;
  assign \V1709(0)  = new_n2950_ | new_n2952_;
  assign new_n2954_ = ~\V280(0)  & new_n591_;
  assign new_n2955_ = ~new_n1304_ & ~new_n1311_;
  assign new_n2956_ = new_n2254_ & new_n2955_;
  assign new_n2957_ = ~new_n2954_ & new_n2956_;
  assign new_n2958_ = \V240(0)  & new_n2957_;
  assign new_n2959_ = ~\V172(0)  & new_n2958_;
  assign new_n2960_ = ~new_n591_ & ~new_n1421_;
  assign new_n2961_ = \V802(0)  & ~new_n2960_;
  assign \V1717(0)  = new_n2959_ | new_n2961_;
  assign new_n2963_ = \V14(0)  & \V242(0) ;
  assign new_n2964_ = new_n566_ & new_n2963_;
  assign new_n2965_ = ~new_n567_ & new_n1858_;
  assign new_n2966_ = ~\V1536(0)  & new_n2965_;
  assign \V1726(0)  = new_n2964_ | new_n2966_;
  assign new_n2968_ = new_n1604_ & new_n2902_;
  assign new_n2969_ = ~\V802(0)  & new_n2968_;
  assign V1736 = ~\V290(0)  & new_n2969_;
  assign new_n2971_ = \V33(0)  & ~new_n499_;
  assign new_n2972_ = \V289(0)  & new_n2971_;
  assign \V1745(0)  = new_n485_ | ~new_n2972_;
  assign new_n2974_ = \V16(0)  & ~\V15(0) ;
  assign \V1758(0)  = new_n1474_ | new_n2974_;
  assign new_n2976_ = new_n485_ & new_n2974_;
  assign new_n2977_ = new_n487_ & new_n2974_;
  assign new_n2978_ = \V56(0)  & new_n2278_;
  assign new_n2979_ = \V101(0)  & ~new_n2978_;
  assign new_n2980_ = \V14(0)  & new_n2979_;
  assign new_n2981_ = ~new_n2976_ & ~new_n2977_;
  assign \V1759(0)  = new_n2980_ | ~new_n2981_;
  assign new_n2983_ = ~\V88(3)  & new_n598_;
  assign new_n2984_ = new_n598_ & new_n2983_;
  assign new_n2985_ = ~\V134(1)  & ~new_n598_;
  assign new_n2986_ = ~new_n598_ & new_n2985_;
  assign \V1771(1)  = new_n2984_ | new_n2986_;
  assign new_n2988_ = ~\V88(2)  & new_n598_;
  assign new_n2989_ = new_n598_ & new_n2988_;
  assign new_n2990_ = ~\V134(0)  & ~new_n598_;
  assign new_n2991_ = ~new_n598_ & new_n2990_;
  assign \V1771(0)  = new_n2989_ | new_n2991_;
  assign new_n2993_ = ~new_n598_ & ~\V1213(11) ;
  assign new_n2994_ = ~new_n598_ & new_n2993_;
  assign new_n2995_ = ~\V78(3)  & new_n598_;
  assign new_n2996_ = new_n598_ & new_n2995_;
  assign \V1781(1)  = new_n2994_ | new_n2996_;
  assign new_n2998_ = ~new_n598_ & ~\V1213(10) ;
  assign new_n2999_ = ~new_n598_ & new_n2998_;
  assign new_n3000_ = ~\V78(2)  & new_n598_;
  assign new_n3001_ = new_n598_ & new_n3000_;
  assign \V1781(0)  = new_n2999_ | new_n3001_;
  assign new_n3003_ = \V37(0)  & ~\V1243(9) ;
  assign new_n3004_ = \V37(0)  & new_n3003_;
  assign new_n3005_ = ~\V37(0)  & \V321(2) ;
  assign new_n3006_ = ~\V37(0)  & new_n3005_;
  assign \V1829(9)  = new_n3004_ | new_n3006_;
  assign new_n3008_ = \V37(0)  & ~\V1243(8) ;
  assign new_n3009_ = \V37(0)  & new_n3008_;
  assign new_n3010_ = ~\V37(0)  & ~\V1213(11) ;
  assign new_n3011_ = ~\V37(0)  & new_n3010_;
  assign \V1829(8)  = new_n3009_ | new_n3011_;
  assign new_n3013_ = \V37(0)  & ~\V1243(7) ;
  assign new_n3014_ = \V37(0)  & new_n3013_;
  assign new_n3015_ = ~\V37(0)  & ~\V1213(10) ;
  assign new_n3016_ = ~\V37(0)  & new_n3015_;
  assign \V1829(7)  = new_n3014_ | new_n3016_;
  assign new_n3018_ = \V37(0)  & ~\V1243(6) ;
  assign new_n3019_ = \V37(0)  & new_n3018_;
  assign new_n3020_ = ~\V37(0)  & ~\V1213(9) ;
  assign new_n3021_ = ~\V37(0)  & new_n3020_;
  assign \V1829(6)  = new_n3019_ | new_n3021_;
  assign new_n3023_ = \V37(0)  & ~\V1243(5) ;
  assign new_n3024_ = \V37(0)  & new_n3023_;
  assign new_n3025_ = ~\V37(0)  & ~\V1213(8) ;
  assign new_n3026_ = ~\V37(0)  & new_n3025_;
  assign \V1829(5)  = new_n3024_ | new_n3026_;
  assign new_n3028_ = \V37(0)  & ~\V1243(4) ;
  assign new_n3029_ = \V37(0)  & new_n3028_;
  assign new_n3030_ = ~\V37(0)  & ~\V1213(7) ;
  assign new_n3031_ = ~\V37(0)  & new_n3030_;
  assign \V1829(4)  = new_n3029_ | new_n3031_;
  assign new_n3033_ = \V37(0)  & ~\V1243(3) ;
  assign new_n3034_ = \V37(0)  & new_n3033_;
  assign new_n3035_ = ~\V37(0)  & ~\V1213(6) ;
  assign new_n3036_ = ~\V37(0)  & new_n3035_;
  assign \V1829(3)  = new_n3034_ | new_n3036_;
  assign new_n3038_ = \V37(0)  & ~\V1243(2) ;
  assign new_n3039_ = \V37(0)  & new_n3038_;
  assign new_n3040_ = ~\V37(0)  & ~\V1213(5) ;
  assign new_n3041_ = ~\V37(0)  & new_n3040_;
  assign \V1829(2)  = new_n3039_ | new_n3041_;
  assign new_n3043_ = \V37(0)  & ~\V1243(1) ;
  assign new_n3044_ = \V37(0)  & new_n3043_;
  assign new_n3045_ = ~\V37(0)  & ~\V1213(4) ;
  assign new_n3046_ = ~\V37(0)  & new_n3045_;
  assign \V1829(1)  = new_n3044_ | new_n3046_;
  assign new_n3048_ = \V37(0)  & ~\V1213(2) ;
  assign new_n3049_ = \V37(0)  & new_n3048_;
  assign \V1829(0)  = new_n3006_ | new_n3049_;
  assign new_n3051_ = \V262(0)  & ~new_n2884_;
  assign new_n3052_ = ~new_n2508_ & new_n3051_;
  assign new_n3053_ = \V261(0)  & ~new_n3052_;
  assign new_n3054_ = ~new_n2535_ & ~new_n3053_;
  assign V1832 = \V14(0)  & ~new_n3054_;
  assign new_n3056_ = \V56(0)  & new_n2277_;
  assign new_n3057_ = \V108(0)  & ~new_n3056_;
  assign new_n3058_ = ~new_n1584_ & ~new_n3057_;
  assign \V1896(0)  = new_n1475_ | ~new_n3058_;
  assign new_n3060_ = new_n538_ & new_n1584_;
  assign new_n3061_ = \V108(1)  & ~new_n3056_;
  assign \V1897(0)  = new_n3060_ | new_n3061_;
  assign new_n3063_ = new_n485_ & new_n2221_;
  assign new_n3064_ = \V108(2)  & ~new_n3056_;
  assign \V1898(0)  = new_n3063_ | new_n3064_;
  assign new_n3066_ = new_n487_ & new_n2221_;
  assign new_n3067_ = \V108(3)  & ~new_n3056_;
  assign \V1899(0)  = new_n3066_ | new_n3067_;
  assign new_n3069_ = \V108(4)  & ~new_n3056_;
  assign \V1900(0)  = new_n1474_ | new_n3069_;
  assign new_n3071_ = \V108(5)  & ~new_n2978_;
  assign \V1901(0)  = new_n2974_ | new_n3071_;
  assign new_n3073_ = ~\V108(4)  & new_n1474_;
  assign new_n3074_ = \V101(0)  & new_n3073_;
  assign new_n3075_ = \V56(0)  & new_n2307_;
  assign new_n3076_ = \V110(0)  & ~new_n3074_;
  assign new_n3077_ = ~new_n3075_ & new_n3076_;
  assign new_n3078_ = \V14(0)  & new_n3077_;
  assign new_n3079_ = ~\V102(0)  & ~\V1758(0) ;
  assign new_n3080_ = ~\V110(0)  & ~new_n3079_;
  assign new_n3081_ = new_n487_ & new_n3080_;
  assign \V1968(0)  = new_n3078_ | new_n3081_;
  assign new_n3083_ = ~new_n1860_ & ~new_n2481_;
  assign new_n3084_ = ~\V134(1)  & ~new_n2481_;
  assign new_n3085_ = new_n1860_ & new_n3084_;
  assign new_n3086_ = ~new_n3083_ & new_n3085_;
  assign new_n3087_ = new_n1860_ & ~new_n2481_;
  assign new_n3088_ = \V134(1)  & ~new_n1860_;
  assign new_n3089_ = ~new_n2481_ & new_n3088_;
  assign new_n3090_ = ~new_n3087_ & new_n3089_;
  assign \V1992(1)  = new_n3086_ | new_n3090_;
  assign new_n3092_ = \V134(1)  & ~\V134(0) ;
  assign new_n3093_ = ~\V134(1)  & \V134(0) ;
  assign new_n3094_ = ~new_n3092_ & ~new_n3093_;
  assign new_n3095_ = ~new_n2481_ & ~new_n3094_;
  assign new_n3096_ = new_n1860_ & new_n3095_;
  assign new_n3097_ = ~new_n3083_ & new_n3096_;
  assign new_n3098_ = \V134(0)  & ~new_n1860_;
  assign new_n3099_ = ~new_n2481_ & new_n3098_;
  assign new_n3100_ = ~new_n3087_ & new_n3099_;
  assign \V1992(0)  = new_n3097_ | new_n3100_;
  assign new_n3102_ = \V257(7)  & \V257(5) ;
  assign new_n3103_ = \V257(3)  & new_n3102_;
  assign new_n3104_ = \V257(1)  & new_n3103_;
  assign new_n3105_ = \V257(2)  & new_n3104_;
  assign new_n3106_ = \V257(4)  & new_n3105_;
  assign new_n3107_ = \V257(6)  & new_n3106_;
  assign new_n3108_ = \V257(0)  & ~new_n3107_;
  assign new_n3109_ = ~\V257(0)  & new_n3107_;
  assign V650 = new_n3108_ | new_n3109_;
  assign new_n3111_ = \V257(2)  & new_n3103_;
  assign new_n3112_ = \V257(4)  & new_n3111_;
  assign new_n3113_ = \V257(6)  & new_n3112_;
  assign new_n3114_ = \V257(1)  & ~new_n3113_;
  assign new_n3115_ = ~\V257(1)  & new_n3113_;
  assign V651 = new_n3114_ | new_n3115_;
  assign new_n3117_ = \V257(4)  & new_n3103_;
  assign new_n3118_ = \V257(6)  & new_n3117_;
  assign new_n3119_ = \V257(2)  & ~new_n3118_;
  assign new_n3120_ = ~\V257(2)  & new_n3118_;
  assign V652 = new_n3119_ | new_n3120_;
  assign new_n3122_ = \V257(4)  & new_n3102_;
  assign new_n3123_ = \V257(6)  & new_n3122_;
  assign new_n3124_ = \V257(3)  & ~new_n3123_;
  assign new_n3125_ = ~\V257(3)  & new_n3123_;
  assign V653 = new_n3124_ | new_n3125_;
  assign new_n3127_ = \V257(6)  & new_n3102_;
  assign new_n3128_ = \V257(4)  & ~new_n3127_;
  assign new_n3129_ = ~\V257(4)  & new_n3127_;
  assign V654 = new_n3128_ | new_n3129_;
  assign new_n3131_ = \V257(7)  & \V257(6) ;
  assign new_n3132_ = \V257(5)  & ~new_n3131_;
  assign new_n3133_ = ~\V257(5)  & new_n3131_;
  assign V655 = new_n3132_ | new_n3133_;
  assign new_n3135_ = ~\V257(7)  & \V257(6) ;
  assign new_n3136_ = \V257(7)  & ~\V257(6) ;
  assign V656 = new_n3135_ | new_n3136_;
  assign new_n3138_ = \V268(0)  & ~new_n2534_;
  assign new_n3139_ = ~\V268(0)  & new_n2534_;
  assign V1370 = new_n3138_ | new_n3139_;
  assign new_n3141_ = \V268(2)  & new_n2531_;
  assign new_n3142_ = \V268(4)  & new_n3141_;
  assign new_n3143_ = \V268(1)  & ~new_n3142_;
  assign new_n3144_ = ~\V268(1)  & new_n3142_;
  assign V1371 = new_n3143_ | new_n3144_;
  assign new_n3146_ = \V268(4)  & new_n2531_;
  assign new_n3147_ = \V268(2)  & ~new_n3146_;
  assign new_n3148_ = ~\V268(2)  & new_n3146_;
  assign V1372 = new_n3147_ | new_n3148_;
  assign new_n3150_ = \V268(5)  & \V268(4) ;
  assign new_n3151_ = \V268(3)  & ~new_n3150_;
  assign new_n3152_ = ~\V268(3)  & new_n3150_;
  assign V1373 = new_n3151_ | new_n3152_;
  assign new_n3154_ = ~\V268(5)  & \V268(4) ;
  assign new_n3155_ = \V268(5)  & ~\V268(4) ;
  assign V1374 = new_n3154_ | new_n3155_;
  assign \V585(0)  = ~\V34(0) ;
  assign V657 = ~\V257(7) ;
  assign \V1243(0)  = ~\V321(2) ;
  assign V1375 = ~\V268(5) ;
  assign \V1481(0)  = ~\V214(0) ;
  assign \V1495(0)  = ~\V175(0) ;
  assign \V1671(0)  = ~\V205(0) ;
  assign \V1760(0)  = ~\V101(0) ;
  assign \V1833(0)  = ~\V261(0) ;
  assign \V1863(0)  = ~\V301(0) ;
  assign \V1864(0)  = ~\V302(0) ;
endmodule


