// Benchmark "arbiter" written by ABC on Mon Sep 11 23:39:30 2023

module arbiter ( 
    \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ,
    \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] , \grant[5] ,
    \grant[6] , \grant[7] , \grant[8] , \grant[9] , \grant[10] ,
    \grant[11] , \grant[12] , \grant[13] , \grant[14] , \grant[15] ,
    \grant[16] , \grant[17] , \grant[18] , \grant[19] , \grant[20] ,
    \grant[21] , \grant[22] , \grant[23] , \grant[24] , \grant[25] ,
    \grant[26] , \grant[27] , \grant[28] , \grant[29] , \grant[30] ,
    \grant[31] , \grant[32] , \grant[33] , \grant[34] , \grant[35] ,
    \grant[36] , \grant[37] , \grant[38] , \grant[39] , \grant[40] ,
    \grant[41] , \grant[42] , \grant[43] , \grant[44] , \grant[45] ,
    \grant[46] , \grant[47] , \grant[48] , \grant[49] , \grant[50] ,
    \grant[51] , \grant[52] , \grant[53] , \grant[54] , \grant[55] ,
    \grant[56] , \grant[57] , \grant[58] , \grant[59] , \grant[60] ,
    \grant[61] , \grant[62] , \grant[63] , \grant[64] , \grant[65] ,
    \grant[66] , \grant[67] , \grant[68] , \grant[69] , \grant[70] ,
    \grant[71] , \grant[72] , \grant[73] , \grant[74] , \grant[75] ,
    \grant[76] , \grant[77] , \grant[78] , \grant[79] , \grant[80] ,
    \grant[81] , \grant[82] , \grant[83] , \grant[84] , \grant[85] ,
    \grant[86] , \grant[87] , \grant[88] , \grant[89] , \grant[90] ,
    \grant[91] , \grant[92] , \grant[93] , \grant[94] , \grant[95] ,
    \grant[96] , \grant[97] , \grant[98] , \grant[99] , \grant[100] ,
    \grant[101] , \grant[102] , \grant[103] , \grant[104] , \grant[105] ,
    \grant[106] , \grant[107] , \grant[108] , \grant[109] , \grant[110] ,
    \grant[111] , \grant[112] , \grant[113] , \grant[114] , \grant[115] ,
    \grant[116] , \grant[117] , \grant[118] , \grant[119] , \grant[120] ,
    \grant[121] , \grant[122] , \grant[123] , \grant[124] , \grant[125] ,
    \grant[126] , \grant[127] , anyGrant  );
  input  \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ;
  output \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] ,
    \grant[5] , \grant[6] , \grant[7] , \grant[8] , \grant[9] ,
    \grant[10] , \grant[11] , \grant[12] , \grant[13] , \grant[14] ,
    \grant[15] , \grant[16] , \grant[17] , \grant[18] , \grant[19] ,
    \grant[20] , \grant[21] , \grant[22] , \grant[23] , \grant[24] ,
    \grant[25] , \grant[26] , \grant[27] , \grant[28] , \grant[29] ,
    \grant[30] , \grant[31] , \grant[32] , \grant[33] , \grant[34] ,
    \grant[35] , \grant[36] , \grant[37] , \grant[38] , \grant[39] ,
    \grant[40] , \grant[41] , \grant[42] , \grant[43] , \grant[44] ,
    \grant[45] , \grant[46] , \grant[47] , \grant[48] , \grant[49] ,
    \grant[50] , \grant[51] , \grant[52] , \grant[53] , \grant[54] ,
    \grant[55] , \grant[56] , \grant[57] , \grant[58] , \grant[59] ,
    \grant[60] , \grant[61] , \grant[62] , \grant[63] , \grant[64] ,
    \grant[65] , \grant[66] , \grant[67] , \grant[68] , \grant[69] ,
    \grant[70] , \grant[71] , \grant[72] , \grant[73] , \grant[74] ,
    \grant[75] , \grant[76] , \grant[77] , \grant[78] , \grant[79] ,
    \grant[80] , \grant[81] , \grant[82] , \grant[83] , \grant[84] ,
    \grant[85] , \grant[86] , \grant[87] , \grant[88] , \grant[89] ,
    \grant[90] , \grant[91] , \grant[92] , \grant[93] , \grant[94] ,
    \grant[95] , \grant[96] , \grant[97] , \grant[98] , \grant[99] ,
    \grant[100] , \grant[101] , \grant[102] , \grant[103] , \grant[104] ,
    \grant[105] , \grant[106] , \grant[107] , \grant[108] , \grant[109] ,
    \grant[110] , \grant[111] , \grant[112] , \grant[113] , \grant[114] ,
    \grant[115] , \grant[116] , \grant[117] , \grant[118] , \grant[119] ,
    \grant[120] , \grant[121] , \grant[122] , \grant[123] , \grant[124] ,
    \grant[125] , \grant[126] , \grant[127] , anyGrant;
  wire new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2144_, new_n2145_,
    new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_,
    new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_,
    new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_,
    new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_,
    new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_,
    new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_,
    new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_,
    new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_,
    new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_,
    new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_,
    new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_,
    new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_,
    new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_,
    new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_,
    new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_,
    new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_,
    new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_,
    new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_,
    new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_,
    new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_,
    new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2408_, new_n2409_,
    new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_,
    new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_,
    new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_,
    new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2549_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_,
    new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_,
    new_n2565_, new_n2566_, new_n2567_, new_n2569_, new_n2570_, new_n2571_,
    new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_,
    new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2640_, new_n2641_,
    new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_,
    new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_,
    new_n2654_, new_n2655_, new_n2657_, new_n2658_, new_n2659_, new_n2660_,
    new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_,
    new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_,
    new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_,
    new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_,
    new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_,
    new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2799_, new_n2800_,
    new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_,
    new_n2813_, new_n2814_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2851_,
    new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2869_, new_n2870_,
    new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_,
    new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_,
    new_n2883_, new_n2884_, new_n2885_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_,
    new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_,
    new_n2966_, new_n2967_, new_n2968_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_,
    new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_,
    new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3017_, new_n3018_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_,
    new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3054_, new_n3055_,
    new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_,
    new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_,
    new_n3068_, new_n3069_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3104_, new_n3105_, new_n3106_,
    new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_,
    new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3136_, new_n3137_, new_n3138_,
    new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_,
    new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_,
    new_n3151_, new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_,
    new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_,
    new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_,
    new_n3202_, new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_,
    new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_,
    new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3238_, new_n3239_, new_n3240_,
    new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_,
    new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_,
    new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_,
    new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_,
    new_n3266_, new_n3267_, new_n3268_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3303_, new_n3304_,
    new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_,
    new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_,
    new_n3317_, new_n3318_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3354_, new_n3355_,
    new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_,
    new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_,
    new_n3368_, new_n3369_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3404_, new_n3405_, new_n3406_,
    new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_,
    new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3436_, new_n3437_, new_n3438_,
    new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_,
    new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_,
    new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3470_,
    new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_,
    new_n3483_, new_n3484_, new_n3485_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_,
    new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_,
    new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3538_, new_n3539_, new_n3540_,
    new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_,
    new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_,
    new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_,
    new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_,
    new_n3566_, new_n3567_, new_n3568_, new_n3570_, new_n3571_, new_n3572_,
    new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_,
    new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3603_, new_n3604_,
    new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_,
    new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_,
    new_n3617_, new_n3618_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_,
    new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_,
    new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3654_, new_n3655_,
    new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_,
    new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_,
    new_n3668_, new_n3669_, new_n3671_, new_n3672_, new_n3673_, new_n3674_,
    new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_,
    new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_,
    new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_,
    new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_,
    new_n3700_, new_n3701_, new_n3702_, new_n3704_, new_n3705_, new_n3706_,
    new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_,
    new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3736_, new_n3737_, new_n3738_,
    new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_,
    new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_,
    new_n3751_, new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_,
    new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_,
    new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3770_,
    new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_,
    new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_,
    new_n3783_, new_n3784_, new_n3785_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3802_, new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_,
    new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_,
    new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3838_, new_n3839_, new_n3840_,
    new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_,
    new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_,
    new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_,
    new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_,
    new_n3866_, new_n3867_, new_n3868_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_,
    new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3903_, new_n3904_,
    new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_,
    new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_,
    new_n3917_, new_n3918_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_,
    new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_,
    new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3954_, new_n3955_,
    new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_,
    new_n3968_, new_n3969_, new_n3971_, new_n3972_, new_n3973_, new_n3974_,
    new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_,
    new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_,
    new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_,
    new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_,
    new_n4000_, new_n4001_, new_n4002_, new_n4004_, new_n4005_, new_n4006_,
    new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_,
    new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4036_, new_n4037_, new_n4038_,
    new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_,
    new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_,
    new_n4051_, new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_,
    new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_,
    new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4070_,
    new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_,
    new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_,
    new_n4083_, new_n4084_, new_n4085_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_,
    new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_,
    new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4138_, new_n4139_, new_n4140_,
    new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4159_,
    new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_, new_n4165_,
    new_n4166_, new_n4167_, new_n4168_, new_n4170_, new_n4171_, new_n4172_,
    new_n4173_, new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_,
    new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_,
    new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_,
    new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_,
    new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4203_, new_n4204_,
    new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_,
    new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_,
    new_n4217_, new_n4218_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4254_, new_n4255_,
    new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_,
    new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_,
    new_n4268_, new_n4269_, new_n4271_, new_n4272_, new_n4273_, new_n4274_,
    new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_,
    new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_,
    new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4304_, new_n4305_, new_n4306_,
    new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_,
    new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4336_, new_n4337_, new_n4338_,
    new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_,
    new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_,
    new_n4351_, new_n4352_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4372_, new_n4373_, new_n4374_, new_n4375_, new_n4376_,
    new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_, new_n4382_,
    new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4389_,
    new_n4390_, new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_,
    new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_,
    new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_,
    new_n4408_;
  INV_X1     g0000(.I(\priority[4] ), .ZN(new_n386_));
  INV_X1     g0001(.I(\priority[5] ), .ZN(new_n387_));
  INV_X1     g0002(.I(\req[3] ), .ZN(new_n388_));
  NAND2_X1   g0003(.A1(new_n388_), .A2(\priority[3] ), .ZN(new_n389_));
  NAND3_X1   g0004(.A1(new_n389_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n390_));
  INV_X1     g0005(.I(\priority[1] ), .ZN(new_n391_));
  NOR2_X1    g0006(.A1(new_n391_), .A2(\req[1] ), .ZN(new_n392_));
  NOR2_X1    g0007(.A1(new_n392_), .A2(\priority[2] ), .ZN(new_n393_));
  NOR2_X1    g0008(.A1(\req[5] ), .A2(\req[6] ), .ZN(new_n394_));
  OAI21_X1   g0009(.A1(new_n387_), .A2(\req[4] ), .B(new_n394_), .ZN(new_n395_));
  NOR2_X1    g0010(.A1(\req[2] ), .A2(\req[3] ), .ZN(new_n396_));
  INV_X1     g0011(.I(new_n396_), .ZN(new_n397_));
  NOR4_X1    g0012(.A1(new_n390_), .A2(new_n393_), .A3(new_n395_), .A4(new_n397_), .ZN(new_n398_));
  INV_X1     g0013(.I(\priority[7] ), .ZN(new_n399_));
  INV_X1     g0014(.I(\priority[8] ), .ZN(new_n400_));
  INV_X1     g0015(.I(\req[6] ), .ZN(new_n401_));
  NAND2_X1   g0016(.A1(new_n401_), .A2(\priority[6] ), .ZN(new_n402_));
  NAND3_X1   g0017(.A1(new_n402_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n403_));
  INV_X1     g0018(.I(\priority[9] ), .ZN(new_n404_));
  NOR2_X1    g0019(.A1(new_n404_), .A2(\req[9] ), .ZN(new_n405_));
  NOR3_X1    g0020(.A1(new_n405_), .A2(\priority[10] ), .A3(\priority[11] ), .ZN(new_n406_));
  NOR2_X1    g0021(.A1(new_n400_), .A2(\req[7] ), .ZN(new_n407_));
  NOR2_X1    g0022(.A1(\req[8] ), .A2(\req[9] ), .ZN(new_n408_));
  INV_X1     g0023(.I(new_n408_), .ZN(new_n409_));
  NOR2_X1    g0024(.A1(new_n409_), .A2(new_n407_), .ZN(new_n410_));
  NAND3_X1   g0025(.A1(new_n406_), .A2(new_n410_), .A3(new_n403_), .ZN(new_n411_));
  INV_X1     g0026(.I(\priority[13] ), .ZN(new_n412_));
  INV_X1     g0027(.I(\priority[14] ), .ZN(new_n413_));
  INV_X1     g0028(.I(\req[12] ), .ZN(new_n414_));
  NAND2_X1   g0029(.A1(new_n414_), .A2(\priority[12] ), .ZN(new_n415_));
  NAND3_X1   g0030(.A1(new_n415_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n416_));
  NOR2_X1    g0031(.A1(\req[14] ), .A2(\req[15] ), .ZN(new_n417_));
  OAI21_X1   g0032(.A1(new_n413_), .A2(\req[13] ), .B(new_n417_), .ZN(new_n418_));
  INV_X1     g0033(.I(\priority[11] ), .ZN(new_n419_));
  NOR2_X1    g0034(.A1(new_n419_), .A2(\req[10] ), .ZN(new_n420_));
  NOR2_X1    g0035(.A1(\req[11] ), .A2(\req[12] ), .ZN(new_n421_));
  INV_X1     g0036(.I(new_n421_), .ZN(new_n422_));
  NOR2_X1    g0037(.A1(new_n422_), .A2(new_n420_), .ZN(new_n423_));
  NOR3_X1    g0038(.A1(new_n423_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n424_));
  OAI21_X1   g0039(.A1(new_n411_), .A2(new_n398_), .B(new_n424_), .ZN(new_n425_));
  INV_X1     g0040(.I(\priority[16] ), .ZN(new_n426_));
  INV_X1     g0041(.I(\priority[17] ), .ZN(new_n427_));
  INV_X1     g0042(.I(\req[15] ), .ZN(new_n428_));
  NAND2_X1   g0043(.A1(new_n428_), .A2(\priority[15] ), .ZN(new_n429_));
  NAND3_X1   g0044(.A1(new_n429_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n430_));
  INV_X1     g0045(.I(\priority[18] ), .ZN(new_n431_));
  NOR2_X1    g0046(.A1(new_n431_), .A2(\req[18] ), .ZN(new_n432_));
  NOR3_X1    g0047(.A1(new_n432_), .A2(\priority[19] ), .A3(\priority[20] ), .ZN(new_n433_));
  NOR2_X1    g0048(.A1(new_n427_), .A2(\req[16] ), .ZN(new_n434_));
  NOR2_X1    g0049(.A1(\req[17] ), .A2(\req[18] ), .ZN(new_n435_));
  INV_X1     g0050(.I(new_n435_), .ZN(new_n436_));
  NOR2_X1    g0051(.A1(new_n436_), .A2(new_n434_), .ZN(new_n437_));
  NAND3_X1   g0052(.A1(new_n433_), .A2(new_n437_), .A3(new_n430_), .ZN(new_n438_));
  INV_X1     g0053(.I(new_n438_), .ZN(new_n439_));
  INV_X1     g0054(.I(\priority[22] ), .ZN(new_n440_));
  INV_X1     g0055(.I(\priority[23] ), .ZN(new_n441_));
  INV_X1     g0056(.I(\req[21] ), .ZN(new_n442_));
  NAND2_X1   g0057(.A1(new_n442_), .A2(\priority[21] ), .ZN(new_n443_));
  NAND3_X1   g0058(.A1(new_n443_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n444_));
  NOR2_X1    g0059(.A1(\req[23] ), .A2(\req[24] ), .ZN(new_n445_));
  OAI21_X1   g0060(.A1(new_n441_), .A2(\req[22] ), .B(new_n445_), .ZN(new_n446_));
  INV_X1     g0061(.I(\priority[20] ), .ZN(new_n447_));
  NOR2_X1    g0062(.A1(new_n447_), .A2(\req[19] ), .ZN(new_n448_));
  NOR2_X1    g0063(.A1(\req[20] ), .A2(\req[21] ), .ZN(new_n449_));
  INV_X1     g0064(.I(new_n449_), .ZN(new_n450_));
  NOR2_X1    g0065(.A1(new_n450_), .A2(new_n448_), .ZN(new_n451_));
  NOR3_X1    g0066(.A1(new_n451_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n452_));
  INV_X1     g0067(.I(new_n452_), .ZN(new_n453_));
  AOI21_X1   g0068(.A1(new_n425_), .A2(new_n439_), .B(new_n453_), .ZN(new_n454_));
  INV_X1     g0069(.I(\priority[25] ), .ZN(new_n455_));
  INV_X1     g0070(.I(\priority[26] ), .ZN(new_n456_));
  INV_X1     g0071(.I(\req[24] ), .ZN(new_n457_));
  NAND2_X1   g0072(.A1(new_n457_), .A2(\priority[24] ), .ZN(new_n458_));
  NAND3_X1   g0073(.A1(new_n458_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n459_));
  INV_X1     g0074(.I(\priority[27] ), .ZN(new_n460_));
  NOR2_X1    g0075(.A1(new_n460_), .A2(\req[27] ), .ZN(new_n461_));
  NOR3_X1    g0076(.A1(new_n461_), .A2(\priority[28] ), .A3(\priority[29] ), .ZN(new_n462_));
  NOR2_X1    g0077(.A1(new_n456_), .A2(\req[25] ), .ZN(new_n463_));
  NOR2_X1    g0078(.A1(\req[26] ), .A2(\req[27] ), .ZN(new_n464_));
  INV_X1     g0079(.I(new_n464_), .ZN(new_n465_));
  NOR2_X1    g0080(.A1(new_n465_), .A2(new_n463_), .ZN(new_n466_));
  NAND3_X1   g0081(.A1(new_n462_), .A2(new_n466_), .A3(new_n459_), .ZN(new_n467_));
  INV_X1     g0082(.I(\priority[31] ), .ZN(new_n468_));
  INV_X1     g0083(.I(\priority[32] ), .ZN(new_n469_));
  INV_X1     g0084(.I(\req[30] ), .ZN(new_n470_));
  NAND2_X1   g0085(.A1(new_n470_), .A2(\priority[30] ), .ZN(new_n471_));
  NAND3_X1   g0086(.A1(new_n471_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n472_));
  NOR2_X1    g0087(.A1(\req[32] ), .A2(\req[33] ), .ZN(new_n473_));
  OAI21_X1   g0088(.A1(new_n469_), .A2(\req[31] ), .B(new_n473_), .ZN(new_n474_));
  INV_X1     g0089(.I(\priority[29] ), .ZN(new_n475_));
  NOR2_X1    g0090(.A1(new_n475_), .A2(\req[28] ), .ZN(new_n476_));
  NOR2_X1    g0091(.A1(\req[29] ), .A2(\req[30] ), .ZN(new_n477_));
  INV_X1     g0092(.I(new_n477_), .ZN(new_n478_));
  NOR2_X1    g0093(.A1(new_n478_), .A2(new_n476_), .ZN(new_n479_));
  NOR3_X1    g0094(.A1(new_n479_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n480_));
  OAI21_X1   g0095(.A1(new_n454_), .A2(new_n467_), .B(new_n480_), .ZN(new_n481_));
  INV_X1     g0096(.I(\priority[34] ), .ZN(new_n482_));
  INV_X1     g0097(.I(\priority[35] ), .ZN(new_n483_));
  INV_X1     g0098(.I(\req[33] ), .ZN(new_n484_));
  NAND2_X1   g0099(.A1(new_n484_), .A2(\priority[33] ), .ZN(new_n485_));
  NAND3_X1   g0100(.A1(new_n485_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n486_));
  INV_X1     g0101(.I(\priority[36] ), .ZN(new_n487_));
  NOR2_X1    g0102(.A1(new_n487_), .A2(\req[36] ), .ZN(new_n488_));
  NOR3_X1    g0103(.A1(new_n488_), .A2(\priority[37] ), .A3(\priority[38] ), .ZN(new_n489_));
  NOR2_X1    g0104(.A1(new_n483_), .A2(\req[34] ), .ZN(new_n490_));
  NOR2_X1    g0105(.A1(\req[35] ), .A2(\req[36] ), .ZN(new_n491_));
  INV_X1     g0106(.I(new_n491_), .ZN(new_n492_));
  NOR2_X1    g0107(.A1(new_n492_), .A2(new_n490_), .ZN(new_n493_));
  NAND3_X1   g0108(.A1(new_n489_), .A2(new_n493_), .A3(new_n486_), .ZN(new_n494_));
  INV_X1     g0109(.I(new_n494_), .ZN(new_n495_));
  INV_X1     g0110(.I(\priority[40] ), .ZN(new_n496_));
  INV_X1     g0111(.I(\priority[41] ), .ZN(new_n497_));
  INV_X1     g0112(.I(\req[39] ), .ZN(new_n498_));
  NAND2_X1   g0113(.A1(new_n498_), .A2(\priority[39] ), .ZN(new_n499_));
  NAND3_X1   g0114(.A1(new_n499_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n500_));
  NOR2_X1    g0115(.A1(\req[41] ), .A2(\req[42] ), .ZN(new_n501_));
  OAI21_X1   g0116(.A1(new_n497_), .A2(\req[40] ), .B(new_n501_), .ZN(new_n502_));
  INV_X1     g0117(.I(\priority[38] ), .ZN(new_n503_));
  NOR2_X1    g0118(.A1(new_n503_), .A2(\req[37] ), .ZN(new_n504_));
  NOR2_X1    g0119(.A1(\req[38] ), .A2(\req[39] ), .ZN(new_n505_));
  INV_X1     g0120(.I(new_n505_), .ZN(new_n506_));
  NOR2_X1    g0121(.A1(new_n506_), .A2(new_n504_), .ZN(new_n507_));
  NOR3_X1    g0122(.A1(new_n507_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n508_));
  INV_X1     g0123(.I(new_n508_), .ZN(new_n509_));
  AOI21_X1   g0124(.A1(new_n481_), .A2(new_n495_), .B(new_n509_), .ZN(new_n510_));
  INV_X1     g0125(.I(\priority[43] ), .ZN(new_n511_));
  INV_X1     g0126(.I(\priority[44] ), .ZN(new_n512_));
  INV_X1     g0127(.I(\req[42] ), .ZN(new_n513_));
  NAND2_X1   g0128(.A1(new_n513_), .A2(\priority[42] ), .ZN(new_n514_));
  NAND3_X1   g0129(.A1(new_n514_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n515_));
  INV_X1     g0130(.I(\priority[45] ), .ZN(new_n516_));
  NOR2_X1    g0131(.A1(new_n516_), .A2(\req[45] ), .ZN(new_n517_));
  NOR3_X1    g0132(.A1(new_n517_), .A2(\priority[46] ), .A3(\priority[47] ), .ZN(new_n518_));
  NOR2_X1    g0133(.A1(new_n512_), .A2(\req[43] ), .ZN(new_n519_));
  NOR2_X1    g0134(.A1(\req[44] ), .A2(\req[45] ), .ZN(new_n520_));
  INV_X1     g0135(.I(new_n520_), .ZN(new_n521_));
  NOR2_X1    g0136(.A1(new_n521_), .A2(new_n519_), .ZN(new_n522_));
  NAND3_X1   g0137(.A1(new_n518_), .A2(new_n522_), .A3(new_n515_), .ZN(new_n523_));
  INV_X1     g0138(.I(\priority[49] ), .ZN(new_n524_));
  INV_X1     g0139(.I(\priority[50] ), .ZN(new_n525_));
  INV_X1     g0140(.I(\req[48] ), .ZN(new_n526_));
  NAND2_X1   g0141(.A1(new_n526_), .A2(\priority[48] ), .ZN(new_n527_));
  NAND3_X1   g0142(.A1(new_n527_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n528_));
  NOR2_X1    g0143(.A1(\req[50] ), .A2(\req[51] ), .ZN(new_n529_));
  OAI21_X1   g0144(.A1(new_n525_), .A2(\req[49] ), .B(new_n529_), .ZN(new_n530_));
  INV_X1     g0145(.I(\priority[47] ), .ZN(new_n531_));
  NOR2_X1    g0146(.A1(new_n531_), .A2(\req[46] ), .ZN(new_n532_));
  NOR2_X1    g0147(.A1(\req[47] ), .A2(\req[48] ), .ZN(new_n533_));
  INV_X1     g0148(.I(new_n533_), .ZN(new_n534_));
  NOR2_X1    g0149(.A1(new_n534_), .A2(new_n532_), .ZN(new_n535_));
  NOR3_X1    g0150(.A1(new_n535_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n536_));
  OAI21_X1   g0151(.A1(new_n510_), .A2(new_n523_), .B(new_n536_), .ZN(new_n537_));
  INV_X1     g0152(.I(\priority[52] ), .ZN(new_n538_));
  INV_X1     g0153(.I(\priority[53] ), .ZN(new_n539_));
  INV_X1     g0154(.I(\req[51] ), .ZN(new_n540_));
  NAND2_X1   g0155(.A1(new_n540_), .A2(\priority[51] ), .ZN(new_n541_));
  NAND3_X1   g0156(.A1(new_n541_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n542_));
  INV_X1     g0157(.I(\priority[54] ), .ZN(new_n543_));
  NOR2_X1    g0158(.A1(new_n543_), .A2(\req[54] ), .ZN(new_n544_));
  NOR3_X1    g0159(.A1(new_n544_), .A2(\priority[55] ), .A3(\priority[56] ), .ZN(new_n545_));
  NOR2_X1    g0160(.A1(new_n539_), .A2(\req[52] ), .ZN(new_n546_));
  NOR2_X1    g0161(.A1(\req[53] ), .A2(\req[54] ), .ZN(new_n547_));
  INV_X1     g0162(.I(new_n547_), .ZN(new_n548_));
  NOR2_X1    g0163(.A1(new_n548_), .A2(new_n546_), .ZN(new_n549_));
  NAND3_X1   g0164(.A1(new_n545_), .A2(new_n549_), .A3(new_n542_), .ZN(new_n550_));
  INV_X1     g0165(.I(new_n550_), .ZN(new_n551_));
  INV_X1     g0166(.I(\priority[58] ), .ZN(new_n552_));
  INV_X1     g0167(.I(\priority[59] ), .ZN(new_n553_));
  INV_X1     g0168(.I(\req[57] ), .ZN(new_n554_));
  NAND2_X1   g0169(.A1(new_n554_), .A2(\priority[57] ), .ZN(new_n555_));
  NAND3_X1   g0170(.A1(new_n555_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n556_));
  NOR2_X1    g0171(.A1(\req[59] ), .A2(\req[60] ), .ZN(new_n557_));
  OAI21_X1   g0172(.A1(new_n553_), .A2(\req[58] ), .B(new_n557_), .ZN(new_n558_));
  INV_X1     g0173(.I(\priority[56] ), .ZN(new_n559_));
  NOR2_X1    g0174(.A1(new_n559_), .A2(\req[55] ), .ZN(new_n560_));
  NOR2_X1    g0175(.A1(\req[56] ), .A2(\req[57] ), .ZN(new_n561_));
  INV_X1     g0176(.I(new_n561_), .ZN(new_n562_));
  NOR2_X1    g0177(.A1(new_n562_), .A2(new_n560_), .ZN(new_n563_));
  NOR3_X1    g0178(.A1(new_n563_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n564_));
  INV_X1     g0179(.I(new_n564_), .ZN(new_n565_));
  AOI21_X1   g0180(.A1(new_n537_), .A2(new_n551_), .B(new_n565_), .ZN(new_n566_));
  INV_X1     g0181(.I(\priority[61] ), .ZN(new_n567_));
  INV_X1     g0182(.I(\priority[62] ), .ZN(new_n568_));
  INV_X1     g0183(.I(\req[60] ), .ZN(new_n569_));
  NAND2_X1   g0184(.A1(new_n569_), .A2(\priority[60] ), .ZN(new_n570_));
  NAND3_X1   g0185(.A1(new_n570_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n571_));
  INV_X1     g0186(.I(\priority[63] ), .ZN(new_n572_));
  NOR2_X1    g0187(.A1(new_n572_), .A2(\req[63] ), .ZN(new_n573_));
  NOR3_X1    g0188(.A1(new_n573_), .A2(\priority[64] ), .A3(\priority[65] ), .ZN(new_n574_));
  NOR2_X1    g0189(.A1(new_n568_), .A2(\req[61] ), .ZN(new_n575_));
  NOR2_X1    g0190(.A1(\req[62] ), .A2(\req[63] ), .ZN(new_n576_));
  INV_X1     g0191(.I(new_n576_), .ZN(new_n577_));
  NOR2_X1    g0192(.A1(new_n577_), .A2(new_n575_), .ZN(new_n578_));
  NAND3_X1   g0193(.A1(new_n574_), .A2(new_n578_), .A3(new_n571_), .ZN(new_n579_));
  INV_X1     g0194(.I(\priority[67] ), .ZN(new_n580_));
  INV_X1     g0195(.I(\priority[68] ), .ZN(new_n581_));
  INV_X1     g0196(.I(\req[66] ), .ZN(new_n582_));
  NAND2_X1   g0197(.A1(new_n582_), .A2(\priority[66] ), .ZN(new_n583_));
  NAND3_X1   g0198(.A1(new_n583_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n584_));
  NOR2_X1    g0199(.A1(\req[68] ), .A2(\req[69] ), .ZN(new_n585_));
  OAI21_X1   g0200(.A1(new_n581_), .A2(\req[67] ), .B(new_n585_), .ZN(new_n586_));
  INV_X1     g0201(.I(\priority[65] ), .ZN(new_n587_));
  NOR2_X1    g0202(.A1(new_n587_), .A2(\req[64] ), .ZN(new_n588_));
  NOR2_X1    g0203(.A1(\req[65] ), .A2(\req[66] ), .ZN(new_n589_));
  INV_X1     g0204(.I(new_n589_), .ZN(new_n590_));
  NOR2_X1    g0205(.A1(new_n590_), .A2(new_n588_), .ZN(new_n591_));
  NOR3_X1    g0206(.A1(new_n591_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n592_));
  OAI21_X1   g0207(.A1(new_n566_), .A2(new_n579_), .B(new_n592_), .ZN(new_n593_));
  INV_X1     g0208(.I(\priority[70] ), .ZN(new_n594_));
  INV_X1     g0209(.I(\priority[71] ), .ZN(new_n595_));
  INV_X1     g0210(.I(\req[69] ), .ZN(new_n596_));
  NAND2_X1   g0211(.A1(new_n596_), .A2(\priority[69] ), .ZN(new_n597_));
  NAND3_X1   g0212(.A1(new_n597_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n598_));
  INV_X1     g0213(.I(\priority[72] ), .ZN(new_n599_));
  NOR2_X1    g0214(.A1(new_n599_), .A2(\req[72] ), .ZN(new_n600_));
  NOR3_X1    g0215(.A1(new_n600_), .A2(\priority[73] ), .A3(\priority[74] ), .ZN(new_n601_));
  NOR2_X1    g0216(.A1(new_n595_), .A2(\req[70] ), .ZN(new_n602_));
  NOR2_X1    g0217(.A1(\req[71] ), .A2(\req[72] ), .ZN(new_n603_));
  INV_X1     g0218(.I(new_n603_), .ZN(new_n604_));
  NOR2_X1    g0219(.A1(new_n604_), .A2(new_n602_), .ZN(new_n605_));
  NAND3_X1   g0220(.A1(new_n601_), .A2(new_n605_), .A3(new_n598_), .ZN(new_n606_));
  INV_X1     g0221(.I(new_n606_), .ZN(new_n607_));
  INV_X1     g0222(.I(\priority[76] ), .ZN(new_n608_));
  INV_X1     g0223(.I(\priority[77] ), .ZN(new_n609_));
  INV_X1     g0224(.I(\req[75] ), .ZN(new_n610_));
  NAND2_X1   g0225(.A1(new_n610_), .A2(\priority[75] ), .ZN(new_n611_));
  NAND3_X1   g0226(.A1(new_n611_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n612_));
  NOR2_X1    g0227(.A1(\req[77] ), .A2(\req[78] ), .ZN(new_n613_));
  OAI21_X1   g0228(.A1(new_n609_), .A2(\req[76] ), .B(new_n613_), .ZN(new_n614_));
  INV_X1     g0229(.I(\priority[74] ), .ZN(new_n615_));
  NOR2_X1    g0230(.A1(new_n615_), .A2(\req[73] ), .ZN(new_n616_));
  NOR2_X1    g0231(.A1(\req[74] ), .A2(\req[75] ), .ZN(new_n617_));
  INV_X1     g0232(.I(new_n617_), .ZN(new_n618_));
  NOR2_X1    g0233(.A1(new_n618_), .A2(new_n616_), .ZN(new_n619_));
  NOR3_X1    g0234(.A1(new_n619_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n620_));
  INV_X1     g0235(.I(new_n620_), .ZN(new_n621_));
  AOI21_X1   g0236(.A1(new_n593_), .A2(new_n607_), .B(new_n621_), .ZN(new_n622_));
  INV_X1     g0237(.I(\priority[79] ), .ZN(new_n623_));
  INV_X1     g0238(.I(\priority[80] ), .ZN(new_n624_));
  INV_X1     g0239(.I(\req[78] ), .ZN(new_n625_));
  NAND2_X1   g0240(.A1(new_n625_), .A2(\priority[78] ), .ZN(new_n626_));
  NAND3_X1   g0241(.A1(new_n626_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n627_));
  INV_X1     g0242(.I(\priority[81] ), .ZN(new_n628_));
  NOR2_X1    g0243(.A1(new_n628_), .A2(\req[81] ), .ZN(new_n629_));
  NOR3_X1    g0244(.A1(new_n629_), .A2(\priority[82] ), .A3(\priority[83] ), .ZN(new_n630_));
  NOR2_X1    g0245(.A1(new_n624_), .A2(\req[79] ), .ZN(new_n631_));
  NOR2_X1    g0246(.A1(\req[80] ), .A2(\req[81] ), .ZN(new_n632_));
  INV_X1     g0247(.I(new_n632_), .ZN(new_n633_));
  NOR2_X1    g0248(.A1(new_n633_), .A2(new_n631_), .ZN(new_n634_));
  NAND3_X1   g0249(.A1(new_n630_), .A2(new_n634_), .A3(new_n627_), .ZN(new_n635_));
  INV_X1     g0250(.I(\priority[85] ), .ZN(new_n636_));
  INV_X1     g0251(.I(\priority[86] ), .ZN(new_n637_));
  INV_X1     g0252(.I(\req[84] ), .ZN(new_n638_));
  NAND2_X1   g0253(.A1(new_n638_), .A2(\priority[84] ), .ZN(new_n639_));
  NAND3_X1   g0254(.A1(new_n639_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n640_));
  NOR2_X1    g0255(.A1(\req[86] ), .A2(\req[87] ), .ZN(new_n641_));
  OAI21_X1   g0256(.A1(new_n637_), .A2(\req[85] ), .B(new_n641_), .ZN(new_n642_));
  INV_X1     g0257(.I(\priority[83] ), .ZN(new_n643_));
  NOR2_X1    g0258(.A1(new_n643_), .A2(\req[82] ), .ZN(new_n644_));
  NOR2_X1    g0259(.A1(\req[83] ), .A2(\req[84] ), .ZN(new_n645_));
  INV_X1     g0260(.I(new_n645_), .ZN(new_n646_));
  NOR2_X1    g0261(.A1(new_n646_), .A2(new_n644_), .ZN(new_n647_));
  NOR3_X1    g0262(.A1(new_n647_), .A2(new_n640_), .A3(new_n642_), .ZN(new_n648_));
  OAI21_X1   g0263(.A1(new_n622_), .A2(new_n635_), .B(new_n648_), .ZN(new_n649_));
  INV_X1     g0264(.I(\priority[88] ), .ZN(new_n650_));
  INV_X1     g0265(.I(\priority[89] ), .ZN(new_n651_));
  INV_X1     g0266(.I(\req[87] ), .ZN(new_n652_));
  NAND2_X1   g0267(.A1(new_n652_), .A2(\priority[87] ), .ZN(new_n653_));
  NAND3_X1   g0268(.A1(new_n653_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n654_));
  INV_X1     g0269(.I(\priority[90] ), .ZN(new_n655_));
  NOR2_X1    g0270(.A1(new_n655_), .A2(\req[90] ), .ZN(new_n656_));
  NOR3_X1    g0271(.A1(new_n656_), .A2(\priority[91] ), .A3(\priority[92] ), .ZN(new_n657_));
  NOR2_X1    g0272(.A1(new_n651_), .A2(\req[88] ), .ZN(new_n658_));
  NOR2_X1    g0273(.A1(\req[89] ), .A2(\req[90] ), .ZN(new_n659_));
  INV_X1     g0274(.I(new_n659_), .ZN(new_n660_));
  NOR2_X1    g0275(.A1(new_n660_), .A2(new_n658_), .ZN(new_n661_));
  NAND3_X1   g0276(.A1(new_n657_), .A2(new_n661_), .A3(new_n654_), .ZN(new_n662_));
  INV_X1     g0277(.I(new_n662_), .ZN(new_n663_));
  INV_X1     g0278(.I(\priority[94] ), .ZN(new_n664_));
  INV_X1     g0279(.I(\priority[95] ), .ZN(new_n665_));
  INV_X1     g0280(.I(\req[93] ), .ZN(new_n666_));
  NAND2_X1   g0281(.A1(new_n666_), .A2(\priority[93] ), .ZN(new_n667_));
  NAND3_X1   g0282(.A1(new_n667_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n668_));
  NOR2_X1    g0283(.A1(\req[95] ), .A2(\req[96] ), .ZN(new_n669_));
  OAI21_X1   g0284(.A1(new_n665_), .A2(\req[94] ), .B(new_n669_), .ZN(new_n670_));
  INV_X1     g0285(.I(\priority[92] ), .ZN(new_n671_));
  NOR2_X1    g0286(.A1(new_n671_), .A2(\req[91] ), .ZN(new_n672_));
  NOR2_X1    g0287(.A1(\req[92] ), .A2(\req[93] ), .ZN(new_n673_));
  INV_X1     g0288(.I(new_n673_), .ZN(new_n674_));
  NOR2_X1    g0289(.A1(new_n674_), .A2(new_n672_), .ZN(new_n675_));
  NOR3_X1    g0290(.A1(new_n675_), .A2(new_n668_), .A3(new_n670_), .ZN(new_n676_));
  INV_X1     g0291(.I(new_n676_), .ZN(new_n677_));
  AOI21_X1   g0292(.A1(new_n649_), .A2(new_n663_), .B(new_n677_), .ZN(new_n678_));
  INV_X1     g0293(.I(\priority[97] ), .ZN(new_n679_));
  INV_X1     g0294(.I(\priority[98] ), .ZN(new_n680_));
  INV_X1     g0295(.I(\req[96] ), .ZN(new_n681_));
  NAND2_X1   g0296(.A1(new_n681_), .A2(\priority[96] ), .ZN(new_n682_));
  NAND3_X1   g0297(.A1(new_n682_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n683_));
  INV_X1     g0298(.I(\priority[99] ), .ZN(new_n684_));
  NOR2_X1    g0299(.A1(new_n684_), .A2(\req[99] ), .ZN(new_n685_));
  NOR3_X1    g0300(.A1(new_n685_), .A2(\priority[100] ), .A3(\priority[101] ), .ZN(new_n686_));
  NOR2_X1    g0301(.A1(new_n680_), .A2(\req[97] ), .ZN(new_n687_));
  NOR2_X1    g0302(.A1(\req[98] ), .A2(\req[99] ), .ZN(new_n688_));
  INV_X1     g0303(.I(new_n688_), .ZN(new_n689_));
  NOR2_X1    g0304(.A1(new_n689_), .A2(new_n687_), .ZN(new_n690_));
  NAND3_X1   g0305(.A1(new_n686_), .A2(new_n690_), .A3(new_n683_), .ZN(new_n691_));
  INV_X1     g0306(.I(\priority[103] ), .ZN(new_n692_));
  INV_X1     g0307(.I(\priority[104] ), .ZN(new_n693_));
  INV_X1     g0308(.I(\req[102] ), .ZN(new_n694_));
  NAND2_X1   g0309(.A1(new_n694_), .A2(\priority[102] ), .ZN(new_n695_));
  NAND3_X1   g0310(.A1(new_n695_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n696_));
  NOR2_X1    g0311(.A1(\req[104] ), .A2(\req[105] ), .ZN(new_n697_));
  OAI21_X1   g0312(.A1(new_n693_), .A2(\req[103] ), .B(new_n697_), .ZN(new_n698_));
  INV_X1     g0313(.I(\priority[101] ), .ZN(new_n699_));
  NOR2_X1    g0314(.A1(new_n699_), .A2(\req[100] ), .ZN(new_n700_));
  NOR2_X1    g0315(.A1(\req[101] ), .A2(\req[102] ), .ZN(new_n701_));
  INV_X1     g0316(.I(new_n701_), .ZN(new_n702_));
  NOR2_X1    g0317(.A1(new_n702_), .A2(new_n700_), .ZN(new_n703_));
  NOR3_X1    g0318(.A1(new_n703_), .A2(new_n696_), .A3(new_n698_), .ZN(new_n704_));
  OAI21_X1   g0319(.A1(new_n678_), .A2(new_n691_), .B(new_n704_), .ZN(new_n705_));
  INV_X1     g0320(.I(\priority[106] ), .ZN(new_n706_));
  INV_X1     g0321(.I(\priority[107] ), .ZN(new_n707_));
  INV_X1     g0322(.I(\req[105] ), .ZN(new_n708_));
  NAND2_X1   g0323(.A1(new_n708_), .A2(\priority[105] ), .ZN(new_n709_));
  NAND3_X1   g0324(.A1(new_n709_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n710_));
  INV_X1     g0325(.I(\priority[108] ), .ZN(new_n711_));
  NOR2_X1    g0326(.A1(new_n711_), .A2(\req[108] ), .ZN(new_n712_));
  NOR3_X1    g0327(.A1(new_n712_), .A2(\priority[109] ), .A3(\priority[110] ), .ZN(new_n713_));
  NOR2_X1    g0328(.A1(new_n707_), .A2(\req[106] ), .ZN(new_n714_));
  NOR2_X1    g0329(.A1(\req[107] ), .A2(\req[108] ), .ZN(new_n715_));
  INV_X1     g0330(.I(new_n715_), .ZN(new_n716_));
  NOR2_X1    g0331(.A1(new_n716_), .A2(new_n714_), .ZN(new_n717_));
  NAND3_X1   g0332(.A1(new_n713_), .A2(new_n717_), .A3(new_n710_), .ZN(new_n718_));
  INV_X1     g0333(.I(new_n718_), .ZN(new_n719_));
  INV_X1     g0334(.I(\priority[112] ), .ZN(new_n720_));
  INV_X1     g0335(.I(\priority[113] ), .ZN(new_n721_));
  INV_X1     g0336(.I(\req[111] ), .ZN(new_n722_));
  NAND2_X1   g0337(.A1(new_n722_), .A2(\priority[111] ), .ZN(new_n723_));
  NAND3_X1   g0338(.A1(new_n723_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n724_));
  NOR2_X1    g0339(.A1(\req[113] ), .A2(\req[114] ), .ZN(new_n725_));
  OAI21_X1   g0340(.A1(new_n721_), .A2(\req[112] ), .B(new_n725_), .ZN(new_n726_));
  INV_X1     g0341(.I(\priority[110] ), .ZN(new_n727_));
  NOR2_X1    g0342(.A1(new_n727_), .A2(\req[109] ), .ZN(new_n728_));
  NOR2_X1    g0343(.A1(\req[110] ), .A2(\req[111] ), .ZN(new_n729_));
  INV_X1     g0344(.I(new_n729_), .ZN(new_n730_));
  NOR2_X1    g0345(.A1(new_n730_), .A2(new_n728_), .ZN(new_n731_));
  NOR3_X1    g0346(.A1(new_n731_), .A2(new_n724_), .A3(new_n726_), .ZN(new_n732_));
  INV_X1     g0347(.I(new_n732_), .ZN(new_n733_));
  AOI21_X1   g0348(.A1(new_n705_), .A2(new_n719_), .B(new_n733_), .ZN(new_n734_));
  INV_X1     g0349(.I(\priority[115] ), .ZN(new_n735_));
  INV_X1     g0350(.I(\priority[116] ), .ZN(new_n736_));
  INV_X1     g0351(.I(\req[114] ), .ZN(new_n737_));
  NAND2_X1   g0352(.A1(new_n737_), .A2(\priority[114] ), .ZN(new_n738_));
  NAND3_X1   g0353(.A1(new_n738_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n739_));
  INV_X1     g0354(.I(\priority[117] ), .ZN(new_n740_));
  NOR2_X1    g0355(.A1(new_n740_), .A2(\req[117] ), .ZN(new_n741_));
  NOR3_X1    g0356(.A1(new_n741_), .A2(\priority[118] ), .A3(\priority[119] ), .ZN(new_n742_));
  NOR2_X1    g0357(.A1(new_n736_), .A2(\req[115] ), .ZN(new_n743_));
  NOR2_X1    g0358(.A1(\req[116] ), .A2(\req[117] ), .ZN(new_n744_));
  INV_X1     g0359(.I(new_n744_), .ZN(new_n745_));
  NOR2_X1    g0360(.A1(new_n745_), .A2(new_n743_), .ZN(new_n746_));
  NAND3_X1   g0361(.A1(new_n742_), .A2(new_n746_), .A3(new_n739_), .ZN(new_n747_));
  INV_X1     g0362(.I(\priority[121] ), .ZN(new_n748_));
  INV_X1     g0363(.I(\priority[122] ), .ZN(new_n749_));
  INV_X1     g0364(.I(\req[120] ), .ZN(new_n750_));
  NAND2_X1   g0365(.A1(new_n750_), .A2(\priority[120] ), .ZN(new_n751_));
  NAND3_X1   g0366(.A1(new_n751_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n752_));
  NOR2_X1    g0367(.A1(\req[122] ), .A2(\req[123] ), .ZN(new_n753_));
  OAI21_X1   g0368(.A1(new_n749_), .A2(\req[121] ), .B(new_n753_), .ZN(new_n754_));
  INV_X1     g0369(.I(\priority[119] ), .ZN(new_n755_));
  NOR2_X1    g0370(.A1(new_n755_), .A2(\req[118] ), .ZN(new_n756_));
  NOR2_X1    g0371(.A1(\req[119] ), .A2(\req[120] ), .ZN(new_n757_));
  INV_X1     g0372(.I(new_n757_), .ZN(new_n758_));
  NOR2_X1    g0373(.A1(new_n758_), .A2(new_n756_), .ZN(new_n759_));
  NOR3_X1    g0374(.A1(new_n759_), .A2(new_n752_), .A3(new_n754_), .ZN(new_n760_));
  OAI21_X1   g0375(.A1(new_n734_), .A2(new_n747_), .B(new_n760_), .ZN(new_n761_));
  INV_X1     g0376(.I(\priority[124] ), .ZN(new_n762_));
  INV_X1     g0377(.I(\priority[125] ), .ZN(new_n763_));
  INV_X1     g0378(.I(\req[123] ), .ZN(new_n764_));
  NAND2_X1   g0379(.A1(new_n764_), .A2(\priority[123] ), .ZN(new_n765_));
  NAND3_X1   g0380(.A1(new_n765_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n766_));
  INV_X1     g0381(.I(\priority[126] ), .ZN(new_n767_));
  NOR2_X1    g0382(.A1(new_n767_), .A2(\req[126] ), .ZN(new_n768_));
  NOR3_X1    g0383(.A1(new_n768_), .A2(\priority[0] ), .A3(\priority[127] ), .ZN(new_n769_));
  NOR2_X1    g0384(.A1(new_n763_), .A2(\req[124] ), .ZN(new_n770_));
  NOR2_X1    g0385(.A1(\req[125] ), .A2(\req[126] ), .ZN(new_n771_));
  INV_X1     g0386(.I(new_n771_), .ZN(new_n772_));
  NOR2_X1    g0387(.A1(new_n772_), .A2(new_n770_), .ZN(new_n773_));
  NAND3_X1   g0388(.A1(new_n769_), .A2(new_n773_), .A3(new_n766_), .ZN(new_n774_));
  INV_X1     g0389(.I(new_n774_), .ZN(new_n775_));
  INV_X1     g0390(.I(\req[0] ), .ZN(new_n776_));
  INV_X1     g0391(.I(\priority[0] ), .ZN(new_n777_));
  NOR2_X1    g0392(.A1(new_n777_), .A2(\req[127] ), .ZN(new_n778_));
  NAND2_X1   g0393(.A1(new_n778_), .A2(new_n776_), .ZN(new_n779_));
  AOI21_X1   g0394(.A1(new_n761_), .A2(new_n775_), .B(new_n779_), .ZN(\grant[0] ));
  INV_X1     g0395(.I(\priority[6] ), .ZN(new_n781_));
  INV_X1     g0396(.I(\req[4] ), .ZN(new_n782_));
  NAND2_X1   g0397(.A1(new_n782_), .A2(\priority[4] ), .ZN(new_n783_));
  NAND3_X1   g0398(.A1(new_n783_), .A2(new_n387_), .A3(new_n781_), .ZN(new_n784_));
  INV_X1     g0399(.I(\priority[2] ), .ZN(new_n785_));
  NOR2_X1    g0400(.A1(new_n785_), .A2(\req[2] ), .ZN(new_n786_));
  NOR2_X1    g0401(.A1(new_n786_), .A2(\priority[3] ), .ZN(new_n787_));
  NOR2_X1    g0402(.A1(\req[6] ), .A2(\req[7] ), .ZN(new_n788_));
  OAI21_X1   g0403(.A1(new_n781_), .A2(\req[5] ), .B(new_n788_), .ZN(new_n789_));
  NOR2_X1    g0404(.A1(\req[3] ), .A2(\req[4] ), .ZN(new_n790_));
  INV_X1     g0405(.I(new_n790_), .ZN(new_n791_));
  NOR4_X1    g0406(.A1(new_n784_), .A2(new_n787_), .A3(new_n789_), .A4(new_n791_), .ZN(new_n792_));
  INV_X1     g0407(.I(\req[7] ), .ZN(new_n793_));
  NAND2_X1   g0408(.A1(new_n793_), .A2(\priority[7] ), .ZN(new_n794_));
  NAND3_X1   g0409(.A1(new_n794_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n795_));
  INV_X1     g0410(.I(\priority[10] ), .ZN(new_n796_));
  NOR2_X1    g0411(.A1(new_n796_), .A2(\req[10] ), .ZN(new_n797_));
  NOR3_X1    g0412(.A1(new_n797_), .A2(\priority[11] ), .A3(\priority[12] ), .ZN(new_n798_));
  NOR2_X1    g0413(.A1(new_n404_), .A2(\req[8] ), .ZN(new_n799_));
  NOR2_X1    g0414(.A1(\req[9] ), .A2(\req[10] ), .ZN(new_n800_));
  INV_X1     g0415(.I(new_n800_), .ZN(new_n801_));
  NOR2_X1    g0416(.A1(new_n801_), .A2(new_n799_), .ZN(new_n802_));
  NAND3_X1   g0417(.A1(new_n798_), .A2(new_n802_), .A3(new_n795_), .ZN(new_n803_));
  INV_X1     g0418(.I(\priority[15] ), .ZN(new_n804_));
  INV_X1     g0419(.I(\req[13] ), .ZN(new_n805_));
  NAND2_X1   g0420(.A1(new_n805_), .A2(\priority[13] ), .ZN(new_n806_));
  NAND3_X1   g0421(.A1(new_n806_), .A2(new_n413_), .A3(new_n804_), .ZN(new_n807_));
  NOR2_X1    g0422(.A1(\req[15] ), .A2(\req[16] ), .ZN(new_n808_));
  OAI21_X1   g0423(.A1(new_n804_), .A2(\req[14] ), .B(new_n808_), .ZN(new_n809_));
  INV_X1     g0424(.I(\priority[12] ), .ZN(new_n810_));
  NOR2_X1    g0425(.A1(new_n810_), .A2(\req[11] ), .ZN(new_n811_));
  NOR2_X1    g0426(.A1(\req[12] ), .A2(\req[13] ), .ZN(new_n812_));
  INV_X1     g0427(.I(new_n812_), .ZN(new_n813_));
  NOR2_X1    g0428(.A1(new_n813_), .A2(new_n811_), .ZN(new_n814_));
  NOR3_X1    g0429(.A1(new_n814_), .A2(new_n807_), .A3(new_n809_), .ZN(new_n815_));
  OAI21_X1   g0430(.A1(new_n803_), .A2(new_n792_), .B(new_n815_), .ZN(new_n816_));
  INV_X1     g0431(.I(\req[16] ), .ZN(new_n817_));
  NAND2_X1   g0432(.A1(new_n817_), .A2(\priority[16] ), .ZN(new_n818_));
  NAND3_X1   g0433(.A1(new_n818_), .A2(new_n427_), .A3(new_n431_), .ZN(new_n819_));
  INV_X1     g0434(.I(\priority[19] ), .ZN(new_n820_));
  NOR2_X1    g0435(.A1(new_n820_), .A2(\req[19] ), .ZN(new_n821_));
  NOR3_X1    g0436(.A1(new_n821_), .A2(\priority[20] ), .A3(\priority[21] ), .ZN(new_n822_));
  NOR2_X1    g0437(.A1(new_n431_), .A2(\req[17] ), .ZN(new_n823_));
  NOR2_X1    g0438(.A1(\req[18] ), .A2(\req[19] ), .ZN(new_n824_));
  INV_X1     g0439(.I(new_n824_), .ZN(new_n825_));
  NOR2_X1    g0440(.A1(new_n825_), .A2(new_n823_), .ZN(new_n826_));
  NAND3_X1   g0441(.A1(new_n822_), .A2(new_n826_), .A3(new_n819_), .ZN(new_n827_));
  INV_X1     g0442(.I(new_n827_), .ZN(new_n828_));
  INV_X1     g0443(.I(\priority[24] ), .ZN(new_n829_));
  INV_X1     g0444(.I(\req[22] ), .ZN(new_n830_));
  NAND2_X1   g0445(.A1(new_n830_), .A2(\priority[22] ), .ZN(new_n831_));
  NAND3_X1   g0446(.A1(new_n831_), .A2(new_n441_), .A3(new_n829_), .ZN(new_n832_));
  NOR2_X1    g0447(.A1(\req[24] ), .A2(\req[25] ), .ZN(new_n833_));
  OAI21_X1   g0448(.A1(new_n829_), .A2(\req[23] ), .B(new_n833_), .ZN(new_n834_));
  INV_X1     g0449(.I(\priority[21] ), .ZN(new_n835_));
  NOR2_X1    g0450(.A1(new_n835_), .A2(\req[20] ), .ZN(new_n836_));
  NOR2_X1    g0451(.A1(\req[21] ), .A2(\req[22] ), .ZN(new_n837_));
  INV_X1     g0452(.I(new_n837_), .ZN(new_n838_));
  NOR2_X1    g0453(.A1(new_n838_), .A2(new_n836_), .ZN(new_n839_));
  NOR3_X1    g0454(.A1(new_n839_), .A2(new_n832_), .A3(new_n834_), .ZN(new_n840_));
  INV_X1     g0455(.I(new_n840_), .ZN(new_n841_));
  AOI21_X1   g0456(.A1(new_n816_), .A2(new_n828_), .B(new_n841_), .ZN(new_n842_));
  INV_X1     g0457(.I(\req[25] ), .ZN(new_n843_));
  NAND2_X1   g0458(.A1(new_n843_), .A2(\priority[25] ), .ZN(new_n844_));
  NAND3_X1   g0459(.A1(new_n844_), .A2(new_n456_), .A3(new_n460_), .ZN(new_n845_));
  INV_X1     g0460(.I(\priority[28] ), .ZN(new_n846_));
  NOR2_X1    g0461(.A1(new_n846_), .A2(\req[28] ), .ZN(new_n847_));
  NOR3_X1    g0462(.A1(new_n847_), .A2(\priority[29] ), .A3(\priority[30] ), .ZN(new_n848_));
  NOR2_X1    g0463(.A1(new_n460_), .A2(\req[26] ), .ZN(new_n849_));
  NOR2_X1    g0464(.A1(\req[27] ), .A2(\req[28] ), .ZN(new_n850_));
  INV_X1     g0465(.I(new_n850_), .ZN(new_n851_));
  NOR2_X1    g0466(.A1(new_n851_), .A2(new_n849_), .ZN(new_n852_));
  NAND3_X1   g0467(.A1(new_n848_), .A2(new_n852_), .A3(new_n845_), .ZN(new_n853_));
  INV_X1     g0468(.I(\priority[33] ), .ZN(new_n854_));
  INV_X1     g0469(.I(\req[31] ), .ZN(new_n855_));
  NAND2_X1   g0470(.A1(new_n855_), .A2(\priority[31] ), .ZN(new_n856_));
  NAND3_X1   g0471(.A1(new_n856_), .A2(new_n469_), .A3(new_n854_), .ZN(new_n857_));
  NOR2_X1    g0472(.A1(\req[33] ), .A2(\req[34] ), .ZN(new_n858_));
  OAI21_X1   g0473(.A1(new_n854_), .A2(\req[32] ), .B(new_n858_), .ZN(new_n859_));
  INV_X1     g0474(.I(\priority[30] ), .ZN(new_n860_));
  NOR2_X1    g0475(.A1(new_n860_), .A2(\req[29] ), .ZN(new_n861_));
  NOR2_X1    g0476(.A1(\req[30] ), .A2(\req[31] ), .ZN(new_n862_));
  INV_X1     g0477(.I(new_n862_), .ZN(new_n863_));
  NOR2_X1    g0478(.A1(new_n863_), .A2(new_n861_), .ZN(new_n864_));
  NOR3_X1    g0479(.A1(new_n864_), .A2(new_n857_), .A3(new_n859_), .ZN(new_n865_));
  OAI21_X1   g0480(.A1(new_n842_), .A2(new_n853_), .B(new_n865_), .ZN(new_n866_));
  INV_X1     g0481(.I(\req[34] ), .ZN(new_n867_));
  NAND2_X1   g0482(.A1(new_n867_), .A2(\priority[34] ), .ZN(new_n868_));
  NAND3_X1   g0483(.A1(new_n868_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n869_));
  INV_X1     g0484(.I(\priority[37] ), .ZN(new_n870_));
  NOR2_X1    g0485(.A1(new_n870_), .A2(\req[37] ), .ZN(new_n871_));
  NOR3_X1    g0486(.A1(new_n871_), .A2(\priority[38] ), .A3(\priority[39] ), .ZN(new_n872_));
  NOR2_X1    g0487(.A1(new_n487_), .A2(\req[35] ), .ZN(new_n873_));
  NOR2_X1    g0488(.A1(\req[36] ), .A2(\req[37] ), .ZN(new_n874_));
  INV_X1     g0489(.I(new_n874_), .ZN(new_n875_));
  NOR2_X1    g0490(.A1(new_n875_), .A2(new_n873_), .ZN(new_n876_));
  NAND3_X1   g0491(.A1(new_n872_), .A2(new_n876_), .A3(new_n869_), .ZN(new_n877_));
  INV_X1     g0492(.I(new_n877_), .ZN(new_n878_));
  INV_X1     g0493(.I(\priority[42] ), .ZN(new_n879_));
  INV_X1     g0494(.I(\req[40] ), .ZN(new_n880_));
  NAND2_X1   g0495(.A1(new_n880_), .A2(\priority[40] ), .ZN(new_n881_));
  NAND3_X1   g0496(.A1(new_n881_), .A2(new_n497_), .A3(new_n879_), .ZN(new_n882_));
  NOR2_X1    g0497(.A1(\req[42] ), .A2(\req[43] ), .ZN(new_n883_));
  OAI21_X1   g0498(.A1(new_n879_), .A2(\req[41] ), .B(new_n883_), .ZN(new_n884_));
  INV_X1     g0499(.I(\priority[39] ), .ZN(new_n885_));
  NOR2_X1    g0500(.A1(new_n885_), .A2(\req[38] ), .ZN(new_n886_));
  NOR2_X1    g0501(.A1(\req[39] ), .A2(\req[40] ), .ZN(new_n887_));
  INV_X1     g0502(.I(new_n887_), .ZN(new_n888_));
  NOR2_X1    g0503(.A1(new_n888_), .A2(new_n886_), .ZN(new_n889_));
  NOR3_X1    g0504(.A1(new_n889_), .A2(new_n882_), .A3(new_n884_), .ZN(new_n890_));
  INV_X1     g0505(.I(new_n890_), .ZN(new_n891_));
  AOI21_X1   g0506(.A1(new_n866_), .A2(new_n878_), .B(new_n891_), .ZN(new_n892_));
  INV_X1     g0507(.I(\req[43] ), .ZN(new_n893_));
  NAND2_X1   g0508(.A1(new_n893_), .A2(\priority[43] ), .ZN(new_n894_));
  NAND3_X1   g0509(.A1(new_n894_), .A2(new_n512_), .A3(new_n516_), .ZN(new_n895_));
  INV_X1     g0510(.I(\priority[46] ), .ZN(new_n896_));
  NOR2_X1    g0511(.A1(new_n896_), .A2(\req[46] ), .ZN(new_n897_));
  NOR3_X1    g0512(.A1(new_n897_), .A2(\priority[47] ), .A3(\priority[48] ), .ZN(new_n898_));
  NOR2_X1    g0513(.A1(new_n516_), .A2(\req[44] ), .ZN(new_n899_));
  NOR2_X1    g0514(.A1(\req[45] ), .A2(\req[46] ), .ZN(new_n900_));
  INV_X1     g0515(.I(new_n900_), .ZN(new_n901_));
  NOR2_X1    g0516(.A1(new_n901_), .A2(new_n899_), .ZN(new_n902_));
  NAND3_X1   g0517(.A1(new_n898_), .A2(new_n902_), .A3(new_n895_), .ZN(new_n903_));
  INV_X1     g0518(.I(\priority[51] ), .ZN(new_n904_));
  INV_X1     g0519(.I(\req[49] ), .ZN(new_n905_));
  NAND2_X1   g0520(.A1(new_n905_), .A2(\priority[49] ), .ZN(new_n906_));
  NAND3_X1   g0521(.A1(new_n906_), .A2(new_n525_), .A3(new_n904_), .ZN(new_n907_));
  NOR2_X1    g0522(.A1(\req[51] ), .A2(\req[52] ), .ZN(new_n908_));
  OAI21_X1   g0523(.A1(new_n904_), .A2(\req[50] ), .B(new_n908_), .ZN(new_n909_));
  INV_X1     g0524(.I(\priority[48] ), .ZN(new_n910_));
  NOR2_X1    g0525(.A1(new_n910_), .A2(\req[47] ), .ZN(new_n911_));
  NOR2_X1    g0526(.A1(\req[48] ), .A2(\req[49] ), .ZN(new_n912_));
  INV_X1     g0527(.I(new_n912_), .ZN(new_n913_));
  NOR2_X1    g0528(.A1(new_n913_), .A2(new_n911_), .ZN(new_n914_));
  NOR3_X1    g0529(.A1(new_n914_), .A2(new_n907_), .A3(new_n909_), .ZN(new_n915_));
  OAI21_X1   g0530(.A1(new_n892_), .A2(new_n903_), .B(new_n915_), .ZN(new_n916_));
  INV_X1     g0531(.I(\req[52] ), .ZN(new_n917_));
  NAND2_X1   g0532(.A1(new_n917_), .A2(\priority[52] ), .ZN(new_n918_));
  NAND3_X1   g0533(.A1(new_n918_), .A2(new_n539_), .A3(new_n543_), .ZN(new_n919_));
  INV_X1     g0534(.I(\priority[55] ), .ZN(new_n920_));
  NOR2_X1    g0535(.A1(new_n920_), .A2(\req[55] ), .ZN(new_n921_));
  NOR3_X1    g0536(.A1(new_n921_), .A2(\priority[56] ), .A3(\priority[57] ), .ZN(new_n922_));
  NOR2_X1    g0537(.A1(new_n543_), .A2(\req[53] ), .ZN(new_n923_));
  NOR2_X1    g0538(.A1(\req[54] ), .A2(\req[55] ), .ZN(new_n924_));
  INV_X1     g0539(.I(new_n924_), .ZN(new_n925_));
  NOR2_X1    g0540(.A1(new_n925_), .A2(new_n923_), .ZN(new_n926_));
  NAND3_X1   g0541(.A1(new_n922_), .A2(new_n926_), .A3(new_n919_), .ZN(new_n927_));
  INV_X1     g0542(.I(new_n927_), .ZN(new_n928_));
  INV_X1     g0543(.I(\priority[60] ), .ZN(new_n929_));
  INV_X1     g0544(.I(\req[58] ), .ZN(new_n930_));
  NAND2_X1   g0545(.A1(new_n930_), .A2(\priority[58] ), .ZN(new_n931_));
  NAND3_X1   g0546(.A1(new_n931_), .A2(new_n553_), .A3(new_n929_), .ZN(new_n932_));
  NOR2_X1    g0547(.A1(\req[60] ), .A2(\req[61] ), .ZN(new_n933_));
  OAI21_X1   g0548(.A1(new_n929_), .A2(\req[59] ), .B(new_n933_), .ZN(new_n934_));
  INV_X1     g0549(.I(\priority[57] ), .ZN(new_n935_));
  NOR2_X1    g0550(.A1(new_n935_), .A2(\req[56] ), .ZN(new_n936_));
  NOR2_X1    g0551(.A1(\req[57] ), .A2(\req[58] ), .ZN(new_n937_));
  INV_X1     g0552(.I(new_n937_), .ZN(new_n938_));
  NOR2_X1    g0553(.A1(new_n938_), .A2(new_n936_), .ZN(new_n939_));
  NOR3_X1    g0554(.A1(new_n939_), .A2(new_n932_), .A3(new_n934_), .ZN(new_n940_));
  INV_X1     g0555(.I(new_n940_), .ZN(new_n941_));
  AOI21_X1   g0556(.A1(new_n916_), .A2(new_n928_), .B(new_n941_), .ZN(new_n942_));
  INV_X1     g0557(.I(\req[61] ), .ZN(new_n943_));
  NAND2_X1   g0558(.A1(new_n943_), .A2(\priority[61] ), .ZN(new_n944_));
  NAND3_X1   g0559(.A1(new_n944_), .A2(new_n568_), .A3(new_n572_), .ZN(new_n945_));
  INV_X1     g0560(.I(\priority[64] ), .ZN(new_n946_));
  NOR2_X1    g0561(.A1(new_n946_), .A2(\req[64] ), .ZN(new_n947_));
  NOR3_X1    g0562(.A1(new_n947_), .A2(\priority[65] ), .A3(\priority[66] ), .ZN(new_n948_));
  NOR2_X1    g0563(.A1(new_n572_), .A2(\req[62] ), .ZN(new_n949_));
  NOR2_X1    g0564(.A1(\req[63] ), .A2(\req[64] ), .ZN(new_n950_));
  INV_X1     g0565(.I(new_n950_), .ZN(new_n951_));
  NOR2_X1    g0566(.A1(new_n951_), .A2(new_n949_), .ZN(new_n952_));
  NAND3_X1   g0567(.A1(new_n948_), .A2(new_n952_), .A3(new_n945_), .ZN(new_n953_));
  INV_X1     g0568(.I(\priority[69] ), .ZN(new_n954_));
  INV_X1     g0569(.I(\req[67] ), .ZN(new_n955_));
  NAND2_X1   g0570(.A1(new_n955_), .A2(\priority[67] ), .ZN(new_n956_));
  NAND3_X1   g0571(.A1(new_n956_), .A2(new_n581_), .A3(new_n954_), .ZN(new_n957_));
  NOR2_X1    g0572(.A1(\req[69] ), .A2(\req[70] ), .ZN(new_n958_));
  OAI21_X1   g0573(.A1(new_n954_), .A2(\req[68] ), .B(new_n958_), .ZN(new_n959_));
  INV_X1     g0574(.I(\priority[66] ), .ZN(new_n960_));
  NOR2_X1    g0575(.A1(new_n960_), .A2(\req[65] ), .ZN(new_n961_));
  NOR2_X1    g0576(.A1(\req[66] ), .A2(\req[67] ), .ZN(new_n962_));
  INV_X1     g0577(.I(new_n962_), .ZN(new_n963_));
  NOR2_X1    g0578(.A1(new_n963_), .A2(new_n961_), .ZN(new_n964_));
  NOR3_X1    g0579(.A1(new_n964_), .A2(new_n957_), .A3(new_n959_), .ZN(new_n965_));
  OAI21_X1   g0580(.A1(new_n942_), .A2(new_n953_), .B(new_n965_), .ZN(new_n966_));
  INV_X1     g0581(.I(\req[70] ), .ZN(new_n967_));
  NAND2_X1   g0582(.A1(new_n967_), .A2(\priority[70] ), .ZN(new_n968_));
  NAND3_X1   g0583(.A1(new_n968_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n969_));
  INV_X1     g0584(.I(\priority[73] ), .ZN(new_n970_));
  NOR2_X1    g0585(.A1(new_n970_), .A2(\req[73] ), .ZN(new_n971_));
  NOR3_X1    g0586(.A1(new_n971_), .A2(\priority[74] ), .A3(\priority[75] ), .ZN(new_n972_));
  NOR2_X1    g0587(.A1(new_n599_), .A2(\req[71] ), .ZN(new_n973_));
  NOR2_X1    g0588(.A1(\req[72] ), .A2(\req[73] ), .ZN(new_n974_));
  INV_X1     g0589(.I(new_n974_), .ZN(new_n975_));
  NOR2_X1    g0590(.A1(new_n975_), .A2(new_n973_), .ZN(new_n976_));
  NAND3_X1   g0591(.A1(new_n972_), .A2(new_n976_), .A3(new_n969_), .ZN(new_n977_));
  INV_X1     g0592(.I(new_n977_), .ZN(new_n978_));
  INV_X1     g0593(.I(\priority[78] ), .ZN(new_n979_));
  INV_X1     g0594(.I(\req[76] ), .ZN(new_n980_));
  NAND2_X1   g0595(.A1(new_n980_), .A2(\priority[76] ), .ZN(new_n981_));
  NAND3_X1   g0596(.A1(new_n981_), .A2(new_n609_), .A3(new_n979_), .ZN(new_n982_));
  NOR2_X1    g0597(.A1(\req[78] ), .A2(\req[79] ), .ZN(new_n983_));
  OAI21_X1   g0598(.A1(new_n979_), .A2(\req[77] ), .B(new_n983_), .ZN(new_n984_));
  INV_X1     g0599(.I(\priority[75] ), .ZN(new_n985_));
  NOR2_X1    g0600(.A1(new_n985_), .A2(\req[74] ), .ZN(new_n986_));
  NOR2_X1    g0601(.A1(\req[75] ), .A2(\req[76] ), .ZN(new_n987_));
  INV_X1     g0602(.I(new_n987_), .ZN(new_n988_));
  NOR2_X1    g0603(.A1(new_n988_), .A2(new_n986_), .ZN(new_n989_));
  NOR3_X1    g0604(.A1(new_n989_), .A2(new_n982_), .A3(new_n984_), .ZN(new_n990_));
  INV_X1     g0605(.I(new_n990_), .ZN(new_n991_));
  AOI21_X1   g0606(.A1(new_n966_), .A2(new_n978_), .B(new_n991_), .ZN(new_n992_));
  INV_X1     g0607(.I(\req[79] ), .ZN(new_n993_));
  NAND2_X1   g0608(.A1(new_n993_), .A2(\priority[79] ), .ZN(new_n994_));
  NAND3_X1   g0609(.A1(new_n994_), .A2(new_n624_), .A3(new_n628_), .ZN(new_n995_));
  INV_X1     g0610(.I(\priority[82] ), .ZN(new_n996_));
  NOR2_X1    g0611(.A1(new_n996_), .A2(\req[82] ), .ZN(new_n997_));
  NOR3_X1    g0612(.A1(new_n997_), .A2(\priority[83] ), .A3(\priority[84] ), .ZN(new_n998_));
  NOR2_X1    g0613(.A1(new_n628_), .A2(\req[80] ), .ZN(new_n999_));
  NOR2_X1    g0614(.A1(\req[81] ), .A2(\req[82] ), .ZN(new_n1000_));
  INV_X1     g0615(.I(new_n1000_), .ZN(new_n1001_));
  NOR2_X1    g0616(.A1(new_n1001_), .A2(new_n999_), .ZN(new_n1002_));
  NAND3_X1   g0617(.A1(new_n998_), .A2(new_n1002_), .A3(new_n995_), .ZN(new_n1003_));
  INV_X1     g0618(.I(\priority[87] ), .ZN(new_n1004_));
  INV_X1     g0619(.I(\req[85] ), .ZN(new_n1005_));
  NAND2_X1   g0620(.A1(new_n1005_), .A2(\priority[85] ), .ZN(new_n1006_));
  NAND3_X1   g0621(.A1(new_n1006_), .A2(new_n637_), .A3(new_n1004_), .ZN(new_n1007_));
  NOR2_X1    g0622(.A1(\req[87] ), .A2(\req[88] ), .ZN(new_n1008_));
  OAI21_X1   g0623(.A1(new_n1004_), .A2(\req[86] ), .B(new_n1008_), .ZN(new_n1009_));
  INV_X1     g0624(.I(\priority[84] ), .ZN(new_n1010_));
  NOR2_X1    g0625(.A1(new_n1010_), .A2(\req[83] ), .ZN(new_n1011_));
  NOR2_X1    g0626(.A1(\req[84] ), .A2(\req[85] ), .ZN(new_n1012_));
  INV_X1     g0627(.I(new_n1012_), .ZN(new_n1013_));
  NOR2_X1    g0628(.A1(new_n1013_), .A2(new_n1011_), .ZN(new_n1014_));
  NOR3_X1    g0629(.A1(new_n1014_), .A2(new_n1007_), .A3(new_n1009_), .ZN(new_n1015_));
  OAI21_X1   g0630(.A1(new_n992_), .A2(new_n1003_), .B(new_n1015_), .ZN(new_n1016_));
  INV_X1     g0631(.I(\req[88] ), .ZN(new_n1017_));
  NAND2_X1   g0632(.A1(new_n1017_), .A2(\priority[88] ), .ZN(new_n1018_));
  NAND3_X1   g0633(.A1(new_n1018_), .A2(new_n651_), .A3(new_n655_), .ZN(new_n1019_));
  INV_X1     g0634(.I(\priority[91] ), .ZN(new_n1020_));
  NOR2_X1    g0635(.A1(new_n1020_), .A2(\req[91] ), .ZN(new_n1021_));
  NOR3_X1    g0636(.A1(new_n1021_), .A2(\priority[92] ), .A3(\priority[93] ), .ZN(new_n1022_));
  NOR2_X1    g0637(.A1(new_n655_), .A2(\req[89] ), .ZN(new_n1023_));
  NOR2_X1    g0638(.A1(\req[90] ), .A2(\req[91] ), .ZN(new_n1024_));
  INV_X1     g0639(.I(new_n1024_), .ZN(new_n1025_));
  NOR2_X1    g0640(.A1(new_n1025_), .A2(new_n1023_), .ZN(new_n1026_));
  NAND3_X1   g0641(.A1(new_n1022_), .A2(new_n1026_), .A3(new_n1019_), .ZN(new_n1027_));
  INV_X1     g0642(.I(new_n1027_), .ZN(new_n1028_));
  INV_X1     g0643(.I(\priority[96] ), .ZN(new_n1029_));
  INV_X1     g0644(.I(\req[94] ), .ZN(new_n1030_));
  NAND2_X1   g0645(.A1(new_n1030_), .A2(\priority[94] ), .ZN(new_n1031_));
  NAND3_X1   g0646(.A1(new_n1031_), .A2(new_n665_), .A3(new_n1029_), .ZN(new_n1032_));
  NOR2_X1    g0647(.A1(\req[96] ), .A2(\req[97] ), .ZN(new_n1033_));
  OAI21_X1   g0648(.A1(new_n1029_), .A2(\req[95] ), .B(new_n1033_), .ZN(new_n1034_));
  INV_X1     g0649(.I(\priority[93] ), .ZN(new_n1035_));
  NOR2_X1    g0650(.A1(new_n1035_), .A2(\req[92] ), .ZN(new_n1036_));
  NOR2_X1    g0651(.A1(\req[93] ), .A2(\req[94] ), .ZN(new_n1037_));
  INV_X1     g0652(.I(new_n1037_), .ZN(new_n1038_));
  NOR2_X1    g0653(.A1(new_n1038_), .A2(new_n1036_), .ZN(new_n1039_));
  NOR3_X1    g0654(.A1(new_n1039_), .A2(new_n1032_), .A3(new_n1034_), .ZN(new_n1040_));
  INV_X1     g0655(.I(new_n1040_), .ZN(new_n1041_));
  AOI21_X1   g0656(.A1(new_n1016_), .A2(new_n1028_), .B(new_n1041_), .ZN(new_n1042_));
  INV_X1     g0657(.I(\req[97] ), .ZN(new_n1043_));
  NAND2_X1   g0658(.A1(new_n1043_), .A2(\priority[97] ), .ZN(new_n1044_));
  NAND3_X1   g0659(.A1(new_n1044_), .A2(new_n680_), .A3(new_n684_), .ZN(new_n1045_));
  INV_X1     g0660(.I(\priority[100] ), .ZN(new_n1046_));
  NOR2_X1    g0661(.A1(new_n1046_), .A2(\req[100] ), .ZN(new_n1047_));
  NOR3_X1    g0662(.A1(new_n1047_), .A2(\priority[101] ), .A3(\priority[102] ), .ZN(new_n1048_));
  NOR2_X1    g0663(.A1(new_n684_), .A2(\req[98] ), .ZN(new_n1049_));
  NOR2_X1    g0664(.A1(\req[99] ), .A2(\req[100] ), .ZN(new_n1050_));
  INV_X1     g0665(.I(new_n1050_), .ZN(new_n1051_));
  NOR2_X1    g0666(.A1(new_n1051_), .A2(new_n1049_), .ZN(new_n1052_));
  NAND3_X1   g0667(.A1(new_n1048_), .A2(new_n1052_), .A3(new_n1045_), .ZN(new_n1053_));
  INV_X1     g0668(.I(\priority[105] ), .ZN(new_n1054_));
  INV_X1     g0669(.I(\req[103] ), .ZN(new_n1055_));
  NAND2_X1   g0670(.A1(new_n1055_), .A2(\priority[103] ), .ZN(new_n1056_));
  NAND3_X1   g0671(.A1(new_n1056_), .A2(new_n693_), .A3(new_n1054_), .ZN(new_n1057_));
  NOR2_X1    g0672(.A1(\req[105] ), .A2(\req[106] ), .ZN(new_n1058_));
  OAI21_X1   g0673(.A1(new_n1054_), .A2(\req[104] ), .B(new_n1058_), .ZN(new_n1059_));
  INV_X1     g0674(.I(\priority[102] ), .ZN(new_n1060_));
  NOR2_X1    g0675(.A1(new_n1060_), .A2(\req[101] ), .ZN(new_n1061_));
  NOR2_X1    g0676(.A1(\req[102] ), .A2(\req[103] ), .ZN(new_n1062_));
  INV_X1     g0677(.I(new_n1062_), .ZN(new_n1063_));
  NOR2_X1    g0678(.A1(new_n1063_), .A2(new_n1061_), .ZN(new_n1064_));
  NOR3_X1    g0679(.A1(new_n1064_), .A2(new_n1057_), .A3(new_n1059_), .ZN(new_n1065_));
  OAI21_X1   g0680(.A1(new_n1042_), .A2(new_n1053_), .B(new_n1065_), .ZN(new_n1066_));
  INV_X1     g0681(.I(\req[106] ), .ZN(new_n1067_));
  NAND2_X1   g0682(.A1(new_n1067_), .A2(\priority[106] ), .ZN(new_n1068_));
  NAND3_X1   g0683(.A1(new_n1068_), .A2(new_n707_), .A3(new_n711_), .ZN(new_n1069_));
  INV_X1     g0684(.I(\priority[109] ), .ZN(new_n1070_));
  NOR2_X1    g0685(.A1(new_n1070_), .A2(\req[109] ), .ZN(new_n1071_));
  NOR3_X1    g0686(.A1(new_n1071_), .A2(\priority[110] ), .A3(\priority[111] ), .ZN(new_n1072_));
  NOR2_X1    g0687(.A1(new_n711_), .A2(\req[107] ), .ZN(new_n1073_));
  NOR2_X1    g0688(.A1(\req[108] ), .A2(\req[109] ), .ZN(new_n1074_));
  INV_X1     g0689(.I(new_n1074_), .ZN(new_n1075_));
  NOR2_X1    g0690(.A1(new_n1075_), .A2(new_n1073_), .ZN(new_n1076_));
  NAND3_X1   g0691(.A1(new_n1072_), .A2(new_n1076_), .A3(new_n1069_), .ZN(new_n1077_));
  INV_X1     g0692(.I(new_n1077_), .ZN(new_n1078_));
  INV_X1     g0693(.I(\priority[114] ), .ZN(new_n1079_));
  INV_X1     g0694(.I(\req[112] ), .ZN(new_n1080_));
  NAND2_X1   g0695(.A1(new_n1080_), .A2(\priority[112] ), .ZN(new_n1081_));
  NAND3_X1   g0696(.A1(new_n1081_), .A2(new_n721_), .A3(new_n1079_), .ZN(new_n1082_));
  NOR2_X1    g0697(.A1(\req[114] ), .A2(\req[115] ), .ZN(new_n1083_));
  OAI21_X1   g0698(.A1(new_n1079_), .A2(\req[113] ), .B(new_n1083_), .ZN(new_n1084_));
  INV_X1     g0699(.I(\priority[111] ), .ZN(new_n1085_));
  NOR2_X1    g0700(.A1(new_n1085_), .A2(\req[110] ), .ZN(new_n1086_));
  NOR2_X1    g0701(.A1(\req[111] ), .A2(\req[112] ), .ZN(new_n1087_));
  INV_X1     g0702(.I(new_n1087_), .ZN(new_n1088_));
  NOR2_X1    g0703(.A1(new_n1088_), .A2(new_n1086_), .ZN(new_n1089_));
  NOR3_X1    g0704(.A1(new_n1089_), .A2(new_n1082_), .A3(new_n1084_), .ZN(new_n1090_));
  INV_X1     g0705(.I(new_n1090_), .ZN(new_n1091_));
  AOI21_X1   g0706(.A1(new_n1066_), .A2(new_n1078_), .B(new_n1091_), .ZN(new_n1092_));
  INV_X1     g0707(.I(\req[115] ), .ZN(new_n1093_));
  NAND2_X1   g0708(.A1(new_n1093_), .A2(\priority[115] ), .ZN(new_n1094_));
  NAND3_X1   g0709(.A1(new_n1094_), .A2(new_n736_), .A3(new_n740_), .ZN(new_n1095_));
  INV_X1     g0710(.I(\priority[118] ), .ZN(new_n1096_));
  NOR2_X1    g0711(.A1(new_n1096_), .A2(\req[118] ), .ZN(new_n1097_));
  NOR3_X1    g0712(.A1(new_n1097_), .A2(\priority[119] ), .A3(\priority[120] ), .ZN(new_n1098_));
  NOR2_X1    g0713(.A1(new_n740_), .A2(\req[116] ), .ZN(new_n1099_));
  NOR2_X1    g0714(.A1(\req[117] ), .A2(\req[118] ), .ZN(new_n1100_));
  INV_X1     g0715(.I(new_n1100_), .ZN(new_n1101_));
  NOR2_X1    g0716(.A1(new_n1101_), .A2(new_n1099_), .ZN(new_n1102_));
  NAND3_X1   g0717(.A1(new_n1098_), .A2(new_n1102_), .A3(new_n1095_), .ZN(new_n1103_));
  INV_X1     g0718(.I(\priority[123] ), .ZN(new_n1104_));
  INV_X1     g0719(.I(\req[121] ), .ZN(new_n1105_));
  NAND2_X1   g0720(.A1(new_n1105_), .A2(\priority[121] ), .ZN(new_n1106_));
  NAND3_X1   g0721(.A1(new_n1106_), .A2(new_n749_), .A3(new_n1104_), .ZN(new_n1107_));
  NOR2_X1    g0722(.A1(\req[123] ), .A2(\req[124] ), .ZN(new_n1108_));
  OAI21_X1   g0723(.A1(new_n1104_), .A2(\req[122] ), .B(new_n1108_), .ZN(new_n1109_));
  INV_X1     g0724(.I(\priority[120] ), .ZN(new_n1110_));
  NOR2_X1    g0725(.A1(new_n1110_), .A2(\req[119] ), .ZN(new_n1111_));
  NOR2_X1    g0726(.A1(\req[120] ), .A2(\req[121] ), .ZN(new_n1112_));
  INV_X1     g0727(.I(new_n1112_), .ZN(new_n1113_));
  NOR2_X1    g0728(.A1(new_n1113_), .A2(new_n1111_), .ZN(new_n1114_));
  NOR3_X1    g0729(.A1(new_n1114_), .A2(new_n1107_), .A3(new_n1109_), .ZN(new_n1115_));
  OAI21_X1   g0730(.A1(new_n1092_), .A2(new_n1103_), .B(new_n1115_), .ZN(new_n1116_));
  INV_X1     g0731(.I(\req[124] ), .ZN(new_n1117_));
  NAND2_X1   g0732(.A1(new_n1117_), .A2(\priority[124] ), .ZN(new_n1118_));
  NAND3_X1   g0733(.A1(new_n1118_), .A2(new_n763_), .A3(new_n767_), .ZN(new_n1119_));
  INV_X1     g0734(.I(\priority[127] ), .ZN(new_n1120_));
  NOR2_X1    g0735(.A1(new_n1120_), .A2(\req[127] ), .ZN(new_n1121_));
  NOR3_X1    g0736(.A1(new_n1121_), .A2(\priority[0] ), .A3(\priority[1] ), .ZN(new_n1122_));
  NOR2_X1    g0737(.A1(new_n767_), .A2(\req[125] ), .ZN(new_n1123_));
  NOR2_X1    g0738(.A1(\req[126] ), .A2(\req[127] ), .ZN(new_n1124_));
  INV_X1     g0739(.I(new_n1124_), .ZN(new_n1125_));
  NOR2_X1    g0740(.A1(new_n1125_), .A2(new_n1123_), .ZN(new_n1126_));
  NAND3_X1   g0741(.A1(new_n1122_), .A2(new_n1126_), .A3(new_n1119_), .ZN(new_n1127_));
  INV_X1     g0742(.I(new_n1127_), .ZN(new_n1128_));
  INV_X1     g0743(.I(\req[1] ), .ZN(new_n1129_));
  NOR2_X1    g0744(.A1(new_n391_), .A2(\req[0] ), .ZN(new_n1130_));
  NAND2_X1   g0745(.A1(new_n1130_), .A2(new_n1129_), .ZN(new_n1131_));
  AOI21_X1   g0746(.A1(new_n1116_), .A2(new_n1128_), .B(new_n1131_), .ZN(\grant[1] ));
  INV_X1     g0747(.I(\req[5] ), .ZN(new_n1133_));
  NAND2_X1   g0748(.A1(new_n1133_), .A2(\priority[5] ), .ZN(new_n1134_));
  NAND3_X1   g0749(.A1(new_n1134_), .A2(new_n781_), .A3(new_n399_), .ZN(new_n1135_));
  NOR2_X1    g0750(.A1(\req[7] ), .A2(\req[8] ), .ZN(new_n1136_));
  OAI21_X1   g0751(.A1(new_n399_), .A2(\req[6] ), .B(new_n1136_), .ZN(new_n1137_));
  INV_X1     g0752(.I(\priority[3] ), .ZN(new_n1138_));
  NOR2_X1    g0753(.A1(new_n1138_), .A2(\req[3] ), .ZN(new_n1139_));
  NOR2_X1    g0754(.A1(\req[4] ), .A2(\req[5] ), .ZN(new_n1140_));
  OAI21_X1   g0755(.A1(new_n1139_), .A2(\priority[4] ), .B(new_n1140_), .ZN(new_n1141_));
  NOR3_X1    g0756(.A1(new_n1141_), .A2(new_n1135_), .A3(new_n1137_), .ZN(new_n1142_));
  INV_X1     g0757(.I(\req[8] ), .ZN(new_n1143_));
  NAND2_X1   g0758(.A1(new_n1143_), .A2(\priority[8] ), .ZN(new_n1144_));
  NAND3_X1   g0759(.A1(new_n1144_), .A2(new_n404_), .A3(new_n796_), .ZN(new_n1145_));
  NOR2_X1    g0760(.A1(new_n419_), .A2(\req[11] ), .ZN(new_n1146_));
  NOR3_X1    g0761(.A1(new_n1146_), .A2(\priority[12] ), .A3(\priority[13] ), .ZN(new_n1147_));
  NOR2_X1    g0762(.A1(new_n796_), .A2(\req[9] ), .ZN(new_n1148_));
  NOR3_X1    g0763(.A1(new_n1148_), .A2(\req[10] ), .A3(\req[11] ), .ZN(new_n1149_));
  NAND3_X1   g0764(.A1(new_n1147_), .A2(new_n1149_), .A3(new_n1145_), .ZN(new_n1150_));
  INV_X1     g0765(.I(\req[14] ), .ZN(new_n1151_));
  NAND2_X1   g0766(.A1(new_n1151_), .A2(\priority[14] ), .ZN(new_n1152_));
  NAND3_X1   g0767(.A1(new_n1152_), .A2(new_n804_), .A3(new_n426_), .ZN(new_n1153_));
  NOR2_X1    g0768(.A1(\req[16] ), .A2(\req[17] ), .ZN(new_n1154_));
  OAI21_X1   g0769(.A1(new_n426_), .A2(\req[15] ), .B(new_n1154_), .ZN(new_n1155_));
  NOR2_X1    g0770(.A1(new_n412_), .A2(\req[12] ), .ZN(new_n1156_));
  NOR3_X1    g0771(.A1(new_n1156_), .A2(\req[13] ), .A3(\req[14] ), .ZN(new_n1157_));
  NOR3_X1    g0772(.A1(new_n1157_), .A2(new_n1153_), .A3(new_n1155_), .ZN(new_n1158_));
  OAI21_X1   g0773(.A1(new_n1150_), .A2(new_n1142_), .B(new_n1158_), .ZN(new_n1159_));
  INV_X1     g0774(.I(\req[17] ), .ZN(new_n1160_));
  NAND2_X1   g0775(.A1(new_n1160_), .A2(\priority[17] ), .ZN(new_n1161_));
  NAND3_X1   g0776(.A1(new_n1161_), .A2(new_n431_), .A3(new_n820_), .ZN(new_n1162_));
  NOR2_X1    g0777(.A1(new_n447_), .A2(\req[20] ), .ZN(new_n1163_));
  NOR3_X1    g0778(.A1(new_n1163_), .A2(\priority[21] ), .A3(\priority[22] ), .ZN(new_n1164_));
  NOR2_X1    g0779(.A1(new_n820_), .A2(\req[18] ), .ZN(new_n1165_));
  NOR3_X1    g0780(.A1(new_n1165_), .A2(\req[19] ), .A3(\req[20] ), .ZN(new_n1166_));
  NAND3_X1   g0781(.A1(new_n1164_), .A2(new_n1166_), .A3(new_n1162_), .ZN(new_n1167_));
  INV_X1     g0782(.I(new_n1167_), .ZN(new_n1168_));
  INV_X1     g0783(.I(\req[23] ), .ZN(new_n1169_));
  NAND2_X1   g0784(.A1(new_n1169_), .A2(\priority[23] ), .ZN(new_n1170_));
  NAND3_X1   g0785(.A1(new_n1170_), .A2(new_n829_), .A3(new_n455_), .ZN(new_n1171_));
  NOR2_X1    g0786(.A1(\req[25] ), .A2(\req[26] ), .ZN(new_n1172_));
  OAI21_X1   g0787(.A1(new_n455_), .A2(\req[24] ), .B(new_n1172_), .ZN(new_n1173_));
  NOR2_X1    g0788(.A1(new_n440_), .A2(\req[21] ), .ZN(new_n1174_));
  NOR3_X1    g0789(.A1(new_n1174_), .A2(\req[22] ), .A3(\req[23] ), .ZN(new_n1175_));
  NOR3_X1    g0790(.A1(new_n1175_), .A2(new_n1171_), .A3(new_n1173_), .ZN(new_n1176_));
  INV_X1     g0791(.I(new_n1176_), .ZN(new_n1177_));
  AOI21_X1   g0792(.A1(new_n1159_), .A2(new_n1168_), .B(new_n1177_), .ZN(new_n1178_));
  INV_X1     g0793(.I(\req[26] ), .ZN(new_n1179_));
  NAND2_X1   g0794(.A1(new_n1179_), .A2(\priority[26] ), .ZN(new_n1180_));
  NAND3_X1   g0795(.A1(new_n1180_), .A2(new_n460_), .A3(new_n846_), .ZN(new_n1181_));
  NOR2_X1    g0796(.A1(new_n475_), .A2(\req[29] ), .ZN(new_n1182_));
  NOR3_X1    g0797(.A1(new_n1182_), .A2(\priority[30] ), .A3(\priority[31] ), .ZN(new_n1183_));
  NOR2_X1    g0798(.A1(new_n846_), .A2(\req[27] ), .ZN(new_n1184_));
  NOR3_X1    g0799(.A1(new_n1184_), .A2(\req[28] ), .A3(\req[29] ), .ZN(new_n1185_));
  NAND3_X1   g0800(.A1(new_n1183_), .A2(new_n1185_), .A3(new_n1181_), .ZN(new_n1186_));
  INV_X1     g0801(.I(\req[32] ), .ZN(new_n1187_));
  NAND2_X1   g0802(.A1(new_n1187_), .A2(\priority[32] ), .ZN(new_n1188_));
  NAND3_X1   g0803(.A1(new_n1188_), .A2(new_n854_), .A3(new_n482_), .ZN(new_n1189_));
  NOR2_X1    g0804(.A1(\req[34] ), .A2(\req[35] ), .ZN(new_n1190_));
  OAI21_X1   g0805(.A1(new_n482_), .A2(\req[33] ), .B(new_n1190_), .ZN(new_n1191_));
  NOR2_X1    g0806(.A1(new_n468_), .A2(\req[30] ), .ZN(new_n1192_));
  NOR3_X1    g0807(.A1(new_n1192_), .A2(\req[31] ), .A3(\req[32] ), .ZN(new_n1193_));
  NOR3_X1    g0808(.A1(new_n1193_), .A2(new_n1189_), .A3(new_n1191_), .ZN(new_n1194_));
  OAI21_X1   g0809(.A1(new_n1178_), .A2(new_n1186_), .B(new_n1194_), .ZN(new_n1195_));
  INV_X1     g0810(.I(\req[35] ), .ZN(new_n1196_));
  NAND2_X1   g0811(.A1(new_n1196_), .A2(\priority[35] ), .ZN(new_n1197_));
  NAND3_X1   g0812(.A1(new_n1197_), .A2(new_n487_), .A3(new_n870_), .ZN(new_n1198_));
  NOR2_X1    g0813(.A1(new_n503_), .A2(\req[38] ), .ZN(new_n1199_));
  NOR3_X1    g0814(.A1(new_n1199_), .A2(\priority[39] ), .A3(\priority[40] ), .ZN(new_n1200_));
  NOR2_X1    g0815(.A1(new_n870_), .A2(\req[36] ), .ZN(new_n1201_));
  NOR3_X1    g0816(.A1(new_n1201_), .A2(\req[37] ), .A3(\req[38] ), .ZN(new_n1202_));
  NAND3_X1   g0817(.A1(new_n1200_), .A2(new_n1202_), .A3(new_n1198_), .ZN(new_n1203_));
  INV_X1     g0818(.I(new_n1203_), .ZN(new_n1204_));
  INV_X1     g0819(.I(\req[41] ), .ZN(new_n1205_));
  NAND2_X1   g0820(.A1(new_n1205_), .A2(\priority[41] ), .ZN(new_n1206_));
  NAND3_X1   g0821(.A1(new_n1206_), .A2(new_n879_), .A3(new_n511_), .ZN(new_n1207_));
  NOR2_X1    g0822(.A1(\req[43] ), .A2(\req[44] ), .ZN(new_n1208_));
  OAI21_X1   g0823(.A1(new_n511_), .A2(\req[42] ), .B(new_n1208_), .ZN(new_n1209_));
  NOR2_X1    g0824(.A1(new_n496_), .A2(\req[39] ), .ZN(new_n1210_));
  NOR3_X1    g0825(.A1(new_n1210_), .A2(\req[40] ), .A3(\req[41] ), .ZN(new_n1211_));
  NOR3_X1    g0826(.A1(new_n1211_), .A2(new_n1207_), .A3(new_n1209_), .ZN(new_n1212_));
  INV_X1     g0827(.I(new_n1212_), .ZN(new_n1213_));
  AOI21_X1   g0828(.A1(new_n1195_), .A2(new_n1204_), .B(new_n1213_), .ZN(new_n1214_));
  INV_X1     g0829(.I(\req[44] ), .ZN(new_n1215_));
  NAND2_X1   g0830(.A1(new_n1215_), .A2(\priority[44] ), .ZN(new_n1216_));
  NAND3_X1   g0831(.A1(new_n1216_), .A2(new_n516_), .A3(new_n896_), .ZN(new_n1217_));
  NOR2_X1    g0832(.A1(new_n531_), .A2(\req[47] ), .ZN(new_n1218_));
  NOR3_X1    g0833(.A1(new_n1218_), .A2(\priority[48] ), .A3(\priority[49] ), .ZN(new_n1219_));
  NOR2_X1    g0834(.A1(new_n896_), .A2(\req[45] ), .ZN(new_n1220_));
  NOR3_X1    g0835(.A1(new_n1220_), .A2(\req[46] ), .A3(\req[47] ), .ZN(new_n1221_));
  NAND3_X1   g0836(.A1(new_n1219_), .A2(new_n1221_), .A3(new_n1217_), .ZN(new_n1222_));
  INV_X1     g0837(.I(\req[50] ), .ZN(new_n1223_));
  NAND2_X1   g0838(.A1(new_n1223_), .A2(\priority[50] ), .ZN(new_n1224_));
  NAND3_X1   g0839(.A1(new_n1224_), .A2(new_n904_), .A3(new_n538_), .ZN(new_n1225_));
  NOR2_X1    g0840(.A1(\req[52] ), .A2(\req[53] ), .ZN(new_n1226_));
  OAI21_X1   g0841(.A1(new_n538_), .A2(\req[51] ), .B(new_n1226_), .ZN(new_n1227_));
  NOR2_X1    g0842(.A1(new_n524_), .A2(\req[48] ), .ZN(new_n1228_));
  NOR3_X1    g0843(.A1(new_n1228_), .A2(\req[49] ), .A3(\req[50] ), .ZN(new_n1229_));
  NOR3_X1    g0844(.A1(new_n1229_), .A2(new_n1225_), .A3(new_n1227_), .ZN(new_n1230_));
  OAI21_X1   g0845(.A1(new_n1214_), .A2(new_n1222_), .B(new_n1230_), .ZN(new_n1231_));
  INV_X1     g0846(.I(\req[53] ), .ZN(new_n1232_));
  NAND2_X1   g0847(.A1(new_n1232_), .A2(\priority[53] ), .ZN(new_n1233_));
  NAND3_X1   g0848(.A1(new_n1233_), .A2(new_n543_), .A3(new_n920_), .ZN(new_n1234_));
  NOR2_X1    g0849(.A1(new_n559_), .A2(\req[56] ), .ZN(new_n1235_));
  NOR3_X1    g0850(.A1(new_n1235_), .A2(\priority[57] ), .A3(\priority[58] ), .ZN(new_n1236_));
  NOR2_X1    g0851(.A1(new_n920_), .A2(\req[54] ), .ZN(new_n1237_));
  NOR3_X1    g0852(.A1(new_n1237_), .A2(\req[55] ), .A3(\req[56] ), .ZN(new_n1238_));
  NAND3_X1   g0853(.A1(new_n1236_), .A2(new_n1238_), .A3(new_n1234_), .ZN(new_n1239_));
  INV_X1     g0854(.I(new_n1239_), .ZN(new_n1240_));
  INV_X1     g0855(.I(\req[59] ), .ZN(new_n1241_));
  NAND2_X1   g0856(.A1(new_n1241_), .A2(\priority[59] ), .ZN(new_n1242_));
  NAND3_X1   g0857(.A1(new_n1242_), .A2(new_n929_), .A3(new_n567_), .ZN(new_n1243_));
  NOR2_X1    g0858(.A1(\req[61] ), .A2(\req[62] ), .ZN(new_n1244_));
  OAI21_X1   g0859(.A1(new_n567_), .A2(\req[60] ), .B(new_n1244_), .ZN(new_n1245_));
  NOR2_X1    g0860(.A1(new_n552_), .A2(\req[57] ), .ZN(new_n1246_));
  NOR3_X1    g0861(.A1(new_n1246_), .A2(\req[58] ), .A3(\req[59] ), .ZN(new_n1247_));
  NOR3_X1    g0862(.A1(new_n1247_), .A2(new_n1243_), .A3(new_n1245_), .ZN(new_n1248_));
  INV_X1     g0863(.I(new_n1248_), .ZN(new_n1249_));
  AOI21_X1   g0864(.A1(new_n1231_), .A2(new_n1240_), .B(new_n1249_), .ZN(new_n1250_));
  INV_X1     g0865(.I(\req[62] ), .ZN(new_n1251_));
  NAND2_X1   g0866(.A1(new_n1251_), .A2(\priority[62] ), .ZN(new_n1252_));
  NAND3_X1   g0867(.A1(new_n1252_), .A2(new_n572_), .A3(new_n946_), .ZN(new_n1253_));
  NOR2_X1    g0868(.A1(new_n587_), .A2(\req[65] ), .ZN(new_n1254_));
  NOR3_X1    g0869(.A1(new_n1254_), .A2(\priority[66] ), .A3(\priority[67] ), .ZN(new_n1255_));
  NOR2_X1    g0870(.A1(new_n946_), .A2(\req[63] ), .ZN(new_n1256_));
  NOR3_X1    g0871(.A1(new_n1256_), .A2(\req[64] ), .A3(\req[65] ), .ZN(new_n1257_));
  NAND3_X1   g0872(.A1(new_n1255_), .A2(new_n1257_), .A3(new_n1253_), .ZN(new_n1258_));
  INV_X1     g0873(.I(\req[68] ), .ZN(new_n1259_));
  NAND2_X1   g0874(.A1(new_n1259_), .A2(\priority[68] ), .ZN(new_n1260_));
  NAND3_X1   g0875(.A1(new_n1260_), .A2(new_n954_), .A3(new_n594_), .ZN(new_n1261_));
  NOR2_X1    g0876(.A1(\req[70] ), .A2(\req[71] ), .ZN(new_n1262_));
  OAI21_X1   g0877(.A1(new_n594_), .A2(\req[69] ), .B(new_n1262_), .ZN(new_n1263_));
  NOR2_X1    g0878(.A1(new_n580_), .A2(\req[66] ), .ZN(new_n1264_));
  NOR3_X1    g0879(.A1(new_n1264_), .A2(\req[67] ), .A3(\req[68] ), .ZN(new_n1265_));
  NOR3_X1    g0880(.A1(new_n1265_), .A2(new_n1261_), .A3(new_n1263_), .ZN(new_n1266_));
  OAI21_X1   g0881(.A1(new_n1250_), .A2(new_n1258_), .B(new_n1266_), .ZN(new_n1267_));
  INV_X1     g0882(.I(\req[71] ), .ZN(new_n1268_));
  NAND2_X1   g0883(.A1(new_n1268_), .A2(\priority[71] ), .ZN(new_n1269_));
  NAND3_X1   g0884(.A1(new_n1269_), .A2(new_n599_), .A3(new_n970_), .ZN(new_n1270_));
  NOR2_X1    g0885(.A1(new_n615_), .A2(\req[74] ), .ZN(new_n1271_));
  NOR3_X1    g0886(.A1(new_n1271_), .A2(\priority[75] ), .A3(\priority[76] ), .ZN(new_n1272_));
  NOR2_X1    g0887(.A1(new_n970_), .A2(\req[72] ), .ZN(new_n1273_));
  NOR3_X1    g0888(.A1(new_n1273_), .A2(\req[73] ), .A3(\req[74] ), .ZN(new_n1274_));
  NAND3_X1   g0889(.A1(new_n1272_), .A2(new_n1274_), .A3(new_n1270_), .ZN(new_n1275_));
  INV_X1     g0890(.I(new_n1275_), .ZN(new_n1276_));
  INV_X1     g0891(.I(\req[77] ), .ZN(new_n1277_));
  NAND2_X1   g0892(.A1(new_n1277_), .A2(\priority[77] ), .ZN(new_n1278_));
  NAND3_X1   g0893(.A1(new_n1278_), .A2(new_n979_), .A3(new_n623_), .ZN(new_n1279_));
  NOR2_X1    g0894(.A1(\req[79] ), .A2(\req[80] ), .ZN(new_n1280_));
  OAI21_X1   g0895(.A1(new_n623_), .A2(\req[78] ), .B(new_n1280_), .ZN(new_n1281_));
  NOR2_X1    g0896(.A1(new_n608_), .A2(\req[75] ), .ZN(new_n1282_));
  NOR3_X1    g0897(.A1(new_n1282_), .A2(\req[76] ), .A3(\req[77] ), .ZN(new_n1283_));
  NOR3_X1    g0898(.A1(new_n1283_), .A2(new_n1279_), .A3(new_n1281_), .ZN(new_n1284_));
  INV_X1     g0899(.I(new_n1284_), .ZN(new_n1285_));
  AOI21_X1   g0900(.A1(new_n1267_), .A2(new_n1276_), .B(new_n1285_), .ZN(new_n1286_));
  INV_X1     g0901(.I(\req[80] ), .ZN(new_n1287_));
  NAND2_X1   g0902(.A1(new_n1287_), .A2(\priority[80] ), .ZN(new_n1288_));
  NAND3_X1   g0903(.A1(new_n1288_), .A2(new_n628_), .A3(new_n996_), .ZN(new_n1289_));
  NOR2_X1    g0904(.A1(new_n643_), .A2(\req[83] ), .ZN(new_n1290_));
  NOR3_X1    g0905(.A1(new_n1290_), .A2(\priority[84] ), .A3(\priority[85] ), .ZN(new_n1291_));
  NOR2_X1    g0906(.A1(new_n996_), .A2(\req[81] ), .ZN(new_n1292_));
  NOR3_X1    g0907(.A1(new_n1292_), .A2(\req[82] ), .A3(\req[83] ), .ZN(new_n1293_));
  NAND3_X1   g0908(.A1(new_n1291_), .A2(new_n1293_), .A3(new_n1289_), .ZN(new_n1294_));
  INV_X1     g0909(.I(\req[86] ), .ZN(new_n1295_));
  NAND2_X1   g0910(.A1(new_n1295_), .A2(\priority[86] ), .ZN(new_n1296_));
  NAND3_X1   g0911(.A1(new_n1296_), .A2(new_n1004_), .A3(new_n650_), .ZN(new_n1297_));
  NOR2_X1    g0912(.A1(\req[88] ), .A2(\req[89] ), .ZN(new_n1298_));
  OAI21_X1   g0913(.A1(new_n650_), .A2(\req[87] ), .B(new_n1298_), .ZN(new_n1299_));
  NOR2_X1    g0914(.A1(new_n636_), .A2(\req[84] ), .ZN(new_n1300_));
  NOR3_X1    g0915(.A1(new_n1300_), .A2(\req[85] ), .A3(\req[86] ), .ZN(new_n1301_));
  NOR3_X1    g0916(.A1(new_n1301_), .A2(new_n1297_), .A3(new_n1299_), .ZN(new_n1302_));
  OAI21_X1   g0917(.A1(new_n1286_), .A2(new_n1294_), .B(new_n1302_), .ZN(new_n1303_));
  INV_X1     g0918(.I(\req[89] ), .ZN(new_n1304_));
  NAND2_X1   g0919(.A1(new_n1304_), .A2(\priority[89] ), .ZN(new_n1305_));
  NAND3_X1   g0920(.A1(new_n1305_), .A2(new_n655_), .A3(new_n1020_), .ZN(new_n1306_));
  NOR2_X1    g0921(.A1(new_n671_), .A2(\req[92] ), .ZN(new_n1307_));
  NOR3_X1    g0922(.A1(new_n1307_), .A2(\priority[93] ), .A3(\priority[94] ), .ZN(new_n1308_));
  NOR2_X1    g0923(.A1(new_n1020_), .A2(\req[90] ), .ZN(new_n1309_));
  NOR3_X1    g0924(.A1(new_n1309_), .A2(\req[91] ), .A3(\req[92] ), .ZN(new_n1310_));
  NAND3_X1   g0925(.A1(new_n1308_), .A2(new_n1310_), .A3(new_n1306_), .ZN(new_n1311_));
  INV_X1     g0926(.I(new_n1311_), .ZN(new_n1312_));
  INV_X1     g0927(.I(\req[95] ), .ZN(new_n1313_));
  NAND2_X1   g0928(.A1(new_n1313_), .A2(\priority[95] ), .ZN(new_n1314_));
  NAND3_X1   g0929(.A1(new_n1314_), .A2(new_n1029_), .A3(new_n679_), .ZN(new_n1315_));
  NOR2_X1    g0930(.A1(\req[97] ), .A2(\req[98] ), .ZN(new_n1316_));
  OAI21_X1   g0931(.A1(new_n679_), .A2(\req[96] ), .B(new_n1316_), .ZN(new_n1317_));
  NOR2_X1    g0932(.A1(new_n664_), .A2(\req[93] ), .ZN(new_n1318_));
  NOR3_X1    g0933(.A1(new_n1318_), .A2(\req[94] ), .A3(\req[95] ), .ZN(new_n1319_));
  NOR3_X1    g0934(.A1(new_n1319_), .A2(new_n1315_), .A3(new_n1317_), .ZN(new_n1320_));
  INV_X1     g0935(.I(new_n1320_), .ZN(new_n1321_));
  AOI21_X1   g0936(.A1(new_n1303_), .A2(new_n1312_), .B(new_n1321_), .ZN(new_n1322_));
  INV_X1     g0937(.I(\req[98] ), .ZN(new_n1323_));
  NAND2_X1   g0938(.A1(new_n1323_), .A2(\priority[98] ), .ZN(new_n1324_));
  NAND3_X1   g0939(.A1(new_n1324_), .A2(new_n684_), .A3(new_n1046_), .ZN(new_n1325_));
  NOR2_X1    g0940(.A1(new_n699_), .A2(\req[101] ), .ZN(new_n1326_));
  NOR3_X1    g0941(.A1(new_n1326_), .A2(\priority[102] ), .A3(\priority[103] ), .ZN(new_n1327_));
  NOR2_X1    g0942(.A1(new_n1046_), .A2(\req[99] ), .ZN(new_n1328_));
  NOR3_X1    g0943(.A1(new_n1328_), .A2(\req[100] ), .A3(\req[101] ), .ZN(new_n1329_));
  NAND3_X1   g0944(.A1(new_n1327_), .A2(new_n1329_), .A3(new_n1325_), .ZN(new_n1330_));
  INV_X1     g0945(.I(\req[104] ), .ZN(new_n1331_));
  NAND2_X1   g0946(.A1(new_n1331_), .A2(\priority[104] ), .ZN(new_n1332_));
  NAND3_X1   g0947(.A1(new_n1332_), .A2(new_n1054_), .A3(new_n706_), .ZN(new_n1333_));
  NOR2_X1    g0948(.A1(\req[106] ), .A2(\req[107] ), .ZN(new_n1334_));
  OAI21_X1   g0949(.A1(new_n706_), .A2(\req[105] ), .B(new_n1334_), .ZN(new_n1335_));
  NOR2_X1    g0950(.A1(new_n692_), .A2(\req[102] ), .ZN(new_n1336_));
  NOR3_X1    g0951(.A1(new_n1336_), .A2(\req[103] ), .A3(\req[104] ), .ZN(new_n1337_));
  NOR3_X1    g0952(.A1(new_n1337_), .A2(new_n1333_), .A3(new_n1335_), .ZN(new_n1338_));
  OAI21_X1   g0953(.A1(new_n1322_), .A2(new_n1330_), .B(new_n1338_), .ZN(new_n1339_));
  INV_X1     g0954(.I(\req[107] ), .ZN(new_n1340_));
  NAND2_X1   g0955(.A1(new_n1340_), .A2(\priority[107] ), .ZN(new_n1341_));
  NAND3_X1   g0956(.A1(new_n1341_), .A2(new_n711_), .A3(new_n1070_), .ZN(new_n1342_));
  NOR2_X1    g0957(.A1(new_n727_), .A2(\req[110] ), .ZN(new_n1343_));
  NOR3_X1    g0958(.A1(new_n1343_), .A2(\priority[111] ), .A3(\priority[112] ), .ZN(new_n1344_));
  NOR2_X1    g0959(.A1(new_n1070_), .A2(\req[108] ), .ZN(new_n1345_));
  NOR3_X1    g0960(.A1(new_n1345_), .A2(\req[109] ), .A3(\req[110] ), .ZN(new_n1346_));
  NAND3_X1   g0961(.A1(new_n1344_), .A2(new_n1346_), .A3(new_n1342_), .ZN(new_n1347_));
  INV_X1     g0962(.I(new_n1347_), .ZN(new_n1348_));
  INV_X1     g0963(.I(\req[113] ), .ZN(new_n1349_));
  NAND2_X1   g0964(.A1(new_n1349_), .A2(\priority[113] ), .ZN(new_n1350_));
  NAND3_X1   g0965(.A1(new_n1350_), .A2(new_n1079_), .A3(new_n735_), .ZN(new_n1351_));
  NOR2_X1    g0966(.A1(\req[115] ), .A2(\req[116] ), .ZN(new_n1352_));
  OAI21_X1   g0967(.A1(new_n735_), .A2(\req[114] ), .B(new_n1352_), .ZN(new_n1353_));
  NOR2_X1    g0968(.A1(new_n720_), .A2(\req[111] ), .ZN(new_n1354_));
  NOR3_X1    g0969(.A1(new_n1354_), .A2(\req[112] ), .A3(\req[113] ), .ZN(new_n1355_));
  NOR3_X1    g0970(.A1(new_n1355_), .A2(new_n1351_), .A3(new_n1353_), .ZN(new_n1356_));
  INV_X1     g0971(.I(new_n1356_), .ZN(new_n1357_));
  AOI21_X1   g0972(.A1(new_n1339_), .A2(new_n1348_), .B(new_n1357_), .ZN(new_n1358_));
  INV_X1     g0973(.I(\req[116] ), .ZN(new_n1359_));
  NAND2_X1   g0974(.A1(new_n1359_), .A2(\priority[116] ), .ZN(new_n1360_));
  NAND3_X1   g0975(.A1(new_n1360_), .A2(new_n740_), .A3(new_n1096_), .ZN(new_n1361_));
  NOR2_X1    g0976(.A1(new_n755_), .A2(\req[119] ), .ZN(new_n1362_));
  NOR3_X1    g0977(.A1(new_n1362_), .A2(\priority[120] ), .A3(\priority[121] ), .ZN(new_n1363_));
  NOR2_X1    g0978(.A1(new_n1096_), .A2(\req[117] ), .ZN(new_n1364_));
  NOR3_X1    g0979(.A1(new_n1364_), .A2(\req[118] ), .A3(\req[119] ), .ZN(new_n1365_));
  NAND3_X1   g0980(.A1(new_n1363_), .A2(new_n1365_), .A3(new_n1361_), .ZN(new_n1366_));
  INV_X1     g0981(.I(\req[122] ), .ZN(new_n1367_));
  NAND2_X1   g0982(.A1(new_n1367_), .A2(\priority[122] ), .ZN(new_n1368_));
  NAND3_X1   g0983(.A1(new_n1368_), .A2(new_n1104_), .A3(new_n762_), .ZN(new_n1369_));
  NOR2_X1    g0984(.A1(\req[124] ), .A2(\req[125] ), .ZN(new_n1370_));
  OAI21_X1   g0985(.A1(new_n762_), .A2(\req[123] ), .B(new_n1370_), .ZN(new_n1371_));
  NOR2_X1    g0986(.A1(new_n748_), .A2(\req[120] ), .ZN(new_n1372_));
  NOR3_X1    g0987(.A1(new_n1372_), .A2(\req[121] ), .A3(\req[122] ), .ZN(new_n1373_));
  NOR3_X1    g0988(.A1(new_n1373_), .A2(new_n1369_), .A3(new_n1371_), .ZN(new_n1374_));
  OAI21_X1   g0989(.A1(new_n1358_), .A2(new_n1366_), .B(new_n1374_), .ZN(new_n1375_));
  INV_X1     g0990(.I(\req[125] ), .ZN(new_n1376_));
  NAND2_X1   g0991(.A1(new_n1376_), .A2(\priority[125] ), .ZN(new_n1377_));
  NAND3_X1   g0992(.A1(new_n1377_), .A2(new_n767_), .A3(new_n1120_), .ZN(new_n1378_));
  NOR2_X1    g0993(.A1(new_n777_), .A2(\req[0] ), .ZN(new_n1379_));
  NOR3_X1    g0994(.A1(new_n1379_), .A2(\priority[1] ), .A3(\priority[2] ), .ZN(new_n1380_));
  NOR2_X1    g0995(.A1(new_n1120_), .A2(\req[126] ), .ZN(new_n1381_));
  NOR2_X1    g0996(.A1(\req[0] ), .A2(\req[127] ), .ZN(new_n1382_));
  INV_X1     g0997(.I(new_n1382_), .ZN(new_n1383_));
  NOR2_X1    g0998(.A1(new_n1383_), .A2(new_n1381_), .ZN(new_n1384_));
  NAND3_X1   g0999(.A1(new_n1380_), .A2(new_n1384_), .A3(new_n1378_), .ZN(new_n1385_));
  INV_X1     g1000(.I(new_n1385_), .ZN(new_n1386_));
  INV_X1     g1001(.I(\req[2] ), .ZN(new_n1387_));
  NOR2_X1    g1002(.A1(new_n785_), .A2(\req[1] ), .ZN(new_n1388_));
  NAND2_X1   g1003(.A1(new_n1388_), .A2(new_n1387_), .ZN(new_n1389_));
  AOI21_X1   g1004(.A1(new_n1375_), .A2(new_n1386_), .B(new_n1389_), .ZN(\grant[2] ));
  INV_X1     g1005(.I(new_n394_), .ZN(new_n1391_));
  OAI21_X1   g1006(.A1(new_n400_), .A2(\req[7] ), .B(new_n408_), .ZN(new_n1392_));
  AOI21_X1   g1007(.A1(new_n782_), .A2(\priority[4] ), .B(\priority[5] ), .ZN(new_n1393_));
  NOR4_X1    g1008(.A1(new_n403_), .A2(new_n1391_), .A3(new_n1392_), .A4(new_n1393_), .ZN(new_n1394_));
  INV_X1     g1009(.I(\req[9] ), .ZN(new_n1395_));
  NAND2_X1   g1010(.A1(new_n1395_), .A2(\priority[9] ), .ZN(new_n1396_));
  NAND3_X1   g1011(.A1(new_n1396_), .A2(new_n796_), .A3(new_n419_), .ZN(new_n1397_));
  NOR2_X1    g1012(.A1(new_n810_), .A2(\req[12] ), .ZN(new_n1398_));
  NOR3_X1    g1013(.A1(new_n1398_), .A2(\priority[13] ), .A3(\priority[14] ), .ZN(new_n1399_));
  NAND3_X1   g1014(.A1(new_n1399_), .A2(new_n423_), .A3(new_n1397_), .ZN(new_n1400_));
  NOR2_X1    g1015(.A1(new_n413_), .A2(\req[13] ), .ZN(new_n1401_));
  INV_X1     g1016(.I(new_n417_), .ZN(new_n1402_));
  NOR2_X1    g1017(.A1(new_n1402_), .A2(new_n1401_), .ZN(new_n1403_));
  OAI21_X1   g1018(.A1(new_n427_), .A2(\req[16] ), .B(new_n435_), .ZN(new_n1404_));
  NOR3_X1    g1019(.A1(new_n1403_), .A2(new_n430_), .A3(new_n1404_), .ZN(new_n1405_));
  OAI21_X1   g1020(.A1(new_n1400_), .A2(new_n1394_), .B(new_n1405_), .ZN(new_n1406_));
  INV_X1     g1021(.I(\req[18] ), .ZN(new_n1407_));
  NAND2_X1   g1022(.A1(new_n1407_), .A2(\priority[18] ), .ZN(new_n1408_));
  NAND3_X1   g1023(.A1(new_n1408_), .A2(new_n820_), .A3(new_n447_), .ZN(new_n1409_));
  NOR2_X1    g1024(.A1(new_n835_), .A2(\req[21] ), .ZN(new_n1410_));
  NOR3_X1    g1025(.A1(new_n1410_), .A2(\priority[22] ), .A3(\priority[23] ), .ZN(new_n1411_));
  NAND3_X1   g1026(.A1(new_n1411_), .A2(new_n451_), .A3(new_n1409_), .ZN(new_n1412_));
  INV_X1     g1027(.I(new_n1412_), .ZN(new_n1413_));
  NOR2_X1    g1028(.A1(new_n441_), .A2(\req[22] ), .ZN(new_n1414_));
  INV_X1     g1029(.I(new_n445_), .ZN(new_n1415_));
  NOR2_X1    g1030(.A1(new_n1415_), .A2(new_n1414_), .ZN(new_n1416_));
  OAI21_X1   g1031(.A1(new_n456_), .A2(\req[25] ), .B(new_n464_), .ZN(new_n1417_));
  NOR3_X1    g1032(.A1(new_n1416_), .A2(new_n459_), .A3(new_n1417_), .ZN(new_n1418_));
  INV_X1     g1033(.I(new_n1418_), .ZN(new_n1419_));
  AOI21_X1   g1034(.A1(new_n1406_), .A2(new_n1413_), .B(new_n1419_), .ZN(new_n1420_));
  INV_X1     g1035(.I(\req[27] ), .ZN(new_n1421_));
  NAND2_X1   g1036(.A1(new_n1421_), .A2(\priority[27] ), .ZN(new_n1422_));
  NAND3_X1   g1037(.A1(new_n1422_), .A2(new_n846_), .A3(new_n475_), .ZN(new_n1423_));
  NOR2_X1    g1038(.A1(new_n860_), .A2(\req[30] ), .ZN(new_n1424_));
  NOR3_X1    g1039(.A1(new_n1424_), .A2(\priority[31] ), .A3(\priority[32] ), .ZN(new_n1425_));
  NAND3_X1   g1040(.A1(new_n1425_), .A2(new_n479_), .A3(new_n1423_), .ZN(new_n1426_));
  NOR2_X1    g1041(.A1(new_n469_), .A2(\req[31] ), .ZN(new_n1427_));
  INV_X1     g1042(.I(new_n473_), .ZN(new_n1428_));
  NOR2_X1    g1043(.A1(new_n1428_), .A2(new_n1427_), .ZN(new_n1429_));
  OAI21_X1   g1044(.A1(new_n483_), .A2(\req[34] ), .B(new_n491_), .ZN(new_n1430_));
  NOR3_X1    g1045(.A1(new_n1429_), .A2(new_n486_), .A3(new_n1430_), .ZN(new_n1431_));
  OAI21_X1   g1046(.A1(new_n1420_), .A2(new_n1426_), .B(new_n1431_), .ZN(new_n1432_));
  INV_X1     g1047(.I(\req[36] ), .ZN(new_n1433_));
  NAND2_X1   g1048(.A1(new_n1433_), .A2(\priority[36] ), .ZN(new_n1434_));
  NAND3_X1   g1049(.A1(new_n1434_), .A2(new_n870_), .A3(new_n503_), .ZN(new_n1435_));
  NOR2_X1    g1050(.A1(new_n885_), .A2(\req[39] ), .ZN(new_n1436_));
  NOR3_X1    g1051(.A1(new_n1436_), .A2(\priority[40] ), .A3(\priority[41] ), .ZN(new_n1437_));
  NAND3_X1   g1052(.A1(new_n1437_), .A2(new_n507_), .A3(new_n1435_), .ZN(new_n1438_));
  INV_X1     g1053(.I(new_n1438_), .ZN(new_n1439_));
  NOR2_X1    g1054(.A1(new_n497_), .A2(\req[40] ), .ZN(new_n1440_));
  INV_X1     g1055(.I(new_n501_), .ZN(new_n1441_));
  NOR2_X1    g1056(.A1(new_n1441_), .A2(new_n1440_), .ZN(new_n1442_));
  OAI21_X1   g1057(.A1(new_n512_), .A2(\req[43] ), .B(new_n520_), .ZN(new_n1443_));
  NOR3_X1    g1058(.A1(new_n1442_), .A2(new_n515_), .A3(new_n1443_), .ZN(new_n1444_));
  INV_X1     g1059(.I(new_n1444_), .ZN(new_n1445_));
  AOI21_X1   g1060(.A1(new_n1432_), .A2(new_n1439_), .B(new_n1445_), .ZN(new_n1446_));
  INV_X1     g1061(.I(\req[45] ), .ZN(new_n1447_));
  NAND2_X1   g1062(.A1(new_n1447_), .A2(\priority[45] ), .ZN(new_n1448_));
  NAND3_X1   g1063(.A1(new_n1448_), .A2(new_n896_), .A3(new_n531_), .ZN(new_n1449_));
  NOR2_X1    g1064(.A1(new_n910_), .A2(\req[48] ), .ZN(new_n1450_));
  NOR3_X1    g1065(.A1(new_n1450_), .A2(\priority[49] ), .A3(\priority[50] ), .ZN(new_n1451_));
  NAND3_X1   g1066(.A1(new_n1451_), .A2(new_n535_), .A3(new_n1449_), .ZN(new_n1452_));
  NOR2_X1    g1067(.A1(new_n525_), .A2(\req[49] ), .ZN(new_n1453_));
  INV_X1     g1068(.I(new_n529_), .ZN(new_n1454_));
  NOR2_X1    g1069(.A1(new_n1454_), .A2(new_n1453_), .ZN(new_n1455_));
  OAI21_X1   g1070(.A1(new_n539_), .A2(\req[52] ), .B(new_n547_), .ZN(new_n1456_));
  NOR3_X1    g1071(.A1(new_n1455_), .A2(new_n542_), .A3(new_n1456_), .ZN(new_n1457_));
  OAI21_X1   g1072(.A1(new_n1446_), .A2(new_n1452_), .B(new_n1457_), .ZN(new_n1458_));
  INV_X1     g1073(.I(\req[54] ), .ZN(new_n1459_));
  NAND2_X1   g1074(.A1(new_n1459_), .A2(\priority[54] ), .ZN(new_n1460_));
  NAND3_X1   g1075(.A1(new_n1460_), .A2(new_n920_), .A3(new_n559_), .ZN(new_n1461_));
  NOR2_X1    g1076(.A1(new_n935_), .A2(\req[57] ), .ZN(new_n1462_));
  NOR3_X1    g1077(.A1(new_n1462_), .A2(\priority[58] ), .A3(\priority[59] ), .ZN(new_n1463_));
  NAND3_X1   g1078(.A1(new_n1463_), .A2(new_n563_), .A3(new_n1461_), .ZN(new_n1464_));
  INV_X1     g1079(.I(new_n1464_), .ZN(new_n1465_));
  NOR2_X1    g1080(.A1(new_n553_), .A2(\req[58] ), .ZN(new_n1466_));
  INV_X1     g1081(.I(new_n557_), .ZN(new_n1467_));
  NOR2_X1    g1082(.A1(new_n1467_), .A2(new_n1466_), .ZN(new_n1468_));
  OAI21_X1   g1083(.A1(new_n568_), .A2(\req[61] ), .B(new_n576_), .ZN(new_n1469_));
  NOR3_X1    g1084(.A1(new_n1468_), .A2(new_n571_), .A3(new_n1469_), .ZN(new_n1470_));
  INV_X1     g1085(.I(new_n1470_), .ZN(new_n1471_));
  AOI21_X1   g1086(.A1(new_n1458_), .A2(new_n1465_), .B(new_n1471_), .ZN(new_n1472_));
  INV_X1     g1087(.I(\req[63] ), .ZN(new_n1473_));
  NAND2_X1   g1088(.A1(new_n1473_), .A2(\priority[63] ), .ZN(new_n1474_));
  NAND3_X1   g1089(.A1(new_n1474_), .A2(new_n946_), .A3(new_n587_), .ZN(new_n1475_));
  NOR2_X1    g1090(.A1(new_n960_), .A2(\req[66] ), .ZN(new_n1476_));
  NOR3_X1    g1091(.A1(new_n1476_), .A2(\priority[67] ), .A3(\priority[68] ), .ZN(new_n1477_));
  NAND3_X1   g1092(.A1(new_n1477_), .A2(new_n591_), .A3(new_n1475_), .ZN(new_n1478_));
  NOR2_X1    g1093(.A1(new_n581_), .A2(\req[67] ), .ZN(new_n1479_));
  INV_X1     g1094(.I(new_n585_), .ZN(new_n1480_));
  NOR2_X1    g1095(.A1(new_n1480_), .A2(new_n1479_), .ZN(new_n1481_));
  OAI21_X1   g1096(.A1(new_n595_), .A2(\req[70] ), .B(new_n603_), .ZN(new_n1482_));
  NOR3_X1    g1097(.A1(new_n1481_), .A2(new_n598_), .A3(new_n1482_), .ZN(new_n1483_));
  OAI21_X1   g1098(.A1(new_n1472_), .A2(new_n1478_), .B(new_n1483_), .ZN(new_n1484_));
  INV_X1     g1099(.I(\req[72] ), .ZN(new_n1485_));
  NAND2_X1   g1100(.A1(new_n1485_), .A2(\priority[72] ), .ZN(new_n1486_));
  NAND3_X1   g1101(.A1(new_n1486_), .A2(new_n970_), .A3(new_n615_), .ZN(new_n1487_));
  NOR2_X1    g1102(.A1(new_n985_), .A2(\req[75] ), .ZN(new_n1488_));
  NOR3_X1    g1103(.A1(new_n1488_), .A2(\priority[76] ), .A3(\priority[77] ), .ZN(new_n1489_));
  NAND3_X1   g1104(.A1(new_n1489_), .A2(new_n619_), .A3(new_n1487_), .ZN(new_n1490_));
  INV_X1     g1105(.I(new_n1490_), .ZN(new_n1491_));
  NOR2_X1    g1106(.A1(new_n609_), .A2(\req[76] ), .ZN(new_n1492_));
  INV_X1     g1107(.I(new_n613_), .ZN(new_n1493_));
  NOR2_X1    g1108(.A1(new_n1493_), .A2(new_n1492_), .ZN(new_n1494_));
  OAI21_X1   g1109(.A1(new_n624_), .A2(\req[79] ), .B(new_n632_), .ZN(new_n1495_));
  NOR3_X1    g1110(.A1(new_n1494_), .A2(new_n627_), .A3(new_n1495_), .ZN(new_n1496_));
  INV_X1     g1111(.I(new_n1496_), .ZN(new_n1497_));
  AOI21_X1   g1112(.A1(new_n1484_), .A2(new_n1491_), .B(new_n1497_), .ZN(new_n1498_));
  INV_X1     g1113(.I(\req[81] ), .ZN(new_n1499_));
  NAND2_X1   g1114(.A1(new_n1499_), .A2(\priority[81] ), .ZN(new_n1500_));
  NAND3_X1   g1115(.A1(new_n1500_), .A2(new_n996_), .A3(new_n643_), .ZN(new_n1501_));
  NOR2_X1    g1116(.A1(new_n1010_), .A2(\req[84] ), .ZN(new_n1502_));
  NOR3_X1    g1117(.A1(new_n1502_), .A2(\priority[85] ), .A3(\priority[86] ), .ZN(new_n1503_));
  NAND3_X1   g1118(.A1(new_n1503_), .A2(new_n647_), .A3(new_n1501_), .ZN(new_n1504_));
  NOR2_X1    g1119(.A1(new_n637_), .A2(\req[85] ), .ZN(new_n1505_));
  INV_X1     g1120(.I(new_n641_), .ZN(new_n1506_));
  NOR2_X1    g1121(.A1(new_n1506_), .A2(new_n1505_), .ZN(new_n1507_));
  OAI21_X1   g1122(.A1(new_n651_), .A2(\req[88] ), .B(new_n659_), .ZN(new_n1508_));
  NOR3_X1    g1123(.A1(new_n1507_), .A2(new_n654_), .A3(new_n1508_), .ZN(new_n1509_));
  OAI21_X1   g1124(.A1(new_n1498_), .A2(new_n1504_), .B(new_n1509_), .ZN(new_n1510_));
  INV_X1     g1125(.I(\req[90] ), .ZN(new_n1511_));
  NAND2_X1   g1126(.A1(new_n1511_), .A2(\priority[90] ), .ZN(new_n1512_));
  NAND3_X1   g1127(.A1(new_n1512_), .A2(new_n1020_), .A3(new_n671_), .ZN(new_n1513_));
  NOR2_X1    g1128(.A1(new_n1035_), .A2(\req[93] ), .ZN(new_n1514_));
  NOR3_X1    g1129(.A1(new_n1514_), .A2(\priority[94] ), .A3(\priority[95] ), .ZN(new_n1515_));
  NAND3_X1   g1130(.A1(new_n1515_), .A2(new_n675_), .A3(new_n1513_), .ZN(new_n1516_));
  INV_X1     g1131(.I(new_n1516_), .ZN(new_n1517_));
  NOR2_X1    g1132(.A1(new_n665_), .A2(\req[94] ), .ZN(new_n1518_));
  INV_X1     g1133(.I(new_n669_), .ZN(new_n1519_));
  NOR2_X1    g1134(.A1(new_n1519_), .A2(new_n1518_), .ZN(new_n1520_));
  OAI21_X1   g1135(.A1(new_n680_), .A2(\req[97] ), .B(new_n688_), .ZN(new_n1521_));
  NOR3_X1    g1136(.A1(new_n1520_), .A2(new_n683_), .A3(new_n1521_), .ZN(new_n1522_));
  INV_X1     g1137(.I(new_n1522_), .ZN(new_n1523_));
  AOI21_X1   g1138(.A1(new_n1510_), .A2(new_n1517_), .B(new_n1523_), .ZN(new_n1524_));
  INV_X1     g1139(.I(\req[99] ), .ZN(new_n1525_));
  NAND2_X1   g1140(.A1(new_n1525_), .A2(\priority[99] ), .ZN(new_n1526_));
  NAND3_X1   g1141(.A1(new_n1526_), .A2(new_n1046_), .A3(new_n699_), .ZN(new_n1527_));
  NOR2_X1    g1142(.A1(new_n1060_), .A2(\req[102] ), .ZN(new_n1528_));
  NOR3_X1    g1143(.A1(new_n1528_), .A2(\priority[103] ), .A3(\priority[104] ), .ZN(new_n1529_));
  NAND3_X1   g1144(.A1(new_n1529_), .A2(new_n703_), .A3(new_n1527_), .ZN(new_n1530_));
  NOR2_X1    g1145(.A1(new_n693_), .A2(\req[103] ), .ZN(new_n1531_));
  INV_X1     g1146(.I(new_n697_), .ZN(new_n1532_));
  NOR2_X1    g1147(.A1(new_n1532_), .A2(new_n1531_), .ZN(new_n1533_));
  OAI21_X1   g1148(.A1(new_n707_), .A2(\req[106] ), .B(new_n715_), .ZN(new_n1534_));
  NOR3_X1    g1149(.A1(new_n1533_), .A2(new_n710_), .A3(new_n1534_), .ZN(new_n1535_));
  OAI21_X1   g1150(.A1(new_n1524_), .A2(new_n1530_), .B(new_n1535_), .ZN(new_n1536_));
  INV_X1     g1151(.I(\req[108] ), .ZN(new_n1537_));
  NAND2_X1   g1152(.A1(new_n1537_), .A2(\priority[108] ), .ZN(new_n1538_));
  NAND3_X1   g1153(.A1(new_n1538_), .A2(new_n1070_), .A3(new_n727_), .ZN(new_n1539_));
  NOR2_X1    g1154(.A1(new_n1085_), .A2(\req[111] ), .ZN(new_n1540_));
  NOR3_X1    g1155(.A1(new_n1540_), .A2(\priority[112] ), .A3(\priority[113] ), .ZN(new_n1541_));
  NAND3_X1   g1156(.A1(new_n1541_), .A2(new_n731_), .A3(new_n1539_), .ZN(new_n1542_));
  INV_X1     g1157(.I(new_n1542_), .ZN(new_n1543_));
  NOR2_X1    g1158(.A1(new_n721_), .A2(\req[112] ), .ZN(new_n1544_));
  INV_X1     g1159(.I(new_n725_), .ZN(new_n1545_));
  NOR2_X1    g1160(.A1(new_n1545_), .A2(new_n1544_), .ZN(new_n1546_));
  OAI21_X1   g1161(.A1(new_n736_), .A2(\req[115] ), .B(new_n744_), .ZN(new_n1547_));
  NOR3_X1    g1162(.A1(new_n1546_), .A2(new_n739_), .A3(new_n1547_), .ZN(new_n1548_));
  INV_X1     g1163(.I(new_n1548_), .ZN(new_n1549_));
  AOI21_X1   g1164(.A1(new_n1536_), .A2(new_n1543_), .B(new_n1549_), .ZN(new_n1550_));
  INV_X1     g1165(.I(\req[117] ), .ZN(new_n1551_));
  NAND2_X1   g1166(.A1(new_n1551_), .A2(\priority[117] ), .ZN(new_n1552_));
  NAND3_X1   g1167(.A1(new_n1552_), .A2(new_n1096_), .A3(new_n755_), .ZN(new_n1553_));
  NOR2_X1    g1168(.A1(new_n1110_), .A2(\req[120] ), .ZN(new_n1554_));
  NOR3_X1    g1169(.A1(new_n1554_), .A2(\priority[121] ), .A3(\priority[122] ), .ZN(new_n1555_));
  NAND3_X1   g1170(.A1(new_n1555_), .A2(new_n759_), .A3(new_n1553_), .ZN(new_n1556_));
  NOR2_X1    g1171(.A1(new_n749_), .A2(\req[121] ), .ZN(new_n1557_));
  INV_X1     g1172(.I(new_n753_), .ZN(new_n1558_));
  NOR2_X1    g1173(.A1(new_n1558_), .A2(new_n1557_), .ZN(new_n1559_));
  OAI21_X1   g1174(.A1(new_n763_), .A2(\req[124] ), .B(new_n771_), .ZN(new_n1560_));
  NOR3_X1    g1175(.A1(new_n1559_), .A2(new_n766_), .A3(new_n1560_), .ZN(new_n1561_));
  OAI21_X1   g1176(.A1(new_n1550_), .A2(new_n1556_), .B(new_n1561_), .ZN(new_n1562_));
  NOR2_X1    g1177(.A1(\priority[0] ), .A2(\priority[127] ), .ZN(new_n1563_));
  OAI21_X1   g1178(.A1(new_n767_), .A2(\req[126] ), .B(new_n1563_), .ZN(new_n1564_));
  NOR3_X1    g1179(.A1(new_n392_), .A2(\priority[2] ), .A3(\priority[3] ), .ZN(new_n1565_));
  NOR2_X1    g1180(.A1(\req[0] ), .A2(\req[1] ), .ZN(new_n1566_));
  INV_X1     g1181(.I(new_n1566_), .ZN(new_n1567_));
  NOR2_X1    g1182(.A1(new_n1567_), .A2(new_n778_), .ZN(new_n1568_));
  NAND3_X1   g1183(.A1(new_n1565_), .A2(new_n1568_), .A3(new_n1564_), .ZN(new_n1569_));
  INV_X1     g1184(.I(new_n1569_), .ZN(new_n1570_));
  NOR2_X1    g1185(.A1(new_n1138_), .A2(\req[2] ), .ZN(new_n1571_));
  NAND2_X1   g1186(.A1(new_n1571_), .A2(new_n388_), .ZN(new_n1572_));
  AOI21_X1   g1187(.A1(new_n1562_), .A2(new_n1570_), .B(new_n1572_), .ZN(\grant[3] ));
  INV_X1     g1188(.I(new_n788_), .ZN(new_n1574_));
  OAI21_X1   g1189(.A1(new_n404_), .A2(\req[8] ), .B(new_n800_), .ZN(new_n1575_));
  AOI21_X1   g1190(.A1(new_n1133_), .A2(\priority[5] ), .B(\priority[6] ), .ZN(new_n1576_));
  NOR4_X1    g1191(.A1(new_n795_), .A2(new_n1574_), .A3(new_n1575_), .A4(new_n1576_), .ZN(new_n1577_));
  INV_X1     g1192(.I(\req[10] ), .ZN(new_n1578_));
  NAND2_X1   g1193(.A1(new_n1578_), .A2(\priority[10] ), .ZN(new_n1579_));
  NAND3_X1   g1194(.A1(new_n1579_), .A2(new_n419_), .A3(new_n810_), .ZN(new_n1580_));
  NOR2_X1    g1195(.A1(new_n412_), .A2(\req[13] ), .ZN(new_n1581_));
  NOR3_X1    g1196(.A1(new_n1581_), .A2(\priority[14] ), .A3(\priority[15] ), .ZN(new_n1582_));
  NAND3_X1   g1197(.A1(new_n1582_), .A2(new_n814_), .A3(new_n1580_), .ZN(new_n1583_));
  NOR2_X1    g1198(.A1(new_n804_), .A2(\req[14] ), .ZN(new_n1584_));
  INV_X1     g1199(.I(new_n808_), .ZN(new_n1585_));
  NOR2_X1    g1200(.A1(new_n1585_), .A2(new_n1584_), .ZN(new_n1586_));
  OAI21_X1   g1201(.A1(new_n431_), .A2(\req[17] ), .B(new_n824_), .ZN(new_n1587_));
  NOR3_X1    g1202(.A1(new_n1586_), .A2(new_n819_), .A3(new_n1587_), .ZN(new_n1588_));
  OAI21_X1   g1203(.A1(new_n1583_), .A2(new_n1577_), .B(new_n1588_), .ZN(new_n1589_));
  INV_X1     g1204(.I(\req[19] ), .ZN(new_n1590_));
  NAND2_X1   g1205(.A1(new_n1590_), .A2(\priority[19] ), .ZN(new_n1591_));
  NAND3_X1   g1206(.A1(new_n1591_), .A2(new_n447_), .A3(new_n835_), .ZN(new_n1592_));
  NOR2_X1    g1207(.A1(new_n440_), .A2(\req[22] ), .ZN(new_n1593_));
  NOR3_X1    g1208(.A1(new_n1593_), .A2(\priority[23] ), .A3(\priority[24] ), .ZN(new_n1594_));
  NAND3_X1   g1209(.A1(new_n1594_), .A2(new_n839_), .A3(new_n1592_), .ZN(new_n1595_));
  INV_X1     g1210(.I(new_n1595_), .ZN(new_n1596_));
  NOR2_X1    g1211(.A1(new_n829_), .A2(\req[23] ), .ZN(new_n1597_));
  INV_X1     g1212(.I(new_n833_), .ZN(new_n1598_));
  NOR2_X1    g1213(.A1(new_n1598_), .A2(new_n1597_), .ZN(new_n1599_));
  OAI21_X1   g1214(.A1(new_n460_), .A2(\req[26] ), .B(new_n850_), .ZN(new_n1600_));
  NOR3_X1    g1215(.A1(new_n1599_), .A2(new_n845_), .A3(new_n1600_), .ZN(new_n1601_));
  INV_X1     g1216(.I(new_n1601_), .ZN(new_n1602_));
  AOI21_X1   g1217(.A1(new_n1589_), .A2(new_n1596_), .B(new_n1602_), .ZN(new_n1603_));
  INV_X1     g1218(.I(\req[28] ), .ZN(new_n1604_));
  NAND2_X1   g1219(.A1(new_n1604_), .A2(\priority[28] ), .ZN(new_n1605_));
  NAND3_X1   g1220(.A1(new_n1605_), .A2(new_n475_), .A3(new_n860_), .ZN(new_n1606_));
  NOR2_X1    g1221(.A1(new_n468_), .A2(\req[31] ), .ZN(new_n1607_));
  NOR3_X1    g1222(.A1(new_n1607_), .A2(\priority[32] ), .A3(\priority[33] ), .ZN(new_n1608_));
  NAND3_X1   g1223(.A1(new_n1608_), .A2(new_n864_), .A3(new_n1606_), .ZN(new_n1609_));
  NOR2_X1    g1224(.A1(new_n854_), .A2(\req[32] ), .ZN(new_n1610_));
  INV_X1     g1225(.I(new_n858_), .ZN(new_n1611_));
  NOR2_X1    g1226(.A1(new_n1611_), .A2(new_n1610_), .ZN(new_n1612_));
  OAI21_X1   g1227(.A1(new_n487_), .A2(\req[35] ), .B(new_n874_), .ZN(new_n1613_));
  NOR3_X1    g1228(.A1(new_n1612_), .A2(new_n869_), .A3(new_n1613_), .ZN(new_n1614_));
  OAI21_X1   g1229(.A1(new_n1603_), .A2(new_n1609_), .B(new_n1614_), .ZN(new_n1615_));
  INV_X1     g1230(.I(\req[37] ), .ZN(new_n1616_));
  NAND2_X1   g1231(.A1(new_n1616_), .A2(\priority[37] ), .ZN(new_n1617_));
  NAND3_X1   g1232(.A1(new_n1617_), .A2(new_n503_), .A3(new_n885_), .ZN(new_n1618_));
  NOR2_X1    g1233(.A1(new_n496_), .A2(\req[40] ), .ZN(new_n1619_));
  NOR3_X1    g1234(.A1(new_n1619_), .A2(\priority[41] ), .A3(\priority[42] ), .ZN(new_n1620_));
  NAND3_X1   g1235(.A1(new_n1620_), .A2(new_n889_), .A3(new_n1618_), .ZN(new_n1621_));
  INV_X1     g1236(.I(new_n1621_), .ZN(new_n1622_));
  NOR2_X1    g1237(.A1(new_n879_), .A2(\req[41] ), .ZN(new_n1623_));
  INV_X1     g1238(.I(new_n883_), .ZN(new_n1624_));
  NOR2_X1    g1239(.A1(new_n1624_), .A2(new_n1623_), .ZN(new_n1625_));
  OAI21_X1   g1240(.A1(new_n516_), .A2(\req[44] ), .B(new_n900_), .ZN(new_n1626_));
  NOR3_X1    g1241(.A1(new_n1625_), .A2(new_n895_), .A3(new_n1626_), .ZN(new_n1627_));
  INV_X1     g1242(.I(new_n1627_), .ZN(new_n1628_));
  AOI21_X1   g1243(.A1(new_n1615_), .A2(new_n1622_), .B(new_n1628_), .ZN(new_n1629_));
  INV_X1     g1244(.I(\req[46] ), .ZN(new_n1630_));
  NAND2_X1   g1245(.A1(new_n1630_), .A2(\priority[46] ), .ZN(new_n1631_));
  NAND3_X1   g1246(.A1(new_n1631_), .A2(new_n531_), .A3(new_n910_), .ZN(new_n1632_));
  NOR2_X1    g1247(.A1(new_n524_), .A2(\req[49] ), .ZN(new_n1633_));
  NOR3_X1    g1248(.A1(new_n1633_), .A2(\priority[50] ), .A3(\priority[51] ), .ZN(new_n1634_));
  NAND3_X1   g1249(.A1(new_n1634_), .A2(new_n914_), .A3(new_n1632_), .ZN(new_n1635_));
  NOR2_X1    g1250(.A1(new_n904_), .A2(\req[50] ), .ZN(new_n1636_));
  INV_X1     g1251(.I(new_n908_), .ZN(new_n1637_));
  NOR2_X1    g1252(.A1(new_n1637_), .A2(new_n1636_), .ZN(new_n1638_));
  OAI21_X1   g1253(.A1(new_n543_), .A2(\req[53] ), .B(new_n924_), .ZN(new_n1639_));
  NOR3_X1    g1254(.A1(new_n1638_), .A2(new_n919_), .A3(new_n1639_), .ZN(new_n1640_));
  OAI21_X1   g1255(.A1(new_n1629_), .A2(new_n1635_), .B(new_n1640_), .ZN(new_n1641_));
  INV_X1     g1256(.I(\req[55] ), .ZN(new_n1642_));
  NAND2_X1   g1257(.A1(new_n1642_), .A2(\priority[55] ), .ZN(new_n1643_));
  NAND3_X1   g1258(.A1(new_n1643_), .A2(new_n559_), .A3(new_n935_), .ZN(new_n1644_));
  NOR2_X1    g1259(.A1(new_n552_), .A2(\req[58] ), .ZN(new_n1645_));
  NOR3_X1    g1260(.A1(new_n1645_), .A2(\priority[59] ), .A3(\priority[60] ), .ZN(new_n1646_));
  NAND3_X1   g1261(.A1(new_n1646_), .A2(new_n939_), .A3(new_n1644_), .ZN(new_n1647_));
  INV_X1     g1262(.I(new_n1647_), .ZN(new_n1648_));
  NOR2_X1    g1263(.A1(new_n929_), .A2(\req[59] ), .ZN(new_n1649_));
  INV_X1     g1264(.I(new_n933_), .ZN(new_n1650_));
  NOR2_X1    g1265(.A1(new_n1650_), .A2(new_n1649_), .ZN(new_n1651_));
  OAI21_X1   g1266(.A1(new_n572_), .A2(\req[62] ), .B(new_n950_), .ZN(new_n1652_));
  NOR3_X1    g1267(.A1(new_n1651_), .A2(new_n945_), .A3(new_n1652_), .ZN(new_n1653_));
  INV_X1     g1268(.I(new_n1653_), .ZN(new_n1654_));
  AOI21_X1   g1269(.A1(new_n1641_), .A2(new_n1648_), .B(new_n1654_), .ZN(new_n1655_));
  INV_X1     g1270(.I(\req[64] ), .ZN(new_n1656_));
  NAND2_X1   g1271(.A1(new_n1656_), .A2(\priority[64] ), .ZN(new_n1657_));
  NAND3_X1   g1272(.A1(new_n1657_), .A2(new_n587_), .A3(new_n960_), .ZN(new_n1658_));
  NOR2_X1    g1273(.A1(new_n580_), .A2(\req[67] ), .ZN(new_n1659_));
  NOR3_X1    g1274(.A1(new_n1659_), .A2(\priority[68] ), .A3(\priority[69] ), .ZN(new_n1660_));
  NAND3_X1   g1275(.A1(new_n1660_), .A2(new_n964_), .A3(new_n1658_), .ZN(new_n1661_));
  NOR2_X1    g1276(.A1(new_n954_), .A2(\req[68] ), .ZN(new_n1662_));
  INV_X1     g1277(.I(new_n958_), .ZN(new_n1663_));
  NOR2_X1    g1278(.A1(new_n1663_), .A2(new_n1662_), .ZN(new_n1664_));
  OAI21_X1   g1279(.A1(new_n599_), .A2(\req[71] ), .B(new_n974_), .ZN(new_n1665_));
  NOR3_X1    g1280(.A1(new_n1664_), .A2(new_n969_), .A3(new_n1665_), .ZN(new_n1666_));
  OAI21_X1   g1281(.A1(new_n1655_), .A2(new_n1661_), .B(new_n1666_), .ZN(new_n1667_));
  INV_X1     g1282(.I(\req[73] ), .ZN(new_n1668_));
  NAND2_X1   g1283(.A1(new_n1668_), .A2(\priority[73] ), .ZN(new_n1669_));
  NAND3_X1   g1284(.A1(new_n1669_), .A2(new_n615_), .A3(new_n985_), .ZN(new_n1670_));
  NOR2_X1    g1285(.A1(new_n608_), .A2(\req[76] ), .ZN(new_n1671_));
  NOR3_X1    g1286(.A1(new_n1671_), .A2(\priority[77] ), .A3(\priority[78] ), .ZN(new_n1672_));
  NAND3_X1   g1287(.A1(new_n1672_), .A2(new_n989_), .A3(new_n1670_), .ZN(new_n1673_));
  INV_X1     g1288(.I(new_n1673_), .ZN(new_n1674_));
  NOR2_X1    g1289(.A1(new_n979_), .A2(\req[77] ), .ZN(new_n1675_));
  INV_X1     g1290(.I(new_n983_), .ZN(new_n1676_));
  NOR2_X1    g1291(.A1(new_n1676_), .A2(new_n1675_), .ZN(new_n1677_));
  OAI21_X1   g1292(.A1(new_n628_), .A2(\req[80] ), .B(new_n1000_), .ZN(new_n1678_));
  NOR3_X1    g1293(.A1(new_n1677_), .A2(new_n995_), .A3(new_n1678_), .ZN(new_n1679_));
  INV_X1     g1294(.I(new_n1679_), .ZN(new_n1680_));
  AOI21_X1   g1295(.A1(new_n1667_), .A2(new_n1674_), .B(new_n1680_), .ZN(new_n1681_));
  INV_X1     g1296(.I(\req[82] ), .ZN(new_n1682_));
  NAND2_X1   g1297(.A1(new_n1682_), .A2(\priority[82] ), .ZN(new_n1683_));
  NAND3_X1   g1298(.A1(new_n1683_), .A2(new_n643_), .A3(new_n1010_), .ZN(new_n1684_));
  NOR2_X1    g1299(.A1(new_n636_), .A2(\req[85] ), .ZN(new_n1685_));
  NOR3_X1    g1300(.A1(new_n1685_), .A2(\priority[86] ), .A3(\priority[87] ), .ZN(new_n1686_));
  NAND3_X1   g1301(.A1(new_n1686_), .A2(new_n1014_), .A3(new_n1684_), .ZN(new_n1687_));
  NOR2_X1    g1302(.A1(new_n1004_), .A2(\req[86] ), .ZN(new_n1688_));
  INV_X1     g1303(.I(new_n1008_), .ZN(new_n1689_));
  NOR2_X1    g1304(.A1(new_n1689_), .A2(new_n1688_), .ZN(new_n1690_));
  OAI21_X1   g1305(.A1(new_n655_), .A2(\req[89] ), .B(new_n1024_), .ZN(new_n1691_));
  NOR3_X1    g1306(.A1(new_n1690_), .A2(new_n1019_), .A3(new_n1691_), .ZN(new_n1692_));
  OAI21_X1   g1307(.A1(new_n1681_), .A2(new_n1687_), .B(new_n1692_), .ZN(new_n1693_));
  INV_X1     g1308(.I(\req[91] ), .ZN(new_n1694_));
  NAND2_X1   g1309(.A1(new_n1694_), .A2(\priority[91] ), .ZN(new_n1695_));
  NAND3_X1   g1310(.A1(new_n1695_), .A2(new_n671_), .A3(new_n1035_), .ZN(new_n1696_));
  NOR2_X1    g1311(.A1(new_n664_), .A2(\req[94] ), .ZN(new_n1697_));
  NOR3_X1    g1312(.A1(new_n1697_), .A2(\priority[95] ), .A3(\priority[96] ), .ZN(new_n1698_));
  NAND3_X1   g1313(.A1(new_n1698_), .A2(new_n1039_), .A3(new_n1696_), .ZN(new_n1699_));
  INV_X1     g1314(.I(new_n1699_), .ZN(new_n1700_));
  NOR2_X1    g1315(.A1(new_n1029_), .A2(\req[95] ), .ZN(new_n1701_));
  INV_X1     g1316(.I(new_n1033_), .ZN(new_n1702_));
  NOR2_X1    g1317(.A1(new_n1702_), .A2(new_n1701_), .ZN(new_n1703_));
  OAI21_X1   g1318(.A1(new_n684_), .A2(\req[98] ), .B(new_n1050_), .ZN(new_n1704_));
  NOR3_X1    g1319(.A1(new_n1703_), .A2(new_n1045_), .A3(new_n1704_), .ZN(new_n1705_));
  INV_X1     g1320(.I(new_n1705_), .ZN(new_n1706_));
  AOI21_X1   g1321(.A1(new_n1693_), .A2(new_n1700_), .B(new_n1706_), .ZN(new_n1707_));
  INV_X1     g1322(.I(\req[100] ), .ZN(new_n1708_));
  NAND2_X1   g1323(.A1(new_n1708_), .A2(\priority[100] ), .ZN(new_n1709_));
  NAND3_X1   g1324(.A1(new_n1709_), .A2(new_n699_), .A3(new_n1060_), .ZN(new_n1710_));
  NOR2_X1    g1325(.A1(new_n692_), .A2(\req[103] ), .ZN(new_n1711_));
  NOR3_X1    g1326(.A1(new_n1711_), .A2(\priority[104] ), .A3(\priority[105] ), .ZN(new_n1712_));
  NAND3_X1   g1327(.A1(new_n1712_), .A2(new_n1064_), .A3(new_n1710_), .ZN(new_n1713_));
  NOR2_X1    g1328(.A1(new_n1054_), .A2(\req[104] ), .ZN(new_n1714_));
  INV_X1     g1329(.I(new_n1058_), .ZN(new_n1715_));
  NOR2_X1    g1330(.A1(new_n1715_), .A2(new_n1714_), .ZN(new_n1716_));
  OAI21_X1   g1331(.A1(new_n711_), .A2(\req[107] ), .B(new_n1074_), .ZN(new_n1717_));
  NOR3_X1    g1332(.A1(new_n1716_), .A2(new_n1069_), .A3(new_n1717_), .ZN(new_n1718_));
  OAI21_X1   g1333(.A1(new_n1707_), .A2(new_n1713_), .B(new_n1718_), .ZN(new_n1719_));
  INV_X1     g1334(.I(\req[109] ), .ZN(new_n1720_));
  NAND2_X1   g1335(.A1(new_n1720_), .A2(\priority[109] ), .ZN(new_n1721_));
  NAND3_X1   g1336(.A1(new_n1721_), .A2(new_n727_), .A3(new_n1085_), .ZN(new_n1722_));
  NOR2_X1    g1337(.A1(new_n720_), .A2(\req[112] ), .ZN(new_n1723_));
  NOR3_X1    g1338(.A1(new_n1723_), .A2(\priority[113] ), .A3(\priority[114] ), .ZN(new_n1724_));
  NAND3_X1   g1339(.A1(new_n1724_), .A2(new_n1089_), .A3(new_n1722_), .ZN(new_n1725_));
  INV_X1     g1340(.I(new_n1725_), .ZN(new_n1726_));
  NOR2_X1    g1341(.A1(new_n1079_), .A2(\req[113] ), .ZN(new_n1727_));
  INV_X1     g1342(.I(new_n1083_), .ZN(new_n1728_));
  NOR2_X1    g1343(.A1(new_n1728_), .A2(new_n1727_), .ZN(new_n1729_));
  OAI21_X1   g1344(.A1(new_n740_), .A2(\req[116] ), .B(new_n1100_), .ZN(new_n1730_));
  NOR3_X1    g1345(.A1(new_n1729_), .A2(new_n1095_), .A3(new_n1730_), .ZN(new_n1731_));
  INV_X1     g1346(.I(new_n1731_), .ZN(new_n1732_));
  AOI21_X1   g1347(.A1(new_n1719_), .A2(new_n1726_), .B(new_n1732_), .ZN(new_n1733_));
  INV_X1     g1348(.I(\req[118] ), .ZN(new_n1734_));
  NAND2_X1   g1349(.A1(new_n1734_), .A2(\priority[118] ), .ZN(new_n1735_));
  NAND3_X1   g1350(.A1(new_n1735_), .A2(new_n755_), .A3(new_n1110_), .ZN(new_n1736_));
  NOR2_X1    g1351(.A1(new_n748_), .A2(\req[121] ), .ZN(new_n1737_));
  NOR3_X1    g1352(.A1(new_n1737_), .A2(\priority[122] ), .A3(\priority[123] ), .ZN(new_n1738_));
  NAND3_X1   g1353(.A1(new_n1738_), .A2(new_n1114_), .A3(new_n1736_), .ZN(new_n1739_));
  NOR2_X1    g1354(.A1(new_n1104_), .A2(\req[122] ), .ZN(new_n1740_));
  INV_X1     g1355(.I(new_n1108_), .ZN(new_n1741_));
  NOR2_X1    g1356(.A1(new_n1741_), .A2(new_n1740_), .ZN(new_n1742_));
  OAI21_X1   g1357(.A1(new_n767_), .A2(\req[125] ), .B(new_n1124_), .ZN(new_n1743_));
  NOR3_X1    g1358(.A1(new_n1742_), .A2(new_n1119_), .A3(new_n1743_), .ZN(new_n1744_));
  OAI21_X1   g1359(.A1(new_n1733_), .A2(new_n1739_), .B(new_n1744_), .ZN(new_n1745_));
  NOR2_X1    g1360(.A1(\priority[0] ), .A2(\priority[1] ), .ZN(new_n1746_));
  OAI21_X1   g1361(.A1(new_n1120_), .A2(\req[127] ), .B(new_n1746_), .ZN(new_n1747_));
  NOR3_X1    g1362(.A1(new_n786_), .A2(\priority[3] ), .A3(\priority[4] ), .ZN(new_n1748_));
  NOR3_X1    g1363(.A1(new_n1130_), .A2(\req[1] ), .A3(\req[2] ), .ZN(new_n1749_));
  NAND3_X1   g1364(.A1(new_n1748_), .A2(new_n1749_), .A3(new_n1747_), .ZN(new_n1750_));
  INV_X1     g1365(.I(new_n1750_), .ZN(new_n1751_));
  NOR2_X1    g1366(.A1(new_n386_), .A2(\req[3] ), .ZN(new_n1752_));
  NAND2_X1   g1367(.A1(new_n1752_), .A2(new_n782_), .ZN(new_n1753_));
  AOI21_X1   g1368(.A1(new_n1745_), .A2(new_n1751_), .B(new_n1753_), .ZN(\grant[4] ));
  NOR2_X1    g1369(.A1(new_n781_), .A2(\req[6] ), .ZN(new_n1755_));
  NOR2_X1    g1370(.A1(new_n1755_), .A2(\priority[7] ), .ZN(new_n1756_));
  INV_X1     g1371(.I(new_n1136_), .ZN(new_n1757_));
  NOR2_X1    g1372(.A1(\req[10] ), .A2(\req[11] ), .ZN(new_n1758_));
  OAI21_X1   g1373(.A1(new_n796_), .A2(\req[9] ), .B(new_n1758_), .ZN(new_n1759_));
  NOR4_X1    g1374(.A1(new_n1145_), .A2(new_n1756_), .A3(new_n1759_), .A4(new_n1757_), .ZN(new_n1760_));
  INV_X1     g1375(.I(\req[11] ), .ZN(new_n1761_));
  NAND2_X1   g1376(.A1(new_n1761_), .A2(\priority[11] ), .ZN(new_n1762_));
  NAND3_X1   g1377(.A1(new_n1762_), .A2(new_n810_), .A3(new_n412_), .ZN(new_n1763_));
  NOR2_X1    g1378(.A1(new_n413_), .A2(\req[14] ), .ZN(new_n1764_));
  NOR3_X1    g1379(.A1(new_n1764_), .A2(\priority[15] ), .A3(\priority[16] ), .ZN(new_n1765_));
  NAND3_X1   g1380(.A1(new_n1765_), .A2(new_n1157_), .A3(new_n1763_), .ZN(new_n1766_));
  NOR2_X1    g1381(.A1(new_n426_), .A2(\req[15] ), .ZN(new_n1767_));
  INV_X1     g1382(.I(new_n1154_), .ZN(new_n1768_));
  NOR2_X1    g1383(.A1(new_n1768_), .A2(new_n1767_), .ZN(new_n1769_));
  NOR2_X1    g1384(.A1(\req[19] ), .A2(\req[20] ), .ZN(new_n1770_));
  OAI21_X1   g1385(.A1(new_n820_), .A2(\req[18] ), .B(new_n1770_), .ZN(new_n1771_));
  NOR3_X1    g1386(.A1(new_n1769_), .A2(new_n1162_), .A3(new_n1771_), .ZN(new_n1772_));
  OAI21_X1   g1387(.A1(new_n1766_), .A2(new_n1760_), .B(new_n1772_), .ZN(new_n1773_));
  INV_X1     g1388(.I(\req[20] ), .ZN(new_n1774_));
  NAND2_X1   g1389(.A1(new_n1774_), .A2(\priority[20] ), .ZN(new_n1775_));
  NAND3_X1   g1390(.A1(new_n1775_), .A2(new_n835_), .A3(new_n440_), .ZN(new_n1776_));
  NOR2_X1    g1391(.A1(new_n441_), .A2(\req[23] ), .ZN(new_n1777_));
  NOR3_X1    g1392(.A1(new_n1777_), .A2(\priority[24] ), .A3(\priority[25] ), .ZN(new_n1778_));
  NAND3_X1   g1393(.A1(new_n1778_), .A2(new_n1175_), .A3(new_n1776_), .ZN(new_n1779_));
  INV_X1     g1394(.I(new_n1779_), .ZN(new_n1780_));
  NOR2_X1    g1395(.A1(new_n455_), .A2(\req[24] ), .ZN(new_n1781_));
  INV_X1     g1396(.I(new_n1172_), .ZN(new_n1782_));
  NOR2_X1    g1397(.A1(new_n1782_), .A2(new_n1781_), .ZN(new_n1783_));
  NOR2_X1    g1398(.A1(\req[28] ), .A2(\req[29] ), .ZN(new_n1784_));
  OAI21_X1   g1399(.A1(new_n846_), .A2(\req[27] ), .B(new_n1784_), .ZN(new_n1785_));
  NOR3_X1    g1400(.A1(new_n1783_), .A2(new_n1181_), .A3(new_n1785_), .ZN(new_n1786_));
  INV_X1     g1401(.I(new_n1786_), .ZN(new_n1787_));
  AOI21_X1   g1402(.A1(new_n1773_), .A2(new_n1780_), .B(new_n1787_), .ZN(new_n1788_));
  INV_X1     g1403(.I(\req[29] ), .ZN(new_n1789_));
  NAND2_X1   g1404(.A1(new_n1789_), .A2(\priority[29] ), .ZN(new_n1790_));
  NAND3_X1   g1405(.A1(new_n1790_), .A2(new_n860_), .A3(new_n468_), .ZN(new_n1791_));
  NOR2_X1    g1406(.A1(new_n469_), .A2(\req[32] ), .ZN(new_n1792_));
  NOR3_X1    g1407(.A1(new_n1792_), .A2(\priority[33] ), .A3(\priority[34] ), .ZN(new_n1793_));
  NAND3_X1   g1408(.A1(new_n1793_), .A2(new_n1193_), .A3(new_n1791_), .ZN(new_n1794_));
  NOR2_X1    g1409(.A1(new_n482_), .A2(\req[33] ), .ZN(new_n1795_));
  INV_X1     g1410(.I(new_n1190_), .ZN(new_n1796_));
  NOR2_X1    g1411(.A1(new_n1796_), .A2(new_n1795_), .ZN(new_n1797_));
  NOR2_X1    g1412(.A1(\req[37] ), .A2(\req[38] ), .ZN(new_n1798_));
  OAI21_X1   g1413(.A1(new_n870_), .A2(\req[36] ), .B(new_n1798_), .ZN(new_n1799_));
  NOR3_X1    g1414(.A1(new_n1797_), .A2(new_n1198_), .A3(new_n1799_), .ZN(new_n1800_));
  OAI21_X1   g1415(.A1(new_n1788_), .A2(new_n1794_), .B(new_n1800_), .ZN(new_n1801_));
  INV_X1     g1416(.I(\req[38] ), .ZN(new_n1802_));
  NAND2_X1   g1417(.A1(new_n1802_), .A2(\priority[38] ), .ZN(new_n1803_));
  NAND3_X1   g1418(.A1(new_n1803_), .A2(new_n885_), .A3(new_n496_), .ZN(new_n1804_));
  NOR2_X1    g1419(.A1(new_n497_), .A2(\req[41] ), .ZN(new_n1805_));
  NOR3_X1    g1420(.A1(new_n1805_), .A2(\priority[42] ), .A3(\priority[43] ), .ZN(new_n1806_));
  NAND3_X1   g1421(.A1(new_n1806_), .A2(new_n1211_), .A3(new_n1804_), .ZN(new_n1807_));
  INV_X1     g1422(.I(new_n1807_), .ZN(new_n1808_));
  NOR2_X1    g1423(.A1(new_n511_), .A2(\req[42] ), .ZN(new_n1809_));
  INV_X1     g1424(.I(new_n1208_), .ZN(new_n1810_));
  NOR2_X1    g1425(.A1(new_n1810_), .A2(new_n1809_), .ZN(new_n1811_));
  NOR2_X1    g1426(.A1(\req[46] ), .A2(\req[47] ), .ZN(new_n1812_));
  OAI21_X1   g1427(.A1(new_n896_), .A2(\req[45] ), .B(new_n1812_), .ZN(new_n1813_));
  NOR3_X1    g1428(.A1(new_n1811_), .A2(new_n1217_), .A3(new_n1813_), .ZN(new_n1814_));
  INV_X1     g1429(.I(new_n1814_), .ZN(new_n1815_));
  AOI21_X1   g1430(.A1(new_n1801_), .A2(new_n1808_), .B(new_n1815_), .ZN(new_n1816_));
  INV_X1     g1431(.I(\req[47] ), .ZN(new_n1817_));
  NAND2_X1   g1432(.A1(new_n1817_), .A2(\priority[47] ), .ZN(new_n1818_));
  NAND3_X1   g1433(.A1(new_n1818_), .A2(new_n910_), .A3(new_n524_), .ZN(new_n1819_));
  NOR2_X1    g1434(.A1(new_n525_), .A2(\req[50] ), .ZN(new_n1820_));
  NOR3_X1    g1435(.A1(new_n1820_), .A2(\priority[51] ), .A3(\priority[52] ), .ZN(new_n1821_));
  NAND3_X1   g1436(.A1(new_n1821_), .A2(new_n1229_), .A3(new_n1819_), .ZN(new_n1822_));
  NOR2_X1    g1437(.A1(new_n538_), .A2(\req[51] ), .ZN(new_n1823_));
  INV_X1     g1438(.I(new_n1226_), .ZN(new_n1824_));
  NOR2_X1    g1439(.A1(new_n1824_), .A2(new_n1823_), .ZN(new_n1825_));
  NOR2_X1    g1440(.A1(\req[55] ), .A2(\req[56] ), .ZN(new_n1826_));
  OAI21_X1   g1441(.A1(new_n920_), .A2(\req[54] ), .B(new_n1826_), .ZN(new_n1827_));
  NOR3_X1    g1442(.A1(new_n1825_), .A2(new_n1234_), .A3(new_n1827_), .ZN(new_n1828_));
  OAI21_X1   g1443(.A1(new_n1816_), .A2(new_n1822_), .B(new_n1828_), .ZN(new_n1829_));
  INV_X1     g1444(.I(\req[56] ), .ZN(new_n1830_));
  NAND2_X1   g1445(.A1(new_n1830_), .A2(\priority[56] ), .ZN(new_n1831_));
  NAND3_X1   g1446(.A1(new_n1831_), .A2(new_n935_), .A3(new_n552_), .ZN(new_n1832_));
  NOR2_X1    g1447(.A1(new_n553_), .A2(\req[59] ), .ZN(new_n1833_));
  NOR3_X1    g1448(.A1(new_n1833_), .A2(\priority[60] ), .A3(\priority[61] ), .ZN(new_n1834_));
  NAND3_X1   g1449(.A1(new_n1834_), .A2(new_n1247_), .A3(new_n1832_), .ZN(new_n1835_));
  INV_X1     g1450(.I(new_n1835_), .ZN(new_n1836_));
  NOR2_X1    g1451(.A1(new_n567_), .A2(\req[60] ), .ZN(new_n1837_));
  INV_X1     g1452(.I(new_n1244_), .ZN(new_n1838_));
  NOR2_X1    g1453(.A1(new_n1838_), .A2(new_n1837_), .ZN(new_n1839_));
  NOR2_X1    g1454(.A1(\req[64] ), .A2(\req[65] ), .ZN(new_n1840_));
  OAI21_X1   g1455(.A1(new_n946_), .A2(\req[63] ), .B(new_n1840_), .ZN(new_n1841_));
  NOR3_X1    g1456(.A1(new_n1839_), .A2(new_n1253_), .A3(new_n1841_), .ZN(new_n1842_));
  INV_X1     g1457(.I(new_n1842_), .ZN(new_n1843_));
  AOI21_X1   g1458(.A1(new_n1829_), .A2(new_n1836_), .B(new_n1843_), .ZN(new_n1844_));
  INV_X1     g1459(.I(\req[65] ), .ZN(new_n1845_));
  NAND2_X1   g1460(.A1(new_n1845_), .A2(\priority[65] ), .ZN(new_n1846_));
  NAND3_X1   g1461(.A1(new_n1846_), .A2(new_n960_), .A3(new_n580_), .ZN(new_n1847_));
  NOR2_X1    g1462(.A1(new_n581_), .A2(\req[68] ), .ZN(new_n1848_));
  NOR3_X1    g1463(.A1(new_n1848_), .A2(\priority[69] ), .A3(\priority[70] ), .ZN(new_n1849_));
  NAND3_X1   g1464(.A1(new_n1849_), .A2(new_n1265_), .A3(new_n1847_), .ZN(new_n1850_));
  NOR2_X1    g1465(.A1(new_n594_), .A2(\req[69] ), .ZN(new_n1851_));
  INV_X1     g1466(.I(new_n1262_), .ZN(new_n1852_));
  NOR2_X1    g1467(.A1(new_n1852_), .A2(new_n1851_), .ZN(new_n1853_));
  NOR2_X1    g1468(.A1(\req[73] ), .A2(\req[74] ), .ZN(new_n1854_));
  OAI21_X1   g1469(.A1(new_n970_), .A2(\req[72] ), .B(new_n1854_), .ZN(new_n1855_));
  NOR3_X1    g1470(.A1(new_n1853_), .A2(new_n1270_), .A3(new_n1855_), .ZN(new_n1856_));
  OAI21_X1   g1471(.A1(new_n1844_), .A2(new_n1850_), .B(new_n1856_), .ZN(new_n1857_));
  INV_X1     g1472(.I(\req[74] ), .ZN(new_n1858_));
  NAND2_X1   g1473(.A1(new_n1858_), .A2(\priority[74] ), .ZN(new_n1859_));
  NAND3_X1   g1474(.A1(new_n1859_), .A2(new_n985_), .A3(new_n608_), .ZN(new_n1860_));
  NOR2_X1    g1475(.A1(new_n609_), .A2(\req[77] ), .ZN(new_n1861_));
  NOR3_X1    g1476(.A1(new_n1861_), .A2(\priority[78] ), .A3(\priority[79] ), .ZN(new_n1862_));
  NAND3_X1   g1477(.A1(new_n1862_), .A2(new_n1283_), .A3(new_n1860_), .ZN(new_n1863_));
  INV_X1     g1478(.I(new_n1863_), .ZN(new_n1864_));
  NOR2_X1    g1479(.A1(new_n623_), .A2(\req[78] ), .ZN(new_n1865_));
  INV_X1     g1480(.I(new_n1280_), .ZN(new_n1866_));
  NOR2_X1    g1481(.A1(new_n1866_), .A2(new_n1865_), .ZN(new_n1867_));
  NOR2_X1    g1482(.A1(\req[82] ), .A2(\req[83] ), .ZN(new_n1868_));
  OAI21_X1   g1483(.A1(new_n996_), .A2(\req[81] ), .B(new_n1868_), .ZN(new_n1869_));
  NOR3_X1    g1484(.A1(new_n1867_), .A2(new_n1289_), .A3(new_n1869_), .ZN(new_n1870_));
  INV_X1     g1485(.I(new_n1870_), .ZN(new_n1871_));
  AOI21_X1   g1486(.A1(new_n1857_), .A2(new_n1864_), .B(new_n1871_), .ZN(new_n1872_));
  INV_X1     g1487(.I(\req[83] ), .ZN(new_n1873_));
  NAND2_X1   g1488(.A1(new_n1873_), .A2(\priority[83] ), .ZN(new_n1874_));
  NAND3_X1   g1489(.A1(new_n1874_), .A2(new_n1010_), .A3(new_n636_), .ZN(new_n1875_));
  NOR2_X1    g1490(.A1(new_n637_), .A2(\req[86] ), .ZN(new_n1876_));
  NOR3_X1    g1491(.A1(new_n1876_), .A2(\priority[87] ), .A3(\priority[88] ), .ZN(new_n1877_));
  NAND3_X1   g1492(.A1(new_n1877_), .A2(new_n1301_), .A3(new_n1875_), .ZN(new_n1878_));
  NOR2_X1    g1493(.A1(new_n650_), .A2(\req[87] ), .ZN(new_n1879_));
  INV_X1     g1494(.I(new_n1298_), .ZN(new_n1880_));
  NOR2_X1    g1495(.A1(new_n1880_), .A2(new_n1879_), .ZN(new_n1881_));
  NOR2_X1    g1496(.A1(\req[91] ), .A2(\req[92] ), .ZN(new_n1882_));
  OAI21_X1   g1497(.A1(new_n1020_), .A2(\req[90] ), .B(new_n1882_), .ZN(new_n1883_));
  NOR3_X1    g1498(.A1(new_n1881_), .A2(new_n1306_), .A3(new_n1883_), .ZN(new_n1884_));
  OAI21_X1   g1499(.A1(new_n1872_), .A2(new_n1878_), .B(new_n1884_), .ZN(new_n1885_));
  INV_X1     g1500(.I(\req[92] ), .ZN(new_n1886_));
  NAND2_X1   g1501(.A1(new_n1886_), .A2(\priority[92] ), .ZN(new_n1887_));
  NAND3_X1   g1502(.A1(new_n1887_), .A2(new_n1035_), .A3(new_n664_), .ZN(new_n1888_));
  NOR2_X1    g1503(.A1(new_n665_), .A2(\req[95] ), .ZN(new_n1889_));
  NOR3_X1    g1504(.A1(new_n1889_), .A2(\priority[96] ), .A3(\priority[97] ), .ZN(new_n1890_));
  NAND3_X1   g1505(.A1(new_n1890_), .A2(new_n1319_), .A3(new_n1888_), .ZN(new_n1891_));
  INV_X1     g1506(.I(new_n1891_), .ZN(new_n1892_));
  NOR2_X1    g1507(.A1(new_n679_), .A2(\req[96] ), .ZN(new_n1893_));
  INV_X1     g1508(.I(new_n1316_), .ZN(new_n1894_));
  NOR2_X1    g1509(.A1(new_n1894_), .A2(new_n1893_), .ZN(new_n1895_));
  NOR2_X1    g1510(.A1(\req[100] ), .A2(\req[101] ), .ZN(new_n1896_));
  OAI21_X1   g1511(.A1(new_n1046_), .A2(\req[99] ), .B(new_n1896_), .ZN(new_n1897_));
  NOR3_X1    g1512(.A1(new_n1895_), .A2(new_n1325_), .A3(new_n1897_), .ZN(new_n1898_));
  INV_X1     g1513(.I(new_n1898_), .ZN(new_n1899_));
  AOI21_X1   g1514(.A1(new_n1885_), .A2(new_n1892_), .B(new_n1899_), .ZN(new_n1900_));
  INV_X1     g1515(.I(\req[101] ), .ZN(new_n1901_));
  NAND2_X1   g1516(.A1(new_n1901_), .A2(\priority[101] ), .ZN(new_n1902_));
  NAND3_X1   g1517(.A1(new_n1902_), .A2(new_n1060_), .A3(new_n692_), .ZN(new_n1903_));
  NOR2_X1    g1518(.A1(new_n693_), .A2(\req[104] ), .ZN(new_n1904_));
  NOR3_X1    g1519(.A1(new_n1904_), .A2(\priority[105] ), .A3(\priority[106] ), .ZN(new_n1905_));
  NAND3_X1   g1520(.A1(new_n1905_), .A2(new_n1337_), .A3(new_n1903_), .ZN(new_n1906_));
  NOR2_X1    g1521(.A1(new_n706_), .A2(\req[105] ), .ZN(new_n1907_));
  INV_X1     g1522(.I(new_n1334_), .ZN(new_n1908_));
  NOR2_X1    g1523(.A1(new_n1908_), .A2(new_n1907_), .ZN(new_n1909_));
  NOR2_X1    g1524(.A1(\req[109] ), .A2(\req[110] ), .ZN(new_n1910_));
  OAI21_X1   g1525(.A1(new_n1070_), .A2(\req[108] ), .B(new_n1910_), .ZN(new_n1911_));
  NOR3_X1    g1526(.A1(new_n1909_), .A2(new_n1342_), .A3(new_n1911_), .ZN(new_n1912_));
  OAI21_X1   g1527(.A1(new_n1900_), .A2(new_n1906_), .B(new_n1912_), .ZN(new_n1913_));
  INV_X1     g1528(.I(\req[110] ), .ZN(new_n1914_));
  NAND2_X1   g1529(.A1(new_n1914_), .A2(\priority[110] ), .ZN(new_n1915_));
  NAND3_X1   g1530(.A1(new_n1915_), .A2(new_n1085_), .A3(new_n720_), .ZN(new_n1916_));
  NOR2_X1    g1531(.A1(new_n721_), .A2(\req[113] ), .ZN(new_n1917_));
  NOR3_X1    g1532(.A1(new_n1917_), .A2(\priority[114] ), .A3(\priority[115] ), .ZN(new_n1918_));
  NAND3_X1   g1533(.A1(new_n1918_), .A2(new_n1355_), .A3(new_n1916_), .ZN(new_n1919_));
  INV_X1     g1534(.I(new_n1919_), .ZN(new_n1920_));
  NOR2_X1    g1535(.A1(new_n735_), .A2(\req[114] ), .ZN(new_n1921_));
  INV_X1     g1536(.I(new_n1352_), .ZN(new_n1922_));
  NOR2_X1    g1537(.A1(new_n1922_), .A2(new_n1921_), .ZN(new_n1923_));
  NOR2_X1    g1538(.A1(\req[118] ), .A2(\req[119] ), .ZN(new_n1924_));
  OAI21_X1   g1539(.A1(new_n1096_), .A2(\req[117] ), .B(new_n1924_), .ZN(new_n1925_));
  NOR3_X1    g1540(.A1(new_n1923_), .A2(new_n1361_), .A3(new_n1925_), .ZN(new_n1926_));
  INV_X1     g1541(.I(new_n1926_), .ZN(new_n1927_));
  AOI21_X1   g1542(.A1(new_n1913_), .A2(new_n1920_), .B(new_n1927_), .ZN(new_n1928_));
  INV_X1     g1543(.I(\req[119] ), .ZN(new_n1929_));
  NAND2_X1   g1544(.A1(new_n1929_), .A2(\priority[119] ), .ZN(new_n1930_));
  NAND3_X1   g1545(.A1(new_n1930_), .A2(new_n1110_), .A3(new_n748_), .ZN(new_n1931_));
  NOR2_X1    g1546(.A1(new_n749_), .A2(\req[122] ), .ZN(new_n1932_));
  NOR3_X1    g1547(.A1(new_n1932_), .A2(\priority[123] ), .A3(\priority[124] ), .ZN(new_n1933_));
  NAND3_X1   g1548(.A1(new_n1933_), .A2(new_n1373_), .A3(new_n1931_), .ZN(new_n1934_));
  NOR2_X1    g1549(.A1(new_n762_), .A2(\req[123] ), .ZN(new_n1935_));
  INV_X1     g1550(.I(new_n1370_), .ZN(new_n1936_));
  NOR2_X1    g1551(.A1(new_n1936_), .A2(new_n1935_), .ZN(new_n1937_));
  OAI21_X1   g1552(.A1(new_n1120_), .A2(\req[126] ), .B(new_n1382_), .ZN(new_n1938_));
  NOR3_X1    g1553(.A1(new_n1937_), .A2(new_n1378_), .A3(new_n1938_), .ZN(new_n1939_));
  OAI21_X1   g1554(.A1(new_n1928_), .A2(new_n1934_), .B(new_n1939_), .ZN(new_n1940_));
  NOR3_X1    g1555(.A1(new_n1139_), .A2(\priority[4] ), .A3(\priority[5] ), .ZN(new_n1941_));
  NAND2_X1   g1556(.A1(new_n776_), .A2(\priority[0] ), .ZN(new_n1942_));
  NAND3_X1   g1557(.A1(new_n1942_), .A2(new_n391_), .A3(new_n785_), .ZN(new_n1943_));
  NOR2_X1    g1558(.A1(new_n397_), .A2(new_n1388_), .ZN(new_n1944_));
  NAND3_X1   g1559(.A1(new_n1941_), .A2(new_n1944_), .A3(new_n1943_), .ZN(new_n1945_));
  INV_X1     g1560(.I(new_n1945_), .ZN(new_n1946_));
  NOR2_X1    g1561(.A1(new_n387_), .A2(\req[4] ), .ZN(new_n1947_));
  NAND2_X1   g1562(.A1(new_n1947_), .A2(new_n1133_), .ZN(new_n1948_));
  AOI21_X1   g1563(.A1(new_n1940_), .A2(new_n1946_), .B(new_n1948_), .ZN(\grant[5] ));
  OAI21_X1   g1564(.A1(new_n419_), .A2(\req[10] ), .B(new_n421_), .ZN(new_n1950_));
  AOI21_X1   g1565(.A1(new_n793_), .A2(\priority[7] ), .B(\priority[8] ), .ZN(new_n1951_));
  NOR4_X1    g1566(.A1(new_n1397_), .A2(new_n409_), .A3(new_n1950_), .A4(new_n1951_), .ZN(new_n1952_));
  NOR2_X1    g1567(.A1(new_n804_), .A2(\req[15] ), .ZN(new_n1953_));
  NOR2_X1    g1568(.A1(new_n1953_), .A2(\priority[16] ), .ZN(new_n1954_));
  NAND4_X1   g1569(.A1(new_n1403_), .A2(new_n416_), .A3(new_n1954_), .A4(new_n427_), .ZN(new_n1955_));
  OAI21_X1   g1570(.A1(new_n447_), .A2(\req[19] ), .B(new_n449_), .ZN(new_n1956_));
  NOR3_X1    g1571(.A1(new_n437_), .A2(new_n1409_), .A3(new_n1956_), .ZN(new_n1957_));
  OAI21_X1   g1572(.A1(new_n1955_), .A2(new_n1952_), .B(new_n1957_), .ZN(new_n1958_));
  NOR2_X1    g1573(.A1(new_n829_), .A2(\req[24] ), .ZN(new_n1959_));
  NOR2_X1    g1574(.A1(new_n1959_), .A2(\priority[25] ), .ZN(new_n1960_));
  NAND4_X1   g1575(.A1(new_n1416_), .A2(new_n444_), .A3(new_n1960_), .A4(new_n456_), .ZN(new_n1961_));
  INV_X1     g1576(.I(new_n1961_), .ZN(new_n1962_));
  OAI21_X1   g1577(.A1(new_n475_), .A2(\req[28] ), .B(new_n477_), .ZN(new_n1963_));
  NOR3_X1    g1578(.A1(new_n466_), .A2(new_n1423_), .A3(new_n1963_), .ZN(new_n1964_));
  INV_X1     g1579(.I(new_n1964_), .ZN(new_n1965_));
  AOI21_X1   g1580(.A1(new_n1958_), .A2(new_n1962_), .B(new_n1965_), .ZN(new_n1966_));
  NOR2_X1    g1581(.A1(new_n854_), .A2(\req[33] ), .ZN(new_n1967_));
  NOR2_X1    g1582(.A1(new_n1967_), .A2(\priority[34] ), .ZN(new_n1968_));
  NAND4_X1   g1583(.A1(new_n1429_), .A2(new_n472_), .A3(new_n1968_), .A4(new_n483_), .ZN(new_n1969_));
  OAI21_X1   g1584(.A1(new_n503_), .A2(\req[37] ), .B(new_n505_), .ZN(new_n1970_));
  NOR3_X1    g1585(.A1(new_n493_), .A2(new_n1435_), .A3(new_n1970_), .ZN(new_n1971_));
  OAI21_X1   g1586(.A1(new_n1966_), .A2(new_n1969_), .B(new_n1971_), .ZN(new_n1972_));
  NOR2_X1    g1587(.A1(new_n879_), .A2(\req[42] ), .ZN(new_n1973_));
  NOR2_X1    g1588(.A1(new_n1973_), .A2(\priority[43] ), .ZN(new_n1974_));
  NAND4_X1   g1589(.A1(new_n1442_), .A2(new_n500_), .A3(new_n1974_), .A4(new_n512_), .ZN(new_n1975_));
  INV_X1     g1590(.I(new_n1975_), .ZN(new_n1976_));
  OAI21_X1   g1591(.A1(new_n531_), .A2(\req[46] ), .B(new_n533_), .ZN(new_n1977_));
  NOR3_X1    g1592(.A1(new_n522_), .A2(new_n1449_), .A3(new_n1977_), .ZN(new_n1978_));
  INV_X1     g1593(.I(new_n1978_), .ZN(new_n1979_));
  AOI21_X1   g1594(.A1(new_n1972_), .A2(new_n1976_), .B(new_n1979_), .ZN(new_n1980_));
  NOR2_X1    g1595(.A1(new_n904_), .A2(\req[51] ), .ZN(new_n1981_));
  NOR2_X1    g1596(.A1(new_n1981_), .A2(\priority[52] ), .ZN(new_n1982_));
  NAND4_X1   g1597(.A1(new_n1455_), .A2(new_n528_), .A3(new_n1982_), .A4(new_n539_), .ZN(new_n1983_));
  OAI21_X1   g1598(.A1(new_n559_), .A2(\req[55] ), .B(new_n561_), .ZN(new_n1984_));
  NOR3_X1    g1599(.A1(new_n549_), .A2(new_n1461_), .A3(new_n1984_), .ZN(new_n1985_));
  OAI21_X1   g1600(.A1(new_n1980_), .A2(new_n1983_), .B(new_n1985_), .ZN(new_n1986_));
  NOR2_X1    g1601(.A1(new_n929_), .A2(\req[60] ), .ZN(new_n1987_));
  NOR2_X1    g1602(.A1(new_n1987_), .A2(\priority[61] ), .ZN(new_n1988_));
  NAND4_X1   g1603(.A1(new_n1468_), .A2(new_n556_), .A3(new_n1988_), .A4(new_n568_), .ZN(new_n1989_));
  INV_X1     g1604(.I(new_n1989_), .ZN(new_n1990_));
  OAI21_X1   g1605(.A1(new_n587_), .A2(\req[64] ), .B(new_n589_), .ZN(new_n1991_));
  NOR3_X1    g1606(.A1(new_n578_), .A2(new_n1475_), .A3(new_n1991_), .ZN(new_n1992_));
  INV_X1     g1607(.I(new_n1992_), .ZN(new_n1993_));
  AOI21_X1   g1608(.A1(new_n1986_), .A2(new_n1990_), .B(new_n1993_), .ZN(new_n1994_));
  NOR2_X1    g1609(.A1(new_n954_), .A2(\req[69] ), .ZN(new_n1995_));
  NOR2_X1    g1610(.A1(new_n1995_), .A2(\priority[70] ), .ZN(new_n1996_));
  NAND4_X1   g1611(.A1(new_n1481_), .A2(new_n584_), .A3(new_n1996_), .A4(new_n595_), .ZN(new_n1997_));
  OAI21_X1   g1612(.A1(new_n615_), .A2(\req[73] ), .B(new_n617_), .ZN(new_n1998_));
  NOR3_X1    g1613(.A1(new_n605_), .A2(new_n1487_), .A3(new_n1998_), .ZN(new_n1999_));
  OAI21_X1   g1614(.A1(new_n1994_), .A2(new_n1997_), .B(new_n1999_), .ZN(new_n2000_));
  NOR2_X1    g1615(.A1(new_n979_), .A2(\req[78] ), .ZN(new_n2001_));
  NOR2_X1    g1616(.A1(new_n2001_), .A2(\priority[79] ), .ZN(new_n2002_));
  NAND4_X1   g1617(.A1(new_n1494_), .A2(new_n612_), .A3(new_n2002_), .A4(new_n624_), .ZN(new_n2003_));
  INV_X1     g1618(.I(new_n2003_), .ZN(new_n2004_));
  OAI21_X1   g1619(.A1(new_n643_), .A2(\req[82] ), .B(new_n645_), .ZN(new_n2005_));
  NOR3_X1    g1620(.A1(new_n634_), .A2(new_n1501_), .A3(new_n2005_), .ZN(new_n2006_));
  INV_X1     g1621(.I(new_n2006_), .ZN(new_n2007_));
  AOI21_X1   g1622(.A1(new_n2000_), .A2(new_n2004_), .B(new_n2007_), .ZN(new_n2008_));
  NOR2_X1    g1623(.A1(new_n1004_), .A2(\req[87] ), .ZN(new_n2009_));
  NOR2_X1    g1624(.A1(new_n2009_), .A2(\priority[88] ), .ZN(new_n2010_));
  NAND4_X1   g1625(.A1(new_n1507_), .A2(new_n640_), .A3(new_n2010_), .A4(new_n651_), .ZN(new_n2011_));
  OAI21_X1   g1626(.A1(new_n671_), .A2(\req[91] ), .B(new_n673_), .ZN(new_n2012_));
  NOR3_X1    g1627(.A1(new_n661_), .A2(new_n1513_), .A3(new_n2012_), .ZN(new_n2013_));
  OAI21_X1   g1628(.A1(new_n2008_), .A2(new_n2011_), .B(new_n2013_), .ZN(new_n2014_));
  NOR2_X1    g1629(.A1(new_n1029_), .A2(\req[96] ), .ZN(new_n2015_));
  NOR2_X1    g1630(.A1(new_n2015_), .A2(\priority[97] ), .ZN(new_n2016_));
  NAND4_X1   g1631(.A1(new_n1520_), .A2(new_n668_), .A3(new_n2016_), .A4(new_n680_), .ZN(new_n2017_));
  INV_X1     g1632(.I(new_n2017_), .ZN(new_n2018_));
  OAI21_X1   g1633(.A1(new_n699_), .A2(\req[100] ), .B(new_n701_), .ZN(new_n2019_));
  NOR3_X1    g1634(.A1(new_n690_), .A2(new_n1527_), .A3(new_n2019_), .ZN(new_n2020_));
  INV_X1     g1635(.I(new_n2020_), .ZN(new_n2021_));
  AOI21_X1   g1636(.A1(new_n2014_), .A2(new_n2018_), .B(new_n2021_), .ZN(new_n2022_));
  NOR2_X1    g1637(.A1(new_n1054_), .A2(\req[105] ), .ZN(new_n2023_));
  NOR2_X1    g1638(.A1(new_n2023_), .A2(\priority[106] ), .ZN(new_n2024_));
  NAND4_X1   g1639(.A1(new_n1533_), .A2(new_n696_), .A3(new_n2024_), .A4(new_n707_), .ZN(new_n2025_));
  OAI21_X1   g1640(.A1(new_n727_), .A2(\req[109] ), .B(new_n729_), .ZN(new_n2026_));
  NOR3_X1    g1641(.A1(new_n717_), .A2(new_n1539_), .A3(new_n2026_), .ZN(new_n2027_));
  OAI21_X1   g1642(.A1(new_n2022_), .A2(new_n2025_), .B(new_n2027_), .ZN(new_n2028_));
  NOR2_X1    g1643(.A1(new_n1079_), .A2(\req[114] ), .ZN(new_n2029_));
  NOR2_X1    g1644(.A1(new_n2029_), .A2(\priority[115] ), .ZN(new_n2030_));
  NAND4_X1   g1645(.A1(new_n1546_), .A2(new_n724_), .A3(new_n2030_), .A4(new_n736_), .ZN(new_n2031_));
  INV_X1     g1646(.I(new_n2031_), .ZN(new_n2032_));
  OAI21_X1   g1647(.A1(new_n755_), .A2(\req[118] ), .B(new_n757_), .ZN(new_n2033_));
  NOR3_X1    g1648(.A1(new_n746_), .A2(new_n1553_), .A3(new_n2033_), .ZN(new_n2034_));
  INV_X1     g1649(.I(new_n2034_), .ZN(new_n2035_));
  AOI21_X1   g1650(.A1(new_n2028_), .A2(new_n2032_), .B(new_n2035_), .ZN(new_n2036_));
  NOR2_X1    g1651(.A1(new_n1104_), .A2(\req[123] ), .ZN(new_n2037_));
  NOR2_X1    g1652(.A1(new_n2037_), .A2(\priority[124] ), .ZN(new_n2038_));
  NAND4_X1   g1653(.A1(new_n1559_), .A2(new_n752_), .A3(new_n2038_), .A4(new_n763_), .ZN(new_n2039_));
  OAI21_X1   g1654(.A1(new_n777_), .A2(\req[127] ), .B(new_n1566_), .ZN(new_n2040_));
  NOR3_X1    g1655(.A1(new_n773_), .A2(new_n1564_), .A3(new_n2040_), .ZN(new_n2041_));
  OAI21_X1   g1656(.A1(new_n2036_), .A2(new_n2039_), .B(new_n2041_), .ZN(new_n2042_));
  NOR2_X1    g1657(.A1(new_n386_), .A2(\req[4] ), .ZN(new_n2043_));
  NOR3_X1    g1658(.A1(new_n2043_), .A2(\priority[5] ), .A3(\priority[6] ), .ZN(new_n2044_));
  NAND2_X1   g1659(.A1(new_n1129_), .A2(\priority[1] ), .ZN(new_n2045_));
  NAND3_X1   g1660(.A1(new_n2045_), .A2(new_n785_), .A3(new_n1138_), .ZN(new_n2046_));
  NOR2_X1    g1661(.A1(new_n791_), .A2(new_n1571_), .ZN(new_n2047_));
  NAND3_X1   g1662(.A1(new_n2044_), .A2(new_n2047_), .A3(new_n2046_), .ZN(new_n2048_));
  INV_X1     g1663(.I(new_n2048_), .ZN(new_n2049_));
  NOR2_X1    g1664(.A1(new_n781_), .A2(\req[5] ), .ZN(new_n2050_));
  NAND2_X1   g1665(.A1(new_n2050_), .A2(new_n401_), .ZN(new_n2051_));
  AOI21_X1   g1666(.A1(new_n2042_), .A2(new_n2049_), .B(new_n2051_), .ZN(\grant[6] ));
  OAI21_X1   g1667(.A1(new_n810_), .A2(\req[11] ), .B(new_n812_), .ZN(new_n2053_));
  AOI21_X1   g1668(.A1(new_n1143_), .A2(\priority[8] ), .B(\priority[9] ), .ZN(new_n2054_));
  NOR4_X1    g1669(.A1(new_n1580_), .A2(new_n801_), .A3(new_n2053_), .A4(new_n2054_), .ZN(new_n2055_));
  AOI21_X1   g1670(.A1(new_n817_), .A2(\priority[16] ), .B(\priority[17] ), .ZN(new_n2056_));
  NAND4_X1   g1671(.A1(new_n1586_), .A2(new_n807_), .A3(new_n431_), .A4(new_n2056_), .ZN(new_n2057_));
  OAI21_X1   g1672(.A1(new_n835_), .A2(\req[20] ), .B(new_n837_), .ZN(new_n2058_));
  NOR3_X1    g1673(.A1(new_n826_), .A2(new_n1592_), .A3(new_n2058_), .ZN(new_n2059_));
  OAI21_X1   g1674(.A1(new_n2057_), .A2(new_n2055_), .B(new_n2059_), .ZN(new_n2060_));
  AOI21_X1   g1675(.A1(new_n843_), .A2(\priority[25] ), .B(\priority[26] ), .ZN(new_n2061_));
  NAND4_X1   g1676(.A1(new_n1599_), .A2(new_n832_), .A3(new_n460_), .A4(new_n2061_), .ZN(new_n2062_));
  INV_X1     g1677(.I(new_n2062_), .ZN(new_n2063_));
  OAI21_X1   g1678(.A1(new_n860_), .A2(\req[29] ), .B(new_n862_), .ZN(new_n2064_));
  NOR3_X1    g1679(.A1(new_n852_), .A2(new_n1606_), .A3(new_n2064_), .ZN(new_n2065_));
  INV_X1     g1680(.I(new_n2065_), .ZN(new_n2066_));
  AOI21_X1   g1681(.A1(new_n2060_), .A2(new_n2063_), .B(new_n2066_), .ZN(new_n2067_));
  AOI21_X1   g1682(.A1(new_n867_), .A2(\priority[34] ), .B(\priority[35] ), .ZN(new_n2068_));
  NAND4_X1   g1683(.A1(new_n1612_), .A2(new_n857_), .A3(new_n487_), .A4(new_n2068_), .ZN(new_n2069_));
  OAI21_X1   g1684(.A1(new_n885_), .A2(\req[38] ), .B(new_n887_), .ZN(new_n2070_));
  NOR3_X1    g1685(.A1(new_n876_), .A2(new_n1618_), .A3(new_n2070_), .ZN(new_n2071_));
  OAI21_X1   g1686(.A1(new_n2067_), .A2(new_n2069_), .B(new_n2071_), .ZN(new_n2072_));
  AOI21_X1   g1687(.A1(new_n893_), .A2(\priority[43] ), .B(\priority[44] ), .ZN(new_n2073_));
  NAND4_X1   g1688(.A1(new_n1625_), .A2(new_n882_), .A3(new_n516_), .A4(new_n2073_), .ZN(new_n2074_));
  INV_X1     g1689(.I(new_n2074_), .ZN(new_n2075_));
  OAI21_X1   g1690(.A1(new_n910_), .A2(\req[47] ), .B(new_n912_), .ZN(new_n2076_));
  NOR3_X1    g1691(.A1(new_n902_), .A2(new_n1632_), .A3(new_n2076_), .ZN(new_n2077_));
  INV_X1     g1692(.I(new_n2077_), .ZN(new_n2078_));
  AOI21_X1   g1693(.A1(new_n2072_), .A2(new_n2075_), .B(new_n2078_), .ZN(new_n2079_));
  AOI21_X1   g1694(.A1(new_n917_), .A2(\priority[52] ), .B(\priority[53] ), .ZN(new_n2080_));
  NAND4_X1   g1695(.A1(new_n1638_), .A2(new_n907_), .A3(new_n543_), .A4(new_n2080_), .ZN(new_n2081_));
  OAI21_X1   g1696(.A1(new_n935_), .A2(\req[56] ), .B(new_n937_), .ZN(new_n2082_));
  NOR3_X1    g1697(.A1(new_n926_), .A2(new_n1644_), .A3(new_n2082_), .ZN(new_n2083_));
  OAI21_X1   g1698(.A1(new_n2079_), .A2(new_n2081_), .B(new_n2083_), .ZN(new_n2084_));
  AOI21_X1   g1699(.A1(new_n943_), .A2(\priority[61] ), .B(\priority[62] ), .ZN(new_n2085_));
  NAND4_X1   g1700(.A1(new_n1651_), .A2(new_n932_), .A3(new_n572_), .A4(new_n2085_), .ZN(new_n2086_));
  INV_X1     g1701(.I(new_n2086_), .ZN(new_n2087_));
  OAI21_X1   g1702(.A1(new_n960_), .A2(\req[65] ), .B(new_n962_), .ZN(new_n2088_));
  NOR3_X1    g1703(.A1(new_n952_), .A2(new_n1658_), .A3(new_n2088_), .ZN(new_n2089_));
  INV_X1     g1704(.I(new_n2089_), .ZN(new_n2090_));
  AOI21_X1   g1705(.A1(new_n2084_), .A2(new_n2087_), .B(new_n2090_), .ZN(new_n2091_));
  AOI21_X1   g1706(.A1(new_n967_), .A2(\priority[70] ), .B(\priority[71] ), .ZN(new_n2092_));
  NAND4_X1   g1707(.A1(new_n1664_), .A2(new_n957_), .A3(new_n599_), .A4(new_n2092_), .ZN(new_n2093_));
  OAI21_X1   g1708(.A1(new_n985_), .A2(\req[74] ), .B(new_n987_), .ZN(new_n2094_));
  NOR3_X1    g1709(.A1(new_n976_), .A2(new_n1670_), .A3(new_n2094_), .ZN(new_n2095_));
  OAI21_X1   g1710(.A1(new_n2091_), .A2(new_n2093_), .B(new_n2095_), .ZN(new_n2096_));
  AOI21_X1   g1711(.A1(new_n993_), .A2(\priority[79] ), .B(\priority[80] ), .ZN(new_n2097_));
  NAND4_X1   g1712(.A1(new_n1677_), .A2(new_n982_), .A3(new_n628_), .A4(new_n2097_), .ZN(new_n2098_));
  INV_X1     g1713(.I(new_n2098_), .ZN(new_n2099_));
  OAI21_X1   g1714(.A1(new_n1010_), .A2(\req[83] ), .B(new_n1012_), .ZN(new_n2100_));
  NOR3_X1    g1715(.A1(new_n1002_), .A2(new_n1684_), .A3(new_n2100_), .ZN(new_n2101_));
  INV_X1     g1716(.I(new_n2101_), .ZN(new_n2102_));
  AOI21_X1   g1717(.A1(new_n2096_), .A2(new_n2099_), .B(new_n2102_), .ZN(new_n2103_));
  AOI21_X1   g1718(.A1(new_n1017_), .A2(\priority[88] ), .B(\priority[89] ), .ZN(new_n2104_));
  NAND4_X1   g1719(.A1(new_n1690_), .A2(new_n1007_), .A3(new_n655_), .A4(new_n2104_), .ZN(new_n2105_));
  OAI21_X1   g1720(.A1(new_n1035_), .A2(\req[92] ), .B(new_n1037_), .ZN(new_n2106_));
  NOR3_X1    g1721(.A1(new_n1026_), .A2(new_n1696_), .A3(new_n2106_), .ZN(new_n2107_));
  OAI21_X1   g1722(.A1(new_n2103_), .A2(new_n2105_), .B(new_n2107_), .ZN(new_n2108_));
  AOI21_X1   g1723(.A1(new_n1043_), .A2(\priority[97] ), .B(\priority[98] ), .ZN(new_n2109_));
  NAND4_X1   g1724(.A1(new_n1703_), .A2(new_n1032_), .A3(new_n684_), .A4(new_n2109_), .ZN(new_n2110_));
  INV_X1     g1725(.I(new_n2110_), .ZN(new_n2111_));
  OAI21_X1   g1726(.A1(new_n1060_), .A2(\req[101] ), .B(new_n1062_), .ZN(new_n2112_));
  NOR3_X1    g1727(.A1(new_n1052_), .A2(new_n1710_), .A3(new_n2112_), .ZN(new_n2113_));
  INV_X1     g1728(.I(new_n2113_), .ZN(new_n2114_));
  AOI21_X1   g1729(.A1(new_n2108_), .A2(new_n2111_), .B(new_n2114_), .ZN(new_n2115_));
  AOI21_X1   g1730(.A1(new_n1067_), .A2(\priority[106] ), .B(\priority[107] ), .ZN(new_n2116_));
  NAND4_X1   g1731(.A1(new_n1716_), .A2(new_n1057_), .A3(new_n711_), .A4(new_n2116_), .ZN(new_n2117_));
  OAI21_X1   g1732(.A1(new_n1085_), .A2(\req[110] ), .B(new_n1087_), .ZN(new_n2118_));
  NOR3_X1    g1733(.A1(new_n1076_), .A2(new_n1722_), .A3(new_n2118_), .ZN(new_n2119_));
  OAI21_X1   g1734(.A1(new_n2115_), .A2(new_n2117_), .B(new_n2119_), .ZN(new_n2120_));
  AOI21_X1   g1735(.A1(new_n1093_), .A2(\priority[115] ), .B(\priority[116] ), .ZN(new_n2121_));
  NAND4_X1   g1736(.A1(new_n1729_), .A2(new_n1082_), .A3(new_n740_), .A4(new_n2121_), .ZN(new_n2122_));
  INV_X1     g1737(.I(new_n2122_), .ZN(new_n2123_));
  OAI21_X1   g1738(.A1(new_n1110_), .A2(\req[119] ), .B(new_n1112_), .ZN(new_n2124_));
  NOR3_X1    g1739(.A1(new_n1102_), .A2(new_n1736_), .A3(new_n2124_), .ZN(new_n2125_));
  INV_X1     g1740(.I(new_n2125_), .ZN(new_n2126_));
  AOI21_X1   g1741(.A1(new_n2120_), .A2(new_n2123_), .B(new_n2126_), .ZN(new_n2127_));
  AOI21_X1   g1742(.A1(new_n1117_), .A2(\priority[124] ), .B(\priority[125] ), .ZN(new_n2128_));
  NAND4_X1   g1743(.A1(new_n1742_), .A2(new_n1107_), .A3(new_n767_), .A4(new_n2128_), .ZN(new_n2129_));
  NOR2_X1    g1744(.A1(\req[1] ), .A2(\req[2] ), .ZN(new_n2130_));
  OAI21_X1   g1745(.A1(new_n391_), .A2(\req[0] ), .B(new_n2130_), .ZN(new_n2131_));
  NOR3_X1    g1746(.A1(new_n1126_), .A2(new_n1747_), .A3(new_n2131_), .ZN(new_n2132_));
  OAI21_X1   g1747(.A1(new_n2127_), .A2(new_n2129_), .B(new_n2132_), .ZN(new_n2133_));
  NOR2_X1    g1748(.A1(new_n387_), .A2(\req[5] ), .ZN(new_n2134_));
  NOR3_X1    g1749(.A1(new_n2134_), .A2(\priority[6] ), .A3(\priority[7] ), .ZN(new_n2135_));
  NAND2_X1   g1750(.A1(new_n1387_), .A2(\priority[2] ), .ZN(new_n2136_));
  NAND3_X1   g1751(.A1(new_n2136_), .A2(new_n1138_), .A3(new_n386_), .ZN(new_n2137_));
  NOR3_X1    g1752(.A1(new_n1752_), .A2(\req[4] ), .A3(\req[5] ), .ZN(new_n2138_));
  NAND3_X1   g1753(.A1(new_n2135_), .A2(new_n2138_), .A3(new_n2137_), .ZN(new_n2139_));
  INV_X1     g1754(.I(new_n2139_), .ZN(new_n2140_));
  NOR2_X1    g1755(.A1(new_n399_), .A2(\req[6] ), .ZN(new_n2141_));
  NAND2_X1   g1756(.A1(new_n2141_), .A2(new_n793_), .ZN(new_n2142_));
  AOI21_X1   g1757(.A1(new_n2133_), .A2(new_n2140_), .B(new_n2142_), .ZN(\grant[7] ));
  NOR2_X1    g1758(.A1(\req[13] ), .A2(\req[14] ), .ZN(new_n2144_));
  OAI21_X1   g1759(.A1(new_n412_), .A2(\req[12] ), .B(new_n2144_), .ZN(new_n2145_));
  OAI21_X1   g1760(.A1(new_n405_), .A2(\priority[10] ), .B(new_n1758_), .ZN(new_n2146_));
  NOR3_X1    g1761(.A1(new_n2146_), .A2(new_n1763_), .A3(new_n2145_), .ZN(new_n2147_));
  AOI21_X1   g1762(.A1(new_n1160_), .A2(\priority[17] ), .B(\priority[18] ), .ZN(new_n2148_));
  NAND4_X1   g1763(.A1(new_n1769_), .A2(new_n1153_), .A3(new_n820_), .A4(new_n2148_), .ZN(new_n2149_));
  NOR2_X1    g1764(.A1(\req[22] ), .A2(\req[23] ), .ZN(new_n2150_));
  OAI21_X1   g1765(.A1(new_n440_), .A2(\req[21] ), .B(new_n2150_), .ZN(new_n2151_));
  NOR3_X1    g1766(.A1(new_n1166_), .A2(new_n1776_), .A3(new_n2151_), .ZN(new_n2152_));
  OAI21_X1   g1767(.A1(new_n2149_), .A2(new_n2147_), .B(new_n2152_), .ZN(new_n2153_));
  AOI21_X1   g1768(.A1(new_n1179_), .A2(\priority[26] ), .B(\priority[27] ), .ZN(new_n2154_));
  NAND4_X1   g1769(.A1(new_n1783_), .A2(new_n1171_), .A3(new_n846_), .A4(new_n2154_), .ZN(new_n2155_));
  INV_X1     g1770(.I(new_n2155_), .ZN(new_n2156_));
  NOR2_X1    g1771(.A1(\req[31] ), .A2(\req[32] ), .ZN(new_n2157_));
  OAI21_X1   g1772(.A1(new_n468_), .A2(\req[30] ), .B(new_n2157_), .ZN(new_n2158_));
  NOR3_X1    g1773(.A1(new_n1185_), .A2(new_n1791_), .A3(new_n2158_), .ZN(new_n2159_));
  INV_X1     g1774(.I(new_n2159_), .ZN(new_n2160_));
  AOI21_X1   g1775(.A1(new_n2153_), .A2(new_n2156_), .B(new_n2160_), .ZN(new_n2161_));
  AOI21_X1   g1776(.A1(new_n1196_), .A2(\priority[35] ), .B(\priority[36] ), .ZN(new_n2162_));
  NAND4_X1   g1777(.A1(new_n1797_), .A2(new_n1189_), .A3(new_n870_), .A4(new_n2162_), .ZN(new_n2163_));
  NOR2_X1    g1778(.A1(\req[40] ), .A2(\req[41] ), .ZN(new_n2164_));
  OAI21_X1   g1779(.A1(new_n496_), .A2(\req[39] ), .B(new_n2164_), .ZN(new_n2165_));
  NOR3_X1    g1780(.A1(new_n1202_), .A2(new_n1804_), .A3(new_n2165_), .ZN(new_n2166_));
  OAI21_X1   g1781(.A1(new_n2161_), .A2(new_n2163_), .B(new_n2166_), .ZN(new_n2167_));
  AOI21_X1   g1782(.A1(new_n1215_), .A2(\priority[44] ), .B(\priority[45] ), .ZN(new_n2168_));
  NAND4_X1   g1783(.A1(new_n1811_), .A2(new_n1207_), .A3(new_n896_), .A4(new_n2168_), .ZN(new_n2169_));
  INV_X1     g1784(.I(new_n2169_), .ZN(new_n2170_));
  NOR2_X1    g1785(.A1(\req[49] ), .A2(\req[50] ), .ZN(new_n2171_));
  OAI21_X1   g1786(.A1(new_n524_), .A2(\req[48] ), .B(new_n2171_), .ZN(new_n2172_));
  NOR3_X1    g1787(.A1(new_n1221_), .A2(new_n1819_), .A3(new_n2172_), .ZN(new_n2173_));
  INV_X1     g1788(.I(new_n2173_), .ZN(new_n2174_));
  AOI21_X1   g1789(.A1(new_n2167_), .A2(new_n2170_), .B(new_n2174_), .ZN(new_n2175_));
  AOI21_X1   g1790(.A1(new_n1232_), .A2(\priority[53] ), .B(\priority[54] ), .ZN(new_n2176_));
  NAND4_X1   g1791(.A1(new_n1825_), .A2(new_n1225_), .A3(new_n920_), .A4(new_n2176_), .ZN(new_n2177_));
  NOR2_X1    g1792(.A1(\req[58] ), .A2(\req[59] ), .ZN(new_n2178_));
  OAI21_X1   g1793(.A1(new_n552_), .A2(\req[57] ), .B(new_n2178_), .ZN(new_n2179_));
  NOR3_X1    g1794(.A1(new_n1238_), .A2(new_n1832_), .A3(new_n2179_), .ZN(new_n2180_));
  OAI21_X1   g1795(.A1(new_n2175_), .A2(new_n2177_), .B(new_n2180_), .ZN(new_n2181_));
  AOI21_X1   g1796(.A1(new_n1251_), .A2(\priority[62] ), .B(\priority[63] ), .ZN(new_n2182_));
  NAND4_X1   g1797(.A1(new_n1839_), .A2(new_n1243_), .A3(new_n946_), .A4(new_n2182_), .ZN(new_n2183_));
  INV_X1     g1798(.I(new_n2183_), .ZN(new_n2184_));
  NOR2_X1    g1799(.A1(\req[67] ), .A2(\req[68] ), .ZN(new_n2185_));
  OAI21_X1   g1800(.A1(new_n580_), .A2(\req[66] ), .B(new_n2185_), .ZN(new_n2186_));
  NOR3_X1    g1801(.A1(new_n1257_), .A2(new_n1847_), .A3(new_n2186_), .ZN(new_n2187_));
  INV_X1     g1802(.I(new_n2187_), .ZN(new_n2188_));
  AOI21_X1   g1803(.A1(new_n2181_), .A2(new_n2184_), .B(new_n2188_), .ZN(new_n2189_));
  AOI21_X1   g1804(.A1(new_n1268_), .A2(\priority[71] ), .B(\priority[72] ), .ZN(new_n2190_));
  NAND4_X1   g1805(.A1(new_n1853_), .A2(new_n1261_), .A3(new_n970_), .A4(new_n2190_), .ZN(new_n2191_));
  NOR2_X1    g1806(.A1(\req[76] ), .A2(\req[77] ), .ZN(new_n2192_));
  OAI21_X1   g1807(.A1(new_n608_), .A2(\req[75] ), .B(new_n2192_), .ZN(new_n2193_));
  NOR3_X1    g1808(.A1(new_n1274_), .A2(new_n1860_), .A3(new_n2193_), .ZN(new_n2194_));
  OAI21_X1   g1809(.A1(new_n2189_), .A2(new_n2191_), .B(new_n2194_), .ZN(new_n2195_));
  AOI21_X1   g1810(.A1(new_n1287_), .A2(\priority[80] ), .B(\priority[81] ), .ZN(new_n2196_));
  NAND4_X1   g1811(.A1(new_n1867_), .A2(new_n1279_), .A3(new_n996_), .A4(new_n2196_), .ZN(new_n2197_));
  INV_X1     g1812(.I(new_n2197_), .ZN(new_n2198_));
  NOR2_X1    g1813(.A1(\req[85] ), .A2(\req[86] ), .ZN(new_n2199_));
  OAI21_X1   g1814(.A1(new_n636_), .A2(\req[84] ), .B(new_n2199_), .ZN(new_n2200_));
  NOR3_X1    g1815(.A1(new_n1293_), .A2(new_n1875_), .A3(new_n2200_), .ZN(new_n2201_));
  INV_X1     g1816(.I(new_n2201_), .ZN(new_n2202_));
  AOI21_X1   g1817(.A1(new_n2195_), .A2(new_n2198_), .B(new_n2202_), .ZN(new_n2203_));
  AOI21_X1   g1818(.A1(new_n1304_), .A2(\priority[89] ), .B(\priority[90] ), .ZN(new_n2204_));
  NAND4_X1   g1819(.A1(new_n1881_), .A2(new_n1297_), .A3(new_n1020_), .A4(new_n2204_), .ZN(new_n2205_));
  NOR2_X1    g1820(.A1(\req[94] ), .A2(\req[95] ), .ZN(new_n2206_));
  OAI21_X1   g1821(.A1(new_n664_), .A2(\req[93] ), .B(new_n2206_), .ZN(new_n2207_));
  NOR3_X1    g1822(.A1(new_n1310_), .A2(new_n1888_), .A3(new_n2207_), .ZN(new_n2208_));
  OAI21_X1   g1823(.A1(new_n2203_), .A2(new_n2205_), .B(new_n2208_), .ZN(new_n2209_));
  AOI21_X1   g1824(.A1(new_n1323_), .A2(\priority[98] ), .B(\priority[99] ), .ZN(new_n2210_));
  NAND4_X1   g1825(.A1(new_n1895_), .A2(new_n1315_), .A3(new_n1046_), .A4(new_n2210_), .ZN(new_n2211_));
  INV_X1     g1826(.I(new_n2211_), .ZN(new_n2212_));
  NOR2_X1    g1827(.A1(\req[103] ), .A2(\req[104] ), .ZN(new_n2213_));
  OAI21_X1   g1828(.A1(new_n692_), .A2(\req[102] ), .B(new_n2213_), .ZN(new_n2214_));
  NOR3_X1    g1829(.A1(new_n1329_), .A2(new_n1903_), .A3(new_n2214_), .ZN(new_n2215_));
  INV_X1     g1830(.I(new_n2215_), .ZN(new_n2216_));
  AOI21_X1   g1831(.A1(new_n2209_), .A2(new_n2212_), .B(new_n2216_), .ZN(new_n2217_));
  AOI21_X1   g1832(.A1(new_n1340_), .A2(\priority[107] ), .B(\priority[108] ), .ZN(new_n2218_));
  NAND4_X1   g1833(.A1(new_n1909_), .A2(new_n1333_), .A3(new_n1070_), .A4(new_n2218_), .ZN(new_n2219_));
  NOR2_X1    g1834(.A1(\req[112] ), .A2(\req[113] ), .ZN(new_n2220_));
  OAI21_X1   g1835(.A1(new_n720_), .A2(\req[111] ), .B(new_n2220_), .ZN(new_n2221_));
  NOR3_X1    g1836(.A1(new_n1346_), .A2(new_n1916_), .A3(new_n2221_), .ZN(new_n2222_));
  OAI21_X1   g1837(.A1(new_n2217_), .A2(new_n2219_), .B(new_n2222_), .ZN(new_n2223_));
  AOI21_X1   g1838(.A1(new_n1359_), .A2(\priority[116] ), .B(\priority[117] ), .ZN(new_n2224_));
  NAND4_X1   g1839(.A1(new_n1923_), .A2(new_n1351_), .A3(new_n1096_), .A4(new_n2224_), .ZN(new_n2225_));
  INV_X1     g1840(.I(new_n2225_), .ZN(new_n2226_));
  NOR2_X1    g1841(.A1(\req[121] ), .A2(\req[122] ), .ZN(new_n2227_));
  OAI21_X1   g1842(.A1(new_n748_), .A2(\req[120] ), .B(new_n2227_), .ZN(new_n2228_));
  NOR3_X1    g1843(.A1(new_n1365_), .A2(new_n1931_), .A3(new_n2228_), .ZN(new_n2229_));
  INV_X1     g1844(.I(new_n2229_), .ZN(new_n2230_));
  AOI21_X1   g1845(.A1(new_n2223_), .A2(new_n2226_), .B(new_n2230_), .ZN(new_n2231_));
  AOI21_X1   g1846(.A1(new_n1376_), .A2(\priority[125] ), .B(\priority[126] ), .ZN(new_n2232_));
  NAND4_X1   g1847(.A1(new_n1937_), .A2(new_n1369_), .A3(new_n1120_), .A4(new_n2232_), .ZN(new_n2233_));
  OAI21_X1   g1848(.A1(new_n785_), .A2(\req[1] ), .B(new_n396_), .ZN(new_n2234_));
  NOR3_X1    g1849(.A1(new_n1384_), .A2(new_n1943_), .A3(new_n2234_), .ZN(new_n2235_));
  OAI21_X1   g1850(.A1(new_n2231_), .A2(new_n2233_), .B(new_n2235_), .ZN(new_n2236_));
  NOR2_X1    g1851(.A1(new_n1391_), .A2(new_n1947_), .ZN(new_n2237_));
  NOR3_X1    g1852(.A1(new_n1755_), .A2(\priority[7] ), .A3(\priority[8] ), .ZN(new_n2238_));
  NAND3_X1   g1853(.A1(new_n2237_), .A2(new_n2238_), .A3(new_n390_), .ZN(new_n2239_));
  INV_X1     g1854(.I(new_n2239_), .ZN(new_n2240_));
  NAND2_X1   g1855(.A1(new_n407_), .A2(new_n1143_), .ZN(new_n2241_));
  AOI21_X1   g1856(.A1(new_n2236_), .A2(new_n2240_), .B(new_n2241_), .ZN(\grant[8] ));
  INV_X1     g1857(.I(new_n747_), .ZN(new_n2243_));
  INV_X1     g1858(.I(new_n760_), .ZN(new_n2244_));
  INV_X1     g1859(.I(new_n691_), .ZN(new_n2245_));
  INV_X1     g1860(.I(new_n704_), .ZN(new_n2246_));
  INV_X1     g1861(.I(new_n635_), .ZN(new_n2247_));
  INV_X1     g1862(.I(new_n648_), .ZN(new_n2248_));
  INV_X1     g1863(.I(new_n579_), .ZN(new_n2249_));
  INV_X1     g1864(.I(new_n592_), .ZN(new_n2250_));
  INV_X1     g1865(.I(new_n523_), .ZN(new_n2251_));
  INV_X1     g1866(.I(new_n536_), .ZN(new_n2252_));
  INV_X1     g1867(.I(new_n467_), .ZN(new_n2253_));
  INV_X1     g1868(.I(new_n480_), .ZN(new_n2254_));
  AOI21_X1   g1869(.A1(new_n1578_), .A2(\priority[10] ), .B(\priority[11] ), .ZN(new_n2255_));
  NOR4_X1    g1870(.A1(new_n416_), .A2(new_n418_), .A3(new_n422_), .A4(new_n2255_), .ZN(new_n2256_));
  OAI21_X1   g1871(.A1(new_n438_), .A2(new_n2256_), .B(new_n452_), .ZN(new_n2257_));
  AOI21_X1   g1872(.A1(new_n2257_), .A2(new_n2253_), .B(new_n2254_), .ZN(new_n2258_));
  OAI21_X1   g1873(.A1(new_n2258_), .A2(new_n494_), .B(new_n508_), .ZN(new_n2259_));
  AOI21_X1   g1874(.A1(new_n2259_), .A2(new_n2251_), .B(new_n2252_), .ZN(new_n2260_));
  OAI21_X1   g1875(.A1(new_n2260_), .A2(new_n550_), .B(new_n564_), .ZN(new_n2261_));
  AOI21_X1   g1876(.A1(new_n2261_), .A2(new_n2249_), .B(new_n2250_), .ZN(new_n2262_));
  OAI21_X1   g1877(.A1(new_n2262_), .A2(new_n606_), .B(new_n620_), .ZN(new_n2263_));
  AOI21_X1   g1878(.A1(new_n2263_), .A2(new_n2247_), .B(new_n2248_), .ZN(new_n2264_));
  OAI21_X1   g1879(.A1(new_n2264_), .A2(new_n662_), .B(new_n676_), .ZN(new_n2265_));
  AOI21_X1   g1880(.A1(new_n2265_), .A2(new_n2245_), .B(new_n2246_), .ZN(new_n2266_));
  OAI21_X1   g1881(.A1(new_n2266_), .A2(new_n718_), .B(new_n732_), .ZN(new_n2267_));
  AOI21_X1   g1882(.A1(new_n2267_), .A2(new_n2243_), .B(new_n2244_), .ZN(new_n2268_));
  OAI21_X1   g1883(.A1(new_n1138_), .A2(\req[2] ), .B(new_n790_), .ZN(new_n2269_));
  NOR3_X1    g1884(.A1(new_n1568_), .A2(new_n2046_), .A3(new_n2269_), .ZN(new_n2270_));
  OAI21_X1   g1885(.A1(new_n2268_), .A2(new_n774_), .B(new_n2270_), .ZN(new_n2271_));
  NOR2_X1    g1886(.A1(new_n1574_), .A2(new_n2050_), .ZN(new_n2272_));
  NOR2_X1    g1887(.A1(new_n399_), .A2(\req[7] ), .ZN(new_n2273_));
  NOR3_X1    g1888(.A1(new_n2273_), .A2(\priority[8] ), .A3(\priority[9] ), .ZN(new_n2274_));
  NAND3_X1   g1889(.A1(new_n2272_), .A2(new_n2274_), .A3(new_n784_), .ZN(new_n2275_));
  INV_X1     g1890(.I(new_n2275_), .ZN(new_n2276_));
  NAND2_X1   g1891(.A1(new_n799_), .A2(new_n1395_), .ZN(new_n2277_));
  AOI21_X1   g1892(.A1(new_n2271_), .A2(new_n2276_), .B(new_n2277_), .ZN(\grant[9] ));
  INV_X1     g1893(.I(new_n1103_), .ZN(new_n2279_));
  INV_X1     g1894(.I(new_n1115_), .ZN(new_n2280_));
  INV_X1     g1895(.I(new_n1053_), .ZN(new_n2281_));
  INV_X1     g1896(.I(new_n1065_), .ZN(new_n2282_));
  INV_X1     g1897(.I(new_n1003_), .ZN(new_n2283_));
  INV_X1     g1898(.I(new_n1015_), .ZN(new_n2284_));
  INV_X1     g1899(.I(new_n953_), .ZN(new_n2285_));
  INV_X1     g1900(.I(new_n965_), .ZN(new_n2286_));
  INV_X1     g1901(.I(new_n903_), .ZN(new_n2287_));
  INV_X1     g1902(.I(new_n915_), .ZN(new_n2288_));
  INV_X1     g1903(.I(new_n853_), .ZN(new_n2289_));
  INV_X1     g1904(.I(new_n865_), .ZN(new_n2290_));
  AOI21_X1   g1905(.A1(new_n1761_), .A2(\priority[11] ), .B(\priority[12] ), .ZN(new_n2291_));
  NOR4_X1    g1906(.A1(new_n807_), .A2(new_n809_), .A3(new_n813_), .A4(new_n2291_), .ZN(new_n2292_));
  OAI21_X1   g1907(.A1(new_n827_), .A2(new_n2292_), .B(new_n840_), .ZN(new_n2293_));
  AOI21_X1   g1908(.A1(new_n2293_), .A2(new_n2289_), .B(new_n2290_), .ZN(new_n2294_));
  OAI21_X1   g1909(.A1(new_n2294_), .A2(new_n877_), .B(new_n890_), .ZN(new_n2295_));
  AOI21_X1   g1910(.A1(new_n2295_), .A2(new_n2287_), .B(new_n2288_), .ZN(new_n2296_));
  OAI21_X1   g1911(.A1(new_n2296_), .A2(new_n927_), .B(new_n940_), .ZN(new_n2297_));
  AOI21_X1   g1912(.A1(new_n2297_), .A2(new_n2285_), .B(new_n2286_), .ZN(new_n2298_));
  OAI21_X1   g1913(.A1(new_n2298_), .A2(new_n977_), .B(new_n990_), .ZN(new_n2299_));
  AOI21_X1   g1914(.A1(new_n2299_), .A2(new_n2283_), .B(new_n2284_), .ZN(new_n2300_));
  OAI21_X1   g1915(.A1(new_n2300_), .A2(new_n1027_), .B(new_n1040_), .ZN(new_n2301_));
  AOI21_X1   g1916(.A1(new_n2301_), .A2(new_n2281_), .B(new_n2282_), .ZN(new_n2302_));
  OAI21_X1   g1917(.A1(new_n2302_), .A2(new_n1077_), .B(new_n1090_), .ZN(new_n2303_));
  AOI21_X1   g1918(.A1(new_n2303_), .A2(new_n2279_), .B(new_n2280_), .ZN(new_n2304_));
  OAI21_X1   g1919(.A1(new_n386_), .A2(\req[3] ), .B(new_n1140_), .ZN(new_n2305_));
  NOR3_X1    g1920(.A1(new_n1749_), .A2(new_n2137_), .A3(new_n2305_), .ZN(new_n2306_));
  OAI21_X1   g1921(.A1(new_n2304_), .A2(new_n1127_), .B(new_n2306_), .ZN(new_n2307_));
  NOR2_X1    g1922(.A1(new_n1757_), .A2(new_n2141_), .ZN(new_n2308_));
  NOR2_X1    g1923(.A1(new_n400_), .A2(\req[8] ), .ZN(new_n2309_));
  NOR3_X1    g1924(.A1(new_n2309_), .A2(\priority[9] ), .A3(\priority[10] ), .ZN(new_n2310_));
  NAND3_X1   g1925(.A1(new_n2308_), .A2(new_n2310_), .A3(new_n1135_), .ZN(new_n2311_));
  INV_X1     g1926(.I(new_n2311_), .ZN(new_n2312_));
  NAND2_X1   g1927(.A1(new_n1148_), .A2(new_n1578_), .ZN(new_n2313_));
  AOI21_X1   g1928(.A1(new_n2307_), .A2(new_n2312_), .B(new_n2313_), .ZN(\grant[10] ));
  INV_X1     g1929(.I(new_n411_), .ZN(new_n2315_));
  INV_X1     g1930(.I(new_n1366_), .ZN(new_n2316_));
  INV_X1     g1931(.I(new_n1374_), .ZN(new_n2317_));
  INV_X1     g1932(.I(new_n1330_), .ZN(new_n2318_));
  INV_X1     g1933(.I(new_n1338_), .ZN(new_n2319_));
  INV_X1     g1934(.I(new_n1294_), .ZN(new_n2320_));
  INV_X1     g1935(.I(new_n1302_), .ZN(new_n2321_));
  INV_X1     g1936(.I(new_n1258_), .ZN(new_n2322_));
  INV_X1     g1937(.I(new_n1266_), .ZN(new_n2323_));
  INV_X1     g1938(.I(new_n1222_), .ZN(new_n2324_));
  INV_X1     g1939(.I(new_n1230_), .ZN(new_n2325_));
  INV_X1     g1940(.I(new_n1186_), .ZN(new_n2326_));
  INV_X1     g1941(.I(new_n1194_), .ZN(new_n2327_));
  OAI21_X1   g1942(.A1(new_n1398_), .A2(\priority[13] ), .B(new_n2144_), .ZN(new_n2328_));
  NOR3_X1    g1943(.A1(new_n2328_), .A2(new_n1153_), .A3(new_n1155_), .ZN(new_n2329_));
  OAI21_X1   g1944(.A1(new_n1167_), .A2(new_n2329_), .B(new_n1176_), .ZN(new_n2330_));
  AOI21_X1   g1945(.A1(new_n2330_), .A2(new_n2326_), .B(new_n2327_), .ZN(new_n2331_));
  OAI21_X1   g1946(.A1(new_n2331_), .A2(new_n1203_), .B(new_n1212_), .ZN(new_n2332_));
  AOI21_X1   g1947(.A1(new_n2332_), .A2(new_n2324_), .B(new_n2325_), .ZN(new_n2333_));
  OAI21_X1   g1948(.A1(new_n2333_), .A2(new_n1239_), .B(new_n1248_), .ZN(new_n2334_));
  AOI21_X1   g1949(.A1(new_n2334_), .A2(new_n2322_), .B(new_n2323_), .ZN(new_n2335_));
  OAI21_X1   g1950(.A1(new_n2335_), .A2(new_n1275_), .B(new_n1284_), .ZN(new_n2336_));
  AOI21_X1   g1951(.A1(new_n2336_), .A2(new_n2320_), .B(new_n2321_), .ZN(new_n2337_));
  OAI21_X1   g1952(.A1(new_n2337_), .A2(new_n1311_), .B(new_n1320_), .ZN(new_n2338_));
  AOI21_X1   g1953(.A1(new_n2338_), .A2(new_n2318_), .B(new_n2319_), .ZN(new_n2339_));
  OAI21_X1   g1954(.A1(new_n2339_), .A2(new_n1347_), .B(new_n1356_), .ZN(new_n2340_));
  AOI21_X1   g1955(.A1(new_n2340_), .A2(new_n2316_), .B(new_n2317_), .ZN(new_n2341_));
  NOR3_X1    g1956(.A1(new_n1944_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n2342_));
  OAI21_X1   g1957(.A1(new_n2341_), .A2(new_n1385_), .B(new_n2342_), .ZN(new_n2343_));
  NAND2_X1   g1958(.A1(new_n420_), .A2(new_n1761_), .ZN(new_n2344_));
  AOI21_X1   g1959(.A1(new_n2343_), .A2(new_n2315_), .B(new_n2344_), .ZN(\grant[11] ));
  INV_X1     g1960(.I(new_n803_), .ZN(new_n2346_));
  INV_X1     g1961(.I(new_n1556_), .ZN(new_n2347_));
  INV_X1     g1962(.I(new_n1561_), .ZN(new_n2348_));
  INV_X1     g1963(.I(new_n1530_), .ZN(new_n2349_));
  INV_X1     g1964(.I(new_n1535_), .ZN(new_n2350_));
  INV_X1     g1965(.I(new_n1504_), .ZN(new_n2351_));
  INV_X1     g1966(.I(new_n1509_), .ZN(new_n2352_));
  INV_X1     g1967(.I(new_n1478_), .ZN(new_n2353_));
  INV_X1     g1968(.I(new_n1483_), .ZN(new_n2354_));
  INV_X1     g1969(.I(new_n1452_), .ZN(new_n2355_));
  INV_X1     g1970(.I(new_n1457_), .ZN(new_n2356_));
  INV_X1     g1971(.I(new_n1426_), .ZN(new_n2357_));
  INV_X1     g1972(.I(new_n1431_), .ZN(new_n2358_));
  AOI21_X1   g1973(.A1(new_n805_), .A2(\priority[13] ), .B(\priority[14] ), .ZN(new_n2359_));
  NOR4_X1    g1974(.A1(new_n430_), .A2(new_n1402_), .A3(new_n1404_), .A4(new_n2359_), .ZN(new_n2360_));
  OAI21_X1   g1975(.A1(new_n1412_), .A2(new_n2360_), .B(new_n1418_), .ZN(new_n2361_));
  AOI21_X1   g1976(.A1(new_n2361_), .A2(new_n2357_), .B(new_n2358_), .ZN(new_n2362_));
  OAI21_X1   g1977(.A1(new_n2362_), .A2(new_n1438_), .B(new_n1444_), .ZN(new_n2363_));
  AOI21_X1   g1978(.A1(new_n2363_), .A2(new_n2355_), .B(new_n2356_), .ZN(new_n2364_));
  OAI21_X1   g1979(.A1(new_n2364_), .A2(new_n1464_), .B(new_n1470_), .ZN(new_n2365_));
  AOI21_X1   g1980(.A1(new_n2365_), .A2(new_n2353_), .B(new_n2354_), .ZN(new_n2366_));
  OAI21_X1   g1981(.A1(new_n2366_), .A2(new_n1490_), .B(new_n1496_), .ZN(new_n2367_));
  AOI21_X1   g1982(.A1(new_n2367_), .A2(new_n2351_), .B(new_n2352_), .ZN(new_n2368_));
  OAI21_X1   g1983(.A1(new_n2368_), .A2(new_n1516_), .B(new_n1522_), .ZN(new_n2369_));
  AOI21_X1   g1984(.A1(new_n2369_), .A2(new_n2349_), .B(new_n2350_), .ZN(new_n2370_));
  OAI21_X1   g1985(.A1(new_n2370_), .A2(new_n1542_), .B(new_n1548_), .ZN(new_n2371_));
  AOI21_X1   g1986(.A1(new_n2371_), .A2(new_n2347_), .B(new_n2348_), .ZN(new_n2372_));
  NOR3_X1    g1987(.A1(new_n2047_), .A2(new_n784_), .A3(new_n789_), .ZN(new_n2373_));
  OAI21_X1   g1988(.A1(new_n2372_), .A2(new_n1569_), .B(new_n2373_), .ZN(new_n2374_));
  NAND2_X1   g1989(.A1(new_n811_), .A2(new_n414_), .ZN(new_n2375_));
  AOI21_X1   g1990(.A1(new_n2374_), .A2(new_n2346_), .B(new_n2375_), .ZN(\grant[12] ));
  INV_X1     g1991(.I(new_n1150_), .ZN(new_n2377_));
  INV_X1     g1992(.I(new_n1739_), .ZN(new_n2378_));
  INV_X1     g1993(.I(new_n1744_), .ZN(new_n2379_));
  INV_X1     g1994(.I(new_n1713_), .ZN(new_n2380_));
  INV_X1     g1995(.I(new_n1718_), .ZN(new_n2381_));
  INV_X1     g1996(.I(new_n1687_), .ZN(new_n2382_));
  INV_X1     g1997(.I(new_n1692_), .ZN(new_n2383_));
  INV_X1     g1998(.I(new_n1661_), .ZN(new_n2384_));
  INV_X1     g1999(.I(new_n1666_), .ZN(new_n2385_));
  INV_X1     g2000(.I(new_n1635_), .ZN(new_n2386_));
  INV_X1     g2001(.I(new_n1640_), .ZN(new_n2387_));
  INV_X1     g2002(.I(new_n1609_), .ZN(new_n2388_));
  INV_X1     g2003(.I(new_n1614_), .ZN(new_n2389_));
  AOI21_X1   g2004(.A1(new_n1151_), .A2(\priority[14] ), .B(\priority[15] ), .ZN(new_n2390_));
  NOR4_X1    g2005(.A1(new_n819_), .A2(new_n1585_), .A3(new_n1587_), .A4(new_n2390_), .ZN(new_n2391_));
  OAI21_X1   g2006(.A1(new_n1595_), .A2(new_n2391_), .B(new_n1601_), .ZN(new_n2392_));
  AOI21_X1   g2007(.A1(new_n2392_), .A2(new_n2388_), .B(new_n2389_), .ZN(new_n2393_));
  OAI21_X1   g2008(.A1(new_n2393_), .A2(new_n1621_), .B(new_n1627_), .ZN(new_n2394_));
  AOI21_X1   g2009(.A1(new_n2394_), .A2(new_n2386_), .B(new_n2387_), .ZN(new_n2395_));
  OAI21_X1   g2010(.A1(new_n2395_), .A2(new_n1647_), .B(new_n1653_), .ZN(new_n2396_));
  AOI21_X1   g2011(.A1(new_n2396_), .A2(new_n2384_), .B(new_n2385_), .ZN(new_n2397_));
  OAI21_X1   g2012(.A1(new_n2397_), .A2(new_n1673_), .B(new_n1679_), .ZN(new_n2398_));
  AOI21_X1   g2013(.A1(new_n2398_), .A2(new_n2382_), .B(new_n2383_), .ZN(new_n2399_));
  OAI21_X1   g2014(.A1(new_n2399_), .A2(new_n1699_), .B(new_n1705_), .ZN(new_n2400_));
  AOI21_X1   g2015(.A1(new_n2400_), .A2(new_n2380_), .B(new_n2381_), .ZN(new_n2401_));
  OAI21_X1   g2016(.A1(new_n2401_), .A2(new_n1725_), .B(new_n1731_), .ZN(new_n2402_));
  AOI21_X1   g2017(.A1(new_n2402_), .A2(new_n2378_), .B(new_n2379_), .ZN(new_n2403_));
  NOR3_X1    g2018(.A1(new_n2138_), .A2(new_n1135_), .A3(new_n1137_), .ZN(new_n2404_));
  OAI21_X1   g2019(.A1(new_n2403_), .A2(new_n1750_), .B(new_n2404_), .ZN(new_n2405_));
  NAND2_X1   g2020(.A1(new_n1156_), .A2(new_n805_), .ZN(new_n2406_));
  AOI21_X1   g2021(.A1(new_n2405_), .A2(new_n2377_), .B(new_n2406_), .ZN(\grant[13] ));
  INV_X1     g2022(.I(new_n1400_), .ZN(new_n2408_));
  INV_X1     g2023(.I(new_n1934_), .ZN(new_n2409_));
  INV_X1     g2024(.I(new_n1939_), .ZN(new_n2410_));
  INV_X1     g2025(.I(new_n1906_), .ZN(new_n2411_));
  INV_X1     g2026(.I(new_n1912_), .ZN(new_n2412_));
  INV_X1     g2027(.I(new_n1878_), .ZN(new_n2413_));
  INV_X1     g2028(.I(new_n1884_), .ZN(new_n2414_));
  INV_X1     g2029(.I(new_n1850_), .ZN(new_n2415_));
  INV_X1     g2030(.I(new_n1856_), .ZN(new_n2416_));
  INV_X1     g2031(.I(new_n1822_), .ZN(new_n2417_));
  INV_X1     g2032(.I(new_n1828_), .ZN(new_n2418_));
  INV_X1     g2033(.I(new_n1794_), .ZN(new_n2419_));
  INV_X1     g2034(.I(new_n1800_), .ZN(new_n2420_));
  NOR4_X1    g2035(.A1(new_n1162_), .A2(new_n1954_), .A3(new_n1771_), .A4(new_n1768_), .ZN(new_n2421_));
  OAI21_X1   g2036(.A1(new_n1779_), .A2(new_n2421_), .B(new_n1786_), .ZN(new_n2422_));
  AOI21_X1   g2037(.A1(new_n2422_), .A2(new_n2419_), .B(new_n2420_), .ZN(new_n2423_));
  OAI21_X1   g2038(.A1(new_n2423_), .A2(new_n1807_), .B(new_n1814_), .ZN(new_n2424_));
  AOI21_X1   g2039(.A1(new_n2424_), .A2(new_n2417_), .B(new_n2418_), .ZN(new_n2425_));
  OAI21_X1   g2040(.A1(new_n2425_), .A2(new_n1835_), .B(new_n1842_), .ZN(new_n2426_));
  AOI21_X1   g2041(.A1(new_n2426_), .A2(new_n2415_), .B(new_n2416_), .ZN(new_n2427_));
  OAI21_X1   g2042(.A1(new_n2427_), .A2(new_n1863_), .B(new_n1870_), .ZN(new_n2428_));
  AOI21_X1   g2043(.A1(new_n2428_), .A2(new_n2413_), .B(new_n2414_), .ZN(new_n2429_));
  OAI21_X1   g2044(.A1(new_n2429_), .A2(new_n1891_), .B(new_n1898_), .ZN(new_n2430_));
  AOI21_X1   g2045(.A1(new_n2430_), .A2(new_n2411_), .B(new_n2412_), .ZN(new_n2431_));
  OAI21_X1   g2046(.A1(new_n2431_), .A2(new_n1919_), .B(new_n1926_), .ZN(new_n2432_));
  AOI21_X1   g2047(.A1(new_n2432_), .A2(new_n2409_), .B(new_n2410_), .ZN(new_n2433_));
  NOR3_X1    g2048(.A1(new_n2237_), .A2(new_n403_), .A3(new_n1392_), .ZN(new_n2434_));
  OAI21_X1   g2049(.A1(new_n2433_), .A2(new_n1945_), .B(new_n2434_), .ZN(new_n2435_));
  NAND2_X1   g2050(.A1(new_n1401_), .A2(new_n1151_), .ZN(new_n2436_));
  AOI21_X1   g2051(.A1(new_n2435_), .A2(new_n2408_), .B(new_n2436_), .ZN(\grant[14] ));
  INV_X1     g2052(.I(new_n1583_), .ZN(new_n2438_));
  INV_X1     g2053(.I(new_n2039_), .ZN(new_n2439_));
  INV_X1     g2054(.I(new_n2041_), .ZN(new_n2440_));
  INV_X1     g2055(.I(new_n2025_), .ZN(new_n2441_));
  INV_X1     g2056(.I(new_n2027_), .ZN(new_n2442_));
  INV_X1     g2057(.I(new_n2011_), .ZN(new_n2443_));
  INV_X1     g2058(.I(new_n2013_), .ZN(new_n2444_));
  INV_X1     g2059(.I(new_n1997_), .ZN(new_n2445_));
  INV_X1     g2060(.I(new_n1999_), .ZN(new_n2446_));
  INV_X1     g2061(.I(new_n1983_), .ZN(new_n2447_));
  INV_X1     g2062(.I(new_n1985_), .ZN(new_n2448_));
  INV_X1     g2063(.I(new_n1969_), .ZN(new_n2449_));
  INV_X1     g2064(.I(new_n1971_), .ZN(new_n2450_));
  NOR4_X1    g2065(.A1(new_n1409_), .A2(new_n436_), .A3(new_n1956_), .A4(new_n2056_), .ZN(new_n2451_));
  OAI21_X1   g2066(.A1(new_n1961_), .A2(new_n2451_), .B(new_n1964_), .ZN(new_n2452_));
  AOI21_X1   g2067(.A1(new_n2452_), .A2(new_n2449_), .B(new_n2450_), .ZN(new_n2453_));
  OAI21_X1   g2068(.A1(new_n2453_), .A2(new_n1975_), .B(new_n1978_), .ZN(new_n2454_));
  AOI21_X1   g2069(.A1(new_n2454_), .A2(new_n2447_), .B(new_n2448_), .ZN(new_n2455_));
  OAI21_X1   g2070(.A1(new_n2455_), .A2(new_n1989_), .B(new_n1992_), .ZN(new_n2456_));
  AOI21_X1   g2071(.A1(new_n2456_), .A2(new_n2445_), .B(new_n2446_), .ZN(new_n2457_));
  OAI21_X1   g2072(.A1(new_n2457_), .A2(new_n2003_), .B(new_n2006_), .ZN(new_n2458_));
  AOI21_X1   g2073(.A1(new_n2458_), .A2(new_n2443_), .B(new_n2444_), .ZN(new_n2459_));
  OAI21_X1   g2074(.A1(new_n2459_), .A2(new_n2017_), .B(new_n2020_), .ZN(new_n2460_));
  AOI21_X1   g2075(.A1(new_n2460_), .A2(new_n2441_), .B(new_n2442_), .ZN(new_n2461_));
  OAI21_X1   g2076(.A1(new_n2461_), .A2(new_n2031_), .B(new_n2034_), .ZN(new_n2462_));
  AOI21_X1   g2077(.A1(new_n2462_), .A2(new_n2439_), .B(new_n2440_), .ZN(new_n2463_));
  NOR3_X1    g2078(.A1(new_n2272_), .A2(new_n795_), .A3(new_n1575_), .ZN(new_n2464_));
  OAI21_X1   g2079(.A1(new_n2463_), .A2(new_n2048_), .B(new_n2464_), .ZN(new_n2465_));
  NAND2_X1   g2080(.A1(new_n1584_), .A2(new_n428_), .ZN(new_n2466_));
  AOI21_X1   g2081(.A1(new_n2465_), .A2(new_n2438_), .B(new_n2466_), .ZN(\grant[15] ));
  INV_X1     g2082(.I(new_n1766_), .ZN(new_n2468_));
  INV_X1     g2083(.I(new_n2129_), .ZN(new_n2469_));
  INV_X1     g2084(.I(new_n2132_), .ZN(new_n2470_));
  INV_X1     g2085(.I(new_n2117_), .ZN(new_n2471_));
  INV_X1     g2086(.I(new_n2119_), .ZN(new_n2472_));
  INV_X1     g2087(.I(new_n2105_), .ZN(new_n2473_));
  INV_X1     g2088(.I(new_n2107_), .ZN(new_n2474_));
  INV_X1     g2089(.I(new_n2093_), .ZN(new_n2475_));
  INV_X1     g2090(.I(new_n2095_), .ZN(new_n2476_));
  INV_X1     g2091(.I(new_n2081_), .ZN(new_n2477_));
  INV_X1     g2092(.I(new_n2083_), .ZN(new_n2478_));
  INV_X1     g2093(.I(new_n2069_), .ZN(new_n2479_));
  INV_X1     g2094(.I(new_n2071_), .ZN(new_n2480_));
  NOR4_X1    g2095(.A1(new_n1592_), .A2(new_n825_), .A3(new_n2058_), .A4(new_n2148_), .ZN(new_n2481_));
  OAI21_X1   g2096(.A1(new_n2062_), .A2(new_n2481_), .B(new_n2065_), .ZN(new_n2482_));
  AOI21_X1   g2097(.A1(new_n2482_), .A2(new_n2479_), .B(new_n2480_), .ZN(new_n2483_));
  OAI21_X1   g2098(.A1(new_n2483_), .A2(new_n2074_), .B(new_n2077_), .ZN(new_n2484_));
  AOI21_X1   g2099(.A1(new_n2484_), .A2(new_n2477_), .B(new_n2478_), .ZN(new_n2485_));
  OAI21_X1   g2100(.A1(new_n2485_), .A2(new_n2086_), .B(new_n2089_), .ZN(new_n2486_));
  AOI21_X1   g2101(.A1(new_n2486_), .A2(new_n2475_), .B(new_n2476_), .ZN(new_n2487_));
  OAI21_X1   g2102(.A1(new_n2487_), .A2(new_n2098_), .B(new_n2101_), .ZN(new_n2488_));
  AOI21_X1   g2103(.A1(new_n2488_), .A2(new_n2473_), .B(new_n2474_), .ZN(new_n2489_));
  OAI21_X1   g2104(.A1(new_n2489_), .A2(new_n2110_), .B(new_n2113_), .ZN(new_n2490_));
  AOI21_X1   g2105(.A1(new_n2490_), .A2(new_n2471_), .B(new_n2472_), .ZN(new_n2491_));
  OAI21_X1   g2106(.A1(new_n2491_), .A2(new_n2122_), .B(new_n2125_), .ZN(new_n2492_));
  AOI21_X1   g2107(.A1(new_n2492_), .A2(new_n2469_), .B(new_n2470_), .ZN(new_n2493_));
  NOR3_X1    g2108(.A1(new_n2308_), .A2(new_n1145_), .A3(new_n1759_), .ZN(new_n2494_));
  OAI21_X1   g2109(.A1(new_n2493_), .A2(new_n2139_), .B(new_n2494_), .ZN(new_n2495_));
  NAND2_X1   g2110(.A1(new_n1767_), .A2(new_n817_), .ZN(new_n2496_));
  AOI21_X1   g2111(.A1(new_n2495_), .A2(new_n2468_), .B(new_n2496_), .ZN(\grant[16] ));
  INV_X1     g2112(.I(new_n1955_), .ZN(new_n2498_));
  INV_X1     g2113(.I(new_n2233_), .ZN(new_n2499_));
  INV_X1     g2114(.I(new_n2235_), .ZN(new_n2500_));
  INV_X1     g2115(.I(new_n2219_), .ZN(new_n2501_));
  INV_X1     g2116(.I(new_n2222_), .ZN(new_n2502_));
  INV_X1     g2117(.I(new_n2205_), .ZN(new_n2503_));
  INV_X1     g2118(.I(new_n2208_), .ZN(new_n2504_));
  INV_X1     g2119(.I(new_n2191_), .ZN(new_n2505_));
  INV_X1     g2120(.I(new_n2194_), .ZN(new_n2506_));
  INV_X1     g2121(.I(new_n2177_), .ZN(new_n2507_));
  INV_X1     g2122(.I(new_n2180_), .ZN(new_n2508_));
  INV_X1     g2123(.I(new_n2163_), .ZN(new_n2509_));
  INV_X1     g2124(.I(new_n2166_), .ZN(new_n2510_));
  OAI21_X1   g2125(.A1(new_n432_), .A2(\priority[19] ), .B(new_n1770_), .ZN(new_n2511_));
  NOR3_X1    g2126(.A1(new_n2511_), .A2(new_n1776_), .A3(new_n2151_), .ZN(new_n2512_));
  OAI21_X1   g2127(.A1(new_n2155_), .A2(new_n2512_), .B(new_n2159_), .ZN(new_n2513_));
  AOI21_X1   g2128(.A1(new_n2513_), .A2(new_n2509_), .B(new_n2510_), .ZN(new_n2514_));
  OAI21_X1   g2129(.A1(new_n2514_), .A2(new_n2169_), .B(new_n2173_), .ZN(new_n2515_));
  AOI21_X1   g2130(.A1(new_n2515_), .A2(new_n2507_), .B(new_n2508_), .ZN(new_n2516_));
  OAI21_X1   g2131(.A1(new_n2516_), .A2(new_n2183_), .B(new_n2187_), .ZN(new_n2517_));
  AOI21_X1   g2132(.A1(new_n2517_), .A2(new_n2505_), .B(new_n2506_), .ZN(new_n2518_));
  OAI21_X1   g2133(.A1(new_n2518_), .A2(new_n2197_), .B(new_n2201_), .ZN(new_n2519_));
  AOI21_X1   g2134(.A1(new_n2519_), .A2(new_n2503_), .B(new_n2504_), .ZN(new_n2520_));
  OAI21_X1   g2135(.A1(new_n2520_), .A2(new_n2211_), .B(new_n2215_), .ZN(new_n2521_));
  AOI21_X1   g2136(.A1(new_n2521_), .A2(new_n2501_), .B(new_n2502_), .ZN(new_n2522_));
  OAI21_X1   g2137(.A1(new_n2522_), .A2(new_n2225_), .B(new_n2229_), .ZN(new_n2523_));
  AOI21_X1   g2138(.A1(new_n2523_), .A2(new_n2499_), .B(new_n2500_), .ZN(new_n2524_));
  NOR3_X1    g2139(.A1(new_n410_), .A2(new_n1397_), .A3(new_n1950_), .ZN(new_n2525_));
  OAI21_X1   g2140(.A1(new_n2524_), .A2(new_n2239_), .B(new_n2525_), .ZN(new_n2526_));
  NAND2_X1   g2141(.A1(new_n434_), .A2(new_n1160_), .ZN(new_n2527_));
  AOI21_X1   g2142(.A1(new_n2526_), .A2(new_n2498_), .B(new_n2527_), .ZN(\grant[17] ));
  INV_X1     g2143(.I(new_n2057_), .ZN(new_n2529_));
  INV_X1     g2144(.I(new_n2270_), .ZN(new_n2530_));
  AOI21_X1   g2145(.A1(new_n1590_), .A2(\priority[19] ), .B(\priority[20] ), .ZN(new_n2531_));
  NOR4_X1    g2146(.A1(new_n444_), .A2(new_n446_), .A3(new_n450_), .A4(new_n2531_), .ZN(new_n2532_));
  OAI21_X1   g2147(.A1(new_n467_), .A2(new_n2532_), .B(new_n480_), .ZN(new_n2533_));
  AOI21_X1   g2148(.A1(new_n2533_), .A2(new_n495_), .B(new_n509_), .ZN(new_n2534_));
  OAI21_X1   g2149(.A1(new_n2534_), .A2(new_n523_), .B(new_n536_), .ZN(new_n2535_));
  AOI21_X1   g2150(.A1(new_n2535_), .A2(new_n551_), .B(new_n565_), .ZN(new_n2536_));
  OAI21_X1   g2151(.A1(new_n2536_), .A2(new_n579_), .B(new_n592_), .ZN(new_n2537_));
  AOI21_X1   g2152(.A1(new_n2537_), .A2(new_n607_), .B(new_n621_), .ZN(new_n2538_));
  OAI21_X1   g2153(.A1(new_n2538_), .A2(new_n635_), .B(new_n648_), .ZN(new_n2539_));
  AOI21_X1   g2154(.A1(new_n2539_), .A2(new_n663_), .B(new_n677_), .ZN(new_n2540_));
  OAI21_X1   g2155(.A1(new_n2540_), .A2(new_n691_), .B(new_n704_), .ZN(new_n2541_));
  AOI21_X1   g2156(.A1(new_n2541_), .A2(new_n719_), .B(new_n733_), .ZN(new_n2542_));
  OAI21_X1   g2157(.A1(new_n2542_), .A2(new_n747_), .B(new_n760_), .ZN(new_n2543_));
  AOI21_X1   g2158(.A1(new_n2543_), .A2(new_n775_), .B(new_n2530_), .ZN(new_n2544_));
  NOR3_X1    g2159(.A1(new_n802_), .A2(new_n1580_), .A3(new_n2053_), .ZN(new_n2545_));
  OAI21_X1   g2160(.A1(new_n2544_), .A2(new_n2275_), .B(new_n2545_), .ZN(new_n2546_));
  NAND2_X1   g2161(.A1(new_n823_), .A2(new_n1407_), .ZN(new_n2547_));
  AOI21_X1   g2162(.A1(new_n2546_), .A2(new_n2529_), .B(new_n2547_), .ZN(\grant[18] ));
  INV_X1     g2163(.I(new_n2149_), .ZN(new_n2549_));
  INV_X1     g2164(.I(new_n2306_), .ZN(new_n2550_));
  AOI21_X1   g2165(.A1(new_n1774_), .A2(\priority[20] ), .B(\priority[21] ), .ZN(new_n2551_));
  NOR4_X1    g2166(.A1(new_n832_), .A2(new_n834_), .A3(new_n838_), .A4(new_n2551_), .ZN(new_n2552_));
  OAI21_X1   g2167(.A1(new_n853_), .A2(new_n2552_), .B(new_n865_), .ZN(new_n2553_));
  AOI21_X1   g2168(.A1(new_n2553_), .A2(new_n878_), .B(new_n891_), .ZN(new_n2554_));
  OAI21_X1   g2169(.A1(new_n2554_), .A2(new_n903_), .B(new_n915_), .ZN(new_n2555_));
  AOI21_X1   g2170(.A1(new_n2555_), .A2(new_n928_), .B(new_n941_), .ZN(new_n2556_));
  OAI21_X1   g2171(.A1(new_n2556_), .A2(new_n953_), .B(new_n965_), .ZN(new_n2557_));
  AOI21_X1   g2172(.A1(new_n2557_), .A2(new_n978_), .B(new_n991_), .ZN(new_n2558_));
  OAI21_X1   g2173(.A1(new_n2558_), .A2(new_n1003_), .B(new_n1015_), .ZN(new_n2559_));
  AOI21_X1   g2174(.A1(new_n2559_), .A2(new_n1028_), .B(new_n1041_), .ZN(new_n2560_));
  OAI21_X1   g2175(.A1(new_n2560_), .A2(new_n1053_), .B(new_n1065_), .ZN(new_n2561_));
  AOI21_X1   g2176(.A1(new_n2561_), .A2(new_n1078_), .B(new_n1091_), .ZN(new_n2562_));
  OAI21_X1   g2177(.A1(new_n2562_), .A2(new_n1103_), .B(new_n1115_), .ZN(new_n2563_));
  AOI21_X1   g2178(.A1(new_n2563_), .A2(new_n1128_), .B(new_n2550_), .ZN(new_n2564_));
  NOR3_X1    g2179(.A1(new_n1149_), .A2(new_n1763_), .A3(new_n2145_), .ZN(new_n2565_));
  OAI21_X1   g2180(.A1(new_n2564_), .A2(new_n2311_), .B(new_n2565_), .ZN(new_n2566_));
  NAND2_X1   g2181(.A1(new_n1165_), .A2(new_n1590_), .ZN(new_n2567_));
  AOI21_X1   g2182(.A1(new_n2566_), .A2(new_n2549_), .B(new_n2567_), .ZN(\grant[19] ));
  INV_X1     g2183(.I(new_n2342_), .ZN(new_n2569_));
  OAI21_X1   g2184(.A1(new_n1410_), .A2(\priority[22] ), .B(new_n2150_), .ZN(new_n2570_));
  NOR3_X1    g2185(.A1(new_n2570_), .A2(new_n1171_), .A3(new_n1173_), .ZN(new_n2571_));
  OAI21_X1   g2186(.A1(new_n1186_), .A2(new_n2571_), .B(new_n1194_), .ZN(new_n2572_));
  AOI21_X1   g2187(.A1(new_n2572_), .A2(new_n1204_), .B(new_n1213_), .ZN(new_n2573_));
  OAI21_X1   g2188(.A1(new_n2573_), .A2(new_n1222_), .B(new_n1230_), .ZN(new_n2574_));
  AOI21_X1   g2189(.A1(new_n2574_), .A2(new_n1240_), .B(new_n1249_), .ZN(new_n2575_));
  OAI21_X1   g2190(.A1(new_n2575_), .A2(new_n1258_), .B(new_n1266_), .ZN(new_n2576_));
  AOI21_X1   g2191(.A1(new_n2576_), .A2(new_n1276_), .B(new_n1285_), .ZN(new_n2577_));
  OAI21_X1   g2192(.A1(new_n2577_), .A2(new_n1294_), .B(new_n1302_), .ZN(new_n2578_));
  AOI21_X1   g2193(.A1(new_n2578_), .A2(new_n1312_), .B(new_n1321_), .ZN(new_n2579_));
  OAI21_X1   g2194(.A1(new_n2579_), .A2(new_n1330_), .B(new_n1338_), .ZN(new_n2580_));
  AOI21_X1   g2195(.A1(new_n2580_), .A2(new_n1348_), .B(new_n1357_), .ZN(new_n2581_));
  OAI21_X1   g2196(.A1(new_n2581_), .A2(new_n1366_), .B(new_n1374_), .ZN(new_n2582_));
  AOI21_X1   g2197(.A1(new_n2582_), .A2(new_n1386_), .B(new_n2569_), .ZN(new_n2583_));
  OAI21_X1   g2198(.A1(new_n2583_), .A2(new_n411_), .B(new_n424_), .ZN(new_n2584_));
  NAND2_X1   g2199(.A1(new_n448_), .A2(new_n1774_), .ZN(new_n2585_));
  AOI21_X1   g2200(.A1(new_n2584_), .A2(new_n439_), .B(new_n2585_), .ZN(\grant[20] ));
  INV_X1     g2201(.I(new_n2373_), .ZN(new_n2587_));
  AOI21_X1   g2202(.A1(new_n830_), .A2(\priority[22] ), .B(\priority[23] ), .ZN(new_n2588_));
  NOR4_X1    g2203(.A1(new_n459_), .A2(new_n1415_), .A3(new_n1417_), .A4(new_n2588_), .ZN(new_n2589_));
  OAI21_X1   g2204(.A1(new_n1426_), .A2(new_n2589_), .B(new_n1431_), .ZN(new_n2590_));
  AOI21_X1   g2205(.A1(new_n2590_), .A2(new_n1439_), .B(new_n1445_), .ZN(new_n2591_));
  OAI21_X1   g2206(.A1(new_n2591_), .A2(new_n1452_), .B(new_n1457_), .ZN(new_n2592_));
  AOI21_X1   g2207(.A1(new_n2592_), .A2(new_n1465_), .B(new_n1471_), .ZN(new_n2593_));
  OAI21_X1   g2208(.A1(new_n2593_), .A2(new_n1478_), .B(new_n1483_), .ZN(new_n2594_));
  AOI21_X1   g2209(.A1(new_n2594_), .A2(new_n1491_), .B(new_n1497_), .ZN(new_n2595_));
  OAI21_X1   g2210(.A1(new_n2595_), .A2(new_n1504_), .B(new_n1509_), .ZN(new_n2596_));
  AOI21_X1   g2211(.A1(new_n2596_), .A2(new_n1517_), .B(new_n1523_), .ZN(new_n2597_));
  OAI21_X1   g2212(.A1(new_n2597_), .A2(new_n1530_), .B(new_n1535_), .ZN(new_n2598_));
  AOI21_X1   g2213(.A1(new_n2598_), .A2(new_n1543_), .B(new_n1549_), .ZN(new_n2599_));
  OAI21_X1   g2214(.A1(new_n2599_), .A2(new_n1556_), .B(new_n1561_), .ZN(new_n2600_));
  AOI21_X1   g2215(.A1(new_n2600_), .A2(new_n1570_), .B(new_n2587_), .ZN(new_n2601_));
  OAI21_X1   g2216(.A1(new_n2601_), .A2(new_n803_), .B(new_n815_), .ZN(new_n2602_));
  NAND2_X1   g2217(.A1(new_n836_), .A2(new_n442_), .ZN(new_n2603_));
  AOI21_X1   g2218(.A1(new_n2602_), .A2(new_n828_), .B(new_n2603_), .ZN(\grant[21] ));
  INV_X1     g2219(.I(new_n2404_), .ZN(new_n2605_));
  AOI21_X1   g2220(.A1(new_n1169_), .A2(\priority[23] ), .B(\priority[24] ), .ZN(new_n2606_));
  NOR4_X1    g2221(.A1(new_n845_), .A2(new_n1598_), .A3(new_n1600_), .A4(new_n2606_), .ZN(new_n2607_));
  OAI21_X1   g2222(.A1(new_n1609_), .A2(new_n2607_), .B(new_n1614_), .ZN(new_n2608_));
  AOI21_X1   g2223(.A1(new_n2608_), .A2(new_n1622_), .B(new_n1628_), .ZN(new_n2609_));
  OAI21_X1   g2224(.A1(new_n2609_), .A2(new_n1635_), .B(new_n1640_), .ZN(new_n2610_));
  AOI21_X1   g2225(.A1(new_n2610_), .A2(new_n1648_), .B(new_n1654_), .ZN(new_n2611_));
  OAI21_X1   g2226(.A1(new_n2611_), .A2(new_n1661_), .B(new_n1666_), .ZN(new_n2612_));
  AOI21_X1   g2227(.A1(new_n2612_), .A2(new_n1674_), .B(new_n1680_), .ZN(new_n2613_));
  OAI21_X1   g2228(.A1(new_n2613_), .A2(new_n1687_), .B(new_n1692_), .ZN(new_n2614_));
  AOI21_X1   g2229(.A1(new_n2614_), .A2(new_n1700_), .B(new_n1706_), .ZN(new_n2615_));
  OAI21_X1   g2230(.A1(new_n2615_), .A2(new_n1713_), .B(new_n1718_), .ZN(new_n2616_));
  AOI21_X1   g2231(.A1(new_n2616_), .A2(new_n1726_), .B(new_n1732_), .ZN(new_n2617_));
  OAI21_X1   g2232(.A1(new_n2617_), .A2(new_n1739_), .B(new_n1744_), .ZN(new_n2618_));
  AOI21_X1   g2233(.A1(new_n2618_), .A2(new_n1751_), .B(new_n2605_), .ZN(new_n2619_));
  OAI21_X1   g2234(.A1(new_n2619_), .A2(new_n1150_), .B(new_n1158_), .ZN(new_n2620_));
  NAND2_X1   g2235(.A1(new_n1174_), .A2(new_n830_), .ZN(new_n2621_));
  AOI21_X1   g2236(.A1(new_n2620_), .A2(new_n1168_), .B(new_n2621_), .ZN(\grant[22] ));
  INV_X1     g2237(.I(new_n2434_), .ZN(new_n2623_));
  NOR4_X1    g2238(.A1(new_n1181_), .A2(new_n1960_), .A3(new_n1785_), .A4(new_n1782_), .ZN(new_n2624_));
  OAI21_X1   g2239(.A1(new_n1794_), .A2(new_n2624_), .B(new_n1800_), .ZN(new_n2625_));
  AOI21_X1   g2240(.A1(new_n2625_), .A2(new_n1808_), .B(new_n1815_), .ZN(new_n2626_));
  OAI21_X1   g2241(.A1(new_n2626_), .A2(new_n1822_), .B(new_n1828_), .ZN(new_n2627_));
  AOI21_X1   g2242(.A1(new_n2627_), .A2(new_n1836_), .B(new_n1843_), .ZN(new_n2628_));
  OAI21_X1   g2243(.A1(new_n2628_), .A2(new_n1850_), .B(new_n1856_), .ZN(new_n2629_));
  AOI21_X1   g2244(.A1(new_n2629_), .A2(new_n1864_), .B(new_n1871_), .ZN(new_n2630_));
  OAI21_X1   g2245(.A1(new_n2630_), .A2(new_n1878_), .B(new_n1884_), .ZN(new_n2631_));
  AOI21_X1   g2246(.A1(new_n2631_), .A2(new_n1892_), .B(new_n1899_), .ZN(new_n2632_));
  OAI21_X1   g2247(.A1(new_n2632_), .A2(new_n1906_), .B(new_n1912_), .ZN(new_n2633_));
  AOI21_X1   g2248(.A1(new_n2633_), .A2(new_n1920_), .B(new_n1927_), .ZN(new_n2634_));
  OAI21_X1   g2249(.A1(new_n2634_), .A2(new_n1934_), .B(new_n1939_), .ZN(new_n2635_));
  AOI21_X1   g2250(.A1(new_n2635_), .A2(new_n1946_), .B(new_n2623_), .ZN(new_n2636_));
  OAI21_X1   g2251(.A1(new_n2636_), .A2(new_n1400_), .B(new_n1405_), .ZN(new_n2637_));
  NAND2_X1   g2252(.A1(new_n1414_), .A2(new_n1169_), .ZN(new_n2638_));
  AOI21_X1   g2253(.A1(new_n2637_), .A2(new_n1413_), .B(new_n2638_), .ZN(\grant[23] ));
  INV_X1     g2254(.I(new_n2464_), .ZN(new_n2640_));
  NOR4_X1    g2255(.A1(new_n1423_), .A2(new_n465_), .A3(new_n1963_), .A4(new_n2061_), .ZN(new_n2641_));
  OAI21_X1   g2256(.A1(new_n1969_), .A2(new_n2641_), .B(new_n1971_), .ZN(new_n2642_));
  AOI21_X1   g2257(.A1(new_n2642_), .A2(new_n1976_), .B(new_n1979_), .ZN(new_n2643_));
  OAI21_X1   g2258(.A1(new_n2643_), .A2(new_n1983_), .B(new_n1985_), .ZN(new_n2644_));
  AOI21_X1   g2259(.A1(new_n2644_), .A2(new_n1990_), .B(new_n1993_), .ZN(new_n2645_));
  OAI21_X1   g2260(.A1(new_n2645_), .A2(new_n1997_), .B(new_n1999_), .ZN(new_n2646_));
  AOI21_X1   g2261(.A1(new_n2646_), .A2(new_n2004_), .B(new_n2007_), .ZN(new_n2647_));
  OAI21_X1   g2262(.A1(new_n2647_), .A2(new_n2011_), .B(new_n2013_), .ZN(new_n2648_));
  AOI21_X1   g2263(.A1(new_n2648_), .A2(new_n2018_), .B(new_n2021_), .ZN(new_n2649_));
  OAI21_X1   g2264(.A1(new_n2649_), .A2(new_n2025_), .B(new_n2027_), .ZN(new_n2650_));
  AOI21_X1   g2265(.A1(new_n2650_), .A2(new_n2032_), .B(new_n2035_), .ZN(new_n2651_));
  OAI21_X1   g2266(.A1(new_n2651_), .A2(new_n2039_), .B(new_n2041_), .ZN(new_n2652_));
  AOI21_X1   g2267(.A1(new_n2652_), .A2(new_n2049_), .B(new_n2640_), .ZN(new_n2653_));
  OAI21_X1   g2268(.A1(new_n2653_), .A2(new_n1583_), .B(new_n1588_), .ZN(new_n2654_));
  NAND2_X1   g2269(.A1(new_n1597_), .A2(new_n457_), .ZN(new_n2655_));
  AOI21_X1   g2270(.A1(new_n2654_), .A2(new_n1596_), .B(new_n2655_), .ZN(\grant[24] ));
  INV_X1     g2271(.I(new_n2494_), .ZN(new_n2657_));
  NOR4_X1    g2272(.A1(new_n1606_), .A2(new_n851_), .A3(new_n2064_), .A4(new_n2154_), .ZN(new_n2658_));
  OAI21_X1   g2273(.A1(new_n2069_), .A2(new_n2658_), .B(new_n2071_), .ZN(new_n2659_));
  AOI21_X1   g2274(.A1(new_n2659_), .A2(new_n2075_), .B(new_n2078_), .ZN(new_n2660_));
  OAI21_X1   g2275(.A1(new_n2660_), .A2(new_n2081_), .B(new_n2083_), .ZN(new_n2661_));
  AOI21_X1   g2276(.A1(new_n2661_), .A2(new_n2087_), .B(new_n2090_), .ZN(new_n2662_));
  OAI21_X1   g2277(.A1(new_n2662_), .A2(new_n2093_), .B(new_n2095_), .ZN(new_n2663_));
  AOI21_X1   g2278(.A1(new_n2663_), .A2(new_n2099_), .B(new_n2102_), .ZN(new_n2664_));
  OAI21_X1   g2279(.A1(new_n2664_), .A2(new_n2105_), .B(new_n2107_), .ZN(new_n2665_));
  AOI21_X1   g2280(.A1(new_n2665_), .A2(new_n2111_), .B(new_n2114_), .ZN(new_n2666_));
  OAI21_X1   g2281(.A1(new_n2666_), .A2(new_n2117_), .B(new_n2119_), .ZN(new_n2667_));
  AOI21_X1   g2282(.A1(new_n2667_), .A2(new_n2123_), .B(new_n2126_), .ZN(new_n2668_));
  OAI21_X1   g2283(.A1(new_n2668_), .A2(new_n2129_), .B(new_n2132_), .ZN(new_n2669_));
  AOI21_X1   g2284(.A1(new_n2669_), .A2(new_n2140_), .B(new_n2657_), .ZN(new_n2670_));
  OAI21_X1   g2285(.A1(new_n2670_), .A2(new_n1766_), .B(new_n1772_), .ZN(new_n2671_));
  NAND2_X1   g2286(.A1(new_n1781_), .A2(new_n843_), .ZN(new_n2672_));
  AOI21_X1   g2287(.A1(new_n2671_), .A2(new_n1780_), .B(new_n2672_), .ZN(\grant[25] ));
  INV_X1     g2288(.I(new_n2525_), .ZN(new_n2674_));
  OAI21_X1   g2289(.A1(new_n461_), .A2(\priority[28] ), .B(new_n1784_), .ZN(new_n2675_));
  NOR3_X1    g2290(.A1(new_n2675_), .A2(new_n1791_), .A3(new_n2158_), .ZN(new_n2676_));
  OAI21_X1   g2291(.A1(new_n2163_), .A2(new_n2676_), .B(new_n2166_), .ZN(new_n2677_));
  AOI21_X1   g2292(.A1(new_n2677_), .A2(new_n2170_), .B(new_n2174_), .ZN(new_n2678_));
  OAI21_X1   g2293(.A1(new_n2678_), .A2(new_n2177_), .B(new_n2180_), .ZN(new_n2679_));
  AOI21_X1   g2294(.A1(new_n2679_), .A2(new_n2184_), .B(new_n2188_), .ZN(new_n2680_));
  OAI21_X1   g2295(.A1(new_n2680_), .A2(new_n2191_), .B(new_n2194_), .ZN(new_n2681_));
  AOI21_X1   g2296(.A1(new_n2681_), .A2(new_n2198_), .B(new_n2202_), .ZN(new_n2682_));
  OAI21_X1   g2297(.A1(new_n2682_), .A2(new_n2205_), .B(new_n2208_), .ZN(new_n2683_));
  AOI21_X1   g2298(.A1(new_n2683_), .A2(new_n2212_), .B(new_n2216_), .ZN(new_n2684_));
  OAI21_X1   g2299(.A1(new_n2684_), .A2(new_n2219_), .B(new_n2222_), .ZN(new_n2685_));
  AOI21_X1   g2300(.A1(new_n2685_), .A2(new_n2226_), .B(new_n2230_), .ZN(new_n2686_));
  OAI21_X1   g2301(.A1(new_n2686_), .A2(new_n2233_), .B(new_n2235_), .ZN(new_n2687_));
  AOI21_X1   g2302(.A1(new_n2687_), .A2(new_n2240_), .B(new_n2674_), .ZN(new_n2688_));
  OAI21_X1   g2303(.A1(new_n2688_), .A2(new_n1955_), .B(new_n1957_), .ZN(new_n2689_));
  NAND2_X1   g2304(.A1(new_n463_), .A2(new_n1179_), .ZN(new_n2690_));
  AOI21_X1   g2305(.A1(new_n2689_), .A2(new_n1962_), .B(new_n2690_), .ZN(\grant[26] ));
  INV_X1     g2306(.I(new_n2545_), .ZN(new_n2692_));
  AOI21_X1   g2307(.A1(new_n1604_), .A2(\priority[28] ), .B(\priority[29] ), .ZN(new_n2693_));
  NOR4_X1    g2308(.A1(new_n472_), .A2(new_n474_), .A3(new_n478_), .A4(new_n2693_), .ZN(new_n2694_));
  OAI21_X1   g2309(.A1(new_n494_), .A2(new_n2694_), .B(new_n508_), .ZN(new_n2695_));
  AOI21_X1   g2310(.A1(new_n2695_), .A2(new_n2251_), .B(new_n2252_), .ZN(new_n2696_));
  OAI21_X1   g2311(.A1(new_n2696_), .A2(new_n550_), .B(new_n564_), .ZN(new_n2697_));
  AOI21_X1   g2312(.A1(new_n2697_), .A2(new_n2249_), .B(new_n2250_), .ZN(new_n2698_));
  OAI21_X1   g2313(.A1(new_n2698_), .A2(new_n606_), .B(new_n620_), .ZN(new_n2699_));
  AOI21_X1   g2314(.A1(new_n2699_), .A2(new_n2247_), .B(new_n2248_), .ZN(new_n2700_));
  OAI21_X1   g2315(.A1(new_n2700_), .A2(new_n662_), .B(new_n676_), .ZN(new_n2701_));
  AOI21_X1   g2316(.A1(new_n2701_), .A2(new_n2245_), .B(new_n2246_), .ZN(new_n2702_));
  OAI21_X1   g2317(.A1(new_n2702_), .A2(new_n718_), .B(new_n732_), .ZN(new_n2703_));
  AOI21_X1   g2318(.A1(new_n2703_), .A2(new_n2243_), .B(new_n2244_), .ZN(new_n2704_));
  OAI21_X1   g2319(.A1(new_n2704_), .A2(new_n774_), .B(new_n2270_), .ZN(new_n2705_));
  AOI21_X1   g2320(.A1(new_n2705_), .A2(new_n2276_), .B(new_n2692_), .ZN(new_n2706_));
  OAI21_X1   g2321(.A1(new_n2706_), .A2(new_n2057_), .B(new_n2059_), .ZN(new_n2707_));
  NAND2_X1   g2322(.A1(new_n849_), .A2(new_n1421_), .ZN(new_n2708_));
  AOI21_X1   g2323(.A1(new_n2707_), .A2(new_n2063_), .B(new_n2708_), .ZN(\grant[27] ));
  INV_X1     g2324(.I(new_n2565_), .ZN(new_n2710_));
  AOI21_X1   g2325(.A1(new_n1789_), .A2(\priority[29] ), .B(\priority[30] ), .ZN(new_n2711_));
  NOR4_X1    g2326(.A1(new_n857_), .A2(new_n859_), .A3(new_n863_), .A4(new_n2711_), .ZN(new_n2712_));
  OAI21_X1   g2327(.A1(new_n877_), .A2(new_n2712_), .B(new_n890_), .ZN(new_n2713_));
  AOI21_X1   g2328(.A1(new_n2713_), .A2(new_n2287_), .B(new_n2288_), .ZN(new_n2714_));
  OAI21_X1   g2329(.A1(new_n2714_), .A2(new_n927_), .B(new_n940_), .ZN(new_n2715_));
  AOI21_X1   g2330(.A1(new_n2715_), .A2(new_n2285_), .B(new_n2286_), .ZN(new_n2716_));
  OAI21_X1   g2331(.A1(new_n2716_), .A2(new_n977_), .B(new_n990_), .ZN(new_n2717_));
  AOI21_X1   g2332(.A1(new_n2717_), .A2(new_n2283_), .B(new_n2284_), .ZN(new_n2718_));
  OAI21_X1   g2333(.A1(new_n2718_), .A2(new_n1027_), .B(new_n1040_), .ZN(new_n2719_));
  AOI21_X1   g2334(.A1(new_n2719_), .A2(new_n2281_), .B(new_n2282_), .ZN(new_n2720_));
  OAI21_X1   g2335(.A1(new_n2720_), .A2(new_n1077_), .B(new_n1090_), .ZN(new_n2721_));
  AOI21_X1   g2336(.A1(new_n2721_), .A2(new_n2279_), .B(new_n2280_), .ZN(new_n2722_));
  OAI21_X1   g2337(.A1(new_n2722_), .A2(new_n1127_), .B(new_n2306_), .ZN(new_n2723_));
  AOI21_X1   g2338(.A1(new_n2723_), .A2(new_n2312_), .B(new_n2710_), .ZN(new_n2724_));
  OAI21_X1   g2339(.A1(new_n2724_), .A2(new_n2149_), .B(new_n2152_), .ZN(new_n2725_));
  NAND2_X1   g2340(.A1(new_n1184_), .A2(new_n1604_), .ZN(new_n2726_));
  AOI21_X1   g2341(.A1(new_n2725_), .A2(new_n2156_), .B(new_n2726_), .ZN(\grant[28] ));
  INV_X1     g2342(.I(new_n424_), .ZN(new_n2728_));
  OAI21_X1   g2343(.A1(new_n1424_), .A2(\priority[31] ), .B(new_n2157_), .ZN(new_n2729_));
  NOR3_X1    g2344(.A1(new_n2729_), .A2(new_n1189_), .A3(new_n1191_), .ZN(new_n2730_));
  OAI21_X1   g2345(.A1(new_n1203_), .A2(new_n2730_), .B(new_n1212_), .ZN(new_n2731_));
  AOI21_X1   g2346(.A1(new_n2731_), .A2(new_n2324_), .B(new_n2325_), .ZN(new_n2732_));
  OAI21_X1   g2347(.A1(new_n2732_), .A2(new_n1239_), .B(new_n1248_), .ZN(new_n2733_));
  AOI21_X1   g2348(.A1(new_n2733_), .A2(new_n2322_), .B(new_n2323_), .ZN(new_n2734_));
  OAI21_X1   g2349(.A1(new_n2734_), .A2(new_n1275_), .B(new_n1284_), .ZN(new_n2735_));
  AOI21_X1   g2350(.A1(new_n2735_), .A2(new_n2320_), .B(new_n2321_), .ZN(new_n2736_));
  OAI21_X1   g2351(.A1(new_n2736_), .A2(new_n1311_), .B(new_n1320_), .ZN(new_n2737_));
  AOI21_X1   g2352(.A1(new_n2737_), .A2(new_n2318_), .B(new_n2319_), .ZN(new_n2738_));
  OAI21_X1   g2353(.A1(new_n2738_), .A2(new_n1347_), .B(new_n1356_), .ZN(new_n2739_));
  AOI21_X1   g2354(.A1(new_n2739_), .A2(new_n2316_), .B(new_n2317_), .ZN(new_n2740_));
  OAI21_X1   g2355(.A1(new_n2740_), .A2(new_n1385_), .B(new_n2342_), .ZN(new_n2741_));
  AOI21_X1   g2356(.A1(new_n2741_), .A2(new_n2315_), .B(new_n2728_), .ZN(new_n2742_));
  OAI21_X1   g2357(.A1(new_n2742_), .A2(new_n438_), .B(new_n452_), .ZN(new_n2743_));
  NAND2_X1   g2358(.A1(new_n476_), .A2(new_n1789_), .ZN(new_n2744_));
  AOI21_X1   g2359(.A1(new_n2743_), .A2(new_n2253_), .B(new_n2744_), .ZN(\grant[29] ));
  INV_X1     g2360(.I(new_n815_), .ZN(new_n2746_));
  AOI21_X1   g2361(.A1(new_n855_), .A2(\priority[31] ), .B(\priority[32] ), .ZN(new_n2747_));
  NOR4_X1    g2362(.A1(new_n486_), .A2(new_n1428_), .A3(new_n1430_), .A4(new_n2747_), .ZN(new_n2748_));
  OAI21_X1   g2363(.A1(new_n1438_), .A2(new_n2748_), .B(new_n1444_), .ZN(new_n2749_));
  AOI21_X1   g2364(.A1(new_n2749_), .A2(new_n2355_), .B(new_n2356_), .ZN(new_n2750_));
  OAI21_X1   g2365(.A1(new_n2750_), .A2(new_n1464_), .B(new_n1470_), .ZN(new_n2751_));
  AOI21_X1   g2366(.A1(new_n2751_), .A2(new_n2353_), .B(new_n2354_), .ZN(new_n2752_));
  OAI21_X1   g2367(.A1(new_n2752_), .A2(new_n1490_), .B(new_n1496_), .ZN(new_n2753_));
  AOI21_X1   g2368(.A1(new_n2753_), .A2(new_n2351_), .B(new_n2352_), .ZN(new_n2754_));
  OAI21_X1   g2369(.A1(new_n2754_), .A2(new_n1516_), .B(new_n1522_), .ZN(new_n2755_));
  AOI21_X1   g2370(.A1(new_n2755_), .A2(new_n2349_), .B(new_n2350_), .ZN(new_n2756_));
  OAI21_X1   g2371(.A1(new_n2756_), .A2(new_n1542_), .B(new_n1548_), .ZN(new_n2757_));
  AOI21_X1   g2372(.A1(new_n2757_), .A2(new_n2347_), .B(new_n2348_), .ZN(new_n2758_));
  OAI21_X1   g2373(.A1(new_n2758_), .A2(new_n1569_), .B(new_n2373_), .ZN(new_n2759_));
  AOI21_X1   g2374(.A1(new_n2759_), .A2(new_n2346_), .B(new_n2746_), .ZN(new_n2760_));
  OAI21_X1   g2375(.A1(new_n2760_), .A2(new_n827_), .B(new_n840_), .ZN(new_n2761_));
  NAND2_X1   g2376(.A1(new_n861_), .A2(new_n470_), .ZN(new_n2762_));
  AOI21_X1   g2377(.A1(new_n2761_), .A2(new_n2289_), .B(new_n2762_), .ZN(\grant[30] ));
  INV_X1     g2378(.I(new_n1158_), .ZN(new_n2764_));
  AOI21_X1   g2379(.A1(new_n1187_), .A2(\priority[32] ), .B(\priority[33] ), .ZN(new_n2765_));
  NOR4_X1    g2380(.A1(new_n869_), .A2(new_n1611_), .A3(new_n1613_), .A4(new_n2765_), .ZN(new_n2766_));
  OAI21_X1   g2381(.A1(new_n1621_), .A2(new_n2766_), .B(new_n1627_), .ZN(new_n2767_));
  AOI21_X1   g2382(.A1(new_n2767_), .A2(new_n2386_), .B(new_n2387_), .ZN(new_n2768_));
  OAI21_X1   g2383(.A1(new_n2768_), .A2(new_n1647_), .B(new_n1653_), .ZN(new_n2769_));
  AOI21_X1   g2384(.A1(new_n2769_), .A2(new_n2384_), .B(new_n2385_), .ZN(new_n2770_));
  OAI21_X1   g2385(.A1(new_n2770_), .A2(new_n1673_), .B(new_n1679_), .ZN(new_n2771_));
  AOI21_X1   g2386(.A1(new_n2771_), .A2(new_n2382_), .B(new_n2383_), .ZN(new_n2772_));
  OAI21_X1   g2387(.A1(new_n2772_), .A2(new_n1699_), .B(new_n1705_), .ZN(new_n2773_));
  AOI21_X1   g2388(.A1(new_n2773_), .A2(new_n2380_), .B(new_n2381_), .ZN(new_n2774_));
  OAI21_X1   g2389(.A1(new_n2774_), .A2(new_n1725_), .B(new_n1731_), .ZN(new_n2775_));
  AOI21_X1   g2390(.A1(new_n2775_), .A2(new_n2378_), .B(new_n2379_), .ZN(new_n2776_));
  OAI21_X1   g2391(.A1(new_n2776_), .A2(new_n1750_), .B(new_n2404_), .ZN(new_n2777_));
  AOI21_X1   g2392(.A1(new_n2777_), .A2(new_n2377_), .B(new_n2764_), .ZN(new_n2778_));
  OAI21_X1   g2393(.A1(new_n2778_), .A2(new_n1167_), .B(new_n1176_), .ZN(new_n2779_));
  NAND2_X1   g2394(.A1(new_n1192_), .A2(new_n855_), .ZN(new_n2780_));
  AOI21_X1   g2395(.A1(new_n2779_), .A2(new_n2326_), .B(new_n2780_), .ZN(\grant[31] ));
  INV_X1     g2396(.I(new_n1405_), .ZN(new_n2782_));
  NOR4_X1    g2397(.A1(new_n1198_), .A2(new_n1968_), .A3(new_n1799_), .A4(new_n1796_), .ZN(new_n2783_));
  OAI21_X1   g2398(.A1(new_n1807_), .A2(new_n2783_), .B(new_n1814_), .ZN(new_n2784_));
  AOI21_X1   g2399(.A1(new_n2784_), .A2(new_n2417_), .B(new_n2418_), .ZN(new_n2785_));
  OAI21_X1   g2400(.A1(new_n2785_), .A2(new_n1835_), .B(new_n1842_), .ZN(new_n2786_));
  AOI21_X1   g2401(.A1(new_n2786_), .A2(new_n2415_), .B(new_n2416_), .ZN(new_n2787_));
  OAI21_X1   g2402(.A1(new_n2787_), .A2(new_n1863_), .B(new_n1870_), .ZN(new_n2788_));
  AOI21_X1   g2403(.A1(new_n2788_), .A2(new_n2413_), .B(new_n2414_), .ZN(new_n2789_));
  OAI21_X1   g2404(.A1(new_n2789_), .A2(new_n1891_), .B(new_n1898_), .ZN(new_n2790_));
  AOI21_X1   g2405(.A1(new_n2790_), .A2(new_n2411_), .B(new_n2412_), .ZN(new_n2791_));
  OAI21_X1   g2406(.A1(new_n2791_), .A2(new_n1919_), .B(new_n1926_), .ZN(new_n2792_));
  AOI21_X1   g2407(.A1(new_n2792_), .A2(new_n2409_), .B(new_n2410_), .ZN(new_n2793_));
  OAI21_X1   g2408(.A1(new_n2793_), .A2(new_n1945_), .B(new_n2434_), .ZN(new_n2794_));
  AOI21_X1   g2409(.A1(new_n2794_), .A2(new_n2408_), .B(new_n2782_), .ZN(new_n2795_));
  OAI21_X1   g2410(.A1(new_n2795_), .A2(new_n1412_), .B(new_n1418_), .ZN(new_n2796_));
  NAND2_X1   g2411(.A1(new_n1427_), .A2(new_n1187_), .ZN(new_n2797_));
  AOI21_X1   g2412(.A1(new_n2796_), .A2(new_n2357_), .B(new_n2797_), .ZN(\grant[32] ));
  INV_X1     g2413(.I(new_n1588_), .ZN(new_n2799_));
  NOR4_X1    g2414(.A1(new_n1435_), .A2(new_n492_), .A3(new_n1970_), .A4(new_n2068_), .ZN(new_n2800_));
  OAI21_X1   g2415(.A1(new_n1975_), .A2(new_n2800_), .B(new_n1978_), .ZN(new_n2801_));
  AOI21_X1   g2416(.A1(new_n2801_), .A2(new_n2447_), .B(new_n2448_), .ZN(new_n2802_));
  OAI21_X1   g2417(.A1(new_n2802_), .A2(new_n1989_), .B(new_n1992_), .ZN(new_n2803_));
  AOI21_X1   g2418(.A1(new_n2803_), .A2(new_n2445_), .B(new_n2446_), .ZN(new_n2804_));
  OAI21_X1   g2419(.A1(new_n2804_), .A2(new_n2003_), .B(new_n2006_), .ZN(new_n2805_));
  AOI21_X1   g2420(.A1(new_n2805_), .A2(new_n2443_), .B(new_n2444_), .ZN(new_n2806_));
  OAI21_X1   g2421(.A1(new_n2806_), .A2(new_n2017_), .B(new_n2020_), .ZN(new_n2807_));
  AOI21_X1   g2422(.A1(new_n2807_), .A2(new_n2441_), .B(new_n2442_), .ZN(new_n2808_));
  OAI21_X1   g2423(.A1(new_n2808_), .A2(new_n2031_), .B(new_n2034_), .ZN(new_n2809_));
  AOI21_X1   g2424(.A1(new_n2809_), .A2(new_n2439_), .B(new_n2440_), .ZN(new_n2810_));
  OAI21_X1   g2425(.A1(new_n2810_), .A2(new_n2048_), .B(new_n2464_), .ZN(new_n2811_));
  AOI21_X1   g2426(.A1(new_n2811_), .A2(new_n2438_), .B(new_n2799_), .ZN(new_n2812_));
  OAI21_X1   g2427(.A1(new_n2812_), .A2(new_n1595_), .B(new_n1601_), .ZN(new_n2813_));
  NAND2_X1   g2428(.A1(new_n1610_), .A2(new_n484_), .ZN(new_n2814_));
  AOI21_X1   g2429(.A1(new_n2813_), .A2(new_n2388_), .B(new_n2814_), .ZN(\grant[33] ));
  INV_X1     g2430(.I(new_n1772_), .ZN(new_n2816_));
  NOR4_X1    g2431(.A1(new_n1618_), .A2(new_n875_), .A3(new_n2070_), .A4(new_n2162_), .ZN(new_n2817_));
  OAI21_X1   g2432(.A1(new_n2074_), .A2(new_n2817_), .B(new_n2077_), .ZN(new_n2818_));
  AOI21_X1   g2433(.A1(new_n2818_), .A2(new_n2477_), .B(new_n2478_), .ZN(new_n2819_));
  OAI21_X1   g2434(.A1(new_n2819_), .A2(new_n2086_), .B(new_n2089_), .ZN(new_n2820_));
  AOI21_X1   g2435(.A1(new_n2820_), .A2(new_n2475_), .B(new_n2476_), .ZN(new_n2821_));
  OAI21_X1   g2436(.A1(new_n2821_), .A2(new_n2098_), .B(new_n2101_), .ZN(new_n2822_));
  AOI21_X1   g2437(.A1(new_n2822_), .A2(new_n2473_), .B(new_n2474_), .ZN(new_n2823_));
  OAI21_X1   g2438(.A1(new_n2823_), .A2(new_n2110_), .B(new_n2113_), .ZN(new_n2824_));
  AOI21_X1   g2439(.A1(new_n2824_), .A2(new_n2471_), .B(new_n2472_), .ZN(new_n2825_));
  OAI21_X1   g2440(.A1(new_n2825_), .A2(new_n2122_), .B(new_n2125_), .ZN(new_n2826_));
  AOI21_X1   g2441(.A1(new_n2826_), .A2(new_n2469_), .B(new_n2470_), .ZN(new_n2827_));
  OAI21_X1   g2442(.A1(new_n2827_), .A2(new_n2139_), .B(new_n2494_), .ZN(new_n2828_));
  AOI21_X1   g2443(.A1(new_n2828_), .A2(new_n2468_), .B(new_n2816_), .ZN(new_n2829_));
  OAI21_X1   g2444(.A1(new_n2829_), .A2(new_n1779_), .B(new_n1786_), .ZN(new_n2830_));
  NAND2_X1   g2445(.A1(new_n1795_), .A2(new_n867_), .ZN(new_n2831_));
  AOI21_X1   g2446(.A1(new_n2830_), .A2(new_n2419_), .B(new_n2831_), .ZN(\grant[34] ));
  INV_X1     g2447(.I(new_n1957_), .ZN(new_n2833_));
  OAI21_X1   g2448(.A1(new_n488_), .A2(\priority[37] ), .B(new_n1798_), .ZN(new_n2834_));
  NOR3_X1    g2449(.A1(new_n2834_), .A2(new_n1804_), .A3(new_n2165_), .ZN(new_n2835_));
  OAI21_X1   g2450(.A1(new_n2169_), .A2(new_n2835_), .B(new_n2173_), .ZN(new_n2836_));
  AOI21_X1   g2451(.A1(new_n2836_), .A2(new_n2507_), .B(new_n2508_), .ZN(new_n2837_));
  OAI21_X1   g2452(.A1(new_n2837_), .A2(new_n2183_), .B(new_n2187_), .ZN(new_n2838_));
  AOI21_X1   g2453(.A1(new_n2838_), .A2(new_n2505_), .B(new_n2506_), .ZN(new_n2839_));
  OAI21_X1   g2454(.A1(new_n2839_), .A2(new_n2197_), .B(new_n2201_), .ZN(new_n2840_));
  AOI21_X1   g2455(.A1(new_n2840_), .A2(new_n2503_), .B(new_n2504_), .ZN(new_n2841_));
  OAI21_X1   g2456(.A1(new_n2841_), .A2(new_n2211_), .B(new_n2215_), .ZN(new_n2842_));
  AOI21_X1   g2457(.A1(new_n2842_), .A2(new_n2501_), .B(new_n2502_), .ZN(new_n2843_));
  OAI21_X1   g2458(.A1(new_n2843_), .A2(new_n2225_), .B(new_n2229_), .ZN(new_n2844_));
  AOI21_X1   g2459(.A1(new_n2844_), .A2(new_n2499_), .B(new_n2500_), .ZN(new_n2845_));
  OAI21_X1   g2460(.A1(new_n2845_), .A2(new_n2239_), .B(new_n2525_), .ZN(new_n2846_));
  AOI21_X1   g2461(.A1(new_n2846_), .A2(new_n2498_), .B(new_n2833_), .ZN(new_n2847_));
  OAI21_X1   g2462(.A1(new_n2847_), .A2(new_n1961_), .B(new_n1964_), .ZN(new_n2848_));
  NAND2_X1   g2463(.A1(new_n490_), .A2(new_n1196_), .ZN(new_n2849_));
  AOI21_X1   g2464(.A1(new_n2848_), .A2(new_n2449_), .B(new_n2849_), .ZN(\grant[35] ));
  INV_X1     g2465(.I(new_n2059_), .ZN(new_n2851_));
  AOI21_X1   g2466(.A1(new_n1616_), .A2(\priority[37] ), .B(\priority[38] ), .ZN(new_n2852_));
  NOR4_X1    g2467(.A1(new_n500_), .A2(new_n502_), .A3(new_n506_), .A4(new_n2852_), .ZN(new_n2853_));
  OAI21_X1   g2468(.A1(new_n523_), .A2(new_n2853_), .B(new_n536_), .ZN(new_n2854_));
  AOI21_X1   g2469(.A1(new_n2854_), .A2(new_n551_), .B(new_n565_), .ZN(new_n2855_));
  OAI21_X1   g2470(.A1(new_n2855_), .A2(new_n579_), .B(new_n592_), .ZN(new_n2856_));
  AOI21_X1   g2471(.A1(new_n2856_), .A2(new_n607_), .B(new_n621_), .ZN(new_n2857_));
  OAI21_X1   g2472(.A1(new_n2857_), .A2(new_n635_), .B(new_n648_), .ZN(new_n2858_));
  AOI21_X1   g2473(.A1(new_n2858_), .A2(new_n663_), .B(new_n677_), .ZN(new_n2859_));
  OAI21_X1   g2474(.A1(new_n2859_), .A2(new_n691_), .B(new_n704_), .ZN(new_n2860_));
  AOI21_X1   g2475(.A1(new_n2860_), .A2(new_n719_), .B(new_n733_), .ZN(new_n2861_));
  OAI21_X1   g2476(.A1(new_n2861_), .A2(new_n747_), .B(new_n760_), .ZN(new_n2862_));
  AOI21_X1   g2477(.A1(new_n2862_), .A2(new_n775_), .B(new_n2530_), .ZN(new_n2863_));
  OAI21_X1   g2478(.A1(new_n2863_), .A2(new_n2275_), .B(new_n2545_), .ZN(new_n2864_));
  AOI21_X1   g2479(.A1(new_n2864_), .A2(new_n2529_), .B(new_n2851_), .ZN(new_n2865_));
  OAI21_X1   g2480(.A1(new_n2865_), .A2(new_n2062_), .B(new_n2065_), .ZN(new_n2866_));
  NAND2_X1   g2481(.A1(new_n873_), .A2(new_n1433_), .ZN(new_n2867_));
  AOI21_X1   g2482(.A1(new_n2866_), .A2(new_n2479_), .B(new_n2867_), .ZN(\grant[36] ));
  INV_X1     g2483(.I(new_n2152_), .ZN(new_n2869_));
  AOI21_X1   g2484(.A1(new_n1802_), .A2(\priority[38] ), .B(\priority[39] ), .ZN(new_n2870_));
  NOR4_X1    g2485(.A1(new_n882_), .A2(new_n884_), .A3(new_n888_), .A4(new_n2870_), .ZN(new_n2871_));
  OAI21_X1   g2486(.A1(new_n903_), .A2(new_n2871_), .B(new_n915_), .ZN(new_n2872_));
  AOI21_X1   g2487(.A1(new_n2872_), .A2(new_n928_), .B(new_n941_), .ZN(new_n2873_));
  OAI21_X1   g2488(.A1(new_n2873_), .A2(new_n953_), .B(new_n965_), .ZN(new_n2874_));
  AOI21_X1   g2489(.A1(new_n2874_), .A2(new_n978_), .B(new_n991_), .ZN(new_n2875_));
  OAI21_X1   g2490(.A1(new_n2875_), .A2(new_n1003_), .B(new_n1015_), .ZN(new_n2876_));
  AOI21_X1   g2491(.A1(new_n2876_), .A2(new_n1028_), .B(new_n1041_), .ZN(new_n2877_));
  OAI21_X1   g2492(.A1(new_n2877_), .A2(new_n1053_), .B(new_n1065_), .ZN(new_n2878_));
  AOI21_X1   g2493(.A1(new_n2878_), .A2(new_n1078_), .B(new_n1091_), .ZN(new_n2879_));
  OAI21_X1   g2494(.A1(new_n2879_), .A2(new_n1103_), .B(new_n1115_), .ZN(new_n2880_));
  AOI21_X1   g2495(.A1(new_n2880_), .A2(new_n1128_), .B(new_n2550_), .ZN(new_n2881_));
  OAI21_X1   g2496(.A1(new_n2881_), .A2(new_n2311_), .B(new_n2565_), .ZN(new_n2882_));
  AOI21_X1   g2497(.A1(new_n2882_), .A2(new_n2549_), .B(new_n2869_), .ZN(new_n2883_));
  OAI21_X1   g2498(.A1(new_n2883_), .A2(new_n2155_), .B(new_n2159_), .ZN(new_n2884_));
  NAND2_X1   g2499(.A1(new_n1201_), .A2(new_n1616_), .ZN(new_n2885_));
  AOI21_X1   g2500(.A1(new_n2884_), .A2(new_n2509_), .B(new_n2885_), .ZN(\grant[37] ));
  OAI21_X1   g2501(.A1(new_n1436_), .A2(\priority[40] ), .B(new_n2164_), .ZN(new_n2887_));
  NOR3_X1    g2502(.A1(new_n2887_), .A2(new_n1207_), .A3(new_n1209_), .ZN(new_n2888_));
  OAI21_X1   g2503(.A1(new_n1222_), .A2(new_n2888_), .B(new_n1230_), .ZN(new_n2889_));
  AOI21_X1   g2504(.A1(new_n2889_), .A2(new_n1240_), .B(new_n1249_), .ZN(new_n2890_));
  OAI21_X1   g2505(.A1(new_n2890_), .A2(new_n1258_), .B(new_n1266_), .ZN(new_n2891_));
  AOI21_X1   g2506(.A1(new_n2891_), .A2(new_n1276_), .B(new_n1285_), .ZN(new_n2892_));
  OAI21_X1   g2507(.A1(new_n2892_), .A2(new_n1294_), .B(new_n1302_), .ZN(new_n2893_));
  AOI21_X1   g2508(.A1(new_n2893_), .A2(new_n1312_), .B(new_n1321_), .ZN(new_n2894_));
  OAI21_X1   g2509(.A1(new_n2894_), .A2(new_n1330_), .B(new_n1338_), .ZN(new_n2895_));
  AOI21_X1   g2510(.A1(new_n2895_), .A2(new_n1348_), .B(new_n1357_), .ZN(new_n2896_));
  OAI21_X1   g2511(.A1(new_n2896_), .A2(new_n1366_), .B(new_n1374_), .ZN(new_n2897_));
  AOI21_X1   g2512(.A1(new_n2897_), .A2(new_n1386_), .B(new_n2569_), .ZN(new_n2898_));
  OAI21_X1   g2513(.A1(new_n2898_), .A2(new_n411_), .B(new_n424_), .ZN(new_n2899_));
  AOI21_X1   g2514(.A1(new_n2899_), .A2(new_n439_), .B(new_n453_), .ZN(new_n2900_));
  OAI21_X1   g2515(.A1(new_n2900_), .A2(new_n467_), .B(new_n480_), .ZN(new_n2901_));
  NAND2_X1   g2516(.A1(new_n504_), .A2(new_n1802_), .ZN(new_n2902_));
  AOI21_X1   g2517(.A1(new_n2901_), .A2(new_n495_), .B(new_n2902_), .ZN(\grant[38] ));
  AOI21_X1   g2518(.A1(new_n880_), .A2(\priority[40] ), .B(\priority[41] ), .ZN(new_n2904_));
  NOR4_X1    g2519(.A1(new_n515_), .A2(new_n1441_), .A3(new_n1443_), .A4(new_n2904_), .ZN(new_n2905_));
  OAI21_X1   g2520(.A1(new_n1452_), .A2(new_n2905_), .B(new_n1457_), .ZN(new_n2906_));
  AOI21_X1   g2521(.A1(new_n2906_), .A2(new_n1465_), .B(new_n1471_), .ZN(new_n2907_));
  OAI21_X1   g2522(.A1(new_n2907_), .A2(new_n1478_), .B(new_n1483_), .ZN(new_n2908_));
  AOI21_X1   g2523(.A1(new_n2908_), .A2(new_n1491_), .B(new_n1497_), .ZN(new_n2909_));
  OAI21_X1   g2524(.A1(new_n2909_), .A2(new_n1504_), .B(new_n1509_), .ZN(new_n2910_));
  AOI21_X1   g2525(.A1(new_n2910_), .A2(new_n1517_), .B(new_n1523_), .ZN(new_n2911_));
  OAI21_X1   g2526(.A1(new_n2911_), .A2(new_n1530_), .B(new_n1535_), .ZN(new_n2912_));
  AOI21_X1   g2527(.A1(new_n2912_), .A2(new_n1543_), .B(new_n1549_), .ZN(new_n2913_));
  OAI21_X1   g2528(.A1(new_n2913_), .A2(new_n1556_), .B(new_n1561_), .ZN(new_n2914_));
  AOI21_X1   g2529(.A1(new_n2914_), .A2(new_n1570_), .B(new_n2587_), .ZN(new_n2915_));
  OAI21_X1   g2530(.A1(new_n2915_), .A2(new_n803_), .B(new_n815_), .ZN(new_n2916_));
  AOI21_X1   g2531(.A1(new_n2916_), .A2(new_n828_), .B(new_n841_), .ZN(new_n2917_));
  OAI21_X1   g2532(.A1(new_n2917_), .A2(new_n853_), .B(new_n865_), .ZN(new_n2918_));
  NAND2_X1   g2533(.A1(new_n886_), .A2(new_n498_), .ZN(new_n2919_));
  AOI21_X1   g2534(.A1(new_n2918_), .A2(new_n878_), .B(new_n2919_), .ZN(\grant[39] ));
  AOI21_X1   g2535(.A1(new_n1205_), .A2(\priority[41] ), .B(\priority[42] ), .ZN(new_n2921_));
  NOR4_X1    g2536(.A1(new_n895_), .A2(new_n1624_), .A3(new_n1626_), .A4(new_n2921_), .ZN(new_n2922_));
  OAI21_X1   g2537(.A1(new_n1635_), .A2(new_n2922_), .B(new_n1640_), .ZN(new_n2923_));
  AOI21_X1   g2538(.A1(new_n2923_), .A2(new_n1648_), .B(new_n1654_), .ZN(new_n2924_));
  OAI21_X1   g2539(.A1(new_n2924_), .A2(new_n1661_), .B(new_n1666_), .ZN(new_n2925_));
  AOI21_X1   g2540(.A1(new_n2925_), .A2(new_n1674_), .B(new_n1680_), .ZN(new_n2926_));
  OAI21_X1   g2541(.A1(new_n2926_), .A2(new_n1687_), .B(new_n1692_), .ZN(new_n2927_));
  AOI21_X1   g2542(.A1(new_n2927_), .A2(new_n1700_), .B(new_n1706_), .ZN(new_n2928_));
  OAI21_X1   g2543(.A1(new_n2928_), .A2(new_n1713_), .B(new_n1718_), .ZN(new_n2929_));
  AOI21_X1   g2544(.A1(new_n2929_), .A2(new_n1726_), .B(new_n1732_), .ZN(new_n2930_));
  OAI21_X1   g2545(.A1(new_n2930_), .A2(new_n1739_), .B(new_n1744_), .ZN(new_n2931_));
  AOI21_X1   g2546(.A1(new_n2931_), .A2(new_n1751_), .B(new_n2605_), .ZN(new_n2932_));
  OAI21_X1   g2547(.A1(new_n2932_), .A2(new_n1150_), .B(new_n1158_), .ZN(new_n2933_));
  AOI21_X1   g2548(.A1(new_n2933_), .A2(new_n1168_), .B(new_n1177_), .ZN(new_n2934_));
  OAI21_X1   g2549(.A1(new_n2934_), .A2(new_n1186_), .B(new_n1194_), .ZN(new_n2935_));
  NAND2_X1   g2550(.A1(new_n1210_), .A2(new_n880_), .ZN(new_n2936_));
  AOI21_X1   g2551(.A1(new_n2935_), .A2(new_n1204_), .B(new_n2936_), .ZN(\grant[40] ));
  NOR4_X1    g2552(.A1(new_n1217_), .A2(new_n1974_), .A3(new_n1813_), .A4(new_n1810_), .ZN(new_n2938_));
  OAI21_X1   g2553(.A1(new_n1822_), .A2(new_n2938_), .B(new_n1828_), .ZN(new_n2939_));
  AOI21_X1   g2554(.A1(new_n2939_), .A2(new_n1836_), .B(new_n1843_), .ZN(new_n2940_));
  OAI21_X1   g2555(.A1(new_n2940_), .A2(new_n1850_), .B(new_n1856_), .ZN(new_n2941_));
  AOI21_X1   g2556(.A1(new_n2941_), .A2(new_n1864_), .B(new_n1871_), .ZN(new_n2942_));
  OAI21_X1   g2557(.A1(new_n2942_), .A2(new_n1878_), .B(new_n1884_), .ZN(new_n2943_));
  AOI21_X1   g2558(.A1(new_n2943_), .A2(new_n1892_), .B(new_n1899_), .ZN(new_n2944_));
  OAI21_X1   g2559(.A1(new_n2944_), .A2(new_n1906_), .B(new_n1912_), .ZN(new_n2945_));
  AOI21_X1   g2560(.A1(new_n2945_), .A2(new_n1920_), .B(new_n1927_), .ZN(new_n2946_));
  OAI21_X1   g2561(.A1(new_n2946_), .A2(new_n1934_), .B(new_n1939_), .ZN(new_n2947_));
  AOI21_X1   g2562(.A1(new_n2947_), .A2(new_n1946_), .B(new_n2623_), .ZN(new_n2948_));
  OAI21_X1   g2563(.A1(new_n2948_), .A2(new_n1400_), .B(new_n1405_), .ZN(new_n2949_));
  AOI21_X1   g2564(.A1(new_n2949_), .A2(new_n1413_), .B(new_n1419_), .ZN(new_n2950_));
  OAI21_X1   g2565(.A1(new_n2950_), .A2(new_n1426_), .B(new_n1431_), .ZN(new_n2951_));
  NAND2_X1   g2566(.A1(new_n1440_), .A2(new_n1205_), .ZN(new_n2952_));
  AOI21_X1   g2567(.A1(new_n2951_), .A2(new_n1439_), .B(new_n2952_), .ZN(\grant[41] ));
  NOR4_X1    g2568(.A1(new_n1449_), .A2(new_n521_), .A3(new_n1977_), .A4(new_n2073_), .ZN(new_n2954_));
  OAI21_X1   g2569(.A1(new_n1983_), .A2(new_n2954_), .B(new_n1985_), .ZN(new_n2955_));
  AOI21_X1   g2570(.A1(new_n2955_), .A2(new_n1990_), .B(new_n1993_), .ZN(new_n2956_));
  OAI21_X1   g2571(.A1(new_n2956_), .A2(new_n1997_), .B(new_n1999_), .ZN(new_n2957_));
  AOI21_X1   g2572(.A1(new_n2957_), .A2(new_n2004_), .B(new_n2007_), .ZN(new_n2958_));
  OAI21_X1   g2573(.A1(new_n2958_), .A2(new_n2011_), .B(new_n2013_), .ZN(new_n2959_));
  AOI21_X1   g2574(.A1(new_n2959_), .A2(new_n2018_), .B(new_n2021_), .ZN(new_n2960_));
  OAI21_X1   g2575(.A1(new_n2960_), .A2(new_n2025_), .B(new_n2027_), .ZN(new_n2961_));
  AOI21_X1   g2576(.A1(new_n2961_), .A2(new_n2032_), .B(new_n2035_), .ZN(new_n2962_));
  OAI21_X1   g2577(.A1(new_n2962_), .A2(new_n2039_), .B(new_n2041_), .ZN(new_n2963_));
  AOI21_X1   g2578(.A1(new_n2963_), .A2(new_n2049_), .B(new_n2640_), .ZN(new_n2964_));
  OAI21_X1   g2579(.A1(new_n2964_), .A2(new_n1583_), .B(new_n1588_), .ZN(new_n2965_));
  AOI21_X1   g2580(.A1(new_n2965_), .A2(new_n1596_), .B(new_n1602_), .ZN(new_n2966_));
  OAI21_X1   g2581(.A1(new_n2966_), .A2(new_n1609_), .B(new_n1614_), .ZN(new_n2967_));
  NAND2_X1   g2582(.A1(new_n1623_), .A2(new_n513_), .ZN(new_n2968_));
  AOI21_X1   g2583(.A1(new_n2967_), .A2(new_n1622_), .B(new_n2968_), .ZN(\grant[42] ));
  NOR4_X1    g2584(.A1(new_n1632_), .A2(new_n901_), .A3(new_n2076_), .A4(new_n2168_), .ZN(new_n2970_));
  OAI21_X1   g2585(.A1(new_n2081_), .A2(new_n2970_), .B(new_n2083_), .ZN(new_n2971_));
  AOI21_X1   g2586(.A1(new_n2971_), .A2(new_n2087_), .B(new_n2090_), .ZN(new_n2972_));
  OAI21_X1   g2587(.A1(new_n2972_), .A2(new_n2093_), .B(new_n2095_), .ZN(new_n2973_));
  AOI21_X1   g2588(.A1(new_n2973_), .A2(new_n2099_), .B(new_n2102_), .ZN(new_n2974_));
  OAI21_X1   g2589(.A1(new_n2974_), .A2(new_n2105_), .B(new_n2107_), .ZN(new_n2975_));
  AOI21_X1   g2590(.A1(new_n2975_), .A2(new_n2111_), .B(new_n2114_), .ZN(new_n2976_));
  OAI21_X1   g2591(.A1(new_n2976_), .A2(new_n2117_), .B(new_n2119_), .ZN(new_n2977_));
  AOI21_X1   g2592(.A1(new_n2977_), .A2(new_n2123_), .B(new_n2126_), .ZN(new_n2978_));
  OAI21_X1   g2593(.A1(new_n2978_), .A2(new_n2129_), .B(new_n2132_), .ZN(new_n2979_));
  AOI21_X1   g2594(.A1(new_n2979_), .A2(new_n2140_), .B(new_n2657_), .ZN(new_n2980_));
  OAI21_X1   g2595(.A1(new_n2980_), .A2(new_n1766_), .B(new_n1772_), .ZN(new_n2981_));
  AOI21_X1   g2596(.A1(new_n2981_), .A2(new_n1780_), .B(new_n1787_), .ZN(new_n2982_));
  OAI21_X1   g2597(.A1(new_n2982_), .A2(new_n1794_), .B(new_n1800_), .ZN(new_n2983_));
  NAND2_X1   g2598(.A1(new_n1809_), .A2(new_n893_), .ZN(new_n2984_));
  AOI21_X1   g2599(.A1(new_n2983_), .A2(new_n1808_), .B(new_n2984_), .ZN(\grant[43] ));
  OAI21_X1   g2600(.A1(new_n517_), .A2(\priority[46] ), .B(new_n1812_), .ZN(new_n2986_));
  NOR3_X1    g2601(.A1(new_n2986_), .A2(new_n1819_), .A3(new_n2172_), .ZN(new_n2987_));
  OAI21_X1   g2602(.A1(new_n2177_), .A2(new_n2987_), .B(new_n2180_), .ZN(new_n2988_));
  AOI21_X1   g2603(.A1(new_n2988_), .A2(new_n2184_), .B(new_n2188_), .ZN(new_n2989_));
  OAI21_X1   g2604(.A1(new_n2989_), .A2(new_n2191_), .B(new_n2194_), .ZN(new_n2990_));
  AOI21_X1   g2605(.A1(new_n2990_), .A2(new_n2198_), .B(new_n2202_), .ZN(new_n2991_));
  OAI21_X1   g2606(.A1(new_n2991_), .A2(new_n2205_), .B(new_n2208_), .ZN(new_n2992_));
  AOI21_X1   g2607(.A1(new_n2992_), .A2(new_n2212_), .B(new_n2216_), .ZN(new_n2993_));
  OAI21_X1   g2608(.A1(new_n2993_), .A2(new_n2219_), .B(new_n2222_), .ZN(new_n2994_));
  AOI21_X1   g2609(.A1(new_n2994_), .A2(new_n2226_), .B(new_n2230_), .ZN(new_n2995_));
  OAI21_X1   g2610(.A1(new_n2995_), .A2(new_n2233_), .B(new_n2235_), .ZN(new_n2996_));
  AOI21_X1   g2611(.A1(new_n2996_), .A2(new_n2240_), .B(new_n2674_), .ZN(new_n2997_));
  OAI21_X1   g2612(.A1(new_n2997_), .A2(new_n1955_), .B(new_n1957_), .ZN(new_n2998_));
  AOI21_X1   g2613(.A1(new_n2998_), .A2(new_n1962_), .B(new_n1965_), .ZN(new_n2999_));
  OAI21_X1   g2614(.A1(new_n2999_), .A2(new_n1969_), .B(new_n1971_), .ZN(new_n3000_));
  NAND2_X1   g2615(.A1(new_n519_), .A2(new_n1215_), .ZN(new_n3001_));
  AOI21_X1   g2616(.A1(new_n3000_), .A2(new_n1976_), .B(new_n3001_), .ZN(\grant[44] ));
  AOI21_X1   g2617(.A1(new_n1630_), .A2(\priority[46] ), .B(\priority[47] ), .ZN(new_n3003_));
  NOR4_X1    g2618(.A1(new_n528_), .A2(new_n530_), .A3(new_n534_), .A4(new_n3003_), .ZN(new_n3004_));
  OAI21_X1   g2619(.A1(new_n550_), .A2(new_n3004_), .B(new_n564_), .ZN(new_n3005_));
  AOI21_X1   g2620(.A1(new_n3005_), .A2(new_n2249_), .B(new_n2250_), .ZN(new_n3006_));
  OAI21_X1   g2621(.A1(new_n3006_), .A2(new_n606_), .B(new_n620_), .ZN(new_n3007_));
  AOI21_X1   g2622(.A1(new_n3007_), .A2(new_n2247_), .B(new_n2248_), .ZN(new_n3008_));
  OAI21_X1   g2623(.A1(new_n3008_), .A2(new_n662_), .B(new_n676_), .ZN(new_n3009_));
  AOI21_X1   g2624(.A1(new_n3009_), .A2(new_n2245_), .B(new_n2246_), .ZN(new_n3010_));
  OAI21_X1   g2625(.A1(new_n3010_), .A2(new_n718_), .B(new_n732_), .ZN(new_n3011_));
  AOI21_X1   g2626(.A1(new_n3011_), .A2(new_n2243_), .B(new_n2244_), .ZN(new_n3012_));
  OAI21_X1   g2627(.A1(new_n3012_), .A2(new_n774_), .B(new_n2270_), .ZN(new_n3013_));
  AOI21_X1   g2628(.A1(new_n3013_), .A2(new_n2276_), .B(new_n2692_), .ZN(new_n3014_));
  OAI21_X1   g2629(.A1(new_n3014_), .A2(new_n2057_), .B(new_n2059_), .ZN(new_n3015_));
  AOI21_X1   g2630(.A1(new_n3015_), .A2(new_n2063_), .B(new_n2066_), .ZN(new_n3016_));
  OAI21_X1   g2631(.A1(new_n3016_), .A2(new_n2069_), .B(new_n2071_), .ZN(new_n3017_));
  NAND2_X1   g2632(.A1(new_n899_), .A2(new_n1447_), .ZN(new_n3018_));
  AOI21_X1   g2633(.A1(new_n3017_), .A2(new_n2075_), .B(new_n3018_), .ZN(\grant[45] ));
  AOI21_X1   g2634(.A1(new_n1817_), .A2(\priority[47] ), .B(\priority[48] ), .ZN(new_n3020_));
  NOR4_X1    g2635(.A1(new_n907_), .A2(new_n909_), .A3(new_n913_), .A4(new_n3020_), .ZN(new_n3021_));
  OAI21_X1   g2636(.A1(new_n927_), .A2(new_n3021_), .B(new_n940_), .ZN(new_n3022_));
  AOI21_X1   g2637(.A1(new_n3022_), .A2(new_n2285_), .B(new_n2286_), .ZN(new_n3023_));
  OAI21_X1   g2638(.A1(new_n3023_), .A2(new_n977_), .B(new_n990_), .ZN(new_n3024_));
  AOI21_X1   g2639(.A1(new_n3024_), .A2(new_n2283_), .B(new_n2284_), .ZN(new_n3025_));
  OAI21_X1   g2640(.A1(new_n3025_), .A2(new_n1027_), .B(new_n1040_), .ZN(new_n3026_));
  AOI21_X1   g2641(.A1(new_n3026_), .A2(new_n2281_), .B(new_n2282_), .ZN(new_n3027_));
  OAI21_X1   g2642(.A1(new_n3027_), .A2(new_n1077_), .B(new_n1090_), .ZN(new_n3028_));
  AOI21_X1   g2643(.A1(new_n3028_), .A2(new_n2279_), .B(new_n2280_), .ZN(new_n3029_));
  OAI21_X1   g2644(.A1(new_n3029_), .A2(new_n1127_), .B(new_n2306_), .ZN(new_n3030_));
  AOI21_X1   g2645(.A1(new_n3030_), .A2(new_n2312_), .B(new_n2710_), .ZN(new_n3031_));
  OAI21_X1   g2646(.A1(new_n3031_), .A2(new_n2149_), .B(new_n2152_), .ZN(new_n3032_));
  AOI21_X1   g2647(.A1(new_n3032_), .A2(new_n2156_), .B(new_n2160_), .ZN(new_n3033_));
  OAI21_X1   g2648(.A1(new_n3033_), .A2(new_n2163_), .B(new_n2166_), .ZN(new_n3034_));
  NAND2_X1   g2649(.A1(new_n1220_), .A2(new_n1630_), .ZN(new_n3035_));
  AOI21_X1   g2650(.A1(new_n3034_), .A2(new_n2170_), .B(new_n3035_), .ZN(\grant[46] ));
  OAI21_X1   g2651(.A1(new_n1450_), .A2(\priority[49] ), .B(new_n2171_), .ZN(new_n3037_));
  NOR3_X1    g2652(.A1(new_n3037_), .A2(new_n1225_), .A3(new_n1227_), .ZN(new_n3038_));
  OAI21_X1   g2653(.A1(new_n1239_), .A2(new_n3038_), .B(new_n1248_), .ZN(new_n3039_));
  AOI21_X1   g2654(.A1(new_n3039_), .A2(new_n2322_), .B(new_n2323_), .ZN(new_n3040_));
  OAI21_X1   g2655(.A1(new_n3040_), .A2(new_n1275_), .B(new_n1284_), .ZN(new_n3041_));
  AOI21_X1   g2656(.A1(new_n3041_), .A2(new_n2320_), .B(new_n2321_), .ZN(new_n3042_));
  OAI21_X1   g2657(.A1(new_n3042_), .A2(new_n1311_), .B(new_n1320_), .ZN(new_n3043_));
  AOI21_X1   g2658(.A1(new_n3043_), .A2(new_n2318_), .B(new_n2319_), .ZN(new_n3044_));
  OAI21_X1   g2659(.A1(new_n3044_), .A2(new_n1347_), .B(new_n1356_), .ZN(new_n3045_));
  AOI21_X1   g2660(.A1(new_n3045_), .A2(new_n2316_), .B(new_n2317_), .ZN(new_n3046_));
  OAI21_X1   g2661(.A1(new_n3046_), .A2(new_n1385_), .B(new_n2342_), .ZN(new_n3047_));
  AOI21_X1   g2662(.A1(new_n3047_), .A2(new_n2315_), .B(new_n2728_), .ZN(new_n3048_));
  OAI21_X1   g2663(.A1(new_n3048_), .A2(new_n438_), .B(new_n452_), .ZN(new_n3049_));
  AOI21_X1   g2664(.A1(new_n3049_), .A2(new_n2253_), .B(new_n2254_), .ZN(new_n3050_));
  OAI21_X1   g2665(.A1(new_n3050_), .A2(new_n494_), .B(new_n508_), .ZN(new_n3051_));
  NAND2_X1   g2666(.A1(new_n532_), .A2(new_n1817_), .ZN(new_n3052_));
  AOI21_X1   g2667(.A1(new_n3051_), .A2(new_n2251_), .B(new_n3052_), .ZN(\grant[47] ));
  AOI21_X1   g2668(.A1(new_n905_), .A2(\priority[49] ), .B(\priority[50] ), .ZN(new_n3054_));
  NOR4_X1    g2669(.A1(new_n542_), .A2(new_n1454_), .A3(new_n1456_), .A4(new_n3054_), .ZN(new_n3055_));
  OAI21_X1   g2670(.A1(new_n1464_), .A2(new_n3055_), .B(new_n1470_), .ZN(new_n3056_));
  AOI21_X1   g2671(.A1(new_n3056_), .A2(new_n2353_), .B(new_n2354_), .ZN(new_n3057_));
  OAI21_X1   g2672(.A1(new_n3057_), .A2(new_n1490_), .B(new_n1496_), .ZN(new_n3058_));
  AOI21_X1   g2673(.A1(new_n3058_), .A2(new_n2351_), .B(new_n2352_), .ZN(new_n3059_));
  OAI21_X1   g2674(.A1(new_n3059_), .A2(new_n1516_), .B(new_n1522_), .ZN(new_n3060_));
  AOI21_X1   g2675(.A1(new_n3060_), .A2(new_n2349_), .B(new_n2350_), .ZN(new_n3061_));
  OAI21_X1   g2676(.A1(new_n3061_), .A2(new_n1542_), .B(new_n1548_), .ZN(new_n3062_));
  AOI21_X1   g2677(.A1(new_n3062_), .A2(new_n2347_), .B(new_n2348_), .ZN(new_n3063_));
  OAI21_X1   g2678(.A1(new_n3063_), .A2(new_n1569_), .B(new_n2373_), .ZN(new_n3064_));
  AOI21_X1   g2679(.A1(new_n3064_), .A2(new_n2346_), .B(new_n2746_), .ZN(new_n3065_));
  OAI21_X1   g2680(.A1(new_n3065_), .A2(new_n827_), .B(new_n840_), .ZN(new_n3066_));
  AOI21_X1   g2681(.A1(new_n3066_), .A2(new_n2289_), .B(new_n2290_), .ZN(new_n3067_));
  OAI21_X1   g2682(.A1(new_n3067_), .A2(new_n877_), .B(new_n890_), .ZN(new_n3068_));
  NAND2_X1   g2683(.A1(new_n911_), .A2(new_n526_), .ZN(new_n3069_));
  AOI21_X1   g2684(.A1(new_n3068_), .A2(new_n2287_), .B(new_n3069_), .ZN(\grant[48] ));
  AOI21_X1   g2685(.A1(new_n1223_), .A2(\priority[50] ), .B(\priority[51] ), .ZN(new_n3071_));
  NOR4_X1    g2686(.A1(new_n919_), .A2(new_n1637_), .A3(new_n1639_), .A4(new_n3071_), .ZN(new_n3072_));
  OAI21_X1   g2687(.A1(new_n1647_), .A2(new_n3072_), .B(new_n1653_), .ZN(new_n3073_));
  AOI21_X1   g2688(.A1(new_n3073_), .A2(new_n2384_), .B(new_n2385_), .ZN(new_n3074_));
  OAI21_X1   g2689(.A1(new_n3074_), .A2(new_n1673_), .B(new_n1679_), .ZN(new_n3075_));
  AOI21_X1   g2690(.A1(new_n3075_), .A2(new_n2382_), .B(new_n2383_), .ZN(new_n3076_));
  OAI21_X1   g2691(.A1(new_n3076_), .A2(new_n1699_), .B(new_n1705_), .ZN(new_n3077_));
  AOI21_X1   g2692(.A1(new_n3077_), .A2(new_n2380_), .B(new_n2381_), .ZN(new_n3078_));
  OAI21_X1   g2693(.A1(new_n3078_), .A2(new_n1725_), .B(new_n1731_), .ZN(new_n3079_));
  AOI21_X1   g2694(.A1(new_n3079_), .A2(new_n2378_), .B(new_n2379_), .ZN(new_n3080_));
  OAI21_X1   g2695(.A1(new_n3080_), .A2(new_n1750_), .B(new_n2404_), .ZN(new_n3081_));
  AOI21_X1   g2696(.A1(new_n3081_), .A2(new_n2377_), .B(new_n2764_), .ZN(new_n3082_));
  OAI21_X1   g2697(.A1(new_n3082_), .A2(new_n1167_), .B(new_n1176_), .ZN(new_n3083_));
  AOI21_X1   g2698(.A1(new_n3083_), .A2(new_n2326_), .B(new_n2327_), .ZN(new_n3084_));
  OAI21_X1   g2699(.A1(new_n3084_), .A2(new_n1203_), .B(new_n1212_), .ZN(new_n3085_));
  NAND2_X1   g2700(.A1(new_n1228_), .A2(new_n905_), .ZN(new_n3086_));
  AOI21_X1   g2701(.A1(new_n3085_), .A2(new_n2324_), .B(new_n3086_), .ZN(\grant[49] ));
  NOR4_X1    g2702(.A1(new_n1234_), .A2(new_n1982_), .A3(new_n1827_), .A4(new_n1824_), .ZN(new_n3088_));
  OAI21_X1   g2703(.A1(new_n1835_), .A2(new_n3088_), .B(new_n1842_), .ZN(new_n3089_));
  AOI21_X1   g2704(.A1(new_n3089_), .A2(new_n2415_), .B(new_n2416_), .ZN(new_n3090_));
  OAI21_X1   g2705(.A1(new_n3090_), .A2(new_n1863_), .B(new_n1870_), .ZN(new_n3091_));
  AOI21_X1   g2706(.A1(new_n3091_), .A2(new_n2413_), .B(new_n2414_), .ZN(new_n3092_));
  OAI21_X1   g2707(.A1(new_n3092_), .A2(new_n1891_), .B(new_n1898_), .ZN(new_n3093_));
  AOI21_X1   g2708(.A1(new_n3093_), .A2(new_n2411_), .B(new_n2412_), .ZN(new_n3094_));
  OAI21_X1   g2709(.A1(new_n3094_), .A2(new_n1919_), .B(new_n1926_), .ZN(new_n3095_));
  AOI21_X1   g2710(.A1(new_n3095_), .A2(new_n2409_), .B(new_n2410_), .ZN(new_n3096_));
  OAI21_X1   g2711(.A1(new_n3096_), .A2(new_n1945_), .B(new_n2434_), .ZN(new_n3097_));
  AOI21_X1   g2712(.A1(new_n3097_), .A2(new_n2408_), .B(new_n2782_), .ZN(new_n3098_));
  OAI21_X1   g2713(.A1(new_n3098_), .A2(new_n1412_), .B(new_n1418_), .ZN(new_n3099_));
  AOI21_X1   g2714(.A1(new_n3099_), .A2(new_n2357_), .B(new_n2358_), .ZN(new_n3100_));
  OAI21_X1   g2715(.A1(new_n3100_), .A2(new_n1438_), .B(new_n1444_), .ZN(new_n3101_));
  NAND2_X1   g2716(.A1(new_n1453_), .A2(new_n1223_), .ZN(new_n3102_));
  AOI21_X1   g2717(.A1(new_n3101_), .A2(new_n2355_), .B(new_n3102_), .ZN(\grant[50] ));
  NOR4_X1    g2718(.A1(new_n1461_), .A2(new_n548_), .A3(new_n1984_), .A4(new_n2080_), .ZN(new_n3104_));
  OAI21_X1   g2719(.A1(new_n1989_), .A2(new_n3104_), .B(new_n1992_), .ZN(new_n3105_));
  AOI21_X1   g2720(.A1(new_n3105_), .A2(new_n2445_), .B(new_n2446_), .ZN(new_n3106_));
  OAI21_X1   g2721(.A1(new_n3106_), .A2(new_n2003_), .B(new_n2006_), .ZN(new_n3107_));
  AOI21_X1   g2722(.A1(new_n3107_), .A2(new_n2443_), .B(new_n2444_), .ZN(new_n3108_));
  OAI21_X1   g2723(.A1(new_n3108_), .A2(new_n2017_), .B(new_n2020_), .ZN(new_n3109_));
  AOI21_X1   g2724(.A1(new_n3109_), .A2(new_n2441_), .B(new_n2442_), .ZN(new_n3110_));
  OAI21_X1   g2725(.A1(new_n3110_), .A2(new_n2031_), .B(new_n2034_), .ZN(new_n3111_));
  AOI21_X1   g2726(.A1(new_n3111_), .A2(new_n2439_), .B(new_n2440_), .ZN(new_n3112_));
  OAI21_X1   g2727(.A1(new_n3112_), .A2(new_n2048_), .B(new_n2464_), .ZN(new_n3113_));
  AOI21_X1   g2728(.A1(new_n3113_), .A2(new_n2438_), .B(new_n2799_), .ZN(new_n3114_));
  OAI21_X1   g2729(.A1(new_n3114_), .A2(new_n1595_), .B(new_n1601_), .ZN(new_n3115_));
  AOI21_X1   g2730(.A1(new_n3115_), .A2(new_n2388_), .B(new_n2389_), .ZN(new_n3116_));
  OAI21_X1   g2731(.A1(new_n3116_), .A2(new_n1621_), .B(new_n1627_), .ZN(new_n3117_));
  NAND2_X1   g2732(.A1(new_n1636_), .A2(new_n540_), .ZN(new_n3118_));
  AOI21_X1   g2733(.A1(new_n3117_), .A2(new_n2386_), .B(new_n3118_), .ZN(\grant[51] ));
  NOR4_X1    g2734(.A1(new_n1644_), .A2(new_n925_), .A3(new_n2082_), .A4(new_n2176_), .ZN(new_n3120_));
  OAI21_X1   g2735(.A1(new_n2086_), .A2(new_n3120_), .B(new_n2089_), .ZN(new_n3121_));
  AOI21_X1   g2736(.A1(new_n3121_), .A2(new_n2475_), .B(new_n2476_), .ZN(new_n3122_));
  OAI21_X1   g2737(.A1(new_n3122_), .A2(new_n2098_), .B(new_n2101_), .ZN(new_n3123_));
  AOI21_X1   g2738(.A1(new_n3123_), .A2(new_n2473_), .B(new_n2474_), .ZN(new_n3124_));
  OAI21_X1   g2739(.A1(new_n3124_), .A2(new_n2110_), .B(new_n2113_), .ZN(new_n3125_));
  AOI21_X1   g2740(.A1(new_n3125_), .A2(new_n2471_), .B(new_n2472_), .ZN(new_n3126_));
  OAI21_X1   g2741(.A1(new_n3126_), .A2(new_n2122_), .B(new_n2125_), .ZN(new_n3127_));
  AOI21_X1   g2742(.A1(new_n3127_), .A2(new_n2469_), .B(new_n2470_), .ZN(new_n3128_));
  OAI21_X1   g2743(.A1(new_n3128_), .A2(new_n2139_), .B(new_n2494_), .ZN(new_n3129_));
  AOI21_X1   g2744(.A1(new_n3129_), .A2(new_n2468_), .B(new_n2816_), .ZN(new_n3130_));
  OAI21_X1   g2745(.A1(new_n3130_), .A2(new_n1779_), .B(new_n1786_), .ZN(new_n3131_));
  AOI21_X1   g2746(.A1(new_n3131_), .A2(new_n2419_), .B(new_n2420_), .ZN(new_n3132_));
  OAI21_X1   g2747(.A1(new_n3132_), .A2(new_n1807_), .B(new_n1814_), .ZN(new_n3133_));
  NAND2_X1   g2748(.A1(new_n1823_), .A2(new_n917_), .ZN(new_n3134_));
  AOI21_X1   g2749(.A1(new_n3133_), .A2(new_n2417_), .B(new_n3134_), .ZN(\grant[52] ));
  OAI21_X1   g2750(.A1(new_n544_), .A2(\priority[55] ), .B(new_n1826_), .ZN(new_n3136_));
  NOR3_X1    g2751(.A1(new_n3136_), .A2(new_n1832_), .A3(new_n2179_), .ZN(new_n3137_));
  OAI21_X1   g2752(.A1(new_n2183_), .A2(new_n3137_), .B(new_n2187_), .ZN(new_n3138_));
  AOI21_X1   g2753(.A1(new_n3138_), .A2(new_n2505_), .B(new_n2506_), .ZN(new_n3139_));
  OAI21_X1   g2754(.A1(new_n3139_), .A2(new_n2197_), .B(new_n2201_), .ZN(new_n3140_));
  AOI21_X1   g2755(.A1(new_n3140_), .A2(new_n2503_), .B(new_n2504_), .ZN(new_n3141_));
  OAI21_X1   g2756(.A1(new_n3141_), .A2(new_n2211_), .B(new_n2215_), .ZN(new_n3142_));
  AOI21_X1   g2757(.A1(new_n3142_), .A2(new_n2501_), .B(new_n2502_), .ZN(new_n3143_));
  OAI21_X1   g2758(.A1(new_n3143_), .A2(new_n2225_), .B(new_n2229_), .ZN(new_n3144_));
  AOI21_X1   g2759(.A1(new_n3144_), .A2(new_n2499_), .B(new_n2500_), .ZN(new_n3145_));
  OAI21_X1   g2760(.A1(new_n3145_), .A2(new_n2239_), .B(new_n2525_), .ZN(new_n3146_));
  AOI21_X1   g2761(.A1(new_n3146_), .A2(new_n2498_), .B(new_n2833_), .ZN(new_n3147_));
  OAI21_X1   g2762(.A1(new_n3147_), .A2(new_n1961_), .B(new_n1964_), .ZN(new_n3148_));
  AOI21_X1   g2763(.A1(new_n3148_), .A2(new_n2449_), .B(new_n2450_), .ZN(new_n3149_));
  OAI21_X1   g2764(.A1(new_n3149_), .A2(new_n1975_), .B(new_n1978_), .ZN(new_n3150_));
  NAND2_X1   g2765(.A1(new_n546_), .A2(new_n1232_), .ZN(new_n3151_));
  AOI21_X1   g2766(.A1(new_n3150_), .A2(new_n2447_), .B(new_n3151_), .ZN(\grant[53] ));
  AOI21_X1   g2767(.A1(new_n1642_), .A2(\priority[55] ), .B(\priority[56] ), .ZN(new_n3153_));
  NOR4_X1    g2768(.A1(new_n556_), .A2(new_n558_), .A3(new_n562_), .A4(new_n3153_), .ZN(new_n3154_));
  OAI21_X1   g2769(.A1(new_n579_), .A2(new_n3154_), .B(new_n592_), .ZN(new_n3155_));
  AOI21_X1   g2770(.A1(new_n3155_), .A2(new_n607_), .B(new_n621_), .ZN(new_n3156_));
  OAI21_X1   g2771(.A1(new_n3156_), .A2(new_n635_), .B(new_n648_), .ZN(new_n3157_));
  AOI21_X1   g2772(.A1(new_n3157_), .A2(new_n663_), .B(new_n677_), .ZN(new_n3158_));
  OAI21_X1   g2773(.A1(new_n3158_), .A2(new_n691_), .B(new_n704_), .ZN(new_n3159_));
  AOI21_X1   g2774(.A1(new_n3159_), .A2(new_n719_), .B(new_n733_), .ZN(new_n3160_));
  OAI21_X1   g2775(.A1(new_n3160_), .A2(new_n747_), .B(new_n760_), .ZN(new_n3161_));
  AOI21_X1   g2776(.A1(new_n3161_), .A2(new_n775_), .B(new_n2530_), .ZN(new_n3162_));
  OAI21_X1   g2777(.A1(new_n3162_), .A2(new_n2275_), .B(new_n2545_), .ZN(new_n3163_));
  AOI21_X1   g2778(.A1(new_n3163_), .A2(new_n2529_), .B(new_n2851_), .ZN(new_n3164_));
  OAI21_X1   g2779(.A1(new_n3164_), .A2(new_n2062_), .B(new_n2065_), .ZN(new_n3165_));
  AOI21_X1   g2780(.A1(new_n3165_), .A2(new_n2479_), .B(new_n2480_), .ZN(new_n3166_));
  OAI21_X1   g2781(.A1(new_n3166_), .A2(new_n2074_), .B(new_n2077_), .ZN(new_n3167_));
  NAND2_X1   g2782(.A1(new_n923_), .A2(new_n1459_), .ZN(new_n3168_));
  AOI21_X1   g2783(.A1(new_n3167_), .A2(new_n2477_), .B(new_n3168_), .ZN(\grant[54] ));
  AOI21_X1   g2784(.A1(new_n1830_), .A2(\priority[56] ), .B(\priority[57] ), .ZN(new_n3170_));
  NOR4_X1    g2785(.A1(new_n932_), .A2(new_n934_), .A3(new_n938_), .A4(new_n3170_), .ZN(new_n3171_));
  OAI21_X1   g2786(.A1(new_n953_), .A2(new_n3171_), .B(new_n965_), .ZN(new_n3172_));
  AOI21_X1   g2787(.A1(new_n3172_), .A2(new_n978_), .B(new_n991_), .ZN(new_n3173_));
  OAI21_X1   g2788(.A1(new_n3173_), .A2(new_n1003_), .B(new_n1015_), .ZN(new_n3174_));
  AOI21_X1   g2789(.A1(new_n3174_), .A2(new_n1028_), .B(new_n1041_), .ZN(new_n3175_));
  OAI21_X1   g2790(.A1(new_n3175_), .A2(new_n1053_), .B(new_n1065_), .ZN(new_n3176_));
  AOI21_X1   g2791(.A1(new_n3176_), .A2(new_n1078_), .B(new_n1091_), .ZN(new_n3177_));
  OAI21_X1   g2792(.A1(new_n3177_), .A2(new_n1103_), .B(new_n1115_), .ZN(new_n3178_));
  AOI21_X1   g2793(.A1(new_n3178_), .A2(new_n1128_), .B(new_n2550_), .ZN(new_n3179_));
  OAI21_X1   g2794(.A1(new_n3179_), .A2(new_n2311_), .B(new_n2565_), .ZN(new_n3180_));
  AOI21_X1   g2795(.A1(new_n3180_), .A2(new_n2549_), .B(new_n2869_), .ZN(new_n3181_));
  OAI21_X1   g2796(.A1(new_n3181_), .A2(new_n2155_), .B(new_n2159_), .ZN(new_n3182_));
  AOI21_X1   g2797(.A1(new_n3182_), .A2(new_n2509_), .B(new_n2510_), .ZN(new_n3183_));
  OAI21_X1   g2798(.A1(new_n3183_), .A2(new_n2169_), .B(new_n2173_), .ZN(new_n3184_));
  NAND2_X1   g2799(.A1(new_n1237_), .A2(new_n1642_), .ZN(new_n3185_));
  AOI21_X1   g2800(.A1(new_n3184_), .A2(new_n2507_), .B(new_n3185_), .ZN(\grant[55] ));
  OAI21_X1   g2801(.A1(new_n1462_), .A2(\priority[58] ), .B(new_n2178_), .ZN(new_n3187_));
  NOR3_X1    g2802(.A1(new_n3187_), .A2(new_n1243_), .A3(new_n1245_), .ZN(new_n3188_));
  OAI21_X1   g2803(.A1(new_n1258_), .A2(new_n3188_), .B(new_n1266_), .ZN(new_n3189_));
  AOI21_X1   g2804(.A1(new_n3189_), .A2(new_n1276_), .B(new_n1285_), .ZN(new_n3190_));
  OAI21_X1   g2805(.A1(new_n3190_), .A2(new_n1294_), .B(new_n1302_), .ZN(new_n3191_));
  AOI21_X1   g2806(.A1(new_n3191_), .A2(new_n1312_), .B(new_n1321_), .ZN(new_n3192_));
  OAI21_X1   g2807(.A1(new_n3192_), .A2(new_n1330_), .B(new_n1338_), .ZN(new_n3193_));
  AOI21_X1   g2808(.A1(new_n3193_), .A2(new_n1348_), .B(new_n1357_), .ZN(new_n3194_));
  OAI21_X1   g2809(.A1(new_n3194_), .A2(new_n1366_), .B(new_n1374_), .ZN(new_n3195_));
  AOI21_X1   g2810(.A1(new_n3195_), .A2(new_n1386_), .B(new_n2569_), .ZN(new_n3196_));
  OAI21_X1   g2811(.A1(new_n3196_), .A2(new_n411_), .B(new_n424_), .ZN(new_n3197_));
  AOI21_X1   g2812(.A1(new_n3197_), .A2(new_n439_), .B(new_n453_), .ZN(new_n3198_));
  OAI21_X1   g2813(.A1(new_n3198_), .A2(new_n467_), .B(new_n480_), .ZN(new_n3199_));
  AOI21_X1   g2814(.A1(new_n3199_), .A2(new_n495_), .B(new_n509_), .ZN(new_n3200_));
  OAI21_X1   g2815(.A1(new_n3200_), .A2(new_n523_), .B(new_n536_), .ZN(new_n3201_));
  NAND2_X1   g2816(.A1(new_n560_), .A2(new_n1830_), .ZN(new_n3202_));
  AOI21_X1   g2817(.A1(new_n3201_), .A2(new_n551_), .B(new_n3202_), .ZN(\grant[56] ));
  AOI21_X1   g2818(.A1(new_n930_), .A2(\priority[58] ), .B(\priority[59] ), .ZN(new_n3204_));
  NOR4_X1    g2819(.A1(new_n571_), .A2(new_n1467_), .A3(new_n1469_), .A4(new_n3204_), .ZN(new_n3205_));
  OAI21_X1   g2820(.A1(new_n1478_), .A2(new_n3205_), .B(new_n1483_), .ZN(new_n3206_));
  AOI21_X1   g2821(.A1(new_n3206_), .A2(new_n1491_), .B(new_n1497_), .ZN(new_n3207_));
  OAI21_X1   g2822(.A1(new_n3207_), .A2(new_n1504_), .B(new_n1509_), .ZN(new_n3208_));
  AOI21_X1   g2823(.A1(new_n3208_), .A2(new_n1517_), .B(new_n1523_), .ZN(new_n3209_));
  OAI21_X1   g2824(.A1(new_n3209_), .A2(new_n1530_), .B(new_n1535_), .ZN(new_n3210_));
  AOI21_X1   g2825(.A1(new_n3210_), .A2(new_n1543_), .B(new_n1549_), .ZN(new_n3211_));
  OAI21_X1   g2826(.A1(new_n3211_), .A2(new_n1556_), .B(new_n1561_), .ZN(new_n3212_));
  AOI21_X1   g2827(.A1(new_n3212_), .A2(new_n1570_), .B(new_n2587_), .ZN(new_n3213_));
  OAI21_X1   g2828(.A1(new_n3213_), .A2(new_n803_), .B(new_n815_), .ZN(new_n3214_));
  AOI21_X1   g2829(.A1(new_n3214_), .A2(new_n828_), .B(new_n841_), .ZN(new_n3215_));
  OAI21_X1   g2830(.A1(new_n3215_), .A2(new_n853_), .B(new_n865_), .ZN(new_n3216_));
  AOI21_X1   g2831(.A1(new_n3216_), .A2(new_n878_), .B(new_n891_), .ZN(new_n3217_));
  OAI21_X1   g2832(.A1(new_n3217_), .A2(new_n903_), .B(new_n915_), .ZN(new_n3218_));
  NAND2_X1   g2833(.A1(new_n936_), .A2(new_n554_), .ZN(new_n3219_));
  AOI21_X1   g2834(.A1(new_n3218_), .A2(new_n928_), .B(new_n3219_), .ZN(\grant[57] ));
  AOI21_X1   g2835(.A1(new_n1241_), .A2(\priority[59] ), .B(\priority[60] ), .ZN(new_n3221_));
  NOR4_X1    g2836(.A1(new_n945_), .A2(new_n1650_), .A3(new_n1652_), .A4(new_n3221_), .ZN(new_n3222_));
  OAI21_X1   g2837(.A1(new_n1661_), .A2(new_n3222_), .B(new_n1666_), .ZN(new_n3223_));
  AOI21_X1   g2838(.A1(new_n3223_), .A2(new_n1674_), .B(new_n1680_), .ZN(new_n3224_));
  OAI21_X1   g2839(.A1(new_n3224_), .A2(new_n1687_), .B(new_n1692_), .ZN(new_n3225_));
  AOI21_X1   g2840(.A1(new_n3225_), .A2(new_n1700_), .B(new_n1706_), .ZN(new_n3226_));
  OAI21_X1   g2841(.A1(new_n3226_), .A2(new_n1713_), .B(new_n1718_), .ZN(new_n3227_));
  AOI21_X1   g2842(.A1(new_n3227_), .A2(new_n1726_), .B(new_n1732_), .ZN(new_n3228_));
  OAI21_X1   g2843(.A1(new_n3228_), .A2(new_n1739_), .B(new_n1744_), .ZN(new_n3229_));
  AOI21_X1   g2844(.A1(new_n3229_), .A2(new_n1751_), .B(new_n2605_), .ZN(new_n3230_));
  OAI21_X1   g2845(.A1(new_n3230_), .A2(new_n1150_), .B(new_n1158_), .ZN(new_n3231_));
  AOI21_X1   g2846(.A1(new_n3231_), .A2(new_n1168_), .B(new_n1177_), .ZN(new_n3232_));
  OAI21_X1   g2847(.A1(new_n3232_), .A2(new_n1186_), .B(new_n1194_), .ZN(new_n3233_));
  AOI21_X1   g2848(.A1(new_n3233_), .A2(new_n1204_), .B(new_n1213_), .ZN(new_n3234_));
  OAI21_X1   g2849(.A1(new_n3234_), .A2(new_n1222_), .B(new_n1230_), .ZN(new_n3235_));
  NAND2_X1   g2850(.A1(new_n1246_), .A2(new_n930_), .ZN(new_n3236_));
  AOI21_X1   g2851(.A1(new_n3235_), .A2(new_n1240_), .B(new_n3236_), .ZN(\grant[58] ));
  NOR4_X1    g2852(.A1(new_n1253_), .A2(new_n1988_), .A3(new_n1841_), .A4(new_n1838_), .ZN(new_n3238_));
  OAI21_X1   g2853(.A1(new_n1850_), .A2(new_n3238_), .B(new_n1856_), .ZN(new_n3239_));
  AOI21_X1   g2854(.A1(new_n3239_), .A2(new_n1864_), .B(new_n1871_), .ZN(new_n3240_));
  OAI21_X1   g2855(.A1(new_n3240_), .A2(new_n1878_), .B(new_n1884_), .ZN(new_n3241_));
  AOI21_X1   g2856(.A1(new_n3241_), .A2(new_n1892_), .B(new_n1899_), .ZN(new_n3242_));
  OAI21_X1   g2857(.A1(new_n3242_), .A2(new_n1906_), .B(new_n1912_), .ZN(new_n3243_));
  AOI21_X1   g2858(.A1(new_n3243_), .A2(new_n1920_), .B(new_n1927_), .ZN(new_n3244_));
  OAI21_X1   g2859(.A1(new_n3244_), .A2(new_n1934_), .B(new_n1939_), .ZN(new_n3245_));
  AOI21_X1   g2860(.A1(new_n3245_), .A2(new_n1946_), .B(new_n2623_), .ZN(new_n3246_));
  OAI21_X1   g2861(.A1(new_n3246_), .A2(new_n1400_), .B(new_n1405_), .ZN(new_n3247_));
  AOI21_X1   g2862(.A1(new_n3247_), .A2(new_n1413_), .B(new_n1419_), .ZN(new_n3248_));
  OAI21_X1   g2863(.A1(new_n3248_), .A2(new_n1426_), .B(new_n1431_), .ZN(new_n3249_));
  AOI21_X1   g2864(.A1(new_n3249_), .A2(new_n1439_), .B(new_n1445_), .ZN(new_n3250_));
  OAI21_X1   g2865(.A1(new_n3250_), .A2(new_n1452_), .B(new_n1457_), .ZN(new_n3251_));
  NAND2_X1   g2866(.A1(new_n1466_), .A2(new_n1241_), .ZN(new_n3252_));
  AOI21_X1   g2867(.A1(new_n3251_), .A2(new_n1465_), .B(new_n3252_), .ZN(\grant[59] ));
  NOR4_X1    g2868(.A1(new_n1475_), .A2(new_n577_), .A3(new_n1991_), .A4(new_n2085_), .ZN(new_n3254_));
  OAI21_X1   g2869(.A1(new_n1997_), .A2(new_n3254_), .B(new_n1999_), .ZN(new_n3255_));
  AOI21_X1   g2870(.A1(new_n3255_), .A2(new_n2004_), .B(new_n2007_), .ZN(new_n3256_));
  OAI21_X1   g2871(.A1(new_n3256_), .A2(new_n2011_), .B(new_n2013_), .ZN(new_n3257_));
  AOI21_X1   g2872(.A1(new_n3257_), .A2(new_n2018_), .B(new_n2021_), .ZN(new_n3258_));
  OAI21_X1   g2873(.A1(new_n3258_), .A2(new_n2025_), .B(new_n2027_), .ZN(new_n3259_));
  AOI21_X1   g2874(.A1(new_n3259_), .A2(new_n2032_), .B(new_n2035_), .ZN(new_n3260_));
  OAI21_X1   g2875(.A1(new_n3260_), .A2(new_n2039_), .B(new_n2041_), .ZN(new_n3261_));
  AOI21_X1   g2876(.A1(new_n3261_), .A2(new_n2049_), .B(new_n2640_), .ZN(new_n3262_));
  OAI21_X1   g2877(.A1(new_n3262_), .A2(new_n1583_), .B(new_n1588_), .ZN(new_n3263_));
  AOI21_X1   g2878(.A1(new_n3263_), .A2(new_n1596_), .B(new_n1602_), .ZN(new_n3264_));
  OAI21_X1   g2879(.A1(new_n3264_), .A2(new_n1609_), .B(new_n1614_), .ZN(new_n3265_));
  AOI21_X1   g2880(.A1(new_n3265_), .A2(new_n1622_), .B(new_n1628_), .ZN(new_n3266_));
  OAI21_X1   g2881(.A1(new_n3266_), .A2(new_n1635_), .B(new_n1640_), .ZN(new_n3267_));
  NAND2_X1   g2882(.A1(new_n1649_), .A2(new_n569_), .ZN(new_n3268_));
  AOI21_X1   g2883(.A1(new_n3267_), .A2(new_n1648_), .B(new_n3268_), .ZN(\grant[60] ));
  NOR4_X1    g2884(.A1(new_n1658_), .A2(new_n951_), .A3(new_n2088_), .A4(new_n2182_), .ZN(new_n3270_));
  OAI21_X1   g2885(.A1(new_n2093_), .A2(new_n3270_), .B(new_n2095_), .ZN(new_n3271_));
  AOI21_X1   g2886(.A1(new_n3271_), .A2(new_n2099_), .B(new_n2102_), .ZN(new_n3272_));
  OAI21_X1   g2887(.A1(new_n3272_), .A2(new_n2105_), .B(new_n2107_), .ZN(new_n3273_));
  AOI21_X1   g2888(.A1(new_n3273_), .A2(new_n2111_), .B(new_n2114_), .ZN(new_n3274_));
  OAI21_X1   g2889(.A1(new_n3274_), .A2(new_n2117_), .B(new_n2119_), .ZN(new_n3275_));
  AOI21_X1   g2890(.A1(new_n3275_), .A2(new_n2123_), .B(new_n2126_), .ZN(new_n3276_));
  OAI21_X1   g2891(.A1(new_n3276_), .A2(new_n2129_), .B(new_n2132_), .ZN(new_n3277_));
  AOI21_X1   g2892(.A1(new_n3277_), .A2(new_n2140_), .B(new_n2657_), .ZN(new_n3278_));
  OAI21_X1   g2893(.A1(new_n3278_), .A2(new_n1766_), .B(new_n1772_), .ZN(new_n3279_));
  AOI21_X1   g2894(.A1(new_n3279_), .A2(new_n1780_), .B(new_n1787_), .ZN(new_n3280_));
  OAI21_X1   g2895(.A1(new_n3280_), .A2(new_n1794_), .B(new_n1800_), .ZN(new_n3281_));
  AOI21_X1   g2896(.A1(new_n3281_), .A2(new_n1808_), .B(new_n1815_), .ZN(new_n3282_));
  OAI21_X1   g2897(.A1(new_n3282_), .A2(new_n1822_), .B(new_n1828_), .ZN(new_n3283_));
  NAND2_X1   g2898(.A1(new_n1837_), .A2(new_n943_), .ZN(new_n3284_));
  AOI21_X1   g2899(.A1(new_n3283_), .A2(new_n1836_), .B(new_n3284_), .ZN(\grant[61] ));
  OAI21_X1   g2900(.A1(new_n573_), .A2(\priority[64] ), .B(new_n1840_), .ZN(new_n3286_));
  NOR3_X1    g2901(.A1(new_n3286_), .A2(new_n1847_), .A3(new_n2186_), .ZN(new_n3287_));
  OAI21_X1   g2902(.A1(new_n2191_), .A2(new_n3287_), .B(new_n2194_), .ZN(new_n3288_));
  AOI21_X1   g2903(.A1(new_n3288_), .A2(new_n2198_), .B(new_n2202_), .ZN(new_n3289_));
  OAI21_X1   g2904(.A1(new_n3289_), .A2(new_n2205_), .B(new_n2208_), .ZN(new_n3290_));
  AOI21_X1   g2905(.A1(new_n3290_), .A2(new_n2212_), .B(new_n2216_), .ZN(new_n3291_));
  OAI21_X1   g2906(.A1(new_n3291_), .A2(new_n2219_), .B(new_n2222_), .ZN(new_n3292_));
  AOI21_X1   g2907(.A1(new_n3292_), .A2(new_n2226_), .B(new_n2230_), .ZN(new_n3293_));
  OAI21_X1   g2908(.A1(new_n3293_), .A2(new_n2233_), .B(new_n2235_), .ZN(new_n3294_));
  AOI21_X1   g2909(.A1(new_n3294_), .A2(new_n2240_), .B(new_n2674_), .ZN(new_n3295_));
  OAI21_X1   g2910(.A1(new_n3295_), .A2(new_n1955_), .B(new_n1957_), .ZN(new_n3296_));
  AOI21_X1   g2911(.A1(new_n3296_), .A2(new_n1962_), .B(new_n1965_), .ZN(new_n3297_));
  OAI21_X1   g2912(.A1(new_n3297_), .A2(new_n1969_), .B(new_n1971_), .ZN(new_n3298_));
  AOI21_X1   g2913(.A1(new_n3298_), .A2(new_n1976_), .B(new_n1979_), .ZN(new_n3299_));
  OAI21_X1   g2914(.A1(new_n3299_), .A2(new_n1983_), .B(new_n1985_), .ZN(new_n3300_));
  NAND2_X1   g2915(.A1(new_n575_), .A2(new_n1251_), .ZN(new_n3301_));
  AOI21_X1   g2916(.A1(new_n3300_), .A2(new_n1990_), .B(new_n3301_), .ZN(\grant[62] ));
  AOI21_X1   g2917(.A1(new_n1656_), .A2(\priority[64] ), .B(\priority[65] ), .ZN(new_n3303_));
  NOR4_X1    g2918(.A1(new_n584_), .A2(new_n586_), .A3(new_n590_), .A4(new_n3303_), .ZN(new_n3304_));
  OAI21_X1   g2919(.A1(new_n606_), .A2(new_n3304_), .B(new_n620_), .ZN(new_n3305_));
  AOI21_X1   g2920(.A1(new_n3305_), .A2(new_n2247_), .B(new_n2248_), .ZN(new_n3306_));
  OAI21_X1   g2921(.A1(new_n3306_), .A2(new_n662_), .B(new_n676_), .ZN(new_n3307_));
  AOI21_X1   g2922(.A1(new_n3307_), .A2(new_n2245_), .B(new_n2246_), .ZN(new_n3308_));
  OAI21_X1   g2923(.A1(new_n3308_), .A2(new_n718_), .B(new_n732_), .ZN(new_n3309_));
  AOI21_X1   g2924(.A1(new_n3309_), .A2(new_n2243_), .B(new_n2244_), .ZN(new_n3310_));
  OAI21_X1   g2925(.A1(new_n3310_), .A2(new_n774_), .B(new_n2270_), .ZN(new_n3311_));
  AOI21_X1   g2926(.A1(new_n3311_), .A2(new_n2276_), .B(new_n2692_), .ZN(new_n3312_));
  OAI21_X1   g2927(.A1(new_n3312_), .A2(new_n2057_), .B(new_n2059_), .ZN(new_n3313_));
  AOI21_X1   g2928(.A1(new_n3313_), .A2(new_n2063_), .B(new_n2066_), .ZN(new_n3314_));
  OAI21_X1   g2929(.A1(new_n3314_), .A2(new_n2069_), .B(new_n2071_), .ZN(new_n3315_));
  AOI21_X1   g2930(.A1(new_n3315_), .A2(new_n2075_), .B(new_n2078_), .ZN(new_n3316_));
  OAI21_X1   g2931(.A1(new_n3316_), .A2(new_n2081_), .B(new_n2083_), .ZN(new_n3317_));
  NAND2_X1   g2932(.A1(new_n949_), .A2(new_n1473_), .ZN(new_n3318_));
  AOI21_X1   g2933(.A1(new_n3317_), .A2(new_n2087_), .B(new_n3318_), .ZN(\grant[63] ));
  AOI21_X1   g2934(.A1(new_n1845_), .A2(\priority[65] ), .B(\priority[66] ), .ZN(new_n3320_));
  NOR4_X1    g2935(.A1(new_n957_), .A2(new_n959_), .A3(new_n963_), .A4(new_n3320_), .ZN(new_n3321_));
  OAI21_X1   g2936(.A1(new_n977_), .A2(new_n3321_), .B(new_n990_), .ZN(new_n3322_));
  AOI21_X1   g2937(.A1(new_n3322_), .A2(new_n2283_), .B(new_n2284_), .ZN(new_n3323_));
  OAI21_X1   g2938(.A1(new_n3323_), .A2(new_n1027_), .B(new_n1040_), .ZN(new_n3324_));
  AOI21_X1   g2939(.A1(new_n3324_), .A2(new_n2281_), .B(new_n2282_), .ZN(new_n3325_));
  OAI21_X1   g2940(.A1(new_n3325_), .A2(new_n1077_), .B(new_n1090_), .ZN(new_n3326_));
  AOI21_X1   g2941(.A1(new_n3326_), .A2(new_n2279_), .B(new_n2280_), .ZN(new_n3327_));
  OAI21_X1   g2942(.A1(new_n3327_), .A2(new_n1127_), .B(new_n2306_), .ZN(new_n3328_));
  AOI21_X1   g2943(.A1(new_n3328_), .A2(new_n2312_), .B(new_n2710_), .ZN(new_n3329_));
  OAI21_X1   g2944(.A1(new_n3329_), .A2(new_n2149_), .B(new_n2152_), .ZN(new_n3330_));
  AOI21_X1   g2945(.A1(new_n3330_), .A2(new_n2156_), .B(new_n2160_), .ZN(new_n3331_));
  OAI21_X1   g2946(.A1(new_n3331_), .A2(new_n2163_), .B(new_n2166_), .ZN(new_n3332_));
  AOI21_X1   g2947(.A1(new_n3332_), .A2(new_n2170_), .B(new_n2174_), .ZN(new_n3333_));
  OAI21_X1   g2948(.A1(new_n3333_), .A2(new_n2177_), .B(new_n2180_), .ZN(new_n3334_));
  NAND2_X1   g2949(.A1(new_n1256_), .A2(new_n1656_), .ZN(new_n3335_));
  AOI21_X1   g2950(.A1(new_n3334_), .A2(new_n2184_), .B(new_n3335_), .ZN(\grant[64] ));
  OAI21_X1   g2951(.A1(new_n1476_), .A2(\priority[67] ), .B(new_n2185_), .ZN(new_n3337_));
  NOR3_X1    g2952(.A1(new_n3337_), .A2(new_n1261_), .A3(new_n1263_), .ZN(new_n3338_));
  OAI21_X1   g2953(.A1(new_n1275_), .A2(new_n3338_), .B(new_n1284_), .ZN(new_n3339_));
  AOI21_X1   g2954(.A1(new_n3339_), .A2(new_n2320_), .B(new_n2321_), .ZN(new_n3340_));
  OAI21_X1   g2955(.A1(new_n3340_), .A2(new_n1311_), .B(new_n1320_), .ZN(new_n3341_));
  AOI21_X1   g2956(.A1(new_n3341_), .A2(new_n2318_), .B(new_n2319_), .ZN(new_n3342_));
  OAI21_X1   g2957(.A1(new_n3342_), .A2(new_n1347_), .B(new_n1356_), .ZN(new_n3343_));
  AOI21_X1   g2958(.A1(new_n3343_), .A2(new_n2316_), .B(new_n2317_), .ZN(new_n3344_));
  OAI21_X1   g2959(.A1(new_n3344_), .A2(new_n1385_), .B(new_n2342_), .ZN(new_n3345_));
  AOI21_X1   g2960(.A1(new_n3345_), .A2(new_n2315_), .B(new_n2728_), .ZN(new_n3346_));
  OAI21_X1   g2961(.A1(new_n3346_), .A2(new_n438_), .B(new_n452_), .ZN(new_n3347_));
  AOI21_X1   g2962(.A1(new_n3347_), .A2(new_n2253_), .B(new_n2254_), .ZN(new_n3348_));
  OAI21_X1   g2963(.A1(new_n3348_), .A2(new_n494_), .B(new_n508_), .ZN(new_n3349_));
  AOI21_X1   g2964(.A1(new_n3349_), .A2(new_n2251_), .B(new_n2252_), .ZN(new_n3350_));
  OAI21_X1   g2965(.A1(new_n3350_), .A2(new_n550_), .B(new_n564_), .ZN(new_n3351_));
  NAND2_X1   g2966(.A1(new_n588_), .A2(new_n1845_), .ZN(new_n3352_));
  AOI21_X1   g2967(.A1(new_n3351_), .A2(new_n2249_), .B(new_n3352_), .ZN(\grant[65] ));
  AOI21_X1   g2968(.A1(new_n955_), .A2(\priority[67] ), .B(\priority[68] ), .ZN(new_n3354_));
  NOR4_X1    g2969(.A1(new_n598_), .A2(new_n1480_), .A3(new_n1482_), .A4(new_n3354_), .ZN(new_n3355_));
  OAI21_X1   g2970(.A1(new_n1490_), .A2(new_n3355_), .B(new_n1496_), .ZN(new_n3356_));
  AOI21_X1   g2971(.A1(new_n3356_), .A2(new_n2351_), .B(new_n2352_), .ZN(new_n3357_));
  OAI21_X1   g2972(.A1(new_n3357_), .A2(new_n1516_), .B(new_n1522_), .ZN(new_n3358_));
  AOI21_X1   g2973(.A1(new_n3358_), .A2(new_n2349_), .B(new_n2350_), .ZN(new_n3359_));
  OAI21_X1   g2974(.A1(new_n3359_), .A2(new_n1542_), .B(new_n1548_), .ZN(new_n3360_));
  AOI21_X1   g2975(.A1(new_n3360_), .A2(new_n2347_), .B(new_n2348_), .ZN(new_n3361_));
  OAI21_X1   g2976(.A1(new_n3361_), .A2(new_n1569_), .B(new_n2373_), .ZN(new_n3362_));
  AOI21_X1   g2977(.A1(new_n3362_), .A2(new_n2346_), .B(new_n2746_), .ZN(new_n3363_));
  OAI21_X1   g2978(.A1(new_n3363_), .A2(new_n827_), .B(new_n840_), .ZN(new_n3364_));
  AOI21_X1   g2979(.A1(new_n3364_), .A2(new_n2289_), .B(new_n2290_), .ZN(new_n3365_));
  OAI21_X1   g2980(.A1(new_n3365_), .A2(new_n877_), .B(new_n890_), .ZN(new_n3366_));
  AOI21_X1   g2981(.A1(new_n3366_), .A2(new_n2287_), .B(new_n2288_), .ZN(new_n3367_));
  OAI21_X1   g2982(.A1(new_n3367_), .A2(new_n927_), .B(new_n940_), .ZN(new_n3368_));
  NAND2_X1   g2983(.A1(new_n961_), .A2(new_n582_), .ZN(new_n3369_));
  AOI21_X1   g2984(.A1(new_n3368_), .A2(new_n2285_), .B(new_n3369_), .ZN(\grant[66] ));
  AOI21_X1   g2985(.A1(new_n1259_), .A2(\priority[68] ), .B(\priority[69] ), .ZN(new_n3371_));
  NOR4_X1    g2986(.A1(new_n969_), .A2(new_n1663_), .A3(new_n1665_), .A4(new_n3371_), .ZN(new_n3372_));
  OAI21_X1   g2987(.A1(new_n1673_), .A2(new_n3372_), .B(new_n1679_), .ZN(new_n3373_));
  AOI21_X1   g2988(.A1(new_n3373_), .A2(new_n2382_), .B(new_n2383_), .ZN(new_n3374_));
  OAI21_X1   g2989(.A1(new_n3374_), .A2(new_n1699_), .B(new_n1705_), .ZN(new_n3375_));
  AOI21_X1   g2990(.A1(new_n3375_), .A2(new_n2380_), .B(new_n2381_), .ZN(new_n3376_));
  OAI21_X1   g2991(.A1(new_n3376_), .A2(new_n1725_), .B(new_n1731_), .ZN(new_n3377_));
  AOI21_X1   g2992(.A1(new_n3377_), .A2(new_n2378_), .B(new_n2379_), .ZN(new_n3378_));
  OAI21_X1   g2993(.A1(new_n3378_), .A2(new_n1750_), .B(new_n2404_), .ZN(new_n3379_));
  AOI21_X1   g2994(.A1(new_n3379_), .A2(new_n2377_), .B(new_n2764_), .ZN(new_n3380_));
  OAI21_X1   g2995(.A1(new_n3380_), .A2(new_n1167_), .B(new_n1176_), .ZN(new_n3381_));
  AOI21_X1   g2996(.A1(new_n3381_), .A2(new_n2326_), .B(new_n2327_), .ZN(new_n3382_));
  OAI21_X1   g2997(.A1(new_n3382_), .A2(new_n1203_), .B(new_n1212_), .ZN(new_n3383_));
  AOI21_X1   g2998(.A1(new_n3383_), .A2(new_n2324_), .B(new_n2325_), .ZN(new_n3384_));
  OAI21_X1   g2999(.A1(new_n3384_), .A2(new_n1239_), .B(new_n1248_), .ZN(new_n3385_));
  NAND2_X1   g3000(.A1(new_n1264_), .A2(new_n955_), .ZN(new_n3386_));
  AOI21_X1   g3001(.A1(new_n3385_), .A2(new_n2322_), .B(new_n3386_), .ZN(\grant[67] ));
  NOR4_X1    g3002(.A1(new_n1270_), .A2(new_n1996_), .A3(new_n1855_), .A4(new_n1852_), .ZN(new_n3388_));
  OAI21_X1   g3003(.A1(new_n1863_), .A2(new_n3388_), .B(new_n1870_), .ZN(new_n3389_));
  AOI21_X1   g3004(.A1(new_n3389_), .A2(new_n2413_), .B(new_n2414_), .ZN(new_n3390_));
  OAI21_X1   g3005(.A1(new_n3390_), .A2(new_n1891_), .B(new_n1898_), .ZN(new_n3391_));
  AOI21_X1   g3006(.A1(new_n3391_), .A2(new_n2411_), .B(new_n2412_), .ZN(new_n3392_));
  OAI21_X1   g3007(.A1(new_n3392_), .A2(new_n1919_), .B(new_n1926_), .ZN(new_n3393_));
  AOI21_X1   g3008(.A1(new_n3393_), .A2(new_n2409_), .B(new_n2410_), .ZN(new_n3394_));
  OAI21_X1   g3009(.A1(new_n3394_), .A2(new_n1945_), .B(new_n2434_), .ZN(new_n3395_));
  AOI21_X1   g3010(.A1(new_n3395_), .A2(new_n2408_), .B(new_n2782_), .ZN(new_n3396_));
  OAI21_X1   g3011(.A1(new_n3396_), .A2(new_n1412_), .B(new_n1418_), .ZN(new_n3397_));
  AOI21_X1   g3012(.A1(new_n3397_), .A2(new_n2357_), .B(new_n2358_), .ZN(new_n3398_));
  OAI21_X1   g3013(.A1(new_n3398_), .A2(new_n1438_), .B(new_n1444_), .ZN(new_n3399_));
  AOI21_X1   g3014(.A1(new_n3399_), .A2(new_n2355_), .B(new_n2356_), .ZN(new_n3400_));
  OAI21_X1   g3015(.A1(new_n3400_), .A2(new_n1464_), .B(new_n1470_), .ZN(new_n3401_));
  NAND2_X1   g3016(.A1(new_n1479_), .A2(new_n1259_), .ZN(new_n3402_));
  AOI21_X1   g3017(.A1(new_n3401_), .A2(new_n2353_), .B(new_n3402_), .ZN(\grant[68] ));
  NOR4_X1    g3018(.A1(new_n1487_), .A2(new_n604_), .A3(new_n1998_), .A4(new_n2092_), .ZN(new_n3404_));
  OAI21_X1   g3019(.A1(new_n2003_), .A2(new_n3404_), .B(new_n2006_), .ZN(new_n3405_));
  AOI21_X1   g3020(.A1(new_n3405_), .A2(new_n2443_), .B(new_n2444_), .ZN(new_n3406_));
  OAI21_X1   g3021(.A1(new_n3406_), .A2(new_n2017_), .B(new_n2020_), .ZN(new_n3407_));
  AOI21_X1   g3022(.A1(new_n3407_), .A2(new_n2441_), .B(new_n2442_), .ZN(new_n3408_));
  OAI21_X1   g3023(.A1(new_n3408_), .A2(new_n2031_), .B(new_n2034_), .ZN(new_n3409_));
  AOI21_X1   g3024(.A1(new_n3409_), .A2(new_n2439_), .B(new_n2440_), .ZN(new_n3410_));
  OAI21_X1   g3025(.A1(new_n3410_), .A2(new_n2048_), .B(new_n2464_), .ZN(new_n3411_));
  AOI21_X1   g3026(.A1(new_n3411_), .A2(new_n2438_), .B(new_n2799_), .ZN(new_n3412_));
  OAI21_X1   g3027(.A1(new_n3412_), .A2(new_n1595_), .B(new_n1601_), .ZN(new_n3413_));
  AOI21_X1   g3028(.A1(new_n3413_), .A2(new_n2388_), .B(new_n2389_), .ZN(new_n3414_));
  OAI21_X1   g3029(.A1(new_n3414_), .A2(new_n1621_), .B(new_n1627_), .ZN(new_n3415_));
  AOI21_X1   g3030(.A1(new_n3415_), .A2(new_n2386_), .B(new_n2387_), .ZN(new_n3416_));
  OAI21_X1   g3031(.A1(new_n3416_), .A2(new_n1647_), .B(new_n1653_), .ZN(new_n3417_));
  NAND2_X1   g3032(.A1(new_n1662_), .A2(new_n596_), .ZN(new_n3418_));
  AOI21_X1   g3033(.A1(new_n3417_), .A2(new_n2384_), .B(new_n3418_), .ZN(\grant[69] ));
  NOR4_X1    g3034(.A1(new_n1670_), .A2(new_n975_), .A3(new_n2094_), .A4(new_n2190_), .ZN(new_n3420_));
  OAI21_X1   g3035(.A1(new_n2098_), .A2(new_n3420_), .B(new_n2101_), .ZN(new_n3421_));
  AOI21_X1   g3036(.A1(new_n3421_), .A2(new_n2473_), .B(new_n2474_), .ZN(new_n3422_));
  OAI21_X1   g3037(.A1(new_n3422_), .A2(new_n2110_), .B(new_n2113_), .ZN(new_n3423_));
  AOI21_X1   g3038(.A1(new_n3423_), .A2(new_n2471_), .B(new_n2472_), .ZN(new_n3424_));
  OAI21_X1   g3039(.A1(new_n3424_), .A2(new_n2122_), .B(new_n2125_), .ZN(new_n3425_));
  AOI21_X1   g3040(.A1(new_n3425_), .A2(new_n2469_), .B(new_n2470_), .ZN(new_n3426_));
  OAI21_X1   g3041(.A1(new_n3426_), .A2(new_n2139_), .B(new_n2494_), .ZN(new_n3427_));
  AOI21_X1   g3042(.A1(new_n3427_), .A2(new_n2468_), .B(new_n2816_), .ZN(new_n3428_));
  OAI21_X1   g3043(.A1(new_n3428_), .A2(new_n1779_), .B(new_n1786_), .ZN(new_n3429_));
  AOI21_X1   g3044(.A1(new_n3429_), .A2(new_n2419_), .B(new_n2420_), .ZN(new_n3430_));
  OAI21_X1   g3045(.A1(new_n3430_), .A2(new_n1807_), .B(new_n1814_), .ZN(new_n3431_));
  AOI21_X1   g3046(.A1(new_n3431_), .A2(new_n2417_), .B(new_n2418_), .ZN(new_n3432_));
  OAI21_X1   g3047(.A1(new_n3432_), .A2(new_n1835_), .B(new_n1842_), .ZN(new_n3433_));
  NAND2_X1   g3048(.A1(new_n1851_), .A2(new_n967_), .ZN(new_n3434_));
  AOI21_X1   g3049(.A1(new_n3433_), .A2(new_n2415_), .B(new_n3434_), .ZN(\grant[70] ));
  OAI21_X1   g3050(.A1(new_n600_), .A2(\priority[73] ), .B(new_n1854_), .ZN(new_n3436_));
  NOR3_X1    g3051(.A1(new_n3436_), .A2(new_n1860_), .A3(new_n2193_), .ZN(new_n3437_));
  OAI21_X1   g3052(.A1(new_n2197_), .A2(new_n3437_), .B(new_n2201_), .ZN(new_n3438_));
  AOI21_X1   g3053(.A1(new_n3438_), .A2(new_n2503_), .B(new_n2504_), .ZN(new_n3439_));
  OAI21_X1   g3054(.A1(new_n3439_), .A2(new_n2211_), .B(new_n2215_), .ZN(new_n3440_));
  AOI21_X1   g3055(.A1(new_n3440_), .A2(new_n2501_), .B(new_n2502_), .ZN(new_n3441_));
  OAI21_X1   g3056(.A1(new_n3441_), .A2(new_n2225_), .B(new_n2229_), .ZN(new_n3442_));
  AOI21_X1   g3057(.A1(new_n3442_), .A2(new_n2499_), .B(new_n2500_), .ZN(new_n3443_));
  OAI21_X1   g3058(.A1(new_n3443_), .A2(new_n2239_), .B(new_n2525_), .ZN(new_n3444_));
  AOI21_X1   g3059(.A1(new_n3444_), .A2(new_n2498_), .B(new_n2833_), .ZN(new_n3445_));
  OAI21_X1   g3060(.A1(new_n3445_), .A2(new_n1961_), .B(new_n1964_), .ZN(new_n3446_));
  AOI21_X1   g3061(.A1(new_n3446_), .A2(new_n2449_), .B(new_n2450_), .ZN(new_n3447_));
  OAI21_X1   g3062(.A1(new_n3447_), .A2(new_n1975_), .B(new_n1978_), .ZN(new_n3448_));
  AOI21_X1   g3063(.A1(new_n3448_), .A2(new_n2447_), .B(new_n2448_), .ZN(new_n3449_));
  OAI21_X1   g3064(.A1(new_n3449_), .A2(new_n1989_), .B(new_n1992_), .ZN(new_n3450_));
  NAND2_X1   g3065(.A1(new_n602_), .A2(new_n1268_), .ZN(new_n3451_));
  AOI21_X1   g3066(.A1(new_n3450_), .A2(new_n2445_), .B(new_n3451_), .ZN(\grant[71] ));
  AOI21_X1   g3067(.A1(new_n1668_), .A2(\priority[73] ), .B(\priority[74] ), .ZN(new_n3453_));
  NOR4_X1    g3068(.A1(new_n612_), .A2(new_n614_), .A3(new_n618_), .A4(new_n3453_), .ZN(new_n3454_));
  OAI21_X1   g3069(.A1(new_n635_), .A2(new_n3454_), .B(new_n648_), .ZN(new_n3455_));
  AOI21_X1   g3070(.A1(new_n3455_), .A2(new_n663_), .B(new_n677_), .ZN(new_n3456_));
  OAI21_X1   g3071(.A1(new_n3456_), .A2(new_n691_), .B(new_n704_), .ZN(new_n3457_));
  AOI21_X1   g3072(.A1(new_n3457_), .A2(new_n719_), .B(new_n733_), .ZN(new_n3458_));
  OAI21_X1   g3073(.A1(new_n3458_), .A2(new_n747_), .B(new_n760_), .ZN(new_n3459_));
  AOI21_X1   g3074(.A1(new_n3459_), .A2(new_n775_), .B(new_n2530_), .ZN(new_n3460_));
  OAI21_X1   g3075(.A1(new_n3460_), .A2(new_n2275_), .B(new_n2545_), .ZN(new_n3461_));
  AOI21_X1   g3076(.A1(new_n3461_), .A2(new_n2529_), .B(new_n2851_), .ZN(new_n3462_));
  OAI21_X1   g3077(.A1(new_n3462_), .A2(new_n2062_), .B(new_n2065_), .ZN(new_n3463_));
  AOI21_X1   g3078(.A1(new_n3463_), .A2(new_n2479_), .B(new_n2480_), .ZN(new_n3464_));
  OAI21_X1   g3079(.A1(new_n3464_), .A2(new_n2074_), .B(new_n2077_), .ZN(new_n3465_));
  AOI21_X1   g3080(.A1(new_n3465_), .A2(new_n2477_), .B(new_n2478_), .ZN(new_n3466_));
  OAI21_X1   g3081(.A1(new_n3466_), .A2(new_n2086_), .B(new_n2089_), .ZN(new_n3467_));
  NAND2_X1   g3082(.A1(new_n973_), .A2(new_n1485_), .ZN(new_n3468_));
  AOI21_X1   g3083(.A1(new_n3467_), .A2(new_n2475_), .B(new_n3468_), .ZN(\grant[72] ));
  AOI21_X1   g3084(.A1(new_n1858_), .A2(\priority[74] ), .B(\priority[75] ), .ZN(new_n3470_));
  NOR4_X1    g3085(.A1(new_n982_), .A2(new_n984_), .A3(new_n988_), .A4(new_n3470_), .ZN(new_n3471_));
  OAI21_X1   g3086(.A1(new_n1003_), .A2(new_n3471_), .B(new_n1015_), .ZN(new_n3472_));
  AOI21_X1   g3087(.A1(new_n3472_), .A2(new_n1028_), .B(new_n1041_), .ZN(new_n3473_));
  OAI21_X1   g3088(.A1(new_n3473_), .A2(new_n1053_), .B(new_n1065_), .ZN(new_n3474_));
  AOI21_X1   g3089(.A1(new_n3474_), .A2(new_n1078_), .B(new_n1091_), .ZN(new_n3475_));
  OAI21_X1   g3090(.A1(new_n3475_), .A2(new_n1103_), .B(new_n1115_), .ZN(new_n3476_));
  AOI21_X1   g3091(.A1(new_n3476_), .A2(new_n1128_), .B(new_n2550_), .ZN(new_n3477_));
  OAI21_X1   g3092(.A1(new_n3477_), .A2(new_n2311_), .B(new_n2565_), .ZN(new_n3478_));
  AOI21_X1   g3093(.A1(new_n3478_), .A2(new_n2549_), .B(new_n2869_), .ZN(new_n3479_));
  OAI21_X1   g3094(.A1(new_n3479_), .A2(new_n2155_), .B(new_n2159_), .ZN(new_n3480_));
  AOI21_X1   g3095(.A1(new_n3480_), .A2(new_n2509_), .B(new_n2510_), .ZN(new_n3481_));
  OAI21_X1   g3096(.A1(new_n3481_), .A2(new_n2169_), .B(new_n2173_), .ZN(new_n3482_));
  AOI21_X1   g3097(.A1(new_n3482_), .A2(new_n2507_), .B(new_n2508_), .ZN(new_n3483_));
  OAI21_X1   g3098(.A1(new_n3483_), .A2(new_n2183_), .B(new_n2187_), .ZN(new_n3484_));
  NAND2_X1   g3099(.A1(new_n1273_), .A2(new_n1668_), .ZN(new_n3485_));
  AOI21_X1   g3100(.A1(new_n3484_), .A2(new_n2505_), .B(new_n3485_), .ZN(\grant[73] ));
  OAI21_X1   g3101(.A1(new_n1488_), .A2(\priority[76] ), .B(new_n2192_), .ZN(new_n3487_));
  NOR3_X1    g3102(.A1(new_n3487_), .A2(new_n1279_), .A3(new_n1281_), .ZN(new_n3488_));
  OAI21_X1   g3103(.A1(new_n1294_), .A2(new_n3488_), .B(new_n1302_), .ZN(new_n3489_));
  AOI21_X1   g3104(.A1(new_n3489_), .A2(new_n1312_), .B(new_n1321_), .ZN(new_n3490_));
  OAI21_X1   g3105(.A1(new_n3490_), .A2(new_n1330_), .B(new_n1338_), .ZN(new_n3491_));
  AOI21_X1   g3106(.A1(new_n3491_), .A2(new_n1348_), .B(new_n1357_), .ZN(new_n3492_));
  OAI21_X1   g3107(.A1(new_n3492_), .A2(new_n1366_), .B(new_n1374_), .ZN(new_n3493_));
  AOI21_X1   g3108(.A1(new_n3493_), .A2(new_n1386_), .B(new_n2569_), .ZN(new_n3494_));
  OAI21_X1   g3109(.A1(new_n3494_), .A2(new_n411_), .B(new_n424_), .ZN(new_n3495_));
  AOI21_X1   g3110(.A1(new_n3495_), .A2(new_n439_), .B(new_n453_), .ZN(new_n3496_));
  OAI21_X1   g3111(.A1(new_n3496_), .A2(new_n467_), .B(new_n480_), .ZN(new_n3497_));
  AOI21_X1   g3112(.A1(new_n3497_), .A2(new_n495_), .B(new_n509_), .ZN(new_n3498_));
  OAI21_X1   g3113(.A1(new_n3498_), .A2(new_n523_), .B(new_n536_), .ZN(new_n3499_));
  AOI21_X1   g3114(.A1(new_n3499_), .A2(new_n551_), .B(new_n565_), .ZN(new_n3500_));
  OAI21_X1   g3115(.A1(new_n3500_), .A2(new_n579_), .B(new_n592_), .ZN(new_n3501_));
  NAND2_X1   g3116(.A1(new_n616_), .A2(new_n1858_), .ZN(new_n3502_));
  AOI21_X1   g3117(.A1(new_n3501_), .A2(new_n607_), .B(new_n3502_), .ZN(\grant[74] ));
  AOI21_X1   g3118(.A1(new_n980_), .A2(\priority[76] ), .B(\priority[77] ), .ZN(new_n3504_));
  NOR4_X1    g3119(.A1(new_n627_), .A2(new_n1493_), .A3(new_n1495_), .A4(new_n3504_), .ZN(new_n3505_));
  OAI21_X1   g3120(.A1(new_n1504_), .A2(new_n3505_), .B(new_n1509_), .ZN(new_n3506_));
  AOI21_X1   g3121(.A1(new_n3506_), .A2(new_n1517_), .B(new_n1523_), .ZN(new_n3507_));
  OAI21_X1   g3122(.A1(new_n3507_), .A2(new_n1530_), .B(new_n1535_), .ZN(new_n3508_));
  AOI21_X1   g3123(.A1(new_n3508_), .A2(new_n1543_), .B(new_n1549_), .ZN(new_n3509_));
  OAI21_X1   g3124(.A1(new_n3509_), .A2(new_n1556_), .B(new_n1561_), .ZN(new_n3510_));
  AOI21_X1   g3125(.A1(new_n3510_), .A2(new_n1570_), .B(new_n2587_), .ZN(new_n3511_));
  OAI21_X1   g3126(.A1(new_n3511_), .A2(new_n803_), .B(new_n815_), .ZN(new_n3512_));
  AOI21_X1   g3127(.A1(new_n3512_), .A2(new_n828_), .B(new_n841_), .ZN(new_n3513_));
  OAI21_X1   g3128(.A1(new_n3513_), .A2(new_n853_), .B(new_n865_), .ZN(new_n3514_));
  AOI21_X1   g3129(.A1(new_n3514_), .A2(new_n878_), .B(new_n891_), .ZN(new_n3515_));
  OAI21_X1   g3130(.A1(new_n3515_), .A2(new_n903_), .B(new_n915_), .ZN(new_n3516_));
  AOI21_X1   g3131(.A1(new_n3516_), .A2(new_n928_), .B(new_n941_), .ZN(new_n3517_));
  OAI21_X1   g3132(.A1(new_n3517_), .A2(new_n953_), .B(new_n965_), .ZN(new_n3518_));
  NAND2_X1   g3133(.A1(new_n986_), .A2(new_n610_), .ZN(new_n3519_));
  AOI21_X1   g3134(.A1(new_n3518_), .A2(new_n978_), .B(new_n3519_), .ZN(\grant[75] ));
  AOI21_X1   g3135(.A1(new_n1277_), .A2(\priority[77] ), .B(\priority[78] ), .ZN(new_n3521_));
  NOR4_X1    g3136(.A1(new_n995_), .A2(new_n1676_), .A3(new_n1678_), .A4(new_n3521_), .ZN(new_n3522_));
  OAI21_X1   g3137(.A1(new_n1687_), .A2(new_n3522_), .B(new_n1692_), .ZN(new_n3523_));
  AOI21_X1   g3138(.A1(new_n3523_), .A2(new_n1700_), .B(new_n1706_), .ZN(new_n3524_));
  OAI21_X1   g3139(.A1(new_n3524_), .A2(new_n1713_), .B(new_n1718_), .ZN(new_n3525_));
  AOI21_X1   g3140(.A1(new_n3525_), .A2(new_n1726_), .B(new_n1732_), .ZN(new_n3526_));
  OAI21_X1   g3141(.A1(new_n3526_), .A2(new_n1739_), .B(new_n1744_), .ZN(new_n3527_));
  AOI21_X1   g3142(.A1(new_n3527_), .A2(new_n1751_), .B(new_n2605_), .ZN(new_n3528_));
  OAI21_X1   g3143(.A1(new_n3528_), .A2(new_n1150_), .B(new_n1158_), .ZN(new_n3529_));
  AOI21_X1   g3144(.A1(new_n3529_), .A2(new_n1168_), .B(new_n1177_), .ZN(new_n3530_));
  OAI21_X1   g3145(.A1(new_n3530_), .A2(new_n1186_), .B(new_n1194_), .ZN(new_n3531_));
  AOI21_X1   g3146(.A1(new_n3531_), .A2(new_n1204_), .B(new_n1213_), .ZN(new_n3532_));
  OAI21_X1   g3147(.A1(new_n3532_), .A2(new_n1222_), .B(new_n1230_), .ZN(new_n3533_));
  AOI21_X1   g3148(.A1(new_n3533_), .A2(new_n1240_), .B(new_n1249_), .ZN(new_n3534_));
  OAI21_X1   g3149(.A1(new_n3534_), .A2(new_n1258_), .B(new_n1266_), .ZN(new_n3535_));
  NAND2_X1   g3150(.A1(new_n1282_), .A2(new_n980_), .ZN(new_n3536_));
  AOI21_X1   g3151(.A1(new_n3535_), .A2(new_n1276_), .B(new_n3536_), .ZN(\grant[76] ));
  NOR4_X1    g3152(.A1(new_n1289_), .A2(new_n2002_), .A3(new_n1869_), .A4(new_n1866_), .ZN(new_n3538_));
  OAI21_X1   g3153(.A1(new_n1878_), .A2(new_n3538_), .B(new_n1884_), .ZN(new_n3539_));
  AOI21_X1   g3154(.A1(new_n3539_), .A2(new_n1892_), .B(new_n1899_), .ZN(new_n3540_));
  OAI21_X1   g3155(.A1(new_n3540_), .A2(new_n1906_), .B(new_n1912_), .ZN(new_n3541_));
  AOI21_X1   g3156(.A1(new_n3541_), .A2(new_n1920_), .B(new_n1927_), .ZN(new_n3542_));
  OAI21_X1   g3157(.A1(new_n3542_), .A2(new_n1934_), .B(new_n1939_), .ZN(new_n3543_));
  AOI21_X1   g3158(.A1(new_n3543_), .A2(new_n1946_), .B(new_n2623_), .ZN(new_n3544_));
  OAI21_X1   g3159(.A1(new_n3544_), .A2(new_n1400_), .B(new_n1405_), .ZN(new_n3545_));
  AOI21_X1   g3160(.A1(new_n3545_), .A2(new_n1413_), .B(new_n1419_), .ZN(new_n3546_));
  OAI21_X1   g3161(.A1(new_n3546_), .A2(new_n1426_), .B(new_n1431_), .ZN(new_n3547_));
  AOI21_X1   g3162(.A1(new_n3547_), .A2(new_n1439_), .B(new_n1445_), .ZN(new_n3548_));
  OAI21_X1   g3163(.A1(new_n3548_), .A2(new_n1452_), .B(new_n1457_), .ZN(new_n3549_));
  AOI21_X1   g3164(.A1(new_n3549_), .A2(new_n1465_), .B(new_n1471_), .ZN(new_n3550_));
  OAI21_X1   g3165(.A1(new_n3550_), .A2(new_n1478_), .B(new_n1483_), .ZN(new_n3551_));
  NAND2_X1   g3166(.A1(new_n1492_), .A2(new_n1277_), .ZN(new_n3552_));
  AOI21_X1   g3167(.A1(new_n3551_), .A2(new_n1491_), .B(new_n3552_), .ZN(\grant[77] ));
  NOR4_X1    g3168(.A1(new_n1501_), .A2(new_n633_), .A3(new_n2005_), .A4(new_n2097_), .ZN(new_n3554_));
  OAI21_X1   g3169(.A1(new_n2011_), .A2(new_n3554_), .B(new_n2013_), .ZN(new_n3555_));
  AOI21_X1   g3170(.A1(new_n3555_), .A2(new_n2018_), .B(new_n2021_), .ZN(new_n3556_));
  OAI21_X1   g3171(.A1(new_n3556_), .A2(new_n2025_), .B(new_n2027_), .ZN(new_n3557_));
  AOI21_X1   g3172(.A1(new_n3557_), .A2(new_n2032_), .B(new_n2035_), .ZN(new_n3558_));
  OAI21_X1   g3173(.A1(new_n3558_), .A2(new_n2039_), .B(new_n2041_), .ZN(new_n3559_));
  AOI21_X1   g3174(.A1(new_n3559_), .A2(new_n2049_), .B(new_n2640_), .ZN(new_n3560_));
  OAI21_X1   g3175(.A1(new_n3560_), .A2(new_n1583_), .B(new_n1588_), .ZN(new_n3561_));
  AOI21_X1   g3176(.A1(new_n3561_), .A2(new_n1596_), .B(new_n1602_), .ZN(new_n3562_));
  OAI21_X1   g3177(.A1(new_n3562_), .A2(new_n1609_), .B(new_n1614_), .ZN(new_n3563_));
  AOI21_X1   g3178(.A1(new_n3563_), .A2(new_n1622_), .B(new_n1628_), .ZN(new_n3564_));
  OAI21_X1   g3179(.A1(new_n3564_), .A2(new_n1635_), .B(new_n1640_), .ZN(new_n3565_));
  AOI21_X1   g3180(.A1(new_n3565_), .A2(new_n1648_), .B(new_n1654_), .ZN(new_n3566_));
  OAI21_X1   g3181(.A1(new_n3566_), .A2(new_n1661_), .B(new_n1666_), .ZN(new_n3567_));
  NAND2_X1   g3182(.A1(new_n1675_), .A2(new_n625_), .ZN(new_n3568_));
  AOI21_X1   g3183(.A1(new_n3567_), .A2(new_n1674_), .B(new_n3568_), .ZN(\grant[78] ));
  NOR4_X1    g3184(.A1(new_n1684_), .A2(new_n1001_), .A3(new_n2100_), .A4(new_n2196_), .ZN(new_n3570_));
  OAI21_X1   g3185(.A1(new_n2105_), .A2(new_n3570_), .B(new_n2107_), .ZN(new_n3571_));
  AOI21_X1   g3186(.A1(new_n3571_), .A2(new_n2111_), .B(new_n2114_), .ZN(new_n3572_));
  OAI21_X1   g3187(.A1(new_n3572_), .A2(new_n2117_), .B(new_n2119_), .ZN(new_n3573_));
  AOI21_X1   g3188(.A1(new_n3573_), .A2(new_n2123_), .B(new_n2126_), .ZN(new_n3574_));
  OAI21_X1   g3189(.A1(new_n3574_), .A2(new_n2129_), .B(new_n2132_), .ZN(new_n3575_));
  AOI21_X1   g3190(.A1(new_n3575_), .A2(new_n2140_), .B(new_n2657_), .ZN(new_n3576_));
  OAI21_X1   g3191(.A1(new_n3576_), .A2(new_n1766_), .B(new_n1772_), .ZN(new_n3577_));
  AOI21_X1   g3192(.A1(new_n3577_), .A2(new_n1780_), .B(new_n1787_), .ZN(new_n3578_));
  OAI21_X1   g3193(.A1(new_n3578_), .A2(new_n1794_), .B(new_n1800_), .ZN(new_n3579_));
  AOI21_X1   g3194(.A1(new_n3579_), .A2(new_n1808_), .B(new_n1815_), .ZN(new_n3580_));
  OAI21_X1   g3195(.A1(new_n3580_), .A2(new_n1822_), .B(new_n1828_), .ZN(new_n3581_));
  AOI21_X1   g3196(.A1(new_n3581_), .A2(new_n1836_), .B(new_n1843_), .ZN(new_n3582_));
  OAI21_X1   g3197(.A1(new_n3582_), .A2(new_n1850_), .B(new_n1856_), .ZN(new_n3583_));
  NAND2_X1   g3198(.A1(new_n1865_), .A2(new_n993_), .ZN(new_n3584_));
  AOI21_X1   g3199(.A1(new_n3583_), .A2(new_n1864_), .B(new_n3584_), .ZN(\grant[79] ));
  OAI21_X1   g3200(.A1(new_n629_), .A2(\priority[82] ), .B(new_n1868_), .ZN(new_n3586_));
  NOR3_X1    g3201(.A1(new_n3586_), .A2(new_n1875_), .A3(new_n2200_), .ZN(new_n3587_));
  OAI21_X1   g3202(.A1(new_n2205_), .A2(new_n3587_), .B(new_n2208_), .ZN(new_n3588_));
  AOI21_X1   g3203(.A1(new_n3588_), .A2(new_n2212_), .B(new_n2216_), .ZN(new_n3589_));
  OAI21_X1   g3204(.A1(new_n3589_), .A2(new_n2219_), .B(new_n2222_), .ZN(new_n3590_));
  AOI21_X1   g3205(.A1(new_n3590_), .A2(new_n2226_), .B(new_n2230_), .ZN(new_n3591_));
  OAI21_X1   g3206(.A1(new_n3591_), .A2(new_n2233_), .B(new_n2235_), .ZN(new_n3592_));
  AOI21_X1   g3207(.A1(new_n3592_), .A2(new_n2240_), .B(new_n2674_), .ZN(new_n3593_));
  OAI21_X1   g3208(.A1(new_n3593_), .A2(new_n1955_), .B(new_n1957_), .ZN(new_n3594_));
  AOI21_X1   g3209(.A1(new_n3594_), .A2(new_n1962_), .B(new_n1965_), .ZN(new_n3595_));
  OAI21_X1   g3210(.A1(new_n3595_), .A2(new_n1969_), .B(new_n1971_), .ZN(new_n3596_));
  AOI21_X1   g3211(.A1(new_n3596_), .A2(new_n1976_), .B(new_n1979_), .ZN(new_n3597_));
  OAI21_X1   g3212(.A1(new_n3597_), .A2(new_n1983_), .B(new_n1985_), .ZN(new_n3598_));
  AOI21_X1   g3213(.A1(new_n3598_), .A2(new_n1990_), .B(new_n1993_), .ZN(new_n3599_));
  OAI21_X1   g3214(.A1(new_n3599_), .A2(new_n1997_), .B(new_n1999_), .ZN(new_n3600_));
  NAND2_X1   g3215(.A1(new_n631_), .A2(new_n1287_), .ZN(new_n3601_));
  AOI21_X1   g3216(.A1(new_n3600_), .A2(new_n2004_), .B(new_n3601_), .ZN(\grant[80] ));
  AOI21_X1   g3217(.A1(new_n1682_), .A2(\priority[82] ), .B(\priority[83] ), .ZN(new_n3603_));
  NOR4_X1    g3218(.A1(new_n640_), .A2(new_n642_), .A3(new_n646_), .A4(new_n3603_), .ZN(new_n3604_));
  OAI21_X1   g3219(.A1(new_n662_), .A2(new_n3604_), .B(new_n676_), .ZN(new_n3605_));
  AOI21_X1   g3220(.A1(new_n3605_), .A2(new_n2245_), .B(new_n2246_), .ZN(new_n3606_));
  OAI21_X1   g3221(.A1(new_n3606_), .A2(new_n718_), .B(new_n732_), .ZN(new_n3607_));
  AOI21_X1   g3222(.A1(new_n3607_), .A2(new_n2243_), .B(new_n2244_), .ZN(new_n3608_));
  OAI21_X1   g3223(.A1(new_n3608_), .A2(new_n774_), .B(new_n2270_), .ZN(new_n3609_));
  AOI21_X1   g3224(.A1(new_n3609_), .A2(new_n2276_), .B(new_n2692_), .ZN(new_n3610_));
  OAI21_X1   g3225(.A1(new_n3610_), .A2(new_n2057_), .B(new_n2059_), .ZN(new_n3611_));
  AOI21_X1   g3226(.A1(new_n3611_), .A2(new_n2063_), .B(new_n2066_), .ZN(new_n3612_));
  OAI21_X1   g3227(.A1(new_n3612_), .A2(new_n2069_), .B(new_n2071_), .ZN(new_n3613_));
  AOI21_X1   g3228(.A1(new_n3613_), .A2(new_n2075_), .B(new_n2078_), .ZN(new_n3614_));
  OAI21_X1   g3229(.A1(new_n3614_), .A2(new_n2081_), .B(new_n2083_), .ZN(new_n3615_));
  AOI21_X1   g3230(.A1(new_n3615_), .A2(new_n2087_), .B(new_n2090_), .ZN(new_n3616_));
  OAI21_X1   g3231(.A1(new_n3616_), .A2(new_n2093_), .B(new_n2095_), .ZN(new_n3617_));
  NAND2_X1   g3232(.A1(new_n999_), .A2(new_n1499_), .ZN(new_n3618_));
  AOI21_X1   g3233(.A1(new_n3617_), .A2(new_n2099_), .B(new_n3618_), .ZN(\grant[81] ));
  AOI21_X1   g3234(.A1(new_n1873_), .A2(\priority[83] ), .B(\priority[84] ), .ZN(new_n3620_));
  NOR4_X1    g3235(.A1(new_n1007_), .A2(new_n1009_), .A3(new_n1013_), .A4(new_n3620_), .ZN(new_n3621_));
  OAI21_X1   g3236(.A1(new_n1027_), .A2(new_n3621_), .B(new_n1040_), .ZN(new_n3622_));
  AOI21_X1   g3237(.A1(new_n3622_), .A2(new_n2281_), .B(new_n2282_), .ZN(new_n3623_));
  OAI21_X1   g3238(.A1(new_n3623_), .A2(new_n1077_), .B(new_n1090_), .ZN(new_n3624_));
  AOI21_X1   g3239(.A1(new_n3624_), .A2(new_n2279_), .B(new_n2280_), .ZN(new_n3625_));
  OAI21_X1   g3240(.A1(new_n3625_), .A2(new_n1127_), .B(new_n2306_), .ZN(new_n3626_));
  AOI21_X1   g3241(.A1(new_n3626_), .A2(new_n2312_), .B(new_n2710_), .ZN(new_n3627_));
  OAI21_X1   g3242(.A1(new_n3627_), .A2(new_n2149_), .B(new_n2152_), .ZN(new_n3628_));
  AOI21_X1   g3243(.A1(new_n3628_), .A2(new_n2156_), .B(new_n2160_), .ZN(new_n3629_));
  OAI21_X1   g3244(.A1(new_n3629_), .A2(new_n2163_), .B(new_n2166_), .ZN(new_n3630_));
  AOI21_X1   g3245(.A1(new_n3630_), .A2(new_n2170_), .B(new_n2174_), .ZN(new_n3631_));
  OAI21_X1   g3246(.A1(new_n3631_), .A2(new_n2177_), .B(new_n2180_), .ZN(new_n3632_));
  AOI21_X1   g3247(.A1(new_n3632_), .A2(new_n2184_), .B(new_n2188_), .ZN(new_n3633_));
  OAI21_X1   g3248(.A1(new_n3633_), .A2(new_n2191_), .B(new_n2194_), .ZN(new_n3634_));
  NAND2_X1   g3249(.A1(new_n1292_), .A2(new_n1682_), .ZN(new_n3635_));
  AOI21_X1   g3250(.A1(new_n3634_), .A2(new_n2198_), .B(new_n3635_), .ZN(\grant[82] ));
  OAI21_X1   g3251(.A1(new_n1502_), .A2(\priority[85] ), .B(new_n2199_), .ZN(new_n3637_));
  NOR3_X1    g3252(.A1(new_n3637_), .A2(new_n1297_), .A3(new_n1299_), .ZN(new_n3638_));
  OAI21_X1   g3253(.A1(new_n1311_), .A2(new_n3638_), .B(new_n1320_), .ZN(new_n3639_));
  AOI21_X1   g3254(.A1(new_n3639_), .A2(new_n2318_), .B(new_n2319_), .ZN(new_n3640_));
  OAI21_X1   g3255(.A1(new_n3640_), .A2(new_n1347_), .B(new_n1356_), .ZN(new_n3641_));
  AOI21_X1   g3256(.A1(new_n3641_), .A2(new_n2316_), .B(new_n2317_), .ZN(new_n3642_));
  OAI21_X1   g3257(.A1(new_n3642_), .A2(new_n1385_), .B(new_n2342_), .ZN(new_n3643_));
  AOI21_X1   g3258(.A1(new_n3643_), .A2(new_n2315_), .B(new_n2728_), .ZN(new_n3644_));
  OAI21_X1   g3259(.A1(new_n3644_), .A2(new_n438_), .B(new_n452_), .ZN(new_n3645_));
  AOI21_X1   g3260(.A1(new_n3645_), .A2(new_n2253_), .B(new_n2254_), .ZN(new_n3646_));
  OAI21_X1   g3261(.A1(new_n3646_), .A2(new_n494_), .B(new_n508_), .ZN(new_n3647_));
  AOI21_X1   g3262(.A1(new_n3647_), .A2(new_n2251_), .B(new_n2252_), .ZN(new_n3648_));
  OAI21_X1   g3263(.A1(new_n3648_), .A2(new_n550_), .B(new_n564_), .ZN(new_n3649_));
  AOI21_X1   g3264(.A1(new_n3649_), .A2(new_n2249_), .B(new_n2250_), .ZN(new_n3650_));
  OAI21_X1   g3265(.A1(new_n3650_), .A2(new_n606_), .B(new_n620_), .ZN(new_n3651_));
  NAND2_X1   g3266(.A1(new_n644_), .A2(new_n1873_), .ZN(new_n3652_));
  AOI21_X1   g3267(.A1(new_n3651_), .A2(new_n2247_), .B(new_n3652_), .ZN(\grant[83] ));
  AOI21_X1   g3268(.A1(new_n1005_), .A2(\priority[85] ), .B(\priority[86] ), .ZN(new_n3654_));
  NOR4_X1    g3269(.A1(new_n654_), .A2(new_n1506_), .A3(new_n1508_), .A4(new_n3654_), .ZN(new_n3655_));
  OAI21_X1   g3270(.A1(new_n1516_), .A2(new_n3655_), .B(new_n1522_), .ZN(new_n3656_));
  AOI21_X1   g3271(.A1(new_n3656_), .A2(new_n2349_), .B(new_n2350_), .ZN(new_n3657_));
  OAI21_X1   g3272(.A1(new_n3657_), .A2(new_n1542_), .B(new_n1548_), .ZN(new_n3658_));
  AOI21_X1   g3273(.A1(new_n3658_), .A2(new_n2347_), .B(new_n2348_), .ZN(new_n3659_));
  OAI21_X1   g3274(.A1(new_n3659_), .A2(new_n1569_), .B(new_n2373_), .ZN(new_n3660_));
  AOI21_X1   g3275(.A1(new_n3660_), .A2(new_n2346_), .B(new_n2746_), .ZN(new_n3661_));
  OAI21_X1   g3276(.A1(new_n3661_), .A2(new_n827_), .B(new_n840_), .ZN(new_n3662_));
  AOI21_X1   g3277(.A1(new_n3662_), .A2(new_n2289_), .B(new_n2290_), .ZN(new_n3663_));
  OAI21_X1   g3278(.A1(new_n3663_), .A2(new_n877_), .B(new_n890_), .ZN(new_n3664_));
  AOI21_X1   g3279(.A1(new_n3664_), .A2(new_n2287_), .B(new_n2288_), .ZN(new_n3665_));
  OAI21_X1   g3280(.A1(new_n3665_), .A2(new_n927_), .B(new_n940_), .ZN(new_n3666_));
  AOI21_X1   g3281(.A1(new_n3666_), .A2(new_n2285_), .B(new_n2286_), .ZN(new_n3667_));
  OAI21_X1   g3282(.A1(new_n3667_), .A2(new_n977_), .B(new_n990_), .ZN(new_n3668_));
  NAND2_X1   g3283(.A1(new_n1011_), .A2(new_n638_), .ZN(new_n3669_));
  AOI21_X1   g3284(.A1(new_n3668_), .A2(new_n2283_), .B(new_n3669_), .ZN(\grant[84] ));
  AOI21_X1   g3285(.A1(new_n1295_), .A2(\priority[86] ), .B(\priority[87] ), .ZN(new_n3671_));
  NOR4_X1    g3286(.A1(new_n1019_), .A2(new_n1689_), .A3(new_n1691_), .A4(new_n3671_), .ZN(new_n3672_));
  OAI21_X1   g3287(.A1(new_n1699_), .A2(new_n3672_), .B(new_n1705_), .ZN(new_n3673_));
  AOI21_X1   g3288(.A1(new_n3673_), .A2(new_n2380_), .B(new_n2381_), .ZN(new_n3674_));
  OAI21_X1   g3289(.A1(new_n3674_), .A2(new_n1725_), .B(new_n1731_), .ZN(new_n3675_));
  AOI21_X1   g3290(.A1(new_n3675_), .A2(new_n2378_), .B(new_n2379_), .ZN(new_n3676_));
  OAI21_X1   g3291(.A1(new_n3676_), .A2(new_n1750_), .B(new_n2404_), .ZN(new_n3677_));
  AOI21_X1   g3292(.A1(new_n3677_), .A2(new_n2377_), .B(new_n2764_), .ZN(new_n3678_));
  OAI21_X1   g3293(.A1(new_n3678_), .A2(new_n1167_), .B(new_n1176_), .ZN(new_n3679_));
  AOI21_X1   g3294(.A1(new_n3679_), .A2(new_n2326_), .B(new_n2327_), .ZN(new_n3680_));
  OAI21_X1   g3295(.A1(new_n3680_), .A2(new_n1203_), .B(new_n1212_), .ZN(new_n3681_));
  AOI21_X1   g3296(.A1(new_n3681_), .A2(new_n2324_), .B(new_n2325_), .ZN(new_n3682_));
  OAI21_X1   g3297(.A1(new_n3682_), .A2(new_n1239_), .B(new_n1248_), .ZN(new_n3683_));
  AOI21_X1   g3298(.A1(new_n3683_), .A2(new_n2322_), .B(new_n2323_), .ZN(new_n3684_));
  OAI21_X1   g3299(.A1(new_n3684_), .A2(new_n1275_), .B(new_n1284_), .ZN(new_n3685_));
  NAND2_X1   g3300(.A1(new_n1300_), .A2(new_n1005_), .ZN(new_n3686_));
  AOI21_X1   g3301(.A1(new_n3685_), .A2(new_n2320_), .B(new_n3686_), .ZN(\grant[85] ));
  NOR4_X1    g3302(.A1(new_n1306_), .A2(new_n2010_), .A3(new_n1883_), .A4(new_n1880_), .ZN(new_n3688_));
  OAI21_X1   g3303(.A1(new_n1891_), .A2(new_n3688_), .B(new_n1898_), .ZN(new_n3689_));
  AOI21_X1   g3304(.A1(new_n3689_), .A2(new_n2411_), .B(new_n2412_), .ZN(new_n3690_));
  OAI21_X1   g3305(.A1(new_n3690_), .A2(new_n1919_), .B(new_n1926_), .ZN(new_n3691_));
  AOI21_X1   g3306(.A1(new_n3691_), .A2(new_n2409_), .B(new_n2410_), .ZN(new_n3692_));
  OAI21_X1   g3307(.A1(new_n3692_), .A2(new_n1945_), .B(new_n2434_), .ZN(new_n3693_));
  AOI21_X1   g3308(.A1(new_n3693_), .A2(new_n2408_), .B(new_n2782_), .ZN(new_n3694_));
  OAI21_X1   g3309(.A1(new_n3694_), .A2(new_n1412_), .B(new_n1418_), .ZN(new_n3695_));
  AOI21_X1   g3310(.A1(new_n3695_), .A2(new_n2357_), .B(new_n2358_), .ZN(new_n3696_));
  OAI21_X1   g3311(.A1(new_n3696_), .A2(new_n1438_), .B(new_n1444_), .ZN(new_n3697_));
  AOI21_X1   g3312(.A1(new_n3697_), .A2(new_n2355_), .B(new_n2356_), .ZN(new_n3698_));
  OAI21_X1   g3313(.A1(new_n3698_), .A2(new_n1464_), .B(new_n1470_), .ZN(new_n3699_));
  AOI21_X1   g3314(.A1(new_n3699_), .A2(new_n2353_), .B(new_n2354_), .ZN(new_n3700_));
  OAI21_X1   g3315(.A1(new_n3700_), .A2(new_n1490_), .B(new_n1496_), .ZN(new_n3701_));
  NAND2_X1   g3316(.A1(new_n1505_), .A2(new_n1295_), .ZN(new_n3702_));
  AOI21_X1   g3317(.A1(new_n3701_), .A2(new_n2351_), .B(new_n3702_), .ZN(\grant[86] ));
  NOR4_X1    g3318(.A1(new_n1513_), .A2(new_n660_), .A3(new_n2012_), .A4(new_n2104_), .ZN(new_n3704_));
  OAI21_X1   g3319(.A1(new_n2017_), .A2(new_n3704_), .B(new_n2020_), .ZN(new_n3705_));
  AOI21_X1   g3320(.A1(new_n3705_), .A2(new_n2441_), .B(new_n2442_), .ZN(new_n3706_));
  OAI21_X1   g3321(.A1(new_n3706_), .A2(new_n2031_), .B(new_n2034_), .ZN(new_n3707_));
  AOI21_X1   g3322(.A1(new_n3707_), .A2(new_n2439_), .B(new_n2440_), .ZN(new_n3708_));
  OAI21_X1   g3323(.A1(new_n3708_), .A2(new_n2048_), .B(new_n2464_), .ZN(new_n3709_));
  AOI21_X1   g3324(.A1(new_n3709_), .A2(new_n2438_), .B(new_n2799_), .ZN(new_n3710_));
  OAI21_X1   g3325(.A1(new_n3710_), .A2(new_n1595_), .B(new_n1601_), .ZN(new_n3711_));
  AOI21_X1   g3326(.A1(new_n3711_), .A2(new_n2388_), .B(new_n2389_), .ZN(new_n3712_));
  OAI21_X1   g3327(.A1(new_n3712_), .A2(new_n1621_), .B(new_n1627_), .ZN(new_n3713_));
  AOI21_X1   g3328(.A1(new_n3713_), .A2(new_n2386_), .B(new_n2387_), .ZN(new_n3714_));
  OAI21_X1   g3329(.A1(new_n3714_), .A2(new_n1647_), .B(new_n1653_), .ZN(new_n3715_));
  AOI21_X1   g3330(.A1(new_n3715_), .A2(new_n2384_), .B(new_n2385_), .ZN(new_n3716_));
  OAI21_X1   g3331(.A1(new_n3716_), .A2(new_n1673_), .B(new_n1679_), .ZN(new_n3717_));
  NAND2_X1   g3332(.A1(new_n1688_), .A2(new_n652_), .ZN(new_n3718_));
  AOI21_X1   g3333(.A1(new_n3717_), .A2(new_n2382_), .B(new_n3718_), .ZN(\grant[87] ));
  NOR4_X1    g3334(.A1(new_n1696_), .A2(new_n1025_), .A3(new_n2106_), .A4(new_n2204_), .ZN(new_n3720_));
  OAI21_X1   g3335(.A1(new_n2110_), .A2(new_n3720_), .B(new_n2113_), .ZN(new_n3721_));
  AOI21_X1   g3336(.A1(new_n3721_), .A2(new_n2471_), .B(new_n2472_), .ZN(new_n3722_));
  OAI21_X1   g3337(.A1(new_n3722_), .A2(new_n2122_), .B(new_n2125_), .ZN(new_n3723_));
  AOI21_X1   g3338(.A1(new_n3723_), .A2(new_n2469_), .B(new_n2470_), .ZN(new_n3724_));
  OAI21_X1   g3339(.A1(new_n3724_), .A2(new_n2139_), .B(new_n2494_), .ZN(new_n3725_));
  AOI21_X1   g3340(.A1(new_n3725_), .A2(new_n2468_), .B(new_n2816_), .ZN(new_n3726_));
  OAI21_X1   g3341(.A1(new_n3726_), .A2(new_n1779_), .B(new_n1786_), .ZN(new_n3727_));
  AOI21_X1   g3342(.A1(new_n3727_), .A2(new_n2419_), .B(new_n2420_), .ZN(new_n3728_));
  OAI21_X1   g3343(.A1(new_n3728_), .A2(new_n1807_), .B(new_n1814_), .ZN(new_n3729_));
  AOI21_X1   g3344(.A1(new_n3729_), .A2(new_n2417_), .B(new_n2418_), .ZN(new_n3730_));
  OAI21_X1   g3345(.A1(new_n3730_), .A2(new_n1835_), .B(new_n1842_), .ZN(new_n3731_));
  AOI21_X1   g3346(.A1(new_n3731_), .A2(new_n2415_), .B(new_n2416_), .ZN(new_n3732_));
  OAI21_X1   g3347(.A1(new_n3732_), .A2(new_n1863_), .B(new_n1870_), .ZN(new_n3733_));
  NAND2_X1   g3348(.A1(new_n1879_), .A2(new_n1017_), .ZN(new_n3734_));
  AOI21_X1   g3349(.A1(new_n3733_), .A2(new_n2413_), .B(new_n3734_), .ZN(\grant[88] ));
  OAI21_X1   g3350(.A1(new_n656_), .A2(\priority[91] ), .B(new_n1882_), .ZN(new_n3736_));
  NOR3_X1    g3351(.A1(new_n3736_), .A2(new_n1888_), .A3(new_n2207_), .ZN(new_n3737_));
  OAI21_X1   g3352(.A1(new_n2211_), .A2(new_n3737_), .B(new_n2215_), .ZN(new_n3738_));
  AOI21_X1   g3353(.A1(new_n3738_), .A2(new_n2501_), .B(new_n2502_), .ZN(new_n3739_));
  OAI21_X1   g3354(.A1(new_n3739_), .A2(new_n2225_), .B(new_n2229_), .ZN(new_n3740_));
  AOI21_X1   g3355(.A1(new_n3740_), .A2(new_n2499_), .B(new_n2500_), .ZN(new_n3741_));
  OAI21_X1   g3356(.A1(new_n3741_), .A2(new_n2239_), .B(new_n2525_), .ZN(new_n3742_));
  AOI21_X1   g3357(.A1(new_n3742_), .A2(new_n2498_), .B(new_n2833_), .ZN(new_n3743_));
  OAI21_X1   g3358(.A1(new_n3743_), .A2(new_n1961_), .B(new_n1964_), .ZN(new_n3744_));
  AOI21_X1   g3359(.A1(new_n3744_), .A2(new_n2449_), .B(new_n2450_), .ZN(new_n3745_));
  OAI21_X1   g3360(.A1(new_n3745_), .A2(new_n1975_), .B(new_n1978_), .ZN(new_n3746_));
  AOI21_X1   g3361(.A1(new_n3746_), .A2(new_n2447_), .B(new_n2448_), .ZN(new_n3747_));
  OAI21_X1   g3362(.A1(new_n3747_), .A2(new_n1989_), .B(new_n1992_), .ZN(new_n3748_));
  AOI21_X1   g3363(.A1(new_n3748_), .A2(new_n2445_), .B(new_n2446_), .ZN(new_n3749_));
  OAI21_X1   g3364(.A1(new_n3749_), .A2(new_n2003_), .B(new_n2006_), .ZN(new_n3750_));
  NAND2_X1   g3365(.A1(new_n658_), .A2(new_n1304_), .ZN(new_n3751_));
  AOI21_X1   g3366(.A1(new_n3750_), .A2(new_n2443_), .B(new_n3751_), .ZN(\grant[89] ));
  AOI21_X1   g3367(.A1(new_n1694_), .A2(\priority[91] ), .B(\priority[92] ), .ZN(new_n3753_));
  NOR4_X1    g3368(.A1(new_n668_), .A2(new_n670_), .A3(new_n674_), .A4(new_n3753_), .ZN(new_n3754_));
  OAI21_X1   g3369(.A1(new_n691_), .A2(new_n3754_), .B(new_n704_), .ZN(new_n3755_));
  AOI21_X1   g3370(.A1(new_n3755_), .A2(new_n719_), .B(new_n733_), .ZN(new_n3756_));
  OAI21_X1   g3371(.A1(new_n3756_), .A2(new_n747_), .B(new_n760_), .ZN(new_n3757_));
  AOI21_X1   g3372(.A1(new_n3757_), .A2(new_n775_), .B(new_n2530_), .ZN(new_n3758_));
  OAI21_X1   g3373(.A1(new_n3758_), .A2(new_n2275_), .B(new_n2545_), .ZN(new_n3759_));
  AOI21_X1   g3374(.A1(new_n3759_), .A2(new_n2529_), .B(new_n2851_), .ZN(new_n3760_));
  OAI21_X1   g3375(.A1(new_n3760_), .A2(new_n2062_), .B(new_n2065_), .ZN(new_n3761_));
  AOI21_X1   g3376(.A1(new_n3761_), .A2(new_n2479_), .B(new_n2480_), .ZN(new_n3762_));
  OAI21_X1   g3377(.A1(new_n3762_), .A2(new_n2074_), .B(new_n2077_), .ZN(new_n3763_));
  AOI21_X1   g3378(.A1(new_n3763_), .A2(new_n2477_), .B(new_n2478_), .ZN(new_n3764_));
  OAI21_X1   g3379(.A1(new_n3764_), .A2(new_n2086_), .B(new_n2089_), .ZN(new_n3765_));
  AOI21_X1   g3380(.A1(new_n3765_), .A2(new_n2475_), .B(new_n2476_), .ZN(new_n3766_));
  OAI21_X1   g3381(.A1(new_n3766_), .A2(new_n2098_), .B(new_n2101_), .ZN(new_n3767_));
  NAND2_X1   g3382(.A1(new_n1023_), .A2(new_n1511_), .ZN(new_n3768_));
  AOI21_X1   g3383(.A1(new_n3767_), .A2(new_n2473_), .B(new_n3768_), .ZN(\grant[90] ));
  AOI21_X1   g3384(.A1(new_n1886_), .A2(\priority[92] ), .B(\priority[93] ), .ZN(new_n3770_));
  NOR4_X1    g3385(.A1(new_n1032_), .A2(new_n1034_), .A3(new_n1038_), .A4(new_n3770_), .ZN(new_n3771_));
  OAI21_X1   g3386(.A1(new_n1053_), .A2(new_n3771_), .B(new_n1065_), .ZN(new_n3772_));
  AOI21_X1   g3387(.A1(new_n3772_), .A2(new_n1078_), .B(new_n1091_), .ZN(new_n3773_));
  OAI21_X1   g3388(.A1(new_n3773_), .A2(new_n1103_), .B(new_n1115_), .ZN(new_n3774_));
  AOI21_X1   g3389(.A1(new_n3774_), .A2(new_n1128_), .B(new_n2550_), .ZN(new_n3775_));
  OAI21_X1   g3390(.A1(new_n3775_), .A2(new_n2311_), .B(new_n2565_), .ZN(new_n3776_));
  AOI21_X1   g3391(.A1(new_n3776_), .A2(new_n2549_), .B(new_n2869_), .ZN(new_n3777_));
  OAI21_X1   g3392(.A1(new_n3777_), .A2(new_n2155_), .B(new_n2159_), .ZN(new_n3778_));
  AOI21_X1   g3393(.A1(new_n3778_), .A2(new_n2509_), .B(new_n2510_), .ZN(new_n3779_));
  OAI21_X1   g3394(.A1(new_n3779_), .A2(new_n2169_), .B(new_n2173_), .ZN(new_n3780_));
  AOI21_X1   g3395(.A1(new_n3780_), .A2(new_n2507_), .B(new_n2508_), .ZN(new_n3781_));
  OAI21_X1   g3396(.A1(new_n3781_), .A2(new_n2183_), .B(new_n2187_), .ZN(new_n3782_));
  AOI21_X1   g3397(.A1(new_n3782_), .A2(new_n2505_), .B(new_n2506_), .ZN(new_n3783_));
  OAI21_X1   g3398(.A1(new_n3783_), .A2(new_n2197_), .B(new_n2201_), .ZN(new_n3784_));
  NAND2_X1   g3399(.A1(new_n1309_), .A2(new_n1694_), .ZN(new_n3785_));
  AOI21_X1   g3400(.A1(new_n3784_), .A2(new_n2503_), .B(new_n3785_), .ZN(\grant[91] ));
  OAI21_X1   g3401(.A1(new_n1514_), .A2(\priority[94] ), .B(new_n2206_), .ZN(new_n3787_));
  NOR3_X1    g3402(.A1(new_n3787_), .A2(new_n1315_), .A3(new_n1317_), .ZN(new_n3788_));
  OAI21_X1   g3403(.A1(new_n1330_), .A2(new_n3788_), .B(new_n1338_), .ZN(new_n3789_));
  AOI21_X1   g3404(.A1(new_n3789_), .A2(new_n1348_), .B(new_n1357_), .ZN(new_n3790_));
  OAI21_X1   g3405(.A1(new_n3790_), .A2(new_n1366_), .B(new_n1374_), .ZN(new_n3791_));
  AOI21_X1   g3406(.A1(new_n3791_), .A2(new_n1386_), .B(new_n2569_), .ZN(new_n3792_));
  OAI21_X1   g3407(.A1(new_n3792_), .A2(new_n411_), .B(new_n424_), .ZN(new_n3793_));
  AOI21_X1   g3408(.A1(new_n3793_), .A2(new_n439_), .B(new_n453_), .ZN(new_n3794_));
  OAI21_X1   g3409(.A1(new_n3794_), .A2(new_n467_), .B(new_n480_), .ZN(new_n3795_));
  AOI21_X1   g3410(.A1(new_n3795_), .A2(new_n495_), .B(new_n509_), .ZN(new_n3796_));
  OAI21_X1   g3411(.A1(new_n3796_), .A2(new_n523_), .B(new_n536_), .ZN(new_n3797_));
  AOI21_X1   g3412(.A1(new_n3797_), .A2(new_n551_), .B(new_n565_), .ZN(new_n3798_));
  OAI21_X1   g3413(.A1(new_n3798_), .A2(new_n579_), .B(new_n592_), .ZN(new_n3799_));
  AOI21_X1   g3414(.A1(new_n3799_), .A2(new_n607_), .B(new_n621_), .ZN(new_n3800_));
  OAI21_X1   g3415(.A1(new_n3800_), .A2(new_n635_), .B(new_n648_), .ZN(new_n3801_));
  NAND2_X1   g3416(.A1(new_n672_), .A2(new_n1886_), .ZN(new_n3802_));
  AOI21_X1   g3417(.A1(new_n3801_), .A2(new_n663_), .B(new_n3802_), .ZN(\grant[92] ));
  AOI21_X1   g3418(.A1(new_n1030_), .A2(\priority[94] ), .B(\priority[95] ), .ZN(new_n3804_));
  NOR4_X1    g3419(.A1(new_n683_), .A2(new_n1519_), .A3(new_n1521_), .A4(new_n3804_), .ZN(new_n3805_));
  OAI21_X1   g3420(.A1(new_n1530_), .A2(new_n3805_), .B(new_n1535_), .ZN(new_n3806_));
  AOI21_X1   g3421(.A1(new_n3806_), .A2(new_n1543_), .B(new_n1549_), .ZN(new_n3807_));
  OAI21_X1   g3422(.A1(new_n3807_), .A2(new_n1556_), .B(new_n1561_), .ZN(new_n3808_));
  AOI21_X1   g3423(.A1(new_n3808_), .A2(new_n1570_), .B(new_n2587_), .ZN(new_n3809_));
  OAI21_X1   g3424(.A1(new_n3809_), .A2(new_n803_), .B(new_n815_), .ZN(new_n3810_));
  AOI21_X1   g3425(.A1(new_n3810_), .A2(new_n828_), .B(new_n841_), .ZN(new_n3811_));
  OAI21_X1   g3426(.A1(new_n3811_), .A2(new_n853_), .B(new_n865_), .ZN(new_n3812_));
  AOI21_X1   g3427(.A1(new_n3812_), .A2(new_n878_), .B(new_n891_), .ZN(new_n3813_));
  OAI21_X1   g3428(.A1(new_n3813_), .A2(new_n903_), .B(new_n915_), .ZN(new_n3814_));
  AOI21_X1   g3429(.A1(new_n3814_), .A2(new_n928_), .B(new_n941_), .ZN(new_n3815_));
  OAI21_X1   g3430(.A1(new_n3815_), .A2(new_n953_), .B(new_n965_), .ZN(new_n3816_));
  AOI21_X1   g3431(.A1(new_n3816_), .A2(new_n978_), .B(new_n991_), .ZN(new_n3817_));
  OAI21_X1   g3432(.A1(new_n3817_), .A2(new_n1003_), .B(new_n1015_), .ZN(new_n3818_));
  NAND2_X1   g3433(.A1(new_n1036_), .A2(new_n666_), .ZN(new_n3819_));
  AOI21_X1   g3434(.A1(new_n3818_), .A2(new_n1028_), .B(new_n3819_), .ZN(\grant[93] ));
  AOI21_X1   g3435(.A1(new_n1313_), .A2(\priority[95] ), .B(\priority[96] ), .ZN(new_n3821_));
  NOR4_X1    g3436(.A1(new_n1045_), .A2(new_n1702_), .A3(new_n1704_), .A4(new_n3821_), .ZN(new_n3822_));
  OAI21_X1   g3437(.A1(new_n1713_), .A2(new_n3822_), .B(new_n1718_), .ZN(new_n3823_));
  AOI21_X1   g3438(.A1(new_n3823_), .A2(new_n1726_), .B(new_n1732_), .ZN(new_n3824_));
  OAI21_X1   g3439(.A1(new_n3824_), .A2(new_n1739_), .B(new_n1744_), .ZN(new_n3825_));
  AOI21_X1   g3440(.A1(new_n3825_), .A2(new_n1751_), .B(new_n2605_), .ZN(new_n3826_));
  OAI21_X1   g3441(.A1(new_n3826_), .A2(new_n1150_), .B(new_n1158_), .ZN(new_n3827_));
  AOI21_X1   g3442(.A1(new_n3827_), .A2(new_n1168_), .B(new_n1177_), .ZN(new_n3828_));
  OAI21_X1   g3443(.A1(new_n3828_), .A2(new_n1186_), .B(new_n1194_), .ZN(new_n3829_));
  AOI21_X1   g3444(.A1(new_n3829_), .A2(new_n1204_), .B(new_n1213_), .ZN(new_n3830_));
  OAI21_X1   g3445(.A1(new_n3830_), .A2(new_n1222_), .B(new_n1230_), .ZN(new_n3831_));
  AOI21_X1   g3446(.A1(new_n3831_), .A2(new_n1240_), .B(new_n1249_), .ZN(new_n3832_));
  OAI21_X1   g3447(.A1(new_n3832_), .A2(new_n1258_), .B(new_n1266_), .ZN(new_n3833_));
  AOI21_X1   g3448(.A1(new_n3833_), .A2(new_n1276_), .B(new_n1285_), .ZN(new_n3834_));
  OAI21_X1   g3449(.A1(new_n3834_), .A2(new_n1294_), .B(new_n1302_), .ZN(new_n3835_));
  NAND2_X1   g3450(.A1(new_n1318_), .A2(new_n1030_), .ZN(new_n3836_));
  AOI21_X1   g3451(.A1(new_n3835_), .A2(new_n1312_), .B(new_n3836_), .ZN(\grant[94] ));
  NOR4_X1    g3452(.A1(new_n1325_), .A2(new_n2016_), .A3(new_n1897_), .A4(new_n1894_), .ZN(new_n3838_));
  OAI21_X1   g3453(.A1(new_n1906_), .A2(new_n3838_), .B(new_n1912_), .ZN(new_n3839_));
  AOI21_X1   g3454(.A1(new_n3839_), .A2(new_n1920_), .B(new_n1927_), .ZN(new_n3840_));
  OAI21_X1   g3455(.A1(new_n3840_), .A2(new_n1934_), .B(new_n1939_), .ZN(new_n3841_));
  AOI21_X1   g3456(.A1(new_n3841_), .A2(new_n1946_), .B(new_n2623_), .ZN(new_n3842_));
  OAI21_X1   g3457(.A1(new_n3842_), .A2(new_n1400_), .B(new_n1405_), .ZN(new_n3843_));
  AOI21_X1   g3458(.A1(new_n3843_), .A2(new_n1413_), .B(new_n1419_), .ZN(new_n3844_));
  OAI21_X1   g3459(.A1(new_n3844_), .A2(new_n1426_), .B(new_n1431_), .ZN(new_n3845_));
  AOI21_X1   g3460(.A1(new_n3845_), .A2(new_n1439_), .B(new_n1445_), .ZN(new_n3846_));
  OAI21_X1   g3461(.A1(new_n3846_), .A2(new_n1452_), .B(new_n1457_), .ZN(new_n3847_));
  AOI21_X1   g3462(.A1(new_n3847_), .A2(new_n1465_), .B(new_n1471_), .ZN(new_n3848_));
  OAI21_X1   g3463(.A1(new_n3848_), .A2(new_n1478_), .B(new_n1483_), .ZN(new_n3849_));
  AOI21_X1   g3464(.A1(new_n3849_), .A2(new_n1491_), .B(new_n1497_), .ZN(new_n3850_));
  OAI21_X1   g3465(.A1(new_n3850_), .A2(new_n1504_), .B(new_n1509_), .ZN(new_n3851_));
  NAND2_X1   g3466(.A1(new_n1518_), .A2(new_n1313_), .ZN(new_n3852_));
  AOI21_X1   g3467(.A1(new_n3851_), .A2(new_n1517_), .B(new_n3852_), .ZN(\grant[95] ));
  NOR4_X1    g3468(.A1(new_n1527_), .A2(new_n689_), .A3(new_n2019_), .A4(new_n2109_), .ZN(new_n3854_));
  OAI21_X1   g3469(.A1(new_n2025_), .A2(new_n3854_), .B(new_n2027_), .ZN(new_n3855_));
  AOI21_X1   g3470(.A1(new_n3855_), .A2(new_n2032_), .B(new_n2035_), .ZN(new_n3856_));
  OAI21_X1   g3471(.A1(new_n3856_), .A2(new_n2039_), .B(new_n2041_), .ZN(new_n3857_));
  AOI21_X1   g3472(.A1(new_n3857_), .A2(new_n2049_), .B(new_n2640_), .ZN(new_n3858_));
  OAI21_X1   g3473(.A1(new_n3858_), .A2(new_n1583_), .B(new_n1588_), .ZN(new_n3859_));
  AOI21_X1   g3474(.A1(new_n3859_), .A2(new_n1596_), .B(new_n1602_), .ZN(new_n3860_));
  OAI21_X1   g3475(.A1(new_n3860_), .A2(new_n1609_), .B(new_n1614_), .ZN(new_n3861_));
  AOI21_X1   g3476(.A1(new_n3861_), .A2(new_n1622_), .B(new_n1628_), .ZN(new_n3862_));
  OAI21_X1   g3477(.A1(new_n3862_), .A2(new_n1635_), .B(new_n1640_), .ZN(new_n3863_));
  AOI21_X1   g3478(.A1(new_n3863_), .A2(new_n1648_), .B(new_n1654_), .ZN(new_n3864_));
  OAI21_X1   g3479(.A1(new_n3864_), .A2(new_n1661_), .B(new_n1666_), .ZN(new_n3865_));
  AOI21_X1   g3480(.A1(new_n3865_), .A2(new_n1674_), .B(new_n1680_), .ZN(new_n3866_));
  OAI21_X1   g3481(.A1(new_n3866_), .A2(new_n1687_), .B(new_n1692_), .ZN(new_n3867_));
  NAND2_X1   g3482(.A1(new_n1701_), .A2(new_n681_), .ZN(new_n3868_));
  AOI21_X1   g3483(.A1(new_n3867_), .A2(new_n1700_), .B(new_n3868_), .ZN(\grant[96] ));
  NOR4_X1    g3484(.A1(new_n1710_), .A2(new_n1051_), .A3(new_n2112_), .A4(new_n2210_), .ZN(new_n3870_));
  OAI21_X1   g3485(.A1(new_n2117_), .A2(new_n3870_), .B(new_n2119_), .ZN(new_n3871_));
  AOI21_X1   g3486(.A1(new_n3871_), .A2(new_n2123_), .B(new_n2126_), .ZN(new_n3872_));
  OAI21_X1   g3487(.A1(new_n3872_), .A2(new_n2129_), .B(new_n2132_), .ZN(new_n3873_));
  AOI21_X1   g3488(.A1(new_n3873_), .A2(new_n2140_), .B(new_n2657_), .ZN(new_n3874_));
  OAI21_X1   g3489(.A1(new_n3874_), .A2(new_n1766_), .B(new_n1772_), .ZN(new_n3875_));
  AOI21_X1   g3490(.A1(new_n3875_), .A2(new_n1780_), .B(new_n1787_), .ZN(new_n3876_));
  OAI21_X1   g3491(.A1(new_n3876_), .A2(new_n1794_), .B(new_n1800_), .ZN(new_n3877_));
  AOI21_X1   g3492(.A1(new_n3877_), .A2(new_n1808_), .B(new_n1815_), .ZN(new_n3878_));
  OAI21_X1   g3493(.A1(new_n3878_), .A2(new_n1822_), .B(new_n1828_), .ZN(new_n3879_));
  AOI21_X1   g3494(.A1(new_n3879_), .A2(new_n1836_), .B(new_n1843_), .ZN(new_n3880_));
  OAI21_X1   g3495(.A1(new_n3880_), .A2(new_n1850_), .B(new_n1856_), .ZN(new_n3881_));
  AOI21_X1   g3496(.A1(new_n3881_), .A2(new_n1864_), .B(new_n1871_), .ZN(new_n3882_));
  OAI21_X1   g3497(.A1(new_n3882_), .A2(new_n1878_), .B(new_n1884_), .ZN(new_n3883_));
  NAND2_X1   g3498(.A1(new_n1893_), .A2(new_n1043_), .ZN(new_n3884_));
  AOI21_X1   g3499(.A1(new_n3883_), .A2(new_n1892_), .B(new_n3884_), .ZN(\grant[97] ));
  OAI21_X1   g3500(.A1(new_n685_), .A2(\priority[100] ), .B(new_n1896_), .ZN(new_n3886_));
  NOR3_X1    g3501(.A1(new_n3886_), .A2(new_n1903_), .A3(new_n2214_), .ZN(new_n3887_));
  OAI21_X1   g3502(.A1(new_n2219_), .A2(new_n3887_), .B(new_n2222_), .ZN(new_n3888_));
  AOI21_X1   g3503(.A1(new_n3888_), .A2(new_n2226_), .B(new_n2230_), .ZN(new_n3889_));
  OAI21_X1   g3504(.A1(new_n3889_), .A2(new_n2233_), .B(new_n2235_), .ZN(new_n3890_));
  AOI21_X1   g3505(.A1(new_n3890_), .A2(new_n2240_), .B(new_n2674_), .ZN(new_n3891_));
  OAI21_X1   g3506(.A1(new_n3891_), .A2(new_n1955_), .B(new_n1957_), .ZN(new_n3892_));
  AOI21_X1   g3507(.A1(new_n3892_), .A2(new_n1962_), .B(new_n1965_), .ZN(new_n3893_));
  OAI21_X1   g3508(.A1(new_n3893_), .A2(new_n1969_), .B(new_n1971_), .ZN(new_n3894_));
  AOI21_X1   g3509(.A1(new_n3894_), .A2(new_n1976_), .B(new_n1979_), .ZN(new_n3895_));
  OAI21_X1   g3510(.A1(new_n3895_), .A2(new_n1983_), .B(new_n1985_), .ZN(new_n3896_));
  AOI21_X1   g3511(.A1(new_n3896_), .A2(new_n1990_), .B(new_n1993_), .ZN(new_n3897_));
  OAI21_X1   g3512(.A1(new_n3897_), .A2(new_n1997_), .B(new_n1999_), .ZN(new_n3898_));
  AOI21_X1   g3513(.A1(new_n3898_), .A2(new_n2004_), .B(new_n2007_), .ZN(new_n3899_));
  OAI21_X1   g3514(.A1(new_n3899_), .A2(new_n2011_), .B(new_n2013_), .ZN(new_n3900_));
  NAND2_X1   g3515(.A1(new_n687_), .A2(new_n1323_), .ZN(new_n3901_));
  AOI21_X1   g3516(.A1(new_n3900_), .A2(new_n2018_), .B(new_n3901_), .ZN(\grant[98] ));
  AOI21_X1   g3517(.A1(new_n1708_), .A2(\priority[100] ), .B(\priority[101] ), .ZN(new_n3903_));
  NOR4_X1    g3518(.A1(new_n696_), .A2(new_n698_), .A3(new_n702_), .A4(new_n3903_), .ZN(new_n3904_));
  OAI21_X1   g3519(.A1(new_n718_), .A2(new_n3904_), .B(new_n732_), .ZN(new_n3905_));
  AOI21_X1   g3520(.A1(new_n3905_), .A2(new_n2243_), .B(new_n2244_), .ZN(new_n3906_));
  OAI21_X1   g3521(.A1(new_n3906_), .A2(new_n774_), .B(new_n2270_), .ZN(new_n3907_));
  AOI21_X1   g3522(.A1(new_n3907_), .A2(new_n2276_), .B(new_n2692_), .ZN(new_n3908_));
  OAI21_X1   g3523(.A1(new_n3908_), .A2(new_n2057_), .B(new_n2059_), .ZN(new_n3909_));
  AOI21_X1   g3524(.A1(new_n3909_), .A2(new_n2063_), .B(new_n2066_), .ZN(new_n3910_));
  OAI21_X1   g3525(.A1(new_n3910_), .A2(new_n2069_), .B(new_n2071_), .ZN(new_n3911_));
  AOI21_X1   g3526(.A1(new_n3911_), .A2(new_n2075_), .B(new_n2078_), .ZN(new_n3912_));
  OAI21_X1   g3527(.A1(new_n3912_), .A2(new_n2081_), .B(new_n2083_), .ZN(new_n3913_));
  AOI21_X1   g3528(.A1(new_n3913_), .A2(new_n2087_), .B(new_n2090_), .ZN(new_n3914_));
  OAI21_X1   g3529(.A1(new_n3914_), .A2(new_n2093_), .B(new_n2095_), .ZN(new_n3915_));
  AOI21_X1   g3530(.A1(new_n3915_), .A2(new_n2099_), .B(new_n2102_), .ZN(new_n3916_));
  OAI21_X1   g3531(.A1(new_n3916_), .A2(new_n2105_), .B(new_n2107_), .ZN(new_n3917_));
  NAND2_X1   g3532(.A1(new_n1049_), .A2(new_n1525_), .ZN(new_n3918_));
  AOI21_X1   g3533(.A1(new_n3917_), .A2(new_n2111_), .B(new_n3918_), .ZN(\grant[99] ));
  AOI21_X1   g3534(.A1(new_n1901_), .A2(\priority[101] ), .B(\priority[102] ), .ZN(new_n3920_));
  NOR4_X1    g3535(.A1(new_n1057_), .A2(new_n1059_), .A3(new_n1063_), .A4(new_n3920_), .ZN(new_n3921_));
  OAI21_X1   g3536(.A1(new_n1077_), .A2(new_n3921_), .B(new_n1090_), .ZN(new_n3922_));
  AOI21_X1   g3537(.A1(new_n3922_), .A2(new_n2279_), .B(new_n2280_), .ZN(new_n3923_));
  OAI21_X1   g3538(.A1(new_n3923_), .A2(new_n1127_), .B(new_n2306_), .ZN(new_n3924_));
  AOI21_X1   g3539(.A1(new_n3924_), .A2(new_n2312_), .B(new_n2710_), .ZN(new_n3925_));
  OAI21_X1   g3540(.A1(new_n3925_), .A2(new_n2149_), .B(new_n2152_), .ZN(new_n3926_));
  AOI21_X1   g3541(.A1(new_n3926_), .A2(new_n2156_), .B(new_n2160_), .ZN(new_n3927_));
  OAI21_X1   g3542(.A1(new_n3927_), .A2(new_n2163_), .B(new_n2166_), .ZN(new_n3928_));
  AOI21_X1   g3543(.A1(new_n3928_), .A2(new_n2170_), .B(new_n2174_), .ZN(new_n3929_));
  OAI21_X1   g3544(.A1(new_n3929_), .A2(new_n2177_), .B(new_n2180_), .ZN(new_n3930_));
  AOI21_X1   g3545(.A1(new_n3930_), .A2(new_n2184_), .B(new_n2188_), .ZN(new_n3931_));
  OAI21_X1   g3546(.A1(new_n3931_), .A2(new_n2191_), .B(new_n2194_), .ZN(new_n3932_));
  AOI21_X1   g3547(.A1(new_n3932_), .A2(new_n2198_), .B(new_n2202_), .ZN(new_n3933_));
  OAI21_X1   g3548(.A1(new_n3933_), .A2(new_n2205_), .B(new_n2208_), .ZN(new_n3934_));
  NAND2_X1   g3549(.A1(new_n1328_), .A2(new_n1708_), .ZN(new_n3935_));
  AOI21_X1   g3550(.A1(new_n3934_), .A2(new_n2212_), .B(new_n3935_), .ZN(\grant[100] ));
  OAI21_X1   g3551(.A1(new_n1528_), .A2(\priority[103] ), .B(new_n2213_), .ZN(new_n3937_));
  NOR3_X1    g3552(.A1(new_n3937_), .A2(new_n1333_), .A3(new_n1335_), .ZN(new_n3938_));
  OAI21_X1   g3553(.A1(new_n1347_), .A2(new_n3938_), .B(new_n1356_), .ZN(new_n3939_));
  AOI21_X1   g3554(.A1(new_n3939_), .A2(new_n2316_), .B(new_n2317_), .ZN(new_n3940_));
  OAI21_X1   g3555(.A1(new_n3940_), .A2(new_n1385_), .B(new_n2342_), .ZN(new_n3941_));
  AOI21_X1   g3556(.A1(new_n3941_), .A2(new_n2315_), .B(new_n2728_), .ZN(new_n3942_));
  OAI21_X1   g3557(.A1(new_n3942_), .A2(new_n438_), .B(new_n452_), .ZN(new_n3943_));
  AOI21_X1   g3558(.A1(new_n3943_), .A2(new_n2253_), .B(new_n2254_), .ZN(new_n3944_));
  OAI21_X1   g3559(.A1(new_n3944_), .A2(new_n494_), .B(new_n508_), .ZN(new_n3945_));
  AOI21_X1   g3560(.A1(new_n3945_), .A2(new_n2251_), .B(new_n2252_), .ZN(new_n3946_));
  OAI21_X1   g3561(.A1(new_n3946_), .A2(new_n550_), .B(new_n564_), .ZN(new_n3947_));
  AOI21_X1   g3562(.A1(new_n3947_), .A2(new_n2249_), .B(new_n2250_), .ZN(new_n3948_));
  OAI21_X1   g3563(.A1(new_n3948_), .A2(new_n606_), .B(new_n620_), .ZN(new_n3949_));
  AOI21_X1   g3564(.A1(new_n3949_), .A2(new_n2247_), .B(new_n2248_), .ZN(new_n3950_));
  OAI21_X1   g3565(.A1(new_n3950_), .A2(new_n662_), .B(new_n676_), .ZN(new_n3951_));
  NAND2_X1   g3566(.A1(new_n700_), .A2(new_n1901_), .ZN(new_n3952_));
  AOI21_X1   g3567(.A1(new_n3951_), .A2(new_n2245_), .B(new_n3952_), .ZN(\grant[101] ));
  AOI21_X1   g3568(.A1(new_n1055_), .A2(\priority[103] ), .B(\priority[104] ), .ZN(new_n3954_));
  NOR4_X1    g3569(.A1(new_n710_), .A2(new_n1532_), .A3(new_n1534_), .A4(new_n3954_), .ZN(new_n3955_));
  OAI21_X1   g3570(.A1(new_n1542_), .A2(new_n3955_), .B(new_n1548_), .ZN(new_n3956_));
  AOI21_X1   g3571(.A1(new_n3956_), .A2(new_n2347_), .B(new_n2348_), .ZN(new_n3957_));
  OAI21_X1   g3572(.A1(new_n3957_), .A2(new_n1569_), .B(new_n2373_), .ZN(new_n3958_));
  AOI21_X1   g3573(.A1(new_n3958_), .A2(new_n2346_), .B(new_n2746_), .ZN(new_n3959_));
  OAI21_X1   g3574(.A1(new_n3959_), .A2(new_n827_), .B(new_n840_), .ZN(new_n3960_));
  AOI21_X1   g3575(.A1(new_n3960_), .A2(new_n2289_), .B(new_n2290_), .ZN(new_n3961_));
  OAI21_X1   g3576(.A1(new_n3961_), .A2(new_n877_), .B(new_n890_), .ZN(new_n3962_));
  AOI21_X1   g3577(.A1(new_n3962_), .A2(new_n2287_), .B(new_n2288_), .ZN(new_n3963_));
  OAI21_X1   g3578(.A1(new_n3963_), .A2(new_n927_), .B(new_n940_), .ZN(new_n3964_));
  AOI21_X1   g3579(.A1(new_n3964_), .A2(new_n2285_), .B(new_n2286_), .ZN(new_n3965_));
  OAI21_X1   g3580(.A1(new_n3965_), .A2(new_n977_), .B(new_n990_), .ZN(new_n3966_));
  AOI21_X1   g3581(.A1(new_n3966_), .A2(new_n2283_), .B(new_n2284_), .ZN(new_n3967_));
  OAI21_X1   g3582(.A1(new_n3967_), .A2(new_n1027_), .B(new_n1040_), .ZN(new_n3968_));
  NAND2_X1   g3583(.A1(new_n1061_), .A2(new_n694_), .ZN(new_n3969_));
  AOI21_X1   g3584(.A1(new_n3968_), .A2(new_n2281_), .B(new_n3969_), .ZN(\grant[102] ));
  AOI21_X1   g3585(.A1(new_n1331_), .A2(\priority[104] ), .B(\priority[105] ), .ZN(new_n3971_));
  NOR4_X1    g3586(.A1(new_n1069_), .A2(new_n1715_), .A3(new_n1717_), .A4(new_n3971_), .ZN(new_n3972_));
  OAI21_X1   g3587(.A1(new_n1725_), .A2(new_n3972_), .B(new_n1731_), .ZN(new_n3973_));
  AOI21_X1   g3588(.A1(new_n3973_), .A2(new_n2378_), .B(new_n2379_), .ZN(new_n3974_));
  OAI21_X1   g3589(.A1(new_n3974_), .A2(new_n1750_), .B(new_n2404_), .ZN(new_n3975_));
  AOI21_X1   g3590(.A1(new_n3975_), .A2(new_n2377_), .B(new_n2764_), .ZN(new_n3976_));
  OAI21_X1   g3591(.A1(new_n3976_), .A2(new_n1167_), .B(new_n1176_), .ZN(new_n3977_));
  AOI21_X1   g3592(.A1(new_n3977_), .A2(new_n2326_), .B(new_n2327_), .ZN(new_n3978_));
  OAI21_X1   g3593(.A1(new_n3978_), .A2(new_n1203_), .B(new_n1212_), .ZN(new_n3979_));
  AOI21_X1   g3594(.A1(new_n3979_), .A2(new_n2324_), .B(new_n2325_), .ZN(new_n3980_));
  OAI21_X1   g3595(.A1(new_n3980_), .A2(new_n1239_), .B(new_n1248_), .ZN(new_n3981_));
  AOI21_X1   g3596(.A1(new_n3981_), .A2(new_n2322_), .B(new_n2323_), .ZN(new_n3982_));
  OAI21_X1   g3597(.A1(new_n3982_), .A2(new_n1275_), .B(new_n1284_), .ZN(new_n3983_));
  AOI21_X1   g3598(.A1(new_n3983_), .A2(new_n2320_), .B(new_n2321_), .ZN(new_n3984_));
  OAI21_X1   g3599(.A1(new_n3984_), .A2(new_n1311_), .B(new_n1320_), .ZN(new_n3985_));
  NAND2_X1   g3600(.A1(new_n1336_), .A2(new_n1055_), .ZN(new_n3986_));
  AOI21_X1   g3601(.A1(new_n3985_), .A2(new_n2318_), .B(new_n3986_), .ZN(\grant[103] ));
  NOR4_X1    g3602(.A1(new_n1342_), .A2(new_n2024_), .A3(new_n1911_), .A4(new_n1908_), .ZN(new_n3988_));
  OAI21_X1   g3603(.A1(new_n1919_), .A2(new_n3988_), .B(new_n1926_), .ZN(new_n3989_));
  AOI21_X1   g3604(.A1(new_n3989_), .A2(new_n2409_), .B(new_n2410_), .ZN(new_n3990_));
  OAI21_X1   g3605(.A1(new_n3990_), .A2(new_n1945_), .B(new_n2434_), .ZN(new_n3991_));
  AOI21_X1   g3606(.A1(new_n3991_), .A2(new_n2408_), .B(new_n2782_), .ZN(new_n3992_));
  OAI21_X1   g3607(.A1(new_n3992_), .A2(new_n1412_), .B(new_n1418_), .ZN(new_n3993_));
  AOI21_X1   g3608(.A1(new_n3993_), .A2(new_n2357_), .B(new_n2358_), .ZN(new_n3994_));
  OAI21_X1   g3609(.A1(new_n3994_), .A2(new_n1438_), .B(new_n1444_), .ZN(new_n3995_));
  AOI21_X1   g3610(.A1(new_n3995_), .A2(new_n2355_), .B(new_n2356_), .ZN(new_n3996_));
  OAI21_X1   g3611(.A1(new_n3996_), .A2(new_n1464_), .B(new_n1470_), .ZN(new_n3997_));
  AOI21_X1   g3612(.A1(new_n3997_), .A2(new_n2353_), .B(new_n2354_), .ZN(new_n3998_));
  OAI21_X1   g3613(.A1(new_n3998_), .A2(new_n1490_), .B(new_n1496_), .ZN(new_n3999_));
  AOI21_X1   g3614(.A1(new_n3999_), .A2(new_n2351_), .B(new_n2352_), .ZN(new_n4000_));
  OAI21_X1   g3615(.A1(new_n4000_), .A2(new_n1516_), .B(new_n1522_), .ZN(new_n4001_));
  NAND2_X1   g3616(.A1(new_n1531_), .A2(new_n1331_), .ZN(new_n4002_));
  AOI21_X1   g3617(.A1(new_n4001_), .A2(new_n2349_), .B(new_n4002_), .ZN(\grant[104] ));
  NOR4_X1    g3618(.A1(new_n1539_), .A2(new_n716_), .A3(new_n2026_), .A4(new_n2116_), .ZN(new_n4004_));
  OAI21_X1   g3619(.A1(new_n2031_), .A2(new_n4004_), .B(new_n2034_), .ZN(new_n4005_));
  AOI21_X1   g3620(.A1(new_n4005_), .A2(new_n2439_), .B(new_n2440_), .ZN(new_n4006_));
  OAI21_X1   g3621(.A1(new_n4006_), .A2(new_n2048_), .B(new_n2464_), .ZN(new_n4007_));
  AOI21_X1   g3622(.A1(new_n4007_), .A2(new_n2438_), .B(new_n2799_), .ZN(new_n4008_));
  OAI21_X1   g3623(.A1(new_n4008_), .A2(new_n1595_), .B(new_n1601_), .ZN(new_n4009_));
  AOI21_X1   g3624(.A1(new_n4009_), .A2(new_n2388_), .B(new_n2389_), .ZN(new_n4010_));
  OAI21_X1   g3625(.A1(new_n4010_), .A2(new_n1621_), .B(new_n1627_), .ZN(new_n4011_));
  AOI21_X1   g3626(.A1(new_n4011_), .A2(new_n2386_), .B(new_n2387_), .ZN(new_n4012_));
  OAI21_X1   g3627(.A1(new_n4012_), .A2(new_n1647_), .B(new_n1653_), .ZN(new_n4013_));
  AOI21_X1   g3628(.A1(new_n4013_), .A2(new_n2384_), .B(new_n2385_), .ZN(new_n4014_));
  OAI21_X1   g3629(.A1(new_n4014_), .A2(new_n1673_), .B(new_n1679_), .ZN(new_n4015_));
  AOI21_X1   g3630(.A1(new_n4015_), .A2(new_n2382_), .B(new_n2383_), .ZN(new_n4016_));
  OAI21_X1   g3631(.A1(new_n4016_), .A2(new_n1699_), .B(new_n1705_), .ZN(new_n4017_));
  NAND2_X1   g3632(.A1(new_n1714_), .A2(new_n708_), .ZN(new_n4018_));
  AOI21_X1   g3633(.A1(new_n4017_), .A2(new_n2380_), .B(new_n4018_), .ZN(\grant[105] ));
  NOR4_X1    g3634(.A1(new_n1722_), .A2(new_n1075_), .A3(new_n2118_), .A4(new_n2218_), .ZN(new_n4020_));
  OAI21_X1   g3635(.A1(new_n2122_), .A2(new_n4020_), .B(new_n2125_), .ZN(new_n4021_));
  AOI21_X1   g3636(.A1(new_n4021_), .A2(new_n2469_), .B(new_n2470_), .ZN(new_n4022_));
  OAI21_X1   g3637(.A1(new_n4022_), .A2(new_n2139_), .B(new_n2494_), .ZN(new_n4023_));
  AOI21_X1   g3638(.A1(new_n4023_), .A2(new_n2468_), .B(new_n2816_), .ZN(new_n4024_));
  OAI21_X1   g3639(.A1(new_n4024_), .A2(new_n1779_), .B(new_n1786_), .ZN(new_n4025_));
  AOI21_X1   g3640(.A1(new_n4025_), .A2(new_n2419_), .B(new_n2420_), .ZN(new_n4026_));
  OAI21_X1   g3641(.A1(new_n4026_), .A2(new_n1807_), .B(new_n1814_), .ZN(new_n4027_));
  AOI21_X1   g3642(.A1(new_n4027_), .A2(new_n2417_), .B(new_n2418_), .ZN(new_n4028_));
  OAI21_X1   g3643(.A1(new_n4028_), .A2(new_n1835_), .B(new_n1842_), .ZN(new_n4029_));
  AOI21_X1   g3644(.A1(new_n4029_), .A2(new_n2415_), .B(new_n2416_), .ZN(new_n4030_));
  OAI21_X1   g3645(.A1(new_n4030_), .A2(new_n1863_), .B(new_n1870_), .ZN(new_n4031_));
  AOI21_X1   g3646(.A1(new_n4031_), .A2(new_n2413_), .B(new_n2414_), .ZN(new_n4032_));
  OAI21_X1   g3647(.A1(new_n4032_), .A2(new_n1891_), .B(new_n1898_), .ZN(new_n4033_));
  NAND2_X1   g3648(.A1(new_n1907_), .A2(new_n1067_), .ZN(new_n4034_));
  AOI21_X1   g3649(.A1(new_n4033_), .A2(new_n2411_), .B(new_n4034_), .ZN(\grant[106] ));
  OAI21_X1   g3650(.A1(new_n712_), .A2(\priority[109] ), .B(new_n1910_), .ZN(new_n4036_));
  NOR3_X1    g3651(.A1(new_n4036_), .A2(new_n1916_), .A3(new_n2221_), .ZN(new_n4037_));
  OAI21_X1   g3652(.A1(new_n2225_), .A2(new_n4037_), .B(new_n2229_), .ZN(new_n4038_));
  AOI21_X1   g3653(.A1(new_n4038_), .A2(new_n2499_), .B(new_n2500_), .ZN(new_n4039_));
  OAI21_X1   g3654(.A1(new_n4039_), .A2(new_n2239_), .B(new_n2525_), .ZN(new_n4040_));
  AOI21_X1   g3655(.A1(new_n4040_), .A2(new_n2498_), .B(new_n2833_), .ZN(new_n4041_));
  OAI21_X1   g3656(.A1(new_n4041_), .A2(new_n1961_), .B(new_n1964_), .ZN(new_n4042_));
  AOI21_X1   g3657(.A1(new_n4042_), .A2(new_n2449_), .B(new_n2450_), .ZN(new_n4043_));
  OAI21_X1   g3658(.A1(new_n4043_), .A2(new_n1975_), .B(new_n1978_), .ZN(new_n4044_));
  AOI21_X1   g3659(.A1(new_n4044_), .A2(new_n2447_), .B(new_n2448_), .ZN(new_n4045_));
  OAI21_X1   g3660(.A1(new_n4045_), .A2(new_n1989_), .B(new_n1992_), .ZN(new_n4046_));
  AOI21_X1   g3661(.A1(new_n4046_), .A2(new_n2445_), .B(new_n2446_), .ZN(new_n4047_));
  OAI21_X1   g3662(.A1(new_n4047_), .A2(new_n2003_), .B(new_n2006_), .ZN(new_n4048_));
  AOI21_X1   g3663(.A1(new_n4048_), .A2(new_n2443_), .B(new_n2444_), .ZN(new_n4049_));
  OAI21_X1   g3664(.A1(new_n4049_), .A2(new_n2017_), .B(new_n2020_), .ZN(new_n4050_));
  NAND2_X1   g3665(.A1(new_n714_), .A2(new_n1340_), .ZN(new_n4051_));
  AOI21_X1   g3666(.A1(new_n4050_), .A2(new_n2441_), .B(new_n4051_), .ZN(\grant[107] ));
  AOI21_X1   g3667(.A1(new_n1720_), .A2(\priority[109] ), .B(\priority[110] ), .ZN(new_n4053_));
  NOR4_X1    g3668(.A1(new_n724_), .A2(new_n726_), .A3(new_n730_), .A4(new_n4053_), .ZN(new_n4054_));
  OAI21_X1   g3669(.A1(new_n747_), .A2(new_n4054_), .B(new_n760_), .ZN(new_n4055_));
  AOI21_X1   g3670(.A1(new_n4055_), .A2(new_n775_), .B(new_n2530_), .ZN(new_n4056_));
  OAI21_X1   g3671(.A1(new_n4056_), .A2(new_n2275_), .B(new_n2545_), .ZN(new_n4057_));
  AOI21_X1   g3672(.A1(new_n4057_), .A2(new_n2529_), .B(new_n2851_), .ZN(new_n4058_));
  OAI21_X1   g3673(.A1(new_n4058_), .A2(new_n2062_), .B(new_n2065_), .ZN(new_n4059_));
  AOI21_X1   g3674(.A1(new_n4059_), .A2(new_n2479_), .B(new_n2480_), .ZN(new_n4060_));
  OAI21_X1   g3675(.A1(new_n4060_), .A2(new_n2074_), .B(new_n2077_), .ZN(new_n4061_));
  AOI21_X1   g3676(.A1(new_n4061_), .A2(new_n2477_), .B(new_n2478_), .ZN(new_n4062_));
  OAI21_X1   g3677(.A1(new_n4062_), .A2(new_n2086_), .B(new_n2089_), .ZN(new_n4063_));
  AOI21_X1   g3678(.A1(new_n4063_), .A2(new_n2475_), .B(new_n2476_), .ZN(new_n4064_));
  OAI21_X1   g3679(.A1(new_n4064_), .A2(new_n2098_), .B(new_n2101_), .ZN(new_n4065_));
  AOI21_X1   g3680(.A1(new_n4065_), .A2(new_n2473_), .B(new_n2474_), .ZN(new_n4066_));
  OAI21_X1   g3681(.A1(new_n4066_), .A2(new_n2110_), .B(new_n2113_), .ZN(new_n4067_));
  NAND2_X1   g3682(.A1(new_n1073_), .A2(new_n1537_), .ZN(new_n4068_));
  AOI21_X1   g3683(.A1(new_n4067_), .A2(new_n2471_), .B(new_n4068_), .ZN(\grant[108] ));
  AOI21_X1   g3684(.A1(new_n1914_), .A2(\priority[110] ), .B(\priority[111] ), .ZN(new_n4070_));
  NOR4_X1    g3685(.A1(new_n1082_), .A2(new_n1084_), .A3(new_n1088_), .A4(new_n4070_), .ZN(new_n4071_));
  OAI21_X1   g3686(.A1(new_n1103_), .A2(new_n4071_), .B(new_n1115_), .ZN(new_n4072_));
  AOI21_X1   g3687(.A1(new_n4072_), .A2(new_n1128_), .B(new_n2550_), .ZN(new_n4073_));
  OAI21_X1   g3688(.A1(new_n4073_), .A2(new_n2311_), .B(new_n2565_), .ZN(new_n4074_));
  AOI21_X1   g3689(.A1(new_n4074_), .A2(new_n2549_), .B(new_n2869_), .ZN(new_n4075_));
  OAI21_X1   g3690(.A1(new_n4075_), .A2(new_n2155_), .B(new_n2159_), .ZN(new_n4076_));
  AOI21_X1   g3691(.A1(new_n4076_), .A2(new_n2509_), .B(new_n2510_), .ZN(new_n4077_));
  OAI21_X1   g3692(.A1(new_n4077_), .A2(new_n2169_), .B(new_n2173_), .ZN(new_n4078_));
  AOI21_X1   g3693(.A1(new_n4078_), .A2(new_n2507_), .B(new_n2508_), .ZN(new_n4079_));
  OAI21_X1   g3694(.A1(new_n4079_), .A2(new_n2183_), .B(new_n2187_), .ZN(new_n4080_));
  AOI21_X1   g3695(.A1(new_n4080_), .A2(new_n2505_), .B(new_n2506_), .ZN(new_n4081_));
  OAI21_X1   g3696(.A1(new_n4081_), .A2(new_n2197_), .B(new_n2201_), .ZN(new_n4082_));
  AOI21_X1   g3697(.A1(new_n4082_), .A2(new_n2503_), .B(new_n2504_), .ZN(new_n4083_));
  OAI21_X1   g3698(.A1(new_n4083_), .A2(new_n2211_), .B(new_n2215_), .ZN(new_n4084_));
  NAND2_X1   g3699(.A1(new_n1345_), .A2(new_n1720_), .ZN(new_n4085_));
  AOI21_X1   g3700(.A1(new_n4084_), .A2(new_n2501_), .B(new_n4085_), .ZN(\grant[109] ));
  OAI21_X1   g3701(.A1(new_n1540_), .A2(\priority[112] ), .B(new_n2220_), .ZN(new_n4087_));
  NOR3_X1    g3702(.A1(new_n4087_), .A2(new_n1351_), .A3(new_n1353_), .ZN(new_n4088_));
  OAI21_X1   g3703(.A1(new_n1366_), .A2(new_n4088_), .B(new_n1374_), .ZN(new_n4089_));
  AOI21_X1   g3704(.A1(new_n4089_), .A2(new_n1386_), .B(new_n2569_), .ZN(new_n4090_));
  OAI21_X1   g3705(.A1(new_n4090_), .A2(new_n411_), .B(new_n424_), .ZN(new_n4091_));
  AOI21_X1   g3706(.A1(new_n4091_), .A2(new_n439_), .B(new_n453_), .ZN(new_n4092_));
  OAI21_X1   g3707(.A1(new_n4092_), .A2(new_n467_), .B(new_n480_), .ZN(new_n4093_));
  AOI21_X1   g3708(.A1(new_n4093_), .A2(new_n495_), .B(new_n509_), .ZN(new_n4094_));
  OAI21_X1   g3709(.A1(new_n4094_), .A2(new_n523_), .B(new_n536_), .ZN(new_n4095_));
  AOI21_X1   g3710(.A1(new_n4095_), .A2(new_n551_), .B(new_n565_), .ZN(new_n4096_));
  OAI21_X1   g3711(.A1(new_n4096_), .A2(new_n579_), .B(new_n592_), .ZN(new_n4097_));
  AOI21_X1   g3712(.A1(new_n4097_), .A2(new_n607_), .B(new_n621_), .ZN(new_n4098_));
  OAI21_X1   g3713(.A1(new_n4098_), .A2(new_n635_), .B(new_n648_), .ZN(new_n4099_));
  AOI21_X1   g3714(.A1(new_n4099_), .A2(new_n663_), .B(new_n677_), .ZN(new_n4100_));
  OAI21_X1   g3715(.A1(new_n4100_), .A2(new_n691_), .B(new_n704_), .ZN(new_n4101_));
  NAND2_X1   g3716(.A1(new_n728_), .A2(new_n1914_), .ZN(new_n4102_));
  AOI21_X1   g3717(.A1(new_n4101_), .A2(new_n719_), .B(new_n4102_), .ZN(\grant[110] ));
  AOI21_X1   g3718(.A1(new_n1080_), .A2(\priority[112] ), .B(\priority[113] ), .ZN(new_n4104_));
  NOR4_X1    g3719(.A1(new_n739_), .A2(new_n1545_), .A3(new_n1547_), .A4(new_n4104_), .ZN(new_n4105_));
  OAI21_X1   g3720(.A1(new_n1556_), .A2(new_n4105_), .B(new_n1561_), .ZN(new_n4106_));
  AOI21_X1   g3721(.A1(new_n4106_), .A2(new_n1570_), .B(new_n2587_), .ZN(new_n4107_));
  OAI21_X1   g3722(.A1(new_n4107_), .A2(new_n803_), .B(new_n815_), .ZN(new_n4108_));
  AOI21_X1   g3723(.A1(new_n4108_), .A2(new_n828_), .B(new_n841_), .ZN(new_n4109_));
  OAI21_X1   g3724(.A1(new_n4109_), .A2(new_n853_), .B(new_n865_), .ZN(new_n4110_));
  AOI21_X1   g3725(.A1(new_n4110_), .A2(new_n878_), .B(new_n891_), .ZN(new_n4111_));
  OAI21_X1   g3726(.A1(new_n4111_), .A2(new_n903_), .B(new_n915_), .ZN(new_n4112_));
  AOI21_X1   g3727(.A1(new_n4112_), .A2(new_n928_), .B(new_n941_), .ZN(new_n4113_));
  OAI21_X1   g3728(.A1(new_n4113_), .A2(new_n953_), .B(new_n965_), .ZN(new_n4114_));
  AOI21_X1   g3729(.A1(new_n4114_), .A2(new_n978_), .B(new_n991_), .ZN(new_n4115_));
  OAI21_X1   g3730(.A1(new_n4115_), .A2(new_n1003_), .B(new_n1015_), .ZN(new_n4116_));
  AOI21_X1   g3731(.A1(new_n4116_), .A2(new_n1028_), .B(new_n1041_), .ZN(new_n4117_));
  OAI21_X1   g3732(.A1(new_n4117_), .A2(new_n1053_), .B(new_n1065_), .ZN(new_n4118_));
  NAND2_X1   g3733(.A1(new_n1086_), .A2(new_n722_), .ZN(new_n4119_));
  AOI21_X1   g3734(.A1(new_n4118_), .A2(new_n1078_), .B(new_n4119_), .ZN(\grant[111] ));
  AOI21_X1   g3735(.A1(new_n1349_), .A2(\priority[113] ), .B(\priority[114] ), .ZN(new_n4121_));
  NOR4_X1    g3736(.A1(new_n1095_), .A2(new_n1728_), .A3(new_n1730_), .A4(new_n4121_), .ZN(new_n4122_));
  OAI21_X1   g3737(.A1(new_n1739_), .A2(new_n4122_), .B(new_n1744_), .ZN(new_n4123_));
  AOI21_X1   g3738(.A1(new_n4123_), .A2(new_n1751_), .B(new_n2605_), .ZN(new_n4124_));
  OAI21_X1   g3739(.A1(new_n4124_), .A2(new_n1150_), .B(new_n1158_), .ZN(new_n4125_));
  AOI21_X1   g3740(.A1(new_n4125_), .A2(new_n1168_), .B(new_n1177_), .ZN(new_n4126_));
  OAI21_X1   g3741(.A1(new_n4126_), .A2(new_n1186_), .B(new_n1194_), .ZN(new_n4127_));
  AOI21_X1   g3742(.A1(new_n4127_), .A2(new_n1204_), .B(new_n1213_), .ZN(new_n4128_));
  OAI21_X1   g3743(.A1(new_n4128_), .A2(new_n1222_), .B(new_n1230_), .ZN(new_n4129_));
  AOI21_X1   g3744(.A1(new_n4129_), .A2(new_n1240_), .B(new_n1249_), .ZN(new_n4130_));
  OAI21_X1   g3745(.A1(new_n4130_), .A2(new_n1258_), .B(new_n1266_), .ZN(new_n4131_));
  AOI21_X1   g3746(.A1(new_n4131_), .A2(new_n1276_), .B(new_n1285_), .ZN(new_n4132_));
  OAI21_X1   g3747(.A1(new_n4132_), .A2(new_n1294_), .B(new_n1302_), .ZN(new_n4133_));
  AOI21_X1   g3748(.A1(new_n4133_), .A2(new_n1312_), .B(new_n1321_), .ZN(new_n4134_));
  OAI21_X1   g3749(.A1(new_n4134_), .A2(new_n1330_), .B(new_n1338_), .ZN(new_n4135_));
  NAND2_X1   g3750(.A1(new_n1354_), .A2(new_n1080_), .ZN(new_n4136_));
  AOI21_X1   g3751(.A1(new_n4135_), .A2(new_n1348_), .B(new_n4136_), .ZN(\grant[112] ));
  NOR4_X1    g3752(.A1(new_n1361_), .A2(new_n2030_), .A3(new_n1925_), .A4(new_n1922_), .ZN(new_n4138_));
  OAI21_X1   g3753(.A1(new_n1934_), .A2(new_n4138_), .B(new_n1939_), .ZN(new_n4139_));
  AOI21_X1   g3754(.A1(new_n4139_), .A2(new_n1946_), .B(new_n2623_), .ZN(new_n4140_));
  OAI21_X1   g3755(.A1(new_n4140_), .A2(new_n1400_), .B(new_n1405_), .ZN(new_n4141_));
  AOI21_X1   g3756(.A1(new_n4141_), .A2(new_n1413_), .B(new_n1419_), .ZN(new_n4142_));
  OAI21_X1   g3757(.A1(new_n4142_), .A2(new_n1426_), .B(new_n1431_), .ZN(new_n4143_));
  AOI21_X1   g3758(.A1(new_n4143_), .A2(new_n1439_), .B(new_n1445_), .ZN(new_n4144_));
  OAI21_X1   g3759(.A1(new_n4144_), .A2(new_n1452_), .B(new_n1457_), .ZN(new_n4145_));
  AOI21_X1   g3760(.A1(new_n4145_), .A2(new_n1465_), .B(new_n1471_), .ZN(new_n4146_));
  OAI21_X1   g3761(.A1(new_n4146_), .A2(new_n1478_), .B(new_n1483_), .ZN(new_n4147_));
  AOI21_X1   g3762(.A1(new_n4147_), .A2(new_n1491_), .B(new_n1497_), .ZN(new_n4148_));
  OAI21_X1   g3763(.A1(new_n4148_), .A2(new_n1504_), .B(new_n1509_), .ZN(new_n4149_));
  AOI21_X1   g3764(.A1(new_n4149_), .A2(new_n1517_), .B(new_n1523_), .ZN(new_n4150_));
  OAI21_X1   g3765(.A1(new_n4150_), .A2(new_n1530_), .B(new_n1535_), .ZN(new_n4151_));
  NAND2_X1   g3766(.A1(new_n1544_), .A2(new_n1349_), .ZN(new_n4152_));
  AOI21_X1   g3767(.A1(new_n4151_), .A2(new_n1543_), .B(new_n4152_), .ZN(\grant[113] ));
  NOR4_X1    g3768(.A1(new_n1553_), .A2(new_n745_), .A3(new_n2033_), .A4(new_n2121_), .ZN(new_n4154_));
  OAI21_X1   g3769(.A1(new_n2039_), .A2(new_n4154_), .B(new_n2041_), .ZN(new_n4155_));
  AOI21_X1   g3770(.A1(new_n4155_), .A2(new_n2049_), .B(new_n2640_), .ZN(new_n4156_));
  OAI21_X1   g3771(.A1(new_n4156_), .A2(new_n1583_), .B(new_n1588_), .ZN(new_n4157_));
  AOI21_X1   g3772(.A1(new_n4157_), .A2(new_n1596_), .B(new_n1602_), .ZN(new_n4158_));
  OAI21_X1   g3773(.A1(new_n4158_), .A2(new_n1609_), .B(new_n1614_), .ZN(new_n4159_));
  AOI21_X1   g3774(.A1(new_n4159_), .A2(new_n1622_), .B(new_n1628_), .ZN(new_n4160_));
  OAI21_X1   g3775(.A1(new_n4160_), .A2(new_n1635_), .B(new_n1640_), .ZN(new_n4161_));
  AOI21_X1   g3776(.A1(new_n4161_), .A2(new_n1648_), .B(new_n1654_), .ZN(new_n4162_));
  OAI21_X1   g3777(.A1(new_n4162_), .A2(new_n1661_), .B(new_n1666_), .ZN(new_n4163_));
  AOI21_X1   g3778(.A1(new_n4163_), .A2(new_n1674_), .B(new_n1680_), .ZN(new_n4164_));
  OAI21_X1   g3779(.A1(new_n4164_), .A2(new_n1687_), .B(new_n1692_), .ZN(new_n4165_));
  AOI21_X1   g3780(.A1(new_n4165_), .A2(new_n1700_), .B(new_n1706_), .ZN(new_n4166_));
  OAI21_X1   g3781(.A1(new_n4166_), .A2(new_n1713_), .B(new_n1718_), .ZN(new_n4167_));
  NAND2_X1   g3782(.A1(new_n1727_), .A2(new_n737_), .ZN(new_n4168_));
  AOI21_X1   g3783(.A1(new_n4167_), .A2(new_n1726_), .B(new_n4168_), .ZN(\grant[114] ));
  NOR4_X1    g3784(.A1(new_n1736_), .A2(new_n1101_), .A3(new_n2124_), .A4(new_n2224_), .ZN(new_n4170_));
  OAI21_X1   g3785(.A1(new_n2129_), .A2(new_n4170_), .B(new_n2132_), .ZN(new_n4171_));
  AOI21_X1   g3786(.A1(new_n4171_), .A2(new_n2140_), .B(new_n2657_), .ZN(new_n4172_));
  OAI21_X1   g3787(.A1(new_n4172_), .A2(new_n1766_), .B(new_n1772_), .ZN(new_n4173_));
  AOI21_X1   g3788(.A1(new_n4173_), .A2(new_n1780_), .B(new_n1787_), .ZN(new_n4174_));
  OAI21_X1   g3789(.A1(new_n4174_), .A2(new_n1794_), .B(new_n1800_), .ZN(new_n4175_));
  AOI21_X1   g3790(.A1(new_n4175_), .A2(new_n1808_), .B(new_n1815_), .ZN(new_n4176_));
  OAI21_X1   g3791(.A1(new_n4176_), .A2(new_n1822_), .B(new_n1828_), .ZN(new_n4177_));
  AOI21_X1   g3792(.A1(new_n4177_), .A2(new_n1836_), .B(new_n1843_), .ZN(new_n4178_));
  OAI21_X1   g3793(.A1(new_n4178_), .A2(new_n1850_), .B(new_n1856_), .ZN(new_n4179_));
  AOI21_X1   g3794(.A1(new_n4179_), .A2(new_n1864_), .B(new_n1871_), .ZN(new_n4180_));
  OAI21_X1   g3795(.A1(new_n4180_), .A2(new_n1878_), .B(new_n1884_), .ZN(new_n4181_));
  AOI21_X1   g3796(.A1(new_n4181_), .A2(new_n1892_), .B(new_n1899_), .ZN(new_n4182_));
  OAI21_X1   g3797(.A1(new_n4182_), .A2(new_n1906_), .B(new_n1912_), .ZN(new_n4183_));
  NAND2_X1   g3798(.A1(new_n1921_), .A2(new_n1093_), .ZN(new_n4184_));
  AOI21_X1   g3799(.A1(new_n4183_), .A2(new_n1920_), .B(new_n4184_), .ZN(\grant[115] ));
  OAI21_X1   g3800(.A1(new_n741_), .A2(\priority[118] ), .B(new_n1924_), .ZN(new_n4186_));
  NOR3_X1    g3801(.A1(new_n4186_), .A2(new_n1931_), .A3(new_n2228_), .ZN(new_n4187_));
  OAI21_X1   g3802(.A1(new_n2233_), .A2(new_n4187_), .B(new_n2235_), .ZN(new_n4188_));
  AOI21_X1   g3803(.A1(new_n4188_), .A2(new_n2240_), .B(new_n2674_), .ZN(new_n4189_));
  OAI21_X1   g3804(.A1(new_n4189_), .A2(new_n1955_), .B(new_n1957_), .ZN(new_n4190_));
  AOI21_X1   g3805(.A1(new_n4190_), .A2(new_n1962_), .B(new_n1965_), .ZN(new_n4191_));
  OAI21_X1   g3806(.A1(new_n4191_), .A2(new_n1969_), .B(new_n1971_), .ZN(new_n4192_));
  AOI21_X1   g3807(.A1(new_n4192_), .A2(new_n1976_), .B(new_n1979_), .ZN(new_n4193_));
  OAI21_X1   g3808(.A1(new_n4193_), .A2(new_n1983_), .B(new_n1985_), .ZN(new_n4194_));
  AOI21_X1   g3809(.A1(new_n4194_), .A2(new_n1990_), .B(new_n1993_), .ZN(new_n4195_));
  OAI21_X1   g3810(.A1(new_n4195_), .A2(new_n1997_), .B(new_n1999_), .ZN(new_n4196_));
  AOI21_X1   g3811(.A1(new_n4196_), .A2(new_n2004_), .B(new_n2007_), .ZN(new_n4197_));
  OAI21_X1   g3812(.A1(new_n4197_), .A2(new_n2011_), .B(new_n2013_), .ZN(new_n4198_));
  AOI21_X1   g3813(.A1(new_n4198_), .A2(new_n2018_), .B(new_n2021_), .ZN(new_n4199_));
  OAI21_X1   g3814(.A1(new_n4199_), .A2(new_n2025_), .B(new_n2027_), .ZN(new_n4200_));
  NAND2_X1   g3815(.A1(new_n743_), .A2(new_n1359_), .ZN(new_n4201_));
  AOI21_X1   g3816(.A1(new_n4200_), .A2(new_n2032_), .B(new_n4201_), .ZN(\grant[116] ));
  AOI21_X1   g3817(.A1(new_n1734_), .A2(\priority[118] ), .B(\priority[119] ), .ZN(new_n4203_));
  NOR4_X1    g3818(.A1(new_n752_), .A2(new_n754_), .A3(new_n758_), .A4(new_n4203_), .ZN(new_n4204_));
  OAI21_X1   g3819(.A1(new_n774_), .A2(new_n4204_), .B(new_n2270_), .ZN(new_n4205_));
  AOI21_X1   g3820(.A1(new_n4205_), .A2(new_n2276_), .B(new_n2692_), .ZN(new_n4206_));
  OAI21_X1   g3821(.A1(new_n4206_), .A2(new_n2057_), .B(new_n2059_), .ZN(new_n4207_));
  AOI21_X1   g3822(.A1(new_n4207_), .A2(new_n2063_), .B(new_n2066_), .ZN(new_n4208_));
  OAI21_X1   g3823(.A1(new_n4208_), .A2(new_n2069_), .B(new_n2071_), .ZN(new_n4209_));
  AOI21_X1   g3824(.A1(new_n4209_), .A2(new_n2075_), .B(new_n2078_), .ZN(new_n4210_));
  OAI21_X1   g3825(.A1(new_n4210_), .A2(new_n2081_), .B(new_n2083_), .ZN(new_n4211_));
  AOI21_X1   g3826(.A1(new_n4211_), .A2(new_n2087_), .B(new_n2090_), .ZN(new_n4212_));
  OAI21_X1   g3827(.A1(new_n4212_), .A2(new_n2093_), .B(new_n2095_), .ZN(new_n4213_));
  AOI21_X1   g3828(.A1(new_n4213_), .A2(new_n2099_), .B(new_n2102_), .ZN(new_n4214_));
  OAI21_X1   g3829(.A1(new_n4214_), .A2(new_n2105_), .B(new_n2107_), .ZN(new_n4215_));
  AOI21_X1   g3830(.A1(new_n4215_), .A2(new_n2111_), .B(new_n2114_), .ZN(new_n4216_));
  OAI21_X1   g3831(.A1(new_n4216_), .A2(new_n2117_), .B(new_n2119_), .ZN(new_n4217_));
  NAND2_X1   g3832(.A1(new_n1099_), .A2(new_n1551_), .ZN(new_n4218_));
  AOI21_X1   g3833(.A1(new_n4217_), .A2(new_n2123_), .B(new_n4218_), .ZN(\grant[117] ));
  AOI21_X1   g3834(.A1(new_n1929_), .A2(\priority[119] ), .B(\priority[120] ), .ZN(new_n4220_));
  NOR4_X1    g3835(.A1(new_n1107_), .A2(new_n1109_), .A3(new_n1113_), .A4(new_n4220_), .ZN(new_n4221_));
  OAI21_X1   g3836(.A1(new_n1127_), .A2(new_n4221_), .B(new_n2306_), .ZN(new_n4222_));
  AOI21_X1   g3837(.A1(new_n4222_), .A2(new_n2312_), .B(new_n2710_), .ZN(new_n4223_));
  OAI21_X1   g3838(.A1(new_n4223_), .A2(new_n2149_), .B(new_n2152_), .ZN(new_n4224_));
  AOI21_X1   g3839(.A1(new_n4224_), .A2(new_n2156_), .B(new_n2160_), .ZN(new_n4225_));
  OAI21_X1   g3840(.A1(new_n4225_), .A2(new_n2163_), .B(new_n2166_), .ZN(new_n4226_));
  AOI21_X1   g3841(.A1(new_n4226_), .A2(new_n2170_), .B(new_n2174_), .ZN(new_n4227_));
  OAI21_X1   g3842(.A1(new_n4227_), .A2(new_n2177_), .B(new_n2180_), .ZN(new_n4228_));
  AOI21_X1   g3843(.A1(new_n4228_), .A2(new_n2184_), .B(new_n2188_), .ZN(new_n4229_));
  OAI21_X1   g3844(.A1(new_n4229_), .A2(new_n2191_), .B(new_n2194_), .ZN(new_n4230_));
  AOI21_X1   g3845(.A1(new_n4230_), .A2(new_n2198_), .B(new_n2202_), .ZN(new_n4231_));
  OAI21_X1   g3846(.A1(new_n4231_), .A2(new_n2205_), .B(new_n2208_), .ZN(new_n4232_));
  AOI21_X1   g3847(.A1(new_n4232_), .A2(new_n2212_), .B(new_n2216_), .ZN(new_n4233_));
  OAI21_X1   g3848(.A1(new_n4233_), .A2(new_n2219_), .B(new_n2222_), .ZN(new_n4234_));
  NAND2_X1   g3849(.A1(new_n1364_), .A2(new_n1734_), .ZN(new_n4235_));
  AOI21_X1   g3850(.A1(new_n4234_), .A2(new_n2226_), .B(new_n4235_), .ZN(\grant[118] ));
  OAI21_X1   g3851(.A1(new_n1554_), .A2(\priority[121] ), .B(new_n2227_), .ZN(new_n4237_));
  NOR3_X1    g3852(.A1(new_n4237_), .A2(new_n1369_), .A3(new_n1371_), .ZN(new_n4238_));
  OAI21_X1   g3853(.A1(new_n1385_), .A2(new_n4238_), .B(new_n2342_), .ZN(new_n4239_));
  AOI21_X1   g3854(.A1(new_n4239_), .A2(new_n2315_), .B(new_n2728_), .ZN(new_n4240_));
  OAI21_X1   g3855(.A1(new_n4240_), .A2(new_n438_), .B(new_n452_), .ZN(new_n4241_));
  AOI21_X1   g3856(.A1(new_n4241_), .A2(new_n2253_), .B(new_n2254_), .ZN(new_n4242_));
  OAI21_X1   g3857(.A1(new_n4242_), .A2(new_n494_), .B(new_n508_), .ZN(new_n4243_));
  AOI21_X1   g3858(.A1(new_n4243_), .A2(new_n2251_), .B(new_n2252_), .ZN(new_n4244_));
  OAI21_X1   g3859(.A1(new_n4244_), .A2(new_n550_), .B(new_n564_), .ZN(new_n4245_));
  AOI21_X1   g3860(.A1(new_n4245_), .A2(new_n2249_), .B(new_n2250_), .ZN(new_n4246_));
  OAI21_X1   g3861(.A1(new_n4246_), .A2(new_n606_), .B(new_n620_), .ZN(new_n4247_));
  AOI21_X1   g3862(.A1(new_n4247_), .A2(new_n2247_), .B(new_n2248_), .ZN(new_n4248_));
  OAI21_X1   g3863(.A1(new_n4248_), .A2(new_n662_), .B(new_n676_), .ZN(new_n4249_));
  AOI21_X1   g3864(.A1(new_n4249_), .A2(new_n2245_), .B(new_n2246_), .ZN(new_n4250_));
  OAI21_X1   g3865(.A1(new_n4250_), .A2(new_n718_), .B(new_n732_), .ZN(new_n4251_));
  NAND2_X1   g3866(.A1(new_n756_), .A2(new_n1929_), .ZN(new_n4252_));
  AOI21_X1   g3867(.A1(new_n4251_), .A2(new_n2243_), .B(new_n4252_), .ZN(\grant[119] ));
  AOI21_X1   g3868(.A1(new_n1105_), .A2(\priority[121] ), .B(\priority[122] ), .ZN(new_n4254_));
  NOR4_X1    g3869(.A1(new_n766_), .A2(new_n1558_), .A3(new_n1560_), .A4(new_n4254_), .ZN(new_n4255_));
  OAI21_X1   g3870(.A1(new_n1569_), .A2(new_n4255_), .B(new_n2373_), .ZN(new_n4256_));
  AOI21_X1   g3871(.A1(new_n4256_), .A2(new_n2346_), .B(new_n2746_), .ZN(new_n4257_));
  OAI21_X1   g3872(.A1(new_n4257_), .A2(new_n827_), .B(new_n840_), .ZN(new_n4258_));
  AOI21_X1   g3873(.A1(new_n4258_), .A2(new_n2289_), .B(new_n2290_), .ZN(new_n4259_));
  OAI21_X1   g3874(.A1(new_n4259_), .A2(new_n877_), .B(new_n890_), .ZN(new_n4260_));
  AOI21_X1   g3875(.A1(new_n4260_), .A2(new_n2287_), .B(new_n2288_), .ZN(new_n4261_));
  OAI21_X1   g3876(.A1(new_n4261_), .A2(new_n927_), .B(new_n940_), .ZN(new_n4262_));
  AOI21_X1   g3877(.A1(new_n4262_), .A2(new_n2285_), .B(new_n2286_), .ZN(new_n4263_));
  OAI21_X1   g3878(.A1(new_n4263_), .A2(new_n977_), .B(new_n990_), .ZN(new_n4264_));
  AOI21_X1   g3879(.A1(new_n4264_), .A2(new_n2283_), .B(new_n2284_), .ZN(new_n4265_));
  OAI21_X1   g3880(.A1(new_n4265_), .A2(new_n1027_), .B(new_n1040_), .ZN(new_n4266_));
  AOI21_X1   g3881(.A1(new_n4266_), .A2(new_n2281_), .B(new_n2282_), .ZN(new_n4267_));
  OAI21_X1   g3882(.A1(new_n4267_), .A2(new_n1077_), .B(new_n1090_), .ZN(new_n4268_));
  NAND2_X1   g3883(.A1(new_n1111_), .A2(new_n750_), .ZN(new_n4269_));
  AOI21_X1   g3884(.A1(new_n4268_), .A2(new_n2279_), .B(new_n4269_), .ZN(\grant[120] ));
  AOI21_X1   g3885(.A1(new_n1367_), .A2(\priority[122] ), .B(\priority[123] ), .ZN(new_n4271_));
  NOR4_X1    g3886(.A1(new_n1119_), .A2(new_n1741_), .A3(new_n1743_), .A4(new_n4271_), .ZN(new_n4272_));
  OAI21_X1   g3887(.A1(new_n1750_), .A2(new_n4272_), .B(new_n2404_), .ZN(new_n4273_));
  AOI21_X1   g3888(.A1(new_n4273_), .A2(new_n2377_), .B(new_n2764_), .ZN(new_n4274_));
  OAI21_X1   g3889(.A1(new_n4274_), .A2(new_n1167_), .B(new_n1176_), .ZN(new_n4275_));
  AOI21_X1   g3890(.A1(new_n4275_), .A2(new_n2326_), .B(new_n2327_), .ZN(new_n4276_));
  OAI21_X1   g3891(.A1(new_n4276_), .A2(new_n1203_), .B(new_n1212_), .ZN(new_n4277_));
  AOI21_X1   g3892(.A1(new_n4277_), .A2(new_n2324_), .B(new_n2325_), .ZN(new_n4278_));
  OAI21_X1   g3893(.A1(new_n4278_), .A2(new_n1239_), .B(new_n1248_), .ZN(new_n4279_));
  AOI21_X1   g3894(.A1(new_n4279_), .A2(new_n2322_), .B(new_n2323_), .ZN(new_n4280_));
  OAI21_X1   g3895(.A1(new_n4280_), .A2(new_n1275_), .B(new_n1284_), .ZN(new_n4281_));
  AOI21_X1   g3896(.A1(new_n4281_), .A2(new_n2320_), .B(new_n2321_), .ZN(new_n4282_));
  OAI21_X1   g3897(.A1(new_n4282_), .A2(new_n1311_), .B(new_n1320_), .ZN(new_n4283_));
  AOI21_X1   g3898(.A1(new_n4283_), .A2(new_n2318_), .B(new_n2319_), .ZN(new_n4284_));
  OAI21_X1   g3899(.A1(new_n4284_), .A2(new_n1347_), .B(new_n1356_), .ZN(new_n4285_));
  NAND2_X1   g3900(.A1(new_n1372_), .A2(new_n1105_), .ZN(new_n4286_));
  AOI21_X1   g3901(.A1(new_n4285_), .A2(new_n2316_), .B(new_n4286_), .ZN(\grant[121] ));
  NOR4_X1    g3902(.A1(new_n1378_), .A2(new_n2038_), .A3(new_n1938_), .A4(new_n1936_), .ZN(new_n4288_));
  OAI21_X1   g3903(.A1(new_n1945_), .A2(new_n4288_), .B(new_n2434_), .ZN(new_n4289_));
  AOI21_X1   g3904(.A1(new_n4289_), .A2(new_n2408_), .B(new_n2782_), .ZN(new_n4290_));
  OAI21_X1   g3905(.A1(new_n4290_), .A2(new_n1412_), .B(new_n1418_), .ZN(new_n4291_));
  AOI21_X1   g3906(.A1(new_n4291_), .A2(new_n2357_), .B(new_n2358_), .ZN(new_n4292_));
  OAI21_X1   g3907(.A1(new_n4292_), .A2(new_n1438_), .B(new_n1444_), .ZN(new_n4293_));
  AOI21_X1   g3908(.A1(new_n4293_), .A2(new_n2355_), .B(new_n2356_), .ZN(new_n4294_));
  OAI21_X1   g3909(.A1(new_n4294_), .A2(new_n1464_), .B(new_n1470_), .ZN(new_n4295_));
  AOI21_X1   g3910(.A1(new_n4295_), .A2(new_n2353_), .B(new_n2354_), .ZN(new_n4296_));
  OAI21_X1   g3911(.A1(new_n4296_), .A2(new_n1490_), .B(new_n1496_), .ZN(new_n4297_));
  AOI21_X1   g3912(.A1(new_n4297_), .A2(new_n2351_), .B(new_n2352_), .ZN(new_n4298_));
  OAI21_X1   g3913(.A1(new_n4298_), .A2(new_n1516_), .B(new_n1522_), .ZN(new_n4299_));
  AOI21_X1   g3914(.A1(new_n4299_), .A2(new_n2349_), .B(new_n2350_), .ZN(new_n4300_));
  OAI21_X1   g3915(.A1(new_n4300_), .A2(new_n1542_), .B(new_n1548_), .ZN(new_n4301_));
  NAND2_X1   g3916(.A1(new_n1557_), .A2(new_n1367_), .ZN(new_n4302_));
  AOI21_X1   g3917(.A1(new_n4301_), .A2(new_n2347_), .B(new_n4302_), .ZN(\grant[122] ));
  NOR4_X1    g3918(.A1(new_n1564_), .A2(new_n2040_), .A3(new_n772_), .A4(new_n2128_), .ZN(new_n4304_));
  OAI21_X1   g3919(.A1(new_n2048_), .A2(new_n4304_), .B(new_n2464_), .ZN(new_n4305_));
  AOI21_X1   g3920(.A1(new_n4305_), .A2(new_n2438_), .B(new_n2799_), .ZN(new_n4306_));
  OAI21_X1   g3921(.A1(new_n4306_), .A2(new_n1595_), .B(new_n1601_), .ZN(new_n4307_));
  AOI21_X1   g3922(.A1(new_n4307_), .A2(new_n2388_), .B(new_n2389_), .ZN(new_n4308_));
  OAI21_X1   g3923(.A1(new_n4308_), .A2(new_n1621_), .B(new_n1627_), .ZN(new_n4309_));
  AOI21_X1   g3924(.A1(new_n4309_), .A2(new_n2386_), .B(new_n2387_), .ZN(new_n4310_));
  OAI21_X1   g3925(.A1(new_n4310_), .A2(new_n1647_), .B(new_n1653_), .ZN(new_n4311_));
  AOI21_X1   g3926(.A1(new_n4311_), .A2(new_n2384_), .B(new_n2385_), .ZN(new_n4312_));
  OAI21_X1   g3927(.A1(new_n4312_), .A2(new_n1673_), .B(new_n1679_), .ZN(new_n4313_));
  AOI21_X1   g3928(.A1(new_n4313_), .A2(new_n2382_), .B(new_n2383_), .ZN(new_n4314_));
  OAI21_X1   g3929(.A1(new_n4314_), .A2(new_n1699_), .B(new_n1705_), .ZN(new_n4315_));
  AOI21_X1   g3930(.A1(new_n4315_), .A2(new_n2380_), .B(new_n2381_), .ZN(new_n4316_));
  OAI21_X1   g3931(.A1(new_n4316_), .A2(new_n1725_), .B(new_n1731_), .ZN(new_n4317_));
  NAND2_X1   g3932(.A1(new_n1740_), .A2(new_n764_), .ZN(new_n4318_));
  AOI21_X1   g3933(.A1(new_n4317_), .A2(new_n2378_), .B(new_n4318_), .ZN(\grant[123] ));
  NOR4_X1    g3934(.A1(new_n1747_), .A2(new_n2131_), .A3(new_n1125_), .A4(new_n2232_), .ZN(new_n4320_));
  OAI21_X1   g3935(.A1(new_n2139_), .A2(new_n4320_), .B(new_n2494_), .ZN(new_n4321_));
  AOI21_X1   g3936(.A1(new_n4321_), .A2(new_n2468_), .B(new_n2816_), .ZN(new_n4322_));
  OAI21_X1   g3937(.A1(new_n4322_), .A2(new_n1779_), .B(new_n1786_), .ZN(new_n4323_));
  AOI21_X1   g3938(.A1(new_n4323_), .A2(new_n2419_), .B(new_n2420_), .ZN(new_n4324_));
  OAI21_X1   g3939(.A1(new_n4324_), .A2(new_n1807_), .B(new_n1814_), .ZN(new_n4325_));
  AOI21_X1   g3940(.A1(new_n4325_), .A2(new_n2417_), .B(new_n2418_), .ZN(new_n4326_));
  OAI21_X1   g3941(.A1(new_n4326_), .A2(new_n1835_), .B(new_n1842_), .ZN(new_n4327_));
  AOI21_X1   g3942(.A1(new_n4327_), .A2(new_n2415_), .B(new_n2416_), .ZN(new_n4328_));
  OAI21_X1   g3943(.A1(new_n4328_), .A2(new_n1863_), .B(new_n1870_), .ZN(new_n4329_));
  AOI21_X1   g3944(.A1(new_n4329_), .A2(new_n2413_), .B(new_n2414_), .ZN(new_n4330_));
  OAI21_X1   g3945(.A1(new_n4330_), .A2(new_n1891_), .B(new_n1898_), .ZN(new_n4331_));
  AOI21_X1   g3946(.A1(new_n4331_), .A2(new_n2411_), .B(new_n2412_), .ZN(new_n4332_));
  OAI21_X1   g3947(.A1(new_n4332_), .A2(new_n1919_), .B(new_n1926_), .ZN(new_n4333_));
  NAND2_X1   g3948(.A1(new_n1935_), .A2(new_n1117_), .ZN(new_n4334_));
  AOI21_X1   g3949(.A1(new_n4333_), .A2(new_n2409_), .B(new_n4334_), .ZN(\grant[124] ));
  INV_X1     g3950(.I(\req[126] ), .ZN(new_n4336_));
  AOI21_X1   g3951(.A1(new_n4336_), .A2(\priority[126] ), .B(\priority[127] ), .ZN(new_n4337_));
  NOR4_X1    g3952(.A1(new_n1943_), .A2(new_n1383_), .A3(new_n2234_), .A4(new_n4337_), .ZN(new_n4338_));
  OAI21_X1   g3953(.A1(new_n2239_), .A2(new_n4338_), .B(new_n2525_), .ZN(new_n4339_));
  AOI21_X1   g3954(.A1(new_n4339_), .A2(new_n2498_), .B(new_n2833_), .ZN(new_n4340_));
  OAI21_X1   g3955(.A1(new_n4340_), .A2(new_n1961_), .B(new_n1964_), .ZN(new_n4341_));
  AOI21_X1   g3956(.A1(new_n4341_), .A2(new_n2449_), .B(new_n2450_), .ZN(new_n4342_));
  OAI21_X1   g3957(.A1(new_n4342_), .A2(new_n1975_), .B(new_n1978_), .ZN(new_n4343_));
  AOI21_X1   g3958(.A1(new_n4343_), .A2(new_n2447_), .B(new_n2448_), .ZN(new_n4344_));
  OAI21_X1   g3959(.A1(new_n4344_), .A2(new_n1989_), .B(new_n1992_), .ZN(new_n4345_));
  AOI21_X1   g3960(.A1(new_n4345_), .A2(new_n2445_), .B(new_n2446_), .ZN(new_n4346_));
  OAI21_X1   g3961(.A1(new_n4346_), .A2(new_n2003_), .B(new_n2006_), .ZN(new_n4347_));
  AOI21_X1   g3962(.A1(new_n4347_), .A2(new_n2443_), .B(new_n2444_), .ZN(new_n4348_));
  OAI21_X1   g3963(.A1(new_n4348_), .A2(new_n2017_), .B(new_n2020_), .ZN(new_n4349_));
  AOI21_X1   g3964(.A1(new_n4349_), .A2(new_n2441_), .B(new_n2442_), .ZN(new_n4350_));
  OAI21_X1   g3965(.A1(new_n4350_), .A2(new_n2031_), .B(new_n2034_), .ZN(new_n4351_));
  NAND2_X1   g3966(.A1(new_n770_), .A2(new_n1376_), .ZN(new_n4352_));
  AOI21_X1   g3967(.A1(new_n4351_), .A2(new_n2439_), .B(new_n4352_), .ZN(\grant[125] ));
  INV_X1     g3968(.I(\req[127] ), .ZN(new_n4354_));
  AOI21_X1   g3969(.A1(new_n4354_), .A2(\priority[127] ), .B(\priority[0] ), .ZN(new_n4355_));
  NOR4_X1    g3970(.A1(new_n2046_), .A2(new_n1567_), .A3(new_n2269_), .A4(new_n4355_), .ZN(new_n4356_));
  OAI21_X1   g3971(.A1(new_n2275_), .A2(new_n4356_), .B(new_n2545_), .ZN(new_n4357_));
  AOI21_X1   g3972(.A1(new_n4357_), .A2(new_n2529_), .B(new_n2851_), .ZN(new_n4358_));
  OAI21_X1   g3973(.A1(new_n4358_), .A2(new_n2062_), .B(new_n2065_), .ZN(new_n4359_));
  AOI21_X1   g3974(.A1(new_n4359_), .A2(new_n2479_), .B(new_n2480_), .ZN(new_n4360_));
  OAI21_X1   g3975(.A1(new_n4360_), .A2(new_n2074_), .B(new_n2077_), .ZN(new_n4361_));
  AOI21_X1   g3976(.A1(new_n4361_), .A2(new_n2477_), .B(new_n2478_), .ZN(new_n4362_));
  OAI21_X1   g3977(.A1(new_n4362_), .A2(new_n2086_), .B(new_n2089_), .ZN(new_n4363_));
  AOI21_X1   g3978(.A1(new_n4363_), .A2(new_n2475_), .B(new_n2476_), .ZN(new_n4364_));
  OAI21_X1   g3979(.A1(new_n4364_), .A2(new_n2098_), .B(new_n2101_), .ZN(new_n4365_));
  AOI21_X1   g3980(.A1(new_n4365_), .A2(new_n2473_), .B(new_n2474_), .ZN(new_n4366_));
  OAI21_X1   g3981(.A1(new_n4366_), .A2(new_n2110_), .B(new_n2113_), .ZN(new_n4367_));
  AOI21_X1   g3982(.A1(new_n4367_), .A2(new_n2471_), .B(new_n2472_), .ZN(new_n4368_));
  OAI21_X1   g3983(.A1(new_n4368_), .A2(new_n2122_), .B(new_n2125_), .ZN(new_n4369_));
  NAND2_X1   g3984(.A1(new_n1123_), .A2(new_n4336_), .ZN(new_n4370_));
  AOI21_X1   g3985(.A1(new_n4369_), .A2(new_n2469_), .B(new_n4370_), .ZN(\grant[126] ));
  OAI21_X1   g3986(.A1(new_n1379_), .A2(\priority[1] ), .B(new_n2130_), .ZN(new_n4372_));
  NOR3_X1    g3987(.A1(new_n4372_), .A2(new_n2137_), .A3(new_n2305_), .ZN(new_n4373_));
  OAI21_X1   g3988(.A1(new_n2311_), .A2(new_n4373_), .B(new_n2565_), .ZN(new_n4374_));
  AOI21_X1   g3989(.A1(new_n4374_), .A2(new_n2549_), .B(new_n2869_), .ZN(new_n4375_));
  OAI21_X1   g3990(.A1(new_n4375_), .A2(new_n2155_), .B(new_n2159_), .ZN(new_n4376_));
  AOI21_X1   g3991(.A1(new_n4376_), .A2(new_n2509_), .B(new_n2510_), .ZN(new_n4377_));
  OAI21_X1   g3992(.A1(new_n4377_), .A2(new_n2169_), .B(new_n2173_), .ZN(new_n4378_));
  AOI21_X1   g3993(.A1(new_n4378_), .A2(new_n2507_), .B(new_n2508_), .ZN(new_n4379_));
  OAI21_X1   g3994(.A1(new_n4379_), .A2(new_n2183_), .B(new_n2187_), .ZN(new_n4380_));
  AOI21_X1   g3995(.A1(new_n4380_), .A2(new_n2505_), .B(new_n2506_), .ZN(new_n4381_));
  OAI21_X1   g3996(.A1(new_n4381_), .A2(new_n2197_), .B(new_n2201_), .ZN(new_n4382_));
  AOI21_X1   g3997(.A1(new_n4382_), .A2(new_n2503_), .B(new_n2504_), .ZN(new_n4383_));
  OAI21_X1   g3998(.A1(new_n4383_), .A2(new_n2211_), .B(new_n2215_), .ZN(new_n4384_));
  AOI21_X1   g3999(.A1(new_n4384_), .A2(new_n2501_), .B(new_n2502_), .ZN(new_n4385_));
  OAI21_X1   g4000(.A1(new_n4385_), .A2(new_n2225_), .B(new_n2229_), .ZN(new_n4386_));
  NAND2_X1   g4001(.A1(new_n1381_), .A2(new_n4354_), .ZN(new_n4387_));
  AOI21_X1   g4002(.A1(new_n4386_), .A2(new_n2499_), .B(new_n4387_), .ZN(\grant[127] ));
  NAND4_X1   g4003(.A1(new_n729_), .A2(new_n1074_), .A3(new_n1083_), .A4(new_n1124_), .ZN(new_n4389_));
  NAND4_X1   g4004(.A1(new_n505_), .A2(new_n561_), .A3(new_n617_), .A4(new_n673_), .ZN(new_n4390_));
  NAND4_X1   g4005(.A1(new_n874_), .A2(new_n883_), .A3(new_n924_), .A4(new_n933_), .ZN(new_n4391_));
  NAND4_X1   g4006(.A1(new_n974_), .A2(new_n983_), .A3(new_n1024_), .A4(new_n1033_), .ZN(new_n4392_));
  NOR4_X1    g4007(.A1(new_n4389_), .A2(new_n4390_), .A3(new_n4391_), .A4(new_n4392_), .ZN(new_n4393_));
  NAND4_X1   g4008(.A1(new_n576_), .A2(new_n585_), .A3(new_n632_), .A4(new_n641_), .ZN(new_n4394_));
  NAND4_X1   g4009(.A1(new_n688_), .A2(new_n697_), .A3(new_n744_), .A4(new_n753_), .ZN(new_n4395_));
  NAND4_X1   g4010(.A1(new_n396_), .A2(new_n408_), .A3(new_n417_), .A4(new_n449_), .ZN(new_n4396_));
  NAND4_X1   g4011(.A1(new_n464_), .A2(new_n473_), .A3(new_n520_), .A4(new_n529_), .ZN(new_n4397_));
  NOR4_X1    g4012(.A1(new_n4394_), .A2(new_n4395_), .A3(new_n4396_), .A4(new_n4397_), .ZN(new_n4398_));
  NAND4_X1   g4013(.A1(new_n1758_), .A2(new_n1154_), .A3(new_n1784_), .A4(new_n1190_), .ZN(new_n4399_));
  NAND4_X1   g4014(.A1(new_n1812_), .A2(new_n1226_), .A3(new_n1840_), .A4(new_n1262_), .ZN(new_n4400_));
  NAND4_X1   g4015(.A1(new_n2192_), .A2(new_n2206_), .A3(new_n2220_), .A4(new_n1566_), .ZN(new_n4401_));
  NAND4_X1   g4016(.A1(new_n1140_), .A2(new_n2150_), .A3(new_n2164_), .A4(new_n2178_), .ZN(new_n4402_));
  NOR4_X1    g4017(.A1(new_n4399_), .A2(new_n4400_), .A3(new_n4401_), .A4(new_n4402_), .ZN(new_n4403_));
  NAND4_X1   g4018(.A1(new_n862_), .A2(new_n912_), .A3(new_n962_), .A4(new_n1012_), .ZN(new_n4404_));
  NAND4_X1   g4019(.A1(new_n788_), .A2(new_n812_), .A3(new_n824_), .A4(new_n833_), .ZN(new_n4405_));
  NAND4_X1   g4020(.A1(new_n1868_), .A2(new_n1298_), .A3(new_n1896_), .A4(new_n1334_), .ZN(new_n4406_));
  NAND4_X1   g4021(.A1(new_n1062_), .A2(new_n1112_), .A3(new_n1924_), .A4(new_n1370_), .ZN(new_n4407_));
  NOR4_X1    g4022(.A1(new_n4404_), .A2(new_n4405_), .A3(new_n4406_), .A4(new_n4407_), .ZN(new_n4408_));
  AND4_X2    g4023(.A1(new_n4393_), .A2(new_n4398_), .A3(new_n4403_), .A4(new_n4408_), .Z(anyGrant));
endmodule


