// Benchmark "priority" written by ABC on Thu Sep 14 22:44:23 2023

module priority ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] ,
    \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] ;
  output \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F;
  wire new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1319_, new_n1320_, new_n1321_, new_n1323_, new_n1325_,
    new_n1326_, new_n1327_;
  INV_X1     g0000(.I(\A[9] ), .ZN(new_n137_));
  INV_X1     g0001(.I(\A[11] ), .ZN(new_n138_));
  INV_X1     g0002(.I(\A[13] ), .ZN(new_n139_));
  INV_X1     g0003(.I(\A[19] ), .ZN(new_n140_));
  INV_X1     g0004(.I(\A[25] ), .ZN(new_n141_));
  INV_X1     g0005(.I(\A[31] ), .ZN(new_n142_));
  INV_X1     g0006(.I(\A[37] ), .ZN(new_n143_));
  INV_X1     g0007(.I(\A[43] ), .ZN(new_n144_));
  INV_X1     g0008(.I(\A[49] ), .ZN(new_n145_));
  INV_X1     g0009(.I(\A[55] ), .ZN(new_n146_));
  INV_X1     g0010(.I(\A[61] ), .ZN(new_n147_));
  INV_X1     g0011(.I(\A[67] ), .ZN(new_n148_));
  INV_X1     g0012(.I(\A[73] ), .ZN(new_n149_));
  INV_X1     g0013(.I(\A[79] ), .ZN(new_n150_));
  INV_X1     g0014(.I(\A[87] ), .ZN(new_n151_));
  INV_X1     g0015(.I(\A[89] ), .ZN(new_n152_));
  INV_X1     g0016(.I(\A[95] ), .ZN(new_n153_));
  INV_X1     g0017(.I(\A[99] ), .ZN(new_n154_));
  INV_X1     g0018(.I(\A[101] ), .ZN(new_n155_));
  INV_X1     g0019(.I(\A[105] ), .ZN(new_n156_));
  INV_X1     g0020(.I(\A[113] ), .ZN(new_n157_));
  INV_X1     g0021(.I(\A[115] ), .ZN(new_n158_));
  INV_X1     g0022(.I(\A[117] ), .ZN(new_n159_));
  INV_X1     g0023(.I(\A[121] ), .ZN(new_n160_));
  INV_X1     g0024(.I(\A[123] ), .ZN(new_n161_));
  INV_X1     g0025(.I(\A[126] ), .ZN(new_n162_));
  AOI21_X1   g0026(.A1(new_n162_), .A2(\A[125] ), .B(\A[127] ), .ZN(new_n163_));
  NAND2_X1   g0027(.A1(new_n163_), .A2(new_n161_), .ZN(new_n164_));
  AND2_X2    g0028(.A1(\A[126] ), .A2(\A[127] ), .Z(new_n165_));
  OAI21_X1   g0029(.A1(new_n165_), .A2(\A[124] ), .B(\A[125] ), .ZN(new_n166_));
  OAI21_X1   g0030(.A1(new_n161_), .A2(new_n166_), .B(new_n164_), .ZN(new_n167_));
  NAND2_X1   g0031(.A1(new_n167_), .A2(new_n160_), .ZN(new_n168_));
  INV_X1     g0032(.I(\A[125] ), .ZN(new_n169_));
  INV_X1     g0033(.I(\A[127] ), .ZN(new_n170_));
  OAI21_X1   g0034(.A1(new_n169_), .A2(\A[126] ), .B(new_n170_), .ZN(new_n171_));
  AOI21_X1   g0035(.A1(\A[126] ), .A2(\A[127] ), .B(\A[124] ), .ZN(new_n172_));
  NAND2_X1   g0036(.A1(\A[122] ), .A2(\A[123] ), .ZN(new_n173_));
  NOR4_X1    g0037(.A1(new_n171_), .A2(new_n169_), .A3(new_n172_), .A4(new_n173_), .ZN(new_n174_));
  NOR2_X1    g0038(.A1(new_n172_), .A2(new_n169_), .ZN(new_n175_));
  NOR3_X1    g0039(.A1(new_n175_), .A2(new_n163_), .A3(new_n173_), .ZN(new_n176_));
  OAI21_X1   g0040(.A1(new_n176_), .A2(new_n174_), .B(\A[121] ), .ZN(new_n177_));
  AOI21_X1   g0041(.A1(new_n168_), .A2(new_n177_), .B(\A[119] ), .ZN(new_n178_));
  INV_X1     g0042(.I(new_n178_), .ZN(new_n179_));
  NOR2_X1    g0043(.A1(new_n171_), .A2(\A[123] ), .ZN(new_n180_));
  NOR3_X1    g0044(.A1(new_n172_), .A2(new_n161_), .A3(new_n169_), .ZN(new_n181_));
  INV_X1     g0045(.I(\A[120] ), .ZN(new_n182_));
  NOR2_X1    g0046(.A1(new_n182_), .A2(new_n160_), .ZN(new_n183_));
  INV_X1     g0047(.I(new_n183_), .ZN(new_n184_));
  NOR3_X1    g0048(.A1(new_n180_), .A2(new_n181_), .A3(new_n184_), .ZN(new_n185_));
  OAI21_X1   g0049(.A1(new_n176_), .A2(new_n174_), .B(new_n183_), .ZN(new_n186_));
  NOR2_X1    g0050(.A1(new_n186_), .A2(new_n185_), .ZN(new_n187_));
  NOR4_X1    g0051(.A1(new_n167_), .A2(new_n174_), .A3(new_n176_), .A4(new_n184_), .ZN(new_n188_));
  OAI21_X1   g0052(.A1(new_n187_), .A2(new_n188_), .B(\A[119] ), .ZN(new_n189_));
  NAND2_X1   g0053(.A1(new_n179_), .A2(new_n189_), .ZN(new_n190_));
  NAND2_X1   g0054(.A1(new_n190_), .A2(new_n159_), .ZN(new_n191_));
  NOR2_X1    g0055(.A1(new_n180_), .A2(new_n181_), .ZN(new_n192_));
  NOR2_X1    g0056(.A1(new_n192_), .A2(\A[121] ), .ZN(new_n193_));
  INV_X1     g0057(.I(new_n177_), .ZN(new_n194_));
  NAND2_X1   g0058(.A1(\A[118] ), .A2(\A[119] ), .ZN(new_n195_));
  NOR3_X1    g0059(.A1(new_n194_), .A2(new_n193_), .A3(new_n195_), .ZN(new_n196_));
  INV_X1     g0060(.I(new_n195_), .ZN(new_n197_));
  OAI21_X1   g0061(.A1(new_n187_), .A2(new_n188_), .B(new_n197_), .ZN(new_n198_));
  NOR2_X1    g0062(.A1(new_n198_), .A2(new_n196_), .ZN(new_n199_));
  NAND2_X1   g0063(.A1(new_n168_), .A2(new_n177_), .ZN(new_n200_));
  NOR4_X1    g0064(.A1(new_n200_), .A2(new_n187_), .A3(new_n188_), .A4(new_n195_), .ZN(new_n201_));
  OAI21_X1   g0065(.A1(new_n199_), .A2(new_n201_), .B(\A[117] ), .ZN(new_n202_));
  AOI21_X1   g0066(.A1(new_n202_), .A2(new_n191_), .B(\A[115] ), .ZN(new_n203_));
  INV_X1     g0067(.I(new_n203_), .ZN(new_n204_));
  INV_X1     g0068(.I(new_n173_), .ZN(new_n205_));
  NAND3_X1   g0069(.A1(new_n175_), .A2(new_n163_), .A3(new_n205_), .ZN(new_n206_));
  NAND3_X1   g0070(.A1(new_n166_), .A2(new_n171_), .A3(new_n205_), .ZN(new_n207_));
  NAND2_X1   g0071(.A1(new_n207_), .A2(new_n206_), .ZN(new_n208_));
  NAND3_X1   g0072(.A1(new_n208_), .A2(new_n167_), .A3(new_n183_), .ZN(new_n209_));
  NAND2_X1   g0073(.A1(new_n186_), .A2(new_n185_), .ZN(new_n210_));
  NAND2_X1   g0074(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  AOI21_X1   g0075(.A1(new_n211_), .A2(\A[119] ), .B(new_n178_), .ZN(new_n212_));
  NOR2_X1    g0076(.A1(new_n199_), .A2(new_n201_), .ZN(new_n213_));
  NAND2_X1   g0077(.A1(\A[116] ), .A2(\A[117] ), .ZN(new_n214_));
  NOR3_X1    g0078(.A1(new_n213_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n215_));
  NOR4_X1    g0079(.A1(new_n190_), .A2(new_n199_), .A3(new_n201_), .A4(new_n214_), .ZN(new_n216_));
  NOR2_X1    g0080(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1   g0081(.A1(new_n158_), .A2(new_n217_), .B(new_n204_), .ZN(new_n218_));
  NAND2_X1   g0082(.A1(new_n218_), .A2(new_n157_), .ZN(new_n219_));
  NOR2_X1    g0083(.A1(new_n212_), .A2(\A[117] ), .ZN(new_n220_));
  NAND3_X1   g0084(.A1(new_n211_), .A2(new_n200_), .A3(new_n197_), .ZN(new_n221_));
  NAND2_X1   g0085(.A1(new_n198_), .A2(new_n196_), .ZN(new_n222_));
  NAND2_X1   g0086(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  AOI21_X1   g0087(.A1(\A[117] ), .A2(new_n223_), .B(new_n220_), .ZN(new_n224_));
  NAND2_X1   g0088(.A1(\A[114] ), .A2(\A[115] ), .ZN(new_n225_));
  NOR3_X1    g0089(.A1(new_n217_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1   g0090(.A1(new_n202_), .A2(new_n191_), .ZN(new_n227_));
  INV_X1     g0091(.I(new_n214_), .ZN(new_n228_));
  NAND3_X1   g0092(.A1(new_n223_), .A2(new_n190_), .A3(new_n228_), .ZN(new_n229_));
  NAND4_X1   g0093(.A1(new_n212_), .A2(new_n221_), .A3(new_n222_), .A4(new_n228_), .ZN(new_n230_));
  NAND2_X1   g0094(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR3_X1    g0095(.A1(new_n231_), .A2(new_n227_), .A3(new_n225_), .ZN(new_n232_));
  OAI21_X1   g0096(.A1(new_n232_), .A2(new_n226_), .B(\A[113] ), .ZN(new_n233_));
  AOI21_X1   g0097(.A1(new_n233_), .A2(new_n219_), .B(\A[111] ), .ZN(new_n234_));
  INV_X1     g0098(.I(new_n225_), .ZN(new_n235_));
  NAND3_X1   g0099(.A1(new_n231_), .A2(new_n227_), .A3(new_n235_), .ZN(new_n236_));
  NAND4_X1   g0100(.A1(new_n224_), .A2(new_n229_), .A3(new_n230_), .A4(new_n235_), .ZN(new_n237_));
  NAND2_X1   g0101(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1   g0102(.A1(\A[112] ), .A2(\A[113] ), .ZN(new_n239_));
  INV_X1     g0103(.I(new_n239_), .ZN(new_n240_));
  NAND3_X1   g0104(.A1(new_n238_), .A2(new_n218_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1   g0105(.A1(new_n231_), .A2(\A[115] ), .B(new_n203_), .ZN(new_n242_));
  NAND4_X1   g0106(.A1(new_n242_), .A2(new_n236_), .A3(new_n237_), .A4(new_n240_), .ZN(new_n243_));
  NAND2_X1   g0107(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1   g0108(.A1(new_n244_), .A2(\A[111] ), .B(new_n234_), .ZN(new_n245_));
  OR2_X2     g0109(.A1(new_n245_), .A2(\A[109] ), .Z(new_n246_));
  NOR2_X1    g0110(.A1(new_n242_), .A2(\A[113] ), .ZN(new_n247_));
  AOI21_X1   g0111(.A1(\A[113] ), .A2(new_n238_), .B(new_n247_), .ZN(new_n248_));
  NOR2_X1    g0112(.A1(new_n232_), .A2(new_n226_), .ZN(new_n249_));
  NOR3_X1    g0113(.A1(new_n249_), .A2(new_n242_), .A3(new_n239_), .ZN(new_n250_));
  INV_X1     g0114(.I(new_n243_), .ZN(new_n251_));
  NOR2_X1    g0115(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1   g0116(.A1(\A[110] ), .A2(\A[111] ), .ZN(new_n253_));
  NOR3_X1    g0117(.A1(new_n252_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1   g0118(.A1(new_n233_), .A2(new_n219_), .ZN(new_n255_));
  NOR3_X1    g0119(.A1(new_n244_), .A2(new_n255_), .A3(new_n253_), .ZN(new_n256_));
  OAI21_X1   g0120(.A1(new_n254_), .A2(new_n256_), .B(\A[109] ), .ZN(new_n257_));
  AOI21_X1   g0121(.A1(new_n246_), .A2(new_n257_), .B(\A[107] ), .ZN(new_n258_));
  INV_X1     g0122(.I(new_n258_), .ZN(new_n259_));
  OAI21_X1   g0123(.A1(new_n250_), .A2(new_n251_), .B(\A[111] ), .ZN(new_n260_));
  OAI21_X1   g0124(.A1(\A[111] ), .A2(new_n248_), .B(new_n260_), .ZN(new_n261_));
  INV_X1     g0125(.I(new_n253_), .ZN(new_n262_));
  NAND3_X1   g0126(.A1(new_n244_), .A2(new_n255_), .A3(new_n262_), .ZN(new_n263_));
  NAND4_X1   g0127(.A1(new_n248_), .A2(new_n241_), .A3(new_n243_), .A4(new_n262_), .ZN(new_n264_));
  NAND2_X1   g0128(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1   g0129(.A1(\A[108] ), .A2(\A[109] ), .ZN(new_n266_));
  INV_X1     g0130(.I(new_n266_), .ZN(new_n267_));
  NAND3_X1   g0131(.A1(new_n265_), .A2(new_n261_), .A3(new_n267_), .ZN(new_n268_));
  NAND4_X1   g0132(.A1(new_n245_), .A2(new_n263_), .A3(new_n264_), .A4(new_n267_), .ZN(new_n269_));
  NAND2_X1   g0133(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1   g0134(.A1(new_n270_), .A2(\A[107] ), .ZN(new_n271_));
  NAND2_X1   g0135(.A1(new_n271_), .A2(new_n259_), .ZN(new_n272_));
  NAND2_X1   g0136(.A1(new_n272_), .A2(new_n156_), .ZN(new_n273_));
  NAND2_X1   g0137(.A1(new_n246_), .A2(new_n257_), .ZN(new_n274_));
  NAND2_X1   g0138(.A1(\A[106] ), .A2(\A[107] ), .ZN(new_n275_));
  INV_X1     g0139(.I(new_n275_), .ZN(new_n276_));
  NAND3_X1   g0140(.A1(new_n270_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  NOR2_X1    g0141(.A1(new_n245_), .A2(\A[109] ), .ZN(new_n278_));
  AOI21_X1   g0142(.A1(\A[109] ), .A2(new_n265_), .B(new_n278_), .ZN(new_n279_));
  NAND4_X1   g0143(.A1(new_n279_), .A2(new_n268_), .A3(new_n269_), .A4(new_n276_), .ZN(new_n280_));
  NAND2_X1   g0144(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1   g0145(.A1(new_n281_), .A2(\A[105] ), .ZN(new_n282_));
  AOI21_X1   g0146(.A1(new_n282_), .A2(new_n273_), .B(\A[103] ), .ZN(new_n283_));
  INV_X1     g0147(.I(\A[103] ), .ZN(new_n284_));
  NAND2_X1   g0148(.A1(\A[104] ), .A2(\A[105] ), .ZN(new_n285_));
  INV_X1     g0149(.I(new_n285_), .ZN(new_n286_));
  NAND3_X1   g0150(.A1(new_n281_), .A2(new_n272_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1   g0151(.A1(new_n270_), .A2(\A[107] ), .B(new_n258_), .ZN(new_n288_));
  NAND4_X1   g0152(.A1(new_n288_), .A2(new_n277_), .A3(new_n280_), .A4(new_n286_), .ZN(new_n289_));
  AOI21_X1   g0153(.A1(new_n287_), .A2(new_n289_), .B(new_n284_), .ZN(new_n290_));
  OAI21_X1   g0154(.A1(new_n290_), .A2(new_n283_), .B(new_n155_), .ZN(new_n291_));
  NAND2_X1   g0155(.A1(new_n282_), .A2(new_n273_), .ZN(new_n292_));
  NAND2_X1   g0156(.A1(new_n287_), .A2(new_n289_), .ZN(new_n293_));
  INV_X1     g0157(.I(\A[102] ), .ZN(new_n294_));
  NOR2_X1    g0158(.A1(new_n294_), .A2(new_n284_), .ZN(new_n295_));
  NAND3_X1   g0159(.A1(new_n293_), .A2(new_n292_), .A3(new_n295_), .ZN(new_n296_));
  NOR2_X1    g0160(.A1(new_n288_), .A2(\A[105] ), .ZN(new_n297_));
  AOI21_X1   g0161(.A1(\A[105] ), .A2(new_n281_), .B(new_n297_), .ZN(new_n298_));
  NAND4_X1   g0162(.A1(new_n298_), .A2(new_n287_), .A3(new_n289_), .A4(new_n295_), .ZN(new_n299_));
  NAND2_X1   g0163(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1   g0164(.A1(new_n300_), .A2(\A[101] ), .ZN(new_n301_));
  NAND2_X1   g0165(.A1(new_n301_), .A2(new_n291_), .ZN(new_n302_));
  NAND2_X1   g0166(.A1(new_n302_), .A2(new_n154_), .ZN(new_n303_));
  OR2_X2     g0167(.A1(new_n290_), .A2(new_n283_), .Z(new_n304_));
  AND2_X2    g0168(.A1(\A[100] ), .A2(\A[101] ), .Z(new_n305_));
  NAND3_X1   g0169(.A1(new_n300_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NOR2_X1    g0170(.A1(new_n290_), .A2(new_n283_), .ZN(new_n307_));
  NAND4_X1   g0171(.A1(new_n307_), .A2(new_n296_), .A3(new_n299_), .A4(new_n305_), .ZN(new_n308_));
  NAND2_X1   g0172(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1   g0173(.A1(new_n309_), .A2(\A[99] ), .ZN(new_n310_));
  AOI21_X1   g0174(.A1(new_n310_), .A2(new_n303_), .B(\A[97] ), .ZN(new_n311_));
  INV_X1     g0175(.I(\A[97] ), .ZN(new_n312_));
  NAND2_X1   g0176(.A1(\A[98] ), .A2(\A[99] ), .ZN(new_n313_));
  INV_X1     g0177(.I(new_n313_), .ZN(new_n314_));
  NAND3_X1   g0178(.A1(new_n309_), .A2(new_n302_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1     g0179(.I(new_n291_), .ZN(new_n316_));
  AOI21_X1   g0180(.A1(\A[101] ), .A2(new_n300_), .B(new_n316_), .ZN(new_n317_));
  NAND4_X1   g0181(.A1(new_n317_), .A2(new_n306_), .A3(new_n308_), .A4(new_n314_), .ZN(new_n318_));
  AOI21_X1   g0182(.A1(new_n315_), .A2(new_n318_), .B(new_n312_), .ZN(new_n319_));
  OAI21_X1   g0183(.A1(new_n319_), .A2(new_n311_), .B(new_n153_), .ZN(new_n320_));
  INV_X1     g0184(.I(new_n320_), .ZN(new_n321_));
  NAND2_X1   g0185(.A1(new_n310_), .A2(new_n303_), .ZN(new_n322_));
  NAND2_X1   g0186(.A1(new_n315_), .A2(new_n318_), .ZN(new_n323_));
  NAND2_X1   g0187(.A1(\A[96] ), .A2(\A[97] ), .ZN(new_n324_));
  INV_X1     g0188(.I(new_n324_), .ZN(new_n325_));
  NAND3_X1   g0189(.A1(new_n323_), .A2(new_n322_), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1   g0190(.A1(new_n301_), .A2(new_n291_), .B(\A[99] ), .ZN(new_n327_));
  AOI21_X1   g0191(.A1(\A[99] ), .A2(new_n309_), .B(new_n327_), .ZN(new_n328_));
  NAND4_X1   g0192(.A1(new_n328_), .A2(new_n315_), .A3(new_n318_), .A4(new_n325_), .ZN(new_n329_));
  NAND2_X1   g0193(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1   g0194(.A1(\A[95] ), .A2(new_n330_), .B(new_n321_), .ZN(new_n331_));
  NOR2_X1    g0195(.A1(new_n331_), .A2(\A[93] ), .ZN(new_n332_));
  INV_X1     g0196(.I(\A[93] ), .ZN(new_n333_));
  OR2_X2     g0197(.A1(new_n319_), .A2(new_n311_), .Z(new_n334_));
  NAND2_X1   g0198(.A1(\A[94] ), .A2(\A[95] ), .ZN(new_n335_));
  INV_X1     g0199(.I(new_n335_), .ZN(new_n336_));
  NAND3_X1   g0200(.A1(new_n330_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  NOR2_X1    g0201(.A1(new_n319_), .A2(new_n311_), .ZN(new_n338_));
  NAND4_X1   g0202(.A1(new_n338_), .A2(new_n326_), .A3(new_n329_), .A4(new_n336_), .ZN(new_n339_));
  AOI21_X1   g0203(.A1(new_n337_), .A2(new_n339_), .B(new_n333_), .ZN(new_n340_));
  NOR2_X1    g0204(.A1(new_n332_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1    g0205(.A1(new_n341_), .A2(\A[91] ), .ZN(new_n342_));
  INV_X1     g0206(.I(\A[91] ), .ZN(new_n343_));
  NAND2_X1   g0207(.A1(new_n330_), .A2(\A[95] ), .ZN(new_n344_));
  NAND2_X1   g0208(.A1(new_n344_), .A2(new_n320_), .ZN(new_n345_));
  NAND2_X1   g0209(.A1(new_n337_), .A2(new_n339_), .ZN(new_n346_));
  NAND2_X1   g0210(.A1(\A[92] ), .A2(\A[93] ), .ZN(new_n347_));
  INV_X1     g0211(.I(new_n347_), .ZN(new_n348_));
  NAND3_X1   g0212(.A1(new_n346_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n349_));
  NAND4_X1   g0213(.A1(new_n331_), .A2(new_n337_), .A3(new_n339_), .A4(new_n348_), .ZN(new_n350_));
  AOI21_X1   g0214(.A1(new_n349_), .A2(new_n350_), .B(new_n343_), .ZN(new_n351_));
  OAI21_X1   g0215(.A1(new_n342_), .A2(new_n351_), .B(new_n152_), .ZN(new_n352_));
  NAND2_X1   g0216(.A1(new_n345_), .A2(new_n333_), .ZN(new_n353_));
  NAND2_X1   g0217(.A1(new_n346_), .A2(\A[93] ), .ZN(new_n354_));
  NAND2_X1   g0218(.A1(new_n354_), .A2(new_n353_), .ZN(new_n355_));
  NAND2_X1   g0219(.A1(new_n349_), .A2(new_n350_), .ZN(new_n356_));
  NAND2_X1   g0220(.A1(\A[90] ), .A2(\A[91] ), .ZN(new_n357_));
  INV_X1     g0221(.I(new_n357_), .ZN(new_n358_));
  NAND3_X1   g0222(.A1(new_n356_), .A2(new_n355_), .A3(new_n358_), .ZN(new_n359_));
  NAND4_X1   g0223(.A1(new_n341_), .A2(new_n349_), .A3(new_n350_), .A4(new_n358_), .ZN(new_n360_));
  NAND2_X1   g0224(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1   g0225(.A1(new_n361_), .A2(\A[89] ), .ZN(new_n362_));
  NAND2_X1   g0226(.A1(new_n362_), .A2(new_n352_), .ZN(new_n363_));
  NAND2_X1   g0227(.A1(new_n363_), .A2(new_n151_), .ZN(new_n364_));
  NAND2_X1   g0228(.A1(new_n355_), .A2(new_n343_), .ZN(new_n365_));
  NAND2_X1   g0229(.A1(new_n356_), .A2(\A[91] ), .ZN(new_n366_));
  NAND2_X1   g0230(.A1(new_n366_), .A2(new_n365_), .ZN(new_n367_));
  NAND2_X1   g0231(.A1(\A[88] ), .A2(\A[89] ), .ZN(new_n368_));
  INV_X1     g0232(.I(new_n368_), .ZN(new_n369_));
  NAND3_X1   g0233(.A1(new_n361_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  NOR2_X1    g0234(.A1(new_n342_), .A2(new_n351_), .ZN(new_n371_));
  NAND4_X1   g0235(.A1(new_n371_), .A2(new_n359_), .A3(new_n360_), .A4(new_n369_), .ZN(new_n372_));
  NAND2_X1   g0236(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1   g0237(.A1(new_n373_), .A2(\A[87] ), .ZN(new_n374_));
  AOI21_X1   g0238(.A1(new_n374_), .A2(new_n364_), .B(\A[85] ), .ZN(new_n375_));
  INV_X1     g0239(.I(\A[85] ), .ZN(new_n376_));
  NAND2_X1   g0240(.A1(\A[86] ), .A2(\A[87] ), .ZN(new_n377_));
  INV_X1     g0241(.I(new_n377_), .ZN(new_n378_));
  NAND3_X1   g0242(.A1(new_n373_), .A2(new_n363_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1     g0243(.I(new_n352_), .ZN(new_n380_));
  AOI21_X1   g0244(.A1(new_n359_), .A2(new_n360_), .B(new_n152_), .ZN(new_n381_));
  NOR2_X1    g0245(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1   g0246(.A1(new_n382_), .A2(new_n370_), .A3(new_n372_), .A4(new_n378_), .ZN(new_n383_));
  AOI21_X1   g0247(.A1(new_n379_), .A2(new_n383_), .B(new_n376_), .ZN(new_n384_));
  NOR2_X1    g0248(.A1(new_n384_), .A2(new_n375_), .ZN(new_n385_));
  NOR2_X1    g0249(.A1(new_n385_), .A2(\A[83] ), .ZN(new_n386_));
  INV_X1     g0250(.I(\A[83] ), .ZN(new_n387_));
  NAND2_X1   g0251(.A1(new_n374_), .A2(new_n364_), .ZN(new_n388_));
  NAND2_X1   g0252(.A1(new_n379_), .A2(new_n383_), .ZN(new_n389_));
  NAND2_X1   g0253(.A1(\A[84] ), .A2(\A[85] ), .ZN(new_n390_));
  INV_X1     g0254(.I(new_n390_), .ZN(new_n391_));
  NAND3_X1   g0255(.A1(new_n389_), .A2(new_n388_), .A3(new_n391_), .ZN(new_n392_));
  NOR2_X1    g0256(.A1(new_n382_), .A2(\A[87] ), .ZN(new_n393_));
  AOI21_X1   g0257(.A1(new_n370_), .A2(new_n372_), .B(new_n151_), .ZN(new_n394_));
  NOR2_X1    g0258(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND4_X1   g0259(.A1(new_n395_), .A2(new_n379_), .A3(new_n383_), .A4(new_n391_), .ZN(new_n396_));
  AOI21_X1   g0260(.A1(new_n392_), .A2(new_n396_), .B(new_n387_), .ZN(new_n397_));
  NOR2_X1    g0261(.A1(new_n397_), .A2(new_n386_), .ZN(new_n398_));
  NOR2_X1    g0262(.A1(new_n398_), .A2(\A[81] ), .ZN(new_n399_));
  INV_X1     g0263(.I(\A[81] ), .ZN(new_n400_));
  OR2_X2     g0264(.A1(new_n384_), .A2(new_n375_), .Z(new_n401_));
  NAND2_X1   g0265(.A1(new_n392_), .A2(new_n396_), .ZN(new_n402_));
  NAND2_X1   g0266(.A1(\A[82] ), .A2(\A[83] ), .ZN(new_n403_));
  INV_X1     g0267(.I(new_n403_), .ZN(new_n404_));
  NAND3_X1   g0268(.A1(new_n402_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n405_));
  NAND4_X1   g0269(.A1(new_n385_), .A2(new_n392_), .A3(new_n396_), .A4(new_n404_), .ZN(new_n406_));
  AOI21_X1   g0270(.A1(new_n405_), .A2(new_n406_), .B(new_n400_), .ZN(new_n407_));
  OAI21_X1   g0271(.A1(new_n407_), .A2(new_n399_), .B(new_n150_), .ZN(new_n408_));
  INV_X1     g0272(.I(new_n408_), .ZN(new_n409_));
  OR2_X2     g0273(.A1(new_n397_), .A2(new_n386_), .Z(new_n410_));
  NAND2_X1   g0274(.A1(new_n405_), .A2(new_n406_), .ZN(new_n411_));
  NAND2_X1   g0275(.A1(\A[80] ), .A2(\A[81] ), .ZN(new_n412_));
  INV_X1     g0276(.I(new_n412_), .ZN(new_n413_));
  NAND3_X1   g0277(.A1(new_n411_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n414_));
  NAND4_X1   g0278(.A1(new_n398_), .A2(new_n405_), .A3(new_n406_), .A4(new_n413_), .ZN(new_n415_));
  AOI21_X1   g0279(.A1(new_n414_), .A2(new_n415_), .B(new_n150_), .ZN(new_n416_));
  NOR2_X1    g0280(.A1(new_n416_), .A2(new_n409_), .ZN(new_n417_));
  NOR2_X1    g0281(.A1(new_n417_), .A2(\A[77] ), .ZN(new_n418_));
  INV_X1     g0282(.I(\A[77] ), .ZN(new_n419_));
  OR2_X2     g0283(.A1(new_n407_), .A2(new_n399_), .Z(new_n420_));
  NAND2_X1   g0284(.A1(new_n414_), .A2(new_n415_), .ZN(new_n421_));
  AND2_X2    g0285(.A1(\A[78] ), .A2(\A[79] ), .Z(new_n422_));
  NAND3_X1   g0286(.A1(new_n421_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  NOR2_X1    g0287(.A1(new_n407_), .A2(new_n399_), .ZN(new_n424_));
  NAND4_X1   g0288(.A1(new_n424_), .A2(new_n414_), .A3(new_n415_), .A4(new_n422_), .ZN(new_n425_));
  AOI21_X1   g0289(.A1(new_n423_), .A2(new_n425_), .B(new_n419_), .ZN(new_n426_));
  NOR2_X1    g0290(.A1(new_n418_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1    g0291(.A1(new_n427_), .A2(\A[75] ), .ZN(new_n428_));
  INV_X1     g0292(.I(\A[75] ), .ZN(new_n429_));
  NAND2_X1   g0293(.A1(new_n421_), .A2(\A[79] ), .ZN(new_n430_));
  NAND2_X1   g0294(.A1(new_n430_), .A2(new_n408_), .ZN(new_n431_));
  NAND2_X1   g0295(.A1(new_n423_), .A2(new_n425_), .ZN(new_n432_));
  AND2_X2    g0296(.A1(\A[76] ), .A2(\A[77] ), .Z(new_n433_));
  NAND3_X1   g0297(.A1(new_n432_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  NAND4_X1   g0298(.A1(new_n417_), .A2(new_n423_), .A3(new_n425_), .A4(new_n433_), .ZN(new_n435_));
  AOI21_X1   g0299(.A1(new_n434_), .A2(new_n435_), .B(new_n429_), .ZN(new_n436_));
  OAI21_X1   g0300(.A1(new_n428_), .A2(new_n436_), .B(new_n149_), .ZN(new_n437_));
  INV_X1     g0301(.I(new_n437_), .ZN(new_n438_));
  NAND2_X1   g0302(.A1(new_n431_), .A2(new_n419_), .ZN(new_n439_));
  NAND2_X1   g0303(.A1(new_n432_), .A2(\A[77] ), .ZN(new_n440_));
  NAND2_X1   g0304(.A1(new_n440_), .A2(new_n439_), .ZN(new_n441_));
  NAND2_X1   g0305(.A1(new_n434_), .A2(new_n435_), .ZN(new_n442_));
  NAND2_X1   g0306(.A1(\A[74] ), .A2(\A[75] ), .ZN(new_n443_));
  INV_X1     g0307(.I(new_n443_), .ZN(new_n444_));
  NAND3_X1   g0308(.A1(new_n442_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  NAND4_X1   g0309(.A1(new_n427_), .A2(new_n434_), .A3(new_n435_), .A4(new_n444_), .ZN(new_n446_));
  AOI21_X1   g0310(.A1(new_n445_), .A2(new_n446_), .B(new_n149_), .ZN(new_n447_));
  NOR2_X1    g0311(.A1(new_n438_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1    g0312(.A1(new_n448_), .A2(\A[71] ), .ZN(new_n449_));
  INV_X1     g0313(.I(\A[71] ), .ZN(new_n450_));
  NAND2_X1   g0314(.A1(new_n441_), .A2(new_n429_), .ZN(new_n451_));
  NAND2_X1   g0315(.A1(new_n442_), .A2(\A[75] ), .ZN(new_n452_));
  NAND2_X1   g0316(.A1(new_n452_), .A2(new_n451_), .ZN(new_n453_));
  NAND2_X1   g0317(.A1(new_n445_), .A2(new_n446_), .ZN(new_n454_));
  NAND2_X1   g0318(.A1(\A[72] ), .A2(\A[73] ), .ZN(new_n455_));
  INV_X1     g0319(.I(new_n455_), .ZN(new_n456_));
  NAND3_X1   g0320(.A1(new_n454_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  NOR2_X1    g0321(.A1(new_n428_), .A2(new_n436_), .ZN(new_n458_));
  NAND4_X1   g0322(.A1(new_n458_), .A2(new_n445_), .A3(new_n446_), .A4(new_n456_), .ZN(new_n459_));
  AOI21_X1   g0323(.A1(new_n457_), .A2(new_n459_), .B(new_n450_), .ZN(new_n460_));
  NOR2_X1    g0324(.A1(new_n449_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1    g0325(.A1(new_n461_), .A2(\A[69] ), .ZN(new_n462_));
  INV_X1     g0326(.I(\A[69] ), .ZN(new_n463_));
  NAND2_X1   g0327(.A1(new_n454_), .A2(\A[73] ), .ZN(new_n464_));
  NAND2_X1   g0328(.A1(new_n464_), .A2(new_n437_), .ZN(new_n465_));
  NAND2_X1   g0329(.A1(new_n457_), .A2(new_n459_), .ZN(new_n466_));
  NAND2_X1   g0330(.A1(\A[70] ), .A2(\A[71] ), .ZN(new_n467_));
  INV_X1     g0331(.I(new_n467_), .ZN(new_n468_));
  NAND3_X1   g0332(.A1(new_n466_), .A2(new_n465_), .A3(new_n468_), .ZN(new_n469_));
  NAND4_X1   g0333(.A1(new_n448_), .A2(new_n457_), .A3(new_n459_), .A4(new_n468_), .ZN(new_n470_));
  AOI21_X1   g0334(.A1(new_n469_), .A2(new_n470_), .B(new_n463_), .ZN(new_n471_));
  OAI21_X1   g0335(.A1(new_n462_), .A2(new_n471_), .B(new_n148_), .ZN(new_n472_));
  INV_X1     g0336(.I(new_n472_), .ZN(new_n473_));
  NAND2_X1   g0337(.A1(new_n465_), .A2(new_n450_), .ZN(new_n474_));
  NAND2_X1   g0338(.A1(new_n466_), .A2(\A[71] ), .ZN(new_n475_));
  NAND2_X1   g0339(.A1(new_n475_), .A2(new_n474_), .ZN(new_n476_));
  NAND2_X1   g0340(.A1(new_n469_), .A2(new_n470_), .ZN(new_n477_));
  NAND2_X1   g0341(.A1(\A[68] ), .A2(\A[69] ), .ZN(new_n478_));
  INV_X1     g0342(.I(new_n478_), .ZN(new_n479_));
  NAND3_X1   g0343(.A1(new_n477_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  NAND4_X1   g0344(.A1(new_n461_), .A2(new_n469_), .A3(new_n470_), .A4(new_n479_), .ZN(new_n481_));
  AOI21_X1   g0345(.A1(new_n480_), .A2(new_n481_), .B(new_n148_), .ZN(new_n482_));
  NOR2_X1    g0346(.A1(new_n473_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1    g0347(.A1(new_n483_), .A2(\A[65] ), .ZN(new_n484_));
  INV_X1     g0348(.I(\A[65] ), .ZN(new_n485_));
  NAND2_X1   g0349(.A1(new_n476_), .A2(new_n463_), .ZN(new_n486_));
  NAND2_X1   g0350(.A1(new_n477_), .A2(\A[69] ), .ZN(new_n487_));
  NAND2_X1   g0351(.A1(new_n487_), .A2(new_n486_), .ZN(new_n488_));
  NAND2_X1   g0352(.A1(new_n480_), .A2(new_n481_), .ZN(new_n489_));
  NAND2_X1   g0353(.A1(\A[66] ), .A2(\A[67] ), .ZN(new_n490_));
  INV_X1     g0354(.I(new_n490_), .ZN(new_n491_));
  NAND3_X1   g0355(.A1(new_n489_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  NOR2_X1    g0356(.A1(new_n462_), .A2(new_n471_), .ZN(new_n493_));
  NAND4_X1   g0357(.A1(new_n493_), .A2(new_n480_), .A3(new_n481_), .A4(new_n491_), .ZN(new_n494_));
  AOI21_X1   g0358(.A1(new_n492_), .A2(new_n494_), .B(new_n485_), .ZN(new_n495_));
  NOR2_X1    g0359(.A1(new_n484_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1    g0360(.A1(new_n496_), .A2(\A[63] ), .ZN(new_n497_));
  INV_X1     g0361(.I(\A[63] ), .ZN(new_n498_));
  NAND2_X1   g0362(.A1(new_n489_), .A2(\A[67] ), .ZN(new_n499_));
  NAND2_X1   g0363(.A1(new_n499_), .A2(new_n472_), .ZN(new_n500_));
  NAND2_X1   g0364(.A1(new_n492_), .A2(new_n494_), .ZN(new_n501_));
  NAND2_X1   g0365(.A1(\A[64] ), .A2(\A[65] ), .ZN(new_n502_));
  INV_X1     g0366(.I(new_n502_), .ZN(new_n503_));
  NAND3_X1   g0367(.A1(new_n501_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n504_));
  NAND4_X1   g0368(.A1(new_n483_), .A2(new_n492_), .A3(new_n494_), .A4(new_n503_), .ZN(new_n505_));
  AOI21_X1   g0369(.A1(new_n504_), .A2(new_n505_), .B(new_n498_), .ZN(new_n506_));
  OAI21_X1   g0370(.A1(new_n497_), .A2(new_n506_), .B(new_n147_), .ZN(new_n507_));
  INV_X1     g0371(.I(new_n507_), .ZN(new_n508_));
  NAND2_X1   g0372(.A1(new_n500_), .A2(new_n485_), .ZN(new_n509_));
  NAND2_X1   g0373(.A1(new_n501_), .A2(\A[65] ), .ZN(new_n510_));
  NAND2_X1   g0374(.A1(new_n510_), .A2(new_n509_), .ZN(new_n511_));
  NAND2_X1   g0375(.A1(new_n504_), .A2(new_n505_), .ZN(new_n512_));
  NAND2_X1   g0376(.A1(\A[62] ), .A2(\A[63] ), .ZN(new_n513_));
  INV_X1     g0377(.I(new_n513_), .ZN(new_n514_));
  NAND3_X1   g0378(.A1(new_n512_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n515_));
  NAND4_X1   g0379(.A1(new_n496_), .A2(new_n504_), .A3(new_n505_), .A4(new_n514_), .ZN(new_n516_));
  AOI21_X1   g0380(.A1(new_n515_), .A2(new_n516_), .B(new_n147_), .ZN(new_n517_));
  NOR2_X1    g0381(.A1(new_n508_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1    g0382(.A1(new_n518_), .A2(\A[59] ), .ZN(new_n519_));
  INV_X1     g0383(.I(\A[59] ), .ZN(new_n520_));
  NAND2_X1   g0384(.A1(new_n511_), .A2(new_n498_), .ZN(new_n521_));
  NAND2_X1   g0385(.A1(new_n512_), .A2(\A[63] ), .ZN(new_n522_));
  NAND2_X1   g0386(.A1(new_n522_), .A2(new_n521_), .ZN(new_n523_));
  NAND2_X1   g0387(.A1(new_n515_), .A2(new_n516_), .ZN(new_n524_));
  NAND2_X1   g0388(.A1(\A[60] ), .A2(\A[61] ), .ZN(new_n525_));
  INV_X1     g0389(.I(new_n525_), .ZN(new_n526_));
  NAND3_X1   g0390(.A1(new_n524_), .A2(new_n523_), .A3(new_n526_), .ZN(new_n527_));
  NOR2_X1    g0391(.A1(new_n497_), .A2(new_n506_), .ZN(new_n528_));
  NAND4_X1   g0392(.A1(new_n528_), .A2(new_n515_), .A3(new_n516_), .A4(new_n526_), .ZN(new_n529_));
  AOI21_X1   g0393(.A1(new_n527_), .A2(new_n529_), .B(new_n520_), .ZN(new_n530_));
  NOR2_X1    g0394(.A1(new_n519_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1    g0395(.A1(new_n531_), .A2(\A[57] ), .ZN(new_n532_));
  INV_X1     g0396(.I(\A[57] ), .ZN(new_n533_));
  NAND2_X1   g0397(.A1(new_n524_), .A2(\A[61] ), .ZN(new_n534_));
  NAND2_X1   g0398(.A1(new_n534_), .A2(new_n507_), .ZN(new_n535_));
  NAND2_X1   g0399(.A1(new_n527_), .A2(new_n529_), .ZN(new_n536_));
  NAND2_X1   g0400(.A1(\A[58] ), .A2(\A[59] ), .ZN(new_n537_));
  INV_X1     g0401(.I(new_n537_), .ZN(new_n538_));
  NAND3_X1   g0402(.A1(new_n536_), .A2(new_n535_), .A3(new_n538_), .ZN(new_n539_));
  NAND4_X1   g0403(.A1(new_n518_), .A2(new_n527_), .A3(new_n529_), .A4(new_n538_), .ZN(new_n540_));
  AOI21_X1   g0404(.A1(new_n539_), .A2(new_n540_), .B(new_n533_), .ZN(new_n541_));
  OAI21_X1   g0405(.A1(new_n532_), .A2(new_n541_), .B(new_n146_), .ZN(new_n542_));
  INV_X1     g0406(.I(new_n542_), .ZN(new_n543_));
  NAND2_X1   g0407(.A1(new_n535_), .A2(new_n520_), .ZN(new_n544_));
  NAND2_X1   g0408(.A1(new_n536_), .A2(\A[59] ), .ZN(new_n545_));
  NAND2_X1   g0409(.A1(new_n545_), .A2(new_n544_), .ZN(new_n546_));
  NAND2_X1   g0410(.A1(new_n539_), .A2(new_n540_), .ZN(new_n547_));
  NAND2_X1   g0411(.A1(\A[56] ), .A2(\A[57] ), .ZN(new_n548_));
  INV_X1     g0412(.I(new_n548_), .ZN(new_n549_));
  NAND3_X1   g0413(.A1(new_n547_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  NAND4_X1   g0414(.A1(new_n531_), .A2(new_n539_), .A3(new_n540_), .A4(new_n549_), .ZN(new_n551_));
  AOI21_X1   g0415(.A1(new_n550_), .A2(new_n551_), .B(new_n146_), .ZN(new_n552_));
  NOR2_X1    g0416(.A1(new_n543_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1    g0417(.A1(new_n553_), .A2(\A[53] ), .ZN(new_n554_));
  INV_X1     g0418(.I(\A[53] ), .ZN(new_n555_));
  NAND2_X1   g0419(.A1(new_n546_), .A2(new_n533_), .ZN(new_n556_));
  NAND2_X1   g0420(.A1(new_n547_), .A2(\A[57] ), .ZN(new_n557_));
  NAND2_X1   g0421(.A1(new_n557_), .A2(new_n556_), .ZN(new_n558_));
  NAND2_X1   g0422(.A1(new_n550_), .A2(new_n551_), .ZN(new_n559_));
  NAND2_X1   g0423(.A1(\A[54] ), .A2(\A[55] ), .ZN(new_n560_));
  INV_X1     g0424(.I(new_n560_), .ZN(new_n561_));
  NAND3_X1   g0425(.A1(new_n559_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_));
  NOR2_X1    g0426(.A1(new_n532_), .A2(new_n541_), .ZN(new_n563_));
  NAND4_X1   g0427(.A1(new_n563_), .A2(new_n550_), .A3(new_n551_), .A4(new_n561_), .ZN(new_n564_));
  AOI21_X1   g0428(.A1(new_n562_), .A2(new_n564_), .B(new_n555_), .ZN(new_n565_));
  NOR2_X1    g0429(.A1(new_n554_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1    g0430(.A1(new_n566_), .A2(\A[51] ), .ZN(new_n567_));
  INV_X1     g0431(.I(\A[51] ), .ZN(new_n568_));
  NAND2_X1   g0432(.A1(new_n559_), .A2(\A[55] ), .ZN(new_n569_));
  NAND2_X1   g0433(.A1(new_n569_), .A2(new_n542_), .ZN(new_n570_));
  NAND2_X1   g0434(.A1(new_n562_), .A2(new_n564_), .ZN(new_n571_));
  NAND2_X1   g0435(.A1(\A[52] ), .A2(\A[53] ), .ZN(new_n572_));
  INV_X1     g0436(.I(new_n572_), .ZN(new_n573_));
  NAND3_X1   g0437(.A1(new_n571_), .A2(new_n570_), .A3(new_n573_), .ZN(new_n574_));
  NAND4_X1   g0438(.A1(new_n553_), .A2(new_n562_), .A3(new_n564_), .A4(new_n573_), .ZN(new_n575_));
  AOI21_X1   g0439(.A1(new_n574_), .A2(new_n575_), .B(new_n568_), .ZN(new_n576_));
  OAI21_X1   g0440(.A1(new_n567_), .A2(new_n576_), .B(new_n145_), .ZN(new_n577_));
  INV_X1     g0441(.I(new_n577_), .ZN(new_n578_));
  NAND2_X1   g0442(.A1(new_n570_), .A2(new_n555_), .ZN(new_n579_));
  NAND2_X1   g0443(.A1(new_n571_), .A2(\A[53] ), .ZN(new_n580_));
  NAND2_X1   g0444(.A1(new_n580_), .A2(new_n579_), .ZN(new_n581_));
  NAND2_X1   g0445(.A1(new_n574_), .A2(new_n575_), .ZN(new_n582_));
  NAND2_X1   g0446(.A1(\A[50] ), .A2(\A[51] ), .ZN(new_n583_));
  INV_X1     g0447(.I(new_n583_), .ZN(new_n584_));
  NAND3_X1   g0448(.A1(new_n582_), .A2(new_n581_), .A3(new_n584_), .ZN(new_n585_));
  NAND4_X1   g0449(.A1(new_n566_), .A2(new_n574_), .A3(new_n575_), .A4(new_n584_), .ZN(new_n586_));
  AOI21_X1   g0450(.A1(new_n585_), .A2(new_n586_), .B(new_n145_), .ZN(new_n587_));
  NOR2_X1    g0451(.A1(new_n578_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1    g0452(.A1(new_n588_), .A2(\A[47] ), .ZN(new_n589_));
  INV_X1     g0453(.I(\A[47] ), .ZN(new_n590_));
  NAND2_X1   g0454(.A1(new_n581_), .A2(new_n568_), .ZN(new_n591_));
  NAND2_X1   g0455(.A1(new_n582_), .A2(\A[51] ), .ZN(new_n592_));
  NAND2_X1   g0456(.A1(new_n592_), .A2(new_n591_), .ZN(new_n593_));
  NAND2_X1   g0457(.A1(new_n585_), .A2(new_n586_), .ZN(new_n594_));
  NAND2_X1   g0458(.A1(\A[48] ), .A2(\A[49] ), .ZN(new_n595_));
  INV_X1     g0459(.I(new_n595_), .ZN(new_n596_));
  NAND3_X1   g0460(.A1(new_n594_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n597_));
  NOR2_X1    g0461(.A1(new_n567_), .A2(new_n576_), .ZN(new_n598_));
  NAND4_X1   g0462(.A1(new_n598_), .A2(new_n585_), .A3(new_n586_), .A4(new_n596_), .ZN(new_n599_));
  AOI21_X1   g0463(.A1(new_n597_), .A2(new_n599_), .B(new_n590_), .ZN(new_n600_));
  NOR2_X1    g0464(.A1(new_n589_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1    g0465(.A1(new_n601_), .A2(\A[45] ), .ZN(new_n602_));
  INV_X1     g0466(.I(\A[45] ), .ZN(new_n603_));
  NAND2_X1   g0467(.A1(new_n594_), .A2(\A[49] ), .ZN(new_n604_));
  NAND2_X1   g0468(.A1(new_n604_), .A2(new_n577_), .ZN(new_n605_));
  NAND2_X1   g0469(.A1(new_n597_), .A2(new_n599_), .ZN(new_n606_));
  NAND2_X1   g0470(.A1(\A[46] ), .A2(\A[47] ), .ZN(new_n607_));
  INV_X1     g0471(.I(new_n607_), .ZN(new_n608_));
  NAND3_X1   g0472(.A1(new_n606_), .A2(new_n605_), .A3(new_n608_), .ZN(new_n609_));
  NAND4_X1   g0473(.A1(new_n588_), .A2(new_n597_), .A3(new_n599_), .A4(new_n608_), .ZN(new_n610_));
  AOI21_X1   g0474(.A1(new_n609_), .A2(new_n610_), .B(new_n603_), .ZN(new_n611_));
  OAI21_X1   g0475(.A1(new_n602_), .A2(new_n611_), .B(new_n144_), .ZN(new_n612_));
  INV_X1     g0476(.I(new_n612_), .ZN(new_n613_));
  NAND2_X1   g0477(.A1(new_n605_), .A2(new_n590_), .ZN(new_n614_));
  NAND2_X1   g0478(.A1(new_n606_), .A2(\A[47] ), .ZN(new_n615_));
  NAND2_X1   g0479(.A1(new_n615_), .A2(new_n614_), .ZN(new_n616_));
  NAND2_X1   g0480(.A1(new_n609_), .A2(new_n610_), .ZN(new_n617_));
  NAND2_X1   g0481(.A1(\A[44] ), .A2(\A[45] ), .ZN(new_n618_));
  INV_X1     g0482(.I(new_n618_), .ZN(new_n619_));
  NAND3_X1   g0483(.A1(new_n617_), .A2(new_n616_), .A3(new_n619_), .ZN(new_n620_));
  NAND4_X1   g0484(.A1(new_n601_), .A2(new_n609_), .A3(new_n610_), .A4(new_n619_), .ZN(new_n621_));
  AOI21_X1   g0485(.A1(new_n620_), .A2(new_n621_), .B(new_n144_), .ZN(new_n622_));
  NOR2_X1    g0486(.A1(new_n613_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1    g0487(.A1(new_n623_), .A2(\A[41] ), .ZN(new_n624_));
  INV_X1     g0488(.I(\A[41] ), .ZN(new_n625_));
  NAND2_X1   g0489(.A1(new_n616_), .A2(new_n603_), .ZN(new_n626_));
  NAND2_X1   g0490(.A1(new_n617_), .A2(\A[45] ), .ZN(new_n627_));
  NAND2_X1   g0491(.A1(new_n627_), .A2(new_n626_), .ZN(new_n628_));
  NAND2_X1   g0492(.A1(new_n620_), .A2(new_n621_), .ZN(new_n629_));
  NAND2_X1   g0493(.A1(\A[42] ), .A2(\A[43] ), .ZN(new_n630_));
  INV_X1     g0494(.I(new_n630_), .ZN(new_n631_));
  NAND3_X1   g0495(.A1(new_n629_), .A2(new_n628_), .A3(new_n631_), .ZN(new_n632_));
  NOR2_X1    g0496(.A1(new_n602_), .A2(new_n611_), .ZN(new_n633_));
  NAND4_X1   g0497(.A1(new_n633_), .A2(new_n620_), .A3(new_n621_), .A4(new_n631_), .ZN(new_n634_));
  AOI21_X1   g0498(.A1(new_n632_), .A2(new_n634_), .B(new_n625_), .ZN(new_n635_));
  NOR2_X1    g0499(.A1(new_n624_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1    g0500(.A1(new_n636_), .A2(\A[39] ), .ZN(new_n637_));
  INV_X1     g0501(.I(\A[39] ), .ZN(new_n638_));
  NAND2_X1   g0502(.A1(new_n629_), .A2(\A[43] ), .ZN(new_n639_));
  NAND2_X1   g0503(.A1(new_n639_), .A2(new_n612_), .ZN(new_n640_));
  NAND2_X1   g0504(.A1(new_n632_), .A2(new_n634_), .ZN(new_n641_));
  NAND2_X1   g0505(.A1(\A[40] ), .A2(\A[41] ), .ZN(new_n642_));
  INV_X1     g0506(.I(new_n642_), .ZN(new_n643_));
  NAND3_X1   g0507(.A1(new_n641_), .A2(new_n640_), .A3(new_n643_), .ZN(new_n644_));
  NAND4_X1   g0508(.A1(new_n623_), .A2(new_n632_), .A3(new_n634_), .A4(new_n643_), .ZN(new_n645_));
  AOI21_X1   g0509(.A1(new_n644_), .A2(new_n645_), .B(new_n638_), .ZN(new_n646_));
  OAI21_X1   g0510(.A1(new_n637_), .A2(new_n646_), .B(new_n143_), .ZN(new_n647_));
  INV_X1     g0511(.I(new_n647_), .ZN(new_n648_));
  NAND2_X1   g0512(.A1(new_n640_), .A2(new_n625_), .ZN(new_n649_));
  NAND2_X1   g0513(.A1(new_n641_), .A2(\A[41] ), .ZN(new_n650_));
  NAND2_X1   g0514(.A1(new_n650_), .A2(new_n649_), .ZN(new_n651_));
  NAND2_X1   g0515(.A1(new_n644_), .A2(new_n645_), .ZN(new_n652_));
  NAND2_X1   g0516(.A1(\A[38] ), .A2(\A[39] ), .ZN(new_n653_));
  INV_X1     g0517(.I(new_n653_), .ZN(new_n654_));
  NAND3_X1   g0518(.A1(new_n652_), .A2(new_n651_), .A3(new_n654_), .ZN(new_n655_));
  NAND4_X1   g0519(.A1(new_n636_), .A2(new_n644_), .A3(new_n645_), .A4(new_n654_), .ZN(new_n656_));
  AOI21_X1   g0520(.A1(new_n655_), .A2(new_n656_), .B(new_n143_), .ZN(new_n657_));
  NOR2_X1    g0521(.A1(new_n648_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1    g0522(.A1(new_n658_), .A2(\A[35] ), .ZN(new_n659_));
  INV_X1     g0523(.I(\A[35] ), .ZN(new_n660_));
  NAND2_X1   g0524(.A1(new_n651_), .A2(new_n638_), .ZN(new_n661_));
  NAND2_X1   g0525(.A1(new_n652_), .A2(\A[39] ), .ZN(new_n662_));
  NAND2_X1   g0526(.A1(new_n662_), .A2(new_n661_), .ZN(new_n663_));
  NAND2_X1   g0527(.A1(new_n655_), .A2(new_n656_), .ZN(new_n664_));
  NAND2_X1   g0528(.A1(\A[36] ), .A2(\A[37] ), .ZN(new_n665_));
  INV_X1     g0529(.I(new_n665_), .ZN(new_n666_));
  NAND3_X1   g0530(.A1(new_n664_), .A2(new_n663_), .A3(new_n666_), .ZN(new_n667_));
  NOR2_X1    g0531(.A1(new_n637_), .A2(new_n646_), .ZN(new_n668_));
  NAND4_X1   g0532(.A1(new_n668_), .A2(new_n655_), .A3(new_n656_), .A4(new_n666_), .ZN(new_n669_));
  AOI21_X1   g0533(.A1(new_n667_), .A2(new_n669_), .B(new_n660_), .ZN(new_n670_));
  NOR2_X1    g0534(.A1(new_n659_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1    g0535(.A1(new_n671_), .A2(\A[33] ), .ZN(new_n672_));
  INV_X1     g0536(.I(\A[33] ), .ZN(new_n673_));
  NAND2_X1   g0537(.A1(new_n664_), .A2(\A[37] ), .ZN(new_n674_));
  NAND2_X1   g0538(.A1(new_n674_), .A2(new_n647_), .ZN(new_n675_));
  NAND2_X1   g0539(.A1(new_n667_), .A2(new_n669_), .ZN(new_n676_));
  NAND2_X1   g0540(.A1(\A[34] ), .A2(\A[35] ), .ZN(new_n677_));
  INV_X1     g0541(.I(new_n677_), .ZN(new_n678_));
  NAND3_X1   g0542(.A1(new_n676_), .A2(new_n675_), .A3(new_n678_), .ZN(new_n679_));
  NAND4_X1   g0543(.A1(new_n658_), .A2(new_n667_), .A3(new_n669_), .A4(new_n678_), .ZN(new_n680_));
  AOI21_X1   g0544(.A1(new_n679_), .A2(new_n680_), .B(new_n673_), .ZN(new_n681_));
  OAI21_X1   g0545(.A1(new_n672_), .A2(new_n681_), .B(new_n142_), .ZN(new_n682_));
  INV_X1     g0546(.I(new_n682_), .ZN(new_n683_));
  NAND2_X1   g0547(.A1(new_n675_), .A2(new_n660_), .ZN(new_n684_));
  NAND2_X1   g0548(.A1(new_n676_), .A2(\A[35] ), .ZN(new_n685_));
  NAND2_X1   g0549(.A1(new_n685_), .A2(new_n684_), .ZN(new_n686_));
  NAND2_X1   g0550(.A1(new_n679_), .A2(new_n680_), .ZN(new_n687_));
  NAND2_X1   g0551(.A1(\A[32] ), .A2(\A[33] ), .ZN(new_n688_));
  INV_X1     g0552(.I(new_n688_), .ZN(new_n689_));
  NAND3_X1   g0553(.A1(new_n687_), .A2(new_n686_), .A3(new_n689_), .ZN(new_n690_));
  NAND4_X1   g0554(.A1(new_n671_), .A2(new_n679_), .A3(new_n680_), .A4(new_n689_), .ZN(new_n691_));
  AOI21_X1   g0555(.A1(new_n690_), .A2(new_n691_), .B(new_n142_), .ZN(new_n692_));
  NOR2_X1    g0556(.A1(new_n683_), .A2(new_n692_), .ZN(new_n693_));
  NOR2_X1    g0557(.A1(new_n693_), .A2(\A[29] ), .ZN(new_n694_));
  INV_X1     g0558(.I(\A[29] ), .ZN(new_n695_));
  NAND2_X1   g0559(.A1(new_n686_), .A2(new_n673_), .ZN(new_n696_));
  NAND2_X1   g0560(.A1(new_n687_), .A2(\A[33] ), .ZN(new_n697_));
  NAND2_X1   g0561(.A1(new_n697_), .A2(new_n696_), .ZN(new_n698_));
  NAND2_X1   g0562(.A1(new_n690_), .A2(new_n691_), .ZN(new_n699_));
  NAND2_X1   g0563(.A1(\A[30] ), .A2(\A[31] ), .ZN(new_n700_));
  INV_X1     g0564(.I(new_n700_), .ZN(new_n701_));
  NAND3_X1   g0565(.A1(new_n699_), .A2(new_n698_), .A3(new_n701_), .ZN(new_n702_));
  NOR2_X1    g0566(.A1(new_n672_), .A2(new_n681_), .ZN(new_n703_));
  NAND4_X1   g0567(.A1(new_n703_), .A2(new_n690_), .A3(new_n691_), .A4(new_n701_), .ZN(new_n704_));
  AOI21_X1   g0568(.A1(new_n702_), .A2(new_n704_), .B(new_n695_), .ZN(new_n705_));
  NOR2_X1    g0569(.A1(new_n694_), .A2(new_n705_), .ZN(new_n706_));
  NOR2_X1    g0570(.A1(new_n706_), .A2(\A[27] ), .ZN(new_n707_));
  INV_X1     g0571(.I(\A[27] ), .ZN(new_n708_));
  NAND2_X1   g0572(.A1(new_n699_), .A2(\A[31] ), .ZN(new_n709_));
  NAND2_X1   g0573(.A1(new_n709_), .A2(new_n682_), .ZN(new_n710_));
  NAND2_X1   g0574(.A1(new_n702_), .A2(new_n704_), .ZN(new_n711_));
  NAND2_X1   g0575(.A1(\A[28] ), .A2(\A[29] ), .ZN(new_n712_));
  INV_X1     g0576(.I(new_n712_), .ZN(new_n713_));
  NAND3_X1   g0577(.A1(new_n711_), .A2(new_n710_), .A3(new_n713_), .ZN(new_n714_));
  NAND4_X1   g0578(.A1(new_n693_), .A2(new_n702_), .A3(new_n704_), .A4(new_n713_), .ZN(new_n715_));
  AOI21_X1   g0579(.A1(new_n714_), .A2(new_n715_), .B(new_n708_), .ZN(new_n716_));
  OAI21_X1   g0580(.A1(new_n707_), .A2(new_n716_), .B(new_n141_), .ZN(new_n717_));
  INV_X1     g0581(.I(new_n717_), .ZN(new_n718_));
  NAND2_X1   g0582(.A1(new_n710_), .A2(new_n695_), .ZN(new_n719_));
  NAND2_X1   g0583(.A1(new_n711_), .A2(\A[29] ), .ZN(new_n720_));
  NAND2_X1   g0584(.A1(new_n720_), .A2(new_n719_), .ZN(new_n721_));
  NAND2_X1   g0585(.A1(new_n714_), .A2(new_n715_), .ZN(new_n722_));
  NAND2_X1   g0586(.A1(\A[26] ), .A2(\A[27] ), .ZN(new_n723_));
  INV_X1     g0587(.I(new_n723_), .ZN(new_n724_));
  NAND3_X1   g0588(.A1(new_n722_), .A2(new_n721_), .A3(new_n724_), .ZN(new_n725_));
  NAND4_X1   g0589(.A1(new_n706_), .A2(new_n714_), .A3(new_n715_), .A4(new_n724_), .ZN(new_n726_));
  AOI21_X1   g0590(.A1(new_n725_), .A2(new_n726_), .B(new_n141_), .ZN(new_n727_));
  NOR2_X1    g0591(.A1(new_n718_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1    g0592(.A1(new_n728_), .A2(\A[23] ), .ZN(new_n729_));
  INV_X1     g0593(.I(\A[23] ), .ZN(new_n730_));
  NAND2_X1   g0594(.A1(new_n721_), .A2(new_n708_), .ZN(new_n731_));
  NAND2_X1   g0595(.A1(new_n722_), .A2(\A[27] ), .ZN(new_n732_));
  NAND2_X1   g0596(.A1(new_n732_), .A2(new_n731_), .ZN(new_n733_));
  NAND2_X1   g0597(.A1(new_n725_), .A2(new_n726_), .ZN(new_n734_));
  NAND2_X1   g0598(.A1(\A[24] ), .A2(\A[25] ), .ZN(new_n735_));
  INV_X1     g0599(.I(new_n735_), .ZN(new_n736_));
  NAND3_X1   g0600(.A1(new_n734_), .A2(new_n733_), .A3(new_n736_), .ZN(new_n737_));
  NOR2_X1    g0601(.A1(new_n707_), .A2(new_n716_), .ZN(new_n738_));
  NAND4_X1   g0602(.A1(new_n738_), .A2(new_n725_), .A3(new_n726_), .A4(new_n736_), .ZN(new_n739_));
  AOI21_X1   g0603(.A1(new_n737_), .A2(new_n739_), .B(new_n730_), .ZN(new_n740_));
  NOR2_X1    g0604(.A1(new_n729_), .A2(new_n740_), .ZN(new_n741_));
  NOR2_X1    g0605(.A1(new_n741_), .A2(\A[21] ), .ZN(new_n742_));
  INV_X1     g0606(.I(\A[21] ), .ZN(new_n743_));
  NAND2_X1   g0607(.A1(new_n734_), .A2(\A[25] ), .ZN(new_n744_));
  NAND2_X1   g0608(.A1(new_n744_), .A2(new_n717_), .ZN(new_n745_));
  NAND2_X1   g0609(.A1(new_n737_), .A2(new_n739_), .ZN(new_n746_));
  NAND2_X1   g0610(.A1(\A[22] ), .A2(\A[23] ), .ZN(new_n747_));
  INV_X1     g0611(.I(new_n747_), .ZN(new_n748_));
  NAND3_X1   g0612(.A1(new_n746_), .A2(new_n745_), .A3(new_n748_), .ZN(new_n749_));
  NAND4_X1   g0613(.A1(new_n728_), .A2(new_n737_), .A3(new_n739_), .A4(new_n748_), .ZN(new_n750_));
  AOI21_X1   g0614(.A1(new_n749_), .A2(new_n750_), .B(new_n743_), .ZN(new_n751_));
  OAI21_X1   g0615(.A1(new_n742_), .A2(new_n751_), .B(new_n140_), .ZN(new_n752_));
  INV_X1     g0616(.I(new_n752_), .ZN(new_n753_));
  NAND2_X1   g0617(.A1(new_n745_), .A2(new_n730_), .ZN(new_n754_));
  NAND2_X1   g0618(.A1(new_n746_), .A2(\A[23] ), .ZN(new_n755_));
  NAND2_X1   g0619(.A1(new_n755_), .A2(new_n754_), .ZN(new_n756_));
  NAND2_X1   g0620(.A1(new_n749_), .A2(new_n750_), .ZN(new_n757_));
  NAND2_X1   g0621(.A1(\A[20] ), .A2(\A[21] ), .ZN(new_n758_));
  INV_X1     g0622(.I(new_n758_), .ZN(new_n759_));
  NAND3_X1   g0623(.A1(new_n757_), .A2(new_n756_), .A3(new_n759_), .ZN(new_n760_));
  NAND4_X1   g0624(.A1(new_n741_), .A2(new_n749_), .A3(new_n750_), .A4(new_n759_), .ZN(new_n761_));
  AOI21_X1   g0625(.A1(new_n760_), .A2(new_n761_), .B(new_n140_), .ZN(new_n762_));
  NOR2_X1    g0626(.A1(new_n753_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1    g0627(.A1(new_n763_), .A2(\A[17] ), .ZN(new_n764_));
  INV_X1     g0628(.I(\A[17] ), .ZN(new_n765_));
  NAND2_X1   g0629(.A1(new_n756_), .A2(new_n743_), .ZN(new_n766_));
  NAND2_X1   g0630(.A1(new_n757_), .A2(\A[21] ), .ZN(new_n767_));
  NAND2_X1   g0631(.A1(new_n767_), .A2(new_n766_), .ZN(new_n768_));
  NAND2_X1   g0632(.A1(new_n760_), .A2(new_n761_), .ZN(new_n769_));
  NAND2_X1   g0633(.A1(\A[18] ), .A2(\A[19] ), .ZN(new_n770_));
  INV_X1     g0634(.I(new_n770_), .ZN(new_n771_));
  NAND3_X1   g0635(.A1(new_n769_), .A2(new_n768_), .A3(new_n771_), .ZN(new_n772_));
  NOR2_X1    g0636(.A1(new_n742_), .A2(new_n751_), .ZN(new_n773_));
  NAND4_X1   g0637(.A1(new_n773_), .A2(new_n760_), .A3(new_n761_), .A4(new_n771_), .ZN(new_n774_));
  AOI21_X1   g0638(.A1(new_n772_), .A2(new_n774_), .B(new_n765_), .ZN(new_n775_));
  NOR2_X1    g0639(.A1(new_n764_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1    g0640(.A1(new_n776_), .A2(\A[15] ), .ZN(new_n777_));
  INV_X1     g0641(.I(\A[15] ), .ZN(new_n778_));
  NAND2_X1   g0642(.A1(new_n769_), .A2(\A[19] ), .ZN(new_n779_));
  NAND2_X1   g0643(.A1(new_n779_), .A2(new_n752_), .ZN(new_n780_));
  NAND2_X1   g0644(.A1(new_n772_), .A2(new_n774_), .ZN(new_n781_));
  NAND2_X1   g0645(.A1(\A[16] ), .A2(\A[17] ), .ZN(new_n782_));
  INV_X1     g0646(.I(new_n782_), .ZN(new_n783_));
  NAND3_X1   g0647(.A1(new_n781_), .A2(new_n780_), .A3(new_n783_), .ZN(new_n784_));
  NAND4_X1   g0648(.A1(new_n763_), .A2(new_n772_), .A3(new_n774_), .A4(new_n783_), .ZN(new_n785_));
  AOI21_X1   g0649(.A1(new_n784_), .A2(new_n785_), .B(new_n778_), .ZN(new_n786_));
  OAI21_X1   g0650(.A1(new_n777_), .A2(new_n786_), .B(new_n139_), .ZN(new_n787_));
  NAND2_X1   g0651(.A1(new_n780_), .A2(new_n765_), .ZN(new_n788_));
  NAND2_X1   g0652(.A1(new_n781_), .A2(\A[17] ), .ZN(new_n789_));
  NAND2_X1   g0653(.A1(new_n789_), .A2(new_n788_), .ZN(new_n790_));
  NAND2_X1   g0654(.A1(new_n784_), .A2(new_n785_), .ZN(new_n791_));
  NAND2_X1   g0655(.A1(\A[14] ), .A2(\A[15] ), .ZN(new_n792_));
  INV_X1     g0656(.I(new_n792_), .ZN(new_n793_));
  NAND3_X1   g0657(.A1(new_n791_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n794_));
  NAND4_X1   g0658(.A1(new_n776_), .A2(new_n784_), .A3(new_n785_), .A4(new_n793_), .ZN(new_n795_));
  NAND2_X1   g0659(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1   g0660(.A1(new_n796_), .A2(\A[13] ), .ZN(new_n797_));
  NAND2_X1   g0661(.A1(new_n797_), .A2(new_n787_), .ZN(new_n798_));
  NAND2_X1   g0662(.A1(new_n798_), .A2(new_n138_), .ZN(new_n799_));
  NAND2_X1   g0663(.A1(new_n790_), .A2(new_n778_), .ZN(new_n800_));
  NAND2_X1   g0664(.A1(new_n791_), .A2(\A[15] ), .ZN(new_n801_));
  NAND2_X1   g0665(.A1(new_n801_), .A2(new_n800_), .ZN(new_n802_));
  NAND2_X1   g0666(.A1(\A[12] ), .A2(\A[13] ), .ZN(new_n803_));
  INV_X1     g0667(.I(new_n803_), .ZN(new_n804_));
  NAND3_X1   g0668(.A1(new_n796_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n805_));
  NOR2_X1    g0669(.A1(new_n777_), .A2(new_n786_), .ZN(new_n806_));
  NAND4_X1   g0670(.A1(new_n806_), .A2(new_n794_), .A3(new_n795_), .A4(new_n804_), .ZN(new_n807_));
  NAND2_X1   g0671(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1   g0672(.A1(new_n808_), .A2(\A[11] ), .ZN(new_n809_));
  NAND2_X1   g0673(.A1(new_n809_), .A2(new_n799_), .ZN(new_n810_));
  NAND2_X1   g0674(.A1(new_n810_), .A2(new_n137_), .ZN(new_n811_));
  AND2_X2    g0675(.A1(\A[10] ), .A2(\A[11] ), .Z(new_n812_));
  NAND3_X1   g0676(.A1(new_n808_), .A2(new_n798_), .A3(new_n812_), .ZN(new_n813_));
  INV_X1     g0677(.I(new_n787_), .ZN(new_n814_));
  AOI21_X1   g0678(.A1(new_n794_), .A2(new_n795_), .B(new_n139_), .ZN(new_n815_));
  NOR2_X1    g0679(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1   g0680(.A1(new_n816_), .A2(new_n805_), .A3(new_n807_), .A4(new_n812_), .ZN(new_n817_));
  NAND2_X1   g0681(.A1(new_n813_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1   g0682(.A1(new_n818_), .A2(\A[9] ), .ZN(new_n819_));
  NAND2_X1   g0683(.A1(new_n819_), .A2(new_n811_), .ZN(new_n820_));
  AND2_X2    g0684(.A1(\A[6] ), .A2(\A[7] ), .Z(new_n821_));
  INV_X1     g0685(.I(\A[8] ), .ZN(new_n822_));
  NOR2_X1    g0686(.A1(new_n822_), .A2(new_n137_), .ZN(new_n823_));
  NAND3_X1   g0687(.A1(new_n818_), .A2(new_n810_), .A3(new_n823_), .ZN(new_n824_));
  NOR2_X1    g0688(.A1(new_n816_), .A2(\A[11] ), .ZN(new_n825_));
  AOI21_X1   g0689(.A1(new_n805_), .A2(new_n807_), .B(new_n138_), .ZN(new_n826_));
  NOR2_X1    g0690(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1   g0691(.A1(new_n827_), .A2(new_n813_), .A3(new_n817_), .A4(new_n823_), .ZN(new_n828_));
  NAND2_X1   g0692(.A1(new_n824_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1   g0693(.A1(new_n829_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n830_));
  NOR2_X1    g0694(.A1(new_n827_), .A2(\A[9] ), .ZN(new_n831_));
  AOI21_X1   g0695(.A1(new_n813_), .A2(new_n817_), .B(new_n137_), .ZN(new_n832_));
  NOR2_X1    g0696(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND4_X1   g0697(.A1(new_n833_), .A2(new_n824_), .A3(new_n821_), .A4(new_n828_), .ZN(new_n834_));
  NAND2_X1   g0698(.A1(new_n830_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1     g0699(.I(\A[7] ), .ZN(new_n836_));
  OAI21_X1   g0700(.A1(new_n831_), .A2(new_n832_), .B(new_n836_), .ZN(new_n837_));
  INV_X1     g0701(.I(new_n837_), .ZN(new_n838_));
  AOI21_X1   g0702(.A1(new_n824_), .A2(new_n828_), .B(new_n836_), .ZN(new_n839_));
  NOR2_X1    g0703(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1     g0704(.I(\A[1] ), .ZN(new_n841_));
  INV_X1     g0705(.I(\A[3] ), .ZN(new_n842_));
  NOR3_X1    g0706(.A1(new_n841_), .A2(new_n842_), .A3(\A[2] ), .ZN(new_n843_));
  OAI21_X1   g0707(.A1(new_n840_), .A2(\A[5] ), .B(new_n843_), .ZN(new_n844_));
  AOI21_X1   g0708(.A1(\A[5] ), .A2(new_n835_), .B(new_n844_), .ZN(new_n845_));
  INV_X1     g0709(.I(new_n843_), .ZN(new_n846_));
  NAND2_X1   g0710(.A1(new_n829_), .A2(\A[7] ), .ZN(new_n847_));
  NAND2_X1   g0711(.A1(new_n847_), .A2(new_n837_), .ZN(new_n848_));
  AND2_X2    g0712(.A1(\A[4] ), .A2(\A[5] ), .Z(new_n849_));
  NAND3_X1   g0713(.A1(new_n835_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  NAND4_X1   g0714(.A1(new_n840_), .A2(new_n830_), .A3(new_n834_), .A4(new_n849_), .ZN(new_n851_));
  AOI21_X1   g0715(.A1(new_n850_), .A2(new_n851_), .B(new_n846_), .ZN(new_n852_));
  XOR2_X1    g0716(.A1(new_n852_), .A2(new_n845_), .Z(\P[0] ));
  NOR2_X1    g0717(.A1(\A[76] ), .A2(\A[77] ), .ZN(new_n854_));
  INV_X1     g0718(.I(new_n854_), .ZN(new_n855_));
  NOR2_X1    g0719(.A1(\A[122] ), .A2(\A[123] ), .ZN(new_n856_));
  OR2_X2     g0720(.A1(\A[124] ), .A2(\A[125] ), .Z(new_n857_));
  NAND3_X1   g0721(.A1(new_n857_), .A2(\A[121] ), .A3(new_n856_), .ZN(new_n858_));
  NAND2_X1   g0722(.A1(new_n858_), .A2(\A[120] ), .ZN(new_n859_));
  INV_X1     g0723(.I(new_n857_), .ZN(new_n860_));
  NAND4_X1   g0724(.A1(new_n856_), .A2(new_n162_), .A3(new_n170_), .A4(\A[120] ), .ZN(new_n861_));
  XOR2_X1    g0725(.A1(new_n859_), .A2(new_n861_), .Z(new_n862_));
  NOR2_X1    g0726(.A1(new_n862_), .A2(new_n214_), .ZN(new_n863_));
  NOR2_X1    g0727(.A1(\A[126] ), .A2(\A[127] ), .ZN(new_n864_));
  INV_X1     g0728(.I(new_n864_), .ZN(new_n865_));
  NAND2_X1   g0729(.A1(new_n860_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1   g0730(.A1(new_n866_), .A2(new_n856_), .B(new_n195_), .ZN(new_n867_));
  NAND2_X1   g0731(.A1(new_n862_), .A2(new_n197_), .ZN(new_n868_));
  XOR2_X1    g0732(.A1(new_n868_), .A2(new_n867_), .Z(new_n869_));
  NOR2_X1    g0733(.A1(new_n869_), .A2(new_n214_), .ZN(new_n870_));
  XOR2_X1    g0734(.A1(new_n870_), .A2(new_n863_), .Z(new_n871_));
  OR2_X2     g0735(.A1(new_n871_), .A2(new_n239_), .Z(new_n872_));
  NAND2_X1   g0736(.A1(new_n869_), .A2(new_n235_), .ZN(new_n873_));
  NAND2_X1   g0737(.A1(new_n871_), .A2(new_n235_), .ZN(new_n874_));
  XOR2_X1    g0738(.A1(new_n874_), .A2(new_n873_), .Z(new_n875_));
  NAND2_X1   g0739(.A1(new_n875_), .A2(new_n240_), .ZN(new_n876_));
  XOR2_X1    g0740(.A1(new_n876_), .A2(new_n872_), .Z(new_n877_));
  OR2_X2     g0741(.A1(new_n877_), .A2(new_n266_), .Z(new_n878_));
  OR2_X2     g0742(.A1(new_n875_), .A2(new_n253_), .Z(new_n879_));
  NAND2_X1   g0743(.A1(new_n877_), .A2(new_n262_), .ZN(new_n880_));
  XOR2_X1    g0744(.A1(new_n880_), .A2(new_n879_), .Z(new_n881_));
  NAND2_X1   g0745(.A1(new_n881_), .A2(new_n267_), .ZN(new_n882_));
  XOR2_X1    g0746(.A1(new_n882_), .A2(new_n878_), .Z(new_n883_));
  NOR2_X1    g0747(.A1(new_n883_), .A2(new_n285_), .ZN(new_n884_));
  OR2_X2     g0748(.A1(new_n881_), .A2(new_n275_), .Z(new_n885_));
  NAND2_X1   g0749(.A1(new_n883_), .A2(new_n276_), .ZN(new_n886_));
  XOR2_X1    g0750(.A1(new_n886_), .A2(new_n885_), .Z(new_n887_));
  NAND2_X1   g0751(.A1(new_n887_), .A2(new_n286_), .ZN(new_n888_));
  XOR2_X1    g0752(.A1(new_n888_), .A2(new_n884_), .Z(new_n889_));
  NAND2_X1   g0753(.A1(new_n889_), .A2(new_n305_), .ZN(new_n890_));
  NAND2_X1   g0754(.A1(new_n294_), .A2(new_n284_), .ZN(new_n891_));
  MUX2_X1    g0755(.I0(new_n887_), .I1(new_n889_), .S(new_n891_), .Z(new_n892_));
  NAND2_X1   g0756(.A1(new_n892_), .A2(new_n305_), .ZN(new_n893_));
  XOR2_X1    g0757(.A1(new_n893_), .A2(new_n890_), .Z(new_n894_));
  NOR2_X1    g0758(.A1(new_n894_), .A2(new_n324_), .ZN(new_n895_));
  NOR2_X1    g0759(.A1(new_n892_), .A2(new_n313_), .ZN(new_n896_));
  NAND2_X1   g0760(.A1(new_n894_), .A2(new_n314_), .ZN(new_n897_));
  XNOR2_X1   g0761(.A1(new_n897_), .A2(new_n896_), .ZN(new_n898_));
  NAND2_X1   g0762(.A1(new_n898_), .A2(new_n325_), .ZN(new_n899_));
  XNOR2_X1   g0763(.A1(new_n899_), .A2(new_n895_), .ZN(new_n900_));
  NOR2_X1    g0764(.A1(new_n900_), .A2(new_n347_), .ZN(new_n901_));
  NOR2_X1    g0765(.A1(new_n898_), .A2(new_n335_), .ZN(new_n902_));
  NAND2_X1   g0766(.A1(new_n900_), .A2(new_n336_), .ZN(new_n903_));
  XNOR2_X1   g0767(.A1(new_n903_), .A2(new_n902_), .ZN(new_n904_));
  NAND2_X1   g0768(.A1(new_n904_), .A2(new_n348_), .ZN(new_n905_));
  XNOR2_X1   g0769(.A1(new_n905_), .A2(new_n901_), .ZN(new_n906_));
  OR2_X2     g0770(.A1(new_n906_), .A2(new_n368_), .Z(new_n907_));
  NOR2_X1    g0771(.A1(new_n904_), .A2(new_n357_), .ZN(new_n908_));
  NAND2_X1   g0772(.A1(new_n906_), .A2(new_n358_), .ZN(new_n909_));
  XNOR2_X1   g0773(.A1(new_n909_), .A2(new_n908_), .ZN(new_n910_));
  NAND2_X1   g0774(.A1(new_n910_), .A2(new_n369_), .ZN(new_n911_));
  XOR2_X1    g0775(.A1(new_n911_), .A2(new_n907_), .Z(new_n912_));
  OR2_X2     g0776(.A1(new_n912_), .A2(new_n390_), .Z(new_n913_));
  OR2_X2     g0777(.A1(new_n910_), .A2(new_n377_), .Z(new_n914_));
  NAND2_X1   g0778(.A1(new_n912_), .A2(new_n378_), .ZN(new_n915_));
  XOR2_X1    g0779(.A1(new_n915_), .A2(new_n914_), .Z(new_n916_));
  NAND2_X1   g0780(.A1(new_n916_), .A2(new_n391_), .ZN(new_n917_));
  XOR2_X1    g0781(.A1(new_n917_), .A2(new_n913_), .Z(new_n918_));
  NOR2_X1    g0782(.A1(new_n918_), .A2(new_n412_), .ZN(new_n919_));
  OR2_X2     g0783(.A1(new_n916_), .A2(new_n403_), .Z(new_n920_));
  NAND2_X1   g0784(.A1(new_n918_), .A2(new_n404_), .ZN(new_n921_));
  XOR2_X1    g0785(.A1(new_n921_), .A2(new_n920_), .Z(new_n922_));
  NAND2_X1   g0786(.A1(new_n922_), .A2(new_n413_), .ZN(new_n923_));
  XOR2_X1    g0787(.A1(new_n923_), .A2(new_n919_), .Z(new_n924_));
  NOR2_X1    g0788(.A1(new_n924_), .A2(new_n855_), .ZN(new_n925_));
  NOR2_X1    g0789(.A1(\A[78] ), .A2(\A[79] ), .ZN(new_n926_));
  INV_X1     g0790(.I(new_n926_), .ZN(new_n927_));
  AND2_X2    g0791(.A1(new_n922_), .A2(new_n926_), .Z(new_n928_));
  AOI21_X1   g0792(.A1(new_n924_), .A2(new_n927_), .B(new_n928_), .ZN(new_n929_));
  AOI21_X1   g0793(.A1(new_n929_), .A2(new_n855_), .B(new_n925_), .ZN(new_n930_));
  NOR3_X1    g0794(.A1(new_n930_), .A2(new_n443_), .A3(new_n929_), .ZN(new_n931_));
  AND4_X2    g0795(.A1(new_n444_), .A2(new_n929_), .A3(new_n924_), .A4(new_n854_), .Z(new_n932_));
  NOR2_X1    g0796(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NOR3_X1    g0797(.A1(new_n933_), .A2(new_n455_), .A3(new_n930_), .ZN(new_n934_));
  AND3_X2    g0798(.A1(new_n933_), .A2(new_n456_), .A3(new_n930_), .Z(new_n935_));
  NOR2_X1    g0799(.A1(new_n935_), .A2(new_n934_), .ZN(new_n936_));
  NOR3_X1    g0800(.A1(new_n936_), .A2(new_n467_), .A3(new_n933_), .ZN(new_n937_));
  INV_X1     g0801(.I(new_n933_), .ZN(new_n938_));
  NOR4_X1    g0802(.A1(new_n935_), .A2(new_n467_), .A3(new_n938_), .A4(new_n934_), .ZN(new_n939_));
  NOR2_X1    g0803(.A1(new_n937_), .A2(new_n939_), .ZN(new_n940_));
  NOR4_X1    g0804(.A1(new_n940_), .A2(new_n478_), .A3(new_n490_), .A4(new_n936_), .ZN(new_n941_));
  INV_X1     g0805(.I(new_n940_), .ZN(new_n942_));
  NOR3_X1    g0806(.A1(new_n940_), .A2(new_n478_), .A3(new_n936_), .ZN(new_n943_));
  INV_X1     g0807(.I(new_n936_), .ZN(new_n944_));
  NOR4_X1    g0808(.A1(new_n937_), .A2(new_n478_), .A3(new_n944_), .A4(new_n939_), .ZN(new_n945_));
  NOR4_X1    g0809(.A1(new_n943_), .A2(new_n490_), .A3(new_n942_), .A4(new_n945_), .ZN(new_n946_));
  NOR2_X1    g0810(.A1(new_n946_), .A2(new_n941_), .ZN(new_n947_));
  NOR2_X1    g0811(.A1(new_n943_), .A2(new_n945_), .ZN(new_n948_));
  NOR4_X1    g0812(.A1(new_n948_), .A2(new_n490_), .A3(new_n502_), .A4(new_n940_), .ZN(new_n949_));
  INV_X1     g0813(.I(new_n948_), .ZN(new_n950_));
  NOR4_X1    g0814(.A1(new_n950_), .A2(new_n502_), .A3(new_n941_), .A4(new_n946_), .ZN(new_n951_));
  NOR2_X1    g0815(.A1(new_n951_), .A2(new_n949_), .ZN(new_n952_));
  NOR4_X1    g0816(.A1(new_n952_), .A2(new_n513_), .A3(new_n525_), .A4(new_n947_), .ZN(new_n953_));
  INV_X1     g0817(.I(new_n953_), .ZN(new_n954_));
  NOR4_X1    g0818(.A1(new_n947_), .A2(new_n502_), .A3(new_n513_), .A4(new_n948_), .ZN(new_n955_));
  INV_X1     g0819(.I(new_n947_), .ZN(new_n956_));
  NOR4_X1    g0820(.A1(new_n951_), .A2(new_n956_), .A3(new_n513_), .A4(new_n949_), .ZN(new_n957_));
  NOR2_X1    g0821(.A1(new_n957_), .A2(new_n955_), .ZN(new_n958_));
  NAND3_X1   g0822(.A1(new_n958_), .A2(new_n526_), .A3(new_n952_), .ZN(new_n959_));
  NAND2_X1   g0823(.A1(new_n959_), .A2(new_n954_), .ZN(new_n960_));
  NOR4_X1    g0824(.A1(new_n958_), .A2(new_n525_), .A3(new_n537_), .A4(new_n952_), .ZN(new_n961_));
  INV_X1     g0825(.I(new_n961_), .ZN(new_n962_));
  NAND4_X1   g0826(.A1(new_n959_), .A2(new_n958_), .A3(new_n954_), .A4(new_n538_), .ZN(new_n963_));
  NAND2_X1   g0827(.A1(new_n963_), .A2(new_n962_), .ZN(new_n964_));
  NAND4_X1   g0828(.A1(new_n964_), .A2(new_n549_), .A3(new_n561_), .A4(new_n960_), .ZN(new_n965_));
  INV_X1     g0829(.I(new_n958_), .ZN(new_n966_));
  INV_X1     g0830(.I(new_n952_), .ZN(new_n967_));
  NOR4_X1    g0831(.A1(new_n967_), .A2(new_n957_), .A3(new_n525_), .A4(new_n955_), .ZN(new_n968_));
  NOR4_X1    g0832(.A1(new_n966_), .A2(new_n968_), .A3(new_n537_), .A4(new_n953_), .ZN(new_n969_));
  NOR2_X1    g0833(.A1(new_n969_), .A2(new_n961_), .ZN(new_n970_));
  NOR2_X1    g0834(.A1(new_n968_), .A2(new_n953_), .ZN(new_n971_));
  NOR4_X1    g0835(.A1(new_n971_), .A2(new_n537_), .A3(new_n548_), .A4(new_n958_), .ZN(new_n972_));
  INV_X1     g0836(.I(new_n972_), .ZN(new_n973_));
  NAND4_X1   g0837(.A1(new_n963_), .A2(new_n971_), .A3(new_n962_), .A4(new_n549_), .ZN(new_n974_));
  NAND4_X1   g0838(.A1(new_n973_), .A2(new_n974_), .A3(new_n561_), .A4(new_n970_), .ZN(new_n975_));
  NAND2_X1   g0839(.A1(new_n975_), .A2(new_n965_), .ZN(new_n976_));
  NAND2_X1   g0840(.A1(new_n973_), .A2(new_n974_), .ZN(new_n977_));
  NAND4_X1   g0841(.A1(new_n977_), .A2(new_n561_), .A3(new_n573_), .A4(new_n964_), .ZN(new_n978_));
  NOR4_X1    g0842(.A1(new_n969_), .A2(new_n960_), .A3(new_n548_), .A4(new_n961_), .ZN(new_n979_));
  NOR2_X1    g0843(.A1(new_n979_), .A2(new_n972_), .ZN(new_n980_));
  NAND4_X1   g0844(.A1(new_n975_), .A2(new_n573_), .A3(new_n965_), .A4(new_n980_), .ZN(new_n981_));
  NAND2_X1   g0845(.A1(new_n981_), .A2(new_n978_), .ZN(new_n982_));
  NAND4_X1   g0846(.A1(new_n982_), .A2(new_n584_), .A3(new_n596_), .A4(new_n976_), .ZN(new_n983_));
  NOR4_X1    g0847(.A1(new_n980_), .A2(new_n560_), .A3(new_n572_), .A4(new_n970_), .ZN(new_n984_));
  NOR4_X1    g0848(.A1(new_n970_), .A2(new_n548_), .A3(new_n560_), .A4(new_n971_), .ZN(new_n985_));
  NOR4_X1    g0849(.A1(new_n979_), .A2(new_n964_), .A3(new_n560_), .A4(new_n972_), .ZN(new_n986_));
  NOR4_X1    g0850(.A1(new_n986_), .A2(new_n977_), .A3(new_n572_), .A4(new_n985_), .ZN(new_n987_));
  NOR2_X1    g0851(.A1(new_n987_), .A2(new_n984_), .ZN(new_n988_));
  NAND4_X1   g0852(.A1(new_n976_), .A2(new_n573_), .A3(new_n584_), .A4(new_n977_), .ZN(new_n989_));
  NOR2_X1    g0853(.A1(new_n986_), .A2(new_n985_), .ZN(new_n990_));
  NAND4_X1   g0854(.A1(new_n981_), .A2(new_n584_), .A3(new_n978_), .A4(new_n990_), .ZN(new_n991_));
  NAND4_X1   g0855(.A1(new_n991_), .A2(new_n988_), .A3(new_n989_), .A4(new_n596_), .ZN(new_n992_));
  NAND2_X1   g0856(.A1(new_n992_), .A2(new_n983_), .ZN(new_n993_));
  NAND2_X1   g0857(.A1(new_n991_), .A2(new_n989_), .ZN(new_n994_));
  NAND4_X1   g0858(.A1(new_n994_), .A2(new_n596_), .A3(new_n608_), .A4(new_n982_), .ZN(new_n995_));
  NOR4_X1    g0859(.A1(new_n990_), .A2(new_n572_), .A3(new_n583_), .A4(new_n980_), .ZN(new_n996_));
  NOR4_X1    g0860(.A1(new_n987_), .A2(new_n583_), .A3(new_n976_), .A4(new_n984_), .ZN(new_n997_));
  NOR2_X1    g0861(.A1(new_n997_), .A2(new_n996_), .ZN(new_n998_));
  NAND4_X1   g0862(.A1(new_n992_), .A2(new_n998_), .A3(new_n983_), .A4(new_n608_), .ZN(new_n999_));
  NAND2_X1   g0863(.A1(new_n999_), .A2(new_n995_), .ZN(new_n1000_));
  NAND4_X1   g0864(.A1(new_n1000_), .A2(new_n619_), .A3(new_n631_), .A4(new_n993_), .ZN(new_n1001_));
  NOR4_X1    g0865(.A1(new_n998_), .A2(new_n595_), .A3(new_n607_), .A4(new_n988_), .ZN(new_n1002_));
  NOR4_X1    g0866(.A1(new_n988_), .A2(new_n583_), .A3(new_n595_), .A4(new_n990_), .ZN(new_n1003_));
  NOR4_X1    g0867(.A1(new_n997_), .A2(new_n595_), .A3(new_n982_), .A4(new_n996_), .ZN(new_n1004_));
  NOR4_X1    g0868(.A1(new_n1004_), .A2(new_n607_), .A3(new_n994_), .A4(new_n1003_), .ZN(new_n1005_));
  NOR2_X1    g0869(.A1(new_n1005_), .A2(new_n1002_), .ZN(new_n1006_));
  NAND4_X1   g0870(.A1(new_n993_), .A2(new_n608_), .A3(new_n619_), .A4(new_n994_), .ZN(new_n1007_));
  NOR2_X1    g0871(.A1(new_n1004_), .A2(new_n1003_), .ZN(new_n1008_));
  NAND4_X1   g0872(.A1(new_n999_), .A2(new_n1008_), .A3(new_n995_), .A4(new_n619_), .ZN(new_n1009_));
  NAND4_X1   g0873(.A1(new_n1009_), .A2(new_n1006_), .A3(new_n1007_), .A4(new_n631_), .ZN(new_n1010_));
  NAND2_X1   g0874(.A1(new_n1010_), .A2(new_n1001_), .ZN(new_n1011_));
  NAND2_X1   g0875(.A1(new_n1009_), .A2(new_n1007_), .ZN(new_n1012_));
  NAND4_X1   g0876(.A1(new_n1012_), .A2(new_n631_), .A3(new_n643_), .A4(new_n1000_), .ZN(new_n1013_));
  NOR4_X1    g0877(.A1(new_n1008_), .A2(new_n607_), .A3(new_n618_), .A4(new_n998_), .ZN(new_n1014_));
  NOR4_X1    g0878(.A1(new_n1005_), .A2(new_n618_), .A3(new_n993_), .A4(new_n1002_), .ZN(new_n1015_));
  NOR2_X1    g0879(.A1(new_n1015_), .A2(new_n1014_), .ZN(new_n1016_));
  NAND4_X1   g0880(.A1(new_n1010_), .A2(new_n1016_), .A3(new_n1001_), .A4(new_n643_), .ZN(new_n1017_));
  NAND2_X1   g0881(.A1(new_n1017_), .A2(new_n1013_), .ZN(new_n1018_));
  NAND4_X1   g0882(.A1(new_n1018_), .A2(new_n654_), .A3(new_n666_), .A4(new_n1011_), .ZN(new_n1019_));
  NOR4_X1    g0883(.A1(new_n1016_), .A2(new_n630_), .A3(new_n642_), .A4(new_n1006_), .ZN(new_n1020_));
  NOR4_X1    g0884(.A1(new_n1006_), .A2(new_n618_), .A3(new_n630_), .A4(new_n1008_), .ZN(new_n1021_));
  NOR4_X1    g0885(.A1(new_n1015_), .A2(new_n630_), .A3(new_n1000_), .A4(new_n1014_), .ZN(new_n1022_));
  NOR4_X1    g0886(.A1(new_n1022_), .A2(new_n642_), .A3(new_n1012_), .A4(new_n1021_), .ZN(new_n1023_));
  NOR2_X1    g0887(.A1(new_n1023_), .A2(new_n1020_), .ZN(new_n1024_));
  NAND4_X1   g0888(.A1(new_n1011_), .A2(new_n643_), .A3(new_n654_), .A4(new_n1012_), .ZN(new_n1025_));
  NOR2_X1    g0889(.A1(new_n1022_), .A2(new_n1021_), .ZN(new_n1026_));
  NAND4_X1   g0890(.A1(new_n1017_), .A2(new_n1026_), .A3(new_n654_), .A4(new_n1013_), .ZN(new_n1027_));
  NAND4_X1   g0891(.A1(new_n1027_), .A2(new_n1024_), .A3(new_n666_), .A4(new_n1025_), .ZN(new_n1028_));
  NAND2_X1   g0892(.A1(new_n1028_), .A2(new_n1019_), .ZN(new_n1029_));
  NAND2_X1   g0893(.A1(new_n1027_), .A2(new_n1025_), .ZN(new_n1030_));
  NAND4_X1   g0894(.A1(new_n1030_), .A2(new_n666_), .A3(new_n678_), .A4(new_n1018_), .ZN(new_n1031_));
  NOR4_X1    g0895(.A1(new_n1026_), .A2(new_n642_), .A3(new_n653_), .A4(new_n1016_), .ZN(new_n1032_));
  NOR4_X1    g0896(.A1(new_n1023_), .A2(new_n653_), .A3(new_n1011_), .A4(new_n1020_), .ZN(new_n1033_));
  NOR2_X1    g0897(.A1(new_n1033_), .A2(new_n1032_), .ZN(new_n1034_));
  NAND4_X1   g0898(.A1(new_n1028_), .A2(new_n1034_), .A3(new_n678_), .A4(new_n1019_), .ZN(new_n1035_));
  NAND2_X1   g0899(.A1(new_n1035_), .A2(new_n1031_), .ZN(new_n1036_));
  NAND4_X1   g0900(.A1(new_n1036_), .A2(new_n689_), .A3(new_n701_), .A4(new_n1029_), .ZN(new_n1037_));
  NOR4_X1    g0901(.A1(new_n1034_), .A2(new_n665_), .A3(new_n677_), .A4(new_n1024_), .ZN(new_n1038_));
  NOR4_X1    g0902(.A1(new_n1024_), .A2(new_n653_), .A3(new_n665_), .A4(new_n1026_), .ZN(new_n1039_));
  NOR4_X1    g0903(.A1(new_n1033_), .A2(new_n665_), .A3(new_n1018_), .A4(new_n1032_), .ZN(new_n1040_));
  NOR4_X1    g0904(.A1(new_n1040_), .A2(new_n677_), .A3(new_n1030_), .A4(new_n1039_), .ZN(new_n1041_));
  NOR2_X1    g0905(.A1(new_n1041_), .A2(new_n1038_), .ZN(new_n1042_));
  NAND4_X1   g0906(.A1(new_n1029_), .A2(new_n678_), .A3(new_n689_), .A4(new_n1030_), .ZN(new_n1043_));
  NOR2_X1    g0907(.A1(new_n1040_), .A2(new_n1039_), .ZN(new_n1044_));
  NAND4_X1   g0908(.A1(new_n1035_), .A2(new_n1044_), .A3(new_n689_), .A4(new_n1031_), .ZN(new_n1045_));
  NAND4_X1   g0909(.A1(new_n1045_), .A2(new_n1042_), .A3(new_n701_), .A4(new_n1043_), .ZN(new_n1046_));
  NAND2_X1   g0910(.A1(new_n1046_), .A2(new_n1037_), .ZN(new_n1047_));
  NAND2_X1   g0911(.A1(new_n1045_), .A2(new_n1043_), .ZN(new_n1048_));
  NAND4_X1   g0912(.A1(new_n1048_), .A2(new_n701_), .A3(new_n713_), .A4(new_n1036_), .ZN(new_n1049_));
  NOR4_X1    g0913(.A1(new_n1044_), .A2(new_n677_), .A3(new_n688_), .A4(new_n1034_), .ZN(new_n1050_));
  NOR4_X1    g0914(.A1(new_n1041_), .A2(new_n688_), .A3(new_n1029_), .A4(new_n1038_), .ZN(new_n1051_));
  NOR2_X1    g0915(.A1(new_n1051_), .A2(new_n1050_), .ZN(new_n1052_));
  NAND4_X1   g0916(.A1(new_n1046_), .A2(new_n1052_), .A3(new_n713_), .A4(new_n1037_), .ZN(new_n1053_));
  NAND2_X1   g0917(.A1(new_n1053_), .A2(new_n1049_), .ZN(new_n1054_));
  NAND4_X1   g0918(.A1(new_n1054_), .A2(new_n724_), .A3(new_n736_), .A4(new_n1047_), .ZN(new_n1055_));
  NOR4_X1    g0919(.A1(new_n1052_), .A2(new_n700_), .A3(new_n712_), .A4(new_n1042_), .ZN(new_n1056_));
  NOR4_X1    g0920(.A1(new_n1042_), .A2(new_n688_), .A3(new_n700_), .A4(new_n1044_), .ZN(new_n1057_));
  NOR4_X1    g0921(.A1(new_n1051_), .A2(new_n700_), .A3(new_n1036_), .A4(new_n1050_), .ZN(new_n1058_));
  NOR4_X1    g0922(.A1(new_n1058_), .A2(new_n712_), .A3(new_n1048_), .A4(new_n1057_), .ZN(new_n1059_));
  NOR2_X1    g0923(.A1(new_n1059_), .A2(new_n1056_), .ZN(new_n1060_));
  NAND4_X1   g0924(.A1(new_n1047_), .A2(new_n713_), .A3(new_n724_), .A4(new_n1048_), .ZN(new_n1061_));
  NOR2_X1    g0925(.A1(new_n1058_), .A2(new_n1057_), .ZN(new_n1062_));
  NAND4_X1   g0926(.A1(new_n1053_), .A2(new_n1062_), .A3(new_n724_), .A4(new_n1049_), .ZN(new_n1063_));
  NAND4_X1   g0927(.A1(new_n1063_), .A2(new_n1060_), .A3(new_n736_), .A4(new_n1061_), .ZN(new_n1064_));
  NAND2_X1   g0928(.A1(new_n1064_), .A2(new_n1055_), .ZN(new_n1065_));
  NAND2_X1   g0929(.A1(new_n1063_), .A2(new_n1061_), .ZN(new_n1066_));
  NAND4_X1   g0930(.A1(new_n1066_), .A2(new_n736_), .A3(new_n748_), .A4(new_n1054_), .ZN(new_n1067_));
  NOR4_X1    g0931(.A1(new_n1062_), .A2(new_n712_), .A3(new_n723_), .A4(new_n1052_), .ZN(new_n1068_));
  NOR4_X1    g0932(.A1(new_n1059_), .A2(new_n723_), .A3(new_n1047_), .A4(new_n1056_), .ZN(new_n1069_));
  NOR2_X1    g0933(.A1(new_n1069_), .A2(new_n1068_), .ZN(new_n1070_));
  NAND4_X1   g0934(.A1(new_n1064_), .A2(new_n1070_), .A3(new_n748_), .A4(new_n1055_), .ZN(new_n1071_));
  NAND2_X1   g0935(.A1(new_n1071_), .A2(new_n1067_), .ZN(new_n1072_));
  NAND4_X1   g0936(.A1(new_n1072_), .A2(new_n759_), .A3(new_n771_), .A4(new_n1065_), .ZN(new_n1073_));
  NOR4_X1    g0937(.A1(new_n1070_), .A2(new_n735_), .A3(new_n747_), .A4(new_n1060_), .ZN(new_n1074_));
  NOR4_X1    g0938(.A1(new_n1060_), .A2(new_n723_), .A3(new_n735_), .A4(new_n1062_), .ZN(new_n1075_));
  NOR4_X1    g0939(.A1(new_n1069_), .A2(new_n735_), .A3(new_n1054_), .A4(new_n1068_), .ZN(new_n1076_));
  NOR4_X1    g0940(.A1(new_n1076_), .A2(new_n747_), .A3(new_n1066_), .A4(new_n1075_), .ZN(new_n1077_));
  NOR2_X1    g0941(.A1(new_n1077_), .A2(new_n1074_), .ZN(new_n1078_));
  NAND4_X1   g0942(.A1(new_n1065_), .A2(new_n748_), .A3(new_n759_), .A4(new_n1066_), .ZN(new_n1079_));
  NOR2_X1    g0943(.A1(new_n1076_), .A2(new_n1075_), .ZN(new_n1080_));
  NAND4_X1   g0944(.A1(new_n1071_), .A2(new_n1080_), .A3(new_n759_), .A4(new_n1067_), .ZN(new_n1081_));
  NAND4_X1   g0945(.A1(new_n1081_), .A2(new_n1078_), .A3(new_n771_), .A4(new_n1079_), .ZN(new_n1082_));
  NAND2_X1   g0946(.A1(new_n1082_), .A2(new_n1073_), .ZN(new_n1083_));
  NAND2_X1   g0947(.A1(new_n1081_), .A2(new_n1079_), .ZN(new_n1084_));
  NAND4_X1   g0948(.A1(new_n1084_), .A2(new_n771_), .A3(new_n783_), .A4(new_n1072_), .ZN(new_n1085_));
  NOR4_X1    g0949(.A1(new_n1080_), .A2(new_n747_), .A3(new_n758_), .A4(new_n1070_), .ZN(new_n1086_));
  NOR4_X1    g0950(.A1(new_n1077_), .A2(new_n758_), .A3(new_n1065_), .A4(new_n1074_), .ZN(new_n1087_));
  NOR2_X1    g0951(.A1(new_n1087_), .A2(new_n1086_), .ZN(new_n1088_));
  NAND4_X1   g0952(.A1(new_n1082_), .A2(new_n1088_), .A3(new_n783_), .A4(new_n1073_), .ZN(new_n1089_));
  NAND2_X1   g0953(.A1(new_n1089_), .A2(new_n1085_), .ZN(new_n1090_));
  NAND4_X1   g0954(.A1(new_n1090_), .A2(new_n793_), .A3(new_n804_), .A4(new_n1083_), .ZN(new_n1091_));
  INV_X1     g0955(.I(new_n1090_), .ZN(new_n1092_));
  NAND4_X1   g0956(.A1(new_n1083_), .A2(new_n783_), .A3(new_n793_), .A4(new_n1084_), .ZN(new_n1093_));
  INV_X1     g0957(.I(new_n1073_), .ZN(new_n1094_));
  NOR4_X1    g0958(.A1(new_n1087_), .A2(new_n770_), .A3(new_n1072_), .A4(new_n1086_), .ZN(new_n1095_));
  NOR2_X1    g0959(.A1(new_n1095_), .A2(new_n1094_), .ZN(new_n1096_));
  NAND4_X1   g0960(.A1(new_n1096_), .A2(new_n1089_), .A3(new_n793_), .A4(new_n1085_), .ZN(new_n1097_));
  NAND4_X1   g0961(.A1(new_n1092_), .A2(new_n804_), .A3(new_n1097_), .A4(new_n1093_), .ZN(new_n1098_));
  NAND2_X1   g0962(.A1(new_n1098_), .A2(new_n1091_), .ZN(new_n1099_));
  NOR2_X1    g0963(.A1(\A[10] ), .A2(\A[11] ), .ZN(new_n1100_));
  NAND2_X1   g0964(.A1(new_n1097_), .A2(new_n1093_), .ZN(new_n1101_));
  NAND2_X1   g0965(.A1(new_n1101_), .A2(new_n1100_), .ZN(new_n1102_));
  OAI21_X1   g0966(.A1(new_n1099_), .A2(new_n1100_), .B(new_n1102_), .ZN(new_n1103_));
  NAND4_X1   g0967(.A1(new_n1099_), .A2(new_n823_), .A3(new_n1101_), .A4(new_n1100_), .ZN(new_n1104_));
  INV_X1     g0968(.I(new_n1091_), .ZN(new_n1105_));
  NOR3_X1    g0969(.A1(new_n1101_), .A2(new_n803_), .A3(new_n1090_), .ZN(new_n1106_));
  NOR2_X1    g0970(.A1(new_n1106_), .A2(new_n1105_), .ZN(new_n1107_));
  NAND4_X1   g0971(.A1(new_n1107_), .A2(new_n823_), .A3(new_n1100_), .A4(new_n1102_), .ZN(new_n1108_));
  NAND2_X1   g0972(.A1(new_n1108_), .A2(new_n1104_), .ZN(new_n1109_));
  NOR4_X1    g0973(.A1(\A[2] ), .A2(\A[3] ), .A3(\A[4] ), .A4(\A[5] ), .ZN(new_n1110_));
  NAND4_X1   g0974(.A1(new_n1109_), .A2(new_n821_), .A3(new_n1103_), .A4(new_n1110_), .ZN(new_n1111_));
  INV_X1     g0975(.I(new_n1104_), .ZN(new_n1112_));
  INV_X1     g0976(.I(new_n823_), .ZN(new_n1113_));
  INV_X1     g0977(.I(new_n1100_), .ZN(new_n1114_));
  NOR4_X1    g0978(.A1(new_n1099_), .A2(new_n1113_), .A3(new_n1101_), .A4(new_n1114_), .ZN(new_n1115_));
  NOR2_X1    g0979(.A1(new_n1112_), .A2(new_n1115_), .ZN(new_n1116_));
  NAND4_X1   g0980(.A1(new_n1103_), .A2(new_n821_), .A3(new_n823_), .A4(new_n1099_), .ZN(new_n1117_));
  INV_X1     g0981(.I(new_n1102_), .ZN(new_n1118_));
  AOI21_X1   g0982(.A1(new_n1107_), .A2(new_n1114_), .B(new_n1118_), .ZN(new_n1119_));
  NAND4_X1   g0983(.A1(new_n1108_), .A2(new_n1119_), .A3(new_n1104_), .A4(new_n821_), .ZN(new_n1120_));
  NAND4_X1   g0984(.A1(new_n1120_), .A2(new_n1116_), .A3(new_n1110_), .A4(new_n1117_), .ZN(new_n1121_));
  NAND2_X1   g0985(.A1(new_n1121_), .A2(new_n1111_), .ZN(\P[1] ));
  NOR2_X1    g0986(.A1(new_n677_), .A2(new_n688_), .ZN(new_n1123_));
  NOR2_X1    g0987(.A1(new_n313_), .A2(new_n324_), .ZN(new_n1124_));
  INV_X1     g0988(.I(new_n1124_), .ZN(new_n1125_));
  NAND3_X1   g0989(.A1(new_n856_), .A2(new_n182_), .A3(new_n160_), .ZN(new_n1126_));
  NOR2_X1    g0990(.A1(new_n195_), .A2(new_n214_), .ZN(new_n1127_));
  INV_X1     g0991(.I(new_n1127_), .ZN(new_n1128_));
  NOR2_X1    g0992(.A1(new_n1128_), .A2(new_n158_), .ZN(new_n1129_));
  NOR3_X1    g0993(.A1(\A[112] ), .A2(\A[113] ), .A3(\A[114] ), .ZN(new_n1130_));
  OAI21_X1   g0994(.A1(new_n1129_), .A2(new_n1126_), .B(new_n1130_), .ZN(new_n1131_));
  NOR2_X1    g0995(.A1(new_n865_), .A2(new_n857_), .ZN(new_n1132_));
  INV_X1     g0996(.I(new_n1126_), .ZN(new_n1133_));
  NAND2_X1   g0997(.A1(new_n1128_), .A2(new_n1133_), .ZN(new_n1134_));
  NAND3_X1   g0998(.A1(new_n1134_), .A2(new_n1130_), .A3(new_n1132_), .ZN(new_n1135_));
  XNOR2_X1   g0999(.A1(new_n1135_), .A2(new_n1131_), .ZN(new_n1136_));
  NOR2_X1    g1000(.A1(new_n275_), .A2(new_n285_), .ZN(new_n1137_));
  INV_X1     g1001(.I(new_n1137_), .ZN(new_n1138_));
  NOR2_X1    g1002(.A1(new_n1136_), .A2(new_n1138_), .ZN(new_n1139_));
  NAND2_X1   g1003(.A1(new_n1134_), .A2(new_n1132_), .ZN(new_n1140_));
  NOR2_X1    g1004(.A1(new_n253_), .A2(new_n266_), .ZN(new_n1141_));
  INV_X1     g1005(.I(new_n1141_), .ZN(new_n1142_));
  NAND2_X1   g1006(.A1(new_n1136_), .A2(new_n1142_), .ZN(new_n1143_));
  OAI21_X1   g1007(.A1(new_n1140_), .A2(new_n1142_), .B(new_n1143_), .ZN(new_n1144_));
  NOR2_X1    g1008(.A1(new_n1144_), .A2(new_n1137_), .ZN(new_n1145_));
  NOR2_X1    g1009(.A1(new_n1145_), .A2(new_n1139_), .ZN(new_n1146_));
  NOR3_X1    g1010(.A1(new_n1146_), .A2(new_n313_), .A3(new_n324_), .ZN(new_n1147_));
  NOR3_X1    g1011(.A1(new_n891_), .A2(\A[100] ), .A3(\A[101] ), .ZN(new_n1148_));
  NAND2_X1   g1012(.A1(new_n1144_), .A2(new_n1148_), .ZN(new_n1149_));
  INV_X1     g1013(.I(new_n1149_), .ZN(new_n1150_));
  NOR3_X1    g1014(.A1(new_n1145_), .A2(new_n1139_), .A3(new_n1148_), .ZN(new_n1151_));
  NOR2_X1    g1015(.A1(new_n1151_), .A2(new_n1150_), .ZN(new_n1152_));
  AOI21_X1   g1016(.A1(new_n1152_), .A2(new_n1125_), .B(new_n1147_), .ZN(new_n1153_));
  NOR2_X1    g1017(.A1(new_n357_), .A2(new_n368_), .ZN(new_n1154_));
  INV_X1     g1018(.I(new_n1154_), .ZN(new_n1155_));
  NOR2_X1    g1019(.A1(new_n1153_), .A2(new_n1155_), .ZN(new_n1156_));
  NOR2_X1    g1020(.A1(new_n335_), .A2(new_n347_), .ZN(new_n1157_));
  INV_X1     g1021(.I(new_n1157_), .ZN(new_n1158_));
  NAND2_X1   g1022(.A1(new_n1153_), .A2(new_n1158_), .ZN(new_n1159_));
  OAI21_X1   g1023(.A1(new_n1152_), .A2(new_n1158_), .B(new_n1159_), .ZN(new_n1160_));
  NOR2_X1    g1024(.A1(new_n1160_), .A2(new_n1154_), .ZN(new_n1161_));
  NOR2_X1    g1025(.A1(new_n1161_), .A2(new_n1156_), .ZN(new_n1162_));
  NOR2_X1    g1026(.A1(new_n403_), .A2(new_n412_), .ZN(new_n1163_));
  INV_X1     g1027(.I(new_n1163_), .ZN(new_n1164_));
  NOR2_X1    g1028(.A1(new_n1162_), .A2(new_n1164_), .ZN(new_n1165_));
  NOR2_X1    g1029(.A1(new_n377_), .A2(new_n390_), .ZN(new_n1166_));
  NAND2_X1   g1030(.A1(new_n1160_), .A2(new_n1166_), .ZN(new_n1167_));
  INV_X1     g1031(.I(new_n1166_), .ZN(new_n1168_));
  NAND2_X1   g1032(.A1(new_n1162_), .A2(new_n1168_), .ZN(new_n1169_));
  NAND2_X1   g1033(.A1(new_n1169_), .A2(new_n1167_), .ZN(new_n1170_));
  NOR2_X1    g1034(.A1(new_n1170_), .A2(new_n1163_), .ZN(new_n1171_));
  NOR2_X1    g1035(.A1(new_n1171_), .A2(new_n1165_), .ZN(new_n1172_));
  NOR2_X1    g1036(.A1(new_n443_), .A2(new_n455_), .ZN(new_n1173_));
  INV_X1     g1037(.I(new_n1173_), .ZN(new_n1174_));
  NOR2_X1    g1038(.A1(new_n1172_), .A2(new_n1174_), .ZN(new_n1175_));
  NOR2_X1    g1039(.A1(new_n855_), .A2(new_n927_), .ZN(new_n1176_));
  NAND2_X1   g1040(.A1(new_n1170_), .A2(new_n1176_), .ZN(new_n1177_));
  INV_X1     g1041(.I(new_n1176_), .ZN(new_n1178_));
  NAND2_X1   g1042(.A1(new_n1172_), .A2(new_n1178_), .ZN(new_n1179_));
  NAND2_X1   g1043(.A1(new_n1179_), .A2(new_n1177_), .ZN(new_n1180_));
  NOR2_X1    g1044(.A1(new_n1180_), .A2(new_n1173_), .ZN(new_n1181_));
  NOR2_X1    g1045(.A1(new_n1181_), .A2(new_n1175_), .ZN(new_n1182_));
  NOR2_X1    g1046(.A1(new_n490_), .A2(new_n502_), .ZN(new_n1183_));
  INV_X1     g1047(.I(new_n1183_), .ZN(new_n1184_));
  NOR2_X1    g1048(.A1(new_n1182_), .A2(new_n1184_), .ZN(new_n1185_));
  NOR2_X1    g1049(.A1(new_n467_), .A2(new_n478_), .ZN(new_n1186_));
  NAND2_X1   g1050(.A1(new_n1180_), .A2(new_n1186_), .ZN(new_n1187_));
  INV_X1     g1051(.I(new_n1186_), .ZN(new_n1188_));
  NAND2_X1   g1052(.A1(new_n1182_), .A2(new_n1188_), .ZN(new_n1189_));
  NAND2_X1   g1053(.A1(new_n1189_), .A2(new_n1187_), .ZN(new_n1190_));
  NOR2_X1    g1054(.A1(new_n1190_), .A2(new_n1183_), .ZN(new_n1191_));
  NOR2_X1    g1055(.A1(new_n1191_), .A2(new_n1185_), .ZN(new_n1192_));
  NOR2_X1    g1056(.A1(new_n537_), .A2(new_n548_), .ZN(new_n1193_));
  INV_X1     g1057(.I(new_n1193_), .ZN(new_n1194_));
  NOR2_X1    g1058(.A1(new_n1192_), .A2(new_n1194_), .ZN(new_n1195_));
  NOR2_X1    g1059(.A1(new_n513_), .A2(new_n525_), .ZN(new_n1196_));
  NAND2_X1   g1060(.A1(new_n1190_), .A2(new_n1196_), .ZN(new_n1197_));
  INV_X1     g1061(.I(new_n1196_), .ZN(new_n1198_));
  NAND2_X1   g1062(.A1(new_n1192_), .A2(new_n1198_), .ZN(new_n1199_));
  NAND2_X1   g1063(.A1(new_n1199_), .A2(new_n1197_), .ZN(new_n1200_));
  NOR2_X1    g1064(.A1(new_n1200_), .A2(new_n1193_), .ZN(new_n1201_));
  NOR2_X1    g1065(.A1(new_n583_), .A2(new_n595_), .ZN(new_n1202_));
  OAI21_X1   g1066(.A1(new_n1201_), .A2(new_n1195_), .B(new_n1202_), .ZN(new_n1203_));
  NOR2_X1    g1067(.A1(new_n560_), .A2(new_n572_), .ZN(new_n1204_));
  NAND2_X1   g1068(.A1(new_n1200_), .A2(new_n1204_), .ZN(new_n1205_));
  OR3_X2     g1069(.A1(new_n1201_), .A2(new_n1195_), .A3(new_n1204_), .Z(new_n1206_));
  NAND2_X1   g1070(.A1(new_n1206_), .A2(new_n1205_), .ZN(new_n1207_));
  OR2_X2     g1071(.A1(new_n1207_), .A2(new_n1202_), .Z(new_n1208_));
  NAND2_X1   g1072(.A1(new_n1208_), .A2(new_n1203_), .ZN(new_n1209_));
  NOR2_X1    g1073(.A1(new_n630_), .A2(new_n642_), .ZN(new_n1210_));
  NAND2_X1   g1074(.A1(new_n1209_), .A2(new_n1210_), .ZN(new_n1211_));
  INV_X1     g1075(.I(new_n1210_), .ZN(new_n1212_));
  NOR2_X1    g1076(.A1(new_n607_), .A2(new_n618_), .ZN(new_n1213_));
  NAND2_X1   g1077(.A1(new_n1207_), .A2(new_n1213_), .ZN(new_n1214_));
  INV_X1     g1078(.I(new_n1213_), .ZN(new_n1215_));
  NAND3_X1   g1079(.A1(new_n1208_), .A2(new_n1203_), .A3(new_n1215_), .ZN(new_n1216_));
  NAND3_X1   g1080(.A1(new_n1216_), .A2(new_n1212_), .A3(new_n1214_), .ZN(new_n1217_));
  NAND2_X1   g1081(.A1(new_n1217_), .A2(new_n1211_), .ZN(new_n1218_));
  NAND2_X1   g1082(.A1(new_n1218_), .A2(new_n1123_), .ZN(new_n1219_));
  NAND2_X1   g1083(.A1(new_n1216_), .A2(new_n1214_), .ZN(new_n1220_));
  NOR2_X1    g1084(.A1(new_n653_), .A2(new_n665_), .ZN(new_n1221_));
  NAND2_X1   g1085(.A1(new_n1220_), .A2(new_n1221_), .ZN(new_n1222_));
  INV_X1     g1086(.I(new_n1221_), .ZN(new_n1223_));
  NAND3_X1   g1087(.A1(new_n1217_), .A2(new_n1211_), .A3(new_n1223_), .ZN(new_n1224_));
  NAND2_X1   g1088(.A1(new_n1224_), .A2(new_n1222_), .ZN(new_n1225_));
  OAI21_X1   g1089(.A1(new_n1225_), .A2(new_n1123_), .B(new_n1219_), .ZN(new_n1226_));
  NOR2_X1    g1090(.A1(new_n723_), .A2(new_n735_), .ZN(new_n1227_));
  NOR2_X1    g1091(.A1(new_n700_), .A2(new_n712_), .ZN(new_n1228_));
  NAND2_X1   g1092(.A1(new_n1225_), .A2(new_n1228_), .ZN(new_n1229_));
  OAI21_X1   g1093(.A1(new_n1226_), .A2(new_n1228_), .B(new_n1229_), .ZN(new_n1230_));
  NOR2_X1    g1094(.A1(new_n1230_), .A2(new_n1227_), .ZN(new_n1231_));
  AOI21_X1   g1095(.A1(new_n1226_), .A2(new_n1227_), .B(new_n1231_), .ZN(new_n1232_));
  NOR2_X1    g1096(.A1(new_n770_), .A2(new_n782_), .ZN(new_n1233_));
  INV_X1     g1097(.I(new_n1233_), .ZN(new_n1234_));
  NOR2_X1    g1098(.A1(new_n747_), .A2(new_n758_), .ZN(new_n1235_));
  INV_X1     g1099(.I(new_n1235_), .ZN(new_n1236_));
  AND2_X2    g1100(.A1(new_n1230_), .A2(new_n1235_), .Z(new_n1237_));
  AOI21_X1   g1101(.A1(new_n1232_), .A2(new_n1236_), .B(new_n1237_), .ZN(new_n1238_));
  NAND2_X1   g1102(.A1(new_n1238_), .A2(new_n1234_), .ZN(new_n1239_));
  OAI21_X1   g1103(.A1(new_n1232_), .A2(new_n1234_), .B(new_n1239_), .ZN(new_n1240_));
  NOR4_X1    g1104(.A1(\A[4] ), .A2(\A[5] ), .A3(\A[6] ), .A4(\A[7] ), .ZN(new_n1241_));
  NOR3_X1    g1105(.A1(new_n1114_), .A2(\A[8] ), .A3(\A[9] ), .ZN(new_n1242_));
  NAND2_X1   g1106(.A1(new_n1242_), .A2(new_n1241_), .ZN(new_n1243_));
  NOR2_X1    g1107(.A1(new_n1240_), .A2(new_n1243_), .ZN(new_n1244_));
  NOR2_X1    g1108(.A1(new_n792_), .A2(new_n803_), .ZN(new_n1245_));
  MUX2_X1    g1109(.I0(new_n1240_), .I1(new_n1238_), .S(new_n1245_), .Z(new_n1246_));
  NOR2_X1    g1110(.A1(new_n1246_), .A2(new_n1243_), .ZN(new_n1247_));
  XOR2_X1    g1111(.A1(new_n1247_), .A2(new_n1244_), .Z(\P[2] ));
  INV_X1     g1112(.I(new_n1123_), .ZN(new_n1249_));
  NOR2_X1    g1113(.A1(new_n1249_), .A2(new_n1223_), .ZN(new_n1250_));
  INV_X1     g1114(.I(new_n1250_), .ZN(new_n1251_));
  NAND2_X1   g1115(.A1(new_n1202_), .A2(new_n1204_), .ZN(new_n1252_));
  NOR2_X1    g1116(.A1(new_n1184_), .A2(new_n1188_), .ZN(new_n1253_));
  INV_X1     g1117(.I(new_n1253_), .ZN(new_n1254_));
  NOR2_X1    g1118(.A1(new_n1164_), .A2(new_n1168_), .ZN(new_n1255_));
  INV_X1     g1119(.I(new_n1255_), .ZN(new_n1256_));
  NOR3_X1    g1120(.A1(new_n1128_), .A2(new_n225_), .A3(new_n239_), .ZN(new_n1257_));
  NOR2_X1    g1121(.A1(new_n1138_), .A2(new_n1142_), .ZN(new_n1258_));
  NAND2_X1   g1122(.A1(new_n1258_), .A2(\A[103] ), .ZN(new_n1259_));
  NAND3_X1   g1123(.A1(new_n1124_), .A2(\A[102] ), .A3(new_n305_), .ZN(new_n1260_));
  AOI21_X1   g1124(.A1(new_n1259_), .A2(new_n1257_), .B(new_n1260_), .ZN(new_n1261_));
  NAND2_X1   g1125(.A1(new_n1133_), .A2(new_n1132_), .ZN(new_n1262_));
  INV_X1     g1126(.I(new_n1257_), .ZN(new_n1263_));
  INV_X1     g1127(.I(new_n1262_), .ZN(new_n1264_));
  OAI21_X1   g1128(.A1(new_n1263_), .A2(new_n1258_), .B(new_n1264_), .ZN(new_n1265_));
  NOR3_X1    g1129(.A1(new_n1265_), .A2(new_n1260_), .A3(new_n1262_), .ZN(new_n1266_));
  XNOR2_X1   g1130(.A1(new_n1266_), .A2(new_n1261_), .ZN(new_n1267_));
  NOR2_X1    g1131(.A1(new_n1267_), .A2(new_n1256_), .ZN(new_n1268_));
  NOR2_X1    g1132(.A1(new_n1155_), .A2(new_n1158_), .ZN(new_n1269_));
  INV_X1     g1133(.I(new_n1269_), .ZN(new_n1270_));
  NOR2_X1    g1134(.A1(new_n1265_), .A2(new_n1270_), .ZN(new_n1271_));
  AOI21_X1   g1135(.A1(new_n1267_), .A2(new_n1270_), .B(new_n1271_), .ZN(new_n1272_));
  AOI21_X1   g1136(.A1(new_n1272_), .A2(new_n1256_), .B(new_n1268_), .ZN(new_n1273_));
  NOR2_X1    g1137(.A1(new_n1273_), .A2(new_n1254_), .ZN(new_n1274_));
  NOR2_X1    g1138(.A1(new_n1178_), .A2(new_n1174_), .ZN(new_n1275_));
  INV_X1     g1139(.I(new_n1275_), .ZN(new_n1276_));
  NOR2_X1    g1140(.A1(new_n1272_), .A2(new_n1276_), .ZN(new_n1277_));
  AOI21_X1   g1141(.A1(new_n1273_), .A2(new_n1276_), .B(new_n1277_), .ZN(new_n1278_));
  AOI21_X1   g1142(.A1(new_n1278_), .A2(new_n1254_), .B(new_n1274_), .ZN(new_n1279_));
  NOR2_X1    g1143(.A1(new_n1279_), .A2(new_n1252_), .ZN(new_n1280_));
  NOR2_X1    g1144(.A1(new_n1194_), .A2(new_n1198_), .ZN(new_n1281_));
  INV_X1     g1145(.I(new_n1281_), .ZN(new_n1282_));
  NOR2_X1    g1146(.A1(new_n1278_), .A2(new_n1282_), .ZN(new_n1283_));
  AOI21_X1   g1147(.A1(new_n1279_), .A2(new_n1282_), .B(new_n1283_), .ZN(new_n1284_));
  AOI21_X1   g1148(.A1(new_n1284_), .A2(new_n1252_), .B(new_n1280_), .ZN(new_n1285_));
  NOR2_X1    g1149(.A1(new_n1285_), .A2(new_n1251_), .ZN(new_n1286_));
  NOR2_X1    g1150(.A1(new_n1212_), .A2(new_n1215_), .ZN(new_n1287_));
  INV_X1     g1151(.I(new_n1287_), .ZN(new_n1288_));
  NOR2_X1    g1152(.A1(new_n1284_), .A2(new_n1288_), .ZN(new_n1289_));
  AOI21_X1   g1153(.A1(new_n1285_), .A2(new_n1288_), .B(new_n1289_), .ZN(new_n1290_));
  AOI21_X1   g1154(.A1(new_n1290_), .A2(new_n1251_), .B(new_n1286_), .ZN(new_n1291_));
  NAND2_X1   g1155(.A1(new_n1242_), .A2(new_n1245_), .ZN(new_n1292_));
  NOR3_X1    g1156(.A1(new_n1292_), .A2(new_n1234_), .A3(new_n1236_), .ZN(new_n1293_));
  NAND2_X1   g1157(.A1(new_n1291_), .A2(new_n1293_), .ZN(new_n1294_));
  NAND2_X1   g1158(.A1(new_n1227_), .A2(new_n1228_), .ZN(new_n1295_));
  NOR2_X1    g1159(.A1(new_n1290_), .A2(new_n1295_), .ZN(new_n1296_));
  AND2_X2    g1160(.A1(new_n1291_), .A2(new_n1295_), .Z(new_n1297_));
  OAI21_X1   g1161(.A1(new_n1297_), .A2(new_n1296_), .B(new_n1293_), .ZN(new_n1298_));
  XOR2_X1    g1162(.A1(new_n1298_), .A2(new_n1294_), .Z(\P[3] ));
  NAND3_X1   g1163(.A1(new_n1258_), .A2(new_n1124_), .A3(new_n1148_), .ZN(new_n1300_));
  NOR2_X1    g1164(.A1(new_n1256_), .A2(new_n1270_), .ZN(new_n1301_));
  AOI21_X1   g1165(.A1(new_n1301_), .A2(\A[79] ), .B(new_n1300_), .ZN(new_n1302_));
  NAND4_X1   g1166(.A1(new_n1253_), .A2(\A[78] ), .A3(new_n854_), .A4(new_n1173_), .ZN(new_n1303_));
  NOR2_X1    g1167(.A1(new_n1302_), .A2(new_n1303_), .ZN(new_n1304_));
  NAND2_X1   g1168(.A1(new_n1264_), .A2(new_n1257_), .ZN(new_n1305_));
  NOR2_X1    g1169(.A1(new_n1301_), .A2(new_n1300_), .ZN(new_n1306_));
  NOR3_X1    g1170(.A1(new_n1306_), .A2(new_n1303_), .A3(new_n1305_), .ZN(new_n1307_));
  XNOR2_X1   g1171(.A1(new_n1307_), .A2(new_n1304_), .ZN(new_n1308_));
  NAND4_X1   g1172(.A1(new_n1227_), .A2(new_n1228_), .A3(new_n1233_), .A4(new_n1235_), .ZN(new_n1309_));
  NAND2_X1   g1173(.A1(new_n1250_), .A2(new_n1287_), .ZN(new_n1310_));
  NOR2_X1    g1174(.A1(new_n1310_), .A2(new_n1309_), .ZN(new_n1311_));
  NAND2_X1   g1175(.A1(new_n1308_), .A2(new_n1311_), .ZN(new_n1312_));
  NOR2_X1    g1176(.A1(new_n1282_), .A2(new_n1252_), .ZN(new_n1313_));
  INV_X1     g1177(.I(new_n1313_), .ZN(new_n1314_));
  NOR3_X1    g1178(.A1(new_n1306_), .A2(new_n1305_), .A3(new_n1314_), .ZN(new_n1315_));
  AND2_X2    g1179(.A1(new_n1308_), .A2(new_n1314_), .Z(new_n1316_));
  OAI21_X1   g1180(.A1(new_n1316_), .A2(new_n1315_), .B(new_n1311_), .ZN(new_n1317_));
  XOR2_X1    g1181(.A1(new_n1317_), .A2(new_n1312_), .Z(\P[4] ));
  NOR2_X1    g1182(.A1(new_n1305_), .A2(new_n1300_), .ZN(new_n1319_));
  NOR2_X1    g1183(.A1(new_n1314_), .A2(new_n1310_), .ZN(new_n1320_));
  NAND3_X1   g1184(.A1(new_n1301_), .A2(new_n1253_), .A3(new_n1275_), .ZN(new_n1321_));
  OAI21_X1   g1185(.A1(new_n1320_), .A2(new_n1321_), .B(new_n1319_), .ZN(\P[5] ));
  INV_X1     g1186(.I(new_n1321_), .ZN(new_n1323_));
  NAND2_X1   g1187(.A1(new_n1323_), .A2(new_n1319_), .ZN(\P[6] ));
  INV_X1     g1188(.I(new_n1241_), .ZN(new_n1325_));
  OR4_X2     g1189(.A1(\A[0] ), .A2(\A[1] ), .A3(\A[2] ), .A4(\A[3] ), .Z(new_n1326_));
  NOR4_X1    g1190(.A1(new_n1292_), .A2(new_n1309_), .A3(new_n1325_), .A4(new_n1326_), .ZN(new_n1327_));
  NAND4_X1   g1191(.A1(new_n1323_), .A2(new_n1319_), .A3(new_n1320_), .A4(new_n1327_), .ZN(F));
endmodule


