// Benchmark "c880.blif" written by ABC on Fri Feb 25 15:12:30 2022

module c880  ( 
    G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat,
    G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat,
    G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat,
    G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat,
    G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat,
    G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat,
    G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat,
    G267gat, G268gat,
    G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat,
    G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat,
    G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat,
    G879gat, G880gat  );
  input  G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat,
    G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat,
    G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat,
    G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat,
    G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat,
    G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat,
    G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat,
    G261gat, G267gat, G268gat;
  output G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat,
    G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat,
    G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat,
    G878gat, G879gat, G880gat;
  wire new_n87_, new_n89_, new_n93_, new_n94_, new_n96_, new_n97_, new_n99_,
    new_n101_, new_n104_, new_n108_, new_n109_, new_n110_, new_n112_,
    new_n113_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_;
  assign new_n87_ = G29gat & G75gat;
  assign G388gat = G42gat & new_n87_;
  assign new_n89_ = G29gat & G36gat;
  assign G389gat = G80gat & new_n89_;
  assign G390gat = G42gat & new_n89_;
  assign G391gat = G85gat & G86gat;
  assign new_n93_ = G13gat & G17gat;
  assign new_n94_ = G1gat & G8gat;
  assign G418gat = new_n93_ & new_n94_;
  assign new_n96_ = G1gat & G26gat;
  assign new_n97_ = new_n93_ & new_n96_;
  assign G419gat = G390gat | ~new_n97_;
  assign new_n99_ = G59gat & G75gat;
  assign G420gat = ~G80gat | ~new_n99_;
  assign new_n101_ = G36gat & G59gat;
  assign G421gat = ~G80gat | ~new_n101_;
  assign G422gat = ~G42gat | ~new_n101_;
  assign new_n104_ = ~G87gat & ~G88gat;
  assign G423gat = G90gat & ~new_n104_;
  assign G446gat = ~G390gat | ~new_n97_;
  assign G447gat = G51gat & new_n96_;
  assign new_n108_ = G13gat & G55gat;
  assign new_n109_ = new_n94_ & new_n108_;
  assign new_n110_ = G29gat & G68gat;
  assign G448gat = new_n109_ & new_n110_;
  assign new_n112_ = G59gat & G68gat;
  assign new_n113_ = G74gat & new_n112_;
  assign G449gat = new_n109_ & new_n113_;
  assign G450gat = G89gat & ~new_n104_;
  assign new_n116_ = G91gat & G96gat;
  assign new_n117_ = ~G91gat & ~G96gat;
  assign new_n118_ = ~new_n116_ & ~new_n117_;
  assign new_n119_ = G101gat & G106gat;
  assign new_n120_ = ~G101gat & ~G106gat;
  assign new_n121_ = ~new_n119_ & ~new_n120_;
  assign new_n122_ = ~new_n118_ & ~new_n121_;
  assign new_n123_ = new_n118_ & new_n121_;
  assign new_n124_ = ~new_n122_ & ~new_n123_;
  assign new_n125_ = G130gat & new_n124_;
  assign new_n126_ = ~G130gat & ~new_n124_;
  assign new_n127_ = ~new_n125_ & ~new_n126_;
  assign new_n128_ = G111gat & G116gat;
  assign new_n129_ = ~G111gat & ~G116gat;
  assign new_n130_ = ~new_n128_ & ~new_n129_;
  assign new_n131_ = G121gat & G126gat;
  assign new_n132_ = ~G121gat & ~G126gat;
  assign new_n133_ = ~new_n131_ & ~new_n132_;
  assign new_n134_ = ~new_n130_ & ~new_n133_;
  assign new_n135_ = new_n130_ & new_n133_;
  assign new_n136_ = ~new_n134_ & ~new_n135_;
  assign new_n137_ = G135gat & new_n136_;
  assign new_n138_ = ~G135gat & ~new_n136_;
  assign new_n139_ = ~new_n137_ & ~new_n138_;
  assign new_n140_ = ~new_n127_ & ~new_n139_;
  assign new_n141_ = new_n127_ & new_n139_;
  assign G767gat = ~new_n140_ & ~new_n141_;
  assign new_n143_ = G159gat & G165gat;
  assign new_n144_ = ~G159gat & ~G165gat;
  assign new_n145_ = ~new_n143_ & ~new_n144_;
  assign new_n146_ = G171gat & G177gat;
  assign new_n147_ = ~G171gat & ~G177gat;
  assign new_n148_ = ~new_n146_ & ~new_n147_;
  assign new_n149_ = ~new_n145_ & ~new_n148_;
  assign new_n150_ = new_n145_ & new_n148_;
  assign new_n151_ = ~new_n149_ & ~new_n150_;
  assign new_n152_ = G130gat & new_n151_;
  assign new_n153_ = ~G130gat & ~new_n151_;
  assign new_n154_ = ~new_n152_ & ~new_n153_;
  assign new_n155_ = G183gat & G189gat;
  assign new_n156_ = ~G183gat & ~G189gat;
  assign new_n157_ = ~new_n155_ & ~new_n156_;
  assign new_n158_ = G195gat & G201gat;
  assign new_n159_ = ~G195gat & ~G201gat;
  assign new_n160_ = ~new_n158_ & ~new_n159_;
  assign new_n161_ = ~new_n157_ & ~new_n160_;
  assign new_n162_ = new_n157_ & new_n160_;
  assign new_n163_ = ~new_n161_ & ~new_n162_;
  assign new_n164_ = G207gat & new_n163_;
  assign new_n165_ = ~G207gat & ~new_n163_;
  assign new_n166_ = ~new_n164_ & ~new_n165_;
  assign new_n167_ = ~new_n154_ & ~new_n166_;
  assign new_n168_ = new_n154_ & new_n166_;
  assign G768gat = ~new_n167_ & ~new_n168_;
  assign new_n170_ = G121gat & G210gat;
  assign new_n171_ = G80gat & new_n87_;
  assign new_n172_ = G447gat & new_n171_;
  assign new_n173_ = G55gat & new_n172_;
  assign new_n174_ = ~G268gat & new_n173_;
  assign new_n175_ = G59gat & G156gat;
  assign new_n176_ = G447gat & ~new_n175_;
  assign new_n177_ = G17gat & new_n176_;
  assign new_n178_ = G1gat & ~new_n177_;
  assign new_n179_ = G153gat & ~new_n178_;
  assign new_n180_ = ~G17gat & ~G42gat;
  assign new_n181_ = G17gat & G42gat;
  assign new_n182_ = ~new_n180_ & ~new_n181_;
  assign new_n183_ = G156gat & G447gat;
  assign new_n184_ = G59gat & new_n182_;
  assign new_n185_ = new_n183_ & new_n184_;
  assign new_n186_ = G17gat & G51gat;
  assign new_n187_ = new_n94_ & new_n186_;
  assign new_n188_ = G42gat & new_n99_;
  assign new_n189_ = new_n187_ & ~new_n188_;
  assign new_n190_ = ~new_n185_ & ~new_n189_;
  assign new_n191_ = G126gat & ~new_n190_;
  assign new_n192_ = ~new_n179_ & ~new_n191_;
  assign new_n193_ = ~new_n174_ & new_n192_;
  assign new_n194_ = ~G201gat & new_n193_;
  assign new_n195_ = G201gat & ~new_n193_;
  assign new_n196_ = ~new_n194_ & ~new_n195_;
  assign new_n197_ = ~G261gat & ~new_n196_;
  assign new_n198_ = G261gat & new_n196_;
  assign new_n199_ = ~new_n197_ & ~new_n198_;
  assign new_n200_ = G219gat & new_n199_;
  assign new_n201_ = ~new_n170_ & ~new_n200_;
  assign new_n202_ = G228gat & new_n196_;
  assign new_n203_ = G237gat & new_n195_;
  assign new_n204_ = ~new_n202_ & ~new_n203_;
  assign new_n205_ = G255gat & G267gat;
  assign new_n206_ = G246gat & ~new_n193_;
  assign new_n207_ = ~new_n205_ & ~new_n206_;
  assign new_n208_ = G68gat & G72gat;
  assign new_n209_ = G42gat & G59gat;
  assign new_n210_ = new_n208_ & new_n209_;
  assign new_n211_ = new_n109_ & new_n210_;
  assign new_n212_ = G73gat & new_n211_;
  assign new_n213_ = G201gat & new_n212_;
  assign new_n214_ = new_n207_ & ~new_n213_;
  assign new_n215_ = new_n201_ & new_n204_;
  assign G850gat = ~new_n214_ | ~new_n215_;
  assign new_n217_ = G106gat & G210gat;
  assign new_n218_ = G143gat & ~new_n178_;
  assign new_n219_ = G111gat & ~new_n190_;
  assign new_n220_ = ~new_n218_ & ~new_n219_;
  assign new_n221_ = ~new_n174_ & new_n220_;
  assign new_n222_ = ~G183gat & new_n221_;
  assign new_n223_ = G183gat & ~new_n221_;
  assign new_n224_ = ~new_n222_ & ~new_n223_;
  assign new_n225_ = G146gat & ~new_n178_;
  assign new_n226_ = G116gat & ~new_n190_;
  assign new_n227_ = ~new_n225_ & ~new_n226_;
  assign new_n228_ = ~new_n174_ & new_n227_;
  assign new_n229_ = G189gat & ~new_n228_;
  assign new_n230_ = ~G189gat & new_n228_;
  assign new_n231_ = G149gat & ~new_n178_;
  assign new_n232_ = G121gat & ~new_n190_;
  assign new_n233_ = ~new_n231_ & ~new_n232_;
  assign new_n234_ = ~new_n174_ & new_n233_;
  assign new_n235_ = G195gat & ~new_n234_;
  assign new_n236_ = ~new_n230_ & new_n235_;
  assign new_n237_ = ~G195gat & new_n234_;
  assign new_n238_ = ~new_n230_ & ~new_n237_;
  assign new_n239_ = new_n195_ & new_n238_;
  assign new_n240_ = G261gat & ~new_n194_;
  assign new_n241_ = new_n238_ & new_n240_;
  assign new_n242_ = ~new_n239_ & ~new_n241_;
  assign new_n243_ = ~new_n229_ & ~new_n236_;
  assign new_n244_ = new_n242_ & new_n243_;
  assign new_n245_ = ~new_n224_ & new_n244_;
  assign new_n246_ = new_n224_ & ~new_n244_;
  assign new_n247_ = ~new_n245_ & ~new_n246_;
  assign new_n248_ = G219gat & new_n247_;
  assign new_n249_ = ~new_n217_ & ~new_n248_;
  assign new_n250_ = G228gat & new_n224_;
  assign new_n251_ = G237gat & new_n223_;
  assign new_n252_ = ~new_n250_ & ~new_n251_;
  assign new_n253_ = G246gat & ~new_n221_;
  assign new_n254_ = G183gat & new_n212_;
  assign new_n255_ = ~new_n253_ & ~new_n254_;
  assign new_n256_ = new_n249_ & new_n252_;
  assign G863gat = ~new_n255_ | ~new_n256_;
  assign new_n258_ = G111gat & G210gat;
  assign new_n259_ = ~new_n229_ & ~new_n230_;
  assign new_n260_ = new_n195_ & ~new_n237_;
  assign new_n261_ = ~new_n194_ & ~new_n237_;
  assign new_n262_ = G261gat & new_n261_;
  assign new_n263_ = ~new_n235_ & ~new_n260_;
  assign new_n264_ = ~new_n262_ & new_n263_;
  assign new_n265_ = ~new_n259_ & new_n264_;
  assign new_n266_ = new_n259_ & ~new_n264_;
  assign new_n267_ = ~new_n265_ & ~new_n266_;
  assign new_n268_ = G219gat & new_n267_;
  assign new_n269_ = ~new_n258_ & ~new_n268_;
  assign new_n270_ = G228gat & new_n259_;
  assign new_n271_ = G237gat & new_n229_;
  assign new_n272_ = ~new_n270_ & ~new_n271_;
  assign new_n273_ = G255gat & G259gat;
  assign new_n274_ = G246gat & ~new_n228_;
  assign new_n275_ = ~new_n273_ & ~new_n274_;
  assign new_n276_ = G189gat & new_n212_;
  assign new_n277_ = new_n275_ & ~new_n276_;
  assign new_n278_ = new_n269_ & new_n272_;
  assign G864gat = ~new_n277_ | ~new_n278_;
  assign new_n280_ = G116gat & G210gat;
  assign new_n281_ = ~new_n235_ & ~new_n237_;
  assign new_n282_ = ~new_n195_ & ~new_n240_;
  assign new_n283_ = ~new_n281_ & new_n282_;
  assign new_n284_ = new_n281_ & ~new_n282_;
  assign new_n285_ = ~new_n283_ & ~new_n284_;
  assign new_n286_ = G219gat & new_n285_;
  assign new_n287_ = ~new_n280_ & ~new_n286_;
  assign new_n288_ = G228gat & new_n281_;
  assign new_n289_ = G237gat & new_n235_;
  assign new_n290_ = ~new_n288_ & ~new_n289_;
  assign new_n291_ = G255gat & G260gat;
  assign new_n292_ = G246gat & ~new_n234_;
  assign new_n293_ = ~new_n291_ & ~new_n292_;
  assign new_n294_ = G195gat & new_n212_;
  assign new_n295_ = new_n293_ & ~new_n294_;
  assign new_n296_ = new_n287_ & new_n290_;
  assign G865gat = ~new_n295_ | ~new_n296_;
  assign new_n298_ = G8gat & G138gat;
  assign new_n299_ = G91gat & ~new_n190_;
  assign new_n300_ = ~new_n298_ & ~new_n299_;
  assign new_n301_ = G55gat & new_n176_;
  assign new_n302_ = G143gat & new_n301_;
  assign new_n303_ = G17gat & G447gat;
  assign new_n304_ = new_n171_ & new_n303_;
  assign new_n305_ = ~G268gat & new_n304_;
  assign new_n306_ = ~new_n302_ & ~new_n305_;
  assign new_n307_ = new_n300_ & new_n306_;
  assign new_n308_ = G159gat & ~new_n307_;
  assign new_n309_ = G51gat & G138gat;
  assign new_n310_ = G96gat & ~new_n190_;
  assign new_n311_ = ~new_n309_ & ~new_n310_;
  assign new_n312_ = G146gat & new_n301_;
  assign new_n313_ = ~new_n305_ & ~new_n312_;
  assign new_n314_ = new_n311_ & new_n313_;
  assign new_n315_ = G165gat & ~new_n314_;
  assign new_n316_ = ~G165gat & new_n314_;
  assign new_n317_ = G17gat & G138gat;
  assign new_n318_ = G101gat & ~new_n190_;
  assign new_n319_ = ~new_n317_ & ~new_n318_;
  assign new_n320_ = G149gat & new_n301_;
  assign new_n321_ = ~new_n305_ & ~new_n320_;
  assign new_n322_ = new_n319_ & new_n321_;
  assign new_n323_ = G171gat & ~new_n322_;
  assign new_n324_ = ~new_n316_ & new_n323_;
  assign new_n325_ = ~G171gat & new_n322_;
  assign new_n326_ = G138gat & G152gat;
  assign new_n327_ = G106gat & ~new_n190_;
  assign new_n328_ = ~new_n326_ & ~new_n327_;
  assign new_n329_ = G153gat & new_n301_;
  assign new_n330_ = ~new_n305_ & ~new_n329_;
  assign new_n331_ = new_n328_ & new_n330_;
  assign new_n332_ = G177gat & ~new_n331_;
  assign new_n333_ = ~new_n316_ & ~new_n325_;
  assign new_n334_ = new_n332_ & new_n333_;
  assign new_n335_ = ~G177gat & new_n331_;
  assign new_n336_ = ~new_n222_ & ~new_n244_;
  assign new_n337_ = ~new_n223_ & ~new_n336_;
  assign new_n338_ = ~new_n335_ & ~new_n337_;
  assign new_n339_ = new_n333_ & new_n338_;
  assign new_n340_ = ~new_n334_ & ~new_n339_;
  assign new_n341_ = ~new_n315_ & ~new_n324_;
  assign new_n342_ = new_n340_ & new_n341_;
  assign new_n343_ = ~G159gat & new_n307_;
  assign new_n344_ = ~new_n342_ & ~new_n343_;
  assign G866gat = new_n308_ | new_n344_;
  assign new_n346_ = G101gat & G210gat;
  assign new_n347_ = ~new_n332_ & ~new_n335_;
  assign new_n348_ = new_n337_ & ~new_n347_;
  assign new_n349_ = ~new_n337_ & new_n347_;
  assign new_n350_ = ~new_n348_ & ~new_n349_;
  assign new_n351_ = G219gat & new_n350_;
  assign new_n352_ = ~new_n346_ & ~new_n351_;
  assign new_n353_ = G228gat & new_n347_;
  assign new_n354_ = G237gat & new_n332_;
  assign new_n355_ = ~new_n353_ & ~new_n354_;
  assign new_n356_ = G246gat & ~new_n331_;
  assign new_n357_ = G177gat & new_n212_;
  assign new_n358_ = ~new_n356_ & ~new_n357_;
  assign new_n359_ = new_n352_ & new_n355_;
  assign G874gat = ~new_n358_ | ~new_n359_;
  assign new_n361_ = G210gat & G268gat;
  assign new_n362_ = ~new_n308_ & ~new_n343_;
  assign new_n363_ = new_n342_ & ~new_n362_;
  assign new_n364_ = ~new_n342_ & new_n362_;
  assign new_n365_ = ~new_n363_ & ~new_n364_;
  assign new_n366_ = G219gat & new_n365_;
  assign new_n367_ = ~new_n361_ & ~new_n366_;
  assign new_n368_ = G228gat & new_n362_;
  assign new_n369_ = G237gat & new_n308_;
  assign new_n370_ = ~new_n368_ & ~new_n369_;
  assign new_n371_ = G246gat & ~new_n307_;
  assign new_n372_ = G159gat & new_n212_;
  assign new_n373_ = ~new_n371_ & ~new_n372_;
  assign new_n374_ = new_n367_ & new_n370_;
  assign G878gat = ~new_n373_ | ~new_n374_;
  assign new_n376_ = G91gat & G210gat;
  assign new_n377_ = ~new_n315_ & ~new_n316_;
  assign new_n378_ = ~new_n325_ & new_n332_;
  assign new_n379_ = ~new_n325_ & ~new_n335_;
  assign new_n380_ = ~new_n337_ & new_n379_;
  assign new_n381_ = ~new_n323_ & ~new_n378_;
  assign new_n382_ = ~new_n380_ & new_n381_;
  assign new_n383_ = ~new_n377_ & new_n382_;
  assign new_n384_ = new_n377_ & ~new_n382_;
  assign new_n385_ = ~new_n383_ & ~new_n384_;
  assign new_n386_ = G219gat & new_n385_;
  assign new_n387_ = ~new_n376_ & ~new_n386_;
  assign new_n388_ = G228gat & new_n377_;
  assign new_n389_ = G237gat & new_n315_;
  assign new_n390_ = ~new_n388_ & ~new_n389_;
  assign new_n391_ = G246gat & ~new_n314_;
  assign new_n392_ = G165gat & new_n212_;
  assign new_n393_ = ~new_n391_ & ~new_n392_;
  assign new_n394_ = new_n387_ & new_n390_;
  assign G879gat = ~new_n393_ | ~new_n394_;
  assign new_n396_ = G96gat & G210gat;
  assign new_n397_ = ~new_n323_ & ~new_n325_;
  assign new_n398_ = ~new_n332_ & ~new_n338_;
  assign new_n399_ = ~new_n397_ & new_n398_;
  assign new_n400_ = new_n397_ & ~new_n398_;
  assign new_n401_ = ~new_n399_ & ~new_n400_;
  assign new_n402_ = G219gat & new_n401_;
  assign new_n403_ = ~new_n396_ & ~new_n402_;
  assign new_n404_ = G228gat & new_n397_;
  assign new_n405_ = G237gat & new_n323_;
  assign new_n406_ = ~new_n404_ & ~new_n405_;
  assign new_n407_ = G246gat & ~new_n322_;
  assign new_n408_ = G171gat & new_n212_;
  assign new_n409_ = ~new_n407_ & ~new_n408_;
  assign new_n410_ = new_n403_ & new_n406_;
  assign G880gat = ~new_n409_ | ~new_n410_;
endmodule


