// Benchmark "i2c" written by ABC on Fri Sep 15 11:25:53 2023

module i2c ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n475_, new_n476_,
    new_n477_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n485_, new_n486_, new_n487_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n507_, new_n508_, new_n509_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n518_,
    new_n519_, new_n521_, new_n522_, new_n523_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n541_, new_n542_, new_n543_, new_n544_, new_n546_,
    new_n547_, new_n548_, new_n550_, new_n551_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n869_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n963_, new_n964_, new_n966_,
    new_n967_, new_n969_, new_n970_, new_n972_, new_n973_, new_n974_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_, new_n986_, new_n987_, new_n989_, new_n990_,
    new_n992_, new_n993_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1010_, new_n1011_,
    new_n1013_, new_n1014_, new_n1016_, new_n1017_, new_n1019_, new_n1020_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1027_, new_n1028_,
    new_n1030_, new_n1031_, new_n1033_, new_n1034_, new_n1036_, new_n1037_,
    new_n1039_, new_n1040_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1053_,
    new_n1055_, new_n1057_, new_n1058_, new_n1060_, new_n1061_, new_n1063_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1114_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1139_, new_n1140_, new_n1142_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1149_, new_n1150_, new_n1152_, new_n1153_, new_n1155_,
    new_n1156_, new_n1158_, new_n1161_, new_n1162_, new_n1165_, new_n1171_,
    new_n1173_;
  NOR2_X1    g000(.A1(pi003), .A2(pi129), .ZN(new_n291_));
  INV_X1     g001(.I(pi054), .ZN(new_n292_));
  INV_X1     g002(.I(pi056), .ZN(new_n293_));
  NOR2_X1    g003(.A1(pi005), .A2(pi022), .ZN(new_n294_));
  NOR3_X1    g004(.A1(new_n294_), .A2(pi009), .A3(pi011), .ZN(new_n295_));
  INV_X1     g005(.I(new_n294_), .ZN(new_n296_));
  NOR2_X1    g006(.A1(pi009), .A2(pi011), .ZN(new_n297_));
  NOR2_X1    g007(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OAI21_X1   g008(.A1(new_n298_), .A2(new_n295_), .B(new_n293_), .ZN(new_n299_));
  INV_X1     g009(.I(pi007), .ZN(new_n300_));
  INV_X1     g010(.I(pi008), .ZN(new_n301_));
  INV_X1     g011(.I(pi021), .ZN(new_n302_));
  NAND3_X1   g012(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  NOR3_X1    g013(.A1(new_n303_), .A2(pi013), .A3(pi014), .ZN(new_n304_));
  NAND2_X1   g014(.A1(new_n304_), .A2(pi010), .ZN(new_n305_));
  INV_X1     g015(.I(pi010), .ZN(new_n306_));
  OAI21_X1   g016(.A1(pi008), .A2(pi021), .B(pi013), .ZN(new_n307_));
  INV_X1     g017(.I(pi013), .ZN(new_n308_));
  NOR2_X1    g018(.A1(pi008), .A2(pi021), .ZN(new_n309_));
  NAND2_X1   g019(.A1(new_n309_), .A2(new_n308_), .ZN(new_n310_));
  NAND2_X1   g020(.A1(pi008), .A2(pi021), .ZN(new_n311_));
  NAND4_X1   g021(.A1(new_n310_), .A2(new_n300_), .A3(new_n307_), .A4(new_n311_), .ZN(new_n312_));
  NAND3_X1   g022(.A1(new_n309_), .A2(pi007), .A3(new_n308_), .ZN(new_n313_));
  AOI21_X1   g023(.A1(new_n312_), .A2(new_n313_), .B(pi014), .ZN(new_n314_));
  INV_X1     g024(.I(pi014), .ZN(new_n315_));
  NOR3_X1    g025(.A1(new_n303_), .A2(pi013), .A3(new_n315_), .ZN(new_n316_));
  OAI21_X1   g026(.A1(new_n314_), .A2(new_n316_), .B(new_n306_), .ZN(new_n317_));
  NAND2_X1   g027(.A1(new_n317_), .A2(new_n305_), .ZN(new_n318_));
  INV_X1     g028(.I(pi006), .ZN(new_n319_));
  INV_X1     g029(.I(pi012), .ZN(new_n320_));
  NAND2_X1   g030(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1     g031(.I(pi018), .ZN(new_n322_));
  NOR2_X1    g032(.A1(pi004), .A2(pi019), .ZN(new_n323_));
  NAND2_X1   g033(.A1(new_n323_), .A2(new_n322_), .ZN(new_n324_));
  NOR2_X1    g034(.A1(new_n324_), .A2(pi016), .ZN(new_n325_));
  INV_X1     g035(.I(new_n325_), .ZN(new_n326_));
  NOR4_X1    g036(.A1(new_n326_), .A2(pi017), .A3(new_n296_), .A4(new_n321_), .ZN(new_n327_));
  NAND3_X1   g037(.A1(new_n318_), .A2(new_n297_), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1   g038(.A1(new_n328_), .A2(new_n299_), .B(new_n292_), .ZN(new_n329_));
  NOR3_X1    g039(.A1(new_n296_), .A2(pi013), .A3(pi014), .ZN(new_n330_));
  NOR3_X1    g040(.A1(pi008), .A2(pi017), .A3(pi021), .ZN(new_n331_));
  NAND2_X1   g041(.A1(new_n331_), .A2(new_n300_), .ZN(new_n332_));
  NOR2_X1    g042(.A1(new_n332_), .A2(new_n321_), .ZN(new_n333_));
  NAND4_X1   g043(.A1(new_n333_), .A2(new_n325_), .A3(new_n330_), .A4(new_n297_), .ZN(new_n334_));
  AOI21_X1   g044(.A1(new_n334_), .A2(pi054), .B(pi000), .ZN(new_n335_));
  OAI21_X1   g045(.A1(new_n329_), .A2(new_n335_), .B(new_n291_), .ZN(po015));
  NAND2_X1   g046(.A1(new_n300_), .A2(new_n308_), .ZN(new_n337_));
  NOR4_X1    g047(.A1(new_n337_), .A2(pi005), .A3(pi006), .A4(pi012), .ZN(new_n338_));
  NAND2_X1   g048(.A1(new_n338_), .A2(pi009), .ZN(new_n339_));
  INV_X1     g049(.I(pi009), .ZN(new_n340_));
  NAND2_X1   g050(.A1(new_n321_), .A2(pi007), .ZN(new_n341_));
  NAND3_X1   g051(.A1(new_n319_), .A2(new_n300_), .A3(new_n320_), .ZN(new_n342_));
  AOI21_X1   g052(.A1(pi006), .A2(pi012), .B(pi005), .ZN(new_n343_));
  NAND3_X1   g053(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND4_X1   g054(.A1(new_n319_), .A2(new_n300_), .A3(new_n320_), .A4(pi005), .ZN(new_n345_));
  AOI21_X1   g055(.A1(new_n344_), .A2(new_n345_), .B(pi013), .ZN(new_n346_));
  NOR4_X1    g056(.A1(pi005), .A2(pi006), .A3(pi007), .A4(pi012), .ZN(new_n347_));
  INV_X1     g057(.I(new_n347_), .ZN(new_n348_));
  NOR2_X1    g058(.A1(new_n348_), .A2(new_n308_), .ZN(new_n349_));
  OAI21_X1   g059(.A1(new_n346_), .A2(new_n349_), .B(new_n340_), .ZN(new_n350_));
  NOR2_X1    g060(.A1(pi010), .A2(pi022), .ZN(new_n351_));
  NAND2_X1   g061(.A1(new_n351_), .A2(new_n315_), .ZN(new_n352_));
  NOR2_X1    g062(.A1(new_n352_), .A2(new_n292_), .ZN(new_n353_));
  INV_X1     g063(.I(pi011), .ZN(new_n354_));
  NAND2_X1   g064(.A1(new_n331_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1     g065(.I(new_n355_), .ZN(new_n356_));
  NAND3_X1   g066(.A1(new_n325_), .A2(new_n356_), .A3(new_n353_), .ZN(new_n357_));
  AOI21_X1   g067(.A1(new_n350_), .A2(new_n339_), .B(new_n357_), .ZN(new_n358_));
  NOR4_X1    g068(.A1(pi005), .A2(pi006), .A3(pi007), .A4(pi013), .ZN(new_n359_));
  INV_X1     g069(.I(new_n309_), .ZN(new_n360_));
  NOR2_X1    g070(.A1(pi011), .A2(pi012), .ZN(new_n361_));
  INV_X1     g071(.I(new_n361_), .ZN(new_n362_));
  NOR4_X1    g072(.A1(new_n326_), .A2(new_n360_), .A3(new_n352_), .A4(new_n362_), .ZN(new_n363_));
  AOI21_X1   g073(.A1(new_n363_), .A2(new_n359_), .B(pi017), .ZN(new_n364_));
  AOI21_X1   g074(.A1(new_n364_), .A2(pi054), .B(pi001), .ZN(new_n365_));
  OAI21_X1   g075(.A1(new_n365_), .A2(new_n358_), .B(new_n291_), .ZN(po016));
  NAND2_X1   g076(.A1(pi122), .A2(pi127), .ZN(new_n367_));
  INV_X1     g077(.I(new_n367_), .ZN(new_n368_));
  INV_X1     g078(.I(pi082), .ZN(new_n369_));
  INV_X1     g079(.I(pi044), .ZN(new_n370_));
  NOR2_X1    g080(.A1(pi040), .A2(pi042), .ZN(new_n371_));
  NAND2_X1   g081(.A1(new_n371_), .A2(new_n370_), .ZN(new_n372_));
  INV_X1     g082(.I(new_n372_), .ZN(new_n373_));
  INV_X1     g083(.I(pi043), .ZN(new_n374_));
  INV_X1     g084(.I(pi047), .ZN(new_n375_));
  INV_X1     g085(.I(pi048), .ZN(new_n376_));
  NAND3_X1   g086(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1     g087(.I(pi002), .ZN(new_n378_));
  INV_X1     g088(.I(pi045), .ZN(new_n379_));
  NOR2_X1    g089(.A1(pi024), .A2(pi049), .ZN(new_n380_));
  INV_X1     g090(.I(new_n380_), .ZN(new_n381_));
  NOR3_X1    g091(.A1(new_n381_), .A2(pi015), .A3(pi020), .ZN(new_n382_));
  NAND3_X1   g092(.A1(new_n382_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n383_));
  INV_X1     g093(.I(pi041), .ZN(new_n384_));
  INV_X1     g094(.I(pi046), .ZN(new_n385_));
  NAND2_X1   g095(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1     g096(.I(pi038), .ZN(new_n387_));
  INV_X1     g097(.I(pi050), .ZN(new_n388_));
  NAND2_X1   g098(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR4_X1    g099(.A1(new_n383_), .A2(new_n377_), .A3(new_n386_), .A4(new_n389_), .ZN(new_n390_));
  AOI21_X1   g100(.A1(new_n390_), .A2(new_n373_), .B(new_n369_), .ZN(new_n391_));
  OR3_X2     g101(.A1(new_n391_), .A2(pi065), .A3(new_n368_), .Z(new_n392_));
  NOR2_X1    g102(.A1(new_n368_), .A2(pi082), .ZN(new_n393_));
  NOR2_X1    g103(.A1(pi047), .A2(pi048), .ZN(new_n394_));
  INV_X1     g104(.I(new_n394_), .ZN(new_n395_));
  INV_X1     g105(.I(pi024), .ZN(new_n396_));
  NOR3_X1    g106(.A1(pi015), .A2(pi020), .A3(pi049), .ZN(new_n397_));
  NAND3_X1   g107(.A1(new_n397_), .A2(new_n396_), .A3(new_n379_), .ZN(new_n398_));
  NAND3_X1   g108(.A1(new_n384_), .A2(new_n385_), .A3(new_n388_), .ZN(new_n399_));
  INV_X1     g109(.I(pi040), .ZN(new_n400_));
  NOR2_X1    g110(.A1(pi042), .A2(pi044), .ZN(new_n401_));
  NAND3_X1   g111(.A1(new_n401_), .A2(new_n387_), .A3(new_n400_), .ZN(new_n402_));
  NOR2_X1    g112(.A1(new_n402_), .A2(new_n399_), .ZN(new_n403_));
  NAND2_X1   g113(.A1(new_n403_), .A2(new_n374_), .ZN(new_n404_));
  NOR4_X1    g114(.A1(new_n404_), .A2(new_n369_), .A3(new_n395_), .A4(new_n398_), .ZN(new_n405_));
  OR3_X2     g115(.A1(new_n405_), .A2(new_n378_), .A3(new_n393_), .Z(new_n406_));
  AOI21_X1   g116(.A1(new_n392_), .A2(new_n406_), .B(pi129), .ZN(po017));
  INV_X1     g117(.I(pi113), .ZN(new_n408_));
  INV_X1     g118(.I(pi123), .ZN(new_n409_));
  NAND3_X1   g119(.A1(new_n408_), .A2(new_n409_), .A3(pi000), .ZN(new_n410_));
  INV_X1     g120(.I(new_n359_), .ZN(new_n411_));
  NAND3_X1   g121(.A1(new_n351_), .A2(new_n340_), .A3(new_n315_), .ZN(new_n412_));
  INV_X1     g122(.I(new_n412_), .ZN(new_n413_));
  NAND4_X1   g123(.A1(new_n325_), .A2(new_n413_), .A3(new_n331_), .A4(new_n361_), .ZN(new_n414_));
  NOR2_X1    g124(.A1(pi061), .A2(pi118), .ZN(new_n415_));
  OAI21_X1   g125(.A1(new_n414_), .A2(new_n411_), .B(new_n415_), .ZN(new_n416_));
  AOI21_X1   g126(.A1(new_n416_), .A2(new_n410_), .B(pi129), .ZN(po018));
  INV_X1     g127(.I(new_n291_), .ZN(new_n418_));
  NOR4_X1    g128(.A1(new_n306_), .A2(pi009), .A3(pi014), .A4(pi022), .ZN(new_n419_));
  NOR3_X1    g129(.A1(new_n326_), .A2(new_n292_), .A3(new_n355_), .ZN(new_n420_));
  NAND3_X1   g130(.A1(new_n420_), .A2(new_n338_), .A3(new_n419_), .ZN(new_n421_));
  NAND2_X1   g131(.A1(new_n292_), .A2(pi004), .ZN(new_n422_));
  AOI21_X1   g132(.A1(new_n421_), .A2(new_n422_), .B(new_n418_), .ZN(po019));
  NOR2_X1    g133(.A1(new_n292_), .A2(pi016), .ZN(new_n424_));
  NOR2_X1    g134(.A1(new_n412_), .A2(pi013), .ZN(new_n425_));
  INV_X1     g135(.I(new_n425_), .ZN(new_n426_));
  NOR3_X1    g136(.A1(new_n426_), .A2(pi059), .A3(new_n355_), .ZN(new_n427_));
  INV_X1     g137(.I(pi028), .ZN(new_n428_));
  NOR4_X1    g138(.A1(new_n324_), .A2(pi025), .A3(new_n428_), .A4(pi029), .ZN(new_n429_));
  NAND4_X1   g139(.A1(new_n427_), .A2(new_n347_), .A3(new_n424_), .A4(new_n429_), .ZN(new_n430_));
  NAND2_X1   g140(.A1(new_n292_), .A2(pi005), .ZN(new_n431_));
  AOI21_X1   g141(.A1(new_n430_), .A2(new_n431_), .B(new_n418_), .ZN(po020));
  INV_X1     g142(.I(pi025), .ZN(new_n433_));
  INV_X1     g143(.I(pi029), .ZN(new_n434_));
  INV_X1     g144(.I(new_n324_), .ZN(new_n435_));
  NAND3_X1   g145(.A1(new_n435_), .A2(new_n428_), .A3(new_n434_), .ZN(new_n436_));
  NOR2_X1    g146(.A1(new_n436_), .A2(new_n433_), .ZN(new_n437_));
  NAND4_X1   g147(.A1(new_n427_), .A2(new_n437_), .A3(new_n347_), .A4(new_n424_), .ZN(new_n438_));
  NAND2_X1   g148(.A1(new_n292_), .A2(pi006), .ZN(new_n439_));
  AOI21_X1   g149(.A1(new_n438_), .A2(new_n439_), .B(new_n418_), .ZN(po021));
  NOR4_X1    g150(.A1(new_n301_), .A2(pi005), .A3(pi007), .A4(pi017), .ZN(new_n441_));
  NAND2_X1   g151(.A1(new_n424_), .A2(new_n323_), .ZN(new_n442_));
  NOR3_X1    g152(.A1(new_n442_), .A2(pi006), .A3(new_n362_), .ZN(new_n443_));
  NOR2_X1    g153(.A1(pi018), .A2(pi021), .ZN(new_n444_));
  NAND4_X1   g154(.A1(new_n443_), .A2(new_n425_), .A3(new_n441_), .A4(new_n444_), .ZN(new_n445_));
  NAND2_X1   g155(.A1(new_n292_), .A2(pi007), .ZN(new_n446_));
  AOI21_X1   g156(.A1(new_n445_), .A2(new_n446_), .B(new_n418_), .ZN(po022));
  NAND2_X1   g157(.A1(new_n292_), .A2(pi008), .ZN(new_n448_));
  NAND2_X1   g158(.A1(new_n338_), .A2(new_n413_), .ZN(new_n449_));
  INV_X1     g159(.I(new_n449_), .ZN(new_n450_));
  NOR2_X1    g160(.A1(pi017), .A2(pi018), .ZN(new_n451_));
  NOR4_X1    g161(.A1(new_n442_), .A2(pi008), .A3(pi011), .A4(new_n302_), .ZN(new_n452_));
  NAND3_X1   g162(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1   g163(.A1(new_n453_), .A2(new_n448_), .B(new_n418_), .ZN(po023));
  INV_X1     g164(.I(new_n442_), .ZN(new_n455_));
  NAND2_X1   g165(.A1(new_n309_), .A2(new_n451_), .ZN(new_n456_));
  NOR2_X1    g166(.A1(new_n348_), .A2(new_n456_), .ZN(new_n457_));
  NOR4_X1    g167(.A1(new_n354_), .A2(pi009), .A3(pi013), .A4(pi014), .ZN(new_n458_));
  NAND4_X1   g168(.A1(new_n457_), .A2(new_n455_), .A3(new_n351_), .A4(new_n458_), .ZN(new_n459_));
  NAND2_X1   g169(.A1(new_n292_), .A2(pi009), .ZN(new_n460_));
  AOI21_X1   g170(.A1(new_n459_), .A2(new_n460_), .B(new_n418_), .ZN(po024));
  NOR4_X1    g171(.A1(new_n362_), .A2(pi005), .A3(pi006), .A4(pi007), .ZN(new_n462_));
  INV_X1     g172(.I(new_n424_), .ZN(new_n463_));
  NOR3_X1    g173(.A1(new_n463_), .A2(pi013), .A3(new_n315_), .ZN(new_n464_));
  NOR4_X1    g174(.A1(new_n456_), .A2(pi009), .A3(pi010), .A4(pi022), .ZN(new_n465_));
  NAND4_X1   g175(.A1(new_n464_), .A2(new_n465_), .A3(new_n323_), .A4(new_n462_), .ZN(new_n466_));
  NAND2_X1   g176(.A1(new_n292_), .A2(pi010), .ZN(new_n467_));
  AOI21_X1   g177(.A1(new_n466_), .A2(new_n467_), .B(new_n418_), .ZN(po025));
  INV_X1     g178(.I(pi022), .ZN(new_n469_));
  NOR4_X1    g179(.A1(new_n456_), .A2(pi010), .A3(pi011), .A4(new_n469_), .ZN(new_n470_));
  NOR3_X1    g180(.A1(new_n463_), .A2(pi009), .A3(pi014), .ZN(new_n471_));
  NAND4_X1   g181(.A1(new_n471_), .A2(new_n470_), .A3(new_n323_), .A4(new_n338_), .ZN(new_n472_));
  NAND2_X1   g182(.A1(new_n292_), .A2(pi011), .ZN(new_n473_));
  AOI21_X1   g183(.A1(new_n472_), .A2(new_n473_), .B(new_n418_), .ZN(po026));
  NOR3_X1    g184(.A1(new_n442_), .A2(new_n322_), .A3(new_n362_), .ZN(new_n475_));
  NAND4_X1   g185(.A1(new_n475_), .A2(new_n331_), .A3(new_n359_), .A4(new_n413_), .ZN(new_n476_));
  NAND2_X1   g186(.A1(new_n292_), .A2(pi012), .ZN(new_n477_));
  AOI21_X1   g187(.A1(new_n476_), .A2(new_n477_), .B(new_n418_), .ZN(po027));
  NOR2_X1    g188(.A1(new_n355_), .A2(pi059), .ZN(new_n479_));
  NOR3_X1    g189(.A1(new_n434_), .A2(pi025), .A3(pi028), .ZN(new_n480_));
  NOR2_X1    g190(.A1(new_n449_), .A2(new_n324_), .ZN(new_n481_));
  NAND4_X1   g191(.A1(new_n481_), .A2(new_n424_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n482_));
  NAND2_X1   g192(.A1(new_n292_), .A2(pi013), .ZN(new_n483_));
  AOI21_X1   g193(.A1(new_n482_), .A2(new_n483_), .B(new_n418_), .ZN(po028));
  NOR4_X1    g194(.A1(new_n456_), .A2(pi009), .A3(new_n308_), .A4(pi016), .ZN(new_n485_));
  NAND4_X1   g195(.A1(new_n485_), .A2(new_n323_), .A3(new_n462_), .A4(new_n353_), .ZN(new_n486_));
  NAND2_X1   g196(.A1(new_n292_), .A2(pi014), .ZN(new_n487_));
  AOI21_X1   g197(.A1(new_n486_), .A2(new_n487_), .B(new_n418_), .ZN(po029));
  INV_X1     g198(.I(pi070), .ZN(new_n489_));
  NOR3_X1    g199(.A1(pi038), .A2(pi046), .A3(pi050), .ZN(new_n490_));
  NOR2_X1    g200(.A1(pi041), .A2(pi043), .ZN(new_n491_));
  INV_X1     g201(.I(new_n491_), .ZN(new_n492_));
  NOR4_X1    g202(.A1(new_n395_), .A2(new_n492_), .A3(pi015), .A4(pi045), .ZN(new_n493_));
  NAND4_X1   g203(.A1(new_n493_), .A2(new_n373_), .A3(new_n380_), .A4(new_n490_), .ZN(new_n494_));
  AOI21_X1   g204(.A1(new_n494_), .A2(pi082), .B(new_n368_), .ZN(new_n495_));
  INV_X1     g205(.I(pi015), .ZN(new_n496_));
  NOR2_X1    g206(.A1(new_n367_), .A2(new_n496_), .ZN(new_n497_));
  AOI22_X1   g207(.A1(new_n495_), .A2(new_n489_), .B1(new_n369_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1     g208(.I(pi020), .ZN(new_n499_));
  NAND2_X1   g209(.A1(new_n378_), .A2(new_n499_), .ZN(new_n500_));
  NAND4_X1   g210(.A1(new_n500_), .A2(new_n496_), .A3(new_n379_), .A4(new_n380_), .ZN(new_n501_));
  NOR3_X1    g211(.A1(new_n404_), .A2(new_n395_), .A3(new_n501_), .ZN(new_n502_));
  NOR3_X1    g212(.A1(new_n377_), .A2(new_n381_), .A3(pi045), .ZN(new_n503_));
  AOI21_X1   g213(.A1(new_n503_), .A2(new_n403_), .B(new_n496_), .ZN(new_n504_));
  OAI21_X1   g214(.A1(new_n502_), .A2(new_n504_), .B(pi082), .ZN(new_n505_));
  AOI21_X1   g215(.A1(new_n498_), .A2(new_n505_), .B(pi129), .ZN(po030));
  NOR4_X1    g216(.A1(new_n337_), .A2(pi005), .A3(new_n319_), .A4(pi012), .ZN(new_n507_));
  NAND3_X1   g217(.A1(new_n420_), .A2(new_n413_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1   g218(.A1(new_n292_), .A2(pi016), .ZN(new_n509_));
  AOI21_X1   g219(.A1(new_n508_), .A2(new_n509_), .B(new_n418_), .ZN(po031));
  NOR4_X1    g220(.A1(new_n292_), .A2(pi005), .A3(pi006), .A4(pi017), .ZN(new_n511_));
  NOR4_X1    g221(.A1(pi007), .A2(pi012), .A3(pi016), .A4(pi025), .ZN(new_n512_));
  INV_X1     g222(.I(pi059), .ZN(new_n513_));
  NOR4_X1    g223(.A1(new_n436_), .A2(pi011), .A3(new_n513_), .A4(new_n360_), .ZN(new_n514_));
  NAND4_X1   g224(.A1(new_n514_), .A2(new_n425_), .A3(new_n511_), .A4(new_n512_), .ZN(new_n515_));
  NAND2_X1   g225(.A1(new_n292_), .A2(pi017), .ZN(new_n516_));
  AOI21_X1   g226(.A1(new_n515_), .A2(new_n516_), .B(new_n418_), .ZN(po032));
  NAND4_X1   g227(.A1(new_n481_), .A2(pi016), .A3(pi054), .A4(new_n356_), .ZN(new_n518_));
  NAND2_X1   g228(.A1(new_n292_), .A2(pi018), .ZN(new_n519_));
  AOI21_X1   g229(.A1(new_n518_), .A2(new_n519_), .B(new_n418_), .ZN(po033));
  NAND4_X1   g230(.A1(new_n435_), .A2(new_n354_), .A3(pi017), .A4(new_n424_), .ZN(new_n521_));
  OR3_X2     g231(.A1(new_n449_), .A2(new_n521_), .A3(new_n360_), .Z(new_n522_));
  NAND2_X1   g232(.A1(new_n292_), .A2(pi019), .ZN(new_n523_));
  AOI21_X1   g233(.A1(new_n522_), .A2(new_n523_), .B(new_n418_), .ZN(po034));
  INV_X1     g234(.I(pi071), .ZN(new_n525_));
  NOR3_X1    g235(.A1(new_n492_), .A2(pi046), .A3(pi047), .ZN(new_n526_));
  NOR3_X1    g236(.A1(pi024), .A2(pi045), .A3(pi048), .ZN(new_n527_));
  NOR2_X1    g237(.A1(new_n372_), .A2(new_n389_), .ZN(new_n528_));
  NAND4_X1   g238(.A1(new_n526_), .A2(new_n528_), .A3(new_n397_), .A4(new_n527_), .ZN(new_n529_));
  AOI21_X1   g239(.A1(new_n529_), .A2(pi082), .B(new_n368_), .ZN(new_n530_));
  NOR2_X1    g240(.A1(new_n367_), .A2(new_n499_), .ZN(new_n531_));
  AOI22_X1   g241(.A1(new_n530_), .A2(new_n525_), .B1(new_n369_), .B2(new_n531_), .ZN(new_n532_));
  NOR3_X1    g242(.A1(pi038), .A2(pi040), .A3(pi050), .ZN(new_n533_));
  INV_X1     g243(.I(new_n401_), .ZN(new_n534_));
  NAND2_X1   g244(.A1(new_n526_), .A2(new_n527_), .ZN(new_n535_));
  NOR4_X1    g245(.A1(new_n535_), .A2(pi015), .A3(pi049), .A4(new_n534_), .ZN(new_n536_));
  AOI21_X1   g246(.A1(new_n536_), .A2(new_n533_), .B(new_n499_), .ZN(new_n537_));
  NOR2_X1    g247(.A1(new_n529_), .A2(new_n378_), .ZN(new_n538_));
  OAI21_X1   g248(.A1(new_n537_), .A2(new_n538_), .B(pi082), .ZN(new_n539_));
  AOI21_X1   g249(.A1(new_n539_), .A2(new_n532_), .B(pi129), .ZN(po035));
  AND3_X2    g250(.A1(new_n302_), .A2(pi019), .A3(pi054), .Z(new_n541_));
  NOR4_X1    g251(.A1(pi004), .A2(pi008), .A3(pi011), .A4(pi016), .ZN(new_n542_));
  NAND4_X1   g252(.A1(new_n450_), .A2(new_n451_), .A3(new_n541_), .A4(new_n542_), .ZN(new_n543_));
  NAND2_X1   g253(.A1(new_n292_), .A2(pi021), .ZN(new_n544_));
  AOI21_X1   g254(.A1(new_n543_), .A2(new_n544_), .B(new_n418_), .ZN(po036));
  NOR2_X1    g255(.A1(new_n337_), .A2(pi014), .ZN(new_n546_));
  NAND4_X1   g256(.A1(new_n443_), .A2(new_n465_), .A3(pi005), .A4(new_n546_), .ZN(new_n547_));
  NAND2_X1   g257(.A1(new_n292_), .A2(pi022), .ZN(new_n548_));
  AOI21_X1   g258(.A1(new_n547_), .A2(new_n548_), .B(new_n418_), .ZN(po037));
  INV_X1     g259(.I(pi055), .ZN(new_n550_));
  OAI21_X1   g260(.A1(new_n550_), .A2(pi023), .B(pi061), .ZN(new_n551_));
  NOR2_X1    g261(.A1(new_n551_), .A2(pi129), .ZN(po038));
  INV_X1     g262(.I(pi063), .ZN(new_n553_));
  NOR3_X1    g263(.A1(new_n395_), .A2(pi002), .A3(pi045), .ZN(new_n554_));
  INV_X1     g264(.I(new_n397_), .ZN(new_n555_));
  NOR2_X1    g265(.A1(new_n404_), .A2(new_n555_), .ZN(new_n556_));
  AOI21_X1   g266(.A1(new_n556_), .A2(new_n554_), .B(new_n369_), .ZN(new_n557_));
  NOR3_X1    g267(.A1(new_n557_), .A2(new_n553_), .A3(new_n368_), .ZN(new_n558_));
  INV_X1     g268(.I(new_n533_), .ZN(new_n559_));
  NAND3_X1   g269(.A1(new_n526_), .A2(new_n379_), .A3(new_n376_), .ZN(new_n560_));
  NAND2_X1   g270(.A1(new_n401_), .A2(pi082), .ZN(new_n561_));
  NOR4_X1    g271(.A1(new_n560_), .A2(new_n396_), .A3(new_n559_), .A4(new_n561_), .ZN(new_n562_));
  NAND2_X1   g272(.A1(new_n373_), .A2(new_n490_), .ZN(new_n563_));
  NAND2_X1   g273(.A1(new_n491_), .A2(new_n375_), .ZN(new_n564_));
  OR4_X2     g274(.A1(pi045), .A2(new_n563_), .A3(pi048), .A4(new_n564_), .Z(new_n565_));
  INV_X1     g275(.I(pi049), .ZN(new_n566_));
  NOR3_X1    g276(.A1(pi002), .A2(pi015), .A3(pi020), .ZN(new_n567_));
  NAND2_X1   g277(.A1(new_n567_), .A2(new_n566_), .ZN(new_n568_));
  NAND2_X1   g278(.A1(new_n568_), .A2(pi082), .ZN(new_n569_));
  AOI22_X1   g279(.A1(new_n565_), .A2(pi082), .B1(new_n368_), .B2(new_n569_), .ZN(new_n570_));
  NOR2_X1    g280(.A1(new_n570_), .A2(pi024), .ZN(new_n571_));
  NOR4_X1    g281(.A1(new_n571_), .A2(pi129), .A3(new_n558_), .A4(new_n562_), .ZN(po039));
  INV_X1     g282(.I(pi053), .ZN(new_n573_));
  INV_X1     g283(.I(pi085), .ZN(new_n574_));
  INV_X1     g284(.I(pi026), .ZN(new_n575_));
  NOR3_X1    g285(.A1(pi039), .A2(pi051), .A3(pi052), .ZN(new_n576_));
  INV_X1     g286(.I(pi116), .ZN(new_n577_));
  NOR2_X1    g287(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1     g288(.I(pi110), .ZN(new_n579_));
  OR2_X2     g289(.A1(pi095), .A2(pi100), .Z(new_n580_));
  OAI21_X1   g290(.A1(new_n580_), .A2(pi097), .B(new_n579_), .ZN(new_n581_));
  AOI21_X1   g291(.A1(new_n581_), .A2(pi025), .B(new_n578_), .ZN(new_n582_));
  NAND2_X1   g292(.A1(new_n577_), .A2(pi025), .ZN(new_n583_));
  OAI22_X1   g293(.A1(new_n582_), .A2(new_n576_), .B1(new_n575_), .B2(new_n583_), .ZN(new_n584_));
  NOR2_X1    g294(.A1(new_n574_), .A2(new_n577_), .ZN(new_n585_));
  NOR3_X1    g295(.A1(pi085), .A2(pi096), .A3(pi110), .ZN(new_n586_));
  OAI21_X1   g296(.A1(new_n585_), .A2(new_n586_), .B(pi100), .ZN(new_n587_));
  NAND3_X1   g297(.A1(new_n577_), .A2(pi025), .A3(pi085), .ZN(new_n588_));
  AOI21_X1   g298(.A1(new_n587_), .A2(new_n588_), .B(pi026), .ZN(new_n589_));
  AOI21_X1   g299(.A1(new_n584_), .A2(new_n574_), .B(new_n589_), .ZN(new_n590_));
  INV_X1     g300(.I(pi027), .ZN(new_n591_));
  NAND2_X1   g301(.A1(new_n576_), .A2(pi116), .ZN(new_n592_));
  AOI21_X1   g302(.A1(new_n592_), .A2(new_n583_), .B(new_n591_), .ZN(new_n593_));
  AND3_X2    g303(.A1(new_n581_), .A2(pi025), .A3(new_n576_), .Z(new_n594_));
  NOR2_X1    g304(.A1(pi026), .A2(pi085), .ZN(new_n595_));
  OAI21_X1   g305(.A1(new_n594_), .A2(new_n593_), .B(new_n595_), .ZN(new_n596_));
  OAI21_X1   g306(.A1(new_n590_), .A2(pi027), .B(new_n596_), .ZN(new_n597_));
  NAND2_X1   g307(.A1(new_n573_), .A2(pi058), .ZN(new_n598_));
  INV_X1     g308(.I(pi058), .ZN(new_n599_));
  NAND2_X1   g309(.A1(new_n599_), .A2(pi053), .ZN(new_n600_));
  NAND2_X1   g310(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1   g311(.A1(new_n597_), .A2(new_n573_), .B(new_n601_), .ZN(new_n602_));
  NOR4_X1    g312(.A1(new_n583_), .A2(pi026), .A3(pi027), .A4(pi085), .ZN(new_n603_));
  NOR2_X1    g313(.A1(pi053), .A2(pi058), .ZN(new_n604_));
  NOR2_X1    g314(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR3_X1    g315(.A1(new_n602_), .A2(new_n418_), .A3(new_n605_), .ZN(po040));
  NAND3_X1   g316(.A1(new_n591_), .A2(new_n573_), .A3(new_n599_), .ZN(new_n607_));
  AOI21_X1   g317(.A1(new_n576_), .A2(pi116), .B(new_n575_), .ZN(new_n608_));
  INV_X1     g318(.I(new_n585_), .ZN(new_n609_));
  OAI21_X1   g319(.A1(new_n574_), .A2(pi116), .B(new_n579_), .ZN(new_n610_));
  INV_X1     g320(.I(pi096), .ZN(new_n611_));
  OAI21_X1   g321(.A1(new_n575_), .A2(new_n577_), .B(new_n611_), .ZN(new_n612_));
  OAI22_X1   g322(.A1(new_n609_), .A2(pi026), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  AOI22_X1   g323(.A1(new_n613_), .A2(pi100), .B1(new_n574_), .B2(new_n608_), .ZN(new_n614_));
  NOR3_X1    g324(.A1(new_n614_), .A2(new_n418_), .A3(new_n607_), .ZN(po041));
  NAND3_X1   g325(.A1(new_n592_), .A2(pi027), .A3(new_n574_), .ZN(new_n616_));
  INV_X1     g326(.I(pi100), .ZN(new_n617_));
  INV_X1     g327(.I(pi095), .ZN(new_n618_));
  NOR2_X1    g328(.A1(new_n618_), .A2(pi096), .ZN(new_n619_));
  NAND2_X1   g329(.A1(pi027), .A2(pi116), .ZN(new_n620_));
  NAND2_X1   g330(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI22_X1   g331(.A1(pi027), .A2(new_n609_), .B1(new_n621_), .B2(new_n610_), .ZN(new_n622_));
  NAND2_X1   g332(.A1(new_n622_), .A2(new_n617_), .ZN(new_n623_));
  NOR2_X1    g333(.A1(new_n418_), .A2(pi026), .ZN(new_n624_));
  NAND2_X1   g334(.A1(new_n624_), .A2(new_n604_), .ZN(new_n625_));
  AOI21_X1   g335(.A1(new_n623_), .A2(new_n616_), .B(new_n625_), .ZN(po042));
  INV_X1     g336(.I(new_n598_), .ZN(new_n627_));
  NOR3_X1    g337(.A1(new_n428_), .A2(pi027), .A3(pi116), .ZN(new_n628_));
  NAND3_X1   g338(.A1(new_n627_), .A2(new_n595_), .A3(new_n628_), .ZN(new_n629_));
  AND3_X2    g339(.A1(new_n628_), .A2(pi053), .A3(new_n595_), .Z(new_n630_));
  NAND2_X1   g340(.A1(new_n575_), .A2(new_n591_), .ZN(new_n631_));
  NOR2_X1    g341(.A1(new_n631_), .A2(new_n574_), .ZN(new_n632_));
  NOR2_X1    g342(.A1(new_n577_), .A2(pi100), .ZN(new_n633_));
  NOR2_X1    g343(.A1(new_n428_), .A2(pi116), .ZN(new_n634_));
  OAI21_X1   g344(.A1(new_n633_), .A2(new_n634_), .B(new_n632_), .ZN(new_n635_));
  NOR3_X1    g345(.A1(pi026), .A2(pi100), .A3(pi110), .ZN(new_n636_));
  AOI22_X1   g346(.A1(new_n578_), .A2(new_n576_), .B1(new_n619_), .B2(new_n636_), .ZN(new_n637_));
  NOR2_X1    g347(.A1(new_n576_), .A2(pi026), .ZN(new_n638_));
  INV_X1     g348(.I(new_n638_), .ZN(new_n639_));
  OAI22_X1   g349(.A1(new_n637_), .A2(pi027), .B1(new_n639_), .B2(new_n620_), .ZN(new_n640_));
  NOR4_X1    g350(.A1(pi027), .A2(pi039), .A3(pi051), .A4(pi052), .ZN(new_n641_));
  OAI21_X1   g351(.A1(new_n638_), .A2(new_n641_), .B(new_n581_), .ZN(new_n642_));
  XOR2_X1    g352(.A1(pi026), .A2(pi027), .Z(new_n643_));
  NAND2_X1   g353(.A1(new_n643_), .A2(new_n577_), .ZN(new_n644_));
  AOI21_X1   g354(.A1(new_n642_), .A2(new_n644_), .B(new_n428_), .ZN(new_n645_));
  OAI21_X1   g355(.A1(new_n645_), .A2(new_n640_), .B(new_n574_), .ZN(new_n646_));
  AOI21_X1   g356(.A1(new_n646_), .A2(new_n635_), .B(pi053), .ZN(new_n647_));
  OAI21_X1   g357(.A1(new_n647_), .A2(new_n630_), .B(new_n599_), .ZN(new_n648_));
  AOI21_X1   g358(.A1(new_n648_), .A2(new_n629_), .B(new_n418_), .ZN(po043));
  INV_X1     g359(.I(new_n604_), .ZN(new_n650_));
  NOR4_X1    g360(.A1(new_n650_), .A2(new_n575_), .A3(pi027), .A4(pi085), .ZN(new_n651_));
  NOR2_X1    g361(.A1(new_n434_), .A2(pi116), .ZN(new_n652_));
  NAND2_X1   g362(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1     g363(.I(new_n652_), .ZN(new_n654_));
  NOR3_X1    g364(.A1(new_n654_), .A2(new_n574_), .A3(new_n607_), .ZN(new_n655_));
  INV_X1     g365(.I(pi097), .ZN(new_n656_));
  NAND2_X1   g366(.A1(new_n656_), .A2(pi029), .ZN(new_n657_));
  NAND3_X1   g367(.A1(new_n611_), .A2(new_n579_), .A3(pi097), .ZN(new_n658_));
  AOI21_X1   g368(.A1(new_n658_), .A2(new_n657_), .B(new_n580_), .ZN(new_n659_));
  NOR2_X1    g369(.A1(new_n434_), .A2(new_n579_), .ZN(new_n660_));
  OAI21_X1   g370(.A1(new_n659_), .A2(new_n660_), .B(new_n599_), .ZN(new_n661_));
  NOR2_X1    g371(.A1(new_n656_), .A2(new_n577_), .ZN(new_n662_));
  OAI21_X1   g372(.A1(new_n662_), .A2(new_n652_), .B(pi058), .ZN(new_n663_));
  AOI21_X1   g373(.A1(new_n661_), .A2(new_n663_), .B(pi053), .ZN(new_n664_));
  NOR2_X1    g374(.A1(new_n654_), .A2(new_n600_), .ZN(new_n665_));
  OAI21_X1   g375(.A1(new_n664_), .A2(new_n665_), .B(new_n591_), .ZN(new_n666_));
  NAND3_X1   g376(.A1(new_n652_), .A2(pi027), .A3(new_n604_), .ZN(new_n667_));
  AOI21_X1   g377(.A1(new_n666_), .A2(new_n667_), .B(pi085), .ZN(new_n668_));
  OAI21_X1   g378(.A1(new_n668_), .A2(new_n655_), .B(new_n575_), .ZN(new_n669_));
  AOI21_X1   g379(.A1(new_n669_), .A2(new_n653_), .B(new_n418_), .ZN(po044));
  NAND2_X1   g380(.A1(pi088), .A2(pi106), .ZN(new_n671_));
  NOR2_X1    g381(.A1(pi030), .A2(pi109), .ZN(new_n672_));
  INV_X1     g382(.I(pi109), .ZN(new_n673_));
  NOR2_X1    g383(.A1(new_n673_), .A2(pi060), .ZN(new_n674_));
  OR3_X2     g384(.A1(new_n674_), .A2(pi106), .A3(new_n672_), .Z(new_n675_));
  AOI21_X1   g385(.A1(new_n675_), .A2(new_n671_), .B(pi129), .ZN(po045));
  NAND2_X1   g386(.A1(pi089), .A2(pi106), .ZN(new_n677_));
  INV_X1     g387(.I(pi106), .ZN(new_n678_));
  INV_X1     g388(.I(pi031), .ZN(new_n679_));
  NAND2_X1   g389(.A1(new_n679_), .A2(new_n673_), .ZN(new_n680_));
  INV_X1     g390(.I(pi030), .ZN(new_n681_));
  NAND2_X1   g391(.A1(new_n681_), .A2(pi109), .ZN(new_n682_));
  NAND3_X1   g392(.A1(new_n680_), .A2(new_n682_), .A3(new_n678_), .ZN(new_n683_));
  AOI21_X1   g393(.A1(new_n683_), .A2(new_n677_), .B(pi129), .ZN(po046));
  NAND2_X1   g394(.A1(pi099), .A2(pi106), .ZN(new_n685_));
  INV_X1     g395(.I(pi032), .ZN(new_n686_));
  NAND2_X1   g396(.A1(new_n686_), .A2(new_n673_), .ZN(new_n687_));
  NAND2_X1   g397(.A1(new_n679_), .A2(pi109), .ZN(new_n688_));
  NAND3_X1   g398(.A1(new_n687_), .A2(new_n688_), .A3(new_n678_), .ZN(new_n689_));
  AOI21_X1   g399(.A1(new_n689_), .A2(new_n685_), .B(pi129), .ZN(po047));
  NAND2_X1   g400(.A1(pi090), .A2(pi106), .ZN(new_n691_));
  INV_X1     g401(.I(pi033), .ZN(new_n692_));
  NAND2_X1   g402(.A1(new_n692_), .A2(new_n673_), .ZN(new_n693_));
  NAND2_X1   g403(.A1(new_n686_), .A2(pi109), .ZN(new_n694_));
  NAND3_X1   g404(.A1(new_n693_), .A2(new_n694_), .A3(new_n678_), .ZN(new_n695_));
  AOI21_X1   g405(.A1(new_n695_), .A2(new_n691_), .B(pi129), .ZN(po048));
  NAND2_X1   g406(.A1(pi091), .A2(pi106), .ZN(new_n697_));
  INV_X1     g407(.I(pi034), .ZN(new_n698_));
  NAND2_X1   g408(.A1(new_n698_), .A2(new_n673_), .ZN(new_n699_));
  NAND2_X1   g409(.A1(new_n692_), .A2(pi109), .ZN(new_n700_));
  NAND3_X1   g410(.A1(new_n699_), .A2(new_n700_), .A3(new_n678_), .ZN(new_n701_));
  AOI21_X1   g411(.A1(new_n701_), .A2(new_n697_), .B(pi129), .ZN(po049));
  NAND2_X1   g412(.A1(pi092), .A2(pi106), .ZN(new_n703_));
  INV_X1     g413(.I(pi035), .ZN(new_n704_));
  NAND2_X1   g414(.A1(new_n704_), .A2(new_n673_), .ZN(new_n705_));
  NAND2_X1   g415(.A1(new_n698_), .A2(pi109), .ZN(new_n706_));
  NAND3_X1   g416(.A1(new_n705_), .A2(new_n706_), .A3(new_n678_), .ZN(new_n707_));
  AOI21_X1   g417(.A1(new_n707_), .A2(new_n703_), .B(pi129), .ZN(po050));
  NAND2_X1   g418(.A1(pi098), .A2(pi106), .ZN(new_n709_));
  INV_X1     g419(.I(pi036), .ZN(new_n710_));
  NAND2_X1   g420(.A1(new_n710_), .A2(new_n673_), .ZN(new_n711_));
  NAND2_X1   g421(.A1(new_n704_), .A2(pi109), .ZN(new_n712_));
  NAND3_X1   g422(.A1(new_n711_), .A2(new_n712_), .A3(new_n678_), .ZN(new_n713_));
  AOI21_X1   g423(.A1(new_n713_), .A2(new_n709_), .B(pi129), .ZN(po051));
  NAND2_X1   g424(.A1(pi093), .A2(pi106), .ZN(new_n715_));
  INV_X1     g425(.I(pi037), .ZN(new_n716_));
  NAND2_X1   g426(.A1(new_n716_), .A2(new_n673_), .ZN(new_n717_));
  NAND2_X1   g427(.A1(new_n710_), .A2(pi109), .ZN(new_n718_));
  NAND3_X1   g428(.A1(new_n717_), .A2(new_n718_), .A3(new_n678_), .ZN(new_n719_));
  AOI21_X1   g429(.A1(new_n719_), .A2(new_n715_), .B(pi129), .ZN(po052));
  NAND2_X1   g430(.A1(new_n370_), .A2(pi082), .ZN(new_n721_));
  NOR4_X1    g431(.A1(new_n721_), .A2(new_n387_), .A3(pi040), .A4(pi042), .ZN(new_n722_));
  NOR3_X1    g432(.A1(new_n383_), .A2(new_n377_), .A3(new_n399_), .ZN(new_n723_));
  OAI21_X1   g433(.A1(new_n723_), .A2(new_n369_), .B(new_n368_), .ZN(new_n724_));
  NAND2_X1   g434(.A1(new_n372_), .A2(pi082), .ZN(new_n725_));
  AOI21_X1   g435(.A1(new_n724_), .A2(new_n725_), .B(pi038), .ZN(new_n726_));
  INV_X1     g436(.I(pi074), .ZN(new_n727_));
  NOR2_X1    g437(.A1(new_n372_), .A2(pi050), .ZN(new_n728_));
  NAND3_X1   g438(.A1(new_n397_), .A2(new_n527_), .A3(new_n378_), .ZN(new_n729_));
  NOR4_X1    g439(.A1(new_n729_), .A2(pi046), .A3(pi047), .A4(new_n492_), .ZN(new_n730_));
  AOI21_X1   g440(.A1(new_n730_), .A2(new_n728_), .B(new_n369_), .ZN(new_n731_));
  NOR3_X1    g441(.A1(new_n731_), .A2(new_n727_), .A3(new_n368_), .ZN(new_n732_));
  NOR4_X1    g442(.A1(new_n726_), .A2(pi129), .A3(new_n722_), .A4(new_n732_), .ZN(po053));
  NAND2_X1   g443(.A1(new_n576_), .A2(pi109), .ZN(new_n734_));
  INV_X1     g444(.I(pi052), .ZN(new_n735_));
  NOR2_X1    g445(.A1(new_n673_), .A2(pi051), .ZN(new_n736_));
  NAND2_X1   g446(.A1(new_n736_), .A2(new_n735_), .ZN(new_n737_));
  AOI21_X1   g447(.A1(new_n737_), .A2(pi039), .B(pi106), .ZN(new_n738_));
  AOI21_X1   g448(.A1(new_n738_), .A2(new_n734_), .B(pi129), .ZN(po054));
  INV_X1     g449(.I(pi073), .ZN(new_n740_));
  NOR2_X1    g450(.A1(new_n534_), .A2(new_n389_), .ZN(new_n741_));
  AOI21_X1   g451(.A1(new_n730_), .A2(new_n741_), .B(new_n369_), .ZN(new_n742_));
  NOR3_X1    g452(.A1(new_n742_), .A2(new_n740_), .A3(new_n368_), .ZN(new_n743_));
  NOR2_X1    g453(.A1(new_n561_), .A2(new_n400_), .ZN(new_n744_));
  OAI21_X1   g454(.A1(new_n390_), .A2(new_n369_), .B(new_n368_), .ZN(new_n745_));
  NAND2_X1   g455(.A1(new_n534_), .A2(pi082), .ZN(new_n746_));
  AOI21_X1   g456(.A1(new_n745_), .A2(new_n746_), .B(pi040), .ZN(new_n747_));
  NOR4_X1    g457(.A1(new_n747_), .A2(pi129), .A3(new_n743_), .A4(new_n744_), .ZN(po055));
  INV_X1     g458(.I(pi076), .ZN(new_n749_));
  NOR2_X1    g459(.A1(new_n729_), .A2(new_n402_), .ZN(new_n750_));
  NAND2_X1   g460(.A1(new_n374_), .A2(new_n375_), .ZN(new_n751_));
  NOR3_X1    g461(.A1(new_n751_), .A2(pi046), .A3(pi050), .ZN(new_n752_));
  AOI21_X1   g462(.A1(new_n750_), .A2(new_n752_), .B(new_n369_), .ZN(new_n753_));
  NOR3_X1    g463(.A1(new_n753_), .A2(new_n749_), .A3(new_n368_), .ZN(new_n754_));
  NAND2_X1   g464(.A1(new_n533_), .A2(new_n385_), .ZN(new_n755_));
  NOR3_X1    g465(.A1(new_n755_), .A2(new_n384_), .A3(new_n561_), .ZN(new_n756_));
  NOR2_X1    g466(.A1(new_n383_), .A2(new_n377_), .ZN(new_n757_));
  NAND4_X1   g467(.A1(new_n490_), .A2(new_n370_), .A3(new_n371_), .A4(pi082), .ZN(new_n758_));
  NOR2_X1    g468(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1   g469(.A1(new_n563_), .A2(pi082), .B(new_n368_), .ZN(new_n760_));
  NOR3_X1    g470(.A1(new_n759_), .A2(pi041), .A3(new_n760_), .ZN(new_n761_));
  NOR4_X1    g471(.A1(new_n761_), .A2(pi129), .A3(new_n754_), .A4(new_n756_), .ZN(po056));
  INV_X1     g472(.I(pi072), .ZN(new_n763_));
  NOR2_X1    g473(.A1(new_n559_), .A2(pi044), .ZN(new_n764_));
  AOI21_X1   g474(.A1(new_n730_), .A2(new_n764_), .B(new_n369_), .ZN(new_n765_));
  NOR3_X1    g475(.A1(new_n765_), .A2(new_n763_), .A3(new_n368_), .ZN(new_n766_));
  INV_X1     g476(.I(pi042), .ZN(new_n767_));
  NOR2_X1    g477(.A1(new_n721_), .A2(new_n767_), .ZN(new_n768_));
  NOR2_X1    g478(.A1(new_n370_), .A2(new_n369_), .ZN(new_n769_));
  NOR3_X1    g479(.A1(new_n729_), .A2(new_n564_), .A3(new_n755_), .ZN(new_n770_));
  OAI22_X1   g480(.A1(new_n770_), .A2(new_n721_), .B1(new_n368_), .B2(new_n769_), .ZN(new_n771_));
  NOR2_X1    g481(.A1(new_n771_), .A2(pi042), .ZN(new_n772_));
  NOR4_X1    g482(.A1(new_n766_), .A2(new_n772_), .A3(pi129), .A4(new_n768_), .ZN(po057));
  NAND2_X1   g483(.A1(new_n371_), .A2(new_n387_), .ZN(new_n774_));
  NOR3_X1    g484(.A1(new_n399_), .A2(new_n774_), .A3(new_n721_), .ZN(new_n775_));
  INV_X1     g485(.I(new_n775_), .ZN(new_n776_));
  NOR2_X1    g486(.A1(new_n776_), .A2(new_n374_), .ZN(new_n777_));
  INV_X1     g487(.I(new_n403_), .ZN(new_n778_));
  NAND2_X1   g488(.A1(new_n382_), .A2(new_n554_), .ZN(new_n779_));
  NAND2_X1   g489(.A1(new_n779_), .A2(pi082), .ZN(new_n780_));
  AOI22_X1   g490(.A1(new_n780_), .A2(new_n368_), .B1(pi082), .B2(new_n778_), .ZN(new_n781_));
  NOR2_X1    g491(.A1(new_n781_), .A2(pi043), .ZN(new_n782_));
  INV_X1     g492(.I(new_n729_), .ZN(new_n783_));
  NAND3_X1   g493(.A1(new_n783_), .A2(new_n403_), .A3(new_n375_), .ZN(new_n784_));
  NAND2_X1   g494(.A1(new_n367_), .A2(pi077), .ZN(new_n785_));
  AOI21_X1   g495(.A1(new_n784_), .A2(pi082), .B(new_n785_), .ZN(new_n786_));
  NOR4_X1    g496(.A1(new_n782_), .A2(pi129), .A3(new_n777_), .A4(new_n786_), .ZN(po058));
  NAND4_X1   g497(.A1(new_n730_), .A2(new_n387_), .A3(new_n388_), .A4(new_n371_), .ZN(new_n788_));
  NAND2_X1   g498(.A1(new_n788_), .A2(pi082), .ZN(new_n789_));
  NAND2_X1   g499(.A1(new_n367_), .A2(pi067), .ZN(new_n790_));
  OAI21_X1   g500(.A1(pi044), .A2(new_n367_), .B(new_n790_), .ZN(new_n791_));
  INV_X1     g501(.I(pi129), .ZN(new_n792_));
  OAI21_X1   g502(.A1(new_n370_), .A2(new_n369_), .B(new_n792_), .ZN(new_n793_));
  AOI21_X1   g503(.A1(new_n789_), .A2(new_n791_), .B(new_n793_), .ZN(po059));
  NOR3_X1    g504(.A1(new_n776_), .A2(new_n379_), .A3(new_n377_), .ZN(new_n795_));
  INV_X1     g505(.I(pi068), .ZN(new_n796_));
  INV_X1     g506(.I(new_n404_), .ZN(new_n797_));
  AND3_X2    g507(.A1(new_n382_), .A2(new_n378_), .A3(new_n394_), .Z(new_n798_));
  AOI21_X1   g508(.A1(new_n797_), .A2(new_n798_), .B(new_n369_), .ZN(new_n799_));
  NOR3_X1    g509(.A1(new_n799_), .A2(new_n796_), .A3(new_n368_), .ZN(new_n800_));
  OAI21_X1   g510(.A1(new_n568_), .A2(pi024), .B(pi082), .ZN(new_n801_));
  NAND2_X1   g511(.A1(new_n801_), .A2(new_n368_), .ZN(new_n802_));
  NAND2_X1   g512(.A1(new_n526_), .A2(new_n528_), .ZN(new_n803_));
  OAI21_X1   g513(.A1(new_n803_), .A2(pi048), .B(pi082), .ZN(new_n804_));
  AOI21_X1   g514(.A1(new_n804_), .A2(new_n802_), .B(pi045), .ZN(new_n805_));
  NOR4_X1    g515(.A1(new_n800_), .A2(pi129), .A3(new_n795_), .A4(new_n805_), .ZN(po060));
  INV_X1     g516(.I(pi075), .ZN(new_n807_));
  NOR2_X1    g517(.A1(new_n729_), .A2(new_n564_), .ZN(new_n808_));
  NOR2_X1    g518(.A1(new_n402_), .A2(pi050), .ZN(new_n809_));
  AOI21_X1   g519(.A1(new_n808_), .A2(new_n809_), .B(new_n369_), .ZN(new_n810_));
  NOR3_X1    g520(.A1(new_n810_), .A2(new_n807_), .A3(new_n368_), .ZN(new_n811_));
  NOR4_X1    g521(.A1(new_n402_), .A2(new_n385_), .A3(pi050), .A4(new_n369_), .ZN(new_n812_));
  OAI21_X1   g522(.A1(new_n372_), .A2(new_n389_), .B(pi082), .ZN(new_n813_));
  OAI21_X1   g523(.A1(new_n808_), .A2(new_n369_), .B(new_n368_), .ZN(new_n814_));
  AOI21_X1   g524(.A1(new_n814_), .A2(new_n813_), .B(pi046), .ZN(new_n815_));
  NOR4_X1    g525(.A1(new_n811_), .A2(new_n815_), .A3(pi129), .A4(new_n812_), .ZN(po061));
  NOR3_X1    g526(.A1(new_n758_), .A2(new_n375_), .A3(new_n492_), .ZN(new_n817_));
  NOR3_X1    g527(.A1(new_n404_), .A2(new_n369_), .A3(new_n783_), .ZN(new_n818_));
  AOI21_X1   g528(.A1(new_n404_), .A2(pi082), .B(new_n368_), .ZN(new_n819_));
  NOR3_X1    g529(.A1(new_n818_), .A2(new_n819_), .A3(pi047), .ZN(new_n820_));
  INV_X1     g530(.I(pi064), .ZN(new_n821_));
  AOI21_X1   g531(.A1(new_n797_), .A2(new_n783_), .B(new_n369_), .ZN(new_n822_));
  NOR3_X1    g532(.A1(new_n822_), .A2(new_n821_), .A3(new_n368_), .ZN(new_n823_));
  NOR4_X1    g533(.A1(new_n823_), .A2(pi129), .A3(new_n817_), .A4(new_n820_), .ZN(po062));
  NOR4_X1    g534(.A1(new_n404_), .A2(pi002), .A3(pi047), .A4(new_n398_), .ZN(new_n825_));
  OAI21_X1   g535(.A1(new_n825_), .A2(new_n369_), .B(pi062), .ZN(new_n826_));
  NOR2_X1    g536(.A1(new_n826_), .A2(new_n368_), .ZN(new_n827_));
  NOR3_X1    g537(.A1(new_n776_), .A2(new_n376_), .A3(new_n751_), .ZN(new_n828_));
  NAND2_X1   g538(.A1(new_n383_), .A2(pi082), .ZN(new_n829_));
  AOI22_X1   g539(.A1(new_n829_), .A2(new_n368_), .B1(pi082), .B2(new_n803_), .ZN(new_n830_));
  NOR2_X1    g540(.A1(new_n830_), .A2(pi048), .ZN(new_n831_));
  NOR4_X1    g541(.A1(new_n827_), .A2(pi129), .A3(new_n831_), .A4(new_n828_), .ZN(po063));
  INV_X1     g542(.I(pi069), .ZN(new_n833_));
  NOR3_X1    g543(.A1(new_n560_), .A2(pi050), .A3(new_n402_), .ZN(new_n834_));
  NAND2_X1   g544(.A1(new_n834_), .A2(new_n380_), .ZN(new_n835_));
  AOI21_X1   g545(.A1(new_n835_), .A2(pi082), .B(new_n368_), .ZN(new_n836_));
  NOR2_X1    g546(.A1(new_n367_), .A2(new_n566_), .ZN(new_n837_));
  AOI22_X1   g547(.A1(new_n836_), .A2(new_n833_), .B1(new_n369_), .B2(new_n837_), .ZN(new_n838_));
  NOR4_X1    g548(.A1(new_n560_), .A2(pi024), .A3(new_n534_), .A4(new_n559_), .ZN(new_n839_));
  OAI22_X1   g549(.A1(new_n835_), .A2(new_n567_), .B1(new_n566_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1   g550(.A1(new_n840_), .A2(pi082), .ZN(new_n841_));
  AOI21_X1   g551(.A1(new_n838_), .A2(new_n841_), .B(pi129), .ZN(po064));
  INV_X1     g552(.I(pi066), .ZN(new_n843_));
  INV_X1     g553(.I(new_n402_), .ZN(new_n844_));
  AOI21_X1   g554(.A1(new_n730_), .A2(new_n844_), .B(new_n369_), .ZN(new_n845_));
  NOR3_X1    g555(.A1(new_n845_), .A2(new_n843_), .A3(new_n368_), .ZN(new_n846_));
  NOR3_X1    g556(.A1(new_n774_), .A2(new_n388_), .A3(new_n721_), .ZN(new_n847_));
  NAND4_X1   g557(.A1(new_n394_), .A2(new_n491_), .A3(new_n378_), .A4(new_n385_), .ZN(new_n848_));
  OAI21_X1   g558(.A1(new_n848_), .A2(new_n398_), .B(pi082), .ZN(new_n849_));
  AOI22_X1   g559(.A1(new_n849_), .A2(new_n368_), .B1(pi082), .B2(new_n402_), .ZN(new_n850_));
  NOR2_X1    g560(.A1(new_n850_), .A2(pi050), .ZN(new_n851_));
  NOR4_X1    g561(.A1(new_n846_), .A2(new_n851_), .A3(pi129), .A4(new_n847_), .ZN(po065));
  XNOR2_X1   g562(.A1(pi051), .A2(pi109), .ZN(new_n853_));
  AOI21_X1   g563(.A1(new_n853_), .A2(new_n678_), .B(pi129), .ZN(po066));
  XOR2_X1    g564(.A1(new_n736_), .A2(new_n735_), .Z(new_n855_));
  AOI21_X1   g565(.A1(new_n855_), .A2(new_n678_), .B(pi129), .ZN(po067));
  INV_X1     g566(.I(new_n624_), .ZN(new_n857_));
  NAND2_X1   g567(.A1(pi058), .A2(pi116), .ZN(new_n858_));
  INV_X1     g568(.I(new_n580_), .ZN(new_n859_));
  NAND4_X1   g569(.A1(new_n859_), .A2(new_n599_), .A3(new_n611_), .A4(new_n579_), .ZN(new_n860_));
  AOI21_X1   g570(.A1(new_n860_), .A2(new_n858_), .B(new_n656_), .ZN(new_n861_));
  NAND2_X1   g571(.A1(new_n599_), .A2(new_n577_), .ZN(new_n862_));
  NOR2_X1    g572(.A1(new_n862_), .A2(new_n573_), .ZN(new_n863_));
  AOI21_X1   g573(.A1(new_n861_), .A2(new_n573_), .B(new_n863_), .ZN(new_n864_));
  NOR4_X1    g574(.A1(new_n864_), .A2(pi027), .A3(pi085), .A4(new_n857_), .ZN(po068));
  NOR2_X1    g575(.A1(new_n404_), .A2(new_n779_), .ZN(new_n866_));
  OAI21_X1   g576(.A1(new_n866_), .A2(new_n369_), .B(new_n367_), .ZN(new_n867_));
  NAND2_X1   g577(.A1(new_n867_), .A2(new_n792_), .ZN(po069));
  INV_X1     g578(.I(pi114), .ZN(new_n869_));
  NAND2_X1   g579(.A1(new_n409_), .A2(new_n792_), .ZN(po129));
  NOR3_X1    g580(.A1(po129), .A2(new_n869_), .A3(pi122), .ZN(po070));
  OAI22_X1   g581(.A1(new_n862_), .A2(new_n716_), .B1(pi026), .B2(new_n858_), .ZN(new_n872_));
  NOR2_X1    g582(.A1(new_n578_), .A2(pi058), .ZN(new_n873_));
  OAI21_X1   g583(.A1(new_n575_), .A2(new_n599_), .B(pi094), .ZN(new_n874_));
  NOR2_X1    g584(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1   g585(.A1(new_n875_), .A2(new_n872_), .B(new_n573_), .ZN(new_n876_));
  NAND3_X1   g586(.A1(new_n575_), .A2(new_n599_), .A3(pi037), .ZN(new_n877_));
  AOI21_X1   g587(.A1(new_n876_), .A2(new_n877_), .B(pi085), .ZN(new_n878_));
  NOR3_X1    g588(.A1(new_n650_), .A2(pi026), .A3(new_n716_), .ZN(new_n879_));
  OAI21_X1   g589(.A1(new_n878_), .A2(new_n879_), .B(new_n591_), .ZN(new_n880_));
  NAND2_X1   g590(.A1(new_n879_), .A2(new_n574_), .ZN(new_n881_));
  AOI21_X1   g591(.A1(new_n880_), .A2(new_n881_), .B(new_n418_), .ZN(po071));
  NOR3_X1    g592(.A1(pi026), .A2(pi053), .A3(pi085), .ZN(new_n883_));
  NAND3_X1   g593(.A1(new_n883_), .A2(pi057), .A3(new_n599_), .ZN(new_n884_));
  INV_X1     g594(.I(pi057), .ZN(new_n885_));
  NAND2_X1   g595(.A1(new_n883_), .A2(new_n577_), .ZN(new_n886_));
  OAI21_X1   g596(.A1(pi026), .A2(pi053), .B(pi085), .ZN(new_n887_));
  NAND2_X1   g597(.A1(pi026), .A2(pi053), .ZN(new_n888_));
  NAND3_X1   g598(.A1(new_n887_), .A2(new_n888_), .A3(new_n599_), .ZN(new_n889_));
  AOI21_X1   g599(.A1(new_n889_), .A2(new_n886_), .B(new_n885_), .ZN(new_n890_));
  NAND2_X1   g600(.A1(new_n883_), .A2(pi060), .ZN(new_n891_));
  NOR2_X1    g601(.A1(new_n891_), .A2(new_n858_), .ZN(new_n892_));
  OAI21_X1   g602(.A1(new_n890_), .A2(new_n892_), .B(new_n591_), .ZN(new_n893_));
  AOI21_X1   g603(.A1(new_n893_), .A2(new_n884_), .B(new_n418_), .ZN(po072));
  INV_X1     g604(.I(new_n631_), .ZN(new_n895_));
  NOR2_X1    g605(.A1(new_n599_), .A2(pi116), .ZN(new_n896_));
  NOR2_X1    g606(.A1(new_n592_), .A2(pi058), .ZN(new_n897_));
  AOI22_X1   g607(.A1(new_n897_), .A2(new_n643_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n898_));
  NOR4_X1    g608(.A1(new_n898_), .A2(pi053), .A3(pi085), .A4(new_n418_), .ZN(po073));
  NAND3_X1   g609(.A1(new_n651_), .A2(pi059), .A3(new_n577_), .ZN(new_n900_));
  NAND4_X1   g610(.A1(new_n604_), .A2(pi059), .A3(new_n577_), .A4(pi085), .ZN(new_n901_));
  NOR3_X1    g611(.A1(new_n581_), .A2(new_n611_), .A3(new_n650_), .ZN(new_n902_));
  AOI22_X1   g612(.A1(new_n581_), .A2(new_n604_), .B1(new_n601_), .B2(new_n577_), .ZN(new_n903_));
  NOR2_X1    g613(.A1(new_n903_), .A2(new_n513_), .ZN(new_n904_));
  OAI21_X1   g614(.A1(new_n904_), .A2(new_n902_), .B(new_n574_), .ZN(new_n905_));
  AOI21_X1   g615(.A1(new_n905_), .A2(new_n901_), .B(pi027), .ZN(new_n906_));
  NAND2_X1   g616(.A1(new_n577_), .A2(pi059), .ZN(new_n907_));
  NOR4_X1    g617(.A1(new_n650_), .A2(new_n907_), .A3(new_n591_), .A4(pi085), .ZN(new_n908_));
  OAI21_X1   g618(.A1(new_n906_), .A2(new_n908_), .B(new_n575_), .ZN(new_n909_));
  AOI21_X1   g619(.A1(new_n909_), .A2(new_n900_), .B(new_n418_), .ZN(po074));
  NOR2_X1    g620(.A1(pi117), .A2(pi122), .ZN(new_n911_));
  MUX2_X1    g621(.I0(pi060), .I1(pi123), .S(new_n911_), .Z(po075));
  NOR4_X1    g622(.A1(new_n409_), .A2(pi114), .A3(pi122), .A4(pi129), .ZN(po076));
  INV_X1     g623(.I(pi062), .ZN(new_n914_));
  NAND3_X1   g624(.A1(pi131), .A2(pi132), .A3(pi133), .ZN(new_n915_));
  NOR2_X1    g625(.A1(new_n915_), .A2(pi138), .ZN(new_n916_));
  INV_X1     g626(.I(pi136), .ZN(new_n917_));
  NOR2_X1    g627(.A1(new_n917_), .A2(pi137), .ZN(new_n918_));
  NAND2_X1   g628(.A1(new_n916_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1     g629(.I(new_n919_), .ZN(new_n920_));
  NOR2_X1    g630(.A1(new_n920_), .A2(new_n914_), .ZN(new_n921_));
  NOR2_X1    g631(.A1(new_n919_), .A2(pi140), .ZN(new_n922_));
  OAI21_X1   g632(.A1(new_n921_), .A2(new_n922_), .B(new_n792_), .ZN(po077));
  NOR2_X1    g633(.A1(new_n920_), .A2(new_n553_), .ZN(new_n924_));
  NOR2_X1    g634(.A1(new_n919_), .A2(pi142), .ZN(new_n925_));
  OAI21_X1   g635(.A1(new_n924_), .A2(new_n925_), .B(new_n792_), .ZN(po078));
  NOR2_X1    g636(.A1(new_n920_), .A2(new_n821_), .ZN(new_n927_));
  NOR2_X1    g637(.A1(new_n919_), .A2(pi139), .ZN(new_n928_));
  OAI21_X1   g638(.A1(new_n927_), .A2(new_n928_), .B(new_n792_), .ZN(po079));
  AND2_X2    g639(.A1(new_n919_), .A2(pi065), .Z(new_n930_));
  NOR2_X1    g640(.A1(new_n919_), .A2(pi146), .ZN(new_n931_));
  OAI21_X1   g641(.A1(new_n930_), .A2(new_n931_), .B(new_n792_), .ZN(po080));
  INV_X1     g642(.I(new_n916_), .ZN(new_n933_));
  NOR2_X1    g643(.A1(pi136), .A2(pi137), .ZN(new_n934_));
  INV_X1     g644(.I(new_n934_), .ZN(new_n935_));
  NOR2_X1    g645(.A1(new_n933_), .A2(new_n935_), .ZN(new_n936_));
  INV_X1     g646(.I(new_n936_), .ZN(new_n937_));
  NOR2_X1    g647(.A1(new_n937_), .A2(pi143), .ZN(new_n938_));
  NOR2_X1    g648(.A1(new_n936_), .A2(new_n843_), .ZN(new_n939_));
  OAI21_X1   g649(.A1(new_n938_), .A2(new_n939_), .B(new_n792_), .ZN(po081));
  NOR2_X1    g650(.A1(new_n937_), .A2(pi139), .ZN(new_n941_));
  INV_X1     g651(.I(pi067), .ZN(new_n942_));
  NOR2_X1    g652(.A1(new_n936_), .A2(new_n942_), .ZN(new_n943_));
  OAI21_X1   g653(.A1(new_n941_), .A2(new_n943_), .B(new_n792_), .ZN(po082));
  NOR2_X1    g654(.A1(new_n920_), .A2(new_n796_), .ZN(new_n945_));
  NOR2_X1    g655(.A1(new_n919_), .A2(pi141), .ZN(new_n946_));
  OAI21_X1   g656(.A1(new_n945_), .A2(new_n946_), .B(new_n792_), .ZN(po083));
  NOR2_X1    g657(.A1(new_n920_), .A2(new_n833_), .ZN(new_n948_));
  NOR2_X1    g658(.A1(new_n919_), .A2(pi143), .ZN(new_n949_));
  OAI21_X1   g659(.A1(new_n948_), .A2(new_n949_), .B(new_n792_), .ZN(po084));
  NOR2_X1    g660(.A1(new_n920_), .A2(new_n489_), .ZN(new_n951_));
  NOR2_X1    g661(.A1(new_n919_), .A2(pi144), .ZN(new_n952_));
  OAI21_X1   g662(.A1(new_n951_), .A2(new_n952_), .B(new_n792_), .ZN(po085));
  NOR2_X1    g663(.A1(new_n920_), .A2(new_n525_), .ZN(new_n954_));
  NOR2_X1    g664(.A1(new_n919_), .A2(pi145), .ZN(new_n955_));
  OAI21_X1   g665(.A1(new_n954_), .A2(new_n955_), .B(new_n792_), .ZN(po086));
  NOR2_X1    g666(.A1(new_n937_), .A2(pi140), .ZN(new_n957_));
  NOR2_X1    g667(.A1(new_n936_), .A2(new_n763_), .ZN(new_n958_));
  OAI21_X1   g668(.A1(new_n957_), .A2(new_n958_), .B(new_n792_), .ZN(po087));
  NOR2_X1    g669(.A1(new_n937_), .A2(pi141), .ZN(new_n960_));
  NOR2_X1    g670(.A1(new_n936_), .A2(new_n740_), .ZN(new_n961_));
  OAI21_X1   g671(.A1(new_n960_), .A2(new_n961_), .B(new_n792_), .ZN(po088));
  NOR2_X1    g672(.A1(new_n937_), .A2(pi142), .ZN(new_n963_));
  NOR2_X1    g673(.A1(new_n936_), .A2(new_n727_), .ZN(new_n964_));
  OAI21_X1   g674(.A1(new_n963_), .A2(new_n964_), .B(new_n792_), .ZN(po089));
  NOR2_X1    g675(.A1(new_n937_), .A2(pi144), .ZN(new_n966_));
  NOR2_X1    g676(.A1(new_n936_), .A2(new_n807_), .ZN(new_n967_));
  OAI21_X1   g677(.A1(new_n966_), .A2(new_n967_), .B(new_n792_), .ZN(po090));
  NOR2_X1    g678(.A1(new_n937_), .A2(pi145), .ZN(new_n969_));
  NOR2_X1    g679(.A1(new_n936_), .A2(new_n749_), .ZN(new_n970_));
  OAI21_X1   g680(.A1(new_n969_), .A2(new_n970_), .B(new_n792_), .ZN(po091));
  NOR2_X1    g681(.A1(new_n937_), .A2(pi146), .ZN(new_n972_));
  INV_X1     g682(.I(pi077), .ZN(new_n973_));
  NOR2_X1    g683(.A1(new_n936_), .A2(new_n973_), .ZN(new_n974_));
  OAI21_X1   g684(.A1(new_n972_), .A2(new_n974_), .B(new_n792_), .ZN(po092));
  INV_X1     g685(.I(pi137), .ZN(new_n976_));
  NOR2_X1    g686(.A1(new_n976_), .A2(pi136), .ZN(new_n977_));
  NAND2_X1   g687(.A1(new_n916_), .A2(new_n977_), .ZN(new_n978_));
  INV_X1     g688(.I(new_n978_), .ZN(new_n979_));
  NAND2_X1   g689(.A1(new_n979_), .A2(pi142), .ZN(new_n980_));
  NAND2_X1   g690(.A1(new_n978_), .A2(pi078), .ZN(new_n981_));
  AOI21_X1   g691(.A1(new_n980_), .A2(new_n981_), .B(pi129), .ZN(po093));
  NAND2_X1   g692(.A1(new_n979_), .A2(pi143), .ZN(new_n983_));
  NAND2_X1   g693(.A1(new_n978_), .A2(pi079), .ZN(new_n984_));
  AOI21_X1   g694(.A1(new_n983_), .A2(new_n984_), .B(pi129), .ZN(po094));
  NAND2_X1   g695(.A1(new_n979_), .A2(pi144), .ZN(new_n986_));
  NAND2_X1   g696(.A1(new_n978_), .A2(pi080), .ZN(new_n987_));
  AOI21_X1   g697(.A1(new_n986_), .A2(new_n987_), .B(pi129), .ZN(po095));
  NAND2_X1   g698(.A1(new_n979_), .A2(pi145), .ZN(new_n989_));
  NAND2_X1   g699(.A1(new_n978_), .A2(pi081), .ZN(new_n990_));
  AOI21_X1   g700(.A1(new_n989_), .A2(new_n990_), .B(pi129), .ZN(po096));
  NAND2_X1   g701(.A1(new_n979_), .A2(pi146), .ZN(new_n992_));
  NAND2_X1   g702(.A1(new_n978_), .A2(pi082), .ZN(new_n993_));
  AOI21_X1   g703(.A1(new_n992_), .A2(new_n993_), .B(pi129), .ZN(po097));
  INV_X1     g704(.I(pi115), .ZN(new_n995_));
  INV_X1     g705(.I(pi138), .ZN(new_n996_));
  NOR2_X1    g706(.A1(new_n995_), .A2(new_n996_), .ZN(new_n997_));
  NOR2_X1    g707(.A1(pi087), .A2(pi138), .ZN(new_n998_));
  NOR3_X1    g708(.A1(new_n997_), .A2(pi136), .A3(new_n998_), .ZN(new_n999_));
  NOR3_X1    g709(.A1(new_n679_), .A2(new_n917_), .A3(pi138), .ZN(new_n1000_));
  NOR3_X1    g710(.A1(new_n999_), .A2(new_n976_), .A3(new_n1000_), .ZN(new_n1001_));
  NAND2_X1   g711(.A1(pi089), .A2(pi138), .ZN(new_n1002_));
  NAND2_X1   g712(.A1(new_n914_), .A2(new_n996_), .ZN(new_n1003_));
  AOI21_X1   g713(.A1(new_n1003_), .A2(new_n1002_), .B(new_n917_), .ZN(new_n1004_));
  NAND2_X1   g714(.A1(pi119), .A2(pi138), .ZN(new_n1005_));
  NAND2_X1   g715(.A1(new_n763_), .A2(new_n996_), .ZN(new_n1006_));
  AOI21_X1   g716(.A1(new_n1006_), .A2(new_n1005_), .B(pi136), .ZN(new_n1007_));
  NOR3_X1    g717(.A1(new_n1004_), .A2(new_n1007_), .A3(pi137), .ZN(new_n1008_));
  NOR2_X1    g718(.A1(new_n1008_), .A2(new_n1001_), .ZN(po098));
  NAND2_X1   g719(.A1(new_n979_), .A2(pi141), .ZN(new_n1010_));
  NAND2_X1   g720(.A1(new_n978_), .A2(pi084), .ZN(new_n1011_));
  AOI21_X1   g721(.A1(new_n1010_), .A2(new_n1011_), .B(pi129), .ZN(po099));
  NOR2_X1    g722(.A1(new_n581_), .A2(pi085), .ZN(new_n1013_));
  AOI22_X1   g723(.A1(new_n1013_), .A2(pi096), .B1(pi085), .B2(new_n577_), .ZN(new_n1014_));
  NOR3_X1    g724(.A1(new_n1014_), .A2(new_n607_), .A3(new_n857_), .ZN(po100));
  NAND2_X1   g725(.A1(new_n979_), .A2(pi139), .ZN(new_n1016_));
  NAND2_X1   g726(.A1(new_n978_), .A2(pi086), .ZN(new_n1017_));
  AOI21_X1   g727(.A1(new_n1016_), .A2(new_n1017_), .B(pi129), .ZN(po101));
  NAND2_X1   g728(.A1(new_n979_), .A2(pi140), .ZN(new_n1019_));
  NAND2_X1   g729(.A1(new_n978_), .A2(pi087), .ZN(new_n1020_));
  AOI21_X1   g730(.A1(new_n1019_), .A2(new_n1020_), .B(pi129), .ZN(po102));
  NOR3_X1    g731(.A1(new_n933_), .A2(new_n917_), .A3(new_n976_), .ZN(new_n1022_));
  NAND2_X1   g732(.A1(new_n1022_), .A2(pi139), .ZN(new_n1023_));
  INV_X1     g733(.I(new_n1022_), .ZN(new_n1024_));
  NAND2_X1   g734(.A1(new_n1024_), .A2(pi088), .ZN(new_n1025_));
  AOI21_X1   g735(.A1(new_n1025_), .A2(new_n1023_), .B(pi129), .ZN(po103));
  NAND2_X1   g736(.A1(new_n1022_), .A2(pi140), .ZN(new_n1027_));
  NAND2_X1   g737(.A1(new_n1024_), .A2(pi089), .ZN(new_n1028_));
  AOI21_X1   g738(.A1(new_n1028_), .A2(new_n1027_), .B(pi129), .ZN(po104));
  NAND2_X1   g739(.A1(new_n1022_), .A2(pi142), .ZN(new_n1030_));
  NAND2_X1   g740(.A1(new_n1024_), .A2(pi090), .ZN(new_n1031_));
  AOI21_X1   g741(.A1(new_n1031_), .A2(new_n1030_), .B(pi129), .ZN(po105));
  NAND2_X1   g742(.A1(new_n1022_), .A2(pi143), .ZN(new_n1033_));
  NAND2_X1   g743(.A1(new_n1024_), .A2(pi091), .ZN(new_n1034_));
  AOI21_X1   g744(.A1(new_n1034_), .A2(new_n1033_), .B(pi129), .ZN(po106));
  NAND2_X1   g745(.A1(new_n1022_), .A2(pi144), .ZN(new_n1036_));
  NAND2_X1   g746(.A1(new_n1024_), .A2(pi092), .ZN(new_n1037_));
  AOI21_X1   g747(.A1(new_n1037_), .A2(new_n1036_), .B(pi129), .ZN(po107));
  NAND2_X1   g748(.A1(new_n1022_), .A2(pi146), .ZN(new_n1039_));
  NAND2_X1   g749(.A1(new_n1024_), .A2(pi093), .ZN(new_n1040_));
  AOI21_X1   g750(.A1(new_n1040_), .A2(new_n1039_), .B(pi129), .ZN(po108));
  NAND3_X1   g751(.A1(new_n934_), .A2(pi082), .A3(pi138), .ZN(new_n1042_));
  NOR2_X1    g752(.A1(new_n1042_), .A2(new_n915_), .ZN(new_n1043_));
  NAND2_X1   g753(.A1(new_n1043_), .A2(pi142), .ZN(new_n1044_));
  OAI21_X1   g754(.A1(new_n1042_), .A2(new_n915_), .B(pi094), .ZN(new_n1045_));
  AOI21_X1   g755(.A1(new_n1044_), .A2(new_n1045_), .B(pi129), .ZN(po109));
  INV_X1     g756(.I(pi003), .ZN(new_n1047_));
  INV_X1     g757(.I(new_n915_), .ZN(new_n1048_));
  AOI21_X1   g758(.A1(new_n1047_), .A2(new_n579_), .B(new_n1048_), .ZN(new_n1049_));
  NOR2_X1    g759(.A1(new_n1049_), .A2(new_n1043_), .ZN(new_n1050_));
  AOI22_X1   g760(.A1(new_n1050_), .A2(pi095), .B1(pi143), .B2(new_n1043_), .ZN(new_n1051_));
  NOR2_X1    g761(.A1(new_n1051_), .A2(pi129), .ZN(po110));
  AOI22_X1   g762(.A1(new_n1050_), .A2(pi096), .B1(pi146), .B2(new_n1043_), .ZN(new_n1053_));
  NOR2_X1    g763(.A1(new_n1053_), .A2(pi129), .ZN(po111));
  AOI22_X1   g764(.A1(new_n1050_), .A2(pi097), .B1(pi145), .B2(new_n1043_), .ZN(new_n1055_));
  NOR2_X1    g765(.A1(new_n1055_), .A2(pi129), .ZN(po112));
  NAND2_X1   g766(.A1(new_n1022_), .A2(pi145), .ZN(new_n1057_));
  NAND2_X1   g767(.A1(new_n1024_), .A2(pi098), .ZN(new_n1058_));
  AOI21_X1   g768(.A1(new_n1058_), .A2(new_n1057_), .B(pi129), .ZN(po113));
  NAND2_X1   g769(.A1(new_n1022_), .A2(pi141), .ZN(new_n1060_));
  NAND2_X1   g770(.A1(new_n1024_), .A2(pi099), .ZN(new_n1061_));
  AOI21_X1   g771(.A1(new_n1061_), .A2(new_n1060_), .B(pi129), .ZN(po114));
  AOI22_X1   g772(.A1(new_n1050_), .A2(pi100), .B1(pi144), .B2(new_n1043_), .ZN(new_n1063_));
  NOR2_X1    g773(.A1(new_n1063_), .A2(pi129), .ZN(po115));
  NOR2_X1    g774(.A1(pi082), .A2(pi138), .ZN(new_n1065_));
  AOI21_X1   g775(.A1(new_n611_), .A2(pi138), .B(new_n1065_), .ZN(new_n1066_));
  NOR2_X1    g776(.A1(new_n716_), .A2(new_n917_), .ZN(new_n1067_));
  AOI22_X1   g777(.A1(new_n1066_), .A2(new_n917_), .B1(new_n996_), .B2(new_n1067_), .ZN(new_n1068_));
  AND2_X2    g778(.A1(pi124), .A2(pi138), .Z(new_n1069_));
  NOR2_X1    g779(.A1(pi077), .A2(pi138), .ZN(new_n1070_));
  OAI21_X1   g780(.A1(new_n1069_), .A2(new_n1070_), .B(new_n917_), .ZN(new_n1071_));
  NAND2_X1   g781(.A1(pi093), .A2(pi138), .ZN(new_n1072_));
  OAI21_X1   g782(.A1(pi065), .A2(pi138), .B(new_n1072_), .ZN(new_n1073_));
  AOI21_X1   g783(.A1(new_n1073_), .A2(pi136), .B(pi137), .ZN(new_n1074_));
  AOI22_X1   g784(.A1(new_n1068_), .A2(pi137), .B1(new_n1074_), .B2(new_n1071_), .ZN(po116));
  AOI22_X1   g785(.A1(pi091), .A2(new_n918_), .B1(new_n977_), .B2(pi095), .ZN(new_n1076_));
  NOR2_X1    g786(.A1(new_n698_), .A2(new_n917_), .ZN(new_n1077_));
  INV_X1     g787(.I(pi079), .ZN(new_n1078_));
  NOR2_X1    g788(.A1(new_n1078_), .A2(pi136), .ZN(new_n1079_));
  OAI21_X1   g789(.A1(new_n1077_), .A2(new_n1079_), .B(pi137), .ZN(new_n1080_));
  NAND2_X1   g790(.A1(new_n833_), .A2(pi136), .ZN(new_n1081_));
  OAI21_X1   g791(.A1(pi066), .A2(pi136), .B(new_n1081_), .ZN(new_n1082_));
  AOI21_X1   g792(.A1(new_n1082_), .A2(new_n976_), .B(pi138), .ZN(new_n1083_));
  AOI22_X1   g793(.A1(new_n1083_), .A2(new_n1080_), .B1(pi138), .B2(new_n1076_), .ZN(po117));
  AOI22_X1   g794(.A1(pi090), .A2(new_n918_), .B1(new_n977_), .B2(pi094), .ZN(new_n1085_));
  NOR2_X1    g795(.A1(new_n692_), .A2(new_n917_), .ZN(new_n1086_));
  INV_X1     g796(.I(pi078), .ZN(new_n1087_));
  NOR2_X1    g797(.A1(new_n1087_), .A2(pi136), .ZN(new_n1088_));
  OAI21_X1   g798(.A1(new_n1086_), .A2(new_n1088_), .B(pi137), .ZN(new_n1089_));
  NAND2_X1   g799(.A1(new_n553_), .A2(pi136), .ZN(new_n1090_));
  OAI21_X1   g800(.A1(pi074), .A2(pi136), .B(new_n1090_), .ZN(new_n1091_));
  AOI21_X1   g801(.A1(new_n1091_), .A2(new_n976_), .B(pi138), .ZN(new_n1092_));
  AOI22_X1   g802(.A1(new_n1092_), .A2(new_n1089_), .B1(pi138), .B2(new_n1085_), .ZN(po118));
  INV_X1     g803(.I(pi112), .ZN(new_n1094_));
  AOI22_X1   g804(.A1(pi099), .A2(new_n918_), .B1(new_n977_), .B2(new_n1094_), .ZN(new_n1095_));
  NOR2_X1    g805(.A1(new_n917_), .A2(pi068), .ZN(new_n1096_));
  NOR2_X1    g806(.A1(pi073), .A2(pi136), .ZN(new_n1097_));
  OAI21_X1   g807(.A1(new_n1096_), .A2(new_n1097_), .B(new_n976_), .ZN(new_n1098_));
  NAND2_X1   g808(.A1(new_n917_), .A2(pi084), .ZN(new_n1099_));
  OAI21_X1   g809(.A1(new_n686_), .A2(new_n917_), .B(new_n1099_), .ZN(new_n1100_));
  AOI21_X1   g810(.A1(new_n1100_), .A2(pi137), .B(pi138), .ZN(new_n1101_));
  AOI22_X1   g811(.A1(new_n1101_), .A2(new_n1098_), .B1(new_n1095_), .B2(pi138), .ZN(po119));
  NOR2_X1    g812(.A1(pi080), .A2(pi138), .ZN(new_n1103_));
  AOI21_X1   g813(.A1(new_n617_), .A2(pi138), .B(new_n1103_), .ZN(new_n1104_));
  NOR2_X1    g814(.A1(new_n704_), .A2(new_n917_), .ZN(new_n1105_));
  AOI22_X1   g815(.A1(new_n1104_), .A2(new_n917_), .B1(new_n996_), .B2(new_n1105_), .ZN(new_n1106_));
  AND2_X2    g816(.A1(pi092), .A2(pi138), .Z(new_n1107_));
  NOR2_X1    g817(.A1(pi070), .A2(pi138), .ZN(new_n1108_));
  OAI21_X1   g818(.A1(new_n1107_), .A2(new_n1108_), .B(pi136), .ZN(new_n1109_));
  NAND2_X1   g819(.A1(pi125), .A2(pi138), .ZN(new_n1110_));
  OAI21_X1   g820(.A1(pi075), .A2(pi138), .B(new_n1110_), .ZN(new_n1111_));
  AOI21_X1   g821(.A1(new_n1111_), .A2(new_n917_), .B(pi137), .ZN(new_n1112_));
  AOI22_X1   g822(.A1(new_n1106_), .A2(pi137), .B1(new_n1112_), .B2(new_n1109_), .ZN(po120));
  NAND3_X1   g823(.A1(new_n1013_), .A2(new_n604_), .A3(new_n895_), .ZN(new_n1114_));
  AOI21_X1   g824(.A1(new_n1114_), .A2(new_n609_), .B(new_n418_), .ZN(po121));
  NOR2_X1    g825(.A1(pi081), .A2(pi138), .ZN(new_n1116_));
  AOI21_X1   g826(.A1(new_n656_), .A2(pi138), .B(new_n1116_), .ZN(new_n1117_));
  NOR2_X1    g827(.A1(new_n710_), .A2(new_n917_), .ZN(new_n1118_));
  AOI22_X1   g828(.A1(new_n1117_), .A2(new_n917_), .B1(new_n996_), .B2(new_n1118_), .ZN(new_n1119_));
  AND2_X2    g829(.A1(pi098), .A2(pi138), .Z(new_n1120_));
  NOR2_X1    g830(.A1(pi071), .A2(pi138), .ZN(new_n1121_));
  OAI21_X1   g831(.A1(new_n1120_), .A2(new_n1121_), .B(pi136), .ZN(new_n1122_));
  NAND2_X1   g832(.A1(pi023), .A2(pi138), .ZN(new_n1123_));
  OAI21_X1   g833(.A1(pi076), .A2(pi138), .B(new_n1123_), .ZN(new_n1124_));
  AOI21_X1   g834(.A1(new_n1124_), .A2(new_n917_), .B(pi137), .ZN(new_n1125_));
  AOI22_X1   g835(.A1(new_n1119_), .A2(pi137), .B1(new_n1125_), .B2(new_n1122_), .ZN(po122));
  NOR2_X1    g836(.A1(pi086), .A2(pi138), .ZN(new_n1127_));
  NOR2_X1    g837(.A1(new_n996_), .A2(pi111), .ZN(new_n1128_));
  NOR2_X1    g838(.A1(new_n1128_), .A2(new_n1127_), .ZN(new_n1129_));
  NOR2_X1    g839(.A1(new_n681_), .A2(new_n917_), .ZN(new_n1130_));
  AOI22_X1   g840(.A1(new_n1129_), .A2(new_n917_), .B1(new_n996_), .B2(new_n1130_), .ZN(new_n1131_));
  AND2_X2    g841(.A1(pi088), .A2(pi138), .Z(new_n1132_));
  NOR2_X1    g842(.A1(pi064), .A2(pi138), .ZN(new_n1133_));
  OAI21_X1   g843(.A1(new_n1132_), .A2(new_n1133_), .B(pi136), .ZN(new_n1134_));
  NAND2_X1   g844(.A1(pi120), .A2(pi138), .ZN(new_n1135_));
  OAI21_X1   g845(.A1(pi067), .A2(pi138), .B(new_n1135_), .ZN(new_n1136_));
  AOI21_X1   g846(.A1(new_n1136_), .A2(new_n917_), .B(pi137), .ZN(new_n1137_));
  AOI22_X1   g847(.A1(new_n1131_), .A2(pi137), .B1(new_n1134_), .B2(new_n1137_), .ZN(po123));
  NAND2_X1   g848(.A1(new_n291_), .A2(pi116), .ZN(new_n1139_));
  OAI21_X1   g849(.A1(new_n638_), .A2(new_n591_), .B(new_n631_), .ZN(new_n1140_));
  NOR2_X1    g850(.A1(new_n1140_), .A2(new_n1139_), .ZN(po124));
  NAND2_X1   g851(.A1(new_n627_), .A2(new_n656_), .ZN(new_n1142_));
  AOI21_X1   g852(.A1(new_n1142_), .A2(new_n600_), .B(new_n1139_), .ZN(po125));
  NAND2_X1   g853(.A1(new_n1048_), .A2(new_n792_), .ZN(new_n1144_));
  INV_X1     g854(.I(new_n1042_), .ZN(new_n1145_));
  NAND2_X1   g855(.A1(new_n1145_), .A2(pi139), .ZN(new_n1146_));
  NAND2_X1   g856(.A1(new_n1042_), .A2(pi111), .ZN(new_n1147_));
  AOI21_X1   g857(.A1(new_n1146_), .A2(new_n1147_), .B(new_n1144_), .ZN(po126));
  NAND2_X1   g858(.A1(new_n1145_), .A2(pi141), .ZN(new_n1149_));
  NAND2_X1   g859(.A1(new_n1042_), .A2(new_n1094_), .ZN(new_n1150_));
  AOI21_X1   g860(.A1(new_n1149_), .A2(new_n1150_), .B(new_n1144_), .ZN(po127));
  NOR2_X1    g861(.A1(new_n408_), .A2(pi054), .ZN(new_n1152_));
  NOR3_X1    g862(.A1(new_n292_), .A2(pi011), .A3(pi022), .ZN(new_n1153_));
  NOR3_X1    g863(.A1(new_n1153_), .A2(new_n418_), .A3(new_n1152_), .ZN(po128));
  NAND2_X1   g864(.A1(new_n1145_), .A2(pi140), .ZN(new_n1155_));
  NAND2_X1   g865(.A1(new_n1042_), .A2(new_n995_), .ZN(new_n1156_));
  AOI21_X1   g866(.A1(new_n1155_), .A2(new_n1156_), .B(new_n1144_), .ZN(po130));
  NOR4_X1    g867(.A1(pi004), .A2(pi007), .A3(pi009), .A4(pi012), .ZN(new_n1158_));
  NOR3_X1    g868(.A1(new_n418_), .A2(new_n1158_), .A3(new_n292_), .ZN(po131));
  NAND2_X1   g869(.A1(new_n792_), .A2(pi122), .ZN(po132));
  NAND2_X1   g870(.A1(new_n292_), .A2(pi118), .ZN(new_n1161_));
  NAND3_X1   g871(.A1(new_n480_), .A2(pi054), .A3(new_n513_), .ZN(new_n1162_));
  AOI21_X1   g872(.A1(new_n1162_), .A2(new_n1161_), .B(pi129), .ZN(po133));
  NOR2_X1    g873(.A1(new_n859_), .A2(pi129), .ZN(po134));
  NOR3_X1    g874(.A1(pi003), .A2(pi110), .A3(pi120), .ZN(new_n1165_));
  NOR3_X1    g875(.A1(new_n1165_), .A2(pi111), .A3(pi129), .ZN(po135));
  AND3_X2    g876(.A1(new_n792_), .A2(pi081), .A3(pi120), .Z(po136));
  OR2_X2     g877(.A1(pi129), .A2(pi134), .Z(po137));
  OR2_X2     g878(.A1(pi129), .A2(pi135), .Z(po138));
  NOR2_X1    g879(.A1(new_n885_), .A2(pi129), .ZN(po139));
  NAND2_X1   g880(.A1(new_n611_), .A2(pi125), .ZN(new_n1171_));
  AOI21_X1   g881(.A1(new_n1171_), .A2(new_n1047_), .B(pi129), .ZN(po140));
  INV_X1     g882(.I(pi126), .ZN(new_n1173_));
  AND3_X2    g883(.A1(new_n1173_), .A2(pi132), .A3(pi133), .Z(po141));
  assign     po012 = 1'b1;
  BUF_X16    g884(.I(pi108), .Z(po000));
  BUF_X16    g885(.I(pi083), .Z(po001));
  BUF_X16    g886(.I(pi104), .Z(po002));
  BUF_X16    g887(.I(pi103), .Z(po003));
  BUF_X16    g888(.I(pi102), .Z(po004));
  BUF_X16    g889(.I(pi105), .Z(po005));
  BUF_X16    g890(.I(pi107), .Z(po006));
  BUF_X16    g891(.I(pi101), .Z(po007));
  BUF_X16    g892(.I(pi126), .Z(po008));
  BUF_X16    g893(.I(pi121), .Z(po009));
  BUF_X16    g894(.I(pi001), .Z(po010));
  BUF_X16    g895(.I(pi000), .Z(po011));
  BUF_X16    g896(.I(pi130), .Z(po013));
  BUF_X16    g897(.I(pi128), .Z(po014));
endmodule


