// Benchmark "ADDERFDS" written by ABC on Fri Feb 25 15:13:04 2022

module my_adder ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, b0, c0, d0, e0, f0, g0,
    h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0;
  output h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0;
  wire new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_,
    new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_,
    new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n225_;
  assign new_n51_ = ~f0 & ~g0;
  assign new_n52_ = f0 & g0;
  assign new_n53_ = ~p & ~new_n52_;
  assign new_n54_ = ~new_n51_ & ~new_n53_;
  assign new_n55_ = ~e0 & ~new_n54_;
  assign new_n56_ = e0 & new_n54_;
  assign new_n57_ = ~o & ~new_n56_;
  assign new_n58_ = ~new_n55_ & ~new_n57_;
  assign new_n59_ = ~d0 & ~new_n58_;
  assign new_n60_ = d0 & new_n58_;
  assign new_n61_ = ~n & ~new_n60_;
  assign new_n62_ = ~new_n59_ & ~new_n61_;
  assign new_n63_ = ~c0 & ~new_n62_;
  assign new_n64_ = c0 & new_n62_;
  assign new_n65_ = ~m & ~new_n64_;
  assign new_n66_ = ~new_n63_ & ~new_n65_;
  assign new_n67_ = ~b0 & ~new_n66_;
  assign new_n68_ = b0 & new_n66_;
  assign new_n69_ = ~l & ~new_n68_;
  assign new_n70_ = ~new_n67_ & ~new_n69_;
  assign new_n71_ = ~a0 & ~new_n70_;
  assign new_n72_ = a0 & new_n70_;
  assign new_n73_ = ~k & ~new_n72_;
  assign new_n74_ = ~new_n71_ & ~new_n73_;
  assign new_n75_ = ~z & ~new_n74_;
  assign new_n76_ = z & new_n74_;
  assign new_n77_ = ~j & ~new_n76_;
  assign new_n78_ = ~new_n75_ & ~new_n77_;
  assign new_n79_ = ~y & ~new_n78_;
  assign new_n80_ = y & new_n78_;
  assign new_n81_ = ~i & ~new_n80_;
  assign new_n82_ = ~new_n79_ & ~new_n81_;
  assign new_n83_ = ~x & ~new_n82_;
  assign new_n84_ = x & new_n82_;
  assign new_n85_ = ~h & ~new_n84_;
  assign new_n86_ = ~new_n83_ & ~new_n85_;
  assign new_n87_ = ~w & ~new_n86_;
  assign new_n88_ = w & new_n86_;
  assign new_n89_ = ~g & ~new_n88_;
  assign new_n90_ = ~new_n87_ & ~new_n89_;
  assign new_n91_ = ~v & ~new_n90_;
  assign new_n92_ = v & new_n90_;
  assign new_n93_ = ~f & ~new_n92_;
  assign new_n94_ = ~new_n91_ & ~new_n93_;
  assign new_n95_ = ~u & ~new_n94_;
  assign new_n96_ = u & new_n94_;
  assign new_n97_ = ~e & ~new_n96_;
  assign new_n98_ = ~new_n95_ & ~new_n97_;
  assign new_n99_ = ~t & ~new_n98_;
  assign new_n100_ = t & new_n98_;
  assign new_n101_ = ~d & ~new_n100_;
  assign new_n102_ = ~new_n99_ & ~new_n101_;
  assign new_n103_ = ~s & ~new_n102_;
  assign new_n104_ = s & new_n102_;
  assign new_n105_ = ~c & ~new_n104_;
  assign new_n106_ = ~new_n103_ & ~new_n105_;
  assign new_n107_ = ~r & ~new_n106_;
  assign new_n108_ = r & new_n106_;
  assign new_n109_ = ~b & ~new_n108_;
  assign new_n110_ = ~new_n107_ & ~new_n109_;
  assign new_n111_ = q & ~new_n110_;
  assign new_n112_ = ~q & new_n110_;
  assign new_n113_ = ~new_n111_ & ~new_n112_;
  assign new_n114_ = a & ~new_n113_;
  assign new_n115_ = ~q & ~new_n110_;
  assign new_n116_ = q & new_n110_;
  assign new_n117_ = ~new_n115_ & ~new_n116_;
  assign new_n118_ = ~a & ~new_n117_;
  assign h0 = ~new_n114_ & ~new_n118_;
  assign new_n120_ = r & ~new_n106_;
  assign new_n121_ = ~r & new_n106_;
  assign new_n122_ = ~new_n120_ & ~new_n121_;
  assign new_n123_ = b & ~new_n122_;
  assign new_n124_ = ~new_n107_ & ~new_n108_;
  assign new_n125_ = ~b & ~new_n124_;
  assign i0 = ~new_n123_ & ~new_n125_;
  assign new_n127_ = s & ~new_n102_;
  assign new_n128_ = ~s & new_n102_;
  assign new_n129_ = ~new_n127_ & ~new_n128_;
  assign new_n130_ = c & ~new_n129_;
  assign new_n131_ = ~new_n103_ & ~new_n104_;
  assign new_n132_ = ~c & ~new_n131_;
  assign j0 = ~new_n130_ & ~new_n132_;
  assign new_n134_ = t & ~new_n98_;
  assign new_n135_ = ~t & new_n98_;
  assign new_n136_ = ~new_n134_ & ~new_n135_;
  assign new_n137_ = d & ~new_n136_;
  assign new_n138_ = ~new_n99_ & ~new_n100_;
  assign new_n139_ = ~d & ~new_n138_;
  assign k0 = ~new_n137_ & ~new_n139_;
  assign new_n141_ = u & ~new_n94_;
  assign new_n142_ = ~u & new_n94_;
  assign new_n143_ = ~new_n141_ & ~new_n142_;
  assign new_n144_ = e & ~new_n143_;
  assign new_n145_ = ~new_n95_ & ~new_n96_;
  assign new_n146_ = ~e & ~new_n145_;
  assign l0 = ~new_n144_ & ~new_n146_;
  assign new_n148_ = v & ~new_n90_;
  assign new_n149_ = ~v & new_n90_;
  assign new_n150_ = ~new_n148_ & ~new_n149_;
  assign new_n151_ = f & ~new_n150_;
  assign new_n152_ = ~new_n91_ & ~new_n92_;
  assign new_n153_ = ~f & ~new_n152_;
  assign m0 = ~new_n151_ & ~new_n153_;
  assign new_n155_ = w & ~new_n86_;
  assign new_n156_ = ~w & new_n86_;
  assign new_n157_ = ~new_n155_ & ~new_n156_;
  assign new_n158_ = g & ~new_n157_;
  assign new_n159_ = ~new_n87_ & ~new_n88_;
  assign new_n160_ = ~g & ~new_n159_;
  assign n0 = ~new_n158_ & ~new_n160_;
  assign new_n162_ = x & ~new_n82_;
  assign new_n163_ = ~x & new_n82_;
  assign new_n164_ = ~new_n162_ & ~new_n163_;
  assign new_n165_ = h & ~new_n164_;
  assign new_n166_ = ~new_n83_ & ~new_n84_;
  assign new_n167_ = ~h & ~new_n166_;
  assign o0 = ~new_n165_ & ~new_n167_;
  assign new_n169_ = y & ~new_n78_;
  assign new_n170_ = ~y & new_n78_;
  assign new_n171_ = ~new_n169_ & ~new_n170_;
  assign new_n172_ = i & ~new_n171_;
  assign new_n173_ = ~new_n79_ & ~new_n80_;
  assign new_n174_ = ~i & ~new_n173_;
  assign p0 = ~new_n172_ & ~new_n174_;
  assign new_n176_ = z & ~new_n74_;
  assign new_n177_ = ~z & new_n74_;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign new_n179_ = j & ~new_n178_;
  assign new_n180_ = ~new_n75_ & ~new_n76_;
  assign new_n181_ = ~j & ~new_n180_;
  assign q0 = ~new_n179_ & ~new_n181_;
  assign new_n183_ = a0 & ~new_n70_;
  assign new_n184_ = ~a0 & new_n70_;
  assign new_n185_ = ~new_n183_ & ~new_n184_;
  assign new_n186_ = k & ~new_n185_;
  assign new_n187_ = ~new_n71_ & ~new_n72_;
  assign new_n188_ = ~k & ~new_n187_;
  assign r0 = ~new_n186_ & ~new_n188_;
  assign new_n190_ = b0 & ~new_n66_;
  assign new_n191_ = ~b0 & new_n66_;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign new_n193_ = l & ~new_n192_;
  assign new_n194_ = ~new_n67_ & ~new_n68_;
  assign new_n195_ = ~l & ~new_n194_;
  assign s0 = ~new_n193_ & ~new_n195_;
  assign new_n197_ = c0 & ~new_n62_;
  assign new_n198_ = ~c0 & new_n62_;
  assign new_n199_ = ~new_n197_ & ~new_n198_;
  assign new_n200_ = m & ~new_n199_;
  assign new_n201_ = ~new_n63_ & ~new_n64_;
  assign new_n202_ = ~m & ~new_n201_;
  assign t0 = ~new_n200_ & ~new_n202_;
  assign new_n204_ = d0 & ~new_n58_;
  assign new_n205_ = ~d0 & new_n58_;
  assign new_n206_ = ~new_n204_ & ~new_n205_;
  assign new_n207_ = n & ~new_n206_;
  assign new_n208_ = ~new_n59_ & ~new_n60_;
  assign new_n209_ = ~n & ~new_n208_;
  assign u0 = ~new_n207_ & ~new_n209_;
  assign new_n211_ = e0 & ~new_n54_;
  assign new_n212_ = ~e0 & new_n54_;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = o & ~new_n213_;
  assign new_n215_ = ~new_n55_ & ~new_n56_;
  assign new_n216_ = ~o & ~new_n215_;
  assign v0 = ~new_n214_ & ~new_n216_;
  assign new_n218_ = ~f0 & g0;
  assign new_n219_ = f0 & ~g0;
  assign new_n220_ = ~new_n218_ & ~new_n219_;
  assign new_n221_ = p & ~new_n220_;
  assign new_n222_ = ~new_n51_ & ~new_n52_;
  assign new_n223_ = ~p & ~new_n222_;
  assign w0 = ~new_n221_ & ~new_n223_;
  assign new_n225_ = ~a & ~new_n116_;
  assign x0 = ~new_n115_ & ~new_n225_;
endmodule


