// Benchmark "sqrt" written by ABC on Thu Sep 14 20:29:38 2023

module sqrt ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] ,
    \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] , \asqrt[5] ,
    \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] , \asqrt[10] ,
    \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] , \asqrt[15] ,
    \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] , \asqrt[20] ,
    \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] , \asqrt[25] ,
    \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] , \asqrt[30] ,
    \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] , \asqrt[35] ,
    \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] , \asqrt[40] ,
    \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] , \asqrt[45] ,
    \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] , \asqrt[50] ,
    \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] , \asqrt[55] ,
    \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] , \asqrt[60] ,
    \asqrt[61] , \asqrt[62] , \asqrt[63]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] ;
  output \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] ,
    \asqrt[5] , \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] ,
    \asqrt[10] , \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] ,
    \asqrt[15] , \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] ,
    \asqrt[20] , \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] ,
    \asqrt[25] , \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] ,
    \asqrt[30] , \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] ,
    \asqrt[35] , \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] ,
    \asqrt[40] , \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] ,
    \asqrt[45] , \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] ,
    \asqrt[50] , \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] ,
    \asqrt[55] , \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] ,
    \asqrt[60] , \asqrt[61] , \asqrt[62] , \asqrt[63] ;
  wire new_n193_, new_n194_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1821_,
    new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_,
    new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_,
    new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_,
    new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_,
    new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_,
    new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_,
    new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_,
    new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_,
    new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_,
    new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_,
    new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_,
    new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_,
    new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_,
    new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_,
    new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_,
    new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_,
    new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_,
    new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_,
    new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_,
    new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_,
    new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_,
    new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_,
    new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_,
    new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_,
    new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_,
    new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_,
    new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_,
    new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_,
    new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_,
    new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_,
    new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_,
    new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_,
    new_n2954_, new_n2955_, new_n2957_, new_n2958_, new_n2959_, new_n2960_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_,
    new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_,
    new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_,
    new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_,
    new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_,
    new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_,
    new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_,
    new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_,
    new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_,
    new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_,
    new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_,
    new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_,
    new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_,
    new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_,
    new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_,
    new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_,
    new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_,
    new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_,
    new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_,
    new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_,
    new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_,
    new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3440_, new_n3441_, new_n3442_,
    new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_,
    new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_,
    new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_,
    new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_,
    new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_,
    new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_,
    new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_,
    new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_,
    new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_,
    new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_,
    new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_,
    new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_,
    new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_,
    new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_,
    new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_,
    new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_,
    new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_,
    new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_,
    new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_,
    new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_,
    new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_,
    new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_,
    new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_,
    new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_,
    new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_,
    new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_,
    new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_,
    new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_,
    new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_,
    new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_,
    new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_,
    new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_,
    new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_,
    new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_,
    new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_,
    new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_,
    new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_,
    new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_,
    new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_,
    new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_,
    new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_,
    new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_,
    new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_,
    new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_,
    new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_,
    new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_,
    new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_,
    new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_,
    new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_,
    new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_,
    new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_,
    new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_,
    new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_,
    new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_,
    new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_,
    new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_,
    new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_,
    new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_,
    new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_,
    new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_,
    new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_,
    new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_,
    new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_,
    new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_,
    new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_,
    new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_,
    new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_,
    new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4604_,
    new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_,
    new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_,
    new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_,
    new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_,
    new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_,
    new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_,
    new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_,
    new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_,
    new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_,
    new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_,
    new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_,
    new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_,
    new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_,
    new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_,
    new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_,
    new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_,
    new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_,
    new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_,
    new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_,
    new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_,
    new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_,
    new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_,
    new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_,
    new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_,
    new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_,
    new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_,
    new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_,
    new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_,
    new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_,
    new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_,
    new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_,
    new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_,
    new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_,
    new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_,
    new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_,
    new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_,
    new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_,
    new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_,
    new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_,
    new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_,
    new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_,
    new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_,
    new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_,
    new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_,
    new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_,
    new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_,
    new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_,
    new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_,
    new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_,
    new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_,
    new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_,
    new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_,
    new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_,
    new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_,
    new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_,
    new_n4935_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_,
    new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_,
    new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_,
    new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_,
    new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_,
    new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_,
    new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_,
    new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_,
    new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_,
    new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_,
    new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_,
    new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_,
    new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_,
    new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_,
    new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_,
    new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_,
    new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_,
    new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_,
    new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_,
    new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_,
    new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_,
    new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_,
    new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_,
    new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_,
    new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_,
    new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_,
    new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_,
    new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_,
    new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_,
    new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_,
    new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_,
    new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_,
    new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_,
    new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_,
    new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_,
    new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_,
    new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_,
    new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_,
    new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_,
    new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_,
    new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_,
    new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_,
    new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_,
    new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_,
    new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_,
    new_n5284_, new_n5285_, new_n5287_, new_n5288_, new_n5289_, new_n5290_,
    new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_,
    new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_,
    new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_,
    new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_,
    new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_,
    new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_,
    new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_,
    new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_,
    new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_,
    new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_,
    new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_,
    new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_,
    new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_,
    new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_,
    new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_,
    new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_,
    new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_,
    new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_,
    new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_,
    new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_,
    new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_,
    new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_,
    new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_,
    new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_,
    new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_,
    new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_,
    new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_,
    new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_,
    new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_,
    new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_,
    new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_,
    new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_,
    new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_,
    new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_,
    new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_,
    new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_,
    new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_,
    new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_,
    new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_,
    new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_,
    new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_,
    new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_,
    new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_,
    new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_,
    new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_,
    new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_,
    new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_,
    new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_,
    new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_,
    new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5590_, new_n5591_,
    new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_,
    new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_,
    new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_,
    new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_,
    new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_,
    new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_,
    new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_,
    new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_,
    new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_,
    new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_,
    new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_,
    new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5950_, new_n5951_, new_n5952_,
    new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_,
    new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_,
    new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_,
    new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_,
    new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_,
    new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_,
    new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_,
    new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_,
    new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_,
    new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_,
    new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_,
    new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_,
    new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_,
    new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_,
    new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_,
    new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_,
    new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_,
    new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_,
    new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_,
    new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_,
    new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_,
    new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_,
    new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_,
    new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_,
    new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_,
    new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_,
    new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_,
    new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_,
    new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_,
    new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_,
    new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_,
    new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_,
    new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_,
    new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_,
    new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_,
    new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_,
    new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_,
    new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_,
    new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_,
    new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_,
    new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_,
    new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_,
    new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_,
    new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_,
    new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_,
    new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_,
    new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_,
    new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_,
    new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_,
    new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_,
    new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_,
    new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_,
    new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_,
    new_n6325_, new_n6326_, new_n6327_, new_n6329_, new_n6330_, new_n6331_,
    new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_,
    new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_,
    new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_,
    new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_,
    new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_,
    new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_,
    new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_,
    new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_,
    new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_,
    new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_,
    new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_,
    new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_,
    new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_,
    new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_,
    new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_,
    new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_,
    new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_,
    new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_,
    new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_,
    new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_,
    new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_,
    new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_,
    new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_,
    new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_,
    new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_,
    new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_,
    new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_,
    new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_,
    new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_,
    new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_,
    new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_,
    new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_,
    new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_,
    new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_,
    new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_,
    new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_,
    new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_,
    new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_,
    new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_,
    new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_,
    new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_,
    new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_,
    new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_,
    new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_,
    new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_,
    new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_,
    new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_,
    new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_,
    new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_,
    new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_,
    new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_,
    new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_,
    new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_,
    new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_,
    new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_,
    new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_,
    new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_,
    new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_,
    new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_,
    new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_,
    new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_,
    new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_,
    new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_,
    new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_,
    new_n7071_, new_n7072_, new_n7073_, new_n7075_, new_n7076_, new_n7077_,
    new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_,
    new_n7084_, new_n7085_, new_n7086_, new_n7087_, new_n7088_, new_n7089_,
    new_n7090_, new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_,
    new_n7096_, new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_,
    new_n7102_, new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_,
    new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_,
    new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_,
    new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_,
    new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_, new_n7131_,
    new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_, new_n7137_,
    new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_, new_n7143_,
    new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_, new_n7149_,
    new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_, new_n7155_,
    new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_, new_n7161_,
    new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_, new_n7167_,
    new_n7168_, new_n7169_, new_n7170_, new_n7171_, new_n7172_, new_n7173_,
    new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_, new_n7179_,
    new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_, new_n7185_,
    new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_, new_n7191_,
    new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_, new_n7197_,
    new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_,
    new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_, new_n7209_,
    new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_, new_n7215_,
    new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_, new_n7221_,
    new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_, new_n7227_,
    new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_, new_n7233_,
    new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_, new_n7239_,
    new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_, new_n7245_,
    new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_,
    new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_,
    new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_,
    new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_,
    new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_,
    new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_, new_n7281_,
    new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_, new_n7287_,
    new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_, new_n7293_,
    new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_, new_n7299_,
    new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_, new_n7305_,
    new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_, new_n7311_,
    new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_, new_n7317_,
    new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_, new_n7323_,
    new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_,
    new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_,
    new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7476_, new_n7477_, new_n7478_, new_n7479_, new_n7480_,
    new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_, new_n7486_,
    new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_, new_n7492_,
    new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_, new_n7498_,
    new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_, new_n7504_,
    new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_, new_n7510_,
    new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_, new_n7516_,
    new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_, new_n7522_,
    new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_, new_n7528_,
    new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_, new_n7534_,
    new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_, new_n7540_,
    new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_, new_n7546_,
    new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_,
    new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_,
    new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_,
    new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_,
    new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_,
    new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_,
    new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_,
    new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_,
    new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_,
    new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_,
    new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_,
    new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_,
    new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_,
    new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_,
    new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_,
    new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_,
    new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_,
    new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_,
    new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_,
    new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_,
    new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_,
    new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_,
    new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_,
    new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_,
    new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_,
    new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_,
    new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_,
    new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_,
    new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_,
    new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_,
    new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_,
    new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_,
    new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_,
    new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_,
    new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_,
    new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_,
    new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_,
    new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_,
    new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_,
    new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_,
    new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_,
    new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_,
    new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_,
    new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_,
    new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_,
    new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_,
    new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_,
    new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_,
    new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_,
    new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_,
    new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_,
    new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_,
    new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_,
    new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_,
    new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_,
    new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_,
    new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_,
    new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7895_,
    new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_,
    new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_,
    new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_,
    new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_,
    new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_,
    new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_,
    new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_,
    new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_,
    new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_,
    new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_,
    new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_,
    new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_,
    new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_,
    new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_,
    new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_,
    new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_,
    new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_,
    new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_,
    new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_,
    new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_,
    new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_,
    new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_,
    new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_,
    new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_,
    new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_,
    new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_,
    new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_,
    new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_,
    new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_,
    new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_,
    new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_,
    new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_,
    new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_,
    new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_,
    new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_,
    new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_,
    new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_,
    new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_,
    new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_,
    new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_,
    new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_,
    new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_,
    new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_,
    new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_,
    new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_,
    new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_,
    new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_,
    new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_,
    new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_,
    new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_,
    new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_,
    new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_,
    new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_,
    new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_,
    new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_,
    new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_,
    new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_,
    new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_,
    new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_,
    new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_,
    new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_,
    new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_,
    new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_,
    new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_,
    new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_,
    new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_,
    new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_,
    new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_,
    new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_,
    new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_,
    new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_,
    new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_,
    new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_,
    new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_,
    new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_,
    new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_,
    new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_,
    new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_,
    new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_,
    new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_,
    new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_,
    new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_,
    new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_,
    new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_,
    new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_,
    new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_,
    new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_,
    new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_,
    new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_,
    new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_,
    new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_,
    new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_,
    new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_,
    new_n8725_, new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_,
    new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_,
    new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_,
    new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_,
    new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_,
    new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_,
    new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_, new_n8767_,
    new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_,
    new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_,
    new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_,
    new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_,
    new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_,
    new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_,
    new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_,
    new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_, new_n8821_,
    new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_,
    new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_,
    new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_,
    new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_,
    new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_,
    new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_,
    new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_,
    new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_,
    new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_,
    new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_,
    new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_,
    new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_,
    new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_,
    new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_,
    new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_,
    new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_,
    new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_,
    new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_,
    new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_,
    new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_,
    new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_,
    new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_,
    new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_,
    new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_,
    new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_,
    new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_,
    new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_,
    new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_,
    new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_,
    new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_,
    new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_,
    new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_,
    new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_,
    new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_,
    new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_,
    new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_,
    new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_,
    new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_,
    new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_,
    new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_,
    new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_,
    new_n9375_, new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_,
    new_n9381_, new_n9382_, new_n9383_, new_n9384_, new_n9385_, new_n9386_,
    new_n9387_, new_n9388_, new_n9389_, new_n9390_, new_n9391_, new_n9392_,
    new_n9393_, new_n9394_, new_n9395_, new_n9396_, new_n9397_, new_n9398_,
    new_n9399_, new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_,
    new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_,
    new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_, new_n9416_,
    new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_, new_n9422_,
    new_n9423_, new_n9424_, new_n9425_, new_n9426_, new_n9427_, new_n9428_,
    new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_,
    new_n9435_, new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9440_,
    new_n9441_, new_n9442_, new_n9443_, new_n9444_, new_n9445_, new_n9446_,
    new_n9447_, new_n9448_, new_n9449_, new_n9450_, new_n9451_, new_n9452_,
    new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_, new_n9458_,
    new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9463_, new_n9464_,
    new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_,
    new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_,
    new_n9477_, new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_,
    new_n9483_, new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_,
    new_n9489_, new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_,
    new_n9495_, new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_,
    new_n9501_, new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_,
    new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_,
    new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_,
    new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_,
    new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_,
    new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_,
    new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_,
    new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_,
    new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_,
    new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_,
    new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_,
    new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_,
    new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_,
    new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_,
    new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_,
    new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_,
    new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_,
    new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_,
    new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_,
    new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_,
    new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_,
    new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_,
    new_n9633_, new_n9634_, new_n9636_, new_n9637_, new_n9638_, new_n9639_,
    new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_,
    new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_,
    new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_,
    new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_,
    new_n9664_, new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_,
    new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_,
    new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_,
    new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_,
    new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_,
    new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_,
    new_n9700_, new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_,
    new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_,
    new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_,
    new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_,
    new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_,
    new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_,
    new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_,
    new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_,
    new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_,
    new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_,
    new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_,
    new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_,
    new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_,
    new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_,
    new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_,
    new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_,
    new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_,
    new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_,
    new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_,
    new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_,
    new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_,
    new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_,
    new_n9832_, new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_,
    new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_,
    new_n9844_, new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_,
    new_n9850_, new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_,
    new_n9856_, new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_,
    new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_,
    new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_,
    new_n9874_, new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_,
    new_n9880_, new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_,
    new_n9886_, new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_,
    new_n9892_, new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_,
    new_n9898_, new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_,
    new_n9904_, new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_,
    new_n9910_, new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_,
    new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_,
    new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_,
    new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_,
    new_n9934_, new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_,
    new_n9940_, new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_,
    new_n9946_, new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_,
    new_n9952_, new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_,
    new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_,
    new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_,
    new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_,
    new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_,
    new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_,
    new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_,
    new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10202_, new_n10203_, new_n10204_, new_n10205_,
    new_n10206_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10293_, new_n10294_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10301_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10578_, new_n10579_, new_n10580_, new_n10581_,
    new_n10582_, new_n10583_, new_n10584_, new_n10585_, new_n10586_,
    new_n10587_, new_n10588_, new_n10589_, new_n10590_, new_n10591_,
    new_n10592_, new_n10593_, new_n10594_, new_n10595_, new_n10596_,
    new_n10597_, new_n10598_, new_n10599_, new_n10600_, new_n10601_,
    new_n10602_, new_n10603_, new_n10604_, new_n10605_, new_n10606_,
    new_n10607_, new_n10608_, new_n10609_, new_n10610_, new_n10611_,
    new_n10612_, new_n10613_, new_n10614_, new_n10615_, new_n10616_,
    new_n10617_, new_n10618_, new_n10619_, new_n10620_, new_n10621_,
    new_n10622_, new_n10623_, new_n10624_, new_n10625_, new_n10626_,
    new_n10627_, new_n10628_, new_n10629_, new_n10630_, new_n10631_,
    new_n10632_, new_n10633_, new_n10634_, new_n10635_, new_n10636_,
    new_n10637_, new_n10638_, new_n10639_, new_n10640_, new_n10641_,
    new_n10642_, new_n10643_, new_n10644_, new_n10645_, new_n10646_,
    new_n10647_, new_n10648_, new_n10649_, new_n10650_, new_n10651_,
    new_n10652_, new_n10653_, new_n10654_, new_n10655_, new_n10656_,
    new_n10657_, new_n10658_, new_n10659_, new_n10660_, new_n10661_,
    new_n10662_, new_n10663_, new_n10664_, new_n10665_, new_n10666_,
    new_n10667_, new_n10668_, new_n10669_, new_n10670_, new_n10671_,
    new_n10672_, new_n10673_, new_n10674_, new_n10675_, new_n10676_,
    new_n10677_, new_n10678_, new_n10679_, new_n10680_, new_n10681_,
    new_n10682_, new_n10683_, new_n10684_, new_n10685_, new_n10686_,
    new_n10687_, new_n10688_, new_n10689_, new_n10690_, new_n10691_,
    new_n10692_, new_n10693_, new_n10694_, new_n10695_, new_n10696_,
    new_n10697_, new_n10698_, new_n10699_, new_n10700_, new_n10701_,
    new_n10702_, new_n10703_, new_n10704_, new_n10705_, new_n10706_,
    new_n10707_, new_n10708_, new_n10709_, new_n10710_, new_n10711_,
    new_n10712_, new_n10713_, new_n10714_, new_n10715_, new_n10716_,
    new_n10717_, new_n10718_, new_n10719_, new_n10720_, new_n10721_,
    new_n10722_, new_n10723_, new_n10724_, new_n10725_, new_n10726_,
    new_n10727_, new_n10728_, new_n10729_, new_n10730_, new_n10731_,
    new_n10732_, new_n10733_, new_n10734_, new_n10735_, new_n10736_,
    new_n10737_, new_n10738_, new_n10739_, new_n10740_, new_n10741_,
    new_n10742_, new_n10743_, new_n10744_, new_n10745_, new_n10746_,
    new_n10747_, new_n10748_, new_n10749_, new_n10750_, new_n10751_,
    new_n10752_, new_n10753_, new_n10754_, new_n10755_, new_n10756_,
    new_n10757_, new_n10758_, new_n10759_, new_n10760_, new_n10761_,
    new_n10762_, new_n10763_, new_n10764_, new_n10765_, new_n10766_,
    new_n10767_, new_n10768_, new_n10769_, new_n10770_, new_n10771_,
    new_n10772_, new_n10773_, new_n10774_, new_n10775_, new_n10776_,
    new_n10777_, new_n10778_, new_n10779_, new_n10780_, new_n10781_,
    new_n10782_, new_n10783_, new_n10784_, new_n10785_, new_n10786_,
    new_n10787_, new_n10788_, new_n10789_, new_n10790_, new_n10791_,
    new_n10792_, new_n10793_, new_n10794_, new_n10795_, new_n10796_,
    new_n10797_, new_n10798_, new_n10799_, new_n10800_, new_n10801_,
    new_n10802_, new_n10803_, new_n10804_, new_n10805_, new_n10806_,
    new_n10807_, new_n10808_, new_n10809_, new_n10810_, new_n10811_,
    new_n10812_, new_n10813_, new_n10814_, new_n10815_, new_n10816_,
    new_n10817_, new_n10818_, new_n10819_, new_n10820_, new_n10821_,
    new_n10822_, new_n10823_, new_n10824_, new_n10825_, new_n10826_,
    new_n10827_, new_n10828_, new_n10829_, new_n10830_, new_n10831_,
    new_n10832_, new_n10833_, new_n10834_, new_n10835_, new_n10836_,
    new_n10837_, new_n10838_, new_n10839_, new_n10840_, new_n10841_,
    new_n10842_, new_n10843_, new_n10844_, new_n10845_, new_n10846_,
    new_n10847_, new_n10848_, new_n10849_, new_n10850_, new_n10851_,
    new_n10852_, new_n10853_, new_n10854_, new_n10855_, new_n10856_,
    new_n10857_, new_n10858_, new_n10859_, new_n10860_, new_n10861_,
    new_n10862_, new_n10863_, new_n10864_, new_n10865_, new_n10866_,
    new_n10867_, new_n10868_, new_n10869_, new_n10870_, new_n10871_,
    new_n10872_, new_n10873_, new_n10874_, new_n10875_, new_n10876_,
    new_n10877_, new_n10878_, new_n10879_, new_n10880_, new_n10881_,
    new_n10882_, new_n10883_, new_n10884_, new_n10885_, new_n10886_,
    new_n10887_, new_n10888_, new_n10889_, new_n10890_, new_n10891_,
    new_n10892_, new_n10893_, new_n10894_, new_n10895_, new_n10896_,
    new_n10897_, new_n10898_, new_n10899_, new_n10900_, new_n10901_,
    new_n10902_, new_n10903_, new_n10904_, new_n10905_, new_n10906_,
    new_n10907_, new_n10908_, new_n10909_, new_n10910_, new_n10911_,
    new_n10912_, new_n10913_, new_n10914_, new_n10915_, new_n10916_,
    new_n10917_, new_n10918_, new_n10919_, new_n10920_, new_n10921_,
    new_n10922_, new_n10923_, new_n10924_, new_n10925_, new_n10926_,
    new_n10927_, new_n10928_, new_n10929_, new_n10930_, new_n10931_,
    new_n10932_, new_n10933_, new_n10934_, new_n10935_, new_n10936_,
    new_n10937_, new_n10938_, new_n10939_, new_n10940_, new_n10941_,
    new_n10942_, new_n10943_, new_n10944_, new_n10945_, new_n10946_,
    new_n10947_, new_n10948_, new_n10949_, new_n10950_, new_n10951_,
    new_n10952_, new_n10953_, new_n10954_, new_n10955_, new_n10956_,
    new_n10957_, new_n10958_, new_n10959_, new_n10960_, new_n10961_,
    new_n10962_, new_n10963_, new_n10964_, new_n10965_, new_n10966_,
    new_n10967_, new_n10968_, new_n10969_, new_n10970_, new_n10971_,
    new_n10972_, new_n10973_, new_n10974_, new_n10975_, new_n10976_,
    new_n10977_, new_n10978_, new_n10979_, new_n10980_, new_n10981_,
    new_n10982_, new_n10983_, new_n10984_, new_n10985_, new_n10986_,
    new_n10987_, new_n10988_, new_n10989_, new_n10990_, new_n10991_,
    new_n10992_, new_n10993_, new_n10994_, new_n10995_, new_n10996_,
    new_n10997_, new_n10998_, new_n10999_, new_n11000_, new_n11001_,
    new_n11002_, new_n11003_, new_n11004_, new_n11005_, new_n11006_,
    new_n11007_, new_n11008_, new_n11009_, new_n11010_, new_n11011_,
    new_n11012_, new_n11013_, new_n11014_, new_n11015_, new_n11016_,
    new_n11017_, new_n11018_, new_n11019_, new_n11020_, new_n11021_,
    new_n11022_, new_n11023_, new_n11024_, new_n11025_, new_n11026_,
    new_n11027_, new_n11028_, new_n11029_, new_n11030_, new_n11031_,
    new_n11032_, new_n11033_, new_n11034_, new_n11035_, new_n11036_,
    new_n11037_, new_n11038_, new_n11039_, new_n11040_, new_n11041_,
    new_n11042_, new_n11043_, new_n11044_, new_n11045_, new_n11046_,
    new_n11047_, new_n11048_, new_n11049_, new_n11050_, new_n11051_,
    new_n11052_, new_n11053_, new_n11054_, new_n11055_, new_n11056_,
    new_n11057_, new_n11058_, new_n11059_, new_n11060_, new_n11061_,
    new_n11062_, new_n11064_, new_n11065_, new_n11066_, new_n11067_,
    new_n11068_, new_n11069_, new_n11070_, new_n11071_, new_n11072_,
    new_n11073_, new_n11074_, new_n11075_, new_n11076_, new_n11077_,
    new_n11078_, new_n11079_, new_n11080_, new_n11081_, new_n11082_,
    new_n11083_, new_n11084_, new_n11085_, new_n11086_, new_n11087_,
    new_n11088_, new_n11089_, new_n11090_, new_n11091_, new_n11092_,
    new_n11093_, new_n11094_, new_n11095_, new_n11096_, new_n11097_,
    new_n11098_, new_n11099_, new_n11100_, new_n11101_, new_n11102_,
    new_n11103_, new_n11104_, new_n11105_, new_n11106_, new_n11107_,
    new_n11108_, new_n11109_, new_n11110_, new_n11111_, new_n11112_,
    new_n11113_, new_n11114_, new_n11115_, new_n11116_, new_n11117_,
    new_n11118_, new_n11119_, new_n11120_, new_n11121_, new_n11122_,
    new_n11123_, new_n11124_, new_n11125_, new_n11126_, new_n11127_,
    new_n11128_, new_n11129_, new_n11130_, new_n11131_, new_n11132_,
    new_n11133_, new_n11134_, new_n11135_, new_n11136_, new_n11137_,
    new_n11138_, new_n11139_, new_n11140_, new_n11141_, new_n11142_,
    new_n11143_, new_n11144_, new_n11145_, new_n11146_, new_n11147_,
    new_n11148_, new_n11149_, new_n11150_, new_n11151_, new_n11152_,
    new_n11153_, new_n11154_, new_n11155_, new_n11156_, new_n11157_,
    new_n11158_, new_n11159_, new_n11160_, new_n11161_, new_n11162_,
    new_n11163_, new_n11164_, new_n11165_, new_n11166_, new_n11167_,
    new_n11168_, new_n11169_, new_n11170_, new_n11171_, new_n11172_,
    new_n11173_, new_n11174_, new_n11175_, new_n11176_, new_n11177_,
    new_n11178_, new_n11179_, new_n11180_, new_n11181_, new_n11182_,
    new_n11183_, new_n11184_, new_n11185_, new_n11186_, new_n11187_,
    new_n11188_, new_n11189_, new_n11190_, new_n11191_, new_n11192_,
    new_n11193_, new_n11194_, new_n11195_, new_n11196_, new_n11197_,
    new_n11198_, new_n11199_, new_n11200_, new_n11201_, new_n11202_,
    new_n11203_, new_n11204_, new_n11205_, new_n11206_, new_n11207_,
    new_n11208_, new_n11209_, new_n11210_, new_n11211_, new_n11212_,
    new_n11213_, new_n11214_, new_n11215_, new_n11216_, new_n11217_,
    new_n11218_, new_n11219_, new_n11220_, new_n11221_, new_n11222_,
    new_n11223_, new_n11224_, new_n11225_, new_n11226_, new_n11227_,
    new_n11228_, new_n11229_, new_n11230_, new_n11231_, new_n11232_,
    new_n11233_, new_n11234_, new_n11235_, new_n11236_, new_n11237_,
    new_n11238_, new_n11239_, new_n11240_, new_n11241_, new_n11242_,
    new_n11243_, new_n11244_, new_n11245_, new_n11246_, new_n11247_,
    new_n11248_, new_n11249_, new_n11250_, new_n11251_, new_n11252_,
    new_n11253_, new_n11254_, new_n11255_, new_n11256_, new_n11257_,
    new_n11258_, new_n11259_, new_n11260_, new_n11261_, new_n11262_,
    new_n11263_, new_n11264_, new_n11265_, new_n11266_, new_n11267_,
    new_n11268_, new_n11269_, new_n11270_, new_n11271_, new_n11272_,
    new_n11273_, new_n11274_, new_n11275_, new_n11276_, new_n11277_,
    new_n11278_, new_n11279_, new_n11280_, new_n11281_, new_n11282_,
    new_n11283_, new_n11284_, new_n11285_, new_n11286_, new_n11287_,
    new_n11288_, new_n11289_, new_n11290_, new_n11291_, new_n11292_,
    new_n11293_, new_n11294_, new_n11295_, new_n11296_, new_n11297_,
    new_n11298_, new_n11299_, new_n11300_, new_n11301_, new_n11302_,
    new_n11303_, new_n11304_, new_n11305_, new_n11306_, new_n11307_,
    new_n11308_, new_n11309_, new_n11310_, new_n11311_, new_n11312_,
    new_n11313_, new_n11314_, new_n11315_, new_n11316_, new_n11317_,
    new_n11318_, new_n11319_, new_n11320_, new_n11321_, new_n11322_,
    new_n11323_, new_n11324_, new_n11325_, new_n11326_, new_n11327_,
    new_n11328_, new_n11329_, new_n11330_, new_n11331_, new_n11332_,
    new_n11333_, new_n11334_, new_n11335_, new_n11336_, new_n11337_,
    new_n11338_, new_n11339_, new_n11340_, new_n11341_, new_n11342_,
    new_n11343_, new_n11344_, new_n11345_, new_n11346_, new_n11347_,
    new_n11348_, new_n11349_, new_n11350_, new_n11351_, new_n11352_,
    new_n11353_, new_n11354_, new_n11355_, new_n11356_, new_n11357_,
    new_n11358_, new_n11359_, new_n11360_, new_n11361_, new_n11362_,
    new_n11363_, new_n11364_, new_n11365_, new_n11366_, new_n11367_,
    new_n11368_, new_n11369_, new_n11370_, new_n11371_, new_n11372_,
    new_n11373_, new_n11374_, new_n11375_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11383_, new_n11384_, new_n11385_, new_n11386_, new_n11387_,
    new_n11388_, new_n11389_, new_n11390_, new_n11391_, new_n11392_,
    new_n11393_, new_n11394_, new_n11395_, new_n11396_, new_n11397_,
    new_n11398_, new_n11399_, new_n11400_, new_n11401_, new_n11402_,
    new_n11403_, new_n11404_, new_n11405_, new_n11406_, new_n11407_,
    new_n11408_, new_n11409_, new_n11410_, new_n11411_, new_n11412_,
    new_n11413_, new_n11414_, new_n11415_, new_n11416_, new_n11417_,
    new_n11418_, new_n11419_, new_n11420_, new_n11421_, new_n11422_,
    new_n11423_, new_n11424_, new_n11425_, new_n11426_, new_n11427_,
    new_n11428_, new_n11429_, new_n11430_, new_n11431_, new_n11432_,
    new_n11433_, new_n11434_, new_n11435_, new_n11436_, new_n11437_,
    new_n11438_, new_n11439_, new_n11440_, new_n11441_, new_n11442_,
    new_n11443_, new_n11444_, new_n11445_, new_n11446_, new_n11447_,
    new_n11448_, new_n11449_, new_n11450_, new_n11451_, new_n11452_,
    new_n11453_, new_n11454_, new_n11455_, new_n11456_, new_n11457_,
    new_n11458_, new_n11459_, new_n11460_, new_n11461_, new_n11462_,
    new_n11463_, new_n11464_, new_n11465_, new_n11466_, new_n11467_,
    new_n11468_, new_n11469_, new_n11470_, new_n11471_, new_n11472_,
    new_n11473_, new_n11474_, new_n11475_, new_n11476_, new_n11477_,
    new_n11478_, new_n11479_, new_n11480_, new_n11481_, new_n11482_,
    new_n11483_, new_n11484_, new_n11485_, new_n11486_, new_n11487_,
    new_n11488_, new_n11489_, new_n11490_, new_n11491_, new_n11492_,
    new_n11493_, new_n11494_, new_n11495_, new_n11496_, new_n11497_,
    new_n11498_, new_n11499_, new_n11500_, new_n11501_, new_n11502_,
    new_n11503_, new_n11504_, new_n11505_, new_n11506_, new_n11507_,
    new_n11508_, new_n11509_, new_n11510_, new_n11511_, new_n11512_,
    new_n11513_, new_n11514_, new_n11515_, new_n11516_, new_n11517_,
    new_n11518_, new_n11519_, new_n11520_, new_n11521_, new_n11522_,
    new_n11523_, new_n11524_, new_n11525_, new_n11526_, new_n11527_,
    new_n11528_, new_n11529_, new_n11530_, new_n11531_, new_n11532_,
    new_n11533_, new_n11534_, new_n11535_, new_n11536_, new_n11537_,
    new_n11538_, new_n11539_, new_n11540_, new_n11541_, new_n11542_,
    new_n11543_, new_n11544_, new_n11545_, new_n11546_, new_n11547_,
    new_n11548_, new_n11549_, new_n11550_, new_n11551_, new_n11552_,
    new_n11553_, new_n11554_, new_n11555_, new_n11556_, new_n11557_,
    new_n11558_, new_n11559_, new_n11560_, new_n11561_, new_n11562_,
    new_n11563_, new_n11564_, new_n11565_, new_n11566_, new_n11567_,
    new_n11568_, new_n11569_, new_n11570_, new_n11571_, new_n11572_,
    new_n11573_, new_n11574_, new_n11575_, new_n11576_, new_n11577_,
    new_n11578_, new_n11579_, new_n11580_, new_n11581_, new_n11582_,
    new_n11583_, new_n11584_, new_n11585_, new_n11586_, new_n11587_,
    new_n11588_, new_n11589_, new_n11590_, new_n11591_, new_n11592_,
    new_n11593_, new_n11595_, new_n11596_, new_n11597_, new_n11598_,
    new_n11599_, new_n11600_, new_n11601_, new_n11602_, new_n11603_,
    new_n11604_, new_n11605_, new_n11606_, new_n11607_, new_n11608_,
    new_n11609_, new_n11610_, new_n11611_, new_n11612_, new_n11613_,
    new_n11614_, new_n11615_, new_n11616_, new_n11617_, new_n11618_,
    new_n11619_, new_n11620_, new_n11621_, new_n11622_, new_n11623_,
    new_n11624_, new_n11625_, new_n11626_, new_n11627_, new_n11628_,
    new_n11629_, new_n11630_, new_n11631_, new_n11632_, new_n11633_,
    new_n11634_, new_n11635_, new_n11636_, new_n11637_, new_n11638_,
    new_n11639_, new_n11640_, new_n11641_, new_n11642_, new_n11643_,
    new_n11644_, new_n11645_, new_n11646_, new_n11647_, new_n11648_,
    new_n11649_, new_n11650_, new_n11651_, new_n11652_, new_n11653_,
    new_n11654_, new_n11655_, new_n11656_, new_n11657_, new_n11658_,
    new_n11659_, new_n11660_, new_n11661_, new_n11662_, new_n11663_,
    new_n11664_, new_n11665_, new_n11666_, new_n11667_, new_n11668_,
    new_n11669_, new_n11670_, new_n11671_, new_n11672_, new_n11673_,
    new_n11674_, new_n11675_, new_n11676_, new_n11677_, new_n11678_,
    new_n11679_, new_n11680_, new_n11681_, new_n11682_, new_n11683_,
    new_n11684_, new_n11685_, new_n11686_, new_n11687_, new_n11688_,
    new_n11689_, new_n11690_, new_n11691_, new_n11692_, new_n11693_,
    new_n11694_, new_n11695_, new_n11696_, new_n11697_, new_n11698_,
    new_n11699_, new_n11700_, new_n11701_, new_n11702_, new_n11703_,
    new_n11704_, new_n11705_, new_n11706_, new_n11707_, new_n11708_,
    new_n11709_, new_n11710_, new_n11711_, new_n11712_, new_n11713_,
    new_n11714_, new_n11715_, new_n11716_, new_n11717_, new_n11718_,
    new_n11719_, new_n11720_, new_n11721_, new_n11722_, new_n11723_,
    new_n11724_, new_n11725_, new_n11726_, new_n11727_, new_n11728_,
    new_n11729_, new_n11730_, new_n11731_, new_n11732_, new_n11733_,
    new_n11734_, new_n11735_, new_n11736_, new_n11737_, new_n11738_,
    new_n11739_, new_n11740_, new_n11741_, new_n11742_, new_n11743_,
    new_n11744_, new_n11745_, new_n11746_, new_n11747_, new_n11748_,
    new_n11749_, new_n11750_, new_n11751_, new_n11752_, new_n11753_,
    new_n11754_, new_n11755_, new_n11756_, new_n11757_, new_n11758_,
    new_n11759_, new_n11760_, new_n11761_, new_n11762_, new_n11763_,
    new_n11764_, new_n11765_, new_n11766_, new_n11767_, new_n11768_,
    new_n11769_, new_n11770_, new_n11771_, new_n11772_, new_n11773_,
    new_n11774_, new_n11775_, new_n11776_, new_n11777_, new_n11778_,
    new_n11779_, new_n11780_, new_n11781_, new_n11782_, new_n11783_,
    new_n11784_, new_n11785_, new_n11786_, new_n11787_, new_n11788_,
    new_n11789_, new_n11790_, new_n11791_, new_n11792_, new_n11793_,
    new_n11794_, new_n11795_, new_n11796_, new_n11797_, new_n11798_,
    new_n11799_, new_n11800_, new_n11801_, new_n11802_, new_n11803_,
    new_n11804_, new_n11805_, new_n11806_, new_n11807_, new_n11808_,
    new_n11809_, new_n11810_, new_n11811_, new_n11812_, new_n11813_,
    new_n11814_, new_n11815_, new_n11816_, new_n11817_, new_n11818_,
    new_n11819_, new_n11820_, new_n11821_, new_n11822_, new_n11823_,
    new_n11824_, new_n11825_, new_n11826_, new_n11827_, new_n11828_,
    new_n11829_, new_n11830_, new_n11831_, new_n11832_, new_n11833_,
    new_n11834_, new_n11835_, new_n11836_, new_n11837_, new_n11838_,
    new_n11839_, new_n11840_, new_n11841_, new_n11842_, new_n11843_,
    new_n11844_, new_n11845_, new_n11846_, new_n11847_, new_n11848_,
    new_n11849_, new_n11850_, new_n11851_, new_n11852_, new_n11853_,
    new_n11854_, new_n11855_, new_n11856_, new_n11857_, new_n11858_,
    new_n11859_, new_n11860_, new_n11861_, new_n11862_, new_n11863_,
    new_n11864_, new_n11865_, new_n11866_, new_n11867_, new_n11868_,
    new_n11869_, new_n11870_, new_n11871_, new_n11872_, new_n11873_,
    new_n11874_, new_n11875_, new_n11876_, new_n11877_, new_n11878_,
    new_n11879_, new_n11880_, new_n11881_, new_n11882_, new_n11883_,
    new_n11884_, new_n11885_, new_n11886_, new_n11887_, new_n11888_,
    new_n11889_, new_n11890_, new_n11891_, new_n11892_, new_n11893_,
    new_n11894_, new_n11895_, new_n11896_, new_n11897_, new_n11898_,
    new_n11899_, new_n11900_, new_n11901_, new_n11902_, new_n11903_,
    new_n11904_, new_n11905_, new_n11906_, new_n11907_, new_n11908_,
    new_n11909_, new_n11910_, new_n11911_, new_n11912_, new_n11913_,
    new_n11914_, new_n11915_, new_n11916_, new_n11917_, new_n11918_,
    new_n11919_, new_n11920_, new_n11921_, new_n11922_, new_n11923_,
    new_n11924_, new_n11925_, new_n11926_, new_n11927_, new_n11928_,
    new_n11929_, new_n11930_, new_n11931_, new_n11932_, new_n11933_,
    new_n11934_, new_n11935_, new_n11936_, new_n11937_, new_n11938_,
    new_n11939_, new_n11940_, new_n11941_, new_n11942_, new_n11943_,
    new_n11944_, new_n11945_, new_n11946_, new_n11947_, new_n11948_,
    new_n11949_, new_n11950_, new_n11951_, new_n11952_, new_n11953_,
    new_n11954_, new_n11955_, new_n11956_, new_n11957_, new_n11958_,
    new_n11959_, new_n11960_, new_n11961_, new_n11962_, new_n11963_,
    new_n11964_, new_n11965_, new_n11966_, new_n11967_, new_n11968_,
    new_n11969_, new_n11970_, new_n11971_, new_n11972_, new_n11973_,
    new_n11974_, new_n11975_, new_n11976_, new_n11977_, new_n11978_,
    new_n11979_, new_n11980_, new_n11981_, new_n11982_, new_n11983_,
    new_n11984_, new_n11985_, new_n11986_, new_n11987_, new_n11988_,
    new_n11989_, new_n11990_, new_n11991_, new_n11992_, new_n11993_,
    new_n11994_, new_n11995_, new_n11996_, new_n11997_, new_n11998_,
    new_n11999_, new_n12000_, new_n12001_, new_n12002_, new_n12003_,
    new_n12004_, new_n12005_, new_n12006_, new_n12007_, new_n12008_,
    new_n12009_, new_n12010_, new_n12011_, new_n12012_, new_n12013_,
    new_n12014_, new_n12015_, new_n12016_, new_n12017_, new_n12018_,
    new_n12019_, new_n12020_, new_n12021_, new_n12022_, new_n12023_,
    new_n12024_, new_n12025_, new_n12026_, new_n12027_, new_n12028_,
    new_n12029_, new_n12030_, new_n12031_, new_n12032_, new_n12033_,
    new_n12034_, new_n12035_, new_n12036_, new_n12037_, new_n12038_,
    new_n12039_, new_n12040_, new_n12041_, new_n12042_, new_n12043_,
    new_n12044_, new_n12045_, new_n12046_, new_n12047_, new_n12048_,
    new_n12049_, new_n12050_, new_n12051_, new_n12052_, new_n12053_,
    new_n12054_, new_n12055_, new_n12056_, new_n12057_, new_n12058_,
    new_n12059_, new_n12060_, new_n12061_, new_n12062_, new_n12063_,
    new_n12064_, new_n12065_, new_n12066_, new_n12067_, new_n12068_,
    new_n12069_, new_n12070_, new_n12071_, new_n12072_, new_n12073_,
    new_n12074_, new_n12075_, new_n12076_, new_n12077_, new_n12078_,
    new_n12079_, new_n12080_, new_n12081_, new_n12082_, new_n12083_,
    new_n12084_, new_n12085_, new_n12086_, new_n12087_, new_n12088_,
    new_n12089_, new_n12090_, new_n12091_, new_n12092_, new_n12093_,
    new_n12094_, new_n12095_, new_n12096_, new_n12097_, new_n12098_,
    new_n12099_, new_n12100_, new_n12101_, new_n12102_, new_n12103_,
    new_n12104_, new_n12105_, new_n12106_, new_n12107_, new_n12108_,
    new_n12109_, new_n12110_, new_n12111_, new_n12112_, new_n12113_,
    new_n12114_, new_n12115_, new_n12117_, new_n12118_, new_n12119_,
    new_n12120_, new_n12121_, new_n12122_, new_n12123_, new_n12124_,
    new_n12125_, new_n12126_, new_n12127_, new_n12128_, new_n12129_,
    new_n12130_, new_n12131_, new_n12132_, new_n12133_, new_n12134_,
    new_n12135_, new_n12136_, new_n12137_, new_n12138_, new_n12139_,
    new_n12140_, new_n12141_, new_n12142_, new_n12143_, new_n12144_,
    new_n12145_, new_n12146_, new_n12147_, new_n12148_, new_n12149_,
    new_n12150_, new_n12151_, new_n12152_, new_n12153_, new_n12154_,
    new_n12155_, new_n12156_, new_n12157_, new_n12158_, new_n12159_,
    new_n12160_, new_n12161_, new_n12162_, new_n12163_, new_n12164_,
    new_n12165_, new_n12166_, new_n12167_, new_n12168_, new_n12169_,
    new_n12170_, new_n12171_, new_n12172_, new_n12173_, new_n12174_,
    new_n12175_, new_n12176_, new_n12177_, new_n12178_, new_n12179_,
    new_n12180_, new_n12181_, new_n12182_, new_n12183_, new_n12184_,
    new_n12185_, new_n12186_, new_n12187_, new_n12188_, new_n12189_,
    new_n12190_, new_n12191_, new_n12192_, new_n12193_, new_n12194_,
    new_n12195_, new_n12196_, new_n12197_, new_n12198_, new_n12199_,
    new_n12200_, new_n12201_, new_n12202_, new_n12203_, new_n12204_,
    new_n12205_, new_n12206_, new_n12207_, new_n12208_, new_n12209_,
    new_n12210_, new_n12211_, new_n12212_, new_n12213_, new_n12214_,
    new_n12215_, new_n12216_, new_n12217_, new_n12218_, new_n12219_,
    new_n12220_, new_n12221_, new_n12222_, new_n12223_, new_n12224_,
    new_n12225_, new_n12226_, new_n12227_, new_n12228_, new_n12229_,
    new_n12230_, new_n12231_, new_n12232_, new_n12233_, new_n12234_,
    new_n12235_, new_n12236_, new_n12237_, new_n12238_, new_n12239_,
    new_n12240_, new_n12241_, new_n12242_, new_n12243_, new_n12244_,
    new_n12245_, new_n12246_, new_n12247_, new_n12248_, new_n12249_,
    new_n12250_, new_n12251_, new_n12252_, new_n12253_, new_n12254_,
    new_n12255_, new_n12256_, new_n12257_, new_n12258_, new_n12259_,
    new_n12260_, new_n12261_, new_n12262_, new_n12263_, new_n12264_,
    new_n12265_, new_n12266_, new_n12267_, new_n12268_, new_n12269_,
    new_n12270_, new_n12271_, new_n12272_, new_n12273_, new_n12274_,
    new_n12275_, new_n12276_, new_n12277_, new_n12278_, new_n12279_,
    new_n12280_, new_n12281_, new_n12282_, new_n12283_, new_n12284_,
    new_n12285_, new_n12286_, new_n12287_, new_n12288_, new_n12289_,
    new_n12290_, new_n12291_, new_n12292_, new_n12293_, new_n12294_,
    new_n12295_, new_n12296_, new_n12297_, new_n12298_, new_n12299_,
    new_n12300_, new_n12301_, new_n12302_, new_n12303_, new_n12304_,
    new_n12305_, new_n12306_, new_n12307_, new_n12308_, new_n12309_,
    new_n12310_, new_n12311_, new_n12312_, new_n12313_, new_n12314_,
    new_n12315_, new_n12316_, new_n12317_, new_n12318_, new_n12319_,
    new_n12320_, new_n12321_, new_n12322_, new_n12323_, new_n12324_,
    new_n12325_, new_n12326_, new_n12327_, new_n12328_, new_n12329_,
    new_n12330_, new_n12331_, new_n12332_, new_n12333_, new_n12334_,
    new_n12335_, new_n12336_, new_n12337_, new_n12338_, new_n12339_,
    new_n12340_, new_n12341_, new_n12342_, new_n12343_, new_n12344_,
    new_n12345_, new_n12346_, new_n12347_, new_n12348_, new_n12349_,
    new_n12350_, new_n12351_, new_n12352_, new_n12353_, new_n12354_,
    new_n12355_, new_n12356_, new_n12357_, new_n12358_, new_n12359_,
    new_n12360_, new_n12361_, new_n12362_, new_n12363_, new_n12364_,
    new_n12365_, new_n12366_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12375_, new_n12376_, new_n12377_, new_n12378_, new_n12379_,
    new_n12380_, new_n12381_, new_n12382_, new_n12383_, new_n12384_,
    new_n12385_, new_n12386_, new_n12387_, new_n12388_, new_n12389_,
    new_n12390_, new_n12391_, new_n12392_, new_n12393_, new_n12394_,
    new_n12395_, new_n12396_, new_n12397_, new_n12398_, new_n12399_,
    new_n12400_, new_n12401_, new_n12402_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12409_,
    new_n12410_, new_n12411_, new_n12412_, new_n12413_, new_n12414_,
    new_n12415_, new_n12416_, new_n12417_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12437_, new_n12438_, new_n12439_,
    new_n12440_, new_n12441_, new_n12442_, new_n12443_, new_n12444_,
    new_n12445_, new_n12446_, new_n12447_, new_n12448_, new_n12449_,
    new_n12450_, new_n12451_, new_n12452_, new_n12453_, new_n12454_,
    new_n12455_, new_n12456_, new_n12457_, new_n12458_, new_n12459_,
    new_n12460_, new_n12461_, new_n12462_, new_n12463_, new_n12464_,
    new_n12465_, new_n12466_, new_n12467_, new_n12468_, new_n12469_,
    new_n12470_, new_n12471_, new_n12472_, new_n12473_, new_n12474_,
    new_n12475_, new_n12476_, new_n12477_, new_n12478_, new_n12479_,
    new_n12480_, new_n12481_, new_n12482_, new_n12483_, new_n12484_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12489_,
    new_n12490_, new_n12491_, new_n12492_, new_n12493_, new_n12494_,
    new_n12495_, new_n12496_, new_n12497_, new_n12498_, new_n12499_,
    new_n12500_, new_n12501_, new_n12502_, new_n12503_, new_n12504_,
    new_n12505_, new_n12506_, new_n12507_, new_n12508_, new_n12509_,
    new_n12510_, new_n12511_, new_n12512_, new_n12513_, new_n12514_,
    new_n12515_, new_n12516_, new_n12517_, new_n12518_, new_n12519_,
    new_n12520_, new_n12521_, new_n12522_, new_n12523_, new_n12524_,
    new_n12525_, new_n12526_, new_n12527_, new_n12528_, new_n12529_,
    new_n12530_, new_n12531_, new_n12532_, new_n12533_, new_n12534_,
    new_n12535_, new_n12536_, new_n12537_, new_n12538_, new_n12539_,
    new_n12540_, new_n12541_, new_n12542_, new_n12543_, new_n12544_,
    new_n12545_, new_n12546_, new_n12547_, new_n12548_, new_n12549_,
    new_n12550_, new_n12551_, new_n12552_, new_n12553_, new_n12554_,
    new_n12555_, new_n12556_, new_n12557_, new_n12558_, new_n12559_,
    new_n12560_, new_n12561_, new_n12562_, new_n12563_, new_n12564_,
    new_n12565_, new_n12566_, new_n12567_, new_n12568_, new_n12569_,
    new_n12570_, new_n12571_, new_n12572_, new_n12573_, new_n12574_,
    new_n12575_, new_n12576_, new_n12577_, new_n12578_, new_n12579_,
    new_n12580_, new_n12581_, new_n12582_, new_n12583_, new_n12584_,
    new_n12585_, new_n12586_, new_n12587_, new_n12588_, new_n12589_,
    new_n12590_, new_n12591_, new_n12592_, new_n12593_, new_n12594_,
    new_n12595_, new_n12596_, new_n12597_, new_n12598_, new_n12599_,
    new_n12600_, new_n12601_, new_n12602_, new_n12603_, new_n12604_,
    new_n12605_, new_n12606_, new_n12607_, new_n12608_, new_n12609_,
    new_n12610_, new_n12611_, new_n12612_, new_n12613_, new_n12614_,
    new_n12615_, new_n12616_, new_n12617_, new_n12618_, new_n12619_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12656_, new_n12657_, new_n12658_, new_n12659_, new_n12660_,
    new_n12661_, new_n12662_, new_n12663_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12714_, new_n12715_,
    new_n12716_, new_n12717_, new_n12718_, new_n12719_, new_n12720_,
    new_n12721_, new_n12722_, new_n12723_, new_n12724_, new_n12725_,
    new_n12726_, new_n12727_, new_n12728_, new_n12729_, new_n12730_,
    new_n12731_, new_n12732_, new_n12733_, new_n12734_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12849_, new_n12850_,
    new_n12851_, new_n12852_, new_n12853_, new_n12854_, new_n12855_,
    new_n12856_, new_n12857_, new_n12858_, new_n12859_, new_n12860_,
    new_n12861_, new_n12862_, new_n12863_, new_n12864_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12909_, new_n12910_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12917_, new_n12918_, new_n12919_, new_n12920_,
    new_n12921_, new_n12922_, new_n12923_, new_n12924_, new_n12925_,
    new_n12926_, new_n12927_, new_n12928_, new_n12929_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12960_,
    new_n12961_, new_n12962_, new_n12963_, new_n12964_, new_n12965_,
    new_n12966_, new_n12967_, new_n12968_, new_n12969_, new_n12970_,
    new_n12971_, new_n12972_, new_n12973_, new_n12974_, new_n12975_,
    new_n12976_, new_n12977_, new_n12978_, new_n12979_, new_n12980_,
    new_n12981_, new_n12982_, new_n12983_, new_n12984_, new_n12985_,
    new_n12986_, new_n12987_, new_n12988_, new_n12989_, new_n12990_,
    new_n12991_, new_n12992_, new_n12993_, new_n12994_, new_n12995_,
    new_n12996_, new_n12997_, new_n12998_, new_n12999_, new_n13000_,
    new_n13001_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13151_,
    new_n13152_, new_n13153_, new_n13154_, new_n13155_, new_n13156_,
    new_n13157_, new_n13158_, new_n13159_, new_n13160_, new_n13161_,
    new_n13162_, new_n13163_, new_n13164_, new_n13165_, new_n13166_,
    new_n13167_, new_n13168_, new_n13169_, new_n13170_, new_n13171_,
    new_n13172_, new_n13173_, new_n13174_, new_n13175_, new_n13176_,
    new_n13177_, new_n13178_, new_n13179_, new_n13180_, new_n13181_,
    new_n13182_, new_n13183_, new_n13184_, new_n13185_, new_n13186_,
    new_n13187_, new_n13188_, new_n13189_, new_n13190_, new_n13191_,
    new_n13192_, new_n13193_, new_n13194_, new_n13195_, new_n13196_,
    new_n13197_, new_n13198_, new_n13199_, new_n13200_, new_n13201_,
    new_n13202_, new_n13203_, new_n13204_, new_n13205_, new_n13206_,
    new_n13207_, new_n13208_, new_n13209_, new_n13210_, new_n13211_,
    new_n13212_, new_n13213_, new_n13214_, new_n13215_, new_n13216_,
    new_n13217_, new_n13218_, new_n13219_, new_n13220_, new_n13221_,
    new_n13222_, new_n13223_, new_n13224_, new_n13225_, new_n13226_,
    new_n13227_, new_n13228_, new_n13229_, new_n13230_, new_n13231_,
    new_n13232_, new_n13233_, new_n13234_, new_n13235_, new_n13236_,
    new_n13237_, new_n13238_, new_n13239_, new_n13240_, new_n13241_,
    new_n13242_, new_n13243_, new_n13244_, new_n13245_, new_n13246_,
    new_n13247_, new_n13248_, new_n13249_, new_n13250_, new_n13251_,
    new_n13252_, new_n13253_, new_n13254_, new_n13255_, new_n13256_,
    new_n13257_, new_n13258_, new_n13259_, new_n13260_, new_n13261_,
    new_n13262_, new_n13263_, new_n13264_, new_n13265_, new_n13266_,
    new_n13267_, new_n13268_, new_n13269_, new_n13270_, new_n13271_,
    new_n13272_, new_n13273_, new_n13274_, new_n13275_, new_n13276_,
    new_n13277_, new_n13278_, new_n13279_, new_n13280_, new_n13281_,
    new_n13282_, new_n13283_, new_n13284_, new_n13285_, new_n13286_,
    new_n13287_, new_n13288_, new_n13289_, new_n13290_, new_n13291_,
    new_n13292_, new_n13293_, new_n13294_, new_n13295_, new_n13296_,
    new_n13297_, new_n13298_, new_n13299_, new_n13300_, new_n13301_,
    new_n13302_, new_n13303_, new_n13304_, new_n13305_, new_n13306_,
    new_n13307_, new_n13308_, new_n13309_, new_n13310_, new_n13311_,
    new_n13312_, new_n13313_, new_n13314_, new_n13315_, new_n13316_,
    new_n13317_, new_n13318_, new_n13319_, new_n13320_, new_n13321_,
    new_n13322_, new_n13323_, new_n13324_, new_n13325_, new_n13326_,
    new_n13327_, new_n13328_, new_n13329_, new_n13330_, new_n13331_,
    new_n13332_, new_n13333_, new_n13334_, new_n13335_, new_n13336_,
    new_n13337_, new_n13338_, new_n13339_, new_n13340_, new_n13341_,
    new_n13342_, new_n13343_, new_n13344_, new_n13345_, new_n13346_,
    new_n13347_, new_n13348_, new_n13349_, new_n13350_, new_n13351_,
    new_n13352_, new_n13353_, new_n13354_, new_n13355_, new_n13356_,
    new_n13357_, new_n13358_, new_n13359_, new_n13360_, new_n13361_,
    new_n13362_, new_n13363_, new_n13364_, new_n13365_, new_n13366_,
    new_n13367_, new_n13368_, new_n13369_, new_n13370_, new_n13371_,
    new_n13372_, new_n13373_, new_n13374_, new_n13375_, new_n13376_,
    new_n13377_, new_n13378_, new_n13379_, new_n13380_, new_n13381_,
    new_n13382_, new_n13383_, new_n13384_, new_n13385_, new_n13386_,
    new_n13387_, new_n13388_, new_n13389_, new_n13390_, new_n13391_,
    new_n13392_, new_n13393_, new_n13394_, new_n13395_, new_n13396_,
    new_n13397_, new_n13398_, new_n13399_, new_n13400_, new_n13401_,
    new_n13402_, new_n13403_, new_n13404_, new_n13405_, new_n13406_,
    new_n13407_, new_n13408_, new_n13409_, new_n13410_, new_n13411_,
    new_n13412_, new_n13413_, new_n13414_, new_n13415_, new_n13416_,
    new_n13417_, new_n13418_, new_n13419_, new_n13420_, new_n13421_,
    new_n13422_, new_n13423_, new_n13424_, new_n13425_, new_n13426_,
    new_n13427_, new_n13428_, new_n13429_, new_n13430_, new_n13431_,
    new_n13432_, new_n13433_, new_n13434_, new_n13435_, new_n13436_,
    new_n13437_, new_n13438_, new_n13439_, new_n13440_, new_n13441_,
    new_n13442_, new_n13443_, new_n13444_, new_n13445_, new_n13446_,
    new_n13447_, new_n13448_, new_n13449_, new_n13450_, new_n13451_,
    new_n13452_, new_n13453_, new_n13454_, new_n13455_, new_n13456_,
    new_n13457_, new_n13458_, new_n13459_, new_n13460_, new_n13461_,
    new_n13462_, new_n13463_, new_n13464_, new_n13465_, new_n13466_,
    new_n13467_, new_n13468_, new_n13469_, new_n13470_, new_n13471_,
    new_n13472_, new_n13473_, new_n13474_, new_n13475_, new_n13476_,
    new_n13477_, new_n13478_, new_n13479_, new_n13480_, new_n13481_,
    new_n13482_, new_n13483_, new_n13484_, new_n13485_, new_n13486_,
    new_n13487_, new_n13488_, new_n13489_, new_n13490_, new_n13491_,
    new_n13492_, new_n13493_, new_n13494_, new_n13495_, new_n13496_,
    new_n13497_, new_n13498_, new_n13499_, new_n13500_, new_n13501_,
    new_n13502_, new_n13503_, new_n13504_, new_n13505_, new_n13506_,
    new_n13507_, new_n13508_, new_n13509_, new_n13510_, new_n13511_,
    new_n13512_, new_n13513_, new_n13514_, new_n13515_, new_n13516_,
    new_n13517_, new_n13518_, new_n13519_, new_n13520_, new_n13521_,
    new_n13522_, new_n13523_, new_n13524_, new_n13525_, new_n13526_,
    new_n13527_, new_n13528_, new_n13529_, new_n13530_, new_n13531_,
    new_n13532_, new_n13533_, new_n13534_, new_n13535_, new_n13536_,
    new_n13537_, new_n13538_, new_n13539_, new_n13540_, new_n13541_,
    new_n13542_, new_n13543_, new_n13544_, new_n13545_, new_n13546_,
    new_n13547_, new_n13548_, new_n13549_, new_n13550_, new_n13551_,
    new_n13552_, new_n13553_, new_n13554_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13596_,
    new_n13597_, new_n13598_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13605_, new_n13606_,
    new_n13607_, new_n13608_, new_n13609_, new_n13610_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13637_, new_n13638_, new_n13639_, new_n13640_, new_n13641_,
    new_n13642_, new_n13643_, new_n13644_, new_n13645_, new_n13646_,
    new_n13647_, new_n13648_, new_n13649_, new_n13650_, new_n13651_,
    new_n13652_, new_n13653_, new_n13654_, new_n13655_, new_n13656_,
    new_n13657_, new_n13658_, new_n13659_, new_n13660_, new_n13661_,
    new_n13662_, new_n13663_, new_n13664_, new_n13665_, new_n13666_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13724_, new_n13725_, new_n13726_, new_n13727_,
    new_n13728_, new_n13729_, new_n13730_, new_n13731_, new_n13732_,
    new_n13733_, new_n13734_, new_n13735_, new_n13736_, new_n13737_,
    new_n13738_, new_n13739_, new_n13740_, new_n13741_, new_n13742_,
    new_n13743_, new_n13744_, new_n13745_, new_n13746_, new_n13747_,
    new_n13748_, new_n13749_, new_n13750_, new_n13751_, new_n13752_,
    new_n13753_, new_n13754_, new_n13755_, new_n13756_, new_n13757_,
    new_n13758_, new_n13759_, new_n13760_, new_n13761_, new_n13762_,
    new_n13763_, new_n13764_, new_n13765_, new_n13766_, new_n13767_,
    new_n13768_, new_n13769_, new_n13770_, new_n13771_, new_n13772_,
    new_n13773_, new_n13774_, new_n13775_, new_n13776_, new_n13777_,
    new_n13778_, new_n13779_, new_n13780_, new_n13781_, new_n13782_,
    new_n13783_, new_n13784_, new_n13785_, new_n13786_, new_n13787_,
    new_n13788_, new_n13789_, new_n13790_, new_n13791_, new_n13792_,
    new_n13793_, new_n13794_, new_n13795_, new_n13796_, new_n13797_,
    new_n13798_, new_n13799_, new_n13800_, new_n13801_, new_n13802_,
    new_n13803_, new_n13804_, new_n13805_, new_n13806_, new_n13807_,
    new_n13808_, new_n13809_, new_n13810_, new_n13811_, new_n13812_,
    new_n13813_, new_n13814_, new_n13815_, new_n13816_, new_n13817_,
    new_n13818_, new_n13819_, new_n13820_, new_n13821_, new_n13822_,
    new_n13823_, new_n13824_, new_n13825_, new_n13826_, new_n13827_,
    new_n13828_, new_n13829_, new_n13830_, new_n13831_, new_n13832_,
    new_n13833_, new_n13834_, new_n13835_, new_n13836_, new_n13837_,
    new_n13838_, new_n13839_, new_n13840_, new_n13841_, new_n13842_,
    new_n13843_, new_n13844_, new_n13845_, new_n13846_, new_n13847_,
    new_n13848_, new_n13849_, new_n13850_, new_n13851_, new_n13852_,
    new_n13853_, new_n13854_, new_n13855_, new_n13856_, new_n13857_,
    new_n13858_, new_n13859_, new_n13860_, new_n13861_, new_n13862_,
    new_n13863_, new_n13864_, new_n13865_, new_n13866_, new_n13867_,
    new_n13868_, new_n13869_, new_n13870_, new_n13871_, new_n13872_,
    new_n13873_, new_n13874_, new_n13875_, new_n13876_, new_n13877_,
    new_n13878_, new_n13879_, new_n13880_, new_n13881_, new_n13882_,
    new_n13883_, new_n13884_, new_n13885_, new_n13886_, new_n13887_,
    new_n13888_, new_n13889_, new_n13890_, new_n13891_, new_n13892_,
    new_n13893_, new_n13894_, new_n13895_, new_n13896_, new_n13897_,
    new_n13898_, new_n13899_, new_n13900_, new_n13901_, new_n13902_,
    new_n13903_, new_n13904_, new_n13905_, new_n13906_, new_n13907_,
    new_n13908_, new_n13909_, new_n13910_, new_n13911_, new_n13912_,
    new_n13913_, new_n13914_, new_n13915_, new_n13916_, new_n13917_,
    new_n13918_, new_n13919_, new_n13920_, new_n13921_, new_n13922_,
    new_n13923_, new_n13924_, new_n13925_, new_n13926_, new_n13927_,
    new_n13928_, new_n13929_, new_n13930_, new_n13931_, new_n13932_,
    new_n13933_, new_n13934_, new_n13935_, new_n13936_, new_n13937_,
    new_n13938_, new_n13939_, new_n13940_, new_n13941_, new_n13942_,
    new_n13943_, new_n13944_, new_n13945_, new_n13946_, new_n13947_,
    new_n13948_, new_n13949_, new_n13950_, new_n13951_, new_n13952_,
    new_n13953_, new_n13954_, new_n13955_, new_n13956_, new_n13957_,
    new_n13958_, new_n13959_, new_n13960_, new_n13961_, new_n13962_,
    new_n13963_, new_n13964_, new_n13965_, new_n13966_, new_n13967_,
    new_n13968_, new_n13969_, new_n13970_, new_n13971_, new_n13972_,
    new_n13973_, new_n13974_, new_n13975_, new_n13976_, new_n13977_,
    new_n13978_, new_n13979_, new_n13980_, new_n13981_, new_n13982_,
    new_n13983_, new_n13984_, new_n13985_, new_n13986_, new_n13987_,
    new_n13988_, new_n13989_, new_n13990_, new_n13991_, new_n13992_,
    new_n13993_, new_n13994_, new_n13995_, new_n13996_, new_n13997_,
    new_n13998_, new_n13999_, new_n14000_, new_n14001_, new_n14002_,
    new_n14003_, new_n14004_, new_n14005_, new_n14006_, new_n14007_,
    new_n14008_, new_n14009_, new_n14010_, new_n14011_, new_n14012_,
    new_n14013_, new_n14014_, new_n14015_, new_n14016_, new_n14017_,
    new_n14018_, new_n14019_, new_n14020_, new_n14021_, new_n14022_,
    new_n14023_, new_n14024_, new_n14025_, new_n14026_, new_n14027_,
    new_n14028_, new_n14029_, new_n14030_, new_n14031_, new_n14032_,
    new_n14033_, new_n14034_, new_n14035_, new_n14036_, new_n14037_,
    new_n14038_, new_n14039_, new_n14040_, new_n14041_, new_n14042_,
    new_n14043_, new_n14044_, new_n14045_, new_n14046_, new_n14047_,
    new_n14048_, new_n14049_, new_n14050_, new_n14051_, new_n14052_,
    new_n14053_, new_n14054_, new_n14055_, new_n14056_, new_n14057_,
    new_n14058_, new_n14059_, new_n14060_, new_n14061_, new_n14062_,
    new_n14063_, new_n14064_, new_n14065_, new_n14066_, new_n14067_,
    new_n14068_, new_n14069_, new_n14070_, new_n14071_, new_n14072_,
    new_n14073_, new_n14074_, new_n14075_, new_n14076_, new_n14077_,
    new_n14078_, new_n14079_, new_n14080_, new_n14081_, new_n14082_,
    new_n14083_, new_n14084_, new_n14085_, new_n14086_, new_n14087_,
    new_n14088_, new_n14089_, new_n14090_, new_n14091_, new_n14092_,
    new_n14093_, new_n14094_, new_n14095_, new_n14096_, new_n14097_,
    new_n14098_, new_n14099_, new_n14100_, new_n14101_, new_n14102_,
    new_n14103_, new_n14104_, new_n14105_, new_n14106_, new_n14107_,
    new_n14108_, new_n14109_, new_n14110_, new_n14111_, new_n14112_,
    new_n14113_, new_n14114_, new_n14115_, new_n14116_, new_n14117_,
    new_n14118_, new_n14119_, new_n14120_, new_n14121_, new_n14122_,
    new_n14123_, new_n14124_, new_n14125_, new_n14126_, new_n14127_,
    new_n14128_, new_n14129_, new_n14130_, new_n14131_, new_n14132_,
    new_n14133_, new_n14134_, new_n14135_, new_n14136_, new_n14137_,
    new_n14138_, new_n14139_, new_n14140_, new_n14141_, new_n14142_,
    new_n14143_, new_n14144_, new_n14145_, new_n14146_, new_n14147_,
    new_n14148_, new_n14149_, new_n14150_, new_n14151_, new_n14152_,
    new_n14153_, new_n14154_, new_n14155_, new_n14156_, new_n14157_,
    new_n14158_, new_n14159_, new_n14160_, new_n14161_, new_n14162_,
    new_n14163_, new_n14164_, new_n14165_, new_n14166_, new_n14167_,
    new_n14168_, new_n14169_, new_n14170_, new_n14171_, new_n14172_,
    new_n14173_, new_n14174_, new_n14175_, new_n14176_, new_n14177_,
    new_n14178_, new_n14179_, new_n14180_, new_n14181_, new_n14182_,
    new_n14183_, new_n14184_, new_n14185_, new_n14186_, new_n14187_,
    new_n14188_, new_n14189_, new_n14190_, new_n14191_, new_n14192_,
    new_n14193_, new_n14194_, new_n14195_, new_n14196_, new_n14197_,
    new_n14198_, new_n14199_, new_n14200_, new_n14201_, new_n14202_,
    new_n14203_, new_n14204_, new_n14205_, new_n14206_, new_n14207_,
    new_n14208_, new_n14209_, new_n14210_, new_n14211_, new_n14212_,
    new_n14213_, new_n14214_, new_n14215_, new_n14216_, new_n14217_,
    new_n14218_, new_n14219_, new_n14220_, new_n14221_, new_n14222_,
    new_n14223_, new_n14224_, new_n14225_, new_n14226_, new_n14227_,
    new_n14228_, new_n14229_, new_n14230_, new_n14231_, new_n14232_,
    new_n14233_, new_n14234_, new_n14235_, new_n14236_, new_n14237_,
    new_n14238_, new_n14239_, new_n14240_, new_n14241_, new_n14242_,
    new_n14243_, new_n14244_, new_n14245_, new_n14246_, new_n14247_,
    new_n14248_, new_n14249_, new_n14250_, new_n14251_, new_n14252_,
    new_n14253_, new_n14254_, new_n14255_, new_n14256_, new_n14257_,
    new_n14258_, new_n14259_, new_n14260_, new_n14261_, new_n14262_,
    new_n14263_, new_n14264_, new_n14265_, new_n14266_, new_n14267_,
    new_n14268_, new_n14269_, new_n14270_, new_n14271_, new_n14272_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14289_, new_n14290_, new_n14291_, new_n14292_, new_n14293_,
    new_n14294_, new_n14295_, new_n14296_, new_n14297_, new_n14298_,
    new_n14299_, new_n14300_, new_n14301_, new_n14302_, new_n14303_,
    new_n14304_, new_n14305_, new_n14306_, new_n14307_, new_n14308_,
    new_n14309_, new_n14310_, new_n14311_, new_n14312_, new_n14313_,
    new_n14314_, new_n14315_, new_n14316_, new_n14317_, new_n14318_,
    new_n14319_, new_n14320_, new_n14321_, new_n14322_, new_n14323_,
    new_n14324_, new_n14325_, new_n14326_, new_n14327_, new_n14328_,
    new_n14329_, new_n14330_, new_n14331_, new_n14332_, new_n14333_,
    new_n14334_, new_n14335_, new_n14336_, new_n14337_, new_n14338_,
    new_n14339_, new_n14340_, new_n14341_, new_n14342_, new_n14343_,
    new_n14344_, new_n14345_, new_n14346_, new_n14347_, new_n14348_,
    new_n14349_, new_n14350_, new_n14351_, new_n14352_, new_n14353_,
    new_n14354_, new_n14355_, new_n14356_, new_n14357_, new_n14358_,
    new_n14359_, new_n14360_, new_n14361_, new_n14362_, new_n14363_,
    new_n14364_, new_n14365_, new_n14366_, new_n14367_, new_n14368_,
    new_n14369_, new_n14370_, new_n14371_, new_n14372_, new_n14373_,
    new_n14374_, new_n14375_, new_n14376_, new_n14377_, new_n14378_,
    new_n14379_, new_n14380_, new_n14381_, new_n14382_, new_n14383_,
    new_n14384_, new_n14385_, new_n14386_, new_n14387_, new_n14388_,
    new_n14389_, new_n14390_, new_n14391_, new_n14392_, new_n14393_,
    new_n14394_, new_n14395_, new_n14396_, new_n14397_, new_n14398_,
    new_n14399_, new_n14400_, new_n14401_, new_n14402_, new_n14403_,
    new_n14404_, new_n14405_, new_n14406_, new_n14407_, new_n14408_,
    new_n14409_, new_n14410_, new_n14411_, new_n14412_, new_n14413_,
    new_n14414_, new_n14415_, new_n14416_, new_n14417_, new_n14418_,
    new_n14419_, new_n14420_, new_n14421_, new_n14422_, new_n14423_,
    new_n14424_, new_n14425_, new_n14426_, new_n14427_, new_n14428_,
    new_n14429_, new_n14430_, new_n14431_, new_n14432_, new_n14433_,
    new_n14434_, new_n14435_, new_n14436_, new_n14437_, new_n14438_,
    new_n14439_, new_n14440_, new_n14441_, new_n14442_, new_n14443_,
    new_n14444_, new_n14445_, new_n14446_, new_n14447_, new_n14448_,
    new_n14449_, new_n14450_, new_n14451_, new_n14452_, new_n14453_,
    new_n14454_, new_n14455_, new_n14456_, new_n14457_, new_n14458_,
    new_n14459_, new_n14460_, new_n14461_, new_n14462_, new_n14463_,
    new_n14464_, new_n14465_, new_n14466_, new_n14467_, new_n14468_,
    new_n14469_, new_n14470_, new_n14471_, new_n14472_, new_n14473_,
    new_n14474_, new_n14475_, new_n14476_, new_n14477_, new_n14478_,
    new_n14479_, new_n14480_, new_n14481_, new_n14482_, new_n14483_,
    new_n14484_, new_n14485_, new_n14486_, new_n14487_, new_n14488_,
    new_n14489_, new_n14490_, new_n14491_, new_n14492_, new_n14493_,
    new_n14494_, new_n14495_, new_n14496_, new_n14497_, new_n14498_,
    new_n14499_, new_n14500_, new_n14501_, new_n14502_, new_n14503_,
    new_n14504_, new_n14505_, new_n14506_, new_n14507_, new_n14508_,
    new_n14509_, new_n14510_, new_n14511_, new_n14512_, new_n14513_,
    new_n14514_, new_n14515_, new_n14516_, new_n14517_, new_n14518_,
    new_n14519_, new_n14520_, new_n14521_, new_n14522_, new_n14523_,
    new_n14524_, new_n14525_, new_n14526_, new_n14527_, new_n14528_,
    new_n14529_, new_n14530_, new_n14531_, new_n14532_, new_n14533_,
    new_n14534_, new_n14535_, new_n14536_, new_n14537_, new_n14538_,
    new_n14539_, new_n14540_, new_n14541_, new_n14542_, new_n14543_,
    new_n14544_, new_n14545_, new_n14546_, new_n14547_, new_n14548_,
    new_n14549_, new_n14550_, new_n14551_, new_n14552_, new_n14553_,
    new_n14554_, new_n14555_, new_n14556_, new_n14557_, new_n14558_,
    new_n14559_, new_n14560_, new_n14561_, new_n14562_, new_n14563_,
    new_n14564_, new_n14565_, new_n14566_, new_n14567_, new_n14568_,
    new_n14569_, new_n14570_, new_n14571_, new_n14572_, new_n14573_,
    new_n14574_, new_n14575_, new_n14576_, new_n14577_, new_n14578_,
    new_n14579_, new_n14580_, new_n14581_, new_n14582_, new_n14583_,
    new_n14584_, new_n14585_, new_n14586_, new_n14587_, new_n14588_,
    new_n14589_, new_n14590_, new_n14591_, new_n14592_, new_n14593_,
    new_n14594_, new_n14595_, new_n14596_, new_n14597_, new_n14598_,
    new_n14599_, new_n14600_, new_n14601_, new_n14602_, new_n14603_,
    new_n14604_, new_n14605_, new_n14606_, new_n14607_, new_n14608_,
    new_n14609_, new_n14610_, new_n14611_, new_n14612_, new_n14613_,
    new_n14614_, new_n14615_, new_n14616_, new_n14617_, new_n14618_,
    new_n14619_, new_n14620_, new_n14621_, new_n14622_, new_n14623_,
    new_n14624_, new_n14625_, new_n14626_, new_n14627_, new_n14628_,
    new_n14629_, new_n14630_, new_n14631_, new_n14632_, new_n14633_,
    new_n14634_, new_n14635_, new_n14636_, new_n14637_, new_n14638_,
    new_n14639_, new_n14640_, new_n14641_, new_n14642_, new_n14643_,
    new_n14644_, new_n14645_, new_n14646_, new_n14647_, new_n14648_,
    new_n14649_, new_n14650_, new_n14651_, new_n14652_, new_n14653_,
    new_n14654_, new_n14655_, new_n14656_, new_n14657_, new_n14658_,
    new_n14659_, new_n14660_, new_n14661_, new_n14662_, new_n14663_,
    new_n14664_, new_n14665_, new_n14666_, new_n14667_, new_n14668_,
    new_n14669_, new_n14670_, new_n14671_, new_n14672_, new_n14673_,
    new_n14674_, new_n14675_, new_n14676_, new_n14677_, new_n14678_,
    new_n14679_, new_n14680_, new_n14681_, new_n14682_, new_n14683_,
    new_n14684_, new_n14685_, new_n14686_, new_n14687_, new_n14688_,
    new_n14689_, new_n14690_, new_n14691_, new_n14692_, new_n14693_,
    new_n14694_, new_n14695_, new_n14696_, new_n14697_, new_n14698_,
    new_n14699_, new_n14700_, new_n14701_, new_n14702_, new_n14703_,
    new_n14704_, new_n14705_, new_n14706_, new_n14707_, new_n14708_,
    new_n14709_, new_n14710_, new_n14711_, new_n14712_, new_n14713_,
    new_n14714_, new_n14715_, new_n14716_, new_n14717_, new_n14718_,
    new_n14719_, new_n14720_, new_n14721_, new_n14722_, new_n14723_,
    new_n14724_, new_n14725_, new_n14726_, new_n14727_, new_n14728_,
    new_n14729_, new_n14730_, new_n14731_, new_n14732_, new_n14733_,
    new_n14734_, new_n14735_, new_n14736_, new_n14737_, new_n14738_,
    new_n14739_, new_n14740_, new_n14741_, new_n14742_, new_n14743_,
    new_n14744_, new_n14745_, new_n14746_, new_n14747_, new_n14748_,
    new_n14749_, new_n14750_, new_n14751_, new_n14752_, new_n14753_,
    new_n14754_, new_n14755_, new_n14756_, new_n14757_, new_n14758_,
    new_n14759_, new_n14760_, new_n14761_, new_n14762_, new_n14763_,
    new_n14764_, new_n14765_, new_n14766_, new_n14767_, new_n14768_,
    new_n14769_, new_n14770_, new_n14771_, new_n14772_, new_n14773_,
    new_n14774_, new_n14775_, new_n14776_, new_n14777_, new_n14778_,
    new_n14779_, new_n14780_, new_n14781_, new_n14782_, new_n14783_,
    new_n14784_, new_n14785_, new_n14786_, new_n14787_, new_n14788_,
    new_n14789_, new_n14790_, new_n14791_, new_n14792_, new_n14793_,
    new_n14794_, new_n14795_, new_n14796_, new_n14797_, new_n14798_,
    new_n14799_, new_n14800_, new_n14801_, new_n14802_, new_n14803_,
    new_n14804_, new_n14805_, new_n14806_, new_n14807_, new_n14808_,
    new_n14809_, new_n14810_, new_n14811_, new_n14812_, new_n14813_,
    new_n14814_, new_n14815_, new_n14816_, new_n14817_, new_n14818_,
    new_n14819_, new_n14820_, new_n14821_, new_n14822_, new_n14823_,
    new_n14824_, new_n14825_, new_n14826_, new_n14827_, new_n14828_,
    new_n14829_, new_n14830_, new_n14831_, new_n14832_, new_n14833_,
    new_n14835_, new_n14836_, new_n14837_, new_n14838_, new_n14839_,
    new_n14840_, new_n14841_, new_n14842_, new_n14843_, new_n14844_,
    new_n14845_, new_n14846_, new_n14847_, new_n14848_, new_n14849_,
    new_n14850_, new_n14851_, new_n14852_, new_n14853_, new_n14854_,
    new_n14855_, new_n14856_, new_n14857_, new_n14858_, new_n14859_,
    new_n14860_, new_n14861_, new_n14862_, new_n14863_, new_n14864_,
    new_n14865_, new_n14866_, new_n14867_, new_n14868_, new_n14869_,
    new_n14870_, new_n14871_, new_n14872_, new_n14873_, new_n14874_,
    new_n14875_, new_n14876_, new_n14877_, new_n14878_, new_n14879_,
    new_n14880_, new_n14881_, new_n14882_, new_n14883_, new_n14884_,
    new_n14885_, new_n14886_, new_n14887_, new_n14888_, new_n14889_,
    new_n14890_, new_n14891_, new_n14892_, new_n14893_, new_n14894_,
    new_n14895_, new_n14896_, new_n14897_, new_n14898_, new_n14899_,
    new_n14900_, new_n14901_, new_n14902_, new_n14903_, new_n14904_,
    new_n14905_, new_n14906_, new_n14907_, new_n14908_, new_n14909_,
    new_n14910_, new_n14911_, new_n14912_, new_n14913_, new_n14914_,
    new_n14915_, new_n14916_, new_n14917_, new_n14918_, new_n14919_,
    new_n14920_, new_n14921_, new_n14922_, new_n14923_, new_n14924_,
    new_n14925_, new_n14926_, new_n14927_, new_n14928_, new_n14929_,
    new_n14930_, new_n14931_, new_n14932_, new_n14933_, new_n14934_,
    new_n14935_, new_n14936_, new_n14937_, new_n14938_, new_n14939_,
    new_n14940_, new_n14941_, new_n14942_, new_n14943_, new_n14944_,
    new_n14945_, new_n14946_, new_n14947_, new_n14948_, new_n14949_,
    new_n14950_, new_n14951_, new_n14952_, new_n14953_, new_n14954_,
    new_n14955_, new_n14956_, new_n14957_, new_n14958_, new_n14959_,
    new_n14960_, new_n14961_, new_n14962_, new_n14963_, new_n14964_,
    new_n14965_, new_n14966_, new_n14967_, new_n14968_, new_n14969_,
    new_n14970_, new_n14971_, new_n14972_, new_n14973_, new_n14974_,
    new_n14975_, new_n14976_, new_n14977_, new_n14978_, new_n14979_,
    new_n14980_, new_n14981_, new_n14982_, new_n14983_, new_n14984_,
    new_n14985_, new_n14986_, new_n14987_, new_n14988_, new_n14989_,
    new_n14990_, new_n14991_, new_n14992_, new_n14993_, new_n14994_,
    new_n14995_, new_n14996_, new_n14997_, new_n14998_, new_n14999_,
    new_n15000_, new_n15001_, new_n15002_, new_n15003_, new_n15004_,
    new_n15005_, new_n15006_, new_n15007_, new_n15008_, new_n15009_,
    new_n15010_, new_n15011_, new_n15012_, new_n15013_, new_n15014_,
    new_n15015_, new_n15016_, new_n15017_, new_n15018_, new_n15019_,
    new_n15020_, new_n15021_, new_n15022_, new_n15023_, new_n15024_,
    new_n15025_, new_n15026_, new_n15027_, new_n15028_, new_n15029_,
    new_n15030_, new_n15031_, new_n15032_, new_n15033_, new_n15034_,
    new_n15035_, new_n15036_, new_n15037_, new_n15038_, new_n15039_,
    new_n15040_, new_n15041_, new_n15042_, new_n15043_, new_n15044_,
    new_n15045_, new_n15046_, new_n15047_, new_n15048_, new_n15049_,
    new_n15050_, new_n15051_, new_n15052_, new_n15053_, new_n15054_,
    new_n15055_, new_n15056_, new_n15057_, new_n15058_, new_n15059_,
    new_n15060_, new_n15061_, new_n15062_, new_n15063_, new_n15064_,
    new_n15065_, new_n15066_, new_n15067_, new_n15068_, new_n15069_,
    new_n15070_, new_n15071_, new_n15072_, new_n15073_, new_n15074_,
    new_n15075_, new_n15076_, new_n15077_, new_n15078_, new_n15079_,
    new_n15080_, new_n15081_, new_n15082_, new_n15083_, new_n15084_,
    new_n15085_, new_n15086_, new_n15087_, new_n15088_, new_n15089_,
    new_n15090_, new_n15091_, new_n15092_, new_n15093_, new_n15094_,
    new_n15095_, new_n15096_, new_n15097_, new_n15098_, new_n15099_,
    new_n15100_, new_n15101_, new_n15102_, new_n15103_, new_n15104_,
    new_n15105_, new_n15106_, new_n15107_, new_n15108_, new_n15109_,
    new_n15110_, new_n15111_, new_n15112_, new_n15113_, new_n15114_,
    new_n15115_, new_n15116_, new_n15117_, new_n15118_, new_n15119_,
    new_n15120_, new_n15121_, new_n15122_, new_n15123_, new_n15124_,
    new_n15125_, new_n15126_, new_n15127_, new_n15128_, new_n15129_,
    new_n15130_, new_n15131_, new_n15132_, new_n15133_, new_n15134_,
    new_n15135_, new_n15136_, new_n15137_, new_n15138_, new_n15139_,
    new_n15140_, new_n15141_, new_n15142_, new_n15143_, new_n15144_,
    new_n15145_, new_n15146_, new_n15147_, new_n15148_, new_n15149_,
    new_n15150_, new_n15151_, new_n15152_, new_n15153_, new_n15154_,
    new_n15155_, new_n15156_, new_n15157_, new_n15158_, new_n15159_,
    new_n15160_, new_n15161_, new_n15162_, new_n15163_, new_n15164_,
    new_n15165_, new_n15166_, new_n15167_, new_n15168_, new_n15169_,
    new_n15170_, new_n15171_, new_n15172_, new_n15173_, new_n15174_,
    new_n15175_, new_n15176_, new_n15177_, new_n15178_, new_n15179_,
    new_n15180_, new_n15181_, new_n15182_, new_n15183_, new_n15184_,
    new_n15185_, new_n15186_, new_n15187_, new_n15188_, new_n15189_,
    new_n15190_, new_n15191_, new_n15192_, new_n15193_, new_n15194_,
    new_n15195_, new_n15196_, new_n15197_, new_n15198_, new_n15199_,
    new_n15200_, new_n15201_, new_n15202_, new_n15203_, new_n15204_,
    new_n15205_, new_n15206_, new_n15207_, new_n15208_, new_n15209_,
    new_n15210_, new_n15211_, new_n15212_, new_n15213_, new_n15214_,
    new_n15215_, new_n15216_, new_n15217_, new_n15218_, new_n15219_,
    new_n15220_, new_n15221_, new_n15222_, new_n15223_, new_n15224_,
    new_n15225_, new_n15226_, new_n15227_, new_n15228_, new_n15229_,
    new_n15230_, new_n15231_, new_n15232_, new_n15233_, new_n15234_,
    new_n15235_, new_n15236_, new_n15237_, new_n15238_, new_n15239_,
    new_n15240_, new_n15241_, new_n15242_, new_n15243_, new_n15244_,
    new_n15245_, new_n15246_, new_n15247_, new_n15248_, new_n15249_,
    new_n15250_, new_n15251_, new_n15252_, new_n15253_, new_n15254_,
    new_n15255_, new_n15256_, new_n15257_, new_n15258_, new_n15259_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15266_, new_n15267_, new_n15268_, new_n15269_,
    new_n15270_, new_n15271_, new_n15272_, new_n15273_, new_n15274_,
    new_n15275_, new_n15276_, new_n15277_, new_n15278_, new_n15279_,
    new_n15280_, new_n15281_, new_n15282_, new_n15283_, new_n15284_,
    new_n15285_, new_n15286_, new_n15287_, new_n15288_, new_n15289_,
    new_n15290_, new_n15291_, new_n15292_, new_n15293_, new_n15294_,
    new_n15295_, new_n15296_, new_n15297_, new_n15298_, new_n15299_,
    new_n15300_, new_n15301_, new_n15302_, new_n15303_, new_n15304_,
    new_n15305_, new_n15306_, new_n15307_, new_n15308_, new_n15309_,
    new_n15310_, new_n15311_, new_n15312_, new_n15313_, new_n15314_,
    new_n15315_, new_n15316_, new_n15317_, new_n15318_, new_n15319_,
    new_n15320_, new_n15321_, new_n15322_, new_n15323_, new_n15324_,
    new_n15325_, new_n15326_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15334_,
    new_n15335_, new_n15336_, new_n15337_, new_n15338_, new_n15339_,
    new_n15340_, new_n15341_, new_n15342_, new_n15343_, new_n15344_,
    new_n15345_, new_n15346_, new_n15347_, new_n15348_, new_n15349_,
    new_n15350_, new_n15351_, new_n15352_, new_n15353_, new_n15354_,
    new_n15355_, new_n15356_, new_n15357_, new_n15358_, new_n15359_,
    new_n15360_, new_n15361_, new_n15362_, new_n15363_, new_n15364_,
    new_n15365_, new_n15366_, new_n15367_, new_n15368_, new_n15369_,
    new_n15370_, new_n15371_, new_n15372_, new_n15373_, new_n15374_,
    new_n15375_, new_n15376_, new_n15377_, new_n15378_, new_n15379_,
    new_n15380_, new_n15381_, new_n15382_, new_n15383_, new_n15384_,
    new_n15385_, new_n15386_, new_n15387_, new_n15388_, new_n15389_,
    new_n15390_, new_n15391_, new_n15392_, new_n15393_, new_n15394_,
    new_n15395_, new_n15396_, new_n15397_, new_n15398_, new_n15399_,
    new_n15400_, new_n15401_, new_n15402_, new_n15403_, new_n15404_,
    new_n15406_, new_n15407_, new_n15408_, new_n15409_, new_n15410_,
    new_n15411_, new_n15412_, new_n15413_, new_n15414_, new_n15415_,
    new_n15416_, new_n15417_, new_n15418_, new_n15419_, new_n15420_,
    new_n15421_, new_n15422_, new_n15423_, new_n15424_, new_n15425_,
    new_n15426_, new_n15427_, new_n15428_, new_n15429_, new_n15430_,
    new_n15431_, new_n15432_, new_n15433_, new_n15434_, new_n15435_,
    new_n15436_, new_n15437_, new_n15438_, new_n15439_, new_n15440_,
    new_n15441_, new_n15442_, new_n15443_, new_n15444_, new_n15445_,
    new_n15446_, new_n15447_, new_n15448_, new_n15449_, new_n15450_,
    new_n15451_, new_n15452_, new_n15453_, new_n15454_, new_n15455_,
    new_n15456_, new_n15457_, new_n15458_, new_n15459_, new_n15460_,
    new_n15461_, new_n15462_, new_n15463_, new_n15464_, new_n15465_,
    new_n15466_, new_n15467_, new_n15468_, new_n15469_, new_n15470_,
    new_n15471_, new_n15472_, new_n15473_, new_n15474_, new_n15475_,
    new_n15476_, new_n15477_, new_n15478_, new_n15479_, new_n15480_,
    new_n15481_, new_n15482_, new_n15483_, new_n15484_, new_n15485_,
    new_n15486_, new_n15487_, new_n15488_, new_n15489_, new_n15490_,
    new_n15491_, new_n15492_, new_n15493_, new_n15494_, new_n15495_,
    new_n15496_, new_n15497_, new_n15498_, new_n15499_, new_n15500_,
    new_n15501_, new_n15502_, new_n15503_, new_n15504_, new_n15505_,
    new_n15506_, new_n15507_, new_n15508_, new_n15509_, new_n15510_,
    new_n15511_, new_n15512_, new_n15513_, new_n15514_, new_n15515_,
    new_n15516_, new_n15517_, new_n15518_, new_n15519_, new_n15520_,
    new_n15521_, new_n15522_, new_n15523_, new_n15524_, new_n15525_,
    new_n15526_, new_n15527_, new_n15528_, new_n15529_, new_n15530_,
    new_n15531_, new_n15532_, new_n15533_, new_n15534_, new_n15535_,
    new_n15536_, new_n15537_, new_n15538_, new_n15539_, new_n15540_,
    new_n15541_, new_n15542_, new_n15543_, new_n15544_, new_n15545_,
    new_n15546_, new_n15547_, new_n15548_, new_n15549_, new_n15550_,
    new_n15551_, new_n15552_, new_n15553_, new_n15554_, new_n15555_,
    new_n15556_, new_n15557_, new_n15558_, new_n15559_, new_n15560_,
    new_n15561_, new_n15562_, new_n15563_, new_n15564_, new_n15565_,
    new_n15566_, new_n15567_, new_n15568_, new_n15569_, new_n15570_,
    new_n15571_, new_n15572_, new_n15573_, new_n15574_, new_n15575_,
    new_n15576_, new_n15577_, new_n15578_, new_n15579_, new_n15580_,
    new_n15581_, new_n15582_, new_n15583_, new_n15584_, new_n15585_,
    new_n15586_, new_n15587_, new_n15588_, new_n15589_, new_n15590_,
    new_n15591_, new_n15592_, new_n15593_, new_n15594_, new_n15595_,
    new_n15596_, new_n15597_, new_n15598_, new_n15599_, new_n15600_,
    new_n15601_, new_n15602_, new_n15603_, new_n15604_, new_n15605_,
    new_n15606_, new_n15607_, new_n15608_, new_n15609_, new_n15610_,
    new_n15611_, new_n15612_, new_n15613_, new_n15614_, new_n15615_,
    new_n15616_, new_n15617_, new_n15618_, new_n15619_, new_n15620_,
    new_n15621_, new_n15622_, new_n15623_, new_n15624_, new_n15625_,
    new_n15626_, new_n15627_, new_n15628_, new_n15629_, new_n15630_,
    new_n15631_, new_n15632_, new_n15633_, new_n15634_, new_n15635_,
    new_n15636_, new_n15637_, new_n15638_, new_n15639_, new_n15640_,
    new_n15641_, new_n15642_, new_n15643_, new_n15644_, new_n15645_,
    new_n15646_, new_n15647_, new_n15648_, new_n15649_, new_n15650_,
    new_n15651_, new_n15652_, new_n15653_, new_n15654_, new_n15655_,
    new_n15656_, new_n15657_, new_n15658_, new_n15659_, new_n15660_,
    new_n15661_, new_n15662_, new_n15663_, new_n15664_, new_n15665_,
    new_n15666_, new_n15667_, new_n15668_, new_n15669_, new_n15670_,
    new_n15671_, new_n15672_, new_n15673_, new_n15674_, new_n15675_,
    new_n15676_, new_n15677_, new_n15678_, new_n15679_, new_n15680_,
    new_n15681_, new_n15682_, new_n15683_, new_n15684_, new_n15685_,
    new_n15686_, new_n15687_, new_n15688_, new_n15689_, new_n15690_,
    new_n15691_, new_n15692_, new_n15693_, new_n15694_, new_n15695_,
    new_n15696_, new_n15697_, new_n15698_, new_n15699_, new_n15700_,
    new_n15701_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15741_, new_n15742_, new_n15743_, new_n15744_, new_n15745_,
    new_n15746_, new_n15747_, new_n15748_, new_n15749_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15781_, new_n15782_, new_n15783_, new_n15784_, new_n15785_,
    new_n15786_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15797_, new_n15798_, new_n15799_, new_n15800_,
    new_n15801_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15840_,
    new_n15841_, new_n15842_, new_n15843_, new_n15844_, new_n15845_,
    new_n15846_, new_n15847_, new_n15848_, new_n15849_, new_n15850_,
    new_n15851_, new_n15852_, new_n15853_, new_n15854_, new_n15855_,
    new_n15856_, new_n15857_, new_n15858_, new_n15859_, new_n15860_,
    new_n15861_, new_n15862_, new_n15863_, new_n15864_, new_n15865_,
    new_n15866_, new_n15867_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15879_, new_n15880_,
    new_n15881_, new_n15882_, new_n15883_, new_n15884_, new_n15885_,
    new_n15886_, new_n15887_, new_n15888_, new_n15889_, new_n15890_,
    new_n15891_, new_n15892_, new_n15893_, new_n15894_, new_n15895_,
    new_n15896_, new_n15897_, new_n15898_, new_n15899_, new_n15900_,
    new_n15901_, new_n15902_, new_n15903_, new_n15904_, new_n15905_,
    new_n15906_, new_n15907_, new_n15908_, new_n15909_, new_n15910_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15916_, new_n15917_, new_n15918_, new_n15919_, new_n15920_,
    new_n15921_, new_n15922_, new_n15923_, new_n15924_, new_n15925_,
    new_n15926_, new_n15927_, new_n15928_, new_n15929_, new_n15930_,
    new_n15931_, new_n15932_, new_n15933_, new_n15934_, new_n15935_,
    new_n15936_, new_n15937_, new_n15938_, new_n15939_, new_n15940_,
    new_n15941_, new_n15942_, new_n15943_, new_n15944_, new_n15945_,
    new_n15946_, new_n15947_, new_n15948_, new_n15949_, new_n15950_,
    new_n15951_, new_n15952_, new_n15953_, new_n15954_, new_n15955_,
    new_n15956_, new_n15957_, new_n15958_, new_n15959_, new_n15960_,
    new_n15961_, new_n15962_, new_n15963_, new_n15964_, new_n15965_,
    new_n15966_, new_n15967_, new_n15968_, new_n15969_, new_n15970_,
    new_n15971_, new_n15972_, new_n15973_, new_n15974_, new_n15975_,
    new_n15976_, new_n15977_, new_n15978_, new_n15979_, new_n15980_,
    new_n15981_, new_n15982_, new_n15983_, new_n15984_, new_n15985_,
    new_n15986_, new_n15987_, new_n15988_, new_n15989_, new_n15990_,
    new_n15991_, new_n15992_, new_n15993_, new_n15994_, new_n15995_,
    new_n15996_, new_n15997_, new_n15998_, new_n15999_, new_n16000_,
    new_n16001_, new_n16002_, new_n16003_, new_n16004_, new_n16005_,
    new_n16006_, new_n16007_, new_n16008_, new_n16009_, new_n16010_,
    new_n16011_, new_n16012_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16024_, new_n16025_, new_n16026_,
    new_n16027_, new_n16028_, new_n16029_, new_n16030_, new_n16031_,
    new_n16032_, new_n16033_, new_n16034_, new_n16035_, new_n16036_,
    new_n16037_, new_n16038_, new_n16039_, new_n16040_, new_n16041_,
    new_n16042_, new_n16043_, new_n16044_, new_n16045_, new_n16046_,
    new_n16047_, new_n16048_, new_n16049_, new_n16050_, new_n16051_,
    new_n16052_, new_n16053_, new_n16054_, new_n16055_, new_n16056_,
    new_n16057_, new_n16058_, new_n16059_, new_n16060_, new_n16061_,
    new_n16062_, new_n16063_, new_n16064_, new_n16065_, new_n16066_,
    new_n16067_, new_n16068_, new_n16069_, new_n16070_, new_n16071_,
    new_n16072_, new_n16073_, new_n16074_, new_n16075_, new_n16076_,
    new_n16077_, new_n16078_, new_n16079_, new_n16080_, new_n16081_,
    new_n16082_, new_n16083_, new_n16084_, new_n16085_, new_n16086_,
    new_n16087_, new_n16088_, new_n16089_, new_n16090_, new_n16091_,
    new_n16092_, new_n16093_, new_n16094_, new_n16095_, new_n16096_,
    new_n16097_, new_n16098_, new_n16099_, new_n16100_, new_n16101_,
    new_n16102_, new_n16103_, new_n16104_, new_n16105_, new_n16106_,
    new_n16107_, new_n16108_, new_n16109_, new_n16110_, new_n16111_,
    new_n16112_, new_n16113_, new_n16114_, new_n16115_, new_n16116_,
    new_n16117_, new_n16118_, new_n16119_, new_n16120_, new_n16121_,
    new_n16122_, new_n16123_, new_n16124_, new_n16125_, new_n16126_,
    new_n16127_, new_n16128_, new_n16129_, new_n16130_, new_n16131_,
    new_n16132_, new_n16133_, new_n16134_, new_n16135_, new_n16136_,
    new_n16137_, new_n16138_, new_n16139_, new_n16140_, new_n16141_,
    new_n16142_, new_n16143_, new_n16144_, new_n16145_, new_n16146_,
    new_n16147_, new_n16148_, new_n16149_, new_n16150_, new_n16151_,
    new_n16152_, new_n16153_, new_n16154_, new_n16155_, new_n16156_,
    new_n16157_, new_n16158_, new_n16159_, new_n16160_, new_n16161_,
    new_n16162_, new_n16163_, new_n16164_, new_n16165_, new_n16166_,
    new_n16167_, new_n16168_, new_n16169_, new_n16170_, new_n16171_,
    new_n16172_, new_n16173_, new_n16174_, new_n16175_, new_n16176_,
    new_n16177_, new_n16178_, new_n16179_, new_n16180_, new_n16181_,
    new_n16182_, new_n16183_, new_n16184_, new_n16185_, new_n16186_,
    new_n16187_, new_n16188_, new_n16189_, new_n16190_, new_n16191_,
    new_n16192_, new_n16193_, new_n16194_, new_n16195_, new_n16196_,
    new_n16197_, new_n16198_, new_n16199_, new_n16200_, new_n16201_,
    new_n16202_, new_n16203_, new_n16204_, new_n16205_, new_n16206_,
    new_n16207_, new_n16208_, new_n16209_, new_n16210_, new_n16211_,
    new_n16212_, new_n16213_, new_n16214_, new_n16215_, new_n16216_,
    new_n16217_, new_n16218_, new_n16219_, new_n16220_, new_n16221_,
    new_n16222_, new_n16223_, new_n16224_, new_n16225_, new_n16226_,
    new_n16227_, new_n16228_, new_n16229_, new_n16230_, new_n16231_,
    new_n16232_, new_n16233_, new_n16234_, new_n16235_, new_n16236_,
    new_n16237_, new_n16238_, new_n16239_, new_n16240_, new_n16241_,
    new_n16242_, new_n16243_, new_n16244_, new_n16245_, new_n16246_,
    new_n16247_, new_n16248_, new_n16249_, new_n16250_, new_n16251_,
    new_n16252_, new_n16253_, new_n16254_, new_n16255_, new_n16256_,
    new_n16257_, new_n16258_, new_n16259_, new_n16260_, new_n16261_,
    new_n16262_, new_n16263_, new_n16264_, new_n16265_, new_n16266_,
    new_n16267_, new_n16268_, new_n16269_, new_n16270_, new_n16271_,
    new_n16272_, new_n16273_, new_n16274_, new_n16275_, new_n16276_,
    new_n16277_, new_n16278_, new_n16279_, new_n16280_, new_n16281_,
    new_n16282_, new_n16283_, new_n16284_, new_n16285_, new_n16286_,
    new_n16287_, new_n16288_, new_n16289_, new_n16290_, new_n16291_,
    new_n16292_, new_n16293_, new_n16294_, new_n16295_, new_n16296_,
    new_n16297_, new_n16298_, new_n16299_, new_n16300_, new_n16301_,
    new_n16302_, new_n16303_, new_n16304_, new_n16305_, new_n16306_,
    new_n16307_, new_n16308_, new_n16309_, new_n16310_, new_n16311_,
    new_n16312_, new_n16313_, new_n16314_, new_n16315_, new_n16316_,
    new_n16317_, new_n16318_, new_n16319_, new_n16320_, new_n16321_,
    new_n16322_, new_n16323_, new_n16324_, new_n16325_, new_n16326_,
    new_n16327_, new_n16328_, new_n16329_, new_n16330_, new_n16331_,
    new_n16332_, new_n16333_, new_n16334_, new_n16335_, new_n16336_,
    new_n16337_, new_n16338_, new_n16339_, new_n16340_, new_n16341_,
    new_n16342_, new_n16343_, new_n16344_, new_n16345_, new_n16346_,
    new_n16347_, new_n16348_, new_n16349_, new_n16350_, new_n16351_,
    new_n16352_, new_n16353_, new_n16354_, new_n16355_, new_n16356_,
    new_n16357_, new_n16358_, new_n16359_, new_n16360_, new_n16361_,
    new_n16362_, new_n16363_, new_n16364_, new_n16365_, new_n16366_,
    new_n16367_, new_n16368_, new_n16369_, new_n16370_, new_n16371_,
    new_n16372_, new_n16373_, new_n16374_, new_n16375_, new_n16376_,
    new_n16377_, new_n16378_, new_n16379_, new_n16380_, new_n16381_,
    new_n16382_, new_n16383_, new_n16384_, new_n16385_, new_n16386_,
    new_n16387_, new_n16388_, new_n16389_, new_n16390_, new_n16391_,
    new_n16392_, new_n16393_, new_n16394_, new_n16395_, new_n16396_,
    new_n16397_, new_n16398_, new_n16399_, new_n16400_, new_n16401_,
    new_n16402_, new_n16403_, new_n16404_, new_n16405_, new_n16406_,
    new_n16407_, new_n16408_, new_n16409_, new_n16410_, new_n16411_,
    new_n16412_, new_n16413_, new_n16414_, new_n16415_, new_n16416_,
    new_n16417_, new_n16418_, new_n16419_, new_n16420_, new_n16421_,
    new_n16422_, new_n16423_, new_n16424_, new_n16425_, new_n16426_,
    new_n16427_, new_n16428_, new_n16429_, new_n16430_, new_n16431_,
    new_n16432_, new_n16433_, new_n16434_, new_n16435_, new_n16436_,
    new_n16437_, new_n16438_, new_n16439_, new_n16440_, new_n16441_,
    new_n16442_, new_n16443_, new_n16444_, new_n16445_, new_n16446_,
    new_n16447_, new_n16448_, new_n16449_, new_n16450_, new_n16451_,
    new_n16452_, new_n16453_, new_n16454_, new_n16455_, new_n16456_,
    new_n16457_, new_n16458_, new_n16459_, new_n16460_, new_n16461_,
    new_n16462_, new_n16463_, new_n16464_, new_n16465_, new_n16466_,
    new_n16467_, new_n16468_, new_n16469_, new_n16470_, new_n16471_,
    new_n16472_, new_n16473_, new_n16474_, new_n16475_, new_n16476_,
    new_n16477_, new_n16478_, new_n16479_, new_n16480_, new_n16481_,
    new_n16482_, new_n16483_, new_n16484_, new_n16485_, new_n16486_,
    new_n16487_, new_n16488_, new_n16489_, new_n16490_, new_n16491_,
    new_n16492_, new_n16493_, new_n16494_, new_n16495_, new_n16496_,
    new_n16497_, new_n16498_, new_n16499_, new_n16500_, new_n16501_,
    new_n16502_, new_n16503_, new_n16504_, new_n16505_, new_n16506_,
    new_n16507_, new_n16508_, new_n16509_, new_n16510_, new_n16511_,
    new_n16512_, new_n16513_, new_n16514_, new_n16515_, new_n16516_,
    new_n16517_, new_n16518_, new_n16519_, new_n16520_, new_n16521_,
    new_n16522_, new_n16523_, new_n16524_, new_n16525_, new_n16526_,
    new_n16527_, new_n16528_, new_n16529_, new_n16530_, new_n16531_,
    new_n16532_, new_n16533_, new_n16534_, new_n16535_, new_n16536_,
    new_n16537_, new_n16538_, new_n16539_, new_n16540_, new_n16541_,
    new_n16542_, new_n16543_, new_n16544_, new_n16545_, new_n16546_,
    new_n16547_, new_n16548_, new_n16549_, new_n16550_, new_n16551_,
    new_n16552_, new_n16553_, new_n16554_, new_n16555_, new_n16556_,
    new_n16557_, new_n16558_, new_n16559_, new_n16560_, new_n16561_,
    new_n16562_, new_n16563_, new_n16564_, new_n16565_, new_n16566_,
    new_n16567_, new_n16568_, new_n16569_, new_n16570_, new_n16571_,
    new_n16572_, new_n16573_, new_n16574_, new_n16575_, new_n16576_,
    new_n16577_, new_n16578_, new_n16579_, new_n16580_, new_n16581_,
    new_n16582_, new_n16583_, new_n16584_, new_n16585_, new_n16586_,
    new_n16587_, new_n16588_, new_n16589_, new_n16590_, new_n16591_,
    new_n16592_, new_n16593_, new_n16594_, new_n16595_, new_n16596_,
    new_n16597_, new_n16598_, new_n16599_, new_n16600_, new_n16601_,
    new_n16602_, new_n16603_, new_n16604_, new_n16605_, new_n16606_,
    new_n16607_, new_n16608_, new_n16609_, new_n16610_, new_n16611_,
    new_n16612_, new_n16613_, new_n16614_, new_n16615_, new_n16616_,
    new_n16617_, new_n16618_, new_n16619_, new_n16620_, new_n16621_,
    new_n16622_, new_n16623_, new_n16624_, new_n16625_, new_n16626_,
    new_n16627_, new_n16628_, new_n16629_, new_n16630_, new_n16631_,
    new_n16632_, new_n16633_, new_n16635_, new_n16636_, new_n16637_,
    new_n16638_, new_n16639_, new_n16640_, new_n16641_, new_n16642_,
    new_n16643_, new_n16644_, new_n16645_, new_n16646_, new_n16647_,
    new_n16648_, new_n16649_, new_n16650_, new_n16651_, new_n16652_,
    new_n16653_, new_n16654_, new_n16655_, new_n16656_, new_n16657_,
    new_n16658_, new_n16659_, new_n16660_, new_n16661_, new_n16662_,
    new_n16663_, new_n16664_, new_n16665_, new_n16666_, new_n16667_,
    new_n16668_, new_n16669_, new_n16670_, new_n16671_, new_n16672_,
    new_n16673_, new_n16674_, new_n16675_, new_n16676_, new_n16677_,
    new_n16678_, new_n16679_, new_n16680_, new_n16681_, new_n16682_,
    new_n16683_, new_n16684_, new_n16685_, new_n16686_, new_n16687_,
    new_n16688_, new_n16689_, new_n16690_, new_n16691_, new_n16692_,
    new_n16693_, new_n16694_, new_n16695_, new_n16696_, new_n16697_,
    new_n16698_, new_n16699_, new_n16700_, new_n16701_, new_n16702_,
    new_n16703_, new_n16704_, new_n16705_, new_n16706_, new_n16707_,
    new_n16708_, new_n16709_, new_n16710_, new_n16711_, new_n16712_,
    new_n16713_, new_n16714_, new_n16715_, new_n16716_, new_n16717_,
    new_n16718_, new_n16719_, new_n16720_, new_n16721_, new_n16722_,
    new_n16723_, new_n16724_, new_n16725_, new_n16726_, new_n16727_,
    new_n16728_, new_n16729_, new_n16730_, new_n16731_, new_n16732_,
    new_n16733_, new_n16734_, new_n16735_, new_n16736_, new_n16737_,
    new_n16738_, new_n16739_, new_n16740_, new_n16741_, new_n16742_,
    new_n16743_, new_n16744_, new_n16745_, new_n16746_, new_n16747_,
    new_n16748_, new_n16749_, new_n16750_, new_n16751_, new_n16752_,
    new_n16753_, new_n16754_, new_n16755_, new_n16756_, new_n16757_,
    new_n16758_, new_n16759_, new_n16760_, new_n16761_, new_n16762_,
    new_n16763_, new_n16764_, new_n16765_, new_n16766_, new_n16767_,
    new_n16768_, new_n16769_, new_n16770_, new_n16771_, new_n16772_,
    new_n16773_, new_n16774_, new_n16775_, new_n16776_, new_n16777_,
    new_n16778_, new_n16779_, new_n16780_, new_n16781_, new_n16782_,
    new_n16783_, new_n16784_, new_n16785_, new_n16786_, new_n16787_,
    new_n16788_, new_n16789_, new_n16790_, new_n16791_, new_n16792_,
    new_n16793_, new_n16794_, new_n16795_, new_n16796_, new_n16797_,
    new_n16798_, new_n16799_, new_n16800_, new_n16801_, new_n16802_,
    new_n16803_, new_n16804_, new_n16805_, new_n16806_, new_n16807_,
    new_n16808_, new_n16809_, new_n16810_, new_n16811_, new_n16812_,
    new_n16813_, new_n16814_, new_n16815_, new_n16816_, new_n16817_,
    new_n16818_, new_n16819_, new_n16820_, new_n16821_, new_n16822_,
    new_n16823_, new_n16824_, new_n16825_, new_n16826_, new_n16827_,
    new_n16828_, new_n16829_, new_n16830_, new_n16831_, new_n16832_,
    new_n16833_, new_n16834_, new_n16835_, new_n16836_, new_n16837_,
    new_n16838_, new_n16839_, new_n16840_, new_n16841_, new_n16842_,
    new_n16843_, new_n16844_, new_n16845_, new_n16846_, new_n16847_,
    new_n16848_, new_n16849_, new_n16850_, new_n16851_, new_n16852_,
    new_n16853_, new_n16854_, new_n16855_, new_n16856_, new_n16857_,
    new_n16858_, new_n16859_, new_n16860_, new_n16861_, new_n16862_,
    new_n16863_, new_n16864_, new_n16865_, new_n16866_, new_n16867_,
    new_n16868_, new_n16869_, new_n16870_, new_n16871_, new_n16872_,
    new_n16873_, new_n16874_, new_n16875_, new_n16876_, new_n16877_,
    new_n16878_, new_n16879_, new_n16880_, new_n16881_, new_n16882_,
    new_n16883_, new_n16884_, new_n16885_, new_n16886_, new_n16887_,
    new_n16888_, new_n16889_, new_n16890_, new_n16891_, new_n16892_,
    new_n16893_, new_n16894_, new_n16895_, new_n16896_, new_n16897_,
    new_n16898_, new_n16899_, new_n16900_, new_n16901_, new_n16902_,
    new_n16903_, new_n16904_, new_n16905_, new_n16906_, new_n16907_,
    new_n16908_, new_n16909_, new_n16910_, new_n16911_, new_n16912_,
    new_n16913_, new_n16914_, new_n16915_, new_n16916_, new_n16917_,
    new_n16918_, new_n16919_, new_n16920_, new_n16921_, new_n16922_,
    new_n16923_, new_n16924_, new_n16925_, new_n16926_, new_n16927_,
    new_n16928_, new_n16929_, new_n16930_, new_n16931_, new_n16932_,
    new_n16933_, new_n16934_, new_n16935_, new_n16936_, new_n16937_,
    new_n16938_, new_n16939_, new_n16940_, new_n16941_, new_n16942_,
    new_n16943_, new_n16944_, new_n16945_, new_n16946_, new_n16947_,
    new_n16948_, new_n16949_, new_n16950_, new_n16951_, new_n16952_,
    new_n16953_, new_n16954_, new_n16955_, new_n16956_, new_n16957_,
    new_n16958_, new_n16959_, new_n16960_, new_n16961_, new_n16962_,
    new_n16963_, new_n16964_, new_n16965_, new_n16966_, new_n16967_,
    new_n16968_, new_n16969_, new_n16970_, new_n16971_, new_n16972_,
    new_n16973_, new_n16974_, new_n16975_, new_n16976_, new_n16977_,
    new_n16978_, new_n16979_, new_n16980_, new_n16981_, new_n16982_,
    new_n16983_, new_n16984_, new_n16985_, new_n16986_, new_n16987_,
    new_n16988_, new_n16989_, new_n16990_, new_n16991_, new_n16992_,
    new_n16993_, new_n16994_, new_n16995_, new_n16996_, new_n16997_,
    new_n16998_, new_n16999_, new_n17000_, new_n17001_, new_n17002_,
    new_n17003_, new_n17004_, new_n17005_, new_n17006_, new_n17007_,
    new_n17008_, new_n17009_, new_n17010_, new_n17011_, new_n17012_,
    new_n17013_, new_n17014_, new_n17015_, new_n17016_, new_n17017_,
    new_n17018_, new_n17019_, new_n17020_, new_n17021_, new_n17022_,
    new_n17023_, new_n17024_, new_n17025_, new_n17026_, new_n17027_,
    new_n17028_, new_n17029_, new_n17030_, new_n17031_, new_n17032_,
    new_n17033_, new_n17034_, new_n17035_, new_n17036_, new_n17037_,
    new_n17038_, new_n17039_, new_n17040_, new_n17041_, new_n17042_,
    new_n17043_, new_n17044_, new_n17045_, new_n17046_, new_n17047_,
    new_n17048_, new_n17049_, new_n17050_, new_n17051_, new_n17052_,
    new_n17053_, new_n17054_, new_n17055_, new_n17056_, new_n17057_,
    new_n17058_, new_n17059_, new_n17060_, new_n17061_, new_n17062_,
    new_n17063_, new_n17064_, new_n17065_, new_n17066_, new_n17067_,
    new_n17068_, new_n17069_, new_n17070_, new_n17071_, new_n17072_,
    new_n17073_, new_n17074_, new_n17075_, new_n17076_, new_n17077_,
    new_n17078_, new_n17079_, new_n17080_, new_n17081_, new_n17082_,
    new_n17083_, new_n17084_, new_n17085_, new_n17086_, new_n17087_,
    new_n17088_, new_n17089_, new_n17090_, new_n17091_, new_n17092_,
    new_n17093_, new_n17094_, new_n17095_, new_n17096_, new_n17097_,
    new_n17098_, new_n17099_, new_n17100_, new_n17101_, new_n17102_,
    new_n17103_, new_n17104_, new_n17105_, new_n17106_, new_n17107_,
    new_n17108_, new_n17109_, new_n17110_, new_n17111_, new_n17112_,
    new_n17113_, new_n17114_, new_n17115_, new_n17116_, new_n17117_,
    new_n17118_, new_n17119_, new_n17120_, new_n17121_, new_n17122_,
    new_n17123_, new_n17124_, new_n17125_, new_n17126_, new_n17127_,
    new_n17128_, new_n17129_, new_n17130_, new_n17131_, new_n17132_,
    new_n17133_, new_n17134_, new_n17135_, new_n17136_, new_n17137_,
    new_n17138_, new_n17139_, new_n17140_, new_n17141_, new_n17142_,
    new_n17143_, new_n17144_, new_n17145_, new_n17146_, new_n17147_,
    new_n17148_, new_n17149_, new_n17150_, new_n17151_, new_n17152_,
    new_n17153_, new_n17154_, new_n17155_, new_n17156_, new_n17157_,
    new_n17158_, new_n17159_, new_n17160_, new_n17161_, new_n17162_,
    new_n17163_, new_n17164_, new_n17165_, new_n17166_, new_n17167_,
    new_n17168_, new_n17169_, new_n17170_, new_n17171_, new_n17172_,
    new_n17173_, new_n17174_, new_n17175_, new_n17176_, new_n17177_,
    new_n17178_, new_n17179_, new_n17180_, new_n17181_, new_n17182_,
    new_n17183_, new_n17184_, new_n17185_, new_n17186_, new_n17187_,
    new_n17188_, new_n17189_, new_n17190_, new_n17191_, new_n17192_,
    new_n17193_, new_n17194_, new_n17195_, new_n17196_, new_n17197_,
    new_n17198_, new_n17199_, new_n17200_, new_n17201_, new_n17202_,
    new_n17203_, new_n17204_, new_n17205_, new_n17206_, new_n17207_,
    new_n17208_, new_n17209_, new_n17210_, new_n17211_, new_n17212_,
    new_n17213_, new_n17214_, new_n17215_, new_n17216_, new_n17217_,
    new_n17218_, new_n17219_, new_n17220_, new_n17221_, new_n17222_,
    new_n17223_, new_n17224_, new_n17225_, new_n17226_, new_n17227_,
    new_n17228_, new_n17229_, new_n17230_, new_n17231_, new_n17233_,
    new_n17234_, new_n17235_, new_n17236_, new_n17237_, new_n17238_,
    new_n17239_, new_n17240_, new_n17241_, new_n17242_, new_n17243_,
    new_n17244_, new_n17245_, new_n17246_, new_n17247_, new_n17248_,
    new_n17249_, new_n17250_, new_n17251_, new_n17252_, new_n17253_,
    new_n17254_, new_n17255_, new_n17256_, new_n17257_, new_n17258_,
    new_n17259_, new_n17260_, new_n17261_, new_n17262_, new_n17263_,
    new_n17264_, new_n17265_, new_n17266_, new_n17267_, new_n17268_,
    new_n17269_, new_n17270_, new_n17271_, new_n17272_, new_n17273_,
    new_n17274_, new_n17275_, new_n17276_, new_n17277_, new_n17278_,
    new_n17279_, new_n17280_, new_n17281_, new_n17282_, new_n17283_,
    new_n17284_, new_n17285_, new_n17286_, new_n17287_, new_n17288_,
    new_n17289_, new_n17290_, new_n17291_, new_n17292_, new_n17293_,
    new_n17294_, new_n17295_, new_n17296_, new_n17297_, new_n17298_,
    new_n17299_, new_n17300_, new_n17301_, new_n17302_, new_n17303_,
    new_n17304_, new_n17305_, new_n17306_, new_n17307_, new_n17308_,
    new_n17309_, new_n17310_, new_n17311_, new_n17312_, new_n17313_,
    new_n17314_, new_n17315_, new_n17316_, new_n17317_, new_n17318_,
    new_n17319_, new_n17320_, new_n17321_, new_n17322_, new_n17323_,
    new_n17324_, new_n17325_, new_n17326_, new_n17327_, new_n17328_,
    new_n17329_, new_n17330_, new_n17331_, new_n17332_, new_n17333_,
    new_n17334_, new_n17335_, new_n17336_, new_n17337_, new_n17338_,
    new_n17339_, new_n17340_, new_n17341_, new_n17342_, new_n17343_,
    new_n17344_, new_n17345_, new_n17346_, new_n17347_, new_n17348_,
    new_n17349_, new_n17350_, new_n17351_, new_n17352_, new_n17353_,
    new_n17354_, new_n17355_, new_n17356_, new_n17357_, new_n17358_,
    new_n17359_, new_n17360_, new_n17361_, new_n17362_, new_n17363_,
    new_n17364_, new_n17365_, new_n17366_, new_n17367_, new_n17368_,
    new_n17369_, new_n17370_, new_n17371_, new_n17372_, new_n17373_,
    new_n17374_, new_n17375_, new_n17376_, new_n17377_, new_n17378_,
    new_n17379_, new_n17380_, new_n17381_, new_n17382_, new_n17383_,
    new_n17384_, new_n17385_, new_n17386_, new_n17387_, new_n17388_,
    new_n17389_, new_n17390_, new_n17391_, new_n17392_, new_n17393_,
    new_n17394_, new_n17395_, new_n17396_, new_n17397_, new_n17398_,
    new_n17399_, new_n17400_, new_n17401_, new_n17402_, new_n17403_,
    new_n17404_, new_n17405_, new_n17406_, new_n17407_, new_n17408_,
    new_n17409_, new_n17410_, new_n17411_, new_n17412_, new_n17413_,
    new_n17414_, new_n17415_, new_n17416_, new_n17417_, new_n17418_,
    new_n17419_, new_n17420_, new_n17421_, new_n17422_, new_n17423_,
    new_n17424_, new_n17425_, new_n17426_, new_n17427_, new_n17428_,
    new_n17429_, new_n17430_, new_n17431_, new_n17432_, new_n17433_,
    new_n17434_, new_n17435_, new_n17436_, new_n17437_, new_n17438_,
    new_n17439_, new_n17440_, new_n17441_, new_n17442_, new_n17443_,
    new_n17444_, new_n17445_, new_n17446_, new_n17447_, new_n17448_,
    new_n17449_, new_n17450_, new_n17451_, new_n17452_, new_n17453_,
    new_n17454_, new_n17455_, new_n17456_, new_n17457_, new_n17458_,
    new_n17459_, new_n17460_, new_n17461_, new_n17462_, new_n17463_,
    new_n17464_, new_n17465_, new_n17466_, new_n17467_, new_n17468_,
    new_n17469_, new_n17470_, new_n17471_, new_n17472_, new_n17473_,
    new_n17474_, new_n17475_, new_n17476_, new_n17477_, new_n17478_,
    new_n17479_, new_n17480_, new_n17481_, new_n17482_, new_n17483_,
    new_n17484_, new_n17485_, new_n17486_, new_n17487_, new_n17488_,
    new_n17489_, new_n17490_, new_n17491_, new_n17492_, new_n17493_,
    new_n17494_, new_n17495_, new_n17496_, new_n17497_, new_n17498_,
    new_n17499_, new_n17500_, new_n17501_, new_n17502_, new_n17503_,
    new_n17504_, new_n17505_, new_n17506_, new_n17507_, new_n17508_,
    new_n17509_, new_n17510_, new_n17511_, new_n17512_, new_n17513_,
    new_n17514_, new_n17515_, new_n17516_, new_n17517_, new_n17518_,
    new_n17519_, new_n17520_, new_n17521_, new_n17522_, new_n17523_,
    new_n17524_, new_n17525_, new_n17526_, new_n17527_, new_n17528_,
    new_n17529_, new_n17530_, new_n17531_, new_n17532_, new_n17533_,
    new_n17534_, new_n17535_, new_n17536_, new_n17537_, new_n17538_,
    new_n17539_, new_n17540_, new_n17541_, new_n17542_, new_n17543_,
    new_n17544_, new_n17545_, new_n17546_, new_n17547_, new_n17548_,
    new_n17549_, new_n17550_, new_n17551_, new_n17552_, new_n17553_,
    new_n17554_, new_n17555_, new_n17556_, new_n17557_, new_n17558_,
    new_n17559_, new_n17560_, new_n17561_, new_n17562_, new_n17563_,
    new_n17564_, new_n17565_, new_n17566_, new_n17567_, new_n17568_,
    new_n17569_, new_n17570_, new_n17571_, new_n17572_, new_n17573_,
    new_n17574_, new_n17575_, new_n17576_, new_n17577_, new_n17578_,
    new_n17579_, new_n17580_, new_n17581_, new_n17582_, new_n17583_,
    new_n17584_, new_n17585_, new_n17586_, new_n17587_, new_n17588_,
    new_n17589_, new_n17590_, new_n17591_, new_n17592_, new_n17593_,
    new_n17594_, new_n17595_, new_n17596_, new_n17597_, new_n17598_,
    new_n17599_, new_n17600_, new_n17601_, new_n17602_, new_n17603_,
    new_n17604_, new_n17605_, new_n17606_, new_n17607_, new_n17608_,
    new_n17609_, new_n17610_, new_n17611_, new_n17612_, new_n17613_,
    new_n17614_, new_n17615_, new_n17616_, new_n17617_, new_n17618_,
    new_n17619_, new_n17620_, new_n17621_, new_n17622_, new_n17623_,
    new_n17624_, new_n17625_, new_n17626_, new_n17627_, new_n17628_,
    new_n17629_, new_n17630_, new_n17631_, new_n17632_, new_n17633_,
    new_n17634_, new_n17635_, new_n17636_, new_n17637_, new_n17638_,
    new_n17639_, new_n17640_, new_n17641_, new_n17642_, new_n17643_,
    new_n17644_, new_n17645_, new_n17646_, new_n17647_, new_n17648_,
    new_n17649_, new_n17650_, new_n17651_, new_n17652_, new_n17653_,
    new_n17654_, new_n17655_, new_n17656_, new_n17657_, new_n17658_,
    new_n17659_, new_n17660_, new_n17661_, new_n17662_, new_n17663_,
    new_n17664_, new_n17665_, new_n17666_, new_n17667_, new_n17668_,
    new_n17669_, new_n17670_, new_n17671_, new_n17672_, new_n17673_,
    new_n17674_, new_n17675_, new_n17676_, new_n17677_, new_n17678_,
    new_n17679_, new_n17680_, new_n17681_, new_n17682_, new_n17683_,
    new_n17684_, new_n17685_, new_n17686_, new_n17687_, new_n17688_,
    new_n17689_, new_n17690_, new_n17691_, new_n17692_, new_n17693_,
    new_n17694_, new_n17695_, new_n17696_, new_n17697_, new_n17698_,
    new_n17699_, new_n17700_, new_n17701_, new_n17702_, new_n17703_,
    new_n17704_, new_n17705_, new_n17706_, new_n17707_, new_n17708_,
    new_n17709_, new_n17710_, new_n17711_, new_n17712_, new_n17713_,
    new_n17714_, new_n17715_, new_n17716_, new_n17717_, new_n17718_,
    new_n17719_, new_n17720_, new_n17721_, new_n17722_, new_n17723_,
    new_n17724_, new_n17725_, new_n17726_, new_n17727_, new_n17728_,
    new_n17729_, new_n17730_, new_n17731_, new_n17732_, new_n17733_,
    new_n17734_, new_n17735_, new_n17736_, new_n17737_, new_n17738_,
    new_n17739_, new_n17740_, new_n17741_, new_n17742_, new_n17743_,
    new_n17744_, new_n17745_, new_n17746_, new_n17747_, new_n17748_,
    new_n17749_, new_n17750_, new_n17751_, new_n17752_, new_n17753_,
    new_n17754_, new_n17755_, new_n17756_, new_n17757_, new_n17758_,
    new_n17759_, new_n17760_, new_n17761_, new_n17762_, new_n17763_,
    new_n17764_, new_n17765_, new_n17766_, new_n17767_, new_n17768_,
    new_n17769_, new_n17770_, new_n17771_, new_n17772_, new_n17773_,
    new_n17774_, new_n17775_, new_n17776_, new_n17777_, new_n17778_,
    new_n17779_, new_n17780_, new_n17781_, new_n17782_, new_n17783_,
    new_n17784_, new_n17785_, new_n17786_, new_n17787_, new_n17788_,
    new_n17789_, new_n17790_, new_n17791_, new_n17792_, new_n17793_,
    new_n17794_, new_n17795_, new_n17796_, new_n17797_, new_n17798_,
    new_n17799_, new_n17800_, new_n17801_, new_n17802_, new_n17803_,
    new_n17804_, new_n17805_, new_n17806_, new_n17807_, new_n17808_,
    new_n17809_, new_n17810_, new_n17811_, new_n17812_, new_n17813_,
    new_n17814_, new_n17815_, new_n17816_, new_n17817_, new_n17818_,
    new_n17819_, new_n17820_, new_n17821_, new_n17822_, new_n17823_,
    new_n17824_, new_n17825_, new_n17826_, new_n17827_, new_n17828_,
    new_n17829_, new_n17830_, new_n17831_, new_n17832_, new_n17833_,
    new_n17834_, new_n17835_, new_n17836_, new_n17837_, new_n17838_,
    new_n17839_, new_n17840_, new_n17841_, new_n17842_, new_n17843_,
    new_n17844_, new_n17845_, new_n17846_, new_n17847_, new_n17848_,
    new_n17849_, new_n17850_, new_n17851_, new_n17852_, new_n17854_,
    new_n17855_, new_n17856_, new_n17857_, new_n17858_, new_n17859_,
    new_n17860_, new_n17861_, new_n17862_, new_n17863_, new_n17864_,
    new_n17865_, new_n17866_, new_n17867_, new_n17868_, new_n17869_,
    new_n17870_, new_n17871_, new_n17872_, new_n17873_, new_n17874_,
    new_n17875_, new_n17876_, new_n17877_, new_n17878_, new_n17879_,
    new_n17880_, new_n17881_, new_n17882_, new_n17883_, new_n17884_,
    new_n17885_, new_n17886_, new_n17887_, new_n17888_, new_n17889_,
    new_n17890_, new_n17891_, new_n17892_, new_n17893_, new_n17894_,
    new_n17895_, new_n17896_, new_n17897_, new_n17898_, new_n17899_,
    new_n17900_, new_n17901_, new_n17902_, new_n17903_, new_n17904_,
    new_n17905_, new_n17906_, new_n17907_, new_n17908_, new_n17909_,
    new_n17910_, new_n17911_, new_n17912_, new_n17913_, new_n17914_,
    new_n17915_, new_n17916_, new_n17917_, new_n17918_, new_n17919_,
    new_n17920_, new_n17921_, new_n17922_, new_n17923_, new_n17924_,
    new_n17925_, new_n17926_, new_n17927_, new_n17928_, new_n17929_,
    new_n17930_, new_n17931_, new_n17932_, new_n17933_, new_n17934_,
    new_n17935_, new_n17936_, new_n17937_, new_n17938_, new_n17939_,
    new_n17940_, new_n17941_, new_n17942_, new_n17943_, new_n17944_,
    new_n17945_, new_n17946_, new_n17947_, new_n17948_, new_n17949_,
    new_n17950_, new_n17951_, new_n17952_, new_n17953_, new_n17954_,
    new_n17955_, new_n17956_, new_n17957_, new_n17958_, new_n17959_,
    new_n17960_, new_n17961_, new_n17962_, new_n17963_, new_n17964_,
    new_n17965_, new_n17966_, new_n17967_, new_n17968_, new_n17969_,
    new_n17970_, new_n17971_, new_n17972_, new_n17973_, new_n17974_,
    new_n17975_, new_n17976_, new_n17977_, new_n17978_, new_n17979_,
    new_n17980_, new_n17981_, new_n17982_, new_n17983_, new_n17984_,
    new_n17985_, new_n17986_, new_n17987_, new_n17988_, new_n17989_,
    new_n17990_, new_n17991_, new_n17992_, new_n17993_, new_n17994_,
    new_n17995_, new_n17996_, new_n17997_, new_n17998_, new_n17999_,
    new_n18000_, new_n18001_, new_n18002_, new_n18003_, new_n18004_,
    new_n18005_, new_n18006_, new_n18007_, new_n18008_, new_n18009_,
    new_n18010_, new_n18011_, new_n18012_, new_n18013_, new_n18014_,
    new_n18015_, new_n18016_, new_n18017_, new_n18018_, new_n18019_,
    new_n18020_, new_n18021_, new_n18022_, new_n18023_, new_n18024_,
    new_n18025_, new_n18026_, new_n18027_, new_n18028_, new_n18029_,
    new_n18030_, new_n18031_, new_n18032_, new_n18033_, new_n18034_,
    new_n18035_, new_n18036_, new_n18037_, new_n18038_, new_n18039_,
    new_n18040_, new_n18041_, new_n18042_, new_n18043_, new_n18044_,
    new_n18045_, new_n18046_, new_n18047_, new_n18048_, new_n18049_,
    new_n18050_, new_n18051_, new_n18052_, new_n18053_, new_n18054_,
    new_n18055_, new_n18056_, new_n18057_, new_n18058_, new_n18059_,
    new_n18060_, new_n18061_, new_n18062_, new_n18063_, new_n18064_,
    new_n18065_, new_n18066_, new_n18067_, new_n18068_, new_n18069_,
    new_n18070_, new_n18071_, new_n18072_, new_n18073_, new_n18074_,
    new_n18075_, new_n18076_, new_n18077_, new_n18078_, new_n18079_,
    new_n18080_, new_n18081_, new_n18082_, new_n18083_, new_n18084_,
    new_n18085_, new_n18086_, new_n18087_, new_n18088_, new_n18089_,
    new_n18090_, new_n18091_, new_n18092_, new_n18093_, new_n18094_,
    new_n18095_, new_n18096_, new_n18097_, new_n18098_, new_n18099_,
    new_n18100_, new_n18101_, new_n18102_, new_n18103_, new_n18104_,
    new_n18105_, new_n18106_, new_n18107_, new_n18108_, new_n18109_,
    new_n18110_, new_n18111_, new_n18112_, new_n18113_, new_n18114_,
    new_n18115_, new_n18116_, new_n18117_, new_n18118_, new_n18119_,
    new_n18120_, new_n18121_, new_n18122_, new_n18123_, new_n18124_,
    new_n18125_, new_n18126_, new_n18127_, new_n18128_, new_n18129_,
    new_n18130_, new_n18131_, new_n18132_, new_n18133_, new_n18134_,
    new_n18135_, new_n18136_, new_n18137_, new_n18138_, new_n18139_,
    new_n18140_, new_n18141_, new_n18142_, new_n18143_, new_n18144_,
    new_n18145_, new_n18146_, new_n18147_, new_n18148_, new_n18149_,
    new_n18150_, new_n18151_, new_n18152_, new_n18153_, new_n18154_,
    new_n18155_, new_n18156_, new_n18157_, new_n18158_, new_n18159_,
    new_n18160_, new_n18161_, new_n18162_, new_n18163_, new_n18164_,
    new_n18165_, new_n18166_, new_n18167_, new_n18168_, new_n18169_,
    new_n18170_, new_n18171_, new_n18172_, new_n18173_, new_n18174_,
    new_n18175_, new_n18176_, new_n18177_, new_n18178_, new_n18179_,
    new_n18180_, new_n18181_, new_n18182_, new_n18183_, new_n18184_,
    new_n18185_, new_n18186_, new_n18187_, new_n18188_, new_n18189_,
    new_n18190_, new_n18191_, new_n18192_, new_n18193_, new_n18194_,
    new_n18195_, new_n18196_, new_n18197_, new_n18198_, new_n18199_,
    new_n18200_, new_n18201_, new_n18202_, new_n18203_, new_n18204_,
    new_n18205_, new_n18206_, new_n18207_, new_n18208_, new_n18209_,
    new_n18210_, new_n18211_, new_n18212_, new_n18213_, new_n18214_,
    new_n18215_, new_n18216_, new_n18217_, new_n18218_, new_n18219_,
    new_n18220_, new_n18221_, new_n18222_, new_n18223_, new_n18224_,
    new_n18225_, new_n18226_, new_n18227_, new_n18228_, new_n18229_,
    new_n18230_, new_n18231_, new_n18232_, new_n18233_, new_n18234_,
    new_n18235_, new_n18236_, new_n18237_, new_n18238_, new_n18239_,
    new_n18240_, new_n18241_, new_n18242_, new_n18243_, new_n18244_,
    new_n18245_, new_n18246_, new_n18247_, new_n18248_, new_n18249_,
    new_n18250_, new_n18251_, new_n18252_, new_n18253_, new_n18254_,
    new_n18255_, new_n18256_, new_n18257_, new_n18258_, new_n18259_,
    new_n18260_, new_n18261_, new_n18262_, new_n18263_, new_n18264_,
    new_n18265_, new_n18266_, new_n18267_, new_n18268_, new_n18269_,
    new_n18270_, new_n18271_, new_n18272_, new_n18273_, new_n18274_,
    new_n18275_, new_n18276_, new_n18277_, new_n18278_, new_n18279_,
    new_n18280_, new_n18281_, new_n18282_, new_n18283_, new_n18284_,
    new_n18285_, new_n18286_, new_n18287_, new_n18288_, new_n18289_,
    new_n18290_, new_n18291_, new_n18292_, new_n18293_, new_n18294_,
    new_n18295_, new_n18296_, new_n18297_, new_n18298_, new_n18299_,
    new_n18300_, new_n18301_, new_n18302_, new_n18303_, new_n18304_,
    new_n18305_, new_n18306_, new_n18307_, new_n18308_, new_n18309_,
    new_n18310_, new_n18311_, new_n18312_, new_n18313_, new_n18314_,
    new_n18315_, new_n18316_, new_n18317_, new_n18318_, new_n18319_,
    new_n18320_, new_n18321_, new_n18322_, new_n18323_, new_n18324_,
    new_n18325_, new_n18326_, new_n18327_, new_n18328_, new_n18329_,
    new_n18330_, new_n18331_, new_n18332_, new_n18333_, new_n18334_,
    new_n18335_, new_n18336_, new_n18337_, new_n18338_, new_n18339_,
    new_n18340_, new_n18341_, new_n18342_, new_n18343_, new_n18344_,
    new_n18345_, new_n18346_, new_n18347_, new_n18348_, new_n18349_,
    new_n18350_, new_n18351_, new_n18352_, new_n18353_, new_n18354_,
    new_n18355_, new_n18356_, new_n18357_, new_n18358_, new_n18359_,
    new_n18360_, new_n18361_, new_n18362_, new_n18363_, new_n18364_,
    new_n18365_, new_n18366_, new_n18367_, new_n18368_, new_n18369_,
    new_n18370_, new_n18371_, new_n18372_, new_n18373_, new_n18374_,
    new_n18375_, new_n18376_, new_n18377_, new_n18378_, new_n18379_,
    new_n18380_, new_n18381_, new_n18382_, new_n18383_, new_n18384_,
    new_n18385_, new_n18386_, new_n18387_, new_n18388_, new_n18389_,
    new_n18390_, new_n18391_, new_n18392_, new_n18393_, new_n18394_,
    new_n18395_, new_n18396_, new_n18397_, new_n18398_, new_n18399_,
    new_n18400_, new_n18401_, new_n18402_, new_n18403_, new_n18404_,
    new_n18405_, new_n18406_, new_n18407_, new_n18408_, new_n18409_,
    new_n18410_, new_n18411_, new_n18412_, new_n18413_, new_n18414_,
    new_n18415_, new_n18416_, new_n18417_, new_n18418_, new_n18419_,
    new_n18420_, new_n18421_, new_n18422_, new_n18423_, new_n18424_,
    new_n18425_, new_n18426_, new_n18427_, new_n18428_, new_n18429_,
    new_n18430_, new_n18431_, new_n18432_, new_n18433_, new_n18434_,
    new_n18435_, new_n18436_, new_n18437_, new_n18438_, new_n18439_,
    new_n18440_, new_n18441_, new_n18442_, new_n18443_, new_n18444_,
    new_n18445_, new_n18446_, new_n18447_, new_n18448_, new_n18449_,
    new_n18450_, new_n18451_, new_n18452_, new_n18453_, new_n18454_,
    new_n18455_, new_n18456_, new_n18457_, new_n18458_, new_n18459_,
    new_n18460_, new_n18461_, new_n18462_, new_n18463_, new_n18464_,
    new_n18465_, new_n18466_, new_n18467_, new_n18468_, new_n18469_,
    new_n18470_, new_n18471_, new_n18472_, new_n18473_, new_n18474_,
    new_n18475_, new_n18476_, new_n18477_, new_n18478_, new_n18479_,
    new_n18480_, new_n18481_, new_n18482_, new_n18483_, new_n18484_,
    new_n18485_, new_n18486_, new_n18487_, new_n18488_, new_n18489_,
    new_n18490_, new_n18491_, new_n18492_, new_n18493_, new_n18494_,
    new_n18495_, new_n18496_, new_n18497_, new_n18498_, new_n18499_,
    new_n18500_, new_n18501_, new_n18502_, new_n18503_, new_n18504_,
    new_n18505_, new_n18507_, new_n18508_, new_n18509_, new_n18510_,
    new_n18511_, new_n18512_, new_n18513_, new_n18514_, new_n18515_,
    new_n18516_, new_n18517_, new_n18518_, new_n18519_, new_n18520_,
    new_n18521_, new_n18522_, new_n18523_, new_n18524_, new_n18525_,
    new_n18526_, new_n18527_, new_n18528_, new_n18529_, new_n18530_,
    new_n18531_, new_n18532_, new_n18533_, new_n18534_, new_n18535_,
    new_n18536_, new_n18537_, new_n18538_, new_n18539_, new_n18540_,
    new_n18541_, new_n18542_, new_n18543_, new_n18544_, new_n18545_,
    new_n18546_, new_n18547_, new_n18548_, new_n18549_, new_n18550_,
    new_n18551_, new_n18552_, new_n18553_, new_n18554_, new_n18555_,
    new_n18556_, new_n18557_, new_n18558_, new_n18559_, new_n18560_,
    new_n18561_, new_n18562_, new_n18563_, new_n18564_, new_n18565_,
    new_n18566_, new_n18567_, new_n18568_, new_n18569_, new_n18570_,
    new_n18571_, new_n18572_, new_n18573_, new_n18574_, new_n18575_,
    new_n18576_, new_n18577_, new_n18578_, new_n18579_, new_n18580_,
    new_n18581_, new_n18582_, new_n18583_, new_n18584_, new_n18585_,
    new_n18586_, new_n18587_, new_n18588_, new_n18589_, new_n18590_,
    new_n18591_, new_n18592_, new_n18593_, new_n18594_, new_n18595_,
    new_n18596_, new_n18597_, new_n18598_, new_n18599_, new_n18600_,
    new_n18601_, new_n18602_, new_n18603_, new_n18604_, new_n18605_,
    new_n18606_, new_n18607_, new_n18608_, new_n18609_, new_n18610_,
    new_n18611_, new_n18612_, new_n18613_, new_n18614_, new_n18615_,
    new_n18616_, new_n18617_, new_n18618_, new_n18619_, new_n18620_,
    new_n18621_, new_n18622_, new_n18623_, new_n18624_, new_n18625_,
    new_n18626_, new_n18627_, new_n18628_, new_n18629_, new_n18630_,
    new_n18631_, new_n18632_, new_n18633_, new_n18634_, new_n18635_,
    new_n18636_, new_n18637_, new_n18638_, new_n18639_, new_n18640_,
    new_n18641_, new_n18642_, new_n18643_, new_n18644_, new_n18645_,
    new_n18646_, new_n18647_, new_n18648_, new_n18649_, new_n18650_,
    new_n18651_, new_n18652_, new_n18653_, new_n18654_, new_n18655_,
    new_n18656_, new_n18657_, new_n18658_, new_n18659_, new_n18660_,
    new_n18661_, new_n18662_, new_n18663_, new_n18664_, new_n18665_,
    new_n18666_, new_n18667_, new_n18668_, new_n18669_, new_n18670_,
    new_n18671_, new_n18672_, new_n18673_, new_n18674_, new_n18675_,
    new_n18676_, new_n18677_, new_n18678_, new_n18679_, new_n18680_,
    new_n18681_, new_n18682_, new_n18683_, new_n18684_, new_n18685_,
    new_n18686_, new_n18687_, new_n18688_, new_n18689_, new_n18690_,
    new_n18691_, new_n18692_, new_n18693_, new_n18694_, new_n18695_,
    new_n18696_, new_n18697_, new_n18698_, new_n18699_, new_n18700_,
    new_n18701_, new_n18702_, new_n18703_, new_n18704_, new_n18705_,
    new_n18706_, new_n18707_, new_n18708_, new_n18709_, new_n18710_,
    new_n18711_, new_n18712_, new_n18713_, new_n18714_, new_n18715_,
    new_n18716_, new_n18717_, new_n18718_, new_n18719_, new_n18720_,
    new_n18721_, new_n18722_, new_n18723_, new_n18724_, new_n18725_,
    new_n18726_, new_n18727_, new_n18728_, new_n18729_, new_n18730_,
    new_n18731_, new_n18732_, new_n18733_, new_n18734_, new_n18735_,
    new_n18736_, new_n18737_, new_n18738_, new_n18739_, new_n18740_,
    new_n18741_, new_n18742_, new_n18743_, new_n18744_, new_n18745_,
    new_n18746_, new_n18747_, new_n18748_, new_n18749_, new_n18750_,
    new_n18751_, new_n18752_, new_n18753_, new_n18754_, new_n18755_,
    new_n18756_, new_n18757_, new_n18758_, new_n18759_, new_n18760_,
    new_n18761_, new_n18762_, new_n18763_, new_n18764_, new_n18765_,
    new_n18766_, new_n18767_, new_n18768_, new_n18769_, new_n18770_,
    new_n18771_, new_n18772_, new_n18773_, new_n18774_, new_n18775_,
    new_n18776_, new_n18777_, new_n18778_, new_n18779_, new_n18780_,
    new_n18781_, new_n18782_, new_n18783_, new_n18784_, new_n18785_,
    new_n18786_, new_n18787_, new_n18788_, new_n18789_, new_n18790_,
    new_n18791_, new_n18792_, new_n18793_, new_n18794_, new_n18795_,
    new_n18796_, new_n18797_, new_n18798_, new_n18799_, new_n18800_,
    new_n18801_, new_n18802_, new_n18803_, new_n18804_, new_n18805_,
    new_n18806_, new_n18807_, new_n18808_, new_n18809_, new_n18810_,
    new_n18811_, new_n18812_, new_n18813_, new_n18814_, new_n18815_,
    new_n18816_, new_n18817_, new_n18818_, new_n18819_, new_n18820_,
    new_n18821_, new_n18822_, new_n18823_, new_n18824_, new_n18825_,
    new_n18826_, new_n18827_, new_n18828_, new_n18829_, new_n18830_,
    new_n18831_, new_n18832_, new_n18833_, new_n18834_, new_n18835_,
    new_n18836_, new_n18837_, new_n18838_, new_n18839_, new_n18840_,
    new_n18841_, new_n18842_, new_n18843_, new_n18844_, new_n18845_,
    new_n18846_, new_n18847_, new_n18848_, new_n18849_, new_n18850_,
    new_n18851_, new_n18852_, new_n18853_, new_n18854_, new_n18855_,
    new_n18856_, new_n18857_, new_n18858_, new_n18859_, new_n18860_,
    new_n18861_, new_n18862_, new_n18863_, new_n18864_, new_n18865_,
    new_n18866_, new_n18867_, new_n18868_, new_n18869_, new_n18870_,
    new_n18871_, new_n18872_, new_n18873_, new_n18874_, new_n18875_,
    new_n18876_, new_n18877_, new_n18878_, new_n18879_, new_n18880_,
    new_n18881_, new_n18882_, new_n18883_, new_n18884_, new_n18885_,
    new_n18886_, new_n18887_, new_n18888_, new_n18889_, new_n18890_,
    new_n18891_, new_n18892_, new_n18893_, new_n18894_, new_n18895_,
    new_n18896_, new_n18897_, new_n18898_, new_n18899_, new_n18900_,
    new_n18901_, new_n18902_, new_n18903_, new_n18904_, new_n18905_,
    new_n18906_, new_n18907_, new_n18908_, new_n18909_, new_n18910_,
    new_n18911_, new_n18912_, new_n18913_, new_n18914_, new_n18915_,
    new_n18916_, new_n18917_, new_n18918_, new_n18919_, new_n18920_,
    new_n18921_, new_n18922_, new_n18923_, new_n18924_, new_n18925_,
    new_n18926_, new_n18927_, new_n18928_, new_n18929_, new_n18930_,
    new_n18931_, new_n18932_, new_n18933_, new_n18934_, new_n18935_,
    new_n18936_, new_n18937_, new_n18938_, new_n18939_, new_n18940_,
    new_n18941_, new_n18942_, new_n18943_, new_n18944_, new_n18945_,
    new_n18946_, new_n18947_, new_n18948_, new_n18949_, new_n18950_,
    new_n18951_, new_n18952_, new_n18953_, new_n18954_, new_n18955_,
    new_n18956_, new_n18957_, new_n18958_, new_n18959_, new_n18960_,
    new_n18961_, new_n18962_, new_n18963_, new_n18964_, new_n18965_,
    new_n18966_, new_n18967_, new_n18968_, new_n18969_, new_n18970_,
    new_n18971_, new_n18972_, new_n18973_, new_n18974_, new_n18975_,
    new_n18976_, new_n18977_, new_n18978_, new_n18979_, new_n18980_,
    new_n18981_, new_n18982_, new_n18983_, new_n18984_, new_n18985_,
    new_n18986_, new_n18987_, new_n18988_, new_n18989_, new_n18990_,
    new_n18991_, new_n18992_, new_n18993_, new_n18994_, new_n18995_,
    new_n18996_, new_n18997_, new_n18998_, new_n18999_, new_n19000_,
    new_n19001_, new_n19002_, new_n19003_, new_n19004_, new_n19005_,
    new_n19006_, new_n19007_, new_n19008_, new_n19009_, new_n19010_,
    new_n19011_, new_n19012_, new_n19013_, new_n19014_, new_n19015_,
    new_n19016_, new_n19017_, new_n19018_, new_n19019_, new_n19020_,
    new_n19021_, new_n19022_, new_n19023_, new_n19024_, new_n19025_,
    new_n19026_, new_n19027_, new_n19028_, new_n19029_, new_n19030_,
    new_n19031_, new_n19032_, new_n19033_, new_n19034_, new_n19035_,
    new_n19036_, new_n19037_, new_n19038_, new_n19039_, new_n19040_,
    new_n19041_, new_n19042_, new_n19043_, new_n19044_, new_n19045_,
    new_n19046_, new_n19047_, new_n19048_, new_n19049_, new_n19050_,
    new_n19051_, new_n19052_, new_n19053_, new_n19054_, new_n19055_,
    new_n19056_, new_n19057_, new_n19058_, new_n19059_, new_n19060_,
    new_n19061_, new_n19062_, new_n19063_, new_n19064_, new_n19065_,
    new_n19066_, new_n19067_, new_n19068_, new_n19069_, new_n19070_,
    new_n19071_, new_n19072_, new_n19073_, new_n19074_, new_n19075_,
    new_n19076_, new_n19077_, new_n19078_, new_n19079_, new_n19080_,
    new_n19081_, new_n19082_, new_n19083_, new_n19084_, new_n19085_,
    new_n19086_, new_n19087_, new_n19088_, new_n19089_, new_n19090_,
    new_n19091_, new_n19092_, new_n19093_, new_n19094_, new_n19095_,
    new_n19096_, new_n19097_, new_n19098_, new_n19099_, new_n19100_,
    new_n19101_, new_n19102_, new_n19103_, new_n19104_, new_n19105_,
    new_n19106_, new_n19107_, new_n19108_, new_n19109_, new_n19110_,
    new_n19111_, new_n19113_, new_n19114_, new_n19115_, new_n19116_,
    new_n19117_, new_n19118_, new_n19119_, new_n19120_, new_n19121_,
    new_n19122_, new_n19123_, new_n19124_, new_n19125_, new_n19126_,
    new_n19127_, new_n19128_, new_n19129_, new_n19130_, new_n19131_,
    new_n19132_, new_n19133_, new_n19134_, new_n19135_, new_n19136_,
    new_n19137_, new_n19138_, new_n19139_, new_n19140_, new_n19141_,
    new_n19142_, new_n19143_, new_n19144_, new_n19145_, new_n19146_,
    new_n19147_, new_n19148_, new_n19149_, new_n19150_, new_n19151_,
    new_n19152_, new_n19153_, new_n19154_, new_n19155_, new_n19156_,
    new_n19157_, new_n19158_, new_n19159_, new_n19160_, new_n19161_,
    new_n19162_, new_n19163_, new_n19164_, new_n19165_, new_n19166_,
    new_n19167_, new_n19168_, new_n19169_, new_n19170_, new_n19171_,
    new_n19172_, new_n19173_, new_n19174_, new_n19175_, new_n19176_,
    new_n19177_, new_n19178_, new_n19179_, new_n19180_, new_n19181_,
    new_n19182_, new_n19183_, new_n19184_, new_n19185_, new_n19186_,
    new_n19187_, new_n19188_, new_n19189_, new_n19190_, new_n19191_,
    new_n19192_, new_n19193_, new_n19194_, new_n19195_, new_n19196_,
    new_n19197_, new_n19198_, new_n19199_, new_n19200_, new_n19201_,
    new_n19202_, new_n19203_, new_n19204_, new_n19205_, new_n19206_,
    new_n19207_, new_n19208_, new_n19209_, new_n19210_, new_n19211_,
    new_n19212_, new_n19213_, new_n19214_, new_n19215_, new_n19216_,
    new_n19217_, new_n19218_, new_n19219_, new_n19220_, new_n19221_,
    new_n19222_, new_n19223_, new_n19224_, new_n19225_, new_n19226_,
    new_n19227_, new_n19228_, new_n19229_, new_n19230_, new_n19231_,
    new_n19232_, new_n19233_, new_n19234_, new_n19235_, new_n19236_,
    new_n19237_, new_n19238_, new_n19239_, new_n19240_, new_n19241_,
    new_n19242_, new_n19243_, new_n19244_, new_n19245_, new_n19246_,
    new_n19247_, new_n19248_, new_n19249_, new_n19250_, new_n19251_,
    new_n19252_, new_n19253_, new_n19254_, new_n19255_, new_n19256_,
    new_n19257_, new_n19258_, new_n19259_, new_n19260_, new_n19261_,
    new_n19262_, new_n19263_, new_n19264_, new_n19265_, new_n19266_,
    new_n19267_, new_n19268_, new_n19269_, new_n19270_, new_n19271_,
    new_n19272_, new_n19273_, new_n19274_, new_n19275_, new_n19276_,
    new_n19277_, new_n19278_, new_n19279_, new_n19280_, new_n19281_,
    new_n19282_, new_n19283_, new_n19284_, new_n19285_, new_n19286_,
    new_n19287_, new_n19288_, new_n19289_, new_n19290_, new_n19291_,
    new_n19292_, new_n19293_, new_n19294_, new_n19295_, new_n19296_,
    new_n19297_, new_n19298_, new_n19299_, new_n19300_, new_n19301_,
    new_n19302_, new_n19303_, new_n19304_, new_n19305_, new_n19306_,
    new_n19307_, new_n19308_, new_n19309_, new_n19310_, new_n19311_,
    new_n19312_, new_n19313_, new_n19314_, new_n19315_, new_n19316_,
    new_n19317_, new_n19318_, new_n19319_, new_n19320_, new_n19321_,
    new_n19322_, new_n19323_, new_n19324_, new_n19325_, new_n19326_,
    new_n19327_, new_n19328_, new_n19329_, new_n19330_, new_n19331_,
    new_n19332_, new_n19333_, new_n19334_, new_n19335_, new_n19336_,
    new_n19337_, new_n19338_, new_n19339_, new_n19340_, new_n19341_,
    new_n19342_, new_n19343_, new_n19344_, new_n19345_, new_n19346_,
    new_n19347_, new_n19348_, new_n19349_, new_n19350_, new_n19351_,
    new_n19352_, new_n19353_, new_n19354_, new_n19355_, new_n19356_,
    new_n19357_, new_n19358_, new_n19359_, new_n19360_, new_n19361_,
    new_n19362_, new_n19363_, new_n19364_, new_n19365_, new_n19366_,
    new_n19367_, new_n19368_, new_n19369_, new_n19370_, new_n19371_,
    new_n19372_, new_n19373_, new_n19374_, new_n19375_, new_n19376_,
    new_n19377_, new_n19378_, new_n19379_, new_n19380_, new_n19381_,
    new_n19382_, new_n19383_, new_n19384_, new_n19385_, new_n19386_,
    new_n19387_, new_n19388_, new_n19389_, new_n19390_, new_n19391_,
    new_n19392_, new_n19393_, new_n19394_, new_n19395_, new_n19396_,
    new_n19397_, new_n19398_, new_n19399_, new_n19400_, new_n19401_,
    new_n19402_, new_n19403_, new_n19404_, new_n19405_, new_n19406_,
    new_n19407_, new_n19408_, new_n19409_, new_n19410_, new_n19411_,
    new_n19412_, new_n19413_, new_n19414_, new_n19415_, new_n19416_,
    new_n19417_, new_n19418_, new_n19419_, new_n19420_, new_n19421_,
    new_n19422_, new_n19423_, new_n19424_, new_n19425_, new_n19426_,
    new_n19427_, new_n19428_, new_n19429_, new_n19430_, new_n19431_,
    new_n19432_, new_n19433_, new_n19434_, new_n19435_, new_n19436_,
    new_n19437_, new_n19438_, new_n19439_, new_n19440_, new_n19441_,
    new_n19442_, new_n19443_, new_n19444_, new_n19445_, new_n19446_,
    new_n19447_, new_n19448_, new_n19449_, new_n19450_, new_n19451_,
    new_n19452_, new_n19453_, new_n19454_, new_n19455_, new_n19456_,
    new_n19457_, new_n19458_, new_n19459_, new_n19460_, new_n19461_,
    new_n19462_, new_n19463_, new_n19464_, new_n19465_, new_n19466_,
    new_n19467_, new_n19468_, new_n19469_, new_n19470_, new_n19471_,
    new_n19472_, new_n19473_, new_n19474_, new_n19475_, new_n19476_,
    new_n19477_, new_n19478_, new_n19479_, new_n19480_, new_n19481_,
    new_n19482_, new_n19483_, new_n19484_, new_n19485_, new_n19486_,
    new_n19487_, new_n19488_, new_n19489_, new_n19490_, new_n19491_,
    new_n19492_, new_n19493_, new_n19494_, new_n19495_, new_n19496_,
    new_n19497_, new_n19498_, new_n19499_, new_n19500_, new_n19501_,
    new_n19502_, new_n19503_, new_n19504_, new_n19505_, new_n19506_,
    new_n19507_, new_n19508_, new_n19509_, new_n19510_, new_n19511_,
    new_n19512_, new_n19513_, new_n19514_, new_n19515_, new_n19516_,
    new_n19517_, new_n19518_, new_n19519_, new_n19520_, new_n19521_,
    new_n19522_, new_n19523_, new_n19524_, new_n19525_, new_n19526_,
    new_n19527_, new_n19528_, new_n19529_, new_n19530_, new_n19531_,
    new_n19532_, new_n19533_, new_n19534_, new_n19535_, new_n19536_,
    new_n19537_, new_n19538_, new_n19539_, new_n19540_, new_n19541_,
    new_n19542_, new_n19543_, new_n19544_, new_n19545_, new_n19546_,
    new_n19547_, new_n19548_, new_n19549_, new_n19550_, new_n19551_,
    new_n19552_, new_n19553_, new_n19554_, new_n19555_, new_n19556_,
    new_n19557_, new_n19558_, new_n19559_, new_n19560_, new_n19561_,
    new_n19562_, new_n19563_, new_n19564_, new_n19565_, new_n19566_,
    new_n19567_, new_n19568_, new_n19569_, new_n19570_, new_n19571_,
    new_n19572_, new_n19573_, new_n19574_, new_n19575_, new_n19576_,
    new_n19577_, new_n19578_, new_n19579_, new_n19580_, new_n19581_,
    new_n19582_, new_n19583_, new_n19584_, new_n19585_, new_n19586_,
    new_n19587_, new_n19588_, new_n19589_, new_n19590_, new_n19591_,
    new_n19592_, new_n19593_, new_n19594_, new_n19595_, new_n19596_,
    new_n19597_, new_n19598_, new_n19599_, new_n19600_, new_n19601_,
    new_n19602_, new_n19603_, new_n19604_, new_n19605_, new_n19606_,
    new_n19607_, new_n19608_, new_n19609_, new_n19610_, new_n19611_,
    new_n19612_, new_n19613_, new_n19614_, new_n19615_, new_n19616_,
    new_n19617_, new_n19618_, new_n19619_, new_n19620_, new_n19621_,
    new_n19622_, new_n19623_, new_n19624_, new_n19625_, new_n19626_,
    new_n19627_, new_n19628_, new_n19629_, new_n19630_, new_n19631_,
    new_n19632_, new_n19633_, new_n19634_, new_n19635_, new_n19636_,
    new_n19637_, new_n19638_, new_n19639_, new_n19640_, new_n19641_,
    new_n19642_, new_n19643_, new_n19644_, new_n19645_, new_n19646_,
    new_n19647_, new_n19648_, new_n19649_, new_n19650_, new_n19651_,
    new_n19652_, new_n19653_, new_n19654_, new_n19655_, new_n19656_,
    new_n19657_, new_n19658_, new_n19659_, new_n19660_, new_n19661_,
    new_n19662_, new_n19663_, new_n19664_, new_n19665_, new_n19666_,
    new_n19667_, new_n19668_, new_n19669_, new_n19670_, new_n19671_,
    new_n19672_, new_n19673_, new_n19674_, new_n19675_, new_n19676_,
    new_n19677_, new_n19678_, new_n19679_, new_n19680_, new_n19681_,
    new_n19682_, new_n19683_, new_n19684_, new_n19685_, new_n19686_,
    new_n19687_, new_n19688_, new_n19689_, new_n19690_, new_n19691_,
    new_n19692_, new_n19693_, new_n19694_, new_n19695_, new_n19696_,
    new_n19697_, new_n19698_, new_n19699_, new_n19700_, new_n19701_,
    new_n19702_, new_n19703_, new_n19704_, new_n19705_, new_n19706_,
    new_n19707_, new_n19708_, new_n19709_, new_n19710_, new_n19711_,
    new_n19712_, new_n19713_, new_n19714_, new_n19715_, new_n19716_,
    new_n19717_, new_n19718_, new_n19719_, new_n19720_, new_n19721_,
    new_n19722_, new_n19723_, new_n19724_, new_n19725_, new_n19726_,
    new_n19727_, new_n19728_, new_n19729_, new_n19730_, new_n19731_,
    new_n19732_, new_n19733_, new_n19734_, new_n19735_, new_n19736_,
    new_n19737_, new_n19738_, new_n19739_, new_n19740_, new_n19741_,
    new_n19742_, new_n19743_, new_n19744_, new_n19745_, new_n19746_,
    new_n19747_, new_n19748_, new_n19749_, new_n19750_, new_n19751_,
    new_n19752_, new_n19753_, new_n19754_, new_n19755_, new_n19756_,
    new_n19757_, new_n19758_, new_n19759_, new_n19760_, new_n19761_,
    new_n19762_, new_n19763_, new_n19764_, new_n19765_, new_n19766_,
    new_n19767_, new_n19768_, new_n19769_, new_n19770_, new_n19771_,
    new_n19772_, new_n19773_, new_n19774_, new_n19775_, new_n19776_,
    new_n19777_, new_n19778_, new_n19779_, new_n19780_, new_n19781_,
    new_n19782_, new_n19783_, new_n19784_, new_n19786_, new_n19787_,
    new_n19788_, new_n19789_, new_n19790_, new_n19791_, new_n19792_,
    new_n19793_, new_n19794_, new_n19795_, new_n19796_, new_n19797_,
    new_n19798_, new_n19799_, new_n19800_, new_n19801_, new_n19802_,
    new_n19803_, new_n19804_, new_n19805_, new_n19806_, new_n19807_,
    new_n19808_, new_n19809_, new_n19810_, new_n19811_, new_n19812_,
    new_n19813_, new_n19814_, new_n19815_, new_n19816_, new_n19817_,
    new_n19818_, new_n19819_, new_n19820_, new_n19821_, new_n19822_,
    new_n19823_, new_n19824_, new_n19825_, new_n19826_, new_n19827_,
    new_n19828_, new_n19829_, new_n19830_, new_n19831_, new_n19832_,
    new_n19833_, new_n19834_, new_n19835_, new_n19836_, new_n19837_,
    new_n19838_, new_n19839_, new_n19840_, new_n19841_, new_n19842_,
    new_n19843_, new_n19844_, new_n19845_, new_n19846_, new_n19847_,
    new_n19848_, new_n19849_, new_n19850_, new_n19851_, new_n19852_,
    new_n19853_, new_n19854_, new_n19855_, new_n19856_, new_n19857_,
    new_n19858_, new_n19859_, new_n19860_, new_n19861_, new_n19862_,
    new_n19863_, new_n19864_, new_n19865_, new_n19866_, new_n19867_,
    new_n19868_, new_n19869_, new_n19870_, new_n19871_, new_n19872_,
    new_n19873_, new_n19874_, new_n19875_, new_n19876_, new_n19877_,
    new_n19878_, new_n19879_, new_n19880_, new_n19881_, new_n19882_,
    new_n19883_, new_n19884_, new_n19885_, new_n19886_, new_n19887_,
    new_n19888_, new_n19889_, new_n19890_, new_n19891_, new_n19892_,
    new_n19893_, new_n19894_, new_n19895_, new_n19896_, new_n19897_,
    new_n19898_, new_n19899_, new_n19900_, new_n19901_, new_n19902_,
    new_n19903_, new_n19904_, new_n19905_, new_n19906_, new_n19907_,
    new_n19908_, new_n19909_, new_n19910_, new_n19911_, new_n19912_,
    new_n19913_, new_n19914_, new_n19915_, new_n19916_, new_n19917_,
    new_n19918_, new_n19919_, new_n19920_, new_n19921_, new_n19922_,
    new_n19923_, new_n19924_, new_n19925_, new_n19926_, new_n19927_,
    new_n19928_, new_n19929_, new_n19930_, new_n19931_, new_n19932_,
    new_n19933_, new_n19934_, new_n19935_, new_n19936_, new_n19937_,
    new_n19938_, new_n19939_, new_n19940_, new_n19941_, new_n19942_,
    new_n19943_, new_n19944_, new_n19945_, new_n19946_, new_n19947_,
    new_n19948_, new_n19949_, new_n19950_, new_n19951_, new_n19952_,
    new_n19953_, new_n19954_, new_n19955_, new_n19956_, new_n19957_,
    new_n19958_, new_n19959_, new_n19960_, new_n19961_, new_n19962_,
    new_n19963_, new_n19964_, new_n19965_, new_n19966_, new_n19967_,
    new_n19968_, new_n19969_, new_n19970_, new_n19971_, new_n19972_,
    new_n19973_, new_n19974_, new_n19975_, new_n19976_, new_n19977_,
    new_n19978_, new_n19979_, new_n19980_, new_n19981_, new_n19982_,
    new_n19983_, new_n19984_, new_n19985_, new_n19986_, new_n19987_,
    new_n19988_, new_n19989_, new_n19990_, new_n19991_, new_n19992_,
    new_n19993_, new_n19994_, new_n19995_, new_n19996_, new_n19997_,
    new_n19998_, new_n19999_, new_n20000_, new_n20001_, new_n20002_,
    new_n20003_, new_n20004_, new_n20005_, new_n20006_, new_n20007_,
    new_n20008_, new_n20009_, new_n20010_, new_n20011_, new_n20012_,
    new_n20013_, new_n20014_, new_n20015_, new_n20016_, new_n20017_,
    new_n20018_, new_n20019_, new_n20020_, new_n20021_, new_n20022_,
    new_n20023_, new_n20024_, new_n20025_, new_n20026_, new_n20027_,
    new_n20028_, new_n20029_, new_n20030_, new_n20031_, new_n20032_,
    new_n20033_, new_n20034_, new_n20035_, new_n20036_, new_n20037_,
    new_n20038_, new_n20039_, new_n20040_, new_n20041_, new_n20042_,
    new_n20043_, new_n20044_, new_n20045_, new_n20046_, new_n20047_,
    new_n20048_, new_n20049_, new_n20050_, new_n20051_, new_n20052_,
    new_n20053_, new_n20054_, new_n20055_, new_n20056_, new_n20057_,
    new_n20058_, new_n20059_, new_n20060_, new_n20061_, new_n20062_,
    new_n20063_, new_n20064_, new_n20065_, new_n20066_, new_n20067_,
    new_n20068_, new_n20069_, new_n20070_, new_n20071_, new_n20072_,
    new_n20073_, new_n20074_, new_n20075_, new_n20076_, new_n20077_,
    new_n20078_, new_n20079_, new_n20080_, new_n20081_, new_n20082_,
    new_n20083_, new_n20084_, new_n20085_, new_n20086_, new_n20087_,
    new_n20088_, new_n20089_, new_n20090_, new_n20091_, new_n20092_,
    new_n20093_, new_n20094_, new_n20095_, new_n20096_, new_n20097_,
    new_n20098_, new_n20099_, new_n20100_, new_n20101_, new_n20102_,
    new_n20103_, new_n20104_, new_n20105_, new_n20106_, new_n20107_,
    new_n20108_, new_n20109_, new_n20110_, new_n20111_, new_n20112_,
    new_n20113_, new_n20114_, new_n20115_, new_n20116_, new_n20117_,
    new_n20118_, new_n20119_, new_n20120_, new_n20121_, new_n20122_,
    new_n20123_, new_n20124_, new_n20125_, new_n20126_, new_n20127_,
    new_n20128_, new_n20129_, new_n20130_, new_n20131_, new_n20132_,
    new_n20133_, new_n20134_, new_n20135_, new_n20136_, new_n20137_,
    new_n20138_, new_n20139_, new_n20140_, new_n20141_, new_n20142_,
    new_n20143_, new_n20144_, new_n20145_, new_n20146_, new_n20147_,
    new_n20148_, new_n20149_, new_n20150_, new_n20151_, new_n20152_,
    new_n20153_, new_n20154_, new_n20155_, new_n20156_, new_n20157_,
    new_n20158_, new_n20159_, new_n20160_, new_n20161_, new_n20162_,
    new_n20163_, new_n20164_, new_n20165_, new_n20166_, new_n20167_,
    new_n20168_, new_n20169_, new_n20170_, new_n20171_, new_n20172_,
    new_n20173_, new_n20174_, new_n20175_, new_n20176_, new_n20177_,
    new_n20178_, new_n20179_, new_n20180_, new_n20181_, new_n20182_,
    new_n20183_, new_n20184_, new_n20185_, new_n20186_, new_n20187_,
    new_n20188_, new_n20189_, new_n20190_, new_n20191_, new_n20192_,
    new_n20193_, new_n20194_, new_n20195_, new_n20196_, new_n20197_,
    new_n20198_, new_n20199_, new_n20200_, new_n20201_, new_n20202_,
    new_n20203_, new_n20204_, new_n20205_, new_n20206_, new_n20207_,
    new_n20208_, new_n20209_, new_n20210_, new_n20211_, new_n20212_,
    new_n20213_, new_n20214_, new_n20215_, new_n20216_, new_n20217_,
    new_n20218_, new_n20219_, new_n20220_, new_n20221_, new_n20222_,
    new_n20223_, new_n20224_, new_n20225_, new_n20226_, new_n20227_,
    new_n20228_, new_n20229_, new_n20230_, new_n20231_, new_n20232_,
    new_n20233_, new_n20234_, new_n20235_, new_n20236_, new_n20237_,
    new_n20238_, new_n20239_, new_n20240_, new_n20241_, new_n20242_,
    new_n20243_, new_n20244_, new_n20245_, new_n20246_, new_n20247_,
    new_n20248_, new_n20249_, new_n20250_, new_n20251_, new_n20252_,
    new_n20253_, new_n20254_, new_n20255_, new_n20256_, new_n20257_,
    new_n20258_, new_n20259_, new_n20260_, new_n20261_, new_n20262_,
    new_n20263_, new_n20264_, new_n20265_, new_n20266_, new_n20267_,
    new_n20268_, new_n20269_, new_n20270_, new_n20271_, new_n20272_,
    new_n20273_, new_n20274_, new_n20275_, new_n20276_, new_n20277_,
    new_n20278_, new_n20279_, new_n20280_, new_n20281_, new_n20282_,
    new_n20283_, new_n20284_, new_n20285_, new_n20286_, new_n20287_,
    new_n20288_, new_n20289_, new_n20290_, new_n20291_, new_n20292_,
    new_n20293_, new_n20294_, new_n20295_, new_n20296_, new_n20297_,
    new_n20298_, new_n20299_, new_n20300_, new_n20301_, new_n20302_,
    new_n20303_, new_n20304_, new_n20305_, new_n20306_, new_n20307_,
    new_n20308_, new_n20309_, new_n20310_, new_n20311_, new_n20312_,
    new_n20313_, new_n20314_, new_n20315_, new_n20316_, new_n20317_,
    new_n20318_, new_n20319_, new_n20320_, new_n20321_, new_n20322_,
    new_n20323_, new_n20324_, new_n20325_, new_n20326_, new_n20327_,
    new_n20328_, new_n20329_, new_n20330_, new_n20331_, new_n20332_,
    new_n20333_, new_n20334_, new_n20335_, new_n20336_, new_n20337_,
    new_n20338_, new_n20339_, new_n20340_, new_n20341_, new_n20342_,
    new_n20343_, new_n20344_, new_n20345_, new_n20346_, new_n20347_,
    new_n20348_, new_n20349_, new_n20350_, new_n20351_, new_n20352_,
    new_n20353_, new_n20354_, new_n20355_, new_n20356_, new_n20357_,
    new_n20358_, new_n20359_, new_n20360_, new_n20361_, new_n20362_,
    new_n20363_, new_n20364_, new_n20365_, new_n20366_, new_n20367_,
    new_n20368_, new_n20369_, new_n20370_, new_n20371_, new_n20372_,
    new_n20373_, new_n20374_, new_n20375_, new_n20376_, new_n20377_,
    new_n20378_, new_n20379_, new_n20380_, new_n20381_, new_n20382_,
    new_n20383_, new_n20384_, new_n20385_, new_n20386_, new_n20387_,
    new_n20388_, new_n20389_, new_n20390_, new_n20391_, new_n20392_,
    new_n20393_, new_n20394_, new_n20395_, new_n20396_, new_n20397_,
    new_n20398_, new_n20399_, new_n20400_, new_n20401_, new_n20402_,
    new_n20403_, new_n20404_, new_n20405_, new_n20406_, new_n20407_,
    new_n20408_, new_n20409_, new_n20410_, new_n20411_, new_n20412_,
    new_n20413_, new_n20414_, new_n20415_, new_n20416_, new_n20417_,
    new_n20418_, new_n20419_, new_n20420_, new_n20421_, new_n20422_,
    new_n20423_, new_n20424_, new_n20425_, new_n20426_, new_n20427_,
    new_n20428_, new_n20429_, new_n20430_, new_n20431_, new_n20432_,
    new_n20433_, new_n20434_, new_n20435_, new_n20436_, new_n20437_,
    new_n20438_, new_n20439_, new_n20441_, new_n20442_, new_n20443_,
    new_n20444_, new_n20446_, new_n20447_, new_n20448_, new_n20449_,
    new_n20450_, new_n20451_, new_n20452_, new_n20453_, new_n20454_,
    new_n20455_, new_n20456_, new_n20457_, new_n20458_, new_n20459_,
    new_n20460_, new_n20461_, new_n20462_, new_n20463_, new_n20464_,
    new_n20465_, new_n20466_, new_n20467_, new_n20468_, new_n20469_,
    new_n20470_, new_n20471_, new_n20472_, new_n20473_, new_n20474_,
    new_n20475_, new_n20476_, new_n20477_, new_n20478_, new_n20479_,
    new_n20480_, new_n20481_, new_n20482_, new_n20483_, new_n20484_,
    new_n20485_, new_n20486_, new_n20487_, new_n20488_, new_n20489_,
    new_n20490_, new_n20491_, new_n20492_, new_n20493_, new_n20494_,
    new_n20495_, new_n20496_, new_n20497_, new_n20498_, new_n20499_,
    new_n20500_, new_n20501_, new_n20502_, new_n20503_, new_n20504_,
    new_n20505_, new_n20506_, new_n20507_, new_n20508_, new_n20509_,
    new_n20510_, new_n20511_, new_n20512_, new_n20513_, new_n20514_,
    new_n20515_, new_n20516_, new_n20517_, new_n20518_, new_n20519_,
    new_n20520_, new_n20521_, new_n20522_, new_n20523_, new_n20524_,
    new_n20525_, new_n20526_, new_n20527_, new_n20528_, new_n20529_,
    new_n20530_, new_n20531_, new_n20532_, new_n20533_, new_n20534_,
    new_n20535_, new_n20536_, new_n20537_, new_n20538_, new_n20539_,
    new_n20540_, new_n20541_, new_n20542_, new_n20543_, new_n20544_,
    new_n20545_, new_n20546_, new_n20547_, new_n20548_, new_n20549_,
    new_n20550_, new_n20551_, new_n20552_, new_n20553_, new_n20554_,
    new_n20555_, new_n20556_, new_n20557_, new_n20558_, new_n20559_,
    new_n20560_, new_n20561_, new_n20562_, new_n20563_, new_n20564_,
    new_n20565_, new_n20566_, new_n20567_, new_n20568_, new_n20569_,
    new_n20570_, new_n20571_, new_n20572_, new_n20573_, new_n20574_,
    new_n20575_, new_n20576_, new_n20577_, new_n20578_, new_n20579_,
    new_n20580_, new_n20581_, new_n20582_, new_n20583_, new_n20584_,
    new_n20585_, new_n20586_, new_n20587_, new_n20588_, new_n20589_,
    new_n20590_, new_n20591_, new_n20592_, new_n20593_, new_n20594_,
    new_n20595_, new_n20596_, new_n20597_, new_n20598_, new_n20599_,
    new_n20600_, new_n20601_, new_n20602_, new_n20603_, new_n20604_,
    new_n20605_, new_n20606_, new_n20607_, new_n20608_, new_n20609_,
    new_n20610_, new_n20611_, new_n20612_, new_n20613_, new_n20614_,
    new_n20615_, new_n20616_, new_n20617_, new_n20618_, new_n20619_,
    new_n20620_, new_n20621_, new_n20622_, new_n20623_, new_n20624_,
    new_n20625_, new_n20626_, new_n20627_, new_n20628_, new_n20629_,
    new_n20630_, new_n20631_, new_n20632_, new_n20633_, new_n20634_,
    new_n20635_, new_n20636_, new_n20637_, new_n20638_, new_n20639_,
    new_n20640_, new_n20641_, new_n20642_, new_n20643_, new_n20644_,
    new_n20645_, new_n20646_, new_n20647_, new_n20648_, new_n20649_,
    new_n20650_, new_n20651_, new_n20652_, new_n20653_, new_n20654_,
    new_n20655_, new_n20656_, new_n20657_, new_n20658_, new_n20659_,
    new_n20660_, new_n20661_, new_n20662_, new_n20663_, new_n20664_,
    new_n20665_, new_n20666_, new_n20667_, new_n20668_, new_n20669_,
    new_n20670_, new_n20671_, new_n20672_, new_n20673_, new_n20674_,
    new_n20675_, new_n20676_, new_n20677_, new_n20678_, new_n20679_,
    new_n20680_, new_n20681_, new_n20682_, new_n20683_, new_n20684_,
    new_n20685_, new_n20686_, new_n20687_, new_n20688_, new_n20689_,
    new_n20690_, new_n20691_, new_n20692_, new_n20693_, new_n20694_,
    new_n20695_, new_n20696_, new_n20697_, new_n20698_, new_n20699_,
    new_n20700_, new_n20701_, new_n20702_, new_n20703_, new_n20704_,
    new_n20705_, new_n20706_, new_n20707_, new_n20708_, new_n20709_,
    new_n20710_, new_n20711_, new_n20712_, new_n20713_, new_n20714_,
    new_n20715_, new_n20716_, new_n20717_, new_n20718_, new_n20719_,
    new_n20720_, new_n20721_, new_n20722_, new_n20723_, new_n20724_,
    new_n20725_, new_n20726_, new_n20727_, new_n20728_, new_n20729_,
    new_n20730_, new_n20731_, new_n20732_, new_n20733_, new_n20734_,
    new_n20735_, new_n20736_, new_n20737_, new_n20738_, new_n20739_,
    new_n20740_, new_n20741_, new_n20742_, new_n20743_, new_n20744_,
    new_n20745_, new_n20746_, new_n20747_, new_n20748_, new_n20749_,
    new_n20750_, new_n20751_, new_n20752_, new_n20753_, new_n20754_,
    new_n20755_, new_n20756_, new_n20757_, new_n20758_, new_n20759_,
    new_n20760_, new_n20761_, new_n20762_, new_n20763_, new_n20764_,
    new_n20765_, new_n20766_, new_n20767_, new_n20768_, new_n20769_,
    new_n20770_, new_n20771_, new_n20772_, new_n20773_, new_n20774_,
    new_n20775_, new_n20776_, new_n20777_, new_n20778_, new_n20779_,
    new_n20780_, new_n20781_, new_n20782_, new_n20783_, new_n20784_,
    new_n20785_, new_n20786_, new_n20787_, new_n20788_, new_n20789_,
    new_n20790_, new_n20791_, new_n20792_, new_n20793_, new_n20794_,
    new_n20795_, new_n20796_, new_n20797_, new_n20798_, new_n20799_,
    new_n20800_, new_n20801_, new_n20802_, new_n20803_, new_n20804_,
    new_n20805_, new_n20806_, new_n20807_, new_n20808_, new_n20809_,
    new_n20810_, new_n20811_, new_n20812_, new_n20813_, new_n20814_,
    new_n20815_, new_n20816_, new_n20817_, new_n20818_, new_n20819_,
    new_n20820_, new_n20821_, new_n20822_, new_n20823_, new_n20824_,
    new_n20825_, new_n20826_, new_n20827_, new_n20828_, new_n20829_,
    new_n20830_, new_n20831_, new_n20832_, new_n20833_, new_n20834_,
    new_n20835_, new_n20836_, new_n20837_, new_n20838_, new_n20839_,
    new_n20840_, new_n20841_, new_n20842_, new_n20843_, new_n20844_,
    new_n20845_, new_n20846_, new_n20847_, new_n20848_, new_n20849_,
    new_n20850_, new_n20851_, new_n20852_, new_n20853_, new_n20854_,
    new_n20855_, new_n20856_, new_n20857_, new_n20858_, new_n20859_,
    new_n20860_, new_n20861_, new_n20862_, new_n20863_, new_n20864_,
    new_n20865_, new_n20866_, new_n20867_, new_n20868_, new_n20869_,
    new_n20870_, new_n20871_, new_n20872_, new_n20873_, new_n20874_,
    new_n20875_, new_n20876_, new_n20877_, new_n20878_, new_n20879_,
    new_n20880_, new_n20881_, new_n20882_, new_n20883_, new_n20884_,
    new_n20885_, new_n20886_, new_n20887_, new_n20888_, new_n20889_,
    new_n20890_, new_n20891_, new_n20892_, new_n20893_, new_n20894_,
    new_n20895_, new_n20896_, new_n20897_, new_n20898_, new_n20899_,
    new_n20900_, new_n20901_, new_n20902_, new_n20903_, new_n20904_,
    new_n20905_, new_n20906_, new_n20907_, new_n20908_, new_n20909_,
    new_n20910_, new_n20911_, new_n20912_, new_n20913_, new_n20914_,
    new_n20915_, new_n20916_, new_n20917_, new_n20918_, new_n20919_,
    new_n20920_, new_n20921_, new_n20922_, new_n20923_, new_n20924_,
    new_n20925_, new_n20926_, new_n20927_, new_n20928_, new_n20929_,
    new_n20930_, new_n20931_, new_n20932_, new_n20933_, new_n20934_,
    new_n20935_, new_n20936_, new_n20937_, new_n20938_, new_n20939_,
    new_n20940_, new_n20941_, new_n20942_, new_n20943_, new_n20944_,
    new_n20945_, new_n20946_, new_n20947_, new_n20948_, new_n20949_,
    new_n20950_, new_n20951_, new_n20952_, new_n20953_, new_n20954_,
    new_n20955_, new_n20956_, new_n20957_, new_n20958_, new_n20959_,
    new_n20960_, new_n20961_, new_n20962_, new_n20963_, new_n20964_,
    new_n20965_, new_n20966_, new_n20967_, new_n20968_, new_n20969_,
    new_n20970_, new_n20971_, new_n20972_, new_n20973_, new_n20974_,
    new_n20975_, new_n20976_, new_n20977_, new_n20978_, new_n20979_,
    new_n20980_, new_n20981_, new_n20982_, new_n20983_, new_n20984_,
    new_n20985_, new_n20986_, new_n20987_, new_n20988_, new_n20989_,
    new_n20990_, new_n20991_, new_n20992_, new_n20993_, new_n20994_,
    new_n20995_, new_n20996_, new_n20997_, new_n20998_, new_n20999_,
    new_n21000_, new_n21001_, new_n21002_, new_n21003_, new_n21004_,
    new_n21005_, new_n21006_, new_n21007_, new_n21008_, new_n21009_,
    new_n21010_, new_n21011_, new_n21012_, new_n21013_, new_n21014_,
    new_n21015_, new_n21016_, new_n21017_, new_n21018_, new_n21019_,
    new_n21020_, new_n21021_, new_n21022_, new_n21023_, new_n21024_,
    new_n21025_, new_n21026_, new_n21027_, new_n21028_, new_n21029_,
    new_n21030_, new_n21031_, new_n21032_, new_n21033_, new_n21034_,
    new_n21035_, new_n21036_, new_n21037_, new_n21038_, new_n21039_,
    new_n21040_, new_n21041_, new_n21042_, new_n21043_, new_n21044_,
    new_n21045_, new_n21046_, new_n21047_, new_n21048_, new_n21049_,
    new_n21050_, new_n21051_, new_n21052_, new_n21053_, new_n21054_,
    new_n21055_, new_n21056_, new_n21057_, new_n21058_, new_n21059_,
    new_n21060_, new_n21061_, new_n21062_, new_n21063_, new_n21064_,
    new_n21065_, new_n21066_, new_n21067_, new_n21068_, new_n21069_,
    new_n21070_, new_n21071_, new_n21072_, new_n21073_, new_n21074_,
    new_n21075_, new_n21076_, new_n21077_, new_n21078_, new_n21079_,
    new_n21080_, new_n21081_, new_n21082_, new_n21083_, new_n21084_,
    new_n21085_, new_n21086_, new_n21087_, new_n21088_, new_n21089_,
    new_n21090_, new_n21091_, new_n21092_, new_n21093_, new_n21094_,
    new_n21095_, new_n21096_, new_n21097_, new_n21098_, new_n21099_,
    new_n21100_, new_n21101_, new_n21102_, new_n21103_, new_n21104_,
    new_n21105_, new_n21106_, new_n21107_, new_n21108_, new_n21109_,
    new_n21110_, new_n21111_, new_n21112_, new_n21113_, new_n21114_,
    new_n21115_, new_n21116_, new_n21117_, new_n21118_, new_n21119_,
    new_n21120_, new_n21121_, new_n21122_, new_n21123_, new_n21124_,
    new_n21125_, new_n21126_, new_n21127_, new_n21129_, new_n21130_,
    new_n21131_, new_n21132_, new_n21133_, new_n21134_, new_n21135_,
    new_n21136_, new_n21137_, new_n21138_, new_n21139_, new_n21140_,
    new_n21141_, new_n21142_, new_n21143_, new_n21144_, new_n21145_,
    new_n21146_, new_n21147_, new_n21148_, new_n21149_, new_n21150_,
    new_n21151_, new_n21152_, new_n21153_, new_n21154_, new_n21155_,
    new_n21156_, new_n21157_, new_n21158_, new_n21159_, new_n21160_,
    new_n21161_, new_n21162_, new_n21163_, new_n21164_, new_n21165_,
    new_n21166_, new_n21167_, new_n21168_, new_n21169_, new_n21170_,
    new_n21171_, new_n21172_, new_n21173_, new_n21174_, new_n21175_,
    new_n21176_, new_n21177_, new_n21178_, new_n21179_, new_n21180_,
    new_n21181_, new_n21182_, new_n21183_, new_n21184_, new_n21185_,
    new_n21186_, new_n21187_, new_n21188_, new_n21189_, new_n21190_,
    new_n21191_, new_n21192_, new_n21193_, new_n21194_, new_n21195_,
    new_n21196_, new_n21197_, new_n21198_, new_n21199_, new_n21200_,
    new_n21201_, new_n21202_, new_n21203_, new_n21204_, new_n21205_,
    new_n21206_, new_n21207_, new_n21208_, new_n21209_, new_n21210_,
    new_n21211_, new_n21212_, new_n21213_, new_n21214_, new_n21215_,
    new_n21216_, new_n21217_, new_n21218_, new_n21219_, new_n21220_,
    new_n21221_, new_n21222_, new_n21223_, new_n21224_, new_n21225_,
    new_n21226_, new_n21227_, new_n21228_, new_n21229_, new_n21230_,
    new_n21231_, new_n21232_, new_n21233_, new_n21234_, new_n21235_,
    new_n21236_, new_n21237_, new_n21238_, new_n21239_, new_n21240_,
    new_n21241_, new_n21242_, new_n21243_, new_n21244_, new_n21245_,
    new_n21246_, new_n21247_, new_n21248_, new_n21249_, new_n21250_,
    new_n21251_, new_n21252_, new_n21253_, new_n21254_, new_n21255_,
    new_n21256_, new_n21257_, new_n21258_, new_n21259_, new_n21260_,
    new_n21261_, new_n21262_, new_n21263_, new_n21264_, new_n21265_,
    new_n21266_, new_n21267_, new_n21268_, new_n21269_, new_n21270_,
    new_n21271_, new_n21272_, new_n21273_, new_n21274_, new_n21275_,
    new_n21276_, new_n21277_, new_n21278_, new_n21279_, new_n21280_,
    new_n21281_, new_n21282_, new_n21283_, new_n21284_, new_n21285_,
    new_n21286_, new_n21287_, new_n21288_, new_n21289_, new_n21290_,
    new_n21291_, new_n21292_, new_n21293_, new_n21294_, new_n21295_,
    new_n21296_, new_n21297_, new_n21298_, new_n21299_, new_n21300_,
    new_n21301_, new_n21302_, new_n21303_, new_n21304_, new_n21305_,
    new_n21306_, new_n21307_, new_n21308_, new_n21309_, new_n21310_,
    new_n21311_, new_n21312_, new_n21313_, new_n21314_, new_n21315_,
    new_n21316_, new_n21317_, new_n21318_, new_n21319_, new_n21320_,
    new_n21321_, new_n21322_, new_n21323_, new_n21324_, new_n21325_,
    new_n21326_, new_n21327_, new_n21328_, new_n21329_, new_n21330_,
    new_n21331_, new_n21332_, new_n21333_, new_n21334_, new_n21335_,
    new_n21336_, new_n21337_, new_n21338_, new_n21339_, new_n21340_,
    new_n21341_, new_n21342_, new_n21343_, new_n21344_, new_n21345_,
    new_n21346_, new_n21347_, new_n21348_, new_n21349_, new_n21350_,
    new_n21351_, new_n21352_, new_n21353_, new_n21354_, new_n21355_,
    new_n21356_, new_n21357_, new_n21358_, new_n21359_, new_n21360_,
    new_n21361_, new_n21362_, new_n21363_, new_n21364_, new_n21365_,
    new_n21366_, new_n21367_, new_n21368_, new_n21369_, new_n21370_,
    new_n21371_, new_n21372_, new_n21373_, new_n21374_, new_n21375_,
    new_n21376_, new_n21377_, new_n21378_, new_n21379_, new_n21380_,
    new_n21381_, new_n21382_, new_n21383_, new_n21384_, new_n21385_,
    new_n21386_, new_n21387_, new_n21388_, new_n21389_, new_n21390_,
    new_n21391_, new_n21392_, new_n21393_, new_n21394_, new_n21395_,
    new_n21396_, new_n21397_, new_n21398_, new_n21399_, new_n21400_,
    new_n21401_, new_n21402_, new_n21403_, new_n21404_, new_n21405_,
    new_n21406_, new_n21407_, new_n21408_, new_n21409_, new_n21410_,
    new_n21411_, new_n21412_, new_n21413_, new_n21414_, new_n21415_,
    new_n21416_, new_n21417_, new_n21418_, new_n21419_, new_n21420_,
    new_n21421_, new_n21422_, new_n21423_, new_n21424_, new_n21425_,
    new_n21426_, new_n21427_, new_n21428_, new_n21429_, new_n21430_,
    new_n21431_, new_n21432_, new_n21433_, new_n21434_, new_n21435_,
    new_n21436_, new_n21437_, new_n21438_, new_n21439_, new_n21440_,
    new_n21441_, new_n21442_, new_n21443_, new_n21444_, new_n21445_,
    new_n21446_, new_n21447_, new_n21448_, new_n21449_, new_n21450_,
    new_n21451_, new_n21452_, new_n21453_, new_n21454_, new_n21455_,
    new_n21456_, new_n21457_, new_n21458_, new_n21459_, new_n21460_,
    new_n21461_, new_n21462_, new_n21463_, new_n21464_, new_n21465_,
    new_n21466_, new_n21467_, new_n21468_, new_n21469_, new_n21470_,
    new_n21471_, new_n21472_, new_n21473_, new_n21474_, new_n21475_,
    new_n21476_, new_n21477_, new_n21478_, new_n21479_, new_n21480_,
    new_n21481_, new_n21482_, new_n21483_, new_n21484_, new_n21485_,
    new_n21486_, new_n21487_, new_n21488_, new_n21489_, new_n21490_,
    new_n21491_, new_n21492_, new_n21493_, new_n21494_, new_n21495_,
    new_n21496_, new_n21497_, new_n21498_, new_n21499_, new_n21500_,
    new_n21501_, new_n21502_, new_n21503_, new_n21504_, new_n21505_,
    new_n21506_, new_n21507_, new_n21508_, new_n21509_, new_n21510_,
    new_n21511_, new_n21512_, new_n21513_, new_n21514_, new_n21515_,
    new_n21516_, new_n21517_, new_n21518_, new_n21519_, new_n21520_,
    new_n21521_, new_n21522_, new_n21523_, new_n21524_, new_n21525_,
    new_n21526_, new_n21527_, new_n21528_, new_n21529_, new_n21530_,
    new_n21531_, new_n21532_, new_n21533_, new_n21534_, new_n21535_,
    new_n21536_, new_n21537_, new_n21538_, new_n21539_, new_n21540_,
    new_n21541_, new_n21542_, new_n21543_, new_n21544_, new_n21545_,
    new_n21546_, new_n21547_, new_n21548_, new_n21549_, new_n21550_,
    new_n21551_, new_n21552_, new_n21553_, new_n21554_, new_n21555_,
    new_n21556_, new_n21557_, new_n21558_, new_n21559_, new_n21560_,
    new_n21561_, new_n21562_, new_n21563_, new_n21564_, new_n21565_,
    new_n21566_, new_n21567_, new_n21568_, new_n21569_, new_n21570_,
    new_n21571_, new_n21572_, new_n21573_, new_n21574_, new_n21575_,
    new_n21576_, new_n21577_, new_n21578_, new_n21579_, new_n21580_,
    new_n21581_, new_n21582_, new_n21583_, new_n21584_, new_n21585_,
    new_n21586_, new_n21587_, new_n21588_, new_n21589_, new_n21590_,
    new_n21591_, new_n21592_, new_n21593_, new_n21594_, new_n21595_,
    new_n21596_, new_n21597_, new_n21598_, new_n21599_, new_n21600_,
    new_n21601_, new_n21602_, new_n21603_, new_n21604_, new_n21605_,
    new_n21606_, new_n21607_, new_n21608_, new_n21609_, new_n21610_,
    new_n21611_, new_n21612_, new_n21613_, new_n21614_, new_n21615_,
    new_n21616_, new_n21617_, new_n21618_, new_n21619_, new_n21620_,
    new_n21621_, new_n21622_, new_n21623_, new_n21624_, new_n21625_,
    new_n21626_, new_n21627_, new_n21628_, new_n21629_, new_n21630_,
    new_n21631_, new_n21632_, new_n21633_, new_n21634_, new_n21635_,
    new_n21636_, new_n21637_, new_n21638_, new_n21639_, new_n21640_,
    new_n21641_, new_n21642_, new_n21643_, new_n21644_, new_n21645_,
    new_n21646_, new_n21647_, new_n21648_, new_n21649_, new_n21650_,
    new_n21651_, new_n21652_, new_n21653_, new_n21654_, new_n21655_,
    new_n21656_, new_n21657_, new_n21658_, new_n21659_, new_n21660_,
    new_n21661_, new_n21662_, new_n21663_, new_n21664_, new_n21665_,
    new_n21666_, new_n21667_, new_n21668_, new_n21669_, new_n21670_,
    new_n21671_, new_n21672_, new_n21673_, new_n21674_, new_n21675_,
    new_n21676_, new_n21677_, new_n21678_, new_n21679_, new_n21680_,
    new_n21681_, new_n21682_, new_n21683_, new_n21684_, new_n21685_,
    new_n21686_, new_n21687_, new_n21688_, new_n21689_, new_n21690_,
    new_n21691_, new_n21692_, new_n21693_, new_n21694_, new_n21695_,
    new_n21696_, new_n21697_, new_n21698_, new_n21699_, new_n21700_,
    new_n21701_, new_n21702_, new_n21703_, new_n21704_, new_n21705_,
    new_n21706_, new_n21707_, new_n21708_, new_n21709_, new_n21710_,
    new_n21711_, new_n21712_, new_n21713_, new_n21714_, new_n21715_,
    new_n21716_, new_n21717_, new_n21718_, new_n21719_, new_n21720_,
    new_n21721_, new_n21722_, new_n21723_, new_n21724_, new_n21725_,
    new_n21726_, new_n21727_, new_n21728_, new_n21729_, new_n21730_,
    new_n21731_, new_n21732_, new_n21733_, new_n21734_, new_n21735_,
    new_n21736_, new_n21737_, new_n21738_, new_n21739_, new_n21740_,
    new_n21741_, new_n21742_, new_n21743_, new_n21744_, new_n21745_,
    new_n21746_, new_n21747_, new_n21748_, new_n21749_, new_n21750_,
    new_n21751_, new_n21752_, new_n21753_, new_n21754_, new_n21755_,
    new_n21756_, new_n21757_, new_n21758_, new_n21759_, new_n21760_,
    new_n21761_, new_n21762_, new_n21763_, new_n21764_, new_n21765_,
    new_n21766_, new_n21767_, new_n21768_, new_n21769_, new_n21770_,
    new_n21771_, new_n21772_, new_n21773_, new_n21774_, new_n21775_,
    new_n21776_, new_n21777_, new_n21778_, new_n21779_, new_n21780_,
    new_n21781_, new_n21782_, new_n21783_, new_n21784_, new_n21785_,
    new_n21786_, new_n21787_, new_n21788_, new_n21789_, new_n21790_,
    new_n21791_, new_n21792_, new_n21793_, new_n21794_, new_n21795_,
    new_n21796_, new_n21797_, new_n21798_, new_n21799_, new_n21800_,
    new_n21801_, new_n21802_, new_n21803_, new_n21804_, new_n21805_,
    new_n21806_, new_n21807_, new_n21808_, new_n21809_, new_n21810_,
    new_n21811_, new_n21812_, new_n21814_, new_n21815_, new_n21816_,
    new_n21817_, new_n21818_, new_n21819_, new_n21820_, new_n21821_,
    new_n21822_, new_n21823_, new_n21824_, new_n21825_, new_n21826_,
    new_n21827_, new_n21828_, new_n21829_, new_n21830_, new_n21831_,
    new_n21832_, new_n21833_, new_n21834_, new_n21835_, new_n21836_,
    new_n21837_, new_n21838_, new_n21839_, new_n21840_, new_n21841_,
    new_n21842_, new_n21843_, new_n21844_, new_n21845_, new_n21846_,
    new_n21847_, new_n21848_, new_n21849_, new_n21850_, new_n21851_,
    new_n21852_, new_n21853_, new_n21854_, new_n21855_, new_n21856_,
    new_n21857_, new_n21858_, new_n21859_, new_n21860_, new_n21861_,
    new_n21862_, new_n21863_, new_n21864_, new_n21865_, new_n21866_,
    new_n21867_, new_n21868_, new_n21869_, new_n21870_, new_n21871_,
    new_n21872_, new_n21873_, new_n21874_, new_n21875_, new_n21876_,
    new_n21877_, new_n21878_, new_n21879_, new_n21880_, new_n21881_,
    new_n21882_, new_n21883_, new_n21884_, new_n21885_, new_n21886_,
    new_n21887_, new_n21888_, new_n21889_, new_n21890_, new_n21891_,
    new_n21892_, new_n21893_, new_n21894_, new_n21895_, new_n21896_,
    new_n21897_, new_n21898_, new_n21899_, new_n21900_, new_n21901_,
    new_n21902_, new_n21903_, new_n21904_, new_n21905_, new_n21906_,
    new_n21907_, new_n21908_, new_n21909_, new_n21910_, new_n21911_,
    new_n21912_, new_n21913_, new_n21914_, new_n21915_, new_n21916_,
    new_n21917_, new_n21918_, new_n21919_, new_n21920_, new_n21921_,
    new_n21922_, new_n21923_, new_n21924_, new_n21925_, new_n21926_,
    new_n21927_, new_n21928_, new_n21929_, new_n21930_, new_n21931_,
    new_n21932_, new_n21933_, new_n21934_, new_n21935_, new_n21936_,
    new_n21937_, new_n21938_, new_n21939_, new_n21940_, new_n21941_,
    new_n21942_, new_n21943_, new_n21944_, new_n21945_, new_n21946_,
    new_n21947_, new_n21948_, new_n21949_, new_n21950_, new_n21951_,
    new_n21952_, new_n21953_, new_n21954_, new_n21955_, new_n21956_,
    new_n21957_, new_n21958_, new_n21959_, new_n21960_, new_n21961_,
    new_n21962_, new_n21963_, new_n21964_, new_n21965_, new_n21966_,
    new_n21967_, new_n21968_, new_n21969_, new_n21970_, new_n21971_,
    new_n21972_, new_n21973_, new_n21974_, new_n21975_, new_n21976_,
    new_n21977_, new_n21978_, new_n21979_, new_n21980_, new_n21981_,
    new_n21982_, new_n21983_, new_n21984_, new_n21985_, new_n21986_,
    new_n21987_, new_n21988_, new_n21989_, new_n21990_, new_n21991_,
    new_n21992_, new_n21993_, new_n21994_, new_n21995_, new_n21996_,
    new_n21997_, new_n21998_, new_n21999_, new_n22000_, new_n22001_,
    new_n22002_, new_n22003_, new_n22004_, new_n22005_, new_n22006_,
    new_n22007_, new_n22008_, new_n22009_, new_n22010_, new_n22011_,
    new_n22012_, new_n22013_, new_n22014_, new_n22015_, new_n22016_,
    new_n22017_, new_n22018_, new_n22019_, new_n22020_, new_n22021_,
    new_n22022_, new_n22023_, new_n22024_, new_n22025_, new_n22026_,
    new_n22027_, new_n22028_, new_n22029_, new_n22030_, new_n22031_,
    new_n22032_, new_n22033_, new_n22034_, new_n22035_, new_n22036_,
    new_n22037_, new_n22038_, new_n22039_, new_n22040_, new_n22041_,
    new_n22042_, new_n22043_, new_n22044_, new_n22045_, new_n22046_,
    new_n22047_, new_n22048_, new_n22049_, new_n22050_, new_n22051_,
    new_n22052_, new_n22053_, new_n22054_, new_n22055_, new_n22056_,
    new_n22057_, new_n22058_, new_n22059_, new_n22060_, new_n22061_,
    new_n22062_, new_n22063_, new_n22064_, new_n22065_, new_n22066_,
    new_n22067_, new_n22068_, new_n22069_, new_n22070_, new_n22071_,
    new_n22072_, new_n22073_, new_n22074_, new_n22075_, new_n22076_,
    new_n22077_, new_n22078_, new_n22079_, new_n22080_, new_n22081_,
    new_n22082_, new_n22083_, new_n22084_, new_n22085_, new_n22086_,
    new_n22087_, new_n22088_, new_n22089_, new_n22090_, new_n22091_,
    new_n22092_, new_n22093_, new_n22094_, new_n22095_, new_n22096_,
    new_n22097_, new_n22098_, new_n22099_, new_n22100_, new_n22101_,
    new_n22102_, new_n22103_, new_n22104_, new_n22105_, new_n22106_,
    new_n22107_, new_n22108_, new_n22109_, new_n22110_, new_n22111_,
    new_n22112_, new_n22113_, new_n22114_, new_n22115_, new_n22116_,
    new_n22117_, new_n22118_, new_n22119_, new_n22120_, new_n22121_,
    new_n22122_, new_n22123_, new_n22124_, new_n22125_, new_n22126_,
    new_n22127_, new_n22128_, new_n22129_, new_n22130_, new_n22131_,
    new_n22132_, new_n22133_, new_n22134_, new_n22135_, new_n22136_,
    new_n22137_, new_n22138_, new_n22139_, new_n22140_, new_n22141_,
    new_n22142_, new_n22143_, new_n22144_, new_n22145_, new_n22146_,
    new_n22147_, new_n22148_, new_n22149_, new_n22150_, new_n22151_,
    new_n22152_, new_n22153_, new_n22154_, new_n22155_, new_n22156_,
    new_n22157_, new_n22158_, new_n22159_, new_n22160_, new_n22161_,
    new_n22162_, new_n22163_, new_n22164_, new_n22165_, new_n22166_,
    new_n22167_, new_n22168_, new_n22169_, new_n22170_, new_n22171_,
    new_n22172_, new_n22173_, new_n22174_, new_n22175_, new_n22176_,
    new_n22177_, new_n22178_, new_n22179_, new_n22180_, new_n22181_,
    new_n22182_, new_n22183_, new_n22184_, new_n22185_, new_n22186_,
    new_n22187_, new_n22188_, new_n22189_, new_n22190_, new_n22191_,
    new_n22192_, new_n22193_, new_n22194_, new_n22195_, new_n22196_,
    new_n22197_, new_n22198_, new_n22199_, new_n22200_, new_n22201_,
    new_n22202_, new_n22203_, new_n22204_, new_n22205_, new_n22206_,
    new_n22207_, new_n22208_, new_n22209_, new_n22210_, new_n22211_,
    new_n22212_, new_n22213_, new_n22214_, new_n22215_, new_n22216_,
    new_n22217_, new_n22218_, new_n22219_, new_n22220_, new_n22221_,
    new_n22222_, new_n22223_, new_n22224_, new_n22225_, new_n22226_,
    new_n22227_, new_n22228_, new_n22229_, new_n22230_, new_n22231_,
    new_n22232_, new_n22233_, new_n22234_, new_n22235_, new_n22236_,
    new_n22237_, new_n22238_, new_n22239_, new_n22240_, new_n22241_,
    new_n22242_, new_n22243_, new_n22244_, new_n22245_, new_n22246_,
    new_n22247_, new_n22248_, new_n22249_, new_n22250_, new_n22251_,
    new_n22252_, new_n22253_, new_n22254_, new_n22255_, new_n22256_,
    new_n22257_, new_n22258_, new_n22259_, new_n22260_, new_n22261_,
    new_n22262_, new_n22263_, new_n22264_, new_n22265_, new_n22266_,
    new_n22267_, new_n22268_, new_n22269_, new_n22270_, new_n22271_,
    new_n22272_, new_n22273_, new_n22274_, new_n22275_, new_n22276_,
    new_n22277_, new_n22278_, new_n22279_, new_n22280_, new_n22281_,
    new_n22282_, new_n22283_, new_n22284_, new_n22285_, new_n22286_,
    new_n22287_, new_n22288_, new_n22289_, new_n22290_, new_n22291_,
    new_n22292_, new_n22293_, new_n22294_, new_n22295_, new_n22296_,
    new_n22297_, new_n22298_, new_n22299_, new_n22300_, new_n22301_,
    new_n22302_, new_n22303_, new_n22304_, new_n22305_, new_n22306_,
    new_n22307_, new_n22308_, new_n22309_, new_n22310_, new_n22311_,
    new_n22312_, new_n22313_, new_n22314_, new_n22315_, new_n22316_,
    new_n22317_, new_n22318_, new_n22319_, new_n22320_, new_n22321_,
    new_n22322_, new_n22323_, new_n22324_, new_n22325_, new_n22326_,
    new_n22327_, new_n22328_, new_n22329_, new_n22330_, new_n22331_,
    new_n22332_, new_n22333_, new_n22334_, new_n22335_, new_n22336_,
    new_n22337_, new_n22338_, new_n22339_, new_n22340_, new_n22341_,
    new_n22342_, new_n22343_, new_n22344_, new_n22345_, new_n22346_,
    new_n22347_, new_n22348_, new_n22349_, new_n22350_, new_n22351_,
    new_n22352_, new_n22353_, new_n22354_, new_n22355_, new_n22356_,
    new_n22357_, new_n22358_, new_n22359_, new_n22360_, new_n22361_,
    new_n22362_, new_n22363_, new_n22364_, new_n22365_, new_n22366_,
    new_n22367_, new_n22368_, new_n22369_, new_n22370_, new_n22371_,
    new_n22372_, new_n22373_, new_n22374_, new_n22375_, new_n22376_,
    new_n22377_, new_n22378_, new_n22379_, new_n22380_, new_n22381_,
    new_n22382_, new_n22383_, new_n22384_, new_n22385_, new_n22386_,
    new_n22387_, new_n22388_, new_n22389_, new_n22390_, new_n22391_,
    new_n22392_, new_n22393_, new_n22394_, new_n22395_, new_n22396_,
    new_n22397_, new_n22398_, new_n22399_, new_n22400_, new_n22401_,
    new_n22402_, new_n22403_, new_n22404_, new_n22405_, new_n22406_,
    new_n22407_, new_n22408_, new_n22409_, new_n22410_, new_n22411_,
    new_n22412_, new_n22413_, new_n22414_, new_n22415_, new_n22416_,
    new_n22417_, new_n22418_, new_n22419_, new_n22420_, new_n22421_,
    new_n22422_, new_n22423_, new_n22424_, new_n22425_, new_n22426_,
    new_n22427_, new_n22428_, new_n22429_, new_n22430_, new_n22431_,
    new_n22432_, new_n22433_, new_n22434_, new_n22435_, new_n22436_,
    new_n22437_, new_n22438_, new_n22439_, new_n22440_, new_n22441_,
    new_n22442_, new_n22443_, new_n22444_, new_n22445_, new_n22446_,
    new_n22447_, new_n22448_, new_n22449_, new_n22450_, new_n22451_,
    new_n22452_, new_n22453_, new_n22454_, new_n22455_, new_n22456_,
    new_n22457_, new_n22458_, new_n22459_, new_n22460_, new_n22461_,
    new_n22462_, new_n22463_, new_n22464_, new_n22465_, new_n22466_,
    new_n22467_, new_n22468_, new_n22469_, new_n22470_, new_n22471_,
    new_n22472_, new_n22473_, new_n22474_, new_n22475_, new_n22476_,
    new_n22477_, new_n22478_, new_n22479_, new_n22480_, new_n22481_,
    new_n22482_, new_n22484_, new_n22485_, new_n22486_, new_n22487_,
    new_n22488_, new_n22489_, new_n22490_, new_n22491_, new_n22492_,
    new_n22493_, new_n22494_, new_n22495_, new_n22496_, new_n22497_,
    new_n22498_, new_n22499_, new_n22500_, new_n22501_, new_n22502_,
    new_n22503_, new_n22504_, new_n22505_, new_n22506_, new_n22507_,
    new_n22508_, new_n22509_, new_n22510_, new_n22511_, new_n22512_,
    new_n22513_, new_n22514_, new_n22515_, new_n22516_, new_n22517_,
    new_n22518_, new_n22519_, new_n22520_, new_n22521_, new_n22522_,
    new_n22523_, new_n22524_, new_n22525_, new_n22526_, new_n22527_,
    new_n22528_, new_n22529_, new_n22530_, new_n22531_, new_n22532_,
    new_n22533_, new_n22534_, new_n22535_, new_n22536_, new_n22537_,
    new_n22538_, new_n22539_, new_n22540_, new_n22541_, new_n22542_,
    new_n22543_, new_n22544_, new_n22545_, new_n22546_, new_n22547_,
    new_n22548_, new_n22549_, new_n22550_, new_n22551_, new_n22552_,
    new_n22553_, new_n22554_, new_n22555_, new_n22556_, new_n22557_,
    new_n22558_, new_n22559_, new_n22560_, new_n22561_, new_n22562_,
    new_n22563_, new_n22564_, new_n22565_, new_n22566_, new_n22567_,
    new_n22568_, new_n22569_, new_n22570_, new_n22571_, new_n22572_,
    new_n22573_, new_n22574_, new_n22575_, new_n22576_, new_n22577_,
    new_n22578_, new_n22579_, new_n22580_, new_n22581_, new_n22582_,
    new_n22583_, new_n22584_, new_n22585_, new_n22586_, new_n22587_,
    new_n22588_, new_n22589_, new_n22590_, new_n22591_, new_n22592_,
    new_n22593_, new_n22594_, new_n22595_, new_n22596_, new_n22597_,
    new_n22598_, new_n22599_, new_n22600_, new_n22601_, new_n22602_,
    new_n22603_, new_n22604_, new_n22605_, new_n22606_, new_n22607_,
    new_n22608_, new_n22609_, new_n22610_, new_n22611_, new_n22612_,
    new_n22613_, new_n22614_, new_n22615_, new_n22616_, new_n22617_,
    new_n22618_, new_n22619_, new_n22620_, new_n22621_, new_n22622_,
    new_n22623_, new_n22624_, new_n22625_, new_n22626_, new_n22627_,
    new_n22628_, new_n22629_, new_n22630_, new_n22631_, new_n22632_,
    new_n22633_, new_n22634_, new_n22635_, new_n22636_, new_n22637_,
    new_n22638_, new_n22639_, new_n22640_, new_n22641_, new_n22642_,
    new_n22643_, new_n22644_, new_n22645_, new_n22646_, new_n22647_,
    new_n22648_, new_n22649_, new_n22650_, new_n22651_, new_n22652_,
    new_n22653_, new_n22654_, new_n22655_, new_n22656_, new_n22657_,
    new_n22658_, new_n22659_, new_n22660_, new_n22661_, new_n22662_,
    new_n22663_, new_n22664_, new_n22665_, new_n22666_, new_n22667_,
    new_n22668_, new_n22669_, new_n22670_, new_n22671_, new_n22672_,
    new_n22673_, new_n22674_, new_n22675_, new_n22676_, new_n22677_,
    new_n22678_, new_n22679_, new_n22680_, new_n22681_, new_n22682_,
    new_n22683_, new_n22684_, new_n22685_, new_n22686_, new_n22687_,
    new_n22688_, new_n22689_, new_n22690_, new_n22691_, new_n22692_,
    new_n22693_, new_n22694_, new_n22695_, new_n22696_, new_n22697_,
    new_n22698_, new_n22699_, new_n22700_, new_n22701_, new_n22702_,
    new_n22703_, new_n22704_, new_n22705_, new_n22706_, new_n22707_,
    new_n22708_, new_n22709_, new_n22710_, new_n22711_, new_n22712_,
    new_n22713_, new_n22714_, new_n22715_, new_n22716_, new_n22717_,
    new_n22718_, new_n22719_, new_n22720_, new_n22721_, new_n22722_,
    new_n22723_, new_n22724_, new_n22725_, new_n22726_, new_n22727_,
    new_n22728_, new_n22729_, new_n22730_, new_n22731_, new_n22732_,
    new_n22733_, new_n22734_, new_n22735_, new_n22736_, new_n22737_,
    new_n22738_, new_n22739_, new_n22740_, new_n22741_, new_n22742_,
    new_n22743_, new_n22744_, new_n22745_, new_n22746_, new_n22747_,
    new_n22748_, new_n22749_, new_n22750_, new_n22751_, new_n22752_,
    new_n22753_, new_n22754_, new_n22755_, new_n22756_, new_n22757_,
    new_n22758_, new_n22759_, new_n22760_, new_n22761_, new_n22762_,
    new_n22763_, new_n22764_, new_n22765_, new_n22766_, new_n22767_,
    new_n22768_, new_n22769_, new_n22770_, new_n22771_, new_n22772_,
    new_n22773_, new_n22774_, new_n22775_, new_n22776_, new_n22777_,
    new_n22778_, new_n22779_, new_n22780_, new_n22781_, new_n22782_,
    new_n22783_, new_n22784_, new_n22785_, new_n22786_, new_n22787_,
    new_n22788_, new_n22789_, new_n22790_, new_n22791_, new_n22792_,
    new_n22793_, new_n22794_, new_n22795_, new_n22796_, new_n22797_,
    new_n22798_, new_n22799_, new_n22800_, new_n22801_, new_n22802_,
    new_n22803_, new_n22804_, new_n22805_, new_n22806_, new_n22807_,
    new_n22808_, new_n22809_, new_n22810_, new_n22811_, new_n22812_,
    new_n22813_, new_n22814_, new_n22815_, new_n22816_, new_n22817_,
    new_n22818_, new_n22819_, new_n22820_, new_n22821_, new_n22822_,
    new_n22823_, new_n22824_, new_n22825_, new_n22826_, new_n22827_,
    new_n22828_, new_n22829_, new_n22830_, new_n22831_, new_n22832_,
    new_n22833_, new_n22834_, new_n22835_, new_n22836_, new_n22837_,
    new_n22838_, new_n22839_, new_n22840_, new_n22841_, new_n22842_,
    new_n22843_, new_n22844_, new_n22845_, new_n22846_, new_n22847_,
    new_n22848_, new_n22849_, new_n22850_, new_n22851_, new_n22852_,
    new_n22853_, new_n22854_, new_n22855_, new_n22856_, new_n22857_,
    new_n22858_, new_n22859_, new_n22860_, new_n22861_, new_n22862_,
    new_n22863_, new_n22864_, new_n22865_, new_n22866_, new_n22867_,
    new_n22868_, new_n22869_, new_n22870_, new_n22871_, new_n22872_,
    new_n22873_, new_n22874_, new_n22875_, new_n22876_, new_n22877_,
    new_n22878_, new_n22879_, new_n22880_, new_n22881_, new_n22882_,
    new_n22883_, new_n22884_, new_n22885_, new_n22886_, new_n22887_,
    new_n22888_, new_n22889_, new_n22890_, new_n22891_, new_n22892_,
    new_n22893_, new_n22894_, new_n22895_, new_n22896_, new_n22897_,
    new_n22898_, new_n22899_, new_n22900_, new_n22901_, new_n22902_,
    new_n22903_, new_n22904_, new_n22905_, new_n22906_, new_n22907_,
    new_n22908_, new_n22909_, new_n22910_, new_n22911_, new_n22912_,
    new_n22913_, new_n22914_, new_n22915_, new_n22916_, new_n22917_,
    new_n22918_, new_n22919_, new_n22920_, new_n22921_, new_n22922_,
    new_n22923_, new_n22924_, new_n22925_, new_n22926_, new_n22927_,
    new_n22928_, new_n22929_, new_n22930_, new_n22931_, new_n22932_,
    new_n22933_, new_n22934_, new_n22935_, new_n22936_, new_n22937_,
    new_n22938_, new_n22939_, new_n22940_, new_n22941_, new_n22942_,
    new_n22943_, new_n22944_, new_n22945_, new_n22946_, new_n22947_,
    new_n22948_, new_n22949_, new_n22950_, new_n22951_, new_n22952_,
    new_n22953_, new_n22954_, new_n22955_, new_n22956_, new_n22957_,
    new_n22958_, new_n22959_, new_n22960_, new_n22961_, new_n22962_,
    new_n22963_, new_n22964_, new_n22965_, new_n22966_, new_n22967_,
    new_n22968_, new_n22969_, new_n22970_, new_n22971_, new_n22972_,
    new_n22973_, new_n22974_, new_n22975_, new_n22976_, new_n22977_,
    new_n22978_, new_n22979_, new_n22980_, new_n22981_, new_n22982_,
    new_n22983_, new_n22984_, new_n22985_, new_n22986_, new_n22987_,
    new_n22988_, new_n22989_, new_n22990_, new_n22991_, new_n22992_,
    new_n22993_, new_n22994_, new_n22995_, new_n22996_, new_n22997_,
    new_n22998_, new_n22999_, new_n23000_, new_n23001_, new_n23002_,
    new_n23003_, new_n23004_, new_n23005_, new_n23006_, new_n23007_,
    new_n23008_, new_n23009_, new_n23010_, new_n23011_, new_n23012_,
    new_n23013_, new_n23014_, new_n23015_, new_n23016_, new_n23017_,
    new_n23018_, new_n23019_, new_n23020_, new_n23021_, new_n23022_,
    new_n23023_, new_n23024_, new_n23025_, new_n23026_, new_n23027_,
    new_n23028_, new_n23029_, new_n23030_, new_n23031_, new_n23032_,
    new_n23033_, new_n23034_, new_n23035_, new_n23036_, new_n23037_,
    new_n23038_, new_n23039_, new_n23040_, new_n23041_, new_n23042_,
    new_n23043_, new_n23044_, new_n23045_, new_n23046_, new_n23047_,
    new_n23048_, new_n23049_, new_n23050_, new_n23051_, new_n23052_,
    new_n23053_, new_n23054_, new_n23055_, new_n23056_, new_n23057_,
    new_n23058_, new_n23059_, new_n23060_, new_n23061_, new_n23062_,
    new_n23063_, new_n23064_, new_n23065_, new_n23066_, new_n23067_,
    new_n23068_, new_n23069_, new_n23070_, new_n23071_, new_n23072_,
    new_n23073_, new_n23074_, new_n23075_, new_n23076_, new_n23077_,
    new_n23078_, new_n23079_, new_n23080_, new_n23081_, new_n23082_,
    new_n23083_, new_n23084_, new_n23085_, new_n23086_, new_n23087_,
    new_n23088_, new_n23089_, new_n23090_, new_n23091_, new_n23092_,
    new_n23093_, new_n23094_, new_n23095_, new_n23096_, new_n23097_,
    new_n23098_, new_n23099_, new_n23100_, new_n23101_, new_n23102_,
    new_n23103_, new_n23104_, new_n23105_, new_n23106_, new_n23107_,
    new_n23108_, new_n23109_, new_n23110_, new_n23111_, new_n23112_,
    new_n23113_, new_n23114_, new_n23115_, new_n23116_, new_n23117_,
    new_n23118_, new_n23119_, new_n23120_, new_n23121_, new_n23122_,
    new_n23123_, new_n23124_, new_n23125_, new_n23126_, new_n23127_,
    new_n23128_, new_n23129_, new_n23130_, new_n23131_, new_n23132_,
    new_n23133_, new_n23134_, new_n23135_, new_n23136_, new_n23137_,
    new_n23138_, new_n23139_, new_n23140_, new_n23141_, new_n23142_,
    new_n23143_, new_n23144_, new_n23145_, new_n23146_, new_n23147_,
    new_n23148_, new_n23149_, new_n23150_, new_n23151_, new_n23152_,
    new_n23153_, new_n23154_, new_n23155_, new_n23156_, new_n23157_,
    new_n23158_, new_n23159_, new_n23160_, new_n23161_, new_n23162_,
    new_n23163_, new_n23164_, new_n23165_, new_n23166_, new_n23167_,
    new_n23168_, new_n23169_, new_n23170_, new_n23171_, new_n23172_,
    new_n23173_, new_n23174_, new_n23175_, new_n23176_, new_n23177_,
    new_n23178_, new_n23179_, new_n23180_, new_n23181_, new_n23182_,
    new_n23183_, new_n23184_, new_n23185_, new_n23186_, new_n23187_,
    new_n23188_, new_n23189_, new_n23190_, new_n23191_, new_n23192_,
    new_n23193_, new_n23194_, new_n23195_, new_n23196_, new_n23198_,
    new_n23199_, new_n23200_, new_n23201_, new_n23202_, new_n23203_,
    new_n23204_, new_n23205_, new_n23206_, new_n23207_, new_n23208_,
    new_n23209_, new_n23210_, new_n23211_, new_n23212_, new_n23213_,
    new_n23214_, new_n23215_, new_n23216_, new_n23217_, new_n23218_,
    new_n23219_, new_n23220_, new_n23221_, new_n23222_, new_n23223_,
    new_n23224_, new_n23225_, new_n23226_, new_n23227_, new_n23228_,
    new_n23229_, new_n23230_, new_n23231_, new_n23232_, new_n23233_,
    new_n23234_, new_n23235_, new_n23236_, new_n23237_, new_n23238_,
    new_n23239_, new_n23240_, new_n23241_, new_n23242_, new_n23243_,
    new_n23244_, new_n23245_, new_n23246_, new_n23247_, new_n23248_,
    new_n23249_, new_n23250_, new_n23251_, new_n23252_, new_n23253_,
    new_n23254_, new_n23255_, new_n23256_, new_n23257_, new_n23258_,
    new_n23259_, new_n23260_, new_n23261_, new_n23262_, new_n23263_,
    new_n23264_, new_n23265_, new_n23266_, new_n23267_, new_n23268_,
    new_n23269_, new_n23270_, new_n23271_, new_n23272_, new_n23273_,
    new_n23274_, new_n23275_, new_n23276_, new_n23277_, new_n23278_,
    new_n23279_, new_n23280_, new_n23281_, new_n23282_, new_n23283_,
    new_n23284_, new_n23285_, new_n23286_, new_n23287_, new_n23288_,
    new_n23289_, new_n23290_, new_n23291_, new_n23292_, new_n23293_,
    new_n23294_, new_n23295_, new_n23296_, new_n23297_, new_n23298_,
    new_n23299_, new_n23300_, new_n23301_, new_n23302_, new_n23303_,
    new_n23304_, new_n23305_, new_n23306_, new_n23307_, new_n23308_,
    new_n23309_, new_n23310_, new_n23311_, new_n23312_, new_n23313_,
    new_n23314_, new_n23315_, new_n23316_, new_n23317_, new_n23318_,
    new_n23319_, new_n23320_, new_n23321_, new_n23322_, new_n23323_,
    new_n23324_, new_n23325_, new_n23326_, new_n23327_, new_n23328_,
    new_n23329_, new_n23330_, new_n23331_, new_n23332_, new_n23333_,
    new_n23334_, new_n23335_, new_n23336_, new_n23337_, new_n23338_,
    new_n23339_, new_n23340_, new_n23341_, new_n23342_, new_n23343_,
    new_n23344_, new_n23345_, new_n23346_, new_n23347_, new_n23348_,
    new_n23349_, new_n23350_, new_n23351_, new_n23352_, new_n23353_,
    new_n23354_, new_n23355_, new_n23356_, new_n23357_, new_n23358_,
    new_n23359_, new_n23360_, new_n23361_, new_n23362_, new_n23363_,
    new_n23364_, new_n23365_, new_n23366_, new_n23367_, new_n23368_,
    new_n23369_, new_n23370_, new_n23371_, new_n23372_, new_n23373_,
    new_n23374_, new_n23375_, new_n23376_, new_n23377_, new_n23378_,
    new_n23379_, new_n23380_, new_n23381_, new_n23382_, new_n23383_,
    new_n23384_, new_n23385_, new_n23386_, new_n23387_, new_n23388_,
    new_n23389_, new_n23390_, new_n23391_, new_n23392_, new_n23393_,
    new_n23394_, new_n23395_, new_n23396_, new_n23397_, new_n23398_,
    new_n23399_, new_n23400_, new_n23401_, new_n23402_, new_n23403_,
    new_n23404_, new_n23405_, new_n23406_, new_n23407_, new_n23408_,
    new_n23409_, new_n23410_, new_n23411_, new_n23412_, new_n23413_,
    new_n23414_, new_n23415_, new_n23416_, new_n23417_, new_n23418_,
    new_n23419_, new_n23420_, new_n23421_, new_n23422_, new_n23423_,
    new_n23424_, new_n23425_, new_n23426_, new_n23427_, new_n23428_,
    new_n23429_, new_n23430_, new_n23431_, new_n23432_, new_n23433_,
    new_n23434_, new_n23435_, new_n23436_, new_n23437_, new_n23438_,
    new_n23439_, new_n23440_, new_n23441_, new_n23442_, new_n23443_,
    new_n23444_, new_n23445_, new_n23446_, new_n23447_, new_n23448_,
    new_n23449_, new_n23450_, new_n23451_, new_n23452_, new_n23453_,
    new_n23454_, new_n23455_, new_n23456_, new_n23457_, new_n23458_,
    new_n23459_, new_n23460_, new_n23461_, new_n23462_, new_n23463_,
    new_n23464_, new_n23465_, new_n23466_, new_n23467_, new_n23468_,
    new_n23469_, new_n23470_, new_n23471_, new_n23472_, new_n23473_,
    new_n23474_, new_n23475_, new_n23476_, new_n23477_, new_n23478_,
    new_n23479_, new_n23480_, new_n23481_, new_n23482_, new_n23483_,
    new_n23484_, new_n23485_, new_n23486_, new_n23487_, new_n23488_,
    new_n23489_, new_n23490_, new_n23491_, new_n23492_, new_n23493_,
    new_n23494_, new_n23495_, new_n23496_, new_n23497_, new_n23498_,
    new_n23499_, new_n23500_, new_n23501_, new_n23502_, new_n23503_,
    new_n23504_, new_n23505_, new_n23506_, new_n23507_, new_n23508_,
    new_n23509_, new_n23510_, new_n23511_, new_n23512_, new_n23513_,
    new_n23514_, new_n23515_, new_n23516_, new_n23517_, new_n23518_,
    new_n23519_, new_n23520_, new_n23521_, new_n23522_, new_n23523_,
    new_n23524_, new_n23525_, new_n23526_, new_n23527_, new_n23528_,
    new_n23529_, new_n23530_, new_n23531_, new_n23532_, new_n23533_,
    new_n23534_, new_n23535_, new_n23536_, new_n23537_, new_n23538_,
    new_n23539_, new_n23540_, new_n23541_, new_n23542_, new_n23543_,
    new_n23544_, new_n23545_, new_n23546_, new_n23547_, new_n23548_,
    new_n23549_, new_n23550_, new_n23551_, new_n23552_, new_n23553_,
    new_n23554_, new_n23555_, new_n23556_, new_n23557_, new_n23558_,
    new_n23559_, new_n23560_, new_n23561_, new_n23562_, new_n23563_,
    new_n23564_, new_n23565_, new_n23566_, new_n23567_, new_n23568_,
    new_n23569_, new_n23570_, new_n23571_, new_n23572_, new_n23573_,
    new_n23574_, new_n23575_, new_n23576_, new_n23577_, new_n23578_,
    new_n23579_, new_n23580_, new_n23581_, new_n23582_, new_n23583_,
    new_n23584_, new_n23585_, new_n23586_, new_n23587_, new_n23588_,
    new_n23589_, new_n23590_, new_n23591_, new_n23592_, new_n23593_,
    new_n23594_, new_n23595_, new_n23596_, new_n23597_, new_n23598_,
    new_n23599_, new_n23600_, new_n23601_, new_n23602_, new_n23603_,
    new_n23604_, new_n23605_, new_n23606_, new_n23607_, new_n23608_,
    new_n23609_, new_n23610_, new_n23611_, new_n23612_, new_n23613_,
    new_n23614_, new_n23615_, new_n23616_, new_n23617_, new_n23618_,
    new_n23619_, new_n23620_, new_n23621_, new_n23622_, new_n23623_,
    new_n23624_, new_n23625_, new_n23626_, new_n23627_, new_n23628_,
    new_n23629_, new_n23630_, new_n23631_, new_n23632_, new_n23633_,
    new_n23634_, new_n23635_, new_n23636_, new_n23637_, new_n23638_,
    new_n23639_, new_n23640_, new_n23641_, new_n23642_, new_n23643_,
    new_n23644_, new_n23645_, new_n23646_, new_n23647_, new_n23648_,
    new_n23649_, new_n23650_, new_n23651_, new_n23652_, new_n23653_,
    new_n23654_, new_n23655_, new_n23656_, new_n23657_, new_n23658_,
    new_n23659_, new_n23660_, new_n23661_, new_n23662_, new_n23663_,
    new_n23664_, new_n23665_, new_n23666_, new_n23667_, new_n23668_,
    new_n23669_, new_n23670_, new_n23671_, new_n23672_, new_n23673_,
    new_n23674_, new_n23675_, new_n23676_, new_n23677_, new_n23678_,
    new_n23679_, new_n23680_, new_n23681_, new_n23682_, new_n23683_,
    new_n23684_, new_n23685_, new_n23686_, new_n23687_, new_n23688_,
    new_n23689_, new_n23690_, new_n23691_, new_n23692_, new_n23693_,
    new_n23694_, new_n23695_, new_n23696_, new_n23697_, new_n23698_,
    new_n23699_, new_n23700_, new_n23701_, new_n23702_, new_n23703_,
    new_n23704_, new_n23705_, new_n23706_, new_n23707_, new_n23708_,
    new_n23709_, new_n23710_, new_n23711_, new_n23712_, new_n23713_,
    new_n23714_, new_n23715_, new_n23716_, new_n23717_, new_n23718_,
    new_n23719_, new_n23720_, new_n23721_, new_n23722_, new_n23723_,
    new_n23724_, new_n23725_, new_n23726_, new_n23727_, new_n23728_,
    new_n23729_, new_n23730_, new_n23731_, new_n23732_, new_n23733_,
    new_n23734_, new_n23735_, new_n23736_, new_n23737_, new_n23738_,
    new_n23739_, new_n23740_, new_n23741_, new_n23742_, new_n23743_,
    new_n23744_, new_n23745_, new_n23746_, new_n23747_, new_n23748_,
    new_n23749_, new_n23750_, new_n23751_, new_n23752_, new_n23753_,
    new_n23754_, new_n23755_, new_n23756_, new_n23757_, new_n23758_,
    new_n23759_, new_n23760_, new_n23761_, new_n23762_, new_n23763_,
    new_n23764_, new_n23765_, new_n23766_, new_n23767_, new_n23768_,
    new_n23769_, new_n23770_, new_n23771_, new_n23772_, new_n23773_,
    new_n23774_, new_n23775_, new_n23776_, new_n23777_, new_n23778_,
    new_n23779_, new_n23780_, new_n23781_, new_n23782_, new_n23783_,
    new_n23784_, new_n23785_, new_n23786_, new_n23787_, new_n23788_,
    new_n23789_, new_n23790_, new_n23791_, new_n23792_, new_n23793_,
    new_n23794_, new_n23795_, new_n23796_, new_n23797_, new_n23798_,
    new_n23799_, new_n23800_, new_n23801_, new_n23802_, new_n23803_,
    new_n23804_, new_n23805_, new_n23806_, new_n23807_, new_n23808_,
    new_n23809_, new_n23810_, new_n23811_, new_n23812_, new_n23813_,
    new_n23814_, new_n23815_, new_n23816_, new_n23817_, new_n23818_,
    new_n23819_, new_n23820_, new_n23821_, new_n23822_, new_n23823_,
    new_n23824_, new_n23825_, new_n23826_, new_n23827_, new_n23828_,
    new_n23829_, new_n23830_, new_n23831_, new_n23832_, new_n23833_,
    new_n23834_, new_n23835_, new_n23836_, new_n23837_, new_n23838_,
    new_n23839_, new_n23840_, new_n23841_, new_n23842_, new_n23843_,
    new_n23844_, new_n23845_, new_n23846_, new_n23847_, new_n23848_,
    new_n23849_, new_n23850_, new_n23851_, new_n23852_, new_n23853_,
    new_n23854_, new_n23855_, new_n23856_, new_n23857_, new_n23858_,
    new_n23859_, new_n23860_, new_n23861_, new_n23862_, new_n23863_,
    new_n23864_, new_n23865_, new_n23866_, new_n23867_, new_n23868_,
    new_n23869_, new_n23870_, new_n23871_, new_n23872_, new_n23873_,
    new_n23874_, new_n23875_, new_n23876_, new_n23877_, new_n23878_,
    new_n23879_, new_n23880_, new_n23881_, new_n23882_, new_n23883_,
    new_n23884_, new_n23885_, new_n23886_, new_n23887_, new_n23888_,
    new_n23889_, new_n23890_, new_n23891_, new_n23892_, new_n23893_,
    new_n23894_, new_n23895_, new_n23896_, new_n23897_, new_n23898_,
    new_n23899_, new_n23900_, new_n23901_, new_n23902_, new_n23903_,
    new_n23904_, new_n23905_, new_n23906_, new_n23907_, new_n23908_,
    new_n23909_, new_n23910_, new_n23911_, new_n23912_, new_n23913_,
    new_n23914_, new_n23915_, new_n23916_, new_n23917_, new_n23918_,
    new_n23919_, new_n23920_, new_n23921_, new_n23922_, new_n23923_,
    new_n23924_, new_n23925_, new_n23926_, new_n23927_, new_n23928_,
    new_n23929_, new_n23930_, new_n23931_, new_n23932_, new_n23933_,
    new_n23934_, new_n23935_, new_n23936_, new_n23937_, new_n23938_,
    new_n23939_, new_n23940_, new_n23941_, new_n23942_, new_n23943_,
    new_n23944_, new_n23945_, new_n23946_, new_n23947_, new_n23948_,
    new_n23949_, new_n23950_, new_n23951_, new_n23952_, new_n23953_,
    new_n23954_, new_n23955_, new_n23956_, new_n23957_, new_n23958_,
    new_n23959_, new_n23960_, new_n23961_, new_n23962_, new_n23963_,
    new_n23964_, new_n23965_, new_n23966_, new_n23967_, new_n23968_,
    new_n23969_, new_n23970_, new_n23971_, new_n23972_, new_n23973_,
    new_n23974_, new_n23975_, new_n23976_, new_n23977_, new_n23978_,
    new_n23979_, new_n23980_, new_n23981_, new_n23982_, new_n23983_,
    new_n23984_, new_n23985_, new_n23986_, new_n23987_, new_n23988_,
    new_n23989_, new_n23990_, new_n23992_, new_n23993_, new_n23994_,
    new_n23995_, new_n23996_, new_n23997_, new_n23998_, new_n23999_,
    new_n24000_, new_n24001_, new_n24002_, new_n24003_, new_n24004_,
    new_n24005_, new_n24006_, new_n24007_, new_n24008_, new_n24009_,
    new_n24010_, new_n24011_, new_n24012_, new_n24013_, new_n24014_,
    new_n24015_, new_n24016_, new_n24017_, new_n24018_, new_n24019_,
    new_n24020_, new_n24021_, new_n24022_, new_n24023_, new_n24024_,
    new_n24025_, new_n24026_, new_n24027_, new_n24028_, new_n24029_,
    new_n24030_, new_n24031_, new_n24032_, new_n24033_, new_n24034_,
    new_n24035_, new_n24036_, new_n24037_, new_n24038_, new_n24039_,
    new_n24040_, new_n24041_, new_n24042_, new_n24043_, new_n24044_,
    new_n24045_, new_n24046_, new_n24047_, new_n24048_, new_n24049_,
    new_n24050_, new_n24051_, new_n24052_, new_n24053_, new_n24054_,
    new_n24055_, new_n24056_, new_n24057_, new_n24058_, new_n24059_,
    new_n24060_, new_n24061_, new_n24062_, new_n24063_, new_n24064_,
    new_n24065_, new_n24066_, new_n24067_, new_n24068_, new_n24069_,
    new_n24070_, new_n24071_, new_n24072_, new_n24073_, new_n24074_,
    new_n24075_, new_n24076_, new_n24077_, new_n24078_, new_n24079_,
    new_n24080_, new_n24081_, new_n24082_, new_n24083_, new_n24084_,
    new_n24085_, new_n24086_, new_n24087_, new_n24088_, new_n24089_,
    new_n24090_, new_n24091_, new_n24092_, new_n24093_, new_n24094_,
    new_n24095_, new_n24096_, new_n24097_, new_n24098_, new_n24099_,
    new_n24100_, new_n24101_, new_n24102_, new_n24103_, new_n24104_,
    new_n24105_, new_n24106_, new_n24107_, new_n24108_, new_n24109_,
    new_n24110_, new_n24111_, new_n24112_, new_n24113_, new_n24114_,
    new_n24115_, new_n24116_, new_n24117_, new_n24118_, new_n24119_,
    new_n24120_, new_n24121_, new_n24122_, new_n24123_, new_n24124_,
    new_n24125_, new_n24126_, new_n24127_, new_n24128_, new_n24129_,
    new_n24130_, new_n24131_, new_n24132_, new_n24133_, new_n24134_,
    new_n24135_, new_n24136_, new_n24137_, new_n24138_, new_n24139_,
    new_n24140_, new_n24141_, new_n24142_, new_n24143_, new_n24144_,
    new_n24145_, new_n24146_, new_n24147_, new_n24148_, new_n24149_,
    new_n24150_, new_n24151_, new_n24152_, new_n24153_, new_n24154_,
    new_n24155_, new_n24156_, new_n24157_, new_n24158_, new_n24159_,
    new_n24160_, new_n24161_, new_n24162_, new_n24163_, new_n24164_,
    new_n24165_, new_n24166_, new_n24167_, new_n24168_, new_n24169_,
    new_n24170_, new_n24171_, new_n24172_, new_n24173_, new_n24174_,
    new_n24175_, new_n24176_, new_n24177_, new_n24178_, new_n24179_,
    new_n24180_, new_n24181_, new_n24182_, new_n24183_, new_n24184_,
    new_n24185_, new_n24186_, new_n24187_, new_n24188_, new_n24189_,
    new_n24190_, new_n24191_, new_n24192_, new_n24193_, new_n24194_,
    new_n24195_, new_n24196_, new_n24197_, new_n24198_, new_n24199_,
    new_n24200_, new_n24201_, new_n24202_, new_n24203_, new_n24204_,
    new_n24205_, new_n24206_, new_n24207_, new_n24208_, new_n24209_,
    new_n24210_, new_n24211_, new_n24212_, new_n24213_, new_n24214_,
    new_n24215_, new_n24216_, new_n24217_, new_n24218_, new_n24219_,
    new_n24220_, new_n24221_, new_n24222_, new_n24223_, new_n24224_,
    new_n24225_, new_n24226_, new_n24227_, new_n24228_, new_n24229_,
    new_n24230_, new_n24231_, new_n24232_, new_n24233_, new_n24234_,
    new_n24235_, new_n24236_, new_n24237_, new_n24238_, new_n24239_,
    new_n24240_, new_n24241_, new_n24242_, new_n24243_, new_n24244_,
    new_n24245_, new_n24246_, new_n24247_, new_n24248_, new_n24249_,
    new_n24250_, new_n24251_, new_n24252_, new_n24253_, new_n24254_,
    new_n24255_, new_n24256_, new_n24257_, new_n24258_, new_n24259_,
    new_n24260_, new_n24261_, new_n24262_, new_n24263_, new_n24264_,
    new_n24265_, new_n24266_, new_n24267_, new_n24268_, new_n24269_,
    new_n24270_, new_n24271_, new_n24272_, new_n24273_, new_n24274_,
    new_n24275_, new_n24276_, new_n24277_, new_n24278_, new_n24279_,
    new_n24280_, new_n24281_, new_n24282_, new_n24283_, new_n24284_,
    new_n24285_, new_n24286_, new_n24287_, new_n24288_, new_n24289_,
    new_n24290_, new_n24291_, new_n24292_, new_n24293_, new_n24294_,
    new_n24295_, new_n24296_, new_n24297_, new_n24298_, new_n24299_,
    new_n24300_, new_n24301_, new_n24302_, new_n24303_, new_n24304_,
    new_n24305_, new_n24306_, new_n24307_, new_n24308_, new_n24309_,
    new_n24310_, new_n24311_, new_n24312_, new_n24313_, new_n24314_,
    new_n24315_, new_n24316_, new_n24317_, new_n24318_, new_n24319_,
    new_n24320_, new_n24321_, new_n24322_, new_n24323_, new_n24324_,
    new_n24325_, new_n24326_, new_n24327_, new_n24328_, new_n24329_,
    new_n24330_, new_n24331_, new_n24332_, new_n24333_, new_n24334_,
    new_n24335_, new_n24336_, new_n24337_, new_n24338_, new_n24339_,
    new_n24340_, new_n24341_, new_n24342_, new_n24343_, new_n24344_,
    new_n24345_, new_n24346_, new_n24347_, new_n24348_, new_n24349_,
    new_n24350_, new_n24351_, new_n24352_, new_n24353_, new_n24354_,
    new_n24355_, new_n24356_, new_n24357_, new_n24358_, new_n24359_,
    new_n24360_, new_n24361_, new_n24362_, new_n24363_, new_n24364_,
    new_n24365_, new_n24366_, new_n24367_, new_n24368_, new_n24369_,
    new_n24370_, new_n24371_, new_n24372_, new_n24373_, new_n24374_,
    new_n24375_, new_n24376_, new_n24377_, new_n24378_, new_n24379_,
    new_n24380_, new_n24381_, new_n24382_, new_n24383_, new_n24384_,
    new_n24385_, new_n24386_, new_n24387_, new_n24388_, new_n24389_,
    new_n24390_, new_n24391_, new_n24392_, new_n24393_, new_n24394_,
    new_n24395_, new_n24396_, new_n24397_, new_n24398_, new_n24399_,
    new_n24400_, new_n24401_, new_n24402_, new_n24403_, new_n24404_,
    new_n24405_, new_n24406_, new_n24407_, new_n24408_, new_n24409_,
    new_n24410_, new_n24411_, new_n24412_, new_n24413_, new_n24414_,
    new_n24415_, new_n24416_, new_n24417_, new_n24418_, new_n24419_,
    new_n24420_, new_n24421_, new_n24422_, new_n24423_, new_n24424_,
    new_n24425_, new_n24426_, new_n24427_, new_n24428_, new_n24429_,
    new_n24430_, new_n24431_, new_n24432_, new_n24433_, new_n24434_,
    new_n24435_, new_n24436_, new_n24437_, new_n24438_, new_n24439_,
    new_n24440_, new_n24441_, new_n24442_, new_n24443_, new_n24444_,
    new_n24445_, new_n24446_, new_n24447_, new_n24448_, new_n24449_,
    new_n24450_, new_n24451_, new_n24452_, new_n24453_, new_n24454_,
    new_n24455_, new_n24456_, new_n24457_, new_n24458_, new_n24459_,
    new_n24460_, new_n24461_, new_n24462_, new_n24463_, new_n24464_,
    new_n24465_, new_n24466_, new_n24467_, new_n24468_, new_n24469_,
    new_n24470_, new_n24471_, new_n24472_, new_n24473_, new_n24474_,
    new_n24475_, new_n24476_, new_n24477_, new_n24478_, new_n24479_,
    new_n24480_, new_n24481_, new_n24482_, new_n24483_, new_n24484_,
    new_n24485_, new_n24486_, new_n24487_, new_n24488_, new_n24489_,
    new_n24490_, new_n24491_, new_n24492_, new_n24493_, new_n24494_,
    new_n24495_, new_n24496_, new_n24497_, new_n24498_, new_n24499_,
    new_n24500_, new_n24501_, new_n24502_, new_n24503_, new_n24504_,
    new_n24505_, new_n24506_, new_n24507_, new_n24508_, new_n24509_,
    new_n24510_, new_n24511_, new_n24512_, new_n24513_, new_n24514_,
    new_n24515_, new_n24516_, new_n24517_, new_n24518_, new_n24519_,
    new_n24520_, new_n24521_, new_n24522_, new_n24523_, new_n24524_,
    new_n24525_, new_n24526_, new_n24527_, new_n24528_, new_n24529_,
    new_n24530_, new_n24531_, new_n24532_, new_n24533_, new_n24534_,
    new_n24535_, new_n24536_, new_n24537_, new_n24538_, new_n24539_,
    new_n24540_, new_n24541_, new_n24542_, new_n24543_, new_n24544_,
    new_n24545_, new_n24546_, new_n24547_, new_n24548_, new_n24549_,
    new_n24550_, new_n24551_, new_n24552_, new_n24553_, new_n24554_,
    new_n24555_, new_n24556_, new_n24557_, new_n24558_, new_n24559_,
    new_n24560_, new_n24561_, new_n24562_, new_n24563_, new_n24564_,
    new_n24565_, new_n24566_, new_n24567_, new_n24568_, new_n24569_,
    new_n24570_, new_n24571_, new_n24572_, new_n24573_, new_n24574_,
    new_n24575_, new_n24576_, new_n24577_, new_n24578_, new_n24579_,
    new_n24580_, new_n24581_, new_n24582_, new_n24583_, new_n24584_,
    new_n24585_, new_n24586_, new_n24587_, new_n24588_, new_n24589_,
    new_n24590_, new_n24591_, new_n24592_, new_n24593_;
  NAND2_X1   g00000(.A1(\a[126] ), .A2(\a[127] ), .ZN(new_n193_));
  OAI21_X1   g00001(.A1(\a[124] ), .A2(\a[127] ), .B(\a[125] ), .ZN(new_n194_));
  NAND2_X1   g00002(.A1(new_n194_), .A2(new_n193_), .ZN(\asqrt[62] ));
  INV_X1     g00003(.I(\asqrt[62] ), .ZN(new_n196_));
  OAI21_X1   g00004(.A1(\a[125] ), .A2(\a[126] ), .B(\a[127] ), .ZN(new_n197_));
  INV_X1     g00005(.I(new_n197_), .ZN(new_n198_));
  NOR3_X1    g00006(.A1(\a[122] ), .A2(\a[123] ), .A3(\a[124] ), .ZN(new_n199_));
  INV_X1     g00007(.I(\a[124] ), .ZN(new_n200_));
  INV_X1     g00008(.I(\a[125] ), .ZN(new_n201_));
  INV_X1     g00009(.I(\a[126] ), .ZN(new_n202_));
  NOR4_X1    g00010(.A1(new_n200_), .A2(new_n201_), .A3(new_n202_), .A4(\a[127] ), .ZN(new_n203_));
  OAI21_X1   g00011(.A1(new_n203_), .A2(new_n199_), .B(new_n198_), .ZN(new_n204_));
  INV_X1     g00012(.I(new_n199_), .ZN(new_n205_));
  NOR2_X1    g00013(.A1(new_n193_), .A2(\a[125] ), .ZN(new_n206_));
  AOI21_X1   g00014(.A1(\a[126] ), .A2(\a[127] ), .B(new_n201_), .ZN(new_n207_));
  OAI21_X1   g00015(.A1(new_n207_), .A2(new_n206_), .B(\a[124] ), .ZN(new_n208_));
  OAI21_X1   g00016(.A1(new_n201_), .A2(new_n202_), .B(\a[124] ), .ZN(new_n209_));
  NOR3_X1    g00017(.A1(new_n201_), .A2(new_n202_), .A3(\a[124] ), .ZN(new_n210_));
  INV_X1     g00018(.I(\a[127] ), .ZN(new_n211_));
  NAND2_X1   g00019(.A1(new_n211_), .A2(\a[125] ), .ZN(new_n212_));
  NOR2_X1    g00020(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  AOI21_X1   g00021(.A1(new_n213_), .A2(new_n209_), .B(new_n198_), .ZN(new_n214_));
  AOI21_X1   g00022(.A1(new_n214_), .A2(new_n208_), .B(new_n205_), .ZN(new_n215_));
  NAND2_X1   g00023(.A1(new_n215_), .A2(new_n204_), .ZN(\asqrt[61] ));
  INV_X1     g00024(.I(\a[7] ), .ZN(new_n217_));
  NAND4_X1   g00025(.A1(new_n211_), .A2(\a[124] ), .A3(\a[125] ), .A4(\a[126] ), .ZN(new_n218_));
  AOI21_X1   g00026(.A1(new_n205_), .A2(new_n218_), .B(new_n197_), .ZN(new_n219_));
  NAND3_X1   g00027(.A1(new_n201_), .A2(\a[126] ), .A3(\a[127] ), .ZN(new_n220_));
  NAND2_X1   g00028(.A1(new_n193_), .A2(\a[125] ), .ZN(new_n221_));
  AOI21_X1   g00029(.A1(new_n221_), .A2(new_n220_), .B(new_n200_), .ZN(new_n222_));
  AOI21_X1   g00030(.A1(\a[125] ), .A2(\a[126] ), .B(new_n200_), .ZN(new_n223_));
  NAND3_X1   g00031(.A1(new_n200_), .A2(\a[125] ), .A3(\a[126] ), .ZN(new_n224_));
  NOR2_X1    g00032(.A1(new_n201_), .A2(\a[127] ), .ZN(new_n225_));
  NAND2_X1   g00033(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1   g00034(.A1(new_n226_), .A2(new_n223_), .B(new_n197_), .ZN(new_n227_));
  OAI21_X1   g00035(.A1(new_n227_), .A2(new_n222_), .B(new_n199_), .ZN(new_n228_));
  NOR2_X1    g00036(.A1(new_n228_), .A2(new_n219_), .ZN(new_n229_));
  INV_X1     g00037(.I(\a[115] ), .ZN(new_n230_));
  NOR2_X1    g00038(.A1(\a[126] ), .A2(\a[127] ), .ZN(new_n231_));
  INV_X1     g00039(.I(new_n231_), .ZN(\asqrt[63] ));
  NOR2_X1    g00040(.A1(\a[120] ), .A2(\a[121] ), .ZN(new_n233_));
  NOR2_X1    g00041(.A1(\a[122] ), .A2(\a[123] ), .ZN(new_n234_));
  NOR4_X1    g00042(.A1(new_n200_), .A2(new_n201_), .A3(new_n202_), .A4(\a[127] ), .ZN(new_n235_));
  INV_X1     g00043(.I(new_n234_), .ZN(new_n236_));
  NOR4_X1    g00044(.A1(new_n200_), .A2(new_n201_), .A3(\a[126] ), .A4(\a[127] ), .ZN(new_n237_));
  NOR4_X1    g00045(.A1(new_n228_), .A2(new_n200_), .A3(new_n236_), .A4(new_n219_), .ZN(new_n238_));
  NAND2_X1   g00046(.A1(new_n219_), .A2(new_n237_), .ZN(new_n239_));
  AOI21_X1   g00047(.A1(new_n239_), .A2(new_n200_), .B(new_n236_), .ZN(new_n240_));
  NOR2_X1    g00048(.A1(new_n229_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1    g00049(.A1(new_n241_), .A2(new_n238_), .ZN(new_n242_));
  NAND3_X1   g00050(.A1(new_n209_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n243_));
  NAND3_X1   g00051(.A1(new_n208_), .A2(new_n243_), .A3(new_n197_), .ZN(new_n244_));
  INV_X1     g00052(.I(\a[122] ), .ZN(new_n245_));
  NOR3_X1    g00053(.A1(new_n194_), .A2(new_n245_), .A3(new_n193_), .ZN(new_n246_));
  AOI21_X1   g00054(.A1(new_n244_), .A2(new_n199_), .B(new_n246_), .ZN(new_n247_));
  NOR3_X1    g00055(.A1(new_n247_), .A2(new_n196_), .A3(new_n204_), .ZN(new_n248_));
  NAND4_X1   g00056(.A1(new_n244_), .A2(new_n236_), .A3(new_n199_), .A4(new_n204_), .ZN(new_n249_));
  OAI21_X1   g00057(.A1(new_n228_), .A2(new_n234_), .B(new_n219_), .ZN(new_n250_));
  NAND2_X1   g00058(.A1(new_n250_), .A2(new_n249_), .ZN(new_n251_));
  NAND2_X1   g00059(.A1(new_n204_), .A2(\a[122] ), .ZN(new_n252_));
  INV_X1     g00060(.I(new_n233_), .ZN(new_n253_));
  NOR2_X1    g00061(.A1(new_n253_), .A2(new_n245_), .ZN(new_n254_));
  NAND4_X1   g00062(.A1(new_n244_), .A2(new_n252_), .A3(new_n199_), .A4(new_n254_), .ZN(new_n255_));
  NOR2_X1    g00063(.A1(new_n219_), .A2(new_n245_), .ZN(new_n256_));
  INV_X1     g00064(.I(new_n254_), .ZN(new_n257_));
  OAI21_X1   g00065(.A1(new_n228_), .A2(new_n257_), .B(new_n256_), .ZN(new_n258_));
  NAND2_X1   g00066(.A1(new_n258_), .A2(new_n255_), .ZN(new_n259_));
  AOI21_X1   g00067(.A1(new_n251_), .A2(new_n259_), .B(new_n248_), .ZN(new_n260_));
  INV_X1     g00068(.I(new_n243_), .ZN(new_n261_));
  NAND2_X1   g00069(.A1(new_n205_), .A2(new_n197_), .ZN(new_n262_));
  NOR2_X1    g00070(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1     g00071(.I(new_n263_), .ZN(new_n264_));
  NAND2_X1   g00072(.A1(new_n261_), .A2(new_n262_), .ZN(new_n265_));
  INV_X1     g00073(.I(new_n265_), .ZN(new_n266_));
  NAND2_X1   g00074(.A1(\asqrt[61] ), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1   g00075(.A1(new_n267_), .A2(new_n264_), .B(\asqrt[63] ), .ZN(new_n268_));
  AOI21_X1   g00076(.A1(new_n260_), .A2(new_n268_), .B(new_n242_), .ZN(new_n269_));
  NAND2_X1   g00077(.A1(new_n243_), .A2(new_n262_), .ZN(new_n270_));
  NAND2_X1   g00078(.A1(new_n270_), .A2(new_n222_), .ZN(new_n271_));
  XOR2_X1    g00079(.A1(new_n262_), .A2(new_n231_), .Z(new_n272_));
  NAND2_X1   g00080(.A1(new_n272_), .A2(new_n271_), .ZN(new_n273_));
  NOR3_X1    g00081(.A1(new_n260_), .A2(new_n242_), .A3(new_n273_), .ZN(new_n274_));
  NAND3_X1   g00082(.A1(new_n274_), .A2(new_n269_), .A3(new_n235_), .ZN(new_n275_));
  INV_X1     g00083(.I(new_n235_), .ZN(new_n276_));
  NAND3_X1   g00084(.A1(new_n273_), .A2(\asqrt[61] ), .A3(new_n276_), .ZN(new_n277_));
  INV_X1     g00085(.I(new_n277_), .ZN(new_n278_));
  OAI21_X1   g00086(.A1(new_n260_), .A2(new_n242_), .B(new_n278_), .ZN(new_n279_));
  OAI21_X1   g00087(.A1(new_n279_), .A2(new_n269_), .B(new_n245_), .ZN(new_n280_));
  NAND3_X1   g00088(.A1(new_n280_), .A2(new_n275_), .A3(new_n233_), .ZN(new_n281_));
  INV_X1     g00089(.I(new_n238_), .ZN(new_n282_));
  INV_X1     g00090(.I(new_n240_), .ZN(new_n283_));
  NAND2_X1   g00091(.A1(\asqrt[61] ), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1   g00092(.A1(new_n284_), .A2(new_n282_), .ZN(new_n285_));
  INV_X1     g00093(.I(new_n246_), .ZN(new_n286_));
  AOI21_X1   g00094(.A1(new_n228_), .A2(new_n286_), .B(new_n204_), .ZN(new_n287_));
  NAND2_X1   g00095(.A1(new_n287_), .A2(\asqrt[62] ), .ZN(new_n288_));
  NOR3_X1    g00096(.A1(new_n228_), .A2(new_n234_), .A3(new_n219_), .ZN(new_n289_));
  AOI21_X1   g00097(.A1(new_n215_), .A2(new_n236_), .B(new_n204_), .ZN(new_n290_));
  NOR2_X1    g00098(.A1(new_n290_), .A2(new_n289_), .ZN(new_n291_));
  NOR3_X1    g00099(.A1(new_n228_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n292_));
  AOI21_X1   g00100(.A1(new_n215_), .A2(new_n254_), .B(new_n252_), .ZN(new_n293_));
  NOR2_X1    g00101(.A1(new_n293_), .A2(new_n292_), .ZN(new_n294_));
  OAI21_X1   g00102(.A1(new_n291_), .A2(new_n294_), .B(new_n288_), .ZN(new_n295_));
  AOI21_X1   g00103(.A1(new_n215_), .A2(new_n204_), .B(new_n265_), .ZN(new_n296_));
  OAI21_X1   g00104(.A1(new_n296_), .A2(new_n263_), .B(new_n231_), .ZN(new_n297_));
  OAI21_X1   g00105(.A1(new_n295_), .A2(new_n297_), .B(new_n285_), .ZN(new_n298_));
  INV_X1     g00106(.I(new_n273_), .ZN(new_n299_));
  NAND3_X1   g00107(.A1(new_n295_), .A2(new_n285_), .A3(new_n299_), .ZN(new_n300_));
  NOR3_X1    g00108(.A1(new_n298_), .A2(new_n300_), .A3(new_n276_), .ZN(\asqrt[60] ));
  AOI21_X1   g00109(.A1(new_n295_), .A2(new_n285_), .B(new_n277_), .ZN(new_n302_));
  AOI21_X1   g00110(.A1(new_n302_), .A2(new_n298_), .B(\a[122] ), .ZN(new_n303_));
  OAI21_X1   g00111(.A1(new_n253_), .A2(new_n303_), .B(\asqrt[60] ), .ZN(new_n304_));
  AOI21_X1   g00112(.A1(new_n304_), .A2(new_n281_), .B(new_n196_), .ZN(new_n305_));
  NOR3_X1    g00113(.A1(new_n303_), .A2(\asqrt[60] ), .A3(new_n253_), .ZN(new_n306_));
  AOI21_X1   g00114(.A1(new_n233_), .A2(new_n280_), .B(new_n275_), .ZN(new_n307_));
  NOR3_X1    g00115(.A1(new_n306_), .A2(new_n307_), .A3(\asqrt[62] ), .ZN(new_n308_));
  INV_X1     g00116(.I(\a[121] ), .ZN(new_n309_));
  NOR2_X1    g00117(.A1(\a[118] ), .A2(\a[119] ), .ZN(new_n310_));
  INV_X1     g00118(.I(new_n310_), .ZN(new_n311_));
  NOR2_X1    g00119(.A1(new_n311_), .A2(\a[120] ), .ZN(new_n312_));
  NOR4_X1    g00120(.A1(new_n263_), .A2(new_n219_), .A3(new_n222_), .A4(new_n312_), .ZN(new_n313_));
  XOR2_X1    g00121(.A1(new_n313_), .A2(new_n309_), .Z(new_n314_));
  INV_X1     g00122(.I(new_n314_), .ZN(new_n315_));
  NAND4_X1   g00123(.A1(new_n274_), .A2(new_n269_), .A3(\a[121] ), .A4(new_n235_), .ZN(new_n316_));
  NOR2_X1    g00124(.A1(new_n314_), .A2(\a[120] ), .ZN(new_n317_));
  INV_X1     g00125(.I(new_n317_), .ZN(new_n318_));
  AOI21_X1   g00126(.A1(new_n316_), .A2(new_n318_), .B(new_n315_), .ZN(new_n319_));
  INV_X1     g00127(.I(\a[120] ), .ZN(new_n320_));
  NOR4_X1    g00128(.A1(new_n298_), .A2(new_n300_), .A3(new_n309_), .A4(new_n276_), .ZN(new_n321_));
  NOR3_X1    g00129(.A1(new_n321_), .A2(new_n320_), .A3(new_n314_), .ZN(new_n322_));
  NOR2_X1    g00130(.A1(new_n322_), .A2(new_n319_), .ZN(new_n323_));
  NOR3_X1    g00131(.A1(new_n275_), .A2(new_n320_), .A3(new_n229_), .ZN(new_n324_));
  NOR3_X1    g00132(.A1(\asqrt[60] ), .A2(\a[120] ), .A3(new_n229_), .ZN(new_n325_));
  OAI21_X1   g00133(.A1(new_n325_), .A2(new_n324_), .B(new_n310_), .ZN(new_n326_));
  NOR3_X1    g00134(.A1(new_n308_), .A2(new_n323_), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1   g00135(.A1(new_n294_), .A2(\asqrt[62] ), .B(new_n287_), .ZN(new_n328_));
  NAND4_X1   g00136(.A1(new_n274_), .A2(new_n269_), .A3(new_n235_), .A4(new_n328_), .ZN(new_n329_));
  INV_X1     g00137(.I(new_n328_), .ZN(new_n330_));
  NOR2_X1    g00138(.A1(new_n330_), .A2(new_n291_), .ZN(new_n331_));
  AOI22_X1   g00139(.A1(\asqrt[60] ), .A2(new_n331_), .B1(new_n329_), .B2(new_n291_), .ZN(new_n332_));
  AOI21_X1   g00140(.A1(new_n332_), .A2(new_n285_), .B(new_n260_), .ZN(new_n333_));
  NAND2_X1   g00141(.A1(new_n333_), .A2(\asqrt[60] ), .ZN(new_n334_));
  NOR3_X1    g00142(.A1(new_n327_), .A2(new_n334_), .A3(new_n305_), .ZN(new_n335_));
  NAND2_X1   g00143(.A1(new_n304_), .A2(new_n281_), .ZN(new_n336_));
  NOR4_X1    g00144(.A1(new_n298_), .A2(new_n300_), .A3(new_n276_), .A4(new_n330_), .ZN(new_n337_));
  INV_X1     g00145(.I(new_n331_), .ZN(new_n338_));
  OAI22_X1   g00146(.A1(new_n337_), .A2(new_n251_), .B1(new_n338_), .B2(new_n275_), .ZN(new_n339_));
  AOI22_X1   g00147(.A1(new_n249_), .A2(new_n250_), .B1(new_n258_), .B2(new_n255_), .ZN(new_n340_));
  NOR3_X1    g00148(.A1(new_n340_), .A2(new_n248_), .A3(new_n297_), .ZN(new_n341_));
  NOR4_X1    g00149(.A1(new_n341_), .A2(new_n242_), .A3(new_n260_), .A4(new_n273_), .ZN(new_n342_));
  NAND4_X1   g00150(.A1(new_n342_), .A2(\a[120] ), .A3(\asqrt[61] ), .A4(new_n235_), .ZN(new_n343_));
  NAND3_X1   g00151(.A1(new_n275_), .A2(new_n320_), .A3(\asqrt[61] ), .ZN(new_n344_));
  AOI21_X1   g00152(.A1(new_n344_), .A2(new_n343_), .B(new_n311_), .ZN(new_n345_));
  NOR3_X1    g00153(.A1(new_n345_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n346_));
  NAND4_X1   g00154(.A1(new_n346_), .A2(new_n196_), .A3(new_n336_), .A4(new_n339_), .ZN(new_n347_));
  AOI21_X1   g00155(.A1(new_n242_), .A2(new_n260_), .B(new_n275_), .ZN(new_n348_));
  XOR2_X1    g00156(.A1(new_n260_), .A2(\asqrt[63] ), .Z(new_n349_));
  NOR2_X1    g00157(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1     g00158(.I(new_n350_), .ZN(new_n351_));
  NOR4_X1    g00159(.A1(new_n335_), .A2(\asqrt[63] ), .A3(new_n347_), .A4(new_n351_), .ZN(new_n352_));
  NOR4_X1    g00160(.A1(new_n200_), .A2(new_n201_), .A3(new_n202_), .A4(\a[127] ), .ZN(new_n353_));
  NAND4_X1   g00161(.A1(new_n342_), .A2(new_n234_), .A3(\asqrt[61] ), .A4(new_n353_), .ZN(new_n354_));
  NOR2_X1    g00162(.A1(new_n354_), .A2(new_n291_), .ZN(new_n355_));
  XOR2_X1    g00163(.A1(new_n355_), .A2(new_n330_), .Z(new_n356_));
  NOR2_X1    g00164(.A1(new_n356_), .A2(new_n275_), .ZN(new_n357_));
  NAND2_X1   g00165(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1     g00166(.I(new_n358_), .ZN(new_n359_));
  NAND2_X1   g00167(.A1(new_n323_), .A2(new_n326_), .ZN(new_n360_));
  NAND2_X1   g00168(.A1(new_n360_), .A2(\asqrt[62] ), .ZN(new_n361_));
  NOR2_X1    g00169(.A1(new_n306_), .A2(new_n307_), .ZN(new_n362_));
  OAI21_X1   g00170(.A1(new_n321_), .A2(new_n317_), .B(new_n314_), .ZN(new_n363_));
  NAND3_X1   g00171(.A1(new_n316_), .A2(\a[120] ), .A3(new_n315_), .ZN(new_n364_));
  NAND2_X1   g00172(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NOR4_X1    g00173(.A1(new_n362_), .A2(new_n365_), .A3(new_n345_), .A4(\asqrt[62] ), .ZN(new_n366_));
  INV_X1     g00174(.I(new_n366_), .ZN(new_n367_));
  OAI21_X1   g00175(.A1(new_n306_), .A2(new_n307_), .B(\asqrt[62] ), .ZN(new_n368_));
  NAND3_X1   g00176(.A1(new_n304_), .A2(new_n281_), .A3(new_n196_), .ZN(new_n369_));
  NAND3_X1   g00177(.A1(new_n369_), .A2(new_n365_), .A3(new_n345_), .ZN(new_n370_));
  OAI21_X1   g00178(.A1(new_n339_), .A2(new_n242_), .B(new_n295_), .ZN(new_n371_));
  NOR2_X1    g00179(.A1(new_n371_), .A2(new_n275_), .ZN(new_n372_));
  NAND3_X1   g00180(.A1(new_n372_), .A2(new_n370_), .A3(new_n368_), .ZN(new_n373_));
  NOR2_X1    g00181(.A1(new_n347_), .A2(new_n351_), .ZN(new_n374_));
  INV_X1     g00182(.I(new_n354_), .ZN(new_n375_));
  NAND4_X1   g00183(.A1(new_n374_), .A2(new_n231_), .A3(new_n373_), .A4(new_n375_), .ZN(new_n376_));
  NOR3_X1    g00184(.A1(new_n376_), .A2(new_n361_), .A3(new_n367_), .ZN(new_n377_));
  NOR2_X1    g00185(.A1(new_n360_), .A2(\asqrt[62] ), .ZN(new_n378_));
  NOR2_X1    g00186(.A1(new_n378_), .A2(new_n336_), .ZN(new_n379_));
  AOI21_X1   g00187(.A1(new_n376_), .A2(new_n379_), .B(new_n361_), .ZN(new_n380_));
  NOR2_X1    g00188(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1   g00189(.A1(new_n365_), .A2(new_n345_), .ZN(new_n382_));
  OAI21_X1   g00190(.A1(new_n382_), .A2(new_n308_), .B(new_n368_), .ZN(new_n383_));
  OAI21_X1   g00191(.A1(new_n383_), .A2(new_n334_), .B(new_n231_), .ZN(new_n384_));
  OAI21_X1   g00192(.A1(new_n346_), .A2(new_n196_), .B(new_n332_), .ZN(new_n385_));
  NAND3_X1   g00193(.A1(new_n385_), .A2(new_n366_), .A3(new_n350_), .ZN(new_n386_));
  NOR3_X1    g00194(.A1(new_n384_), .A2(new_n386_), .A3(new_n354_), .ZN(\asqrt[59] ));
  NOR2_X1    g00195(.A1(new_n275_), .A2(\a[120] ), .ZN(new_n388_));
  OAI22_X1   g00196(.A1(new_n388_), .A2(\a[121] ), .B1(\a[120] ), .B2(new_n316_), .ZN(new_n389_));
  NAND2_X1   g00197(.A1(new_n345_), .A2(new_n313_), .ZN(new_n390_));
  AOI21_X1   g00198(.A1(new_n390_), .A2(new_n320_), .B(new_n275_), .ZN(new_n391_));
  AOI21_X1   g00199(.A1(\asqrt[59] ), .A2(new_n391_), .B(new_n389_), .ZN(new_n392_));
  NAND2_X1   g00200(.A1(new_n391_), .A2(new_n389_), .ZN(new_n393_));
  NOR2_X1    g00201(.A1(new_n376_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1    g00202(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1    g00203(.A1(new_n395_), .A2(new_n196_), .ZN(new_n396_));
  INV_X1     g00204(.I(new_n396_), .ZN(new_n397_));
  INV_X1     g00205(.I(\a[119] ), .ZN(new_n398_));
  NOR2_X1    g00206(.A1(\a[116] ), .A2(\a[117] ), .ZN(new_n399_));
  INV_X1     g00207(.I(new_n399_), .ZN(new_n400_));
  NOR2_X1    g00208(.A1(new_n400_), .A2(\a[118] ), .ZN(new_n401_));
  NOR4_X1    g00209(.A1(new_n298_), .A2(new_n300_), .A3(new_n235_), .A4(new_n401_), .ZN(new_n402_));
  XOR2_X1    g00210(.A1(new_n402_), .A2(new_n398_), .Z(new_n403_));
  NOR4_X1    g00211(.A1(new_n384_), .A2(new_n386_), .A3(new_n398_), .A4(new_n354_), .ZN(new_n404_));
  NOR2_X1    g00212(.A1(new_n403_), .A2(\a[118] ), .ZN(new_n405_));
  OAI21_X1   g00213(.A1(new_n404_), .A2(new_n405_), .B(new_n403_), .ZN(new_n406_));
  INV_X1     g00214(.I(new_n403_), .ZN(new_n407_));
  NOR2_X1    g00215(.A1(new_n323_), .A2(new_n326_), .ZN(new_n408_));
  AOI21_X1   g00216(.A1(new_n408_), .A2(new_n369_), .B(new_n305_), .ZN(new_n409_));
  AOI21_X1   g00217(.A1(new_n409_), .A2(new_n372_), .B(\asqrt[63] ), .ZN(new_n410_));
  NAND4_X1   g00218(.A1(new_n410_), .A2(\a[119] ), .A3(new_n374_), .A4(new_n375_), .ZN(new_n411_));
  NAND3_X1   g00219(.A1(new_n411_), .A2(\a[118] ), .A3(new_n407_), .ZN(new_n412_));
  NAND2_X1   g00220(.A1(new_n412_), .A2(new_n406_), .ZN(new_n413_));
  NAND4_X1   g00221(.A1(new_n352_), .A2(\a[118] ), .A3(\asqrt[60] ), .A4(new_n375_), .ZN(new_n414_));
  INV_X1     g00222(.I(\a[118] ), .ZN(new_n415_));
  NAND3_X1   g00223(.A1(new_n376_), .A2(new_n415_), .A3(\asqrt[60] ), .ZN(new_n416_));
  AOI21_X1   g00224(.A1(new_n416_), .A2(new_n414_), .B(new_n400_), .ZN(new_n417_));
  NOR2_X1    g00225(.A1(new_n375_), .A2(new_n275_), .ZN(new_n418_));
  NAND3_X1   g00226(.A1(new_n347_), .A2(new_n351_), .A3(new_n418_), .ZN(new_n419_));
  OAI21_X1   g00227(.A1(new_n410_), .A2(new_n419_), .B(new_n320_), .ZN(new_n420_));
  NAND3_X1   g00228(.A1(new_n420_), .A2(new_n376_), .A3(new_n310_), .ZN(new_n421_));
  NAND2_X1   g00229(.A1(new_n351_), .A2(new_n418_), .ZN(new_n422_));
  AOI21_X1   g00230(.A1(new_n385_), .A2(new_n366_), .B(new_n422_), .ZN(new_n423_));
  AOI21_X1   g00231(.A1(new_n384_), .A2(new_n423_), .B(\a[120] ), .ZN(new_n424_));
  OAI21_X1   g00232(.A1(new_n311_), .A2(new_n424_), .B(\asqrt[59] ), .ZN(new_n425_));
  NAND3_X1   g00233(.A1(new_n425_), .A2(new_n421_), .A3(new_n229_), .ZN(new_n426_));
  OAI21_X1   g00234(.A1(new_n417_), .A2(new_n426_), .B(new_n413_), .ZN(new_n427_));
  NOR4_X1    g00235(.A1(new_n360_), .A2(\asqrt[62] ), .A3(new_n362_), .A4(new_n332_), .ZN(new_n428_));
  NAND4_X1   g00236(.A1(new_n373_), .A2(new_n428_), .A3(new_n231_), .A4(new_n350_), .ZN(new_n429_));
  NOR4_X1    g00237(.A1(new_n429_), .A2(new_n415_), .A3(new_n275_), .A4(new_n354_), .ZN(new_n430_));
  NOR3_X1    g00238(.A1(\asqrt[59] ), .A2(\a[118] ), .A3(new_n275_), .ZN(new_n431_));
  OAI21_X1   g00239(.A1(new_n431_), .A2(new_n430_), .B(new_n399_), .ZN(new_n432_));
  NAND3_X1   g00240(.A1(new_n432_), .A2(new_n406_), .A3(new_n412_), .ZN(new_n433_));
  NOR3_X1    g00241(.A1(new_n392_), .A2(new_n394_), .A3(\asqrt[62] ), .ZN(new_n434_));
  INV_X1     g00242(.I(new_n434_), .ZN(new_n435_));
  NAND3_X1   g00243(.A1(new_n433_), .A2(\asqrt[61] ), .A3(new_n435_), .ZN(new_n436_));
  OAI21_X1   g00244(.A1(new_n436_), .A2(new_n427_), .B(new_n397_), .ZN(new_n437_));
  NOR3_X1    g00245(.A1(\asqrt[59] ), .A2(new_n339_), .A3(new_n428_), .ZN(new_n438_));
  OAI21_X1   g00246(.A1(new_n438_), .A2(new_n409_), .B(new_n231_), .ZN(new_n439_));
  OAI21_X1   g00247(.A1(new_n437_), .A2(new_n439_), .B(new_n381_), .ZN(new_n440_));
  INV_X1     g00248(.I(new_n381_), .ZN(new_n441_));
  OAI21_X1   g00249(.A1(new_n413_), .A2(new_n417_), .B(\asqrt[61] ), .ZN(new_n442_));
  NAND2_X1   g00250(.A1(new_n427_), .A2(new_n442_), .ZN(new_n443_));
  NOR4_X1    g00251(.A1(new_n443_), .A2(\asqrt[62] ), .A3(new_n441_), .A4(new_n395_), .ZN(new_n444_));
  OAI21_X1   g00252(.A1(new_n376_), .A2(new_n409_), .B(new_n332_), .ZN(new_n445_));
  NOR2_X1    g00253(.A1(new_n428_), .A2(new_n231_), .ZN(new_n446_));
  NAND2_X1   g00254(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1     g00255(.I(new_n447_), .ZN(new_n448_));
  NAND2_X1   g00256(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1    g00257(.A1(\a[112] ), .A2(\a[113] ), .ZN(new_n450_));
  INV_X1     g00258(.I(new_n450_), .ZN(new_n451_));
  NOR2_X1    g00259(.A1(new_n451_), .A2(\a[114] ), .ZN(new_n452_));
  NOR4_X1    g00260(.A1(new_n449_), .A2(new_n359_), .A3(new_n440_), .A4(new_n452_), .ZN(new_n453_));
  XOR2_X1    g00261(.A1(new_n453_), .A2(new_n230_), .Z(new_n454_));
  INV_X1     g00262(.I(new_n405_), .ZN(new_n455_));
  AOI21_X1   g00263(.A1(new_n411_), .A2(new_n455_), .B(new_n407_), .ZN(new_n456_));
  NOR3_X1    g00264(.A1(new_n404_), .A2(new_n415_), .A3(new_n403_), .ZN(new_n457_));
  NOR2_X1    g00265(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NOR3_X1    g00266(.A1(new_n424_), .A2(\asqrt[59] ), .A3(new_n311_), .ZN(new_n459_));
  AOI21_X1   g00267(.A1(new_n420_), .A2(new_n310_), .B(new_n376_), .ZN(new_n460_));
  NOR3_X1    g00268(.A1(new_n460_), .A2(new_n459_), .A3(\asqrt[61] ), .ZN(new_n461_));
  AOI21_X1   g00269(.A1(new_n461_), .A2(new_n432_), .B(new_n458_), .ZN(new_n462_));
  AOI21_X1   g00270(.A1(new_n458_), .A2(new_n432_), .B(new_n229_), .ZN(new_n463_));
  NOR2_X1    g00271(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NOR2_X1    g00272(.A1(new_n464_), .A2(new_n196_), .ZN(new_n465_));
  INV_X1     g00273(.I(new_n395_), .ZN(new_n466_));
  NAND4_X1   g00274(.A1(new_n427_), .A2(new_n196_), .A3(new_n442_), .A4(new_n466_), .ZN(new_n467_));
  INV_X1     g00275(.I(new_n467_), .ZN(new_n468_));
  NAND4_X1   g00276(.A1(new_n464_), .A2(new_n196_), .A3(new_n381_), .A4(new_n466_), .ZN(new_n469_));
  NOR4_X1    g00277(.A1(new_n440_), .A2(new_n358_), .A3(new_n469_), .A4(new_n447_), .ZN(\asqrt[58] ));
  NAND3_X1   g00278(.A1(\asqrt[58] ), .A2(new_n465_), .A3(new_n468_), .ZN(new_n471_));
  OAI21_X1   g00279(.A1(new_n443_), .A2(\asqrt[62] ), .B(new_n395_), .ZN(new_n472_));
  OAI21_X1   g00280(.A1(\asqrt[58] ), .A2(new_n472_), .B(new_n465_), .ZN(new_n473_));
  NAND2_X1   g00281(.A1(new_n473_), .A2(new_n471_), .ZN(new_n474_));
  INV_X1     g00282(.I(new_n474_), .ZN(new_n475_));
  NOR3_X1    g00283(.A1(new_n417_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n476_));
  AOI21_X1   g00284(.A1(new_n425_), .A2(new_n421_), .B(\asqrt[61] ), .ZN(new_n477_));
  NAND4_X1   g00285(.A1(\asqrt[58] ), .A2(new_n476_), .A3(new_n442_), .A4(new_n477_), .ZN(new_n478_));
  NAND2_X1   g00286(.A1(new_n433_), .A2(\asqrt[61] ), .ZN(new_n479_));
  NAND2_X1   g00287(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1     g00288(.I(new_n480_), .ZN(new_n481_));
  NOR2_X1    g00289(.A1(new_n481_), .A2(new_n196_), .ZN(new_n482_));
  INV_X1     g00290(.I(new_n482_), .ZN(new_n483_));
  INV_X1     g00291(.I(\a[116] ), .ZN(new_n484_));
  NOR2_X1    g00292(.A1(\a[114] ), .A2(\a[115] ), .ZN(new_n485_));
  AOI21_X1   g00293(.A1(new_n484_), .A2(new_n485_), .B(new_n375_), .ZN(new_n486_));
  NAND2_X1   g00294(.A1(new_n352_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1    g00295(.A1(new_n487_), .A2(\a[117] ), .Z(new_n488_));
  INV_X1     g00296(.I(new_n488_), .ZN(new_n489_));
  NOR3_X1    g00297(.A1(new_n476_), .A2(new_n229_), .A3(new_n434_), .ZN(new_n490_));
  AOI21_X1   g00298(.A1(new_n490_), .A2(new_n462_), .B(new_n396_), .ZN(new_n491_));
  INV_X1     g00299(.I(new_n439_), .ZN(new_n492_));
  AOI21_X1   g00300(.A1(new_n491_), .A2(new_n492_), .B(new_n441_), .ZN(new_n493_));
  AOI21_X1   g00301(.A1(new_n443_), .A2(\asqrt[62] ), .B(new_n381_), .ZN(new_n494_));
  NOR3_X1    g00302(.A1(new_n494_), .A2(new_n467_), .A3(new_n447_), .ZN(new_n495_));
  NAND4_X1   g00303(.A1(new_n495_), .A2(\a[117] ), .A3(new_n493_), .A4(new_n359_), .ZN(new_n496_));
  NOR2_X1    g00304(.A1(new_n488_), .A2(\a[116] ), .ZN(new_n497_));
  INV_X1     g00305(.I(new_n497_), .ZN(new_n498_));
  AOI21_X1   g00306(.A1(new_n496_), .A2(new_n498_), .B(new_n489_), .ZN(new_n499_));
  INV_X1     g00307(.I(\a[117] ), .ZN(new_n500_));
  NOR4_X1    g00308(.A1(new_n449_), .A2(new_n500_), .A3(new_n440_), .A4(new_n358_), .ZN(new_n501_));
  NOR3_X1    g00309(.A1(new_n501_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n502_));
  NOR2_X1    g00310(.A1(new_n502_), .A2(new_n499_), .ZN(new_n503_));
  NAND4_X1   g00311(.A1(new_n493_), .A2(new_n359_), .A3(new_n444_), .A4(new_n448_), .ZN(new_n504_));
  NAND2_X1   g00312(.A1(\asqrt[59] ), .A2(\a[116] ), .ZN(new_n505_));
  AOI21_X1   g00313(.A1(new_n504_), .A2(\asqrt[59] ), .B(new_n505_), .ZN(new_n506_));
  NOR3_X1    g00314(.A1(\asqrt[58] ), .A2(\a[116] ), .A3(new_n376_), .ZN(new_n507_));
  OAI21_X1   g00315(.A1(new_n507_), .A2(new_n506_), .B(new_n485_), .ZN(new_n508_));
  NOR3_X1    g00316(.A1(new_n448_), .A2(new_n359_), .A3(new_n376_), .ZN(new_n509_));
  INV_X1     g00317(.I(new_n509_), .ZN(new_n510_));
  NOR2_X1    g00318(.A1(new_n444_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1   g00319(.A1(new_n511_), .A2(new_n440_), .B(\a[118] ), .ZN(new_n512_));
  NOR3_X1    g00320(.A1(new_n512_), .A2(\asqrt[58] ), .A3(new_n400_), .ZN(new_n513_));
  NAND2_X1   g00321(.A1(new_n469_), .A2(new_n509_), .ZN(new_n514_));
  OAI21_X1   g00322(.A1(new_n514_), .A2(new_n493_), .B(new_n415_), .ZN(new_n515_));
  AOI21_X1   g00323(.A1(new_n515_), .A2(new_n399_), .B(new_n504_), .ZN(new_n516_));
  NOR3_X1    g00324(.A1(new_n516_), .A2(new_n513_), .A3(\asqrt[60] ), .ZN(new_n517_));
  AOI21_X1   g00325(.A1(new_n508_), .A2(new_n517_), .B(new_n503_), .ZN(new_n518_));
  OAI21_X1   g00326(.A1(new_n501_), .A2(new_n497_), .B(new_n488_), .ZN(new_n519_));
  NAND3_X1   g00327(.A1(new_n496_), .A2(\a[116] ), .A3(new_n489_), .ZN(new_n520_));
  NAND2_X1   g00328(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1     g00329(.I(new_n485_), .ZN(new_n522_));
  NOR3_X1    g00330(.A1(new_n427_), .A2(new_n442_), .A3(new_n434_), .ZN(new_n523_));
  NOR3_X1    g00331(.A1(new_n523_), .A2(new_n396_), .A3(new_n439_), .ZN(new_n524_));
  NOR4_X1    g00332(.A1(new_n524_), .A2(new_n469_), .A3(new_n441_), .A4(new_n447_), .ZN(new_n525_));
  NAND4_X1   g00333(.A1(new_n525_), .A2(\a[116] ), .A3(new_n359_), .A4(\asqrt[59] ), .ZN(new_n526_));
  NAND3_X1   g00334(.A1(new_n504_), .A2(new_n484_), .A3(\asqrt[59] ), .ZN(new_n527_));
  AOI21_X1   g00335(.A1(new_n527_), .A2(new_n526_), .B(new_n522_), .ZN(new_n528_));
  OAI21_X1   g00336(.A1(new_n521_), .A2(new_n528_), .B(\asqrt[60] ), .ZN(new_n529_));
  NOR2_X1    g00337(.A1(new_n376_), .A2(\a[118] ), .ZN(new_n530_));
  OAI22_X1   g00338(.A1(new_n530_), .A2(\a[119] ), .B1(\a[118] ), .B2(new_n411_), .ZN(new_n531_));
  NAND2_X1   g00339(.A1(new_n417_), .A2(new_n402_), .ZN(new_n532_));
  NAND2_X1   g00340(.A1(new_n532_), .A2(new_n415_), .ZN(new_n533_));
  NAND2_X1   g00341(.A1(new_n533_), .A2(\asqrt[59] ), .ZN(new_n534_));
  NOR2_X1    g00342(.A1(new_n504_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1    g00343(.A1(new_n535_), .A2(new_n531_), .ZN(new_n536_));
  INV_X1     g00344(.I(new_n531_), .ZN(new_n537_));
  NOR3_X1    g00345(.A1(new_n504_), .A2(new_n537_), .A3(new_n534_), .ZN(new_n538_));
  NOR3_X1    g00346(.A1(new_n536_), .A2(new_n538_), .A3(\asqrt[61] ), .ZN(new_n539_));
  NAND2_X1   g00347(.A1(new_n529_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1   g00348(.A1(new_n540_), .A2(new_n518_), .ZN(new_n541_));
  NAND3_X1   g00349(.A1(new_n515_), .A2(new_n504_), .A3(new_n399_), .ZN(new_n542_));
  OAI21_X1   g00350(.A1(new_n512_), .A2(new_n400_), .B(\asqrt[58] ), .ZN(new_n543_));
  NAND3_X1   g00351(.A1(new_n543_), .A2(new_n542_), .A3(new_n275_), .ZN(new_n544_));
  OAI21_X1   g00352(.A1(new_n528_), .A2(new_n544_), .B(new_n521_), .ZN(new_n545_));
  AOI21_X1   g00353(.A1(new_n545_), .A2(new_n529_), .B(new_n229_), .ZN(new_n546_));
  NOR2_X1    g00354(.A1(new_n480_), .A2(\asqrt[62] ), .ZN(new_n547_));
  INV_X1     g00355(.I(new_n547_), .ZN(new_n548_));
  NAND2_X1   g00356(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  OAI21_X1   g00357(.A1(new_n549_), .A2(new_n541_), .B(new_n483_), .ZN(new_n550_));
  NOR3_X1    g00358(.A1(\asqrt[58] ), .A2(new_n381_), .A3(new_n444_), .ZN(new_n551_));
  OAI21_X1   g00359(.A1(new_n551_), .A2(new_n491_), .B(new_n231_), .ZN(new_n552_));
  OAI21_X1   g00360(.A1(new_n550_), .A2(new_n552_), .B(new_n475_), .ZN(new_n553_));
  NAND2_X1   g00361(.A1(new_n545_), .A2(new_n529_), .ZN(new_n554_));
  AOI22_X1   g00362(.A1(new_n554_), .A2(\asqrt[61] ), .B1(new_n540_), .B2(new_n518_), .ZN(new_n555_));
  OAI21_X1   g00363(.A1(new_n555_), .A2(new_n196_), .B(new_n474_), .ZN(new_n556_));
  AOI21_X1   g00364(.A1(new_n529_), .A2(new_n539_), .B(new_n545_), .ZN(new_n557_));
  NOR4_X1    g00365(.A1(new_n557_), .A2(\asqrt[62] ), .A3(new_n546_), .A4(new_n481_), .ZN(new_n558_));
  AOI21_X1   g00366(.A1(new_n441_), .A2(new_n491_), .B(new_n504_), .ZN(new_n559_));
  XOR2_X1    g00367(.A1(new_n437_), .A2(new_n231_), .Z(new_n560_));
  NOR2_X1    g00368(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1   g00369(.A1(new_n556_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_));
  NAND3_X1   g00370(.A1(new_n525_), .A2(new_n358_), .A3(new_n381_), .ZN(new_n563_));
  NOR4_X1    g00371(.A1(new_n562_), .A2(new_n553_), .A3(new_n230_), .A4(new_n563_), .ZN(new_n564_));
  NOR2_X1    g00372(.A1(new_n454_), .A2(\a[114] ), .ZN(new_n565_));
  OAI21_X1   g00373(.A1(new_n564_), .A2(new_n565_), .B(new_n454_), .ZN(new_n566_));
  INV_X1     g00374(.I(new_n454_), .ZN(new_n567_));
  AOI21_X1   g00375(.A1(new_n503_), .A2(new_n508_), .B(new_n275_), .ZN(new_n568_));
  OAI21_X1   g00376(.A1(new_n518_), .A2(new_n568_), .B(\asqrt[61] ), .ZN(new_n569_));
  NOR2_X1    g00377(.A1(new_n569_), .A2(new_n547_), .ZN(new_n570_));
  AOI21_X1   g00378(.A1(new_n570_), .A2(new_n557_), .B(new_n482_), .ZN(new_n571_));
  INV_X1     g00379(.I(new_n552_), .ZN(new_n572_));
  AOI21_X1   g00380(.A1(new_n571_), .A2(new_n572_), .B(new_n474_), .ZN(new_n573_));
  NAND4_X1   g00381(.A1(new_n555_), .A2(new_n196_), .A3(new_n475_), .A4(new_n480_), .ZN(new_n574_));
  INV_X1     g00382(.I(new_n561_), .ZN(new_n575_));
  NOR2_X1    g00383(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1     g00384(.I(new_n563_), .ZN(new_n577_));
  NAND4_X1   g00385(.A1(new_n576_), .A2(new_n573_), .A3(\a[115] ), .A4(new_n577_), .ZN(new_n578_));
  NAND3_X1   g00386(.A1(new_n578_), .A2(\a[114] ), .A3(new_n567_), .ZN(new_n579_));
  NAND2_X1   g00387(.A1(new_n566_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1    g00388(.A1(new_n562_), .A2(new_n553_), .ZN(new_n581_));
  NOR4_X1    g00389(.A1(new_n449_), .A2(new_n358_), .A3(new_n441_), .A4(new_n524_), .ZN(new_n582_));
  NAND2_X1   g00390(.A1(\asqrt[58] ), .A2(\a[114] ), .ZN(new_n583_));
  XOR2_X1    g00391(.A1(new_n583_), .A2(new_n582_), .Z(new_n584_));
  NOR2_X1    g00392(.A1(new_n584_), .A2(new_n451_), .ZN(new_n585_));
  INV_X1     g00393(.I(new_n585_), .ZN(new_n586_));
  NAND3_X1   g00394(.A1(new_n576_), .A2(new_n573_), .A3(new_n577_), .ZN(new_n587_));
  NOR2_X1    g00395(.A1(new_n577_), .A2(new_n504_), .ZN(new_n588_));
  NAND3_X1   g00396(.A1(new_n574_), .A2(new_n575_), .A3(new_n588_), .ZN(new_n589_));
  OAI21_X1   g00397(.A1(new_n589_), .A2(new_n573_), .B(new_n484_), .ZN(new_n590_));
  NAND3_X1   g00398(.A1(new_n590_), .A2(new_n587_), .A3(new_n485_), .ZN(new_n591_));
  NOR3_X1    g00399(.A1(new_n562_), .A2(new_n553_), .A3(new_n563_), .ZN(\asqrt[57] ));
  NAND2_X1   g00400(.A1(new_n575_), .A2(new_n588_), .ZN(new_n593_));
  AOI21_X1   g00401(.A1(new_n556_), .A2(new_n558_), .B(new_n593_), .ZN(new_n594_));
  AOI21_X1   g00402(.A1(new_n594_), .A2(new_n553_), .B(\a[116] ), .ZN(new_n595_));
  OAI21_X1   g00403(.A1(new_n522_), .A2(new_n595_), .B(\asqrt[57] ), .ZN(new_n596_));
  NAND4_X1   g00404(.A1(new_n596_), .A2(new_n591_), .A3(new_n376_), .A4(new_n586_), .ZN(new_n597_));
  NAND2_X1   g00405(.A1(new_n597_), .A2(new_n580_), .ZN(new_n598_));
  NAND3_X1   g00406(.A1(new_n566_), .A2(new_n579_), .A3(new_n586_), .ZN(new_n599_));
  NOR2_X1    g00407(.A1(new_n504_), .A2(\a[116] ), .ZN(new_n600_));
  OAI22_X1   g00408(.A1(new_n600_), .A2(\a[117] ), .B1(\a[116] ), .B2(new_n496_), .ZN(new_n601_));
  INV_X1     g00409(.I(new_n601_), .ZN(new_n602_));
  OAI21_X1   g00410(.A1(new_n508_), .A2(new_n487_), .B(new_n484_), .ZN(new_n603_));
  NAND2_X1   g00411(.A1(new_n603_), .A2(\asqrt[58] ), .ZN(new_n604_));
  OAI21_X1   g00412(.A1(new_n587_), .A2(new_n604_), .B(new_n602_), .ZN(new_n605_));
  INV_X1     g00413(.I(new_n604_), .ZN(new_n606_));
  NAND3_X1   g00414(.A1(\asqrt[57] ), .A2(new_n601_), .A3(new_n606_), .ZN(new_n607_));
  NAND3_X1   g00415(.A1(new_n605_), .A2(new_n607_), .A3(new_n275_), .ZN(new_n608_));
  AOI21_X1   g00416(.A1(new_n599_), .A2(\asqrt[59] ), .B(new_n608_), .ZN(new_n609_));
  NOR2_X1    g00417(.A1(new_n609_), .A2(new_n598_), .ZN(new_n610_));
  AOI22_X1   g00418(.A1(new_n597_), .A2(new_n580_), .B1(new_n599_), .B2(\asqrt[59] ), .ZN(new_n611_));
  OAI22_X1   g00419(.A1(new_n611_), .A2(new_n275_), .B1(new_n609_), .B2(new_n598_), .ZN(new_n612_));
  NOR2_X1    g00420(.A1(new_n516_), .A2(new_n513_), .ZN(new_n613_));
  NAND2_X1   g00421(.A1(new_n503_), .A2(new_n508_), .ZN(new_n614_));
  NOR4_X1    g00422(.A1(new_n587_), .A2(\asqrt[60] ), .A3(new_n613_), .A4(new_n614_), .ZN(new_n615_));
  OAI21_X1   g00423(.A1(new_n521_), .A2(new_n528_), .B(\asqrt[60] ), .ZN(new_n616_));
  INV_X1     g00424(.I(new_n616_), .ZN(new_n617_));
  NOR3_X1    g00425(.A1(new_n615_), .A2(\asqrt[61] ), .A3(new_n617_), .ZN(new_n618_));
  OAI21_X1   g00426(.A1(new_n611_), .A2(new_n275_), .B(new_n618_), .ZN(new_n619_));
  AOI22_X1   g00427(.A1(new_n612_), .A2(\asqrt[61] ), .B1(new_n619_), .B2(new_n610_), .ZN(new_n620_));
  NOR2_X1    g00428(.A1(new_n620_), .A2(new_n196_), .ZN(new_n621_));
  NOR2_X1    g00429(.A1(new_n536_), .A2(new_n538_), .ZN(new_n622_));
  NOR4_X1    g00430(.A1(new_n587_), .A2(\asqrt[61] ), .A3(new_n622_), .A4(new_n554_), .ZN(new_n623_));
  XOR2_X1    g00431(.A1(new_n623_), .A2(new_n569_), .Z(new_n624_));
  INV_X1     g00432(.I(new_n565_), .ZN(new_n625_));
  AOI21_X1   g00433(.A1(new_n578_), .A2(new_n625_), .B(new_n567_), .ZN(new_n626_));
  INV_X1     g00434(.I(\a[114] ), .ZN(new_n627_));
  NOR3_X1    g00435(.A1(new_n564_), .A2(new_n627_), .A3(new_n454_), .ZN(new_n628_));
  NOR3_X1    g00436(.A1(new_n628_), .A2(new_n626_), .A3(new_n585_), .ZN(new_n629_));
  AOI21_X1   g00437(.A1(\asqrt[57] ), .A2(new_n606_), .B(new_n601_), .ZN(new_n630_));
  NOR3_X1    g00438(.A1(new_n587_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n631_));
  NOR3_X1    g00439(.A1(new_n631_), .A2(new_n630_), .A3(\asqrt[60] ), .ZN(new_n632_));
  OAI21_X1   g00440(.A1(new_n629_), .A2(new_n376_), .B(new_n632_), .ZN(new_n633_));
  NAND3_X1   g00441(.A1(new_n633_), .A2(new_n580_), .A3(new_n597_), .ZN(new_n634_));
  NOR2_X1    g00442(.A1(new_n628_), .A2(new_n626_), .ZN(new_n635_));
  NOR3_X1    g00443(.A1(new_n595_), .A2(\asqrt[57] ), .A3(new_n522_), .ZN(new_n636_));
  AOI21_X1   g00444(.A1(new_n590_), .A2(new_n485_), .B(new_n587_), .ZN(new_n637_));
  NOR4_X1    g00445(.A1(new_n637_), .A2(new_n636_), .A3(\asqrt[59] ), .A4(new_n585_), .ZN(new_n638_));
  OAI22_X1   g00446(.A1(new_n638_), .A2(new_n635_), .B1(new_n629_), .B2(new_n376_), .ZN(new_n639_));
  NAND2_X1   g00447(.A1(new_n639_), .A2(\asqrt[60] ), .ZN(new_n640_));
  AOI21_X1   g00448(.A1(new_n640_), .A2(new_n634_), .B(new_n229_), .ZN(new_n641_));
  INV_X1     g00449(.I(new_n618_), .ZN(new_n642_));
  AOI21_X1   g00450(.A1(new_n639_), .A2(\asqrt[60] ), .B(new_n642_), .ZN(new_n643_));
  NOR2_X1    g00451(.A1(new_n643_), .A2(new_n634_), .ZN(new_n644_));
  NOR4_X1    g00452(.A1(new_n644_), .A2(new_n641_), .A3(\asqrt[62] ), .A4(new_n624_), .ZN(new_n645_));
  NOR2_X1    g00453(.A1(new_n474_), .A2(new_n577_), .ZN(new_n646_));
  NAND2_X1   g00454(.A1(new_n581_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1     g00455(.I(new_n555_), .ZN(new_n648_));
  NAND2_X1   g00456(.A1(new_n648_), .A2(\asqrt[62] ), .ZN(new_n649_));
  INV_X1     g00457(.I(new_n558_), .ZN(new_n650_));
  NOR3_X1    g00458(.A1(new_n587_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  NOR2_X1    g00459(.A1(new_n648_), .A2(\asqrt[62] ), .ZN(new_n652_));
  NOR2_X1    g00460(.A1(new_n652_), .A2(new_n480_), .ZN(new_n653_));
  AOI21_X1   g00461(.A1(new_n587_), .A2(new_n653_), .B(new_n649_), .ZN(new_n654_));
  NOR2_X1    g00462(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1    g00463(.A1(new_n624_), .A2(new_n196_), .ZN(new_n656_));
  INV_X1     g00464(.I(new_n656_), .ZN(new_n657_));
  NAND2_X1   g00465(.A1(new_n599_), .A2(\asqrt[59] ), .ZN(new_n658_));
  AOI21_X1   g00466(.A1(new_n598_), .A2(new_n658_), .B(new_n275_), .ZN(new_n659_));
  OAI21_X1   g00467(.A1(new_n659_), .A2(new_n610_), .B(\asqrt[61] ), .ZN(new_n660_));
  NAND2_X1   g00468(.A1(new_n624_), .A2(new_n196_), .ZN(new_n661_));
  NAND3_X1   g00469(.A1(new_n619_), .A2(new_n610_), .A3(new_n661_), .ZN(new_n662_));
  OAI21_X1   g00470(.A1(new_n662_), .A2(new_n660_), .B(new_n657_), .ZN(new_n663_));
  NAND3_X1   g00471(.A1(new_n587_), .A2(new_n474_), .A3(new_n574_), .ZN(new_n664_));
  AOI21_X1   g00472(.A1(new_n664_), .A2(new_n550_), .B(\asqrt[63] ), .ZN(new_n665_));
  INV_X1     g00473(.I(new_n665_), .ZN(new_n666_));
  OAI21_X1   g00474(.A1(new_n663_), .A2(new_n666_), .B(new_n655_), .ZN(new_n667_));
  XOR2_X1    g00475(.A1(new_n623_), .A2(new_n546_), .Z(new_n668_));
  NAND4_X1   g00476(.A1(new_n620_), .A2(new_n196_), .A3(new_n655_), .A4(new_n668_), .ZN(new_n669_));
  OAI21_X1   g00477(.A1(new_n475_), .A2(new_n550_), .B(\asqrt[57] ), .ZN(new_n670_));
  XOR2_X1    g00478(.A1(new_n550_), .A2(\asqrt[63] ), .Z(new_n671_));
  NAND2_X1   g00479(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NOR4_X1    g00480(.A1(new_n667_), .A2(new_n647_), .A3(new_n669_), .A4(new_n672_), .ZN(\asqrt[56] ));
  NAND3_X1   g00481(.A1(\asqrt[56] ), .A2(new_n621_), .A3(new_n645_), .ZN(new_n674_));
  NAND2_X1   g00482(.A1(new_n619_), .A2(new_n610_), .ZN(new_n675_));
  NAND2_X1   g00483(.A1(new_n675_), .A2(new_n660_), .ZN(new_n676_));
  OAI21_X1   g00484(.A1(new_n676_), .A2(\asqrt[62] ), .B(new_n624_), .ZN(new_n677_));
  OAI21_X1   g00485(.A1(\asqrt[56] ), .A2(new_n677_), .B(new_n621_), .ZN(new_n678_));
  NAND2_X1   g00486(.A1(new_n678_), .A2(new_n674_), .ZN(new_n679_));
  INV_X1     g00487(.I(new_n679_), .ZN(new_n680_));
  NOR2_X1    g00488(.A1(new_n615_), .A2(new_n617_), .ZN(new_n681_));
  NOR3_X1    g00489(.A1(new_n612_), .A2(\asqrt[61] ), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1   g00490(.A1(\asqrt[56] ), .A2(new_n682_), .ZN(new_n683_));
  XOR2_X1    g00491(.A1(new_n683_), .A2(new_n641_), .Z(new_n684_));
  NOR2_X1    g00492(.A1(new_n684_), .A2(new_n196_), .ZN(new_n685_));
  INV_X1     g00493(.I(new_n685_), .ZN(new_n686_));
  INV_X1     g00494(.I(\a[112] ), .ZN(new_n687_));
  NOR2_X1    g00495(.A1(\a[110] ), .A2(\a[111] ), .ZN(new_n688_));
  AOI21_X1   g00496(.A1(new_n687_), .A2(new_n688_), .B(new_n577_), .ZN(new_n689_));
  NAND2_X1   g00497(.A1(new_n581_), .A2(new_n689_), .ZN(new_n690_));
  XOR2_X1    g00498(.A1(new_n690_), .A2(\a[113] ), .Z(new_n691_));
  INV_X1     g00499(.I(new_n691_), .ZN(new_n692_));
  INV_X1     g00500(.I(new_n647_), .ZN(new_n693_));
  INV_X1     g00501(.I(new_n655_), .ZN(new_n694_));
  NOR2_X1    g00502(.A1(new_n668_), .A2(\asqrt[62] ), .ZN(new_n695_));
  NOR3_X1    g00503(.A1(new_n643_), .A2(new_n634_), .A3(new_n695_), .ZN(new_n696_));
  AOI21_X1   g00504(.A1(new_n696_), .A2(new_n641_), .B(new_n656_), .ZN(new_n697_));
  AOI21_X1   g00505(.A1(new_n697_), .A2(new_n665_), .B(new_n694_), .ZN(new_n698_));
  NOR2_X1    g00506(.A1(new_n669_), .A2(new_n672_), .ZN(new_n699_));
  NAND4_X1   g00507(.A1(new_n699_), .A2(\a[113] ), .A3(new_n698_), .A4(new_n693_), .ZN(new_n700_));
  NOR2_X1    g00508(.A1(new_n691_), .A2(\a[112] ), .ZN(new_n701_));
  INV_X1     g00509(.I(new_n701_), .ZN(new_n702_));
  AOI21_X1   g00510(.A1(new_n700_), .A2(new_n702_), .B(new_n692_), .ZN(new_n703_));
  INV_X1     g00511(.I(\a[113] ), .ZN(new_n704_));
  OAI21_X1   g00512(.A1(new_n620_), .A2(new_n196_), .B(new_n694_), .ZN(new_n705_));
  INV_X1     g00513(.I(new_n672_), .ZN(new_n706_));
  NAND3_X1   g00514(.A1(new_n705_), .A2(new_n645_), .A3(new_n706_), .ZN(new_n707_));
  NOR4_X1    g00515(.A1(new_n707_), .A2(new_n704_), .A3(new_n647_), .A4(new_n667_), .ZN(new_n708_));
  NOR3_X1    g00516(.A1(new_n708_), .A2(new_n687_), .A3(new_n691_), .ZN(new_n709_));
  NOR2_X1    g00517(.A1(new_n709_), .A2(new_n703_), .ZN(new_n710_));
  INV_X1     g00518(.I(new_n688_), .ZN(new_n711_));
  NAND2_X1   g00519(.A1(new_n571_), .A2(new_n572_), .ZN(new_n712_));
  NOR2_X1    g00520(.A1(new_n707_), .A2(new_n667_), .ZN(new_n713_));
  NAND4_X1   g00521(.A1(new_n576_), .A2(new_n475_), .A3(new_n712_), .A4(new_n577_), .ZN(new_n714_));
  NOR2_X1    g00522(.A1(new_n587_), .A2(new_n687_), .ZN(new_n715_));
  XOR2_X1    g00523(.A1(new_n715_), .A2(new_n714_), .Z(new_n716_));
  NOR2_X1    g00524(.A1(new_n716_), .A2(new_n711_), .ZN(new_n717_));
  NOR3_X1    g00525(.A1(new_n706_), .A2(new_n693_), .A3(new_n587_), .ZN(new_n718_));
  INV_X1     g00526(.I(new_n718_), .ZN(new_n719_));
  AOI21_X1   g00527(.A1(new_n705_), .A2(new_n645_), .B(new_n719_), .ZN(new_n720_));
  AOI21_X1   g00528(.A1(new_n720_), .A2(new_n667_), .B(\a[114] ), .ZN(new_n721_));
  NOR3_X1    g00529(.A1(new_n721_), .A2(new_n451_), .A3(\asqrt[56] ), .ZN(new_n722_));
  NOR4_X1    g00530(.A1(new_n676_), .A2(\asqrt[62] ), .A3(new_n694_), .A4(new_n624_), .ZN(new_n723_));
  NAND4_X1   g00531(.A1(new_n698_), .A2(new_n693_), .A3(new_n723_), .A4(new_n706_), .ZN(new_n724_));
  NAND2_X1   g00532(.A1(new_n669_), .A2(new_n718_), .ZN(new_n725_));
  OAI21_X1   g00533(.A1(new_n725_), .A2(new_n698_), .B(new_n627_), .ZN(new_n726_));
  AOI21_X1   g00534(.A1(new_n726_), .A2(new_n450_), .B(new_n724_), .ZN(new_n727_));
  NOR4_X1    g00535(.A1(new_n727_), .A2(new_n722_), .A3(\asqrt[58] ), .A4(new_n717_), .ZN(new_n728_));
  NOR2_X1    g00536(.A1(new_n728_), .A2(new_n710_), .ZN(new_n729_));
  NOR3_X1    g00537(.A1(new_n709_), .A2(new_n703_), .A3(new_n717_), .ZN(new_n730_));
  NAND2_X1   g00538(.A1(\asqrt[57] ), .A2(new_n627_), .ZN(new_n731_));
  AOI22_X1   g00539(.A1(new_n731_), .A2(new_n230_), .B1(new_n627_), .B2(new_n564_), .ZN(new_n732_));
  INV_X1     g00540(.I(new_n732_), .ZN(new_n733_));
  AOI21_X1   g00541(.A1(new_n585_), .A2(new_n453_), .B(\a[114] ), .ZN(new_n734_));
  NOR2_X1    g00542(.A1(new_n587_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1   g00543(.A1(\asqrt[56] ), .A2(new_n735_), .B(new_n733_), .ZN(new_n736_));
  INV_X1     g00544(.I(new_n735_), .ZN(new_n737_));
  NOR3_X1    g00545(.A1(new_n724_), .A2(new_n732_), .A3(new_n737_), .ZN(new_n738_));
  NOR3_X1    g00546(.A1(new_n738_), .A2(new_n736_), .A3(\asqrt[59] ), .ZN(new_n739_));
  OAI21_X1   g00547(.A1(new_n730_), .A2(new_n504_), .B(new_n739_), .ZN(new_n740_));
  NAND2_X1   g00548(.A1(new_n740_), .A2(new_n729_), .ZN(new_n741_));
  OAI22_X1   g00549(.A1(new_n710_), .A2(new_n728_), .B1(new_n730_), .B2(new_n504_), .ZN(new_n742_));
  NAND2_X1   g00550(.A1(new_n742_), .A2(\asqrt[59] ), .ZN(new_n743_));
  AOI21_X1   g00551(.A1(new_n596_), .A2(new_n591_), .B(\asqrt[59] ), .ZN(new_n744_));
  AND4_X2    g00552(.A1(new_n629_), .A2(\asqrt[56] ), .A3(new_n658_), .A4(new_n744_), .Z(new_n745_));
  NOR2_X1    g00553(.A1(new_n629_), .A2(new_n376_), .ZN(new_n746_));
  NOR3_X1    g00554(.A1(new_n745_), .A2(new_n746_), .A3(\asqrt[60] ), .ZN(new_n747_));
  AOI21_X1   g00555(.A1(new_n743_), .A2(new_n747_), .B(new_n741_), .ZN(new_n748_));
  AOI21_X1   g00556(.A1(new_n743_), .A2(new_n741_), .B(new_n275_), .ZN(new_n749_));
  OAI21_X1   g00557(.A1(new_n748_), .A2(new_n749_), .B(\asqrt[61] ), .ZN(new_n750_));
  AOI22_X1   g00558(.A1(new_n742_), .A2(\asqrt[59] ), .B1(new_n729_), .B2(new_n740_), .ZN(new_n751_));
  NAND2_X1   g00559(.A1(new_n605_), .A2(new_n607_), .ZN(new_n752_));
  NAND4_X1   g00560(.A1(\asqrt[56] ), .A2(new_n275_), .A3(new_n752_), .A4(new_n611_), .ZN(new_n753_));
  XOR2_X1    g00561(.A1(new_n753_), .A2(new_n659_), .Z(new_n754_));
  NAND2_X1   g00562(.A1(new_n754_), .A2(new_n229_), .ZN(new_n755_));
  INV_X1     g00563(.I(new_n755_), .ZN(new_n756_));
  OAI21_X1   g00564(.A1(new_n751_), .A2(new_n275_), .B(new_n756_), .ZN(new_n757_));
  INV_X1     g00565(.I(new_n684_), .ZN(new_n758_));
  NOR2_X1    g00566(.A1(new_n758_), .A2(\asqrt[62] ), .ZN(new_n759_));
  INV_X1     g00567(.I(new_n759_), .ZN(new_n760_));
  NAND3_X1   g00568(.A1(new_n757_), .A2(new_n748_), .A3(new_n760_), .ZN(new_n761_));
  OAI21_X1   g00569(.A1(new_n761_), .A2(new_n750_), .B(new_n686_), .ZN(new_n762_));
  NAND3_X1   g00570(.A1(new_n724_), .A2(new_n694_), .A3(new_n669_), .ZN(new_n763_));
  AOI21_X1   g00571(.A1(new_n763_), .A2(new_n663_), .B(\asqrt[63] ), .ZN(new_n764_));
  INV_X1     g00572(.I(new_n764_), .ZN(new_n765_));
  OAI21_X1   g00573(.A1(new_n762_), .A2(new_n765_), .B(new_n680_), .ZN(new_n766_));
  OAI21_X1   g00574(.A1(new_n708_), .A2(new_n701_), .B(new_n691_), .ZN(new_n767_));
  NAND3_X1   g00575(.A1(new_n700_), .A2(\a[112] ), .A3(new_n692_), .ZN(new_n768_));
  NAND2_X1   g00576(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1     g00577(.I(new_n717_), .ZN(new_n770_));
  NAND3_X1   g00578(.A1(new_n726_), .A2(new_n724_), .A3(new_n450_), .ZN(new_n771_));
  OAI21_X1   g00579(.A1(new_n721_), .A2(new_n451_), .B(\asqrt[56] ), .ZN(new_n772_));
  NAND4_X1   g00580(.A1(new_n772_), .A2(new_n771_), .A3(new_n504_), .A4(new_n770_), .ZN(new_n773_));
  NAND2_X1   g00581(.A1(new_n773_), .A2(new_n769_), .ZN(new_n774_));
  NAND3_X1   g00582(.A1(new_n767_), .A2(new_n768_), .A3(new_n770_), .ZN(new_n775_));
  OAI21_X1   g00583(.A1(new_n724_), .A2(new_n737_), .B(new_n732_), .ZN(new_n776_));
  NAND3_X1   g00584(.A1(\asqrt[56] ), .A2(new_n733_), .A3(new_n735_), .ZN(new_n777_));
  NAND3_X1   g00585(.A1(new_n776_), .A2(new_n777_), .A3(new_n376_), .ZN(new_n778_));
  AOI21_X1   g00586(.A1(new_n775_), .A2(\asqrt[58] ), .B(new_n778_), .ZN(new_n779_));
  NOR2_X1    g00587(.A1(new_n779_), .A2(new_n774_), .ZN(new_n780_));
  AOI22_X1   g00588(.A1(\asqrt[58] ), .A2(new_n775_), .B1(new_n773_), .B2(new_n769_), .ZN(new_n781_));
  OAI21_X1   g00589(.A1(new_n781_), .A2(new_n376_), .B(new_n747_), .ZN(new_n782_));
  NAND2_X1   g00590(.A1(new_n782_), .A2(new_n780_), .ZN(new_n783_));
  OAI22_X1   g00591(.A1(new_n781_), .A2(new_n376_), .B1(new_n774_), .B2(new_n779_), .ZN(new_n784_));
  AOI22_X1   g00592(.A1(new_n784_), .A2(\asqrt[60] ), .B1(new_n782_), .B2(new_n780_), .ZN(new_n785_));
  AOI21_X1   g00593(.A1(new_n784_), .A2(\asqrt[60] ), .B(new_n755_), .ZN(new_n786_));
  OAI22_X1   g00594(.A1(new_n785_), .A2(new_n229_), .B1(new_n786_), .B2(new_n783_), .ZN(new_n787_));
  NOR4_X1    g00595(.A1(new_n787_), .A2(\asqrt[62] ), .A3(new_n679_), .A4(new_n684_), .ZN(new_n788_));
  AOI21_X1   g00596(.A1(new_n694_), .A2(new_n697_), .B(new_n724_), .ZN(new_n789_));
  XOR2_X1    g00597(.A1(new_n663_), .A2(new_n231_), .Z(new_n790_));
  NOR2_X1    g00598(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1   g00599(.A1(new_n788_), .A2(new_n791_), .ZN(new_n792_));
  NOR2_X1    g00600(.A1(new_n792_), .A2(new_n766_), .ZN(new_n793_));
  INV_X1     g00601(.I(\a[108] ), .ZN(new_n794_));
  INV_X1     g00602(.I(new_n713_), .ZN(new_n795_));
  NOR3_X1    g00603(.A1(new_n795_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n796_));
  NOR2_X1    g00604(.A1(\a[106] ), .A2(\a[107] ), .ZN(new_n797_));
  AOI21_X1   g00605(.A1(new_n794_), .A2(new_n797_), .B(new_n796_), .ZN(new_n798_));
  NAND2_X1   g00606(.A1(new_n793_), .A2(new_n798_), .ZN(new_n799_));
  XOR2_X1    g00607(.A1(new_n799_), .A2(\a[109] ), .Z(new_n800_));
  INV_X1     g00608(.I(\a[109] ), .ZN(new_n801_));
  NOR2_X1    g00609(.A1(new_n679_), .A2(new_n796_), .ZN(new_n802_));
  NAND2_X1   g00610(.A1(new_n793_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1   g00611(.A1(new_n775_), .A2(\asqrt[58] ), .ZN(new_n804_));
  AOI21_X1   g00612(.A1(new_n774_), .A2(new_n804_), .B(new_n376_), .ZN(new_n805_));
  OAI21_X1   g00613(.A1(new_n805_), .A2(new_n780_), .B(\asqrt[60] ), .ZN(new_n806_));
  AOI21_X1   g00614(.A1(new_n783_), .A2(new_n806_), .B(new_n229_), .ZN(new_n807_));
  AOI21_X1   g00615(.A1(new_n748_), .A2(new_n757_), .B(new_n807_), .ZN(new_n808_));
  NOR2_X1    g00616(.A1(new_n808_), .A2(new_n196_), .ZN(new_n809_));
  NAND2_X1   g00617(.A1(new_n757_), .A2(new_n748_), .ZN(new_n810_));
  NAND4_X1   g00618(.A1(new_n810_), .A2(new_n750_), .A3(new_n196_), .A4(new_n758_), .ZN(new_n811_));
  INV_X1     g00619(.I(new_n811_), .ZN(new_n812_));
  NAND4_X1   g00620(.A1(new_n808_), .A2(new_n196_), .A3(new_n680_), .A4(new_n758_), .ZN(new_n813_));
  INV_X1     g00621(.I(new_n791_), .ZN(new_n814_));
  INV_X1     g00622(.I(new_n796_), .ZN(new_n815_));
  NOR4_X1    g00623(.A1(new_n766_), .A2(new_n813_), .A3(new_n814_), .A4(new_n815_), .ZN(\asqrt[55] ));
  NAND3_X1   g00624(.A1(\asqrt[55] ), .A2(new_n809_), .A3(new_n812_), .ZN(new_n817_));
  OAI21_X1   g00625(.A1(new_n787_), .A2(\asqrt[62] ), .B(new_n684_), .ZN(new_n818_));
  OAI21_X1   g00626(.A1(\asqrt[55] ), .A2(new_n818_), .B(new_n809_), .ZN(new_n819_));
  AND2_X2    g00627(.A1(new_n819_), .A2(new_n817_), .Z(new_n820_));
  INV_X1     g00628(.I(new_n785_), .ZN(new_n821_));
  NOR3_X1    g00629(.A1(new_n786_), .A2(new_n783_), .A3(new_n759_), .ZN(new_n822_));
  AOI21_X1   g00630(.A1(new_n822_), .A2(new_n807_), .B(new_n685_), .ZN(new_n823_));
  AOI21_X1   g00631(.A1(new_n823_), .A2(new_n764_), .B(new_n679_), .ZN(new_n824_));
  NAND4_X1   g00632(.A1(new_n824_), .A2(new_n788_), .A3(new_n791_), .A4(new_n796_), .ZN(new_n825_));
  NOR4_X1    g00633(.A1(new_n825_), .A2(\asqrt[61] ), .A3(new_n821_), .A4(new_n754_), .ZN(new_n826_));
  XOR2_X1    g00634(.A1(new_n826_), .A2(new_n750_), .Z(new_n827_));
  NOR2_X1    g00635(.A1(new_n827_), .A2(new_n196_), .ZN(new_n828_));
  INV_X1     g00636(.I(new_n828_), .ZN(new_n829_));
  INV_X1     g00637(.I(\a[110] ), .ZN(new_n830_));
  NOR2_X1    g00638(.A1(\a[108] ), .A2(\a[109] ), .ZN(new_n831_));
  AOI21_X1   g00639(.A1(new_n830_), .A2(new_n831_), .B(new_n693_), .ZN(new_n832_));
  NAND2_X1   g00640(.A1(new_n713_), .A2(new_n832_), .ZN(new_n833_));
  XOR2_X1    g00641(.A1(new_n833_), .A2(\a[111] ), .Z(new_n834_));
  INV_X1     g00642(.I(\a[111] ), .ZN(new_n835_));
  NOR4_X1    g00643(.A1(new_n792_), .A2(new_n835_), .A3(new_n766_), .A4(new_n815_), .ZN(new_n836_));
  NOR2_X1    g00644(.A1(new_n834_), .A2(\a[110] ), .ZN(new_n837_));
  OAI21_X1   g00645(.A1(new_n836_), .A2(new_n837_), .B(new_n834_), .ZN(new_n838_));
  INV_X1     g00646(.I(new_n834_), .ZN(new_n839_));
  AOI21_X1   g00647(.A1(new_n787_), .A2(\asqrt[62] ), .B(new_n680_), .ZN(new_n840_));
  NOR3_X1    g00648(.A1(new_n840_), .A2(new_n811_), .A3(new_n814_), .ZN(new_n841_));
  NAND4_X1   g00649(.A1(new_n841_), .A2(\a[111] ), .A3(new_n824_), .A4(new_n796_), .ZN(new_n842_));
  NAND3_X1   g00650(.A1(new_n842_), .A2(\a[110] ), .A3(new_n839_), .ZN(new_n843_));
  NAND2_X1   g00651(.A1(new_n838_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1     g00652(.I(new_n831_), .ZN(new_n845_));
  NAND2_X1   g00653(.A1(new_n697_), .A2(new_n665_), .ZN(new_n846_));
  NAND4_X1   g00654(.A1(new_n699_), .A2(new_n693_), .A3(new_n655_), .A4(new_n846_), .ZN(new_n847_));
  NOR2_X1    g00655(.A1(new_n724_), .A2(new_n830_), .ZN(new_n848_));
  XOR2_X1    g00656(.A1(new_n848_), .A2(new_n847_), .Z(new_n849_));
  NOR2_X1    g00657(.A1(new_n849_), .A2(new_n845_), .ZN(new_n850_));
  INV_X1     g00658(.I(new_n850_), .ZN(new_n851_));
  NOR3_X1    g00659(.A1(new_n791_), .A2(new_n796_), .A3(new_n724_), .ZN(new_n852_));
  OAI21_X1   g00660(.A1(new_n840_), .A2(new_n811_), .B(new_n852_), .ZN(new_n853_));
  OAI21_X1   g00661(.A1(new_n853_), .A2(new_n824_), .B(new_n687_), .ZN(new_n854_));
  NAND3_X1   g00662(.A1(new_n854_), .A2(new_n688_), .A3(new_n825_), .ZN(new_n855_));
  INV_X1     g00663(.I(new_n852_), .ZN(new_n856_));
  NOR2_X1    g00664(.A1(new_n788_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1   g00665(.A1(new_n857_), .A2(new_n766_), .B(\a[112] ), .ZN(new_n858_));
  OAI21_X1   g00666(.A1(new_n858_), .A2(new_n711_), .B(\asqrt[55] ), .ZN(new_n859_));
  NAND4_X1   g00667(.A1(new_n859_), .A2(new_n855_), .A3(new_n587_), .A4(new_n851_), .ZN(new_n860_));
  NAND2_X1   g00668(.A1(new_n860_), .A2(new_n844_), .ZN(new_n861_));
  NAND3_X1   g00669(.A1(new_n838_), .A2(new_n843_), .A3(new_n851_), .ZN(new_n862_));
  AOI21_X1   g00670(.A1(\asqrt[56] ), .A2(new_n687_), .B(\a[113] ), .ZN(new_n863_));
  NOR2_X1    g00671(.A1(new_n700_), .A2(\a[112] ), .ZN(new_n864_));
  NOR2_X1    g00672(.A1(new_n864_), .A2(new_n863_), .ZN(new_n865_));
  OAI21_X1   g00673(.A1(new_n770_), .A2(new_n690_), .B(new_n687_), .ZN(new_n866_));
  NAND2_X1   g00674(.A1(\asqrt[56] ), .A2(new_n866_), .ZN(new_n867_));
  OAI21_X1   g00675(.A1(new_n825_), .A2(new_n867_), .B(new_n865_), .ZN(new_n868_));
  INV_X1     g00676(.I(new_n865_), .ZN(new_n869_));
  INV_X1     g00677(.I(new_n867_), .ZN(new_n870_));
  NAND3_X1   g00678(.A1(\asqrt[55] ), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  NAND3_X1   g00679(.A1(new_n871_), .A2(new_n868_), .A3(new_n504_), .ZN(new_n872_));
  AOI21_X1   g00680(.A1(new_n862_), .A2(\asqrt[57] ), .B(new_n872_), .ZN(new_n873_));
  NOR2_X1    g00681(.A1(new_n873_), .A2(new_n861_), .ZN(new_n874_));
  AOI22_X1   g00682(.A1(new_n844_), .A2(new_n860_), .B1(new_n862_), .B2(\asqrt[57] ), .ZN(new_n875_));
  AOI21_X1   g00683(.A1(new_n772_), .A2(new_n771_), .B(\asqrt[58] ), .ZN(new_n876_));
  AND4_X2    g00684(.A1(new_n730_), .A2(\asqrt[55] ), .A3(new_n804_), .A4(new_n876_), .Z(new_n877_));
  NOR2_X1    g00685(.A1(new_n730_), .A2(new_n504_), .ZN(new_n878_));
  NOR3_X1    g00686(.A1(new_n877_), .A2(\asqrt[59] ), .A3(new_n878_), .ZN(new_n879_));
  OAI21_X1   g00687(.A1(new_n875_), .A2(new_n504_), .B(new_n879_), .ZN(new_n880_));
  NAND2_X1   g00688(.A1(new_n880_), .A2(new_n874_), .ZN(new_n881_));
  OAI22_X1   g00689(.A1(new_n875_), .A2(new_n504_), .B1(new_n861_), .B2(new_n873_), .ZN(new_n882_));
  NAND2_X1   g00690(.A1(new_n776_), .A2(new_n777_), .ZN(new_n883_));
  NAND4_X1   g00691(.A1(\asqrt[55] ), .A2(new_n376_), .A3(new_n883_), .A4(new_n781_), .ZN(new_n884_));
  XOR2_X1    g00692(.A1(new_n884_), .A2(new_n805_), .Z(new_n885_));
  NAND2_X1   g00693(.A1(new_n885_), .A2(new_n275_), .ZN(new_n886_));
  AOI21_X1   g00694(.A1(new_n882_), .A2(\asqrt[59] ), .B(new_n886_), .ZN(new_n887_));
  NOR2_X1    g00695(.A1(new_n887_), .A2(new_n881_), .ZN(new_n888_));
  NAND2_X1   g00696(.A1(new_n862_), .A2(\asqrt[57] ), .ZN(new_n889_));
  AOI21_X1   g00697(.A1(new_n861_), .A2(new_n889_), .B(new_n504_), .ZN(new_n890_));
  OAI21_X1   g00698(.A1(new_n890_), .A2(new_n874_), .B(\asqrt[59] ), .ZN(new_n891_));
  AOI21_X1   g00699(.A1(new_n881_), .A2(new_n891_), .B(new_n275_), .ZN(new_n892_));
  OAI21_X1   g00700(.A1(new_n888_), .A2(new_n892_), .B(\asqrt[61] ), .ZN(new_n893_));
  AOI22_X1   g00701(.A1(new_n882_), .A2(\asqrt[59] ), .B1(new_n880_), .B2(new_n874_), .ZN(new_n894_));
  OR2_X2     g00702(.A1(new_n745_), .A2(new_n746_), .Z(new_n895_));
  NAND4_X1   g00703(.A1(\asqrt[55] ), .A2(new_n275_), .A3(new_n895_), .A4(new_n751_), .ZN(new_n896_));
  XOR2_X1    g00704(.A1(new_n896_), .A2(new_n749_), .Z(new_n897_));
  NAND2_X1   g00705(.A1(new_n897_), .A2(new_n229_), .ZN(new_n898_));
  INV_X1     g00706(.I(new_n898_), .ZN(new_n899_));
  OAI21_X1   g00707(.A1(new_n894_), .A2(new_n275_), .B(new_n899_), .ZN(new_n900_));
  NAND2_X1   g00708(.A1(new_n827_), .A2(new_n196_), .ZN(new_n901_));
  NAND3_X1   g00709(.A1(new_n900_), .A2(new_n888_), .A3(new_n901_), .ZN(new_n902_));
  OAI21_X1   g00710(.A1(new_n902_), .A2(new_n893_), .B(new_n829_), .ZN(new_n903_));
  NOR3_X1    g00711(.A1(\asqrt[55] ), .A2(new_n680_), .A3(new_n788_), .ZN(new_n904_));
  OAI21_X1   g00712(.A1(new_n904_), .A2(new_n823_), .B(new_n231_), .ZN(new_n905_));
  OAI21_X1   g00713(.A1(new_n903_), .A2(new_n905_), .B(new_n820_), .ZN(new_n906_));
  INV_X1     g00714(.I(new_n820_), .ZN(new_n907_));
  OAI22_X1   g00715(.A1(new_n894_), .A2(new_n275_), .B1(new_n887_), .B2(new_n881_), .ZN(new_n908_));
  AOI22_X1   g00716(.A1(new_n908_), .A2(\asqrt[61] ), .B1(new_n900_), .B2(new_n888_), .ZN(new_n909_));
  OAI21_X1   g00717(.A1(new_n909_), .A2(new_n196_), .B(new_n907_), .ZN(new_n910_));
  INV_X1     g00718(.I(new_n837_), .ZN(new_n911_));
  AOI21_X1   g00719(.A1(new_n842_), .A2(new_n911_), .B(new_n839_), .ZN(new_n912_));
  NOR3_X1    g00720(.A1(new_n836_), .A2(new_n830_), .A3(new_n834_), .ZN(new_n913_));
  NOR2_X1    g00721(.A1(new_n913_), .A2(new_n912_), .ZN(new_n914_));
  NOR3_X1    g00722(.A1(new_n858_), .A2(\asqrt[55] ), .A3(new_n711_), .ZN(new_n915_));
  AOI21_X1   g00723(.A1(new_n854_), .A2(new_n688_), .B(new_n825_), .ZN(new_n916_));
  NOR4_X1    g00724(.A1(new_n915_), .A2(new_n916_), .A3(\asqrt[57] ), .A4(new_n850_), .ZN(new_n917_));
  NOR2_X1    g00725(.A1(new_n917_), .A2(new_n914_), .ZN(new_n918_));
  NOR3_X1    g00726(.A1(new_n913_), .A2(new_n912_), .A3(new_n850_), .ZN(new_n919_));
  AOI21_X1   g00727(.A1(\asqrt[55] ), .A2(new_n870_), .B(new_n869_), .ZN(new_n920_));
  NOR3_X1    g00728(.A1(new_n825_), .A2(new_n865_), .A3(new_n867_), .ZN(new_n921_));
  NOR3_X1    g00729(.A1(new_n920_), .A2(new_n921_), .A3(\asqrt[58] ), .ZN(new_n922_));
  OAI21_X1   g00730(.A1(new_n919_), .A2(new_n587_), .B(new_n922_), .ZN(new_n923_));
  NAND2_X1   g00731(.A1(new_n923_), .A2(new_n918_), .ZN(new_n924_));
  OAI22_X1   g00732(.A1(new_n917_), .A2(new_n914_), .B1(new_n919_), .B2(new_n587_), .ZN(new_n925_));
  INV_X1     g00733(.I(new_n879_), .ZN(new_n926_));
  AOI21_X1   g00734(.A1(new_n925_), .A2(\asqrt[58] ), .B(new_n926_), .ZN(new_n927_));
  NOR2_X1    g00735(.A1(new_n927_), .A2(new_n924_), .ZN(new_n928_));
  NAND2_X1   g00736(.A1(new_n925_), .A2(\asqrt[58] ), .ZN(new_n929_));
  AOI21_X1   g00737(.A1(new_n929_), .A2(new_n924_), .B(new_n376_), .ZN(new_n930_));
  OAI21_X1   g00738(.A1(new_n930_), .A2(new_n886_), .B(new_n928_), .ZN(new_n931_));
  OAI21_X1   g00739(.A1(new_n928_), .A2(new_n930_), .B(\asqrt[60] ), .ZN(new_n932_));
  AOI21_X1   g00740(.A1(new_n931_), .A2(new_n932_), .B(new_n229_), .ZN(new_n933_));
  AOI22_X1   g00741(.A1(new_n925_), .A2(\asqrt[58] ), .B1(new_n918_), .B2(new_n923_), .ZN(new_n934_));
  OAI22_X1   g00742(.A1(new_n934_), .A2(new_n376_), .B1(new_n927_), .B2(new_n924_), .ZN(new_n935_));
  AOI21_X1   g00743(.A1(new_n935_), .A2(\asqrt[60] ), .B(new_n898_), .ZN(new_n936_));
  NOR2_X1    g00744(.A1(new_n936_), .A2(new_n931_), .ZN(new_n937_));
  NOR4_X1    g00745(.A1(new_n937_), .A2(new_n933_), .A3(\asqrt[62] ), .A4(new_n827_), .ZN(new_n938_));
  AOI21_X1   g00746(.A1(new_n679_), .A2(new_n823_), .B(new_n825_), .ZN(new_n939_));
  XOR2_X1    g00747(.A1(new_n823_), .A2(\asqrt[63] ), .Z(new_n940_));
  NOR2_X1    g00748(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND3_X1   g00749(.A1(new_n910_), .A2(new_n938_), .A3(new_n941_), .ZN(new_n942_));
  NOR4_X1    g00750(.A1(new_n942_), .A2(new_n801_), .A3(new_n803_), .A4(new_n906_), .ZN(new_n943_));
  NOR2_X1    g00751(.A1(new_n800_), .A2(\a[108] ), .ZN(new_n944_));
  OAI21_X1   g00752(.A1(new_n943_), .A2(new_n944_), .B(new_n800_), .ZN(new_n945_));
  INV_X1     g00753(.I(new_n800_), .ZN(new_n946_));
  INV_X1     g00754(.I(new_n803_), .ZN(new_n947_));
  INV_X1     g00755(.I(new_n901_), .ZN(new_n948_));
  NOR3_X1    g00756(.A1(new_n936_), .A2(new_n931_), .A3(new_n948_), .ZN(new_n949_));
  AOI21_X1   g00757(.A1(new_n949_), .A2(new_n933_), .B(new_n828_), .ZN(new_n950_));
  INV_X1     g00758(.I(new_n905_), .ZN(new_n951_));
  AOI21_X1   g00759(.A1(new_n950_), .A2(new_n951_), .B(new_n907_), .ZN(new_n952_));
  INV_X1     g00760(.I(new_n827_), .ZN(new_n953_));
  NAND4_X1   g00761(.A1(new_n909_), .A2(new_n196_), .A3(new_n820_), .A4(new_n953_), .ZN(new_n954_));
  INV_X1     g00762(.I(new_n941_), .ZN(new_n955_));
  NOR2_X1    g00763(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  NAND4_X1   g00764(.A1(new_n956_), .A2(\a[109] ), .A3(new_n952_), .A4(new_n947_), .ZN(new_n957_));
  NAND3_X1   g00765(.A1(new_n957_), .A2(\a[108] ), .A3(new_n946_), .ZN(new_n958_));
  NAND2_X1   g00766(.A1(new_n945_), .A2(new_n958_), .ZN(new_n959_));
  INV_X1     g00767(.I(new_n797_), .ZN(new_n960_));
  NOR2_X1    g00768(.A1(new_n762_), .A2(new_n765_), .ZN(new_n961_));
  NOR2_X1    g00769(.A1(new_n942_), .A2(new_n906_), .ZN(new_n962_));
  NOR4_X1    g00770(.A1(new_n792_), .A2(new_n679_), .A3(new_n961_), .A4(new_n815_), .ZN(new_n963_));
  NOR2_X1    g00771(.A1(new_n825_), .A2(new_n794_), .ZN(new_n964_));
  XNOR2_X1   g00772(.A1(new_n964_), .A2(new_n963_), .ZN(new_n965_));
  NOR2_X1    g00773(.A1(new_n965_), .A2(new_n960_), .ZN(new_n966_));
  INV_X1     g00774(.I(new_n966_), .ZN(new_n967_));
  OAI21_X1   g00775(.A1(new_n931_), .A2(new_n936_), .B(new_n893_), .ZN(new_n968_));
  NOR4_X1    g00776(.A1(new_n968_), .A2(\asqrt[62] ), .A3(new_n907_), .A4(new_n827_), .ZN(new_n969_));
  NAND4_X1   g00777(.A1(new_n952_), .A2(new_n969_), .A3(new_n947_), .A4(new_n941_), .ZN(new_n970_));
  NOR3_X1    g00778(.A1(new_n941_), .A2(new_n947_), .A3(new_n825_), .ZN(new_n971_));
  NAND2_X1   g00779(.A1(new_n954_), .A2(new_n971_), .ZN(new_n972_));
  OAI21_X1   g00780(.A1(new_n972_), .A2(new_n952_), .B(new_n830_), .ZN(new_n973_));
  NAND3_X1   g00781(.A1(new_n973_), .A2(new_n970_), .A3(new_n831_), .ZN(new_n974_));
  NOR4_X1    g00782(.A1(new_n906_), .A2(new_n803_), .A3(new_n954_), .A4(new_n955_), .ZN(\asqrt[54] ));
  INV_X1     g00783(.I(new_n971_), .ZN(new_n976_));
  AOI21_X1   g00784(.A1(new_n910_), .A2(new_n938_), .B(new_n976_), .ZN(new_n977_));
  AOI21_X1   g00785(.A1(new_n977_), .A2(new_n906_), .B(\a[110] ), .ZN(new_n978_));
  OAI21_X1   g00786(.A1(new_n978_), .A2(new_n845_), .B(\asqrt[54] ), .ZN(new_n979_));
  NAND4_X1   g00787(.A1(new_n979_), .A2(new_n974_), .A3(new_n724_), .A4(new_n967_), .ZN(new_n980_));
  NAND2_X1   g00788(.A1(new_n980_), .A2(new_n959_), .ZN(new_n981_));
  NAND3_X1   g00789(.A1(new_n945_), .A2(new_n958_), .A3(new_n967_), .ZN(new_n982_));
  AOI21_X1   g00790(.A1(\asqrt[55] ), .A2(new_n830_), .B(\a[111] ), .ZN(new_n983_));
  NOR2_X1    g00791(.A1(new_n842_), .A2(\a[110] ), .ZN(new_n984_));
  NOR2_X1    g00792(.A1(new_n984_), .A2(new_n983_), .ZN(new_n985_));
  OAI21_X1   g00793(.A1(new_n851_), .A2(new_n833_), .B(new_n830_), .ZN(new_n986_));
  NAND2_X1   g00794(.A1(\asqrt[55] ), .A2(new_n986_), .ZN(new_n987_));
  OAI21_X1   g00795(.A1(new_n970_), .A2(new_n987_), .B(new_n985_), .ZN(new_n988_));
  INV_X1     g00796(.I(new_n985_), .ZN(new_n989_));
  INV_X1     g00797(.I(new_n987_), .ZN(new_n990_));
  NAND3_X1   g00798(.A1(\asqrt[54] ), .A2(new_n989_), .A3(new_n990_), .ZN(new_n991_));
  NAND3_X1   g00799(.A1(new_n988_), .A2(new_n991_), .A3(new_n587_), .ZN(new_n992_));
  AOI21_X1   g00800(.A1(new_n982_), .A2(\asqrt[56] ), .B(new_n992_), .ZN(new_n993_));
  NOR2_X1    g00801(.A1(new_n993_), .A2(new_n981_), .ZN(new_n994_));
  AOI22_X1   g00802(.A1(new_n959_), .A2(new_n980_), .B1(new_n982_), .B2(\asqrt[56] ), .ZN(new_n995_));
  AOI21_X1   g00803(.A1(new_n859_), .A2(new_n855_), .B(\asqrt[57] ), .ZN(new_n996_));
  AND4_X2    g00804(.A1(new_n919_), .A2(\asqrt[54] ), .A3(new_n889_), .A4(new_n996_), .Z(new_n997_));
  NOR2_X1    g00805(.A1(new_n919_), .A2(new_n587_), .ZN(new_n998_));
  NOR3_X1    g00806(.A1(new_n997_), .A2(new_n998_), .A3(\asqrt[58] ), .ZN(new_n999_));
  OAI21_X1   g00807(.A1(new_n995_), .A2(new_n587_), .B(new_n999_), .ZN(new_n1000_));
  NAND2_X1   g00808(.A1(new_n1000_), .A2(new_n994_), .ZN(new_n1001_));
  OAI22_X1   g00809(.A1(new_n995_), .A2(new_n587_), .B1(new_n981_), .B2(new_n993_), .ZN(new_n1002_));
  NAND2_X1   g00810(.A1(new_n871_), .A2(new_n868_), .ZN(new_n1003_));
  NAND4_X1   g00811(.A1(\asqrt[54] ), .A2(new_n504_), .A3(new_n1003_), .A4(new_n875_), .ZN(new_n1004_));
  XOR2_X1    g00812(.A1(new_n1004_), .A2(new_n890_), .Z(new_n1005_));
  NAND2_X1   g00813(.A1(new_n1005_), .A2(new_n376_), .ZN(new_n1006_));
  AOI21_X1   g00814(.A1(new_n1002_), .A2(\asqrt[58] ), .B(new_n1006_), .ZN(new_n1007_));
  NOR2_X1    g00815(.A1(new_n1007_), .A2(new_n1001_), .ZN(new_n1008_));
  AOI22_X1   g00816(.A1(new_n1002_), .A2(\asqrt[58] ), .B1(new_n1000_), .B2(new_n994_), .ZN(new_n1009_));
  NOR2_X1    g00817(.A1(new_n877_), .A2(new_n878_), .ZN(new_n1010_));
  NOR4_X1    g00818(.A1(new_n970_), .A2(\asqrt[59] ), .A3(new_n1010_), .A4(new_n882_), .ZN(new_n1011_));
  XOR2_X1    g00819(.A1(new_n1011_), .A2(new_n891_), .Z(new_n1012_));
  NAND2_X1   g00820(.A1(new_n1012_), .A2(new_n275_), .ZN(new_n1013_));
  INV_X1     g00821(.I(new_n1013_), .ZN(new_n1014_));
  OAI21_X1   g00822(.A1(new_n1009_), .A2(new_n376_), .B(new_n1014_), .ZN(new_n1015_));
  NAND2_X1   g00823(.A1(new_n1015_), .A2(new_n1008_), .ZN(new_n1016_));
  OAI22_X1   g00824(.A1(new_n1009_), .A2(new_n376_), .B1(new_n1007_), .B2(new_n1001_), .ZN(new_n1017_));
  NOR4_X1    g00825(.A1(new_n970_), .A2(\asqrt[60] ), .A3(new_n885_), .A4(new_n935_), .ZN(new_n1018_));
  XOR2_X1    g00826(.A1(new_n1018_), .A2(new_n932_), .Z(new_n1019_));
  NAND2_X1   g00827(.A1(new_n1019_), .A2(new_n229_), .ZN(new_n1020_));
  AOI21_X1   g00828(.A1(new_n1017_), .A2(\asqrt[60] ), .B(new_n1020_), .ZN(new_n1021_));
  AOI22_X1   g00829(.A1(new_n1017_), .A2(\asqrt[60] ), .B1(new_n1015_), .B2(new_n1008_), .ZN(new_n1022_));
  OAI22_X1   g00830(.A1(new_n1022_), .A2(new_n229_), .B1(new_n1021_), .B2(new_n1016_), .ZN(new_n1023_));
  INV_X1     g00831(.I(new_n1023_), .ZN(new_n1024_));
  NOR2_X1    g00832(.A1(new_n1024_), .A2(new_n196_), .ZN(new_n1025_));
  NOR3_X1    g00833(.A1(new_n908_), .A2(\asqrt[61] ), .A3(new_n897_), .ZN(new_n1026_));
  NAND2_X1   g00834(.A1(\asqrt[54] ), .A2(new_n1026_), .ZN(new_n1027_));
  XOR2_X1    g00835(.A1(new_n1027_), .A2(new_n933_), .Z(new_n1028_));
  INV_X1     g00836(.I(new_n1028_), .ZN(new_n1029_));
  INV_X1     g00837(.I(new_n944_), .ZN(new_n1030_));
  AOI21_X1   g00838(.A1(new_n957_), .A2(new_n1030_), .B(new_n946_), .ZN(new_n1031_));
  NOR3_X1    g00839(.A1(new_n943_), .A2(new_n794_), .A3(new_n800_), .ZN(new_n1032_));
  NOR2_X1    g00840(.A1(new_n1032_), .A2(new_n1031_), .ZN(new_n1033_));
  NOR3_X1    g00841(.A1(new_n978_), .A2(new_n845_), .A3(\asqrt[54] ), .ZN(new_n1034_));
  AOI21_X1   g00842(.A1(new_n973_), .A2(new_n831_), .B(new_n970_), .ZN(new_n1035_));
  NOR4_X1    g00843(.A1(new_n1035_), .A2(new_n1034_), .A3(\asqrt[56] ), .A4(new_n966_), .ZN(new_n1036_));
  NOR2_X1    g00844(.A1(new_n1036_), .A2(new_n1033_), .ZN(new_n1037_));
  NOR3_X1    g00845(.A1(new_n1032_), .A2(new_n1031_), .A3(new_n966_), .ZN(new_n1038_));
  AOI21_X1   g00846(.A1(\asqrt[54] ), .A2(new_n990_), .B(new_n989_), .ZN(new_n1039_));
  NOR3_X1    g00847(.A1(new_n970_), .A2(new_n985_), .A3(new_n987_), .ZN(new_n1040_));
  NOR3_X1    g00848(.A1(new_n1040_), .A2(new_n1039_), .A3(\asqrt[57] ), .ZN(new_n1041_));
  OAI21_X1   g00849(.A1(new_n1038_), .A2(new_n724_), .B(new_n1041_), .ZN(new_n1042_));
  NAND2_X1   g00850(.A1(new_n1042_), .A2(new_n1037_), .ZN(new_n1043_));
  OAI22_X1   g00851(.A1(new_n1033_), .A2(new_n1036_), .B1(new_n1038_), .B2(new_n724_), .ZN(new_n1044_));
  INV_X1     g00852(.I(new_n999_), .ZN(new_n1045_));
  AOI21_X1   g00853(.A1(new_n1044_), .A2(\asqrt[57] ), .B(new_n1045_), .ZN(new_n1046_));
  NOR2_X1    g00854(.A1(new_n1046_), .A2(new_n1043_), .ZN(new_n1047_));
  AOI22_X1   g00855(.A1(new_n1044_), .A2(\asqrt[57] ), .B1(new_n1037_), .B2(new_n1042_), .ZN(new_n1048_));
  INV_X1     g00856(.I(new_n1006_), .ZN(new_n1049_));
  OAI21_X1   g00857(.A1(new_n1048_), .A2(new_n504_), .B(new_n1049_), .ZN(new_n1050_));
  NAND2_X1   g00858(.A1(new_n1050_), .A2(new_n1047_), .ZN(new_n1051_));
  OAI22_X1   g00859(.A1(new_n1048_), .A2(new_n504_), .B1(new_n1046_), .B2(new_n1043_), .ZN(new_n1052_));
  AOI21_X1   g00860(.A1(new_n1052_), .A2(\asqrt[59] ), .B(new_n1013_), .ZN(new_n1053_));
  NOR2_X1    g00861(.A1(new_n1053_), .A2(new_n1051_), .ZN(new_n1054_));
  NAND2_X1   g00862(.A1(new_n1052_), .A2(\asqrt[59] ), .ZN(new_n1055_));
  AOI21_X1   g00863(.A1(new_n1055_), .A2(new_n1051_), .B(new_n275_), .ZN(new_n1056_));
  OAI21_X1   g00864(.A1(new_n1056_), .A2(new_n1020_), .B(new_n1054_), .ZN(new_n1057_));
  OAI21_X1   g00865(.A1(new_n1054_), .A2(new_n1056_), .B(\asqrt[61] ), .ZN(new_n1058_));
  NAND4_X1   g00866(.A1(new_n1057_), .A2(new_n1058_), .A3(new_n196_), .A4(new_n1029_), .ZN(new_n1059_));
  INV_X1     g00867(.I(new_n1059_), .ZN(new_n1060_));
  NOR2_X1    g00868(.A1(new_n909_), .A2(new_n196_), .ZN(new_n1061_));
  AND3_X2    g00869(.A1(\asqrt[54] ), .A2(new_n1061_), .A3(new_n938_), .Z(new_n1062_));
  NAND2_X1   g00870(.A1(new_n909_), .A2(new_n196_), .ZN(new_n1063_));
  NAND3_X1   g00871(.A1(new_n970_), .A2(new_n827_), .A3(new_n1063_), .ZN(new_n1064_));
  AOI21_X1   g00872(.A1(new_n1061_), .A2(new_n1064_), .B(new_n1062_), .ZN(new_n1065_));
  NOR2_X1    g00873(.A1(new_n1028_), .A2(new_n196_), .ZN(new_n1066_));
  INV_X1     g00874(.I(new_n1066_), .ZN(new_n1067_));
  AOI22_X1   g00875(.A1(new_n1052_), .A2(\asqrt[59] ), .B1(new_n1050_), .B2(new_n1047_), .ZN(new_n1068_));
  OAI22_X1   g00876(.A1(new_n1068_), .A2(new_n275_), .B1(new_n1053_), .B2(new_n1051_), .ZN(new_n1069_));
  NOR2_X1    g00877(.A1(new_n1029_), .A2(\asqrt[62] ), .ZN(new_n1070_));
  INV_X1     g00878(.I(new_n1070_), .ZN(new_n1071_));
  NAND3_X1   g00879(.A1(new_n1069_), .A2(\asqrt[61] ), .A3(new_n1071_), .ZN(new_n1072_));
  OAI21_X1   g00880(.A1(new_n1072_), .A2(new_n1057_), .B(new_n1067_), .ZN(new_n1073_));
  NOR3_X1    g00881(.A1(\asqrt[54] ), .A2(new_n820_), .A3(new_n969_), .ZN(new_n1074_));
  OAI21_X1   g00882(.A1(new_n1074_), .A2(new_n950_), .B(new_n231_), .ZN(new_n1075_));
  OAI21_X1   g00883(.A1(new_n1073_), .A2(new_n1075_), .B(new_n1065_), .ZN(new_n1076_));
  INV_X1     g00884(.I(new_n1065_), .ZN(new_n1077_));
  NOR4_X1    g00885(.A1(new_n1023_), .A2(\asqrt[62] ), .A3(new_n1077_), .A4(new_n1028_), .ZN(new_n1078_));
  AOI21_X1   g00886(.A1(new_n907_), .A2(new_n950_), .B(new_n970_), .ZN(new_n1079_));
  XOR2_X1    g00887(.A1(new_n903_), .A2(new_n231_), .Z(new_n1080_));
  NOR2_X1    g00888(.A1(new_n1079_), .A2(new_n1080_), .ZN(new_n1081_));
  NAND2_X1   g00889(.A1(new_n1078_), .A2(new_n1081_), .ZN(new_n1082_));
  NOR2_X1    g00890(.A1(new_n907_), .A2(new_n947_), .ZN(new_n1083_));
  NAND2_X1   g00891(.A1(new_n962_), .A2(new_n1083_), .ZN(new_n1084_));
  NOR3_X1    g00892(.A1(new_n1082_), .A2(new_n1076_), .A3(new_n1084_), .ZN(\asqrt[53] ));
  NAND3_X1   g00893(.A1(\asqrt[53] ), .A2(new_n1025_), .A3(new_n1060_), .ZN(new_n1086_));
  NOR2_X1    g00894(.A1(new_n1021_), .A2(new_n1016_), .ZN(new_n1087_));
  NOR3_X1    g00895(.A1(new_n1022_), .A2(new_n229_), .A3(new_n1070_), .ZN(new_n1088_));
  AOI21_X1   g00896(.A1(new_n1088_), .A2(new_n1087_), .B(new_n1066_), .ZN(new_n1089_));
  INV_X1     g00897(.I(new_n1075_), .ZN(new_n1090_));
  AOI21_X1   g00898(.A1(new_n1089_), .A2(new_n1090_), .B(new_n1077_), .ZN(new_n1091_));
  AOI21_X1   g00899(.A1(new_n1023_), .A2(\asqrt[62] ), .B(new_n1065_), .ZN(new_n1092_));
  INV_X1     g00900(.I(new_n1081_), .ZN(new_n1093_));
  NOR3_X1    g00901(.A1(new_n1092_), .A2(new_n1059_), .A3(new_n1093_), .ZN(new_n1094_));
  INV_X1     g00902(.I(new_n1084_), .ZN(new_n1095_));
  NAND3_X1   g00903(.A1(new_n1094_), .A2(new_n1091_), .A3(new_n1095_), .ZN(new_n1096_));
  AOI21_X1   g00904(.A1(new_n1024_), .A2(new_n196_), .B(new_n1029_), .ZN(new_n1097_));
  NAND2_X1   g00905(.A1(new_n1096_), .A2(new_n1097_), .ZN(new_n1098_));
  NAND2_X1   g00906(.A1(new_n1098_), .A2(new_n1025_), .ZN(new_n1099_));
  AND2_X2    g00907(.A1(new_n1099_), .A2(new_n1086_), .Z(new_n1100_));
  NOR3_X1    g00908(.A1(new_n1069_), .A2(\asqrt[61] ), .A3(new_n1019_), .ZN(new_n1101_));
  NAND2_X1   g00909(.A1(\asqrt[53] ), .A2(new_n1101_), .ZN(new_n1102_));
  XNOR2_X1   g00910(.A1(new_n1102_), .A2(new_n1058_), .ZN(new_n1103_));
  NOR2_X1    g00911(.A1(new_n1103_), .A2(new_n196_), .ZN(new_n1104_));
  INV_X1     g00912(.I(new_n1104_), .ZN(new_n1105_));
  INV_X1     g00913(.I(\a[106] ), .ZN(new_n1106_));
  NOR2_X1    g00914(.A1(\a[104] ), .A2(\a[105] ), .ZN(new_n1107_));
  AOI21_X1   g00915(.A1(new_n1106_), .A2(new_n1107_), .B(new_n947_), .ZN(new_n1108_));
  NAND2_X1   g00916(.A1(new_n962_), .A2(new_n1108_), .ZN(new_n1109_));
  XOR2_X1    g00917(.A1(new_n1109_), .A2(\a[107] ), .Z(new_n1110_));
  INV_X1     g00918(.I(\a[107] ), .ZN(new_n1111_));
  NOR4_X1    g00919(.A1(new_n1082_), .A2(new_n1076_), .A3(new_n1111_), .A4(new_n1084_), .ZN(new_n1112_));
  NOR2_X1    g00920(.A1(new_n1110_), .A2(\a[106] ), .ZN(new_n1113_));
  OAI21_X1   g00921(.A1(new_n1112_), .A2(new_n1113_), .B(new_n1110_), .ZN(new_n1114_));
  INV_X1     g00922(.I(new_n1110_), .ZN(new_n1115_));
  NAND4_X1   g00923(.A1(new_n1094_), .A2(new_n1091_), .A3(\a[107] ), .A4(new_n1095_), .ZN(new_n1116_));
  NAND3_X1   g00924(.A1(new_n1116_), .A2(\a[106] ), .A3(new_n1115_), .ZN(new_n1117_));
  NAND2_X1   g00925(.A1(new_n1114_), .A2(new_n1117_), .ZN(new_n1118_));
  INV_X1     g00926(.I(new_n1107_), .ZN(new_n1119_));
  NAND2_X1   g00927(.A1(new_n950_), .A2(new_n951_), .ZN(new_n1120_));
  NOR2_X1    g00928(.A1(new_n1082_), .A2(new_n1076_), .ZN(new_n1121_));
  NAND4_X1   g00929(.A1(new_n956_), .A2(new_n947_), .A3(new_n820_), .A4(new_n1120_), .ZN(new_n1122_));
  NOR2_X1    g00930(.A1(new_n970_), .A2(new_n1106_), .ZN(new_n1123_));
  XOR2_X1    g00931(.A1(new_n1123_), .A2(new_n1122_), .Z(new_n1124_));
  NOR2_X1    g00932(.A1(new_n1124_), .A2(new_n1119_), .ZN(new_n1125_));
  INV_X1     g00933(.I(new_n1125_), .ZN(new_n1126_));
  NOR3_X1    g00934(.A1(new_n1081_), .A2(new_n1095_), .A3(new_n970_), .ZN(new_n1127_));
  OAI21_X1   g00935(.A1(new_n1092_), .A2(new_n1059_), .B(new_n1127_), .ZN(new_n1128_));
  OAI21_X1   g00936(.A1(new_n1128_), .A2(new_n1091_), .B(new_n794_), .ZN(new_n1129_));
  NAND3_X1   g00937(.A1(new_n1129_), .A2(new_n1096_), .A3(new_n797_), .ZN(new_n1130_));
  INV_X1     g00938(.I(new_n1127_), .ZN(new_n1131_));
  NOR2_X1    g00939(.A1(new_n1078_), .A2(new_n1131_), .ZN(new_n1132_));
  AOI21_X1   g00940(.A1(new_n1132_), .A2(new_n1076_), .B(\a[108] ), .ZN(new_n1133_));
  OAI21_X1   g00941(.A1(new_n960_), .A2(new_n1133_), .B(\asqrt[53] ), .ZN(new_n1134_));
  NAND4_X1   g00942(.A1(new_n1134_), .A2(new_n1130_), .A3(new_n825_), .A4(new_n1126_), .ZN(new_n1135_));
  NAND2_X1   g00943(.A1(new_n1135_), .A2(new_n1118_), .ZN(new_n1136_));
  NAND3_X1   g00944(.A1(new_n1114_), .A2(new_n1117_), .A3(new_n1126_), .ZN(new_n1137_));
  AOI21_X1   g00945(.A1(\asqrt[54] ), .A2(new_n794_), .B(\a[109] ), .ZN(new_n1138_));
  NOR2_X1    g00946(.A1(new_n957_), .A2(\a[108] ), .ZN(new_n1139_));
  NOR2_X1    g00947(.A1(new_n1139_), .A2(new_n1138_), .ZN(new_n1140_));
  OAI21_X1   g00948(.A1(new_n967_), .A2(new_n799_), .B(new_n794_), .ZN(new_n1141_));
  NAND2_X1   g00949(.A1(\asqrt[54] ), .A2(new_n1141_), .ZN(new_n1142_));
  OAI21_X1   g00950(.A1(new_n1096_), .A2(new_n1142_), .B(new_n1140_), .ZN(new_n1143_));
  INV_X1     g00951(.I(new_n1140_), .ZN(new_n1144_));
  INV_X1     g00952(.I(new_n1142_), .ZN(new_n1145_));
  NAND3_X1   g00953(.A1(\asqrt[53] ), .A2(new_n1144_), .A3(new_n1145_), .ZN(new_n1146_));
  NAND3_X1   g00954(.A1(new_n1143_), .A2(new_n1146_), .A3(new_n724_), .ZN(new_n1147_));
  AOI21_X1   g00955(.A1(new_n1137_), .A2(\asqrt[55] ), .B(new_n1147_), .ZN(new_n1148_));
  NOR2_X1    g00956(.A1(new_n1148_), .A2(new_n1136_), .ZN(new_n1149_));
  AOI22_X1   g00957(.A1(new_n1135_), .A2(new_n1118_), .B1(new_n1137_), .B2(\asqrt[55] ), .ZN(new_n1150_));
  NOR2_X1    g00958(.A1(new_n1035_), .A2(new_n1034_), .ZN(new_n1151_));
  NOR4_X1    g00959(.A1(new_n1096_), .A2(\asqrt[56] ), .A3(new_n1151_), .A4(new_n982_), .ZN(new_n1152_));
  AOI21_X1   g00960(.A1(new_n1033_), .A2(new_n967_), .B(new_n724_), .ZN(new_n1153_));
  NOR3_X1    g00961(.A1(new_n1152_), .A2(\asqrt[57] ), .A3(new_n1153_), .ZN(new_n1154_));
  OAI21_X1   g00962(.A1(new_n1150_), .A2(new_n724_), .B(new_n1154_), .ZN(new_n1155_));
  NAND2_X1   g00963(.A1(new_n1155_), .A2(new_n1149_), .ZN(new_n1156_));
  OAI22_X1   g00964(.A1(new_n1150_), .A2(new_n724_), .B1(new_n1148_), .B2(new_n1136_), .ZN(new_n1157_));
  NAND2_X1   g00965(.A1(new_n1044_), .A2(\asqrt[57] ), .ZN(new_n1158_));
  NAND2_X1   g00966(.A1(new_n988_), .A2(new_n991_), .ZN(new_n1159_));
  NAND4_X1   g00967(.A1(\asqrt[53] ), .A2(new_n587_), .A3(new_n1159_), .A4(new_n995_), .ZN(new_n1160_));
  XNOR2_X1   g00968(.A1(new_n1160_), .A2(new_n1158_), .ZN(new_n1161_));
  NAND2_X1   g00969(.A1(new_n1161_), .A2(new_n504_), .ZN(new_n1162_));
  AOI21_X1   g00970(.A1(new_n1157_), .A2(\asqrt[57] ), .B(new_n1162_), .ZN(new_n1163_));
  NOR2_X1    g00971(.A1(new_n1163_), .A2(new_n1156_), .ZN(new_n1164_));
  AOI22_X1   g00972(.A1(new_n1157_), .A2(\asqrt[57] ), .B1(new_n1155_), .B2(new_n1149_), .ZN(new_n1165_));
  NOR2_X1    g00973(.A1(new_n997_), .A2(new_n998_), .ZN(new_n1166_));
  NOR4_X1    g00974(.A1(new_n1096_), .A2(\asqrt[58] ), .A3(new_n1166_), .A4(new_n1002_), .ZN(new_n1167_));
  AOI21_X1   g00975(.A1(new_n1158_), .A2(new_n1043_), .B(new_n504_), .ZN(new_n1168_));
  NOR2_X1    g00976(.A1(new_n1167_), .A2(new_n1168_), .ZN(new_n1169_));
  NAND2_X1   g00977(.A1(new_n1169_), .A2(new_n376_), .ZN(new_n1170_));
  INV_X1     g00978(.I(new_n1170_), .ZN(new_n1171_));
  OAI21_X1   g00979(.A1(new_n1165_), .A2(new_n504_), .B(new_n1171_), .ZN(new_n1172_));
  NAND2_X1   g00980(.A1(new_n1172_), .A2(new_n1164_), .ZN(new_n1173_));
  OAI22_X1   g00981(.A1(new_n1165_), .A2(new_n504_), .B1(new_n1163_), .B2(new_n1156_), .ZN(new_n1174_));
  NOR4_X1    g00982(.A1(new_n1096_), .A2(\asqrt[59] ), .A3(new_n1005_), .A4(new_n1052_), .ZN(new_n1175_));
  XOR2_X1    g00983(.A1(new_n1175_), .A2(new_n1055_), .Z(new_n1176_));
  NAND2_X1   g00984(.A1(new_n1176_), .A2(new_n275_), .ZN(new_n1177_));
  AOI21_X1   g00985(.A1(new_n1174_), .A2(\asqrt[59] ), .B(new_n1177_), .ZN(new_n1178_));
  NOR2_X1    g00986(.A1(new_n1178_), .A2(new_n1173_), .ZN(new_n1179_));
  AOI22_X1   g00987(.A1(new_n1174_), .A2(\asqrt[59] ), .B1(new_n1172_), .B2(new_n1164_), .ZN(new_n1180_));
  NOR4_X1    g00988(.A1(new_n1096_), .A2(\asqrt[60] ), .A3(new_n1012_), .A4(new_n1017_), .ZN(new_n1181_));
  XNOR2_X1   g00989(.A1(new_n1181_), .A2(new_n1056_), .ZN(new_n1182_));
  NAND2_X1   g00990(.A1(new_n1182_), .A2(new_n229_), .ZN(new_n1183_));
  INV_X1     g00991(.I(new_n1183_), .ZN(new_n1184_));
  OAI21_X1   g00992(.A1(new_n1180_), .A2(new_n275_), .B(new_n1184_), .ZN(new_n1185_));
  NAND2_X1   g00993(.A1(new_n1185_), .A2(new_n1179_), .ZN(new_n1186_));
  OAI22_X1   g00994(.A1(new_n1180_), .A2(new_n275_), .B1(new_n1178_), .B2(new_n1173_), .ZN(new_n1187_));
  INV_X1     g00995(.I(new_n1103_), .ZN(new_n1188_));
  NOR2_X1    g00996(.A1(new_n1188_), .A2(\asqrt[62] ), .ZN(new_n1189_));
  INV_X1     g00997(.I(new_n1189_), .ZN(new_n1190_));
  NAND3_X1   g00998(.A1(new_n1187_), .A2(\asqrt[61] ), .A3(new_n1190_), .ZN(new_n1191_));
  OAI21_X1   g00999(.A1(new_n1191_), .A2(new_n1186_), .B(new_n1105_), .ZN(new_n1192_));
  NOR3_X1    g01000(.A1(\asqrt[53] ), .A2(new_n1065_), .A3(new_n1078_), .ZN(new_n1193_));
  OAI21_X1   g01001(.A1(new_n1193_), .A2(new_n1089_), .B(new_n231_), .ZN(new_n1194_));
  OAI21_X1   g01002(.A1(new_n1192_), .A2(new_n1194_), .B(new_n1100_), .ZN(new_n1195_));
  INV_X1     g01003(.I(new_n1100_), .ZN(new_n1196_));
  AOI22_X1   g01004(.A1(new_n1187_), .A2(\asqrt[61] ), .B1(new_n1185_), .B2(new_n1179_), .ZN(new_n1197_));
  OAI21_X1   g01005(.A1(new_n1197_), .A2(new_n196_), .B(new_n1196_), .ZN(new_n1198_));
  INV_X1     g01006(.I(new_n1113_), .ZN(new_n1199_));
  AOI21_X1   g01007(.A1(new_n1116_), .A2(new_n1199_), .B(new_n1115_), .ZN(new_n1200_));
  NOR3_X1    g01008(.A1(new_n1112_), .A2(new_n1106_), .A3(new_n1110_), .ZN(new_n1201_));
  NOR2_X1    g01009(.A1(new_n1201_), .A2(new_n1200_), .ZN(new_n1202_));
  NOR3_X1    g01010(.A1(new_n1133_), .A2(\asqrt[53] ), .A3(new_n960_), .ZN(new_n1203_));
  AOI21_X1   g01011(.A1(new_n797_), .A2(new_n1129_), .B(new_n1096_), .ZN(new_n1204_));
  NOR4_X1    g01012(.A1(new_n1204_), .A2(new_n1203_), .A3(\asqrt[55] ), .A4(new_n1125_), .ZN(new_n1205_));
  NOR2_X1    g01013(.A1(new_n1205_), .A2(new_n1202_), .ZN(new_n1206_));
  NOR3_X1    g01014(.A1(new_n1201_), .A2(new_n1200_), .A3(new_n1125_), .ZN(new_n1207_));
  AOI21_X1   g01015(.A1(\asqrt[53] ), .A2(new_n1145_), .B(new_n1144_), .ZN(new_n1208_));
  NOR3_X1    g01016(.A1(new_n1096_), .A2(new_n1140_), .A3(new_n1142_), .ZN(new_n1209_));
  NOR3_X1    g01017(.A1(new_n1208_), .A2(new_n1209_), .A3(\asqrt[56] ), .ZN(new_n1210_));
  OAI21_X1   g01018(.A1(new_n1207_), .A2(new_n825_), .B(new_n1210_), .ZN(new_n1211_));
  NAND2_X1   g01019(.A1(new_n1211_), .A2(new_n1206_), .ZN(new_n1212_));
  OAI22_X1   g01020(.A1(new_n1205_), .A2(new_n1202_), .B1(new_n1207_), .B2(new_n825_), .ZN(new_n1213_));
  INV_X1     g01021(.I(new_n1154_), .ZN(new_n1214_));
  AOI21_X1   g01022(.A1(new_n1213_), .A2(\asqrt[56] ), .B(new_n1214_), .ZN(new_n1215_));
  NOR2_X1    g01023(.A1(new_n1215_), .A2(new_n1212_), .ZN(new_n1216_));
  AOI22_X1   g01024(.A1(new_n1213_), .A2(\asqrt[56] ), .B1(new_n1206_), .B2(new_n1211_), .ZN(new_n1217_));
  XOR2_X1    g01025(.A1(new_n1160_), .A2(new_n1158_), .Z(new_n1218_));
  NOR2_X1    g01026(.A1(new_n1218_), .A2(\asqrt[58] ), .ZN(new_n1219_));
  OAI21_X1   g01027(.A1(new_n1217_), .A2(new_n587_), .B(new_n1219_), .ZN(new_n1220_));
  NAND2_X1   g01028(.A1(new_n1220_), .A2(new_n1216_), .ZN(new_n1221_));
  OAI22_X1   g01029(.A1(new_n1217_), .A2(new_n587_), .B1(new_n1215_), .B2(new_n1212_), .ZN(new_n1222_));
  AOI21_X1   g01030(.A1(new_n1222_), .A2(\asqrt[58] ), .B(new_n1170_), .ZN(new_n1223_));
  NOR2_X1    g01031(.A1(new_n1223_), .A2(new_n1221_), .ZN(new_n1224_));
  AOI22_X1   g01032(.A1(new_n1222_), .A2(\asqrt[58] ), .B1(new_n1220_), .B2(new_n1216_), .ZN(new_n1225_));
  INV_X1     g01033(.I(new_n1177_), .ZN(new_n1226_));
  OAI21_X1   g01034(.A1(new_n1225_), .A2(new_n376_), .B(new_n1226_), .ZN(new_n1227_));
  NAND2_X1   g01035(.A1(new_n1227_), .A2(new_n1224_), .ZN(new_n1228_));
  NAND2_X1   g01036(.A1(new_n1222_), .A2(\asqrt[58] ), .ZN(new_n1229_));
  AOI21_X1   g01037(.A1(new_n1229_), .A2(new_n1221_), .B(new_n376_), .ZN(new_n1230_));
  OAI21_X1   g01038(.A1(new_n1224_), .A2(new_n1230_), .B(\asqrt[60] ), .ZN(new_n1231_));
  AOI21_X1   g01039(.A1(new_n1231_), .A2(new_n1184_), .B(new_n1228_), .ZN(new_n1232_));
  AOI21_X1   g01040(.A1(new_n1228_), .A2(new_n1231_), .B(new_n229_), .ZN(new_n1233_));
  NOR4_X1    g01041(.A1(new_n1232_), .A2(new_n1233_), .A3(\asqrt[62] ), .A4(new_n1103_), .ZN(new_n1234_));
  AOI21_X1   g01042(.A1(new_n1077_), .A2(new_n1089_), .B(new_n1096_), .ZN(new_n1235_));
  XOR2_X1    g01043(.A1(new_n1089_), .A2(\asqrt[63] ), .Z(new_n1236_));
  NOR2_X1    g01044(.A1(new_n1235_), .A2(new_n1236_), .ZN(new_n1237_));
  NAND3_X1   g01045(.A1(new_n1198_), .A2(new_n1234_), .A3(new_n1237_), .ZN(new_n1238_));
  NOR2_X1    g01046(.A1(new_n1238_), .A2(new_n1195_), .ZN(new_n1239_));
  INV_X1     g01047(.I(\a[102] ), .ZN(new_n1240_));
  NOR2_X1    g01048(.A1(new_n1077_), .A2(new_n1095_), .ZN(new_n1241_));
  NAND2_X1   g01049(.A1(new_n1121_), .A2(new_n1241_), .ZN(new_n1242_));
  INV_X1     g01050(.I(new_n1242_), .ZN(new_n1243_));
  NOR2_X1    g01051(.A1(\a[100] ), .A2(\a[101] ), .ZN(new_n1244_));
  AOI21_X1   g01052(.A1(new_n1240_), .A2(new_n1244_), .B(new_n1243_), .ZN(new_n1245_));
  NAND2_X1   g01053(.A1(new_n1239_), .A2(new_n1245_), .ZN(new_n1246_));
  XOR2_X1    g01054(.A1(new_n1246_), .A2(\a[103] ), .Z(new_n1247_));
  INV_X1     g01055(.I(\a[103] ), .ZN(new_n1248_));
  OAI21_X1   g01056(.A1(new_n1232_), .A2(new_n1233_), .B(\asqrt[62] ), .ZN(new_n1249_));
  INV_X1     g01057(.I(new_n1234_), .ZN(new_n1250_));
  OAI22_X1   g01058(.A1(new_n1225_), .A2(new_n376_), .B1(new_n1223_), .B2(new_n1221_), .ZN(new_n1251_));
  AOI22_X1   g01059(.A1(new_n1251_), .A2(\asqrt[60] ), .B1(new_n1227_), .B2(new_n1224_), .ZN(new_n1252_));
  NOR3_X1    g01060(.A1(new_n1252_), .A2(new_n229_), .A3(new_n1189_), .ZN(new_n1253_));
  AOI21_X1   g01061(.A1(new_n1253_), .A2(new_n1232_), .B(new_n1104_), .ZN(new_n1254_));
  INV_X1     g01062(.I(new_n1194_), .ZN(new_n1255_));
  AOI21_X1   g01063(.A1(new_n1254_), .A2(new_n1255_), .B(new_n1196_), .ZN(new_n1256_));
  NAND4_X1   g01064(.A1(new_n1197_), .A2(new_n196_), .A3(new_n1100_), .A4(new_n1188_), .ZN(new_n1257_));
  INV_X1     g01065(.I(new_n1237_), .ZN(new_n1258_));
  NOR2_X1    g01066(.A1(new_n1257_), .A2(new_n1258_), .ZN(new_n1259_));
  NAND3_X1   g01067(.A1(new_n1259_), .A2(new_n1256_), .A3(new_n1243_), .ZN(new_n1260_));
  NOR3_X1    g01068(.A1(new_n1260_), .A2(new_n1249_), .A3(new_n1250_), .ZN(new_n1261_));
  AOI21_X1   g01069(.A1(new_n1197_), .A2(new_n196_), .B(new_n1188_), .ZN(new_n1262_));
  AOI21_X1   g01070(.A1(new_n1260_), .A2(new_n1262_), .B(new_n1249_), .ZN(new_n1263_));
  NOR2_X1    g01071(.A1(new_n1261_), .A2(new_n1263_), .ZN(new_n1264_));
  NOR3_X1    g01072(.A1(new_n1238_), .A2(new_n1195_), .A3(new_n1242_), .ZN(\asqrt[52] ));
  NOR3_X1    g01073(.A1(new_n1187_), .A2(\asqrt[61] ), .A3(new_n1182_), .ZN(new_n1266_));
  NAND2_X1   g01074(.A1(\asqrt[52] ), .A2(new_n1266_), .ZN(new_n1267_));
  XOR2_X1    g01075(.A1(new_n1267_), .A2(new_n1233_), .Z(new_n1268_));
  NOR2_X1    g01076(.A1(new_n1268_), .A2(new_n196_), .ZN(new_n1269_));
  INV_X1     g01077(.I(new_n1269_), .ZN(new_n1270_));
  INV_X1     g01078(.I(\a[104] ), .ZN(new_n1271_));
  NOR2_X1    g01079(.A1(\a[102] ), .A2(\a[103] ), .ZN(new_n1272_));
  AOI21_X1   g01080(.A1(new_n1271_), .A2(new_n1272_), .B(new_n1095_), .ZN(new_n1273_));
  NAND2_X1   g01081(.A1(new_n1121_), .A2(new_n1273_), .ZN(new_n1274_));
  XOR2_X1    g01082(.A1(new_n1274_), .A2(\a[105] ), .Z(new_n1275_));
  INV_X1     g01083(.I(new_n1275_), .ZN(new_n1276_));
  NAND4_X1   g01084(.A1(new_n1259_), .A2(new_n1256_), .A3(\a[105] ), .A4(new_n1243_), .ZN(new_n1277_));
  NOR2_X1    g01085(.A1(new_n1275_), .A2(\a[104] ), .ZN(new_n1278_));
  INV_X1     g01086(.I(new_n1278_), .ZN(new_n1279_));
  AOI21_X1   g01087(.A1(new_n1277_), .A2(new_n1279_), .B(new_n1276_), .ZN(new_n1280_));
  INV_X1     g01088(.I(\a[105] ), .ZN(new_n1281_));
  NOR4_X1    g01089(.A1(new_n1238_), .A2(new_n1195_), .A3(new_n1281_), .A4(new_n1242_), .ZN(new_n1282_));
  NOR3_X1    g01090(.A1(new_n1282_), .A2(new_n1271_), .A3(new_n1275_), .ZN(new_n1283_));
  NOR2_X1    g01091(.A1(new_n1283_), .A2(new_n1280_), .ZN(new_n1284_));
  INV_X1     g01092(.I(new_n1272_), .ZN(new_n1285_));
  NOR2_X1    g01093(.A1(new_n1073_), .A2(new_n1075_), .ZN(new_n1286_));
  NOR4_X1    g01094(.A1(new_n1082_), .A2(new_n1077_), .A3(new_n1286_), .A4(new_n1084_), .ZN(new_n1287_));
  NAND2_X1   g01095(.A1(\asqrt[53] ), .A2(\a[104] ), .ZN(new_n1288_));
  XOR2_X1    g01096(.A1(new_n1288_), .A2(new_n1287_), .Z(new_n1289_));
  NOR2_X1    g01097(.A1(new_n1289_), .A2(new_n1285_), .ZN(new_n1290_));
  NOR2_X1    g01098(.A1(new_n1243_), .A2(new_n1096_), .ZN(new_n1291_));
  NAND2_X1   g01099(.A1(new_n1258_), .A2(new_n1291_), .ZN(new_n1292_));
  AOI21_X1   g01100(.A1(new_n1198_), .A2(new_n1234_), .B(new_n1292_), .ZN(new_n1293_));
  AOI21_X1   g01101(.A1(new_n1293_), .A2(new_n1195_), .B(\a[106] ), .ZN(new_n1294_));
  NOR3_X1    g01102(.A1(new_n1294_), .A2(\asqrt[52] ), .A3(new_n1119_), .ZN(new_n1295_));
  NAND3_X1   g01103(.A1(new_n1257_), .A2(new_n1258_), .A3(new_n1291_), .ZN(new_n1296_));
  OAI21_X1   g01104(.A1(new_n1296_), .A2(new_n1256_), .B(new_n1106_), .ZN(new_n1297_));
  AOI21_X1   g01105(.A1(new_n1297_), .A2(new_n1107_), .B(new_n1260_), .ZN(new_n1298_));
  NOR4_X1    g01106(.A1(new_n1298_), .A2(new_n1295_), .A3(\asqrt[54] ), .A4(new_n1290_), .ZN(new_n1299_));
  NOR2_X1    g01107(.A1(new_n1299_), .A2(new_n1284_), .ZN(new_n1300_));
  NOR3_X1    g01108(.A1(new_n1283_), .A2(new_n1280_), .A3(new_n1290_), .ZN(new_n1301_));
  AOI21_X1   g01109(.A1(\asqrt[53] ), .A2(new_n1106_), .B(\a[107] ), .ZN(new_n1302_));
  NOR2_X1    g01110(.A1(new_n1116_), .A2(\a[106] ), .ZN(new_n1303_));
  NOR2_X1    g01111(.A1(new_n1302_), .A2(new_n1303_), .ZN(new_n1304_));
  INV_X1     g01112(.I(new_n1304_), .ZN(new_n1305_));
  OAI21_X1   g01113(.A1(new_n1126_), .A2(new_n1109_), .B(new_n1106_), .ZN(new_n1306_));
  NAND2_X1   g01114(.A1(\asqrt[53] ), .A2(new_n1306_), .ZN(new_n1307_));
  INV_X1     g01115(.I(new_n1307_), .ZN(new_n1308_));
  AOI21_X1   g01116(.A1(\asqrt[52] ), .A2(new_n1308_), .B(new_n1305_), .ZN(new_n1309_));
  NOR3_X1    g01117(.A1(new_n1260_), .A2(new_n1304_), .A3(new_n1307_), .ZN(new_n1310_));
  NOR3_X1    g01118(.A1(new_n1310_), .A2(new_n1309_), .A3(\asqrt[55] ), .ZN(new_n1311_));
  OAI21_X1   g01119(.A1(new_n1301_), .A2(new_n970_), .B(new_n1311_), .ZN(new_n1312_));
  NAND2_X1   g01120(.A1(new_n1312_), .A2(new_n1300_), .ZN(new_n1313_));
  OAI22_X1   g01121(.A1(new_n1299_), .A2(new_n1284_), .B1(new_n1301_), .B2(new_n970_), .ZN(new_n1314_));
  NOR2_X1    g01122(.A1(new_n1204_), .A2(new_n1203_), .ZN(new_n1315_));
  NOR4_X1    g01123(.A1(new_n1260_), .A2(\asqrt[55] ), .A3(new_n1315_), .A4(new_n1137_), .ZN(new_n1316_));
  AOI21_X1   g01124(.A1(new_n1202_), .A2(new_n1126_), .B(new_n825_), .ZN(new_n1317_));
  NOR3_X1    g01125(.A1(new_n1316_), .A2(new_n1317_), .A3(\asqrt[56] ), .ZN(new_n1318_));
  INV_X1     g01126(.I(new_n1318_), .ZN(new_n1319_));
  AOI21_X1   g01127(.A1(new_n1314_), .A2(\asqrt[55] ), .B(new_n1319_), .ZN(new_n1320_));
  NOR2_X1    g01128(.A1(new_n1320_), .A2(new_n1313_), .ZN(new_n1321_));
  AOI22_X1   g01129(.A1(new_n1314_), .A2(\asqrt[55] ), .B1(new_n1300_), .B2(new_n1312_), .ZN(new_n1322_));
  NOR2_X1    g01130(.A1(new_n1150_), .A2(new_n724_), .ZN(new_n1323_));
  NAND2_X1   g01131(.A1(new_n1143_), .A2(new_n1146_), .ZN(new_n1324_));
  NAND4_X1   g01132(.A1(\asqrt[52] ), .A2(new_n724_), .A3(new_n1324_), .A4(new_n1150_), .ZN(new_n1325_));
  XOR2_X1    g01133(.A1(new_n1325_), .A2(new_n1323_), .Z(new_n1326_));
  NAND2_X1   g01134(.A1(new_n1326_), .A2(new_n587_), .ZN(new_n1327_));
  INV_X1     g01135(.I(new_n1327_), .ZN(new_n1328_));
  OAI21_X1   g01136(.A1(new_n1322_), .A2(new_n724_), .B(new_n1328_), .ZN(new_n1329_));
  NAND2_X1   g01137(.A1(new_n1329_), .A2(new_n1321_), .ZN(new_n1330_));
  OAI22_X1   g01138(.A1(new_n1322_), .A2(new_n724_), .B1(new_n1320_), .B2(new_n1313_), .ZN(new_n1331_));
  NOR2_X1    g01139(.A1(new_n1217_), .A2(new_n587_), .ZN(new_n1332_));
  OR2_X2     g01140(.A1(new_n1152_), .A2(new_n1153_), .Z(new_n1333_));
  NAND4_X1   g01141(.A1(\asqrt[52] ), .A2(new_n587_), .A3(new_n1333_), .A4(new_n1217_), .ZN(new_n1334_));
  XOR2_X1    g01142(.A1(new_n1334_), .A2(new_n1332_), .Z(new_n1335_));
  NAND2_X1   g01143(.A1(new_n1335_), .A2(new_n504_), .ZN(new_n1336_));
  AOI21_X1   g01144(.A1(new_n1331_), .A2(\asqrt[57] ), .B(new_n1336_), .ZN(new_n1337_));
  NOR2_X1    g01145(.A1(new_n1337_), .A2(new_n1330_), .ZN(new_n1338_));
  AOI22_X1   g01146(.A1(new_n1331_), .A2(\asqrt[57] ), .B1(new_n1329_), .B2(new_n1321_), .ZN(new_n1339_));
  NOR4_X1    g01147(.A1(new_n1260_), .A2(\asqrt[58] ), .A3(new_n1161_), .A4(new_n1222_), .ZN(new_n1340_));
  XOR2_X1    g01148(.A1(new_n1340_), .A2(new_n1229_), .Z(new_n1341_));
  NAND2_X1   g01149(.A1(new_n1341_), .A2(new_n376_), .ZN(new_n1342_));
  INV_X1     g01150(.I(new_n1342_), .ZN(new_n1343_));
  OAI21_X1   g01151(.A1(new_n1339_), .A2(new_n504_), .B(new_n1343_), .ZN(new_n1344_));
  NAND2_X1   g01152(.A1(new_n1344_), .A2(new_n1338_), .ZN(new_n1345_));
  OAI22_X1   g01153(.A1(new_n1339_), .A2(new_n504_), .B1(new_n1337_), .B2(new_n1330_), .ZN(new_n1346_));
  NOR4_X1    g01154(.A1(new_n1260_), .A2(\asqrt[59] ), .A3(new_n1169_), .A4(new_n1174_), .ZN(new_n1347_));
  XNOR2_X1   g01155(.A1(new_n1347_), .A2(new_n1230_), .ZN(new_n1348_));
  NAND2_X1   g01156(.A1(new_n1348_), .A2(new_n275_), .ZN(new_n1349_));
  AOI21_X1   g01157(.A1(new_n1346_), .A2(\asqrt[59] ), .B(new_n1349_), .ZN(new_n1350_));
  NOR2_X1    g01158(.A1(new_n1350_), .A2(new_n1345_), .ZN(new_n1351_));
  AOI22_X1   g01159(.A1(new_n1346_), .A2(\asqrt[59] ), .B1(new_n1344_), .B2(new_n1338_), .ZN(new_n1352_));
  NOR4_X1    g01160(.A1(new_n1260_), .A2(\asqrt[60] ), .A3(new_n1176_), .A4(new_n1251_), .ZN(new_n1353_));
  XOR2_X1    g01161(.A1(new_n1353_), .A2(new_n1231_), .Z(new_n1354_));
  NAND2_X1   g01162(.A1(new_n1354_), .A2(new_n229_), .ZN(new_n1355_));
  INV_X1     g01163(.I(new_n1355_), .ZN(new_n1356_));
  OAI21_X1   g01164(.A1(new_n1352_), .A2(new_n275_), .B(new_n1356_), .ZN(new_n1357_));
  NAND2_X1   g01165(.A1(new_n1357_), .A2(new_n1351_), .ZN(new_n1358_));
  OAI22_X1   g01166(.A1(new_n1352_), .A2(new_n275_), .B1(new_n1350_), .B2(new_n1345_), .ZN(new_n1359_));
  INV_X1     g01167(.I(new_n1268_), .ZN(new_n1360_));
  NOR2_X1    g01168(.A1(new_n1360_), .A2(\asqrt[62] ), .ZN(new_n1361_));
  INV_X1     g01169(.I(new_n1361_), .ZN(new_n1362_));
  NAND3_X1   g01170(.A1(new_n1359_), .A2(\asqrt[61] ), .A3(new_n1362_), .ZN(new_n1363_));
  OAI21_X1   g01171(.A1(new_n1363_), .A2(new_n1358_), .B(new_n1270_), .ZN(new_n1364_));
  AOI21_X1   g01172(.A1(new_n1198_), .A2(new_n1234_), .B(new_n1100_), .ZN(new_n1365_));
  AOI21_X1   g01173(.A1(new_n1260_), .A2(new_n1365_), .B(new_n1254_), .ZN(new_n1366_));
  NOR2_X1    g01174(.A1(new_n1366_), .A2(\asqrt[63] ), .ZN(new_n1367_));
  INV_X1     g01175(.I(new_n1367_), .ZN(new_n1368_));
  OAI21_X1   g01176(.A1(new_n1364_), .A2(new_n1368_), .B(new_n1264_), .ZN(new_n1369_));
  OAI21_X1   g01177(.A1(new_n1100_), .A2(new_n1192_), .B(\asqrt[52] ), .ZN(new_n1370_));
  XOR2_X1    g01178(.A1(new_n1192_), .A2(\asqrt[63] ), .Z(new_n1371_));
  NAND2_X1   g01179(.A1(new_n1370_), .A2(new_n1371_), .ZN(new_n1372_));
  INV_X1     g01180(.I(new_n1372_), .ZN(new_n1373_));
  INV_X1     g01181(.I(new_n1264_), .ZN(new_n1374_));
  OAI21_X1   g01182(.A1(new_n1282_), .A2(new_n1278_), .B(new_n1275_), .ZN(new_n1375_));
  NAND3_X1   g01183(.A1(new_n1277_), .A2(\a[104] ), .A3(new_n1276_), .ZN(new_n1376_));
  NAND2_X1   g01184(.A1(new_n1375_), .A2(new_n1376_), .ZN(new_n1377_));
  INV_X1     g01185(.I(new_n1290_), .ZN(new_n1378_));
  NAND3_X1   g01186(.A1(new_n1297_), .A2(new_n1260_), .A3(new_n1107_), .ZN(new_n1379_));
  OAI21_X1   g01187(.A1(new_n1119_), .A2(new_n1294_), .B(\asqrt[52] ), .ZN(new_n1380_));
  NAND4_X1   g01188(.A1(new_n1380_), .A2(new_n1379_), .A3(new_n970_), .A4(new_n1378_), .ZN(new_n1381_));
  NAND2_X1   g01189(.A1(new_n1381_), .A2(new_n1377_), .ZN(new_n1382_));
  NAND3_X1   g01190(.A1(new_n1375_), .A2(new_n1376_), .A3(new_n1378_), .ZN(new_n1383_));
  OAI21_X1   g01191(.A1(new_n1260_), .A2(new_n1307_), .B(new_n1304_), .ZN(new_n1384_));
  NAND4_X1   g01192(.A1(new_n1239_), .A2(new_n1243_), .A3(new_n1305_), .A4(new_n1308_), .ZN(new_n1385_));
  NAND3_X1   g01193(.A1(new_n1384_), .A2(new_n1385_), .A3(new_n825_), .ZN(new_n1386_));
  AOI21_X1   g01194(.A1(new_n1383_), .A2(\asqrt[54] ), .B(new_n1386_), .ZN(new_n1387_));
  NOR2_X1    g01195(.A1(new_n1387_), .A2(new_n1382_), .ZN(new_n1388_));
  AOI22_X1   g01196(.A1(new_n1381_), .A2(new_n1377_), .B1(new_n1383_), .B2(\asqrt[54] ), .ZN(new_n1389_));
  OAI21_X1   g01197(.A1(new_n1389_), .A2(new_n825_), .B(new_n1318_), .ZN(new_n1390_));
  NAND2_X1   g01198(.A1(new_n1390_), .A2(new_n1388_), .ZN(new_n1391_));
  OAI22_X1   g01199(.A1(new_n1389_), .A2(new_n825_), .B1(new_n1382_), .B2(new_n1387_), .ZN(new_n1392_));
  AOI21_X1   g01200(.A1(new_n1392_), .A2(\asqrt[56] ), .B(new_n1327_), .ZN(new_n1393_));
  NOR2_X1    g01201(.A1(new_n1393_), .A2(new_n1391_), .ZN(new_n1394_));
  AOI22_X1   g01202(.A1(new_n1392_), .A2(\asqrt[56] ), .B1(new_n1390_), .B2(new_n1388_), .ZN(new_n1395_));
  INV_X1     g01203(.I(new_n1336_), .ZN(new_n1396_));
  OAI21_X1   g01204(.A1(new_n1395_), .A2(new_n587_), .B(new_n1396_), .ZN(new_n1397_));
  NAND2_X1   g01205(.A1(new_n1397_), .A2(new_n1394_), .ZN(new_n1398_));
  OAI22_X1   g01206(.A1(new_n1395_), .A2(new_n587_), .B1(new_n1393_), .B2(new_n1391_), .ZN(new_n1399_));
  AOI21_X1   g01207(.A1(new_n1399_), .A2(\asqrt[58] ), .B(new_n1342_), .ZN(new_n1400_));
  NOR2_X1    g01208(.A1(new_n1400_), .A2(new_n1398_), .ZN(new_n1401_));
  AOI22_X1   g01209(.A1(new_n1399_), .A2(\asqrt[58] ), .B1(new_n1397_), .B2(new_n1394_), .ZN(new_n1402_));
  INV_X1     g01210(.I(new_n1349_), .ZN(new_n1403_));
  OAI21_X1   g01211(.A1(new_n1402_), .A2(new_n376_), .B(new_n1403_), .ZN(new_n1404_));
  NAND2_X1   g01212(.A1(new_n1404_), .A2(new_n1401_), .ZN(new_n1405_));
  OAI22_X1   g01213(.A1(new_n1402_), .A2(new_n376_), .B1(new_n1400_), .B2(new_n1398_), .ZN(new_n1406_));
  AOI21_X1   g01214(.A1(new_n1406_), .A2(\asqrt[60] ), .B(new_n1355_), .ZN(new_n1407_));
  AOI22_X1   g01215(.A1(new_n1406_), .A2(\asqrt[60] ), .B1(new_n1404_), .B2(new_n1401_), .ZN(new_n1408_));
  OAI22_X1   g01216(.A1(new_n1408_), .A2(new_n229_), .B1(new_n1407_), .B2(new_n1405_), .ZN(new_n1409_));
  NOR4_X1    g01217(.A1(new_n1409_), .A2(\asqrt[62] ), .A3(new_n1374_), .A4(new_n1268_), .ZN(new_n1410_));
  NAND2_X1   g01218(.A1(new_n1410_), .A2(new_n1373_), .ZN(new_n1411_));
  NAND3_X1   g01219(.A1(new_n1239_), .A2(new_n1242_), .A3(new_n1100_), .ZN(new_n1412_));
  NOR4_X1    g01220(.A1(new_n1411_), .A2(new_n1369_), .A3(new_n1248_), .A4(new_n1412_), .ZN(new_n1413_));
  NOR2_X1    g01221(.A1(new_n1247_), .A2(\a[102] ), .ZN(new_n1414_));
  OAI21_X1   g01222(.A1(new_n1413_), .A2(new_n1414_), .B(new_n1247_), .ZN(new_n1415_));
  INV_X1     g01223(.I(new_n1247_), .ZN(new_n1416_));
  NOR2_X1    g01224(.A1(new_n1407_), .A2(new_n1405_), .ZN(new_n1417_));
  NOR3_X1    g01225(.A1(new_n1408_), .A2(new_n229_), .A3(new_n1361_), .ZN(new_n1418_));
  AOI21_X1   g01226(.A1(new_n1418_), .A2(new_n1417_), .B(new_n1269_), .ZN(new_n1419_));
  AOI21_X1   g01227(.A1(new_n1419_), .A2(new_n1367_), .B(new_n1374_), .ZN(new_n1420_));
  AOI22_X1   g01228(.A1(new_n1359_), .A2(\asqrt[61] ), .B1(new_n1357_), .B2(new_n1351_), .ZN(new_n1421_));
  NAND4_X1   g01229(.A1(new_n1421_), .A2(new_n196_), .A3(new_n1264_), .A4(new_n1360_), .ZN(new_n1422_));
  NOR2_X1    g01230(.A1(new_n1422_), .A2(new_n1372_), .ZN(new_n1423_));
  INV_X1     g01231(.I(new_n1412_), .ZN(new_n1424_));
  NAND4_X1   g01232(.A1(new_n1423_), .A2(\a[103] ), .A3(new_n1420_), .A4(new_n1424_), .ZN(new_n1425_));
  NAND3_X1   g01233(.A1(new_n1425_), .A2(\a[102] ), .A3(new_n1416_), .ZN(new_n1426_));
  NAND2_X1   g01234(.A1(new_n1415_), .A2(new_n1426_), .ZN(new_n1427_));
  INV_X1     g01235(.I(new_n1244_), .ZN(new_n1428_));
  NAND2_X1   g01236(.A1(new_n1254_), .A2(new_n1255_), .ZN(new_n1429_));
  NOR2_X1    g01237(.A1(new_n1411_), .A2(new_n1369_), .ZN(new_n1430_));
  NAND4_X1   g01238(.A1(new_n1259_), .A2(new_n1243_), .A3(new_n1429_), .A4(new_n1100_), .ZN(new_n1431_));
  NOR2_X1    g01239(.A1(new_n1260_), .A2(new_n1240_), .ZN(new_n1432_));
  XOR2_X1    g01240(.A1(new_n1432_), .A2(new_n1431_), .Z(new_n1433_));
  NOR2_X1    g01241(.A1(new_n1433_), .A2(new_n1428_), .ZN(new_n1434_));
  INV_X1     g01242(.I(new_n1434_), .ZN(new_n1435_));
  NAND3_X1   g01243(.A1(new_n1423_), .A2(new_n1420_), .A3(new_n1424_), .ZN(new_n1436_));
  NAND2_X1   g01244(.A1(new_n1314_), .A2(\asqrt[55] ), .ZN(new_n1437_));
  AOI21_X1   g01245(.A1(new_n1437_), .A2(new_n1313_), .B(new_n724_), .ZN(new_n1438_));
  OAI21_X1   g01246(.A1(new_n1321_), .A2(new_n1438_), .B(\asqrt[57] ), .ZN(new_n1439_));
  AOI21_X1   g01247(.A1(new_n1330_), .A2(new_n1439_), .B(new_n504_), .ZN(new_n1440_));
  OAI21_X1   g01248(.A1(new_n1338_), .A2(new_n1440_), .B(\asqrt[59] ), .ZN(new_n1441_));
  AOI21_X1   g01249(.A1(new_n1345_), .A2(new_n1441_), .B(new_n275_), .ZN(new_n1442_));
  OAI21_X1   g01250(.A1(new_n1351_), .A2(new_n1442_), .B(\asqrt[61] ), .ZN(new_n1443_));
  NOR3_X1    g01251(.A1(new_n1358_), .A2(new_n1443_), .A3(new_n1361_), .ZN(new_n1444_));
  NOR3_X1    g01252(.A1(new_n1444_), .A2(new_n1269_), .A3(new_n1368_), .ZN(new_n1445_));
  OAI21_X1   g01253(.A1(new_n1445_), .A2(new_n1374_), .B(new_n1422_), .ZN(new_n1446_));
  NOR2_X1    g01254(.A1(new_n1373_), .A2(new_n1424_), .ZN(new_n1447_));
  NAND2_X1   g01255(.A1(new_n1447_), .A2(\asqrt[52] ), .ZN(new_n1448_));
  OAI21_X1   g01256(.A1(new_n1446_), .A2(new_n1448_), .B(new_n1271_), .ZN(new_n1449_));
  NAND3_X1   g01257(.A1(new_n1449_), .A2(new_n1272_), .A3(new_n1436_), .ZN(new_n1450_));
  NOR3_X1    g01258(.A1(new_n1411_), .A2(new_n1369_), .A3(new_n1412_), .ZN(\asqrt[51] ));
  NAND2_X1   g01259(.A1(new_n1392_), .A2(\asqrt[56] ), .ZN(new_n1452_));
  AOI21_X1   g01260(.A1(new_n1452_), .A2(new_n1391_), .B(new_n587_), .ZN(new_n1453_));
  OAI21_X1   g01261(.A1(new_n1394_), .A2(new_n1453_), .B(\asqrt[58] ), .ZN(new_n1454_));
  AOI21_X1   g01262(.A1(new_n1398_), .A2(new_n1454_), .B(new_n376_), .ZN(new_n1455_));
  OAI21_X1   g01263(.A1(new_n1401_), .A2(new_n1455_), .B(\asqrt[60] ), .ZN(new_n1456_));
  AOI21_X1   g01264(.A1(new_n1405_), .A2(new_n1456_), .B(new_n229_), .ZN(new_n1457_));
  NAND3_X1   g01265(.A1(new_n1417_), .A2(new_n1457_), .A3(new_n1362_), .ZN(new_n1458_));
  NAND3_X1   g01266(.A1(new_n1458_), .A2(new_n1270_), .A3(new_n1367_), .ZN(new_n1459_));
  AOI21_X1   g01267(.A1(new_n1459_), .A2(new_n1264_), .B(new_n1410_), .ZN(new_n1460_));
  INV_X1     g01268(.I(new_n1448_), .ZN(new_n1461_));
  AOI21_X1   g01269(.A1(new_n1460_), .A2(new_n1461_), .B(\a[104] ), .ZN(new_n1462_));
  OAI21_X1   g01270(.A1(new_n1462_), .A2(new_n1285_), .B(\asqrt[51] ), .ZN(new_n1463_));
  NAND4_X1   g01271(.A1(new_n1450_), .A2(new_n1463_), .A3(new_n1096_), .A4(new_n1435_), .ZN(new_n1464_));
  INV_X1     g01272(.I(new_n1414_), .ZN(new_n1465_));
  AOI21_X1   g01273(.A1(new_n1425_), .A2(new_n1465_), .B(new_n1416_), .ZN(new_n1466_));
  NOR3_X1    g01274(.A1(new_n1413_), .A2(new_n1240_), .A3(new_n1247_), .ZN(new_n1467_));
  NOR3_X1    g01275(.A1(new_n1466_), .A2(new_n1467_), .A3(new_n1434_), .ZN(new_n1468_));
  NAND2_X1   g01276(.A1(\asqrt[52] ), .A2(new_n1271_), .ZN(new_n1469_));
  AOI22_X1   g01277(.A1(new_n1469_), .A2(new_n1281_), .B1(new_n1271_), .B2(new_n1282_), .ZN(new_n1470_));
  INV_X1     g01278(.I(new_n1470_), .ZN(new_n1471_));
  OAI21_X1   g01279(.A1(new_n1378_), .A2(new_n1274_), .B(new_n1271_), .ZN(new_n1472_));
  NAND2_X1   g01280(.A1(\asqrt[52] ), .A2(new_n1472_), .ZN(new_n1473_));
  INV_X1     g01281(.I(new_n1473_), .ZN(new_n1474_));
  AOI21_X1   g01282(.A1(\asqrt[51] ), .A2(new_n1474_), .B(new_n1471_), .ZN(new_n1475_));
  NOR2_X1    g01283(.A1(new_n1470_), .A2(new_n1473_), .ZN(new_n1476_));
  INV_X1     g01284(.I(new_n1476_), .ZN(new_n1477_));
  NOR2_X1    g01285(.A1(new_n1436_), .A2(new_n1477_), .ZN(new_n1478_));
  NOR3_X1    g01286(.A1(new_n1475_), .A2(new_n1478_), .A3(\asqrt[54] ), .ZN(new_n1479_));
  OAI21_X1   g01287(.A1(new_n1468_), .A2(new_n1096_), .B(new_n1479_), .ZN(new_n1480_));
  NAND3_X1   g01288(.A1(new_n1480_), .A2(new_n1427_), .A3(new_n1464_), .ZN(new_n1481_));
  NOR2_X1    g01289(.A1(new_n1466_), .A2(new_n1467_), .ZN(new_n1482_));
  NOR3_X1    g01290(.A1(new_n1462_), .A2(new_n1285_), .A3(\asqrt[51] ), .ZN(new_n1483_));
  AOI21_X1   g01291(.A1(new_n1449_), .A2(new_n1272_), .B(new_n1436_), .ZN(new_n1484_));
  NOR3_X1    g01292(.A1(new_n1484_), .A2(new_n1483_), .A3(\asqrt[53] ), .ZN(new_n1485_));
  AOI21_X1   g01293(.A1(new_n1485_), .A2(new_n1435_), .B(new_n1482_), .ZN(new_n1486_));
  NOR2_X1    g01294(.A1(new_n1468_), .A2(new_n1096_), .ZN(new_n1487_));
  OAI21_X1   g01295(.A1(new_n1486_), .A2(new_n1487_), .B(\asqrt[54] ), .ZN(new_n1488_));
  NOR2_X1    g01296(.A1(new_n1298_), .A2(new_n1295_), .ZN(new_n1489_));
  NOR4_X1    g01297(.A1(new_n1436_), .A2(\asqrt[54] ), .A3(new_n1489_), .A4(new_n1383_), .ZN(new_n1490_));
  AOI21_X1   g01298(.A1(new_n1284_), .A2(new_n1378_), .B(new_n970_), .ZN(new_n1491_));
  NOR3_X1    g01299(.A1(new_n1490_), .A2(\asqrt[55] ), .A3(new_n1491_), .ZN(new_n1492_));
  AOI21_X1   g01300(.A1(new_n1488_), .A2(new_n1492_), .B(new_n1481_), .ZN(new_n1493_));
  AOI21_X1   g01301(.A1(new_n1488_), .A2(new_n1481_), .B(new_n825_), .ZN(new_n1494_));
  NAND2_X1   g01302(.A1(new_n1384_), .A2(new_n1385_), .ZN(new_n1495_));
  NAND4_X1   g01303(.A1(\asqrt[51] ), .A2(new_n825_), .A3(new_n1495_), .A4(new_n1389_), .ZN(new_n1496_));
  XNOR2_X1   g01304(.A1(new_n1496_), .A2(new_n1437_), .ZN(new_n1497_));
  NAND2_X1   g01305(.A1(new_n1497_), .A2(new_n724_), .ZN(new_n1498_));
  OAI21_X1   g01306(.A1(new_n1494_), .A2(new_n1498_), .B(new_n1493_), .ZN(new_n1499_));
  OAI21_X1   g01307(.A1(new_n1493_), .A2(new_n1494_), .B(\asqrt[56] ), .ZN(new_n1500_));
  NOR2_X1    g01308(.A1(new_n1316_), .A2(new_n1317_), .ZN(new_n1501_));
  NOR4_X1    g01309(.A1(new_n1436_), .A2(\asqrt[56] ), .A3(new_n1501_), .A4(new_n1392_), .ZN(new_n1502_));
  XOR2_X1    g01310(.A1(new_n1502_), .A2(new_n1452_), .Z(new_n1503_));
  AND2_X2    g01311(.A1(new_n1503_), .A2(new_n587_), .Z(new_n1504_));
  AOI21_X1   g01312(.A1(new_n1500_), .A2(new_n1504_), .B(new_n1499_), .ZN(new_n1505_));
  AOI21_X1   g01313(.A1(new_n1499_), .A2(new_n1500_), .B(new_n587_), .ZN(new_n1506_));
  NOR4_X1    g01314(.A1(new_n1436_), .A2(\asqrt[57] ), .A3(new_n1326_), .A4(new_n1331_), .ZN(new_n1507_));
  XOR2_X1    g01315(.A1(new_n1507_), .A2(new_n1439_), .Z(new_n1508_));
  NAND2_X1   g01316(.A1(new_n1508_), .A2(new_n504_), .ZN(new_n1509_));
  OAI21_X1   g01317(.A1(new_n1506_), .A2(new_n1509_), .B(new_n1505_), .ZN(new_n1510_));
  OAI21_X1   g01318(.A1(new_n1505_), .A2(new_n1506_), .B(\asqrt[58] ), .ZN(new_n1511_));
  NOR4_X1    g01319(.A1(new_n1436_), .A2(\asqrt[58] ), .A3(new_n1335_), .A4(new_n1399_), .ZN(new_n1512_));
  XOR2_X1    g01320(.A1(new_n1512_), .A2(new_n1454_), .Z(new_n1513_));
  NAND2_X1   g01321(.A1(new_n1513_), .A2(new_n376_), .ZN(new_n1514_));
  INV_X1     g01322(.I(new_n1514_), .ZN(new_n1515_));
  AOI21_X1   g01323(.A1(new_n1511_), .A2(new_n1515_), .B(new_n1510_), .ZN(new_n1516_));
  AOI21_X1   g01324(.A1(new_n1510_), .A2(new_n1511_), .B(new_n376_), .ZN(new_n1517_));
  NOR4_X1    g01325(.A1(new_n1436_), .A2(\asqrt[59] ), .A3(new_n1341_), .A4(new_n1346_), .ZN(new_n1518_));
  XOR2_X1    g01326(.A1(new_n1518_), .A2(new_n1441_), .Z(new_n1519_));
  NAND2_X1   g01327(.A1(new_n1519_), .A2(new_n275_), .ZN(new_n1520_));
  OAI21_X1   g01328(.A1(new_n1517_), .A2(new_n1520_), .B(new_n1516_), .ZN(new_n1521_));
  OAI21_X1   g01329(.A1(new_n1516_), .A2(new_n1517_), .B(\asqrt[60] ), .ZN(new_n1522_));
  AOI21_X1   g01330(.A1(new_n1521_), .A2(new_n1522_), .B(new_n229_), .ZN(new_n1523_));
  NAND2_X1   g01331(.A1(new_n1464_), .A2(new_n1427_), .ZN(new_n1524_));
  NAND3_X1   g01332(.A1(new_n1415_), .A2(new_n1426_), .A3(new_n1435_), .ZN(new_n1525_));
  OAI21_X1   g01333(.A1(new_n1436_), .A2(new_n1473_), .B(new_n1470_), .ZN(new_n1526_));
  NAND2_X1   g01334(.A1(\asqrt[51] ), .A2(new_n1476_), .ZN(new_n1527_));
  NAND3_X1   g01335(.A1(new_n1526_), .A2(new_n1527_), .A3(new_n970_), .ZN(new_n1528_));
  AOI21_X1   g01336(.A1(new_n1525_), .A2(\asqrt[53] ), .B(new_n1528_), .ZN(new_n1529_));
  NOR2_X1    g01337(.A1(new_n1524_), .A2(new_n1529_), .ZN(new_n1530_));
  AOI22_X1   g01338(.A1(new_n1464_), .A2(new_n1427_), .B1(\asqrt[53] ), .B2(new_n1525_), .ZN(new_n1531_));
  OAI21_X1   g01339(.A1(new_n1531_), .A2(new_n970_), .B(new_n1492_), .ZN(new_n1532_));
  NAND2_X1   g01340(.A1(new_n1532_), .A2(new_n1530_), .ZN(new_n1533_));
  OAI22_X1   g01341(.A1(new_n1531_), .A2(new_n970_), .B1(new_n1524_), .B2(new_n1529_), .ZN(new_n1534_));
  AOI21_X1   g01342(.A1(new_n1534_), .A2(\asqrt[55] ), .B(new_n1498_), .ZN(new_n1535_));
  NOR2_X1    g01343(.A1(new_n1535_), .A2(new_n1533_), .ZN(new_n1536_));
  AOI22_X1   g01344(.A1(new_n1534_), .A2(\asqrt[55] ), .B1(new_n1532_), .B2(new_n1530_), .ZN(new_n1537_));
  OAI21_X1   g01345(.A1(new_n1537_), .A2(new_n724_), .B(new_n1504_), .ZN(new_n1538_));
  NAND2_X1   g01346(.A1(new_n1538_), .A2(new_n1536_), .ZN(new_n1539_));
  OAI22_X1   g01347(.A1(new_n1537_), .A2(new_n724_), .B1(new_n1535_), .B2(new_n1533_), .ZN(new_n1540_));
  AOI21_X1   g01348(.A1(new_n1540_), .A2(\asqrt[57] ), .B(new_n1509_), .ZN(new_n1541_));
  NOR2_X1    g01349(.A1(new_n1541_), .A2(new_n1539_), .ZN(new_n1542_));
  AOI22_X1   g01350(.A1(new_n1540_), .A2(\asqrt[57] ), .B1(new_n1538_), .B2(new_n1536_), .ZN(new_n1543_));
  OAI21_X1   g01351(.A1(new_n1543_), .A2(new_n504_), .B(new_n1515_), .ZN(new_n1544_));
  NAND2_X1   g01352(.A1(new_n1544_), .A2(new_n1542_), .ZN(new_n1545_));
  NOR2_X1    g01353(.A1(new_n1531_), .A2(new_n970_), .ZN(new_n1546_));
  OAI21_X1   g01354(.A1(new_n1546_), .A2(new_n1530_), .B(\asqrt[55] ), .ZN(new_n1547_));
  AOI21_X1   g01355(.A1(new_n1547_), .A2(new_n1533_), .B(new_n724_), .ZN(new_n1548_));
  OAI21_X1   g01356(.A1(new_n1536_), .A2(new_n1548_), .B(\asqrt[57] ), .ZN(new_n1549_));
  AOI21_X1   g01357(.A1(new_n1539_), .A2(new_n1549_), .B(new_n504_), .ZN(new_n1550_));
  OAI21_X1   g01358(.A1(new_n1542_), .A2(new_n1550_), .B(\asqrt[59] ), .ZN(new_n1551_));
  AOI21_X1   g01359(.A1(new_n1545_), .A2(new_n1551_), .B(new_n275_), .ZN(new_n1552_));
  NOR4_X1    g01360(.A1(new_n1436_), .A2(\asqrt[60] ), .A3(new_n1348_), .A4(new_n1406_), .ZN(new_n1553_));
  XOR2_X1    g01361(.A1(new_n1553_), .A2(new_n1456_), .Z(new_n1554_));
  NAND2_X1   g01362(.A1(new_n1554_), .A2(new_n229_), .ZN(new_n1555_));
  NOR2_X1    g01363(.A1(new_n1552_), .A2(new_n1555_), .ZN(new_n1556_));
  NOR2_X1    g01364(.A1(new_n1556_), .A2(new_n1521_), .ZN(new_n1557_));
  OAI21_X1   g01365(.A1(new_n1557_), .A2(new_n1523_), .B(\asqrt[62] ), .ZN(new_n1558_));
  NOR3_X1    g01366(.A1(new_n1359_), .A2(\asqrt[61] ), .A3(new_n1354_), .ZN(new_n1559_));
  NAND2_X1   g01367(.A1(\asqrt[51] ), .A2(new_n1559_), .ZN(new_n1560_));
  XOR2_X1    g01368(.A1(new_n1560_), .A2(new_n1457_), .Z(new_n1561_));
  NOR4_X1    g01369(.A1(new_n1557_), .A2(\asqrt[62] ), .A3(new_n1561_), .A4(new_n1523_), .ZN(new_n1562_));
  INV_X1     g01370(.I(new_n1562_), .ZN(new_n1563_));
  NAND3_X1   g01371(.A1(new_n1430_), .A2(new_n1264_), .A3(new_n1412_), .ZN(new_n1564_));
  INV_X1     g01372(.I(new_n1564_), .ZN(new_n1565_));
  NOR2_X1    g01373(.A1(new_n1421_), .A2(new_n196_), .ZN(new_n1566_));
  INV_X1     g01374(.I(new_n1566_), .ZN(new_n1567_));
  NOR2_X1    g01375(.A1(new_n1409_), .A2(\asqrt[62] ), .ZN(new_n1568_));
  NAND4_X1   g01376(.A1(\asqrt[51] ), .A2(new_n1360_), .A3(new_n1566_), .A4(new_n1568_), .ZN(new_n1569_));
  NOR3_X1    g01377(.A1(\asqrt[51] ), .A2(new_n1360_), .A3(new_n1568_), .ZN(new_n1570_));
  OAI21_X1   g01378(.A1(new_n1567_), .A2(new_n1570_), .B(new_n1569_), .ZN(new_n1571_));
  NOR2_X1    g01379(.A1(new_n1561_), .A2(new_n196_), .ZN(new_n1572_));
  INV_X1     g01380(.I(new_n1561_), .ZN(new_n1573_));
  NOR2_X1    g01381(.A1(new_n1573_), .A2(\asqrt[62] ), .ZN(new_n1574_));
  NOR3_X1    g01382(.A1(new_n1556_), .A2(new_n1521_), .A3(new_n1574_), .ZN(new_n1575_));
  AOI21_X1   g01383(.A1(new_n1575_), .A2(new_n1523_), .B(new_n1572_), .ZN(new_n1576_));
  NAND3_X1   g01384(.A1(new_n1436_), .A2(new_n1374_), .A3(new_n1422_), .ZN(new_n1577_));
  AOI21_X1   g01385(.A1(new_n1577_), .A2(new_n1364_), .B(\asqrt[63] ), .ZN(new_n1578_));
  AOI21_X1   g01386(.A1(new_n1576_), .A2(new_n1578_), .B(new_n1571_), .ZN(new_n1579_));
  INV_X1     g01387(.I(new_n1571_), .ZN(new_n1580_));
  OAI22_X1   g01388(.A1(new_n1543_), .A2(new_n504_), .B1(new_n1541_), .B2(new_n1539_), .ZN(new_n1581_));
  AOI21_X1   g01389(.A1(new_n1581_), .A2(\asqrt[59] ), .B(new_n1520_), .ZN(new_n1582_));
  NOR2_X1    g01390(.A1(new_n1582_), .A2(new_n1545_), .ZN(new_n1583_));
  AOI22_X1   g01391(.A1(new_n1581_), .A2(\asqrt[59] ), .B1(new_n1544_), .B2(new_n1542_), .ZN(new_n1584_));
  OAI22_X1   g01392(.A1(new_n1584_), .A2(new_n275_), .B1(new_n1582_), .B2(new_n1545_), .ZN(new_n1585_));
  INV_X1     g01393(.I(new_n1555_), .ZN(new_n1586_));
  OAI21_X1   g01394(.A1(new_n1584_), .A2(new_n275_), .B(new_n1586_), .ZN(new_n1587_));
  AOI22_X1   g01395(.A1(new_n1585_), .A2(\asqrt[61] ), .B1(new_n1587_), .B2(new_n1583_), .ZN(new_n1588_));
  NAND4_X1   g01396(.A1(new_n1588_), .A2(new_n196_), .A3(new_n1580_), .A4(new_n1573_), .ZN(new_n1589_));
  NAND2_X1   g01397(.A1(new_n1419_), .A2(new_n1374_), .ZN(new_n1590_));
  XOR2_X1    g01398(.A1(new_n1419_), .A2(\asqrt[63] ), .Z(new_n1591_));
  AOI21_X1   g01399(.A1(\asqrt[51] ), .A2(new_n1590_), .B(new_n1591_), .ZN(new_n1592_));
  INV_X1     g01400(.I(new_n1592_), .ZN(new_n1593_));
  NOR2_X1    g01401(.A1(new_n1589_), .A2(new_n1593_), .ZN(new_n1594_));
  NAND3_X1   g01402(.A1(new_n1594_), .A2(new_n1579_), .A3(new_n1565_), .ZN(new_n1595_));
  NOR3_X1    g01403(.A1(new_n1595_), .A2(new_n1558_), .A3(new_n1563_), .ZN(new_n1596_));
  AOI21_X1   g01404(.A1(new_n1588_), .A2(new_n196_), .B(new_n1573_), .ZN(new_n1597_));
  AOI21_X1   g01405(.A1(new_n1595_), .A2(new_n1597_), .B(new_n1558_), .ZN(new_n1598_));
  NOR2_X1    g01406(.A1(new_n1596_), .A2(new_n1598_), .ZN(new_n1599_));
  INV_X1     g01407(.I(new_n1572_), .ZN(new_n1600_));
  OAI21_X1   g01408(.A1(new_n1583_), .A2(new_n1552_), .B(\asqrt[61] ), .ZN(new_n1601_));
  INV_X1     g01409(.I(new_n1574_), .ZN(new_n1602_));
  NAND3_X1   g01410(.A1(new_n1587_), .A2(new_n1583_), .A3(new_n1602_), .ZN(new_n1603_));
  OAI21_X1   g01411(.A1(new_n1603_), .A2(new_n1601_), .B(new_n1600_), .ZN(new_n1604_));
  INV_X1     g01412(.I(new_n1578_), .ZN(new_n1605_));
  OAI21_X1   g01413(.A1(new_n1604_), .A2(new_n1605_), .B(new_n1580_), .ZN(new_n1606_));
  OAI21_X1   g01414(.A1(new_n1588_), .A2(new_n196_), .B(new_n1571_), .ZN(new_n1607_));
  NAND3_X1   g01415(.A1(new_n1607_), .A2(new_n1562_), .A3(new_n1592_), .ZN(new_n1608_));
  NOR3_X1    g01416(.A1(new_n1608_), .A2(new_n1564_), .A3(new_n1606_), .ZN(\asqrt[50] ));
  NOR3_X1    g01417(.A1(new_n1585_), .A2(\asqrt[61] ), .A3(new_n1554_), .ZN(new_n1610_));
  NAND2_X1   g01418(.A1(\asqrt[50] ), .A2(new_n1610_), .ZN(new_n1611_));
  XOR2_X1    g01419(.A1(new_n1611_), .A2(new_n1523_), .Z(new_n1612_));
  NOR2_X1    g01420(.A1(new_n1612_), .A2(new_n196_), .ZN(new_n1613_));
  INV_X1     g01421(.I(new_n1613_), .ZN(new_n1614_));
  INV_X1     g01422(.I(\a[100] ), .ZN(new_n1615_));
  NOR2_X1    g01423(.A1(\a[98] ), .A2(\a[99] ), .ZN(new_n1616_));
  INV_X1     g01424(.I(new_n1616_), .ZN(new_n1617_));
  NOR3_X1    g01425(.A1(new_n1447_), .A2(new_n1615_), .A3(new_n1617_), .ZN(new_n1618_));
  NAND2_X1   g01426(.A1(new_n1460_), .A2(new_n1618_), .ZN(new_n1619_));
  XOR2_X1    g01427(.A1(new_n1619_), .A2(\a[101] ), .Z(new_n1620_));
  INV_X1     g01428(.I(\a[101] ), .ZN(new_n1621_));
  NOR4_X1    g01429(.A1(new_n1608_), .A2(new_n1621_), .A3(new_n1564_), .A4(new_n1606_), .ZN(new_n1622_));
  NOR2_X1    g01430(.A1(new_n1621_), .A2(\a[100] ), .ZN(new_n1623_));
  OAI21_X1   g01431(.A1(new_n1622_), .A2(new_n1623_), .B(new_n1620_), .ZN(new_n1624_));
  INV_X1     g01432(.I(new_n1620_), .ZN(new_n1625_));
  NAND4_X1   g01433(.A1(new_n1594_), .A2(new_n1579_), .A3(\a[101] ), .A4(new_n1565_), .ZN(new_n1626_));
  NAND3_X1   g01434(.A1(new_n1626_), .A2(\a[100] ), .A3(new_n1625_), .ZN(new_n1627_));
  NAND2_X1   g01435(.A1(new_n1624_), .A2(new_n1627_), .ZN(new_n1628_));
  NOR2_X1    g01436(.A1(new_n1608_), .A2(new_n1606_), .ZN(new_n1629_));
  NOR4_X1    g01437(.A1(new_n1411_), .A2(new_n1374_), .A3(new_n1445_), .A4(new_n1412_), .ZN(new_n1630_));
  NAND2_X1   g01438(.A1(\asqrt[51] ), .A2(\a[100] ), .ZN(new_n1631_));
  XOR2_X1    g01439(.A1(new_n1631_), .A2(new_n1630_), .Z(new_n1632_));
  NOR2_X1    g01440(.A1(new_n1632_), .A2(new_n1617_), .ZN(new_n1633_));
  INV_X1     g01441(.I(new_n1633_), .ZN(new_n1634_));
  NAND2_X1   g01442(.A1(new_n1593_), .A2(new_n1564_), .ZN(new_n1635_));
  NOR2_X1    g01443(.A1(new_n1635_), .A2(new_n1436_), .ZN(new_n1636_));
  NAND3_X1   g01444(.A1(new_n1606_), .A2(new_n1589_), .A3(new_n1636_), .ZN(new_n1637_));
  NAND2_X1   g01445(.A1(new_n1637_), .A2(new_n1240_), .ZN(new_n1638_));
  NAND3_X1   g01446(.A1(new_n1638_), .A2(new_n1244_), .A3(new_n1595_), .ZN(new_n1639_));
  NAND4_X1   g01447(.A1(new_n1523_), .A2(new_n1583_), .A3(new_n1587_), .A4(new_n1602_), .ZN(new_n1640_));
  NAND3_X1   g01448(.A1(new_n1640_), .A2(new_n1600_), .A3(new_n1578_), .ZN(new_n1641_));
  AOI22_X1   g01449(.A1(new_n1641_), .A2(new_n1580_), .B1(new_n1607_), .B2(new_n1562_), .ZN(new_n1642_));
  AOI21_X1   g01450(.A1(new_n1642_), .A2(new_n1636_), .B(\a[102] ), .ZN(new_n1643_));
  OAI21_X1   g01451(.A1(new_n1643_), .A2(new_n1428_), .B(\asqrt[50] ), .ZN(new_n1644_));
  NAND4_X1   g01452(.A1(new_n1644_), .A2(new_n1639_), .A3(new_n1260_), .A4(new_n1634_), .ZN(new_n1645_));
  NAND2_X1   g01453(.A1(new_n1645_), .A2(new_n1628_), .ZN(new_n1646_));
  NAND3_X1   g01454(.A1(new_n1624_), .A2(new_n1627_), .A3(new_n1634_), .ZN(new_n1647_));
  AOI21_X1   g01455(.A1(\asqrt[51] ), .A2(new_n1240_), .B(\a[103] ), .ZN(new_n1648_));
  NOR2_X1    g01456(.A1(new_n1425_), .A2(\a[102] ), .ZN(new_n1649_));
  NOR2_X1    g01457(.A1(new_n1649_), .A2(new_n1648_), .ZN(new_n1650_));
  OAI21_X1   g01458(.A1(new_n1435_), .A2(new_n1246_), .B(new_n1240_), .ZN(new_n1651_));
  NAND2_X1   g01459(.A1(\asqrt[51] ), .A2(new_n1651_), .ZN(new_n1652_));
  OAI21_X1   g01460(.A1(new_n1595_), .A2(new_n1652_), .B(new_n1650_), .ZN(new_n1653_));
  INV_X1     g01461(.I(new_n1650_), .ZN(new_n1654_));
  INV_X1     g01462(.I(new_n1652_), .ZN(new_n1655_));
  NAND3_X1   g01463(.A1(\asqrt[50] ), .A2(new_n1654_), .A3(new_n1655_), .ZN(new_n1656_));
  NAND3_X1   g01464(.A1(new_n1653_), .A2(new_n1656_), .A3(new_n1096_), .ZN(new_n1657_));
  AOI21_X1   g01465(.A1(new_n1647_), .A2(\asqrt[52] ), .B(new_n1657_), .ZN(new_n1658_));
  NOR2_X1    g01466(.A1(new_n1646_), .A2(new_n1658_), .ZN(new_n1659_));
  AOI22_X1   g01467(.A1(new_n1645_), .A2(new_n1628_), .B1(\asqrt[52] ), .B2(new_n1647_), .ZN(new_n1660_));
  AOI21_X1   g01468(.A1(new_n1450_), .A2(new_n1463_), .B(\asqrt[53] ), .ZN(new_n1661_));
  NAND2_X1   g01469(.A1(new_n1661_), .A2(new_n1468_), .ZN(new_n1662_));
  NOR3_X1    g01470(.A1(new_n1595_), .A2(new_n1487_), .A3(new_n1662_), .ZN(new_n1663_));
  NOR2_X1    g01471(.A1(new_n1468_), .A2(new_n1096_), .ZN(new_n1664_));
  NOR2_X1    g01472(.A1(new_n1663_), .A2(new_n1664_), .ZN(new_n1665_));
  NAND2_X1   g01473(.A1(new_n1665_), .A2(new_n970_), .ZN(new_n1666_));
  INV_X1     g01474(.I(new_n1666_), .ZN(new_n1667_));
  OAI21_X1   g01475(.A1(new_n1660_), .A2(new_n1096_), .B(new_n1667_), .ZN(new_n1668_));
  NAND2_X1   g01476(.A1(new_n1668_), .A2(new_n1659_), .ZN(new_n1669_));
  OAI22_X1   g01477(.A1(new_n1660_), .A2(new_n1096_), .B1(new_n1646_), .B2(new_n1658_), .ZN(new_n1670_));
  NAND2_X1   g01478(.A1(new_n1526_), .A2(new_n1527_), .ZN(new_n1671_));
  NAND4_X1   g01479(.A1(\asqrt[50] ), .A2(new_n970_), .A3(new_n1671_), .A4(new_n1531_), .ZN(new_n1672_));
  XOR2_X1    g01480(.A1(new_n1672_), .A2(new_n1546_), .Z(new_n1673_));
  NAND2_X1   g01481(.A1(new_n1673_), .A2(new_n825_), .ZN(new_n1674_));
  AOI21_X1   g01482(.A1(new_n1670_), .A2(\asqrt[54] ), .B(new_n1674_), .ZN(new_n1675_));
  NOR2_X1    g01483(.A1(new_n1675_), .A2(new_n1669_), .ZN(new_n1676_));
  AOI22_X1   g01484(.A1(new_n1670_), .A2(\asqrt[54] ), .B1(new_n1668_), .B2(new_n1659_), .ZN(new_n1677_));
  NOR2_X1    g01485(.A1(new_n1490_), .A2(new_n1491_), .ZN(new_n1678_));
  NOR4_X1    g01486(.A1(new_n1595_), .A2(\asqrt[55] ), .A3(new_n1678_), .A4(new_n1534_), .ZN(new_n1679_));
  XOR2_X1    g01487(.A1(new_n1679_), .A2(new_n1547_), .Z(new_n1680_));
  NAND2_X1   g01488(.A1(new_n1680_), .A2(new_n724_), .ZN(new_n1681_));
  INV_X1     g01489(.I(new_n1681_), .ZN(new_n1682_));
  OAI21_X1   g01490(.A1(new_n1677_), .A2(new_n825_), .B(new_n1682_), .ZN(new_n1683_));
  NAND2_X1   g01491(.A1(new_n1683_), .A2(new_n1676_), .ZN(new_n1684_));
  OAI22_X1   g01492(.A1(new_n1677_), .A2(new_n825_), .B1(new_n1675_), .B2(new_n1669_), .ZN(new_n1685_));
  INV_X1     g01493(.I(new_n1537_), .ZN(new_n1686_));
  NOR4_X1    g01494(.A1(new_n1595_), .A2(\asqrt[56] ), .A3(new_n1497_), .A4(new_n1686_), .ZN(new_n1687_));
  XOR2_X1    g01495(.A1(new_n1687_), .A2(new_n1500_), .Z(new_n1688_));
  NAND2_X1   g01496(.A1(new_n1688_), .A2(new_n587_), .ZN(new_n1689_));
  AOI21_X1   g01497(.A1(new_n1685_), .A2(\asqrt[56] ), .B(new_n1689_), .ZN(new_n1690_));
  NOR2_X1    g01498(.A1(new_n1690_), .A2(new_n1684_), .ZN(new_n1691_));
  AOI22_X1   g01499(.A1(new_n1685_), .A2(\asqrt[56] ), .B1(new_n1683_), .B2(new_n1676_), .ZN(new_n1692_));
  NOR4_X1    g01500(.A1(new_n1595_), .A2(\asqrt[57] ), .A3(new_n1503_), .A4(new_n1540_), .ZN(new_n1693_));
  XOR2_X1    g01501(.A1(new_n1693_), .A2(new_n1549_), .Z(new_n1694_));
  NAND2_X1   g01502(.A1(new_n1694_), .A2(new_n504_), .ZN(new_n1695_));
  INV_X1     g01503(.I(new_n1695_), .ZN(new_n1696_));
  OAI21_X1   g01504(.A1(new_n1692_), .A2(new_n587_), .B(new_n1696_), .ZN(new_n1697_));
  NAND2_X1   g01505(.A1(new_n1697_), .A2(new_n1691_), .ZN(new_n1698_));
  OAI22_X1   g01506(.A1(new_n1692_), .A2(new_n587_), .B1(new_n1690_), .B2(new_n1684_), .ZN(new_n1699_));
  INV_X1     g01507(.I(new_n1543_), .ZN(new_n1700_));
  NOR4_X1    g01508(.A1(new_n1595_), .A2(\asqrt[58] ), .A3(new_n1508_), .A4(new_n1700_), .ZN(new_n1701_));
  XOR2_X1    g01509(.A1(new_n1701_), .A2(new_n1511_), .Z(new_n1702_));
  NAND2_X1   g01510(.A1(new_n1702_), .A2(new_n376_), .ZN(new_n1703_));
  AOI21_X1   g01511(.A1(new_n1699_), .A2(\asqrt[58] ), .B(new_n1703_), .ZN(new_n1704_));
  NOR2_X1    g01512(.A1(new_n1704_), .A2(new_n1698_), .ZN(new_n1705_));
  AOI22_X1   g01513(.A1(new_n1699_), .A2(\asqrt[58] ), .B1(new_n1697_), .B2(new_n1691_), .ZN(new_n1706_));
  NOR4_X1    g01514(.A1(new_n1595_), .A2(\asqrt[59] ), .A3(new_n1513_), .A4(new_n1581_), .ZN(new_n1707_));
  XOR2_X1    g01515(.A1(new_n1707_), .A2(new_n1551_), .Z(new_n1708_));
  NAND2_X1   g01516(.A1(new_n1708_), .A2(new_n275_), .ZN(new_n1709_));
  INV_X1     g01517(.I(new_n1709_), .ZN(new_n1710_));
  OAI21_X1   g01518(.A1(new_n1706_), .A2(new_n376_), .B(new_n1710_), .ZN(new_n1711_));
  NAND2_X1   g01519(.A1(new_n1711_), .A2(new_n1705_), .ZN(new_n1712_));
  OAI22_X1   g01520(.A1(new_n1706_), .A2(new_n376_), .B1(new_n1704_), .B2(new_n1698_), .ZN(new_n1713_));
  INV_X1     g01521(.I(new_n1584_), .ZN(new_n1714_));
  NOR4_X1    g01522(.A1(new_n1595_), .A2(\asqrt[60] ), .A3(new_n1519_), .A4(new_n1714_), .ZN(new_n1715_));
  XOR2_X1    g01523(.A1(new_n1715_), .A2(new_n1522_), .Z(new_n1716_));
  NAND2_X1   g01524(.A1(new_n1716_), .A2(new_n229_), .ZN(new_n1717_));
  AOI21_X1   g01525(.A1(new_n1713_), .A2(\asqrt[60] ), .B(new_n1717_), .ZN(new_n1718_));
  NOR2_X1    g01526(.A1(new_n1718_), .A2(new_n1712_), .ZN(new_n1719_));
  NOR2_X1    g01527(.A1(new_n1692_), .A2(new_n587_), .ZN(new_n1720_));
  OAI21_X1   g01528(.A1(new_n1720_), .A2(new_n1691_), .B(\asqrt[58] ), .ZN(new_n1721_));
  AOI21_X1   g01529(.A1(new_n1721_), .A2(new_n1698_), .B(new_n376_), .ZN(new_n1722_));
  OAI21_X1   g01530(.A1(new_n1705_), .A2(new_n1722_), .B(\asqrt[60] ), .ZN(new_n1723_));
  AOI21_X1   g01531(.A1(new_n1712_), .A2(new_n1723_), .B(new_n229_), .ZN(new_n1724_));
  INV_X1     g01532(.I(new_n1612_), .ZN(new_n1725_));
  NOR2_X1    g01533(.A1(new_n1725_), .A2(\asqrt[62] ), .ZN(new_n1726_));
  INV_X1     g01534(.I(new_n1726_), .ZN(new_n1727_));
  NAND3_X1   g01535(.A1(new_n1719_), .A2(new_n1724_), .A3(new_n1727_), .ZN(new_n1728_));
  AND3_X2    g01536(.A1(new_n1595_), .A2(new_n1571_), .A3(new_n1589_), .Z(new_n1729_));
  OAI21_X1   g01537(.A1(new_n1729_), .A2(new_n1576_), .B(new_n231_), .ZN(new_n1730_));
  INV_X1     g01538(.I(new_n1730_), .ZN(new_n1731_));
  NAND3_X1   g01539(.A1(new_n1728_), .A2(new_n1614_), .A3(new_n1731_), .ZN(new_n1732_));
  INV_X1     g01540(.I(new_n1599_), .ZN(new_n1733_));
  AOI22_X1   g01541(.A1(new_n1713_), .A2(\asqrt[60] ), .B1(new_n1711_), .B2(new_n1705_), .ZN(new_n1734_));
  OAI22_X1   g01542(.A1(new_n1734_), .A2(new_n229_), .B1(new_n1718_), .B2(new_n1712_), .ZN(new_n1735_));
  NOR4_X1    g01543(.A1(new_n1735_), .A2(\asqrt[62] ), .A3(new_n1733_), .A4(new_n1612_), .ZN(new_n1736_));
  AOI21_X1   g01544(.A1(new_n1732_), .A2(new_n1599_), .B(new_n1736_), .ZN(new_n1737_));
  INV_X1     g01545(.I(\a[96] ), .ZN(new_n1738_));
  OAI21_X1   g01546(.A1(new_n1580_), .A2(new_n1604_), .B(\asqrt[50] ), .ZN(new_n1739_));
  XOR2_X1    g01547(.A1(new_n1604_), .A2(\asqrt[63] ), .Z(new_n1740_));
  NAND2_X1   g01548(.A1(new_n1739_), .A2(new_n1740_), .ZN(new_n1741_));
  INV_X1     g01549(.I(new_n1741_), .ZN(new_n1742_));
  NAND3_X1   g01550(.A1(new_n1629_), .A2(new_n1564_), .A3(new_n1580_), .ZN(new_n1743_));
  INV_X1     g01551(.I(new_n1743_), .ZN(new_n1744_));
  NOR2_X1    g01552(.A1(new_n1742_), .A2(new_n1744_), .ZN(new_n1745_));
  NOR2_X1    g01553(.A1(\a[94] ), .A2(\a[95] ), .ZN(new_n1746_));
  INV_X1     g01554(.I(new_n1746_), .ZN(new_n1747_));
  NOR3_X1    g01555(.A1(new_n1745_), .A2(new_n1738_), .A3(new_n1747_), .ZN(new_n1748_));
  NAND2_X1   g01556(.A1(new_n1737_), .A2(new_n1748_), .ZN(new_n1749_));
  XOR2_X1    g01557(.A1(new_n1749_), .A2(\a[97] ), .Z(new_n1750_));
  INV_X1     g01558(.I(new_n1750_), .ZN(new_n1751_));
  INV_X1     g01559(.I(new_n1623_), .ZN(new_n1752_));
  AOI21_X1   g01560(.A1(new_n1626_), .A2(new_n1752_), .B(new_n1625_), .ZN(new_n1753_));
  NOR3_X1    g01561(.A1(new_n1622_), .A2(new_n1615_), .A3(new_n1620_), .ZN(new_n1754_));
  NOR3_X1    g01562(.A1(new_n1754_), .A2(new_n1753_), .A3(new_n1633_), .ZN(new_n1755_));
  AOI21_X1   g01563(.A1(\asqrt[50] ), .A2(new_n1655_), .B(new_n1654_), .ZN(new_n1756_));
  NOR3_X1    g01564(.A1(new_n1595_), .A2(new_n1650_), .A3(new_n1652_), .ZN(new_n1757_));
  NOR3_X1    g01565(.A1(new_n1756_), .A2(new_n1757_), .A3(\asqrt[53] ), .ZN(new_n1758_));
  OAI21_X1   g01566(.A1(new_n1755_), .A2(new_n1260_), .B(new_n1758_), .ZN(new_n1759_));
  NAND3_X1   g01567(.A1(new_n1759_), .A2(new_n1628_), .A3(new_n1645_), .ZN(new_n1760_));
  NOR2_X1    g01568(.A1(new_n1754_), .A2(new_n1753_), .ZN(new_n1761_));
  NOR3_X1    g01569(.A1(new_n1643_), .A2(new_n1428_), .A3(\asqrt[50] ), .ZN(new_n1762_));
  AOI21_X1   g01570(.A1(new_n1638_), .A2(new_n1244_), .B(new_n1595_), .ZN(new_n1763_));
  NOR3_X1    g01571(.A1(new_n1762_), .A2(new_n1763_), .A3(\asqrt[52] ), .ZN(new_n1764_));
  AOI21_X1   g01572(.A1(new_n1764_), .A2(new_n1634_), .B(new_n1761_), .ZN(new_n1765_));
  NOR2_X1    g01573(.A1(new_n1755_), .A2(new_n1260_), .ZN(new_n1766_));
  OAI21_X1   g01574(.A1(new_n1765_), .A2(new_n1766_), .B(\asqrt[53] ), .ZN(new_n1767_));
  AOI21_X1   g01575(.A1(new_n1767_), .A2(new_n1667_), .B(new_n1760_), .ZN(new_n1768_));
  AOI21_X1   g01576(.A1(new_n1767_), .A2(new_n1760_), .B(new_n970_), .ZN(new_n1769_));
  OAI21_X1   g01577(.A1(new_n1769_), .A2(new_n1674_), .B(new_n1768_), .ZN(new_n1770_));
  OAI21_X1   g01578(.A1(new_n1768_), .A2(new_n1769_), .B(\asqrt[55] ), .ZN(new_n1771_));
  AOI21_X1   g01579(.A1(new_n1771_), .A2(new_n1682_), .B(new_n1770_), .ZN(new_n1772_));
  AOI21_X1   g01580(.A1(new_n1770_), .A2(new_n1771_), .B(new_n724_), .ZN(new_n1773_));
  OAI21_X1   g01581(.A1(new_n1773_), .A2(new_n1689_), .B(new_n1772_), .ZN(new_n1774_));
  OAI21_X1   g01582(.A1(new_n1772_), .A2(new_n1773_), .B(\asqrt[57] ), .ZN(new_n1775_));
  AOI21_X1   g01583(.A1(new_n1775_), .A2(new_n1696_), .B(new_n1774_), .ZN(new_n1776_));
  AOI21_X1   g01584(.A1(new_n1774_), .A2(new_n1775_), .B(new_n504_), .ZN(new_n1777_));
  OAI21_X1   g01585(.A1(new_n1777_), .A2(new_n1703_), .B(new_n1776_), .ZN(new_n1778_));
  OAI21_X1   g01586(.A1(new_n1776_), .A2(new_n1777_), .B(\asqrt[59] ), .ZN(new_n1779_));
  AOI21_X1   g01587(.A1(new_n1779_), .A2(new_n1710_), .B(new_n1778_), .ZN(new_n1780_));
  AOI21_X1   g01588(.A1(new_n1778_), .A2(new_n1779_), .B(new_n275_), .ZN(new_n1781_));
  OAI21_X1   g01589(.A1(new_n1780_), .A2(new_n1781_), .B(\asqrt[61] ), .ZN(new_n1782_));
  NOR4_X1    g01590(.A1(new_n1782_), .A2(new_n1712_), .A3(new_n1718_), .A4(new_n1726_), .ZN(new_n1783_));
  NOR3_X1    g01591(.A1(new_n1783_), .A2(new_n1613_), .A3(new_n1730_), .ZN(new_n1784_));
  NOR4_X1    g01592(.A1(new_n1762_), .A2(new_n1763_), .A3(\asqrt[52] ), .A4(new_n1633_), .ZN(new_n1785_));
  OAI22_X1   g01593(.A1(new_n1785_), .A2(new_n1761_), .B1(new_n1260_), .B2(new_n1755_), .ZN(new_n1786_));
  AOI22_X1   g01594(.A1(new_n1786_), .A2(\asqrt[53] ), .B1(new_n1765_), .B2(new_n1759_), .ZN(new_n1787_));
  INV_X1     g01595(.I(new_n1674_), .ZN(new_n1788_));
  OAI21_X1   g01596(.A1(new_n1787_), .A2(new_n970_), .B(new_n1788_), .ZN(new_n1789_));
  AOI21_X1   g01597(.A1(new_n1786_), .A2(\asqrt[53] ), .B(new_n1666_), .ZN(new_n1790_));
  OAI22_X1   g01598(.A1(new_n1787_), .A2(new_n970_), .B1(new_n1790_), .B2(new_n1760_), .ZN(new_n1791_));
  AOI22_X1   g01599(.A1(new_n1791_), .A2(\asqrt[55] ), .B1(new_n1789_), .B2(new_n1768_), .ZN(new_n1792_));
  INV_X1     g01600(.I(new_n1689_), .ZN(new_n1793_));
  OAI21_X1   g01601(.A1(new_n1792_), .A2(new_n724_), .B(new_n1793_), .ZN(new_n1794_));
  AOI21_X1   g01602(.A1(new_n1791_), .A2(\asqrt[55] ), .B(new_n1681_), .ZN(new_n1795_));
  OAI22_X1   g01603(.A1(new_n1792_), .A2(new_n724_), .B1(new_n1795_), .B2(new_n1770_), .ZN(new_n1796_));
  AOI22_X1   g01604(.A1(new_n1796_), .A2(\asqrt[57] ), .B1(new_n1794_), .B2(new_n1772_), .ZN(new_n1797_));
  INV_X1     g01605(.I(new_n1703_), .ZN(new_n1798_));
  OAI21_X1   g01606(.A1(new_n1797_), .A2(new_n504_), .B(new_n1798_), .ZN(new_n1799_));
  AOI21_X1   g01607(.A1(new_n1796_), .A2(\asqrt[57] ), .B(new_n1695_), .ZN(new_n1800_));
  OAI22_X1   g01608(.A1(new_n1797_), .A2(new_n504_), .B1(new_n1800_), .B2(new_n1774_), .ZN(new_n1801_));
  AOI22_X1   g01609(.A1(new_n1801_), .A2(\asqrt[59] ), .B1(new_n1799_), .B2(new_n1776_), .ZN(new_n1802_));
  INV_X1     g01610(.I(new_n1717_), .ZN(new_n1803_));
  OAI21_X1   g01611(.A1(new_n1802_), .A2(new_n275_), .B(new_n1803_), .ZN(new_n1804_));
  AOI21_X1   g01612(.A1(new_n1801_), .A2(\asqrt[59] ), .B(new_n1709_), .ZN(new_n1805_));
  OAI22_X1   g01613(.A1(new_n1802_), .A2(new_n275_), .B1(new_n1805_), .B2(new_n1778_), .ZN(new_n1806_));
  AOI22_X1   g01614(.A1(new_n1806_), .A2(\asqrt[61] ), .B1(new_n1804_), .B2(new_n1780_), .ZN(new_n1807_));
  NAND4_X1   g01615(.A1(new_n1807_), .A2(new_n196_), .A3(new_n1599_), .A4(new_n1725_), .ZN(new_n1808_));
  NOR4_X1    g01616(.A1(new_n1784_), .A2(new_n1733_), .A3(new_n1808_), .A4(new_n1741_), .ZN(new_n1809_));
  NAND3_X1   g01617(.A1(new_n1809_), .A2(new_n1599_), .A3(new_n1743_), .ZN(new_n1810_));
  INV_X1     g01618(.I(new_n1810_), .ZN(new_n1811_));
  NOR2_X1    g01619(.A1(new_n1807_), .A2(new_n196_), .ZN(new_n1812_));
  INV_X1     g01620(.I(new_n1812_), .ZN(new_n1813_));
  NOR2_X1    g01621(.A1(new_n1735_), .A2(\asqrt[62] ), .ZN(new_n1814_));
  NAND2_X1   g01622(.A1(new_n1804_), .A2(new_n1780_), .ZN(new_n1815_));
  NAND3_X1   g01623(.A1(new_n1806_), .A2(\asqrt[61] ), .A3(new_n1727_), .ZN(new_n1816_));
  OAI21_X1   g01624(.A1(new_n1816_), .A2(new_n1815_), .B(new_n1614_), .ZN(new_n1817_));
  OAI21_X1   g01625(.A1(new_n1817_), .A2(new_n1730_), .B(new_n1599_), .ZN(new_n1818_));
  NAND2_X1   g01626(.A1(new_n1736_), .A2(new_n1742_), .ZN(new_n1819_));
  NOR3_X1    g01627(.A1(new_n1819_), .A2(new_n1818_), .A3(new_n1743_), .ZN(\asqrt[49] ));
  NAND4_X1   g01628(.A1(\asqrt[49] ), .A2(new_n1725_), .A3(new_n1812_), .A4(new_n1814_), .ZN(new_n1821_));
  NOR3_X1    g01629(.A1(\asqrt[49] ), .A2(new_n1725_), .A3(new_n1814_), .ZN(new_n1822_));
  OAI21_X1   g01630(.A1(new_n1813_), .A2(new_n1822_), .B(new_n1821_), .ZN(new_n1823_));
  NOR3_X1    g01631(.A1(new_n1806_), .A2(\asqrt[61] ), .A3(new_n1716_), .ZN(new_n1824_));
  NAND2_X1   g01632(.A1(\asqrt[49] ), .A2(new_n1824_), .ZN(new_n1825_));
  XOR2_X1    g01633(.A1(new_n1825_), .A2(new_n1724_), .Z(new_n1826_));
  NOR2_X1    g01634(.A1(new_n1826_), .A2(new_n196_), .ZN(new_n1827_));
  NOR2_X1    g01635(.A1(\a[96] ), .A2(\a[97] ), .ZN(new_n1828_));
  NAND4_X1   g01636(.A1(new_n1642_), .A2(\a[98] ), .A3(new_n1635_), .A4(new_n1828_), .ZN(new_n1829_));
  XOR2_X1    g01637(.A1(new_n1829_), .A2(\a[99] ), .Z(new_n1830_));
  INV_X1     g01638(.I(new_n1830_), .ZN(new_n1831_));
  NOR3_X1    g01639(.A1(new_n1734_), .A2(new_n229_), .A3(new_n1726_), .ZN(new_n1832_));
  AOI21_X1   g01640(.A1(new_n1832_), .A2(new_n1719_), .B(new_n1613_), .ZN(new_n1833_));
  AOI21_X1   g01641(.A1(new_n1833_), .A2(new_n1731_), .B(new_n1733_), .ZN(new_n1834_));
  NOR2_X1    g01642(.A1(new_n1808_), .A2(new_n1741_), .ZN(new_n1835_));
  NAND4_X1   g01643(.A1(new_n1835_), .A2(\a[99] ), .A3(new_n1834_), .A4(new_n1744_), .ZN(new_n1836_));
  NOR2_X1    g01644(.A1(new_n1830_), .A2(\a[98] ), .ZN(new_n1837_));
  INV_X1     g01645(.I(new_n1837_), .ZN(new_n1838_));
  AOI21_X1   g01646(.A1(new_n1836_), .A2(new_n1838_), .B(new_n1831_), .ZN(new_n1839_));
  INV_X1     g01647(.I(\a[98] ), .ZN(new_n1840_));
  INV_X1     g01648(.I(\a[99] ), .ZN(new_n1841_));
  NOR4_X1    g01649(.A1(new_n1819_), .A2(new_n1818_), .A3(new_n1841_), .A4(new_n1743_), .ZN(new_n1842_));
  NOR3_X1    g01650(.A1(new_n1842_), .A2(new_n1840_), .A3(new_n1830_), .ZN(new_n1843_));
  NOR2_X1    g01651(.A1(new_n1843_), .A2(new_n1839_), .ZN(new_n1844_));
  INV_X1     g01652(.I(new_n1828_), .ZN(new_n1845_));
  NAND4_X1   g01653(.A1(new_n1594_), .A2(new_n1565_), .A3(new_n1580_), .A4(new_n1641_), .ZN(new_n1846_));
  NOR2_X1    g01654(.A1(new_n1595_), .A2(new_n1840_), .ZN(new_n1847_));
  XOR2_X1    g01655(.A1(new_n1847_), .A2(new_n1846_), .Z(new_n1848_));
  NOR2_X1    g01656(.A1(new_n1848_), .A2(new_n1845_), .ZN(new_n1849_));
  NAND2_X1   g01657(.A1(new_n1745_), .A2(\asqrt[50] ), .ZN(new_n1850_));
  INV_X1     g01658(.I(new_n1850_), .ZN(new_n1851_));
  AOI21_X1   g01659(.A1(new_n1737_), .A2(new_n1851_), .B(\a[100] ), .ZN(new_n1852_));
  NOR3_X1    g01660(.A1(new_n1852_), .A2(new_n1617_), .A3(\asqrt[49] ), .ZN(new_n1853_));
  NAND3_X1   g01661(.A1(new_n1835_), .A2(new_n1834_), .A3(new_n1744_), .ZN(new_n1854_));
  OAI21_X1   g01662(.A1(new_n1784_), .A2(new_n1733_), .B(new_n1808_), .ZN(new_n1855_));
  OAI21_X1   g01663(.A1(new_n1855_), .A2(new_n1850_), .B(new_n1615_), .ZN(new_n1856_));
  AOI21_X1   g01664(.A1(new_n1856_), .A2(new_n1616_), .B(new_n1854_), .ZN(new_n1857_));
  NOR4_X1    g01665(.A1(new_n1853_), .A2(new_n1857_), .A3(\asqrt[51] ), .A4(new_n1849_), .ZN(new_n1858_));
  NOR2_X1    g01666(.A1(new_n1858_), .A2(new_n1844_), .ZN(new_n1859_));
  NOR3_X1    g01667(.A1(new_n1843_), .A2(new_n1839_), .A3(new_n1849_), .ZN(new_n1860_));
  AOI21_X1   g01668(.A1(\asqrt[50] ), .A2(new_n1615_), .B(\a[101] ), .ZN(new_n1861_));
  NOR2_X1    g01669(.A1(new_n1626_), .A2(\a[100] ), .ZN(new_n1862_));
  AOI21_X1   g01670(.A1(\asqrt[50] ), .A2(\a[100] ), .B(new_n1619_), .ZN(new_n1863_));
  OAI21_X1   g01671(.A1(new_n1862_), .A2(new_n1861_), .B(new_n1863_), .ZN(new_n1864_));
  NOR3_X1    g01672(.A1(new_n1854_), .A2(new_n1633_), .A3(new_n1864_), .ZN(new_n1865_));
  INV_X1     g01673(.I(new_n1864_), .ZN(new_n1866_));
  AOI21_X1   g01674(.A1(\asqrt[49] ), .A2(new_n1866_), .B(new_n1634_), .ZN(new_n1867_));
  NOR3_X1    g01675(.A1(new_n1867_), .A2(new_n1865_), .A3(\asqrt[52] ), .ZN(new_n1868_));
  OAI21_X1   g01676(.A1(new_n1860_), .A2(new_n1436_), .B(new_n1868_), .ZN(new_n1869_));
  NAND2_X1   g01677(.A1(new_n1859_), .A2(new_n1869_), .ZN(new_n1870_));
  OAI22_X1   g01678(.A1(new_n1858_), .A2(new_n1844_), .B1(new_n1436_), .B2(new_n1860_), .ZN(new_n1871_));
  AOI21_X1   g01679(.A1(new_n1644_), .A2(new_n1639_), .B(\asqrt[52] ), .ZN(new_n1872_));
  NAND2_X1   g01680(.A1(new_n1872_), .A2(new_n1755_), .ZN(new_n1873_));
  NOR3_X1    g01681(.A1(new_n1854_), .A2(new_n1766_), .A3(new_n1873_), .ZN(new_n1874_));
  NOR2_X1    g01682(.A1(new_n1755_), .A2(new_n1260_), .ZN(new_n1875_));
  NOR2_X1    g01683(.A1(new_n1874_), .A2(new_n1875_), .ZN(new_n1876_));
  NAND2_X1   g01684(.A1(new_n1876_), .A2(new_n1096_), .ZN(new_n1877_));
  AOI21_X1   g01685(.A1(new_n1871_), .A2(\asqrt[52] ), .B(new_n1877_), .ZN(new_n1878_));
  NOR2_X1    g01686(.A1(new_n1878_), .A2(new_n1870_), .ZN(new_n1879_));
  AOI22_X1   g01687(.A1(new_n1871_), .A2(\asqrt[52] ), .B1(new_n1859_), .B2(new_n1869_), .ZN(new_n1880_));
  NAND2_X1   g01688(.A1(new_n1653_), .A2(new_n1656_), .ZN(new_n1881_));
  NAND4_X1   g01689(.A1(\asqrt[49] ), .A2(new_n1096_), .A3(new_n1881_), .A4(new_n1660_), .ZN(new_n1882_));
  XNOR2_X1   g01690(.A1(new_n1882_), .A2(new_n1767_), .ZN(new_n1883_));
  NAND2_X1   g01691(.A1(new_n1883_), .A2(new_n970_), .ZN(new_n1884_));
  INV_X1     g01692(.I(new_n1884_), .ZN(new_n1885_));
  OAI21_X1   g01693(.A1(new_n1880_), .A2(new_n1096_), .B(new_n1885_), .ZN(new_n1886_));
  NAND2_X1   g01694(.A1(new_n1886_), .A2(new_n1879_), .ZN(new_n1887_));
  OAI21_X1   g01695(.A1(new_n1842_), .A2(new_n1837_), .B(new_n1830_), .ZN(new_n1888_));
  NAND3_X1   g01696(.A1(new_n1836_), .A2(\a[98] ), .A3(new_n1831_), .ZN(new_n1889_));
  INV_X1     g01697(.I(new_n1849_), .ZN(new_n1890_));
  NAND3_X1   g01698(.A1(new_n1888_), .A2(new_n1889_), .A3(new_n1890_), .ZN(new_n1891_));
  NAND4_X1   g01699(.A1(new_n1809_), .A2(new_n1634_), .A3(new_n1744_), .A4(new_n1866_), .ZN(new_n1892_));
  OAI21_X1   g01700(.A1(new_n1854_), .A2(new_n1864_), .B(new_n1633_), .ZN(new_n1893_));
  NAND3_X1   g01701(.A1(new_n1893_), .A2(new_n1260_), .A3(new_n1892_), .ZN(new_n1894_));
  AOI21_X1   g01702(.A1(new_n1891_), .A2(\asqrt[51] ), .B(new_n1894_), .ZN(new_n1895_));
  NOR3_X1    g01703(.A1(new_n1895_), .A2(new_n1844_), .A3(new_n1858_), .ZN(new_n1896_));
  NAND2_X1   g01704(.A1(new_n1888_), .A2(new_n1889_), .ZN(new_n1897_));
  NAND3_X1   g01705(.A1(new_n1856_), .A2(new_n1616_), .A3(new_n1854_), .ZN(new_n1898_));
  OAI21_X1   g01706(.A1(new_n1852_), .A2(new_n1617_), .B(\asqrt[49] ), .ZN(new_n1899_));
  NAND4_X1   g01707(.A1(new_n1899_), .A2(new_n1898_), .A3(new_n1436_), .A4(new_n1890_), .ZN(new_n1900_));
  NAND2_X1   g01708(.A1(new_n1900_), .A2(new_n1897_), .ZN(new_n1901_));
  NAND2_X1   g01709(.A1(new_n1891_), .A2(\asqrt[51] ), .ZN(new_n1902_));
  AOI21_X1   g01710(.A1(new_n1901_), .A2(new_n1902_), .B(new_n1260_), .ZN(new_n1903_));
  OAI21_X1   g01711(.A1(new_n1903_), .A2(new_n1877_), .B(new_n1896_), .ZN(new_n1904_));
  OAI21_X1   g01712(.A1(new_n1903_), .A2(new_n1896_), .B(\asqrt[53] ), .ZN(new_n1905_));
  AOI21_X1   g01713(.A1(new_n1904_), .A2(new_n1905_), .B(new_n970_), .ZN(new_n1906_));
  INV_X1     g01714(.I(new_n1906_), .ZN(new_n1907_));
  NOR4_X1    g01715(.A1(new_n1854_), .A2(\asqrt[54] ), .A3(new_n1665_), .A4(new_n1670_), .ZN(new_n1908_));
  XNOR2_X1   g01716(.A1(new_n1908_), .A2(new_n1769_), .ZN(new_n1909_));
  NAND2_X1   g01717(.A1(new_n1909_), .A2(new_n825_), .ZN(new_n1910_));
  INV_X1     g01718(.I(new_n1910_), .ZN(new_n1911_));
  AOI21_X1   g01719(.A1(new_n1907_), .A2(new_n1911_), .B(new_n1887_), .ZN(new_n1912_));
  OAI22_X1   g01720(.A1(new_n1880_), .A2(new_n1096_), .B1(new_n1878_), .B2(new_n1870_), .ZN(new_n1913_));
  AOI22_X1   g01721(.A1(new_n1913_), .A2(\asqrt[54] ), .B1(new_n1886_), .B2(new_n1879_), .ZN(new_n1914_));
  NOR4_X1    g01722(.A1(new_n1854_), .A2(\asqrt[55] ), .A3(new_n1673_), .A4(new_n1791_), .ZN(new_n1915_));
  XOR2_X1    g01723(.A1(new_n1915_), .A2(new_n1771_), .Z(new_n1916_));
  NAND2_X1   g01724(.A1(new_n1916_), .A2(new_n724_), .ZN(new_n1917_));
  INV_X1     g01725(.I(new_n1917_), .ZN(new_n1918_));
  OAI21_X1   g01726(.A1(new_n1914_), .A2(new_n825_), .B(new_n1918_), .ZN(new_n1919_));
  NAND2_X1   g01727(.A1(new_n1919_), .A2(new_n1912_), .ZN(new_n1920_));
  AOI21_X1   g01728(.A1(new_n1905_), .A2(new_n1885_), .B(new_n1904_), .ZN(new_n1921_));
  OAI21_X1   g01729(.A1(new_n1906_), .A2(new_n1910_), .B(new_n1921_), .ZN(new_n1922_));
  OAI21_X1   g01730(.A1(new_n1921_), .A2(new_n1906_), .B(\asqrt[55] ), .ZN(new_n1923_));
  NAND2_X1   g01731(.A1(new_n1922_), .A2(new_n1923_), .ZN(new_n1924_));
  NOR4_X1    g01732(.A1(new_n1854_), .A2(\asqrt[56] ), .A3(new_n1680_), .A4(new_n1685_), .ZN(new_n1925_));
  XNOR2_X1   g01733(.A1(new_n1925_), .A2(new_n1773_), .ZN(new_n1926_));
  NAND2_X1   g01734(.A1(new_n1926_), .A2(new_n587_), .ZN(new_n1927_));
  AOI21_X1   g01735(.A1(new_n1924_), .A2(\asqrt[56] ), .B(new_n1927_), .ZN(new_n1928_));
  NOR2_X1    g01736(.A1(new_n1928_), .A2(new_n1920_), .ZN(new_n1929_));
  AOI21_X1   g01737(.A1(new_n1923_), .A2(new_n1918_), .B(new_n1922_), .ZN(new_n1930_));
  AOI21_X1   g01738(.A1(new_n1922_), .A2(new_n1923_), .B(new_n724_), .ZN(new_n1931_));
  OAI21_X1   g01739(.A1(new_n1930_), .A2(new_n1931_), .B(\asqrt[57] ), .ZN(new_n1932_));
  NOR4_X1    g01740(.A1(new_n1854_), .A2(\asqrt[57] ), .A3(new_n1688_), .A4(new_n1796_), .ZN(new_n1933_));
  XOR2_X1    g01741(.A1(new_n1933_), .A2(new_n1775_), .Z(new_n1934_));
  NAND2_X1   g01742(.A1(new_n1934_), .A2(new_n504_), .ZN(new_n1935_));
  INV_X1     g01743(.I(new_n1935_), .ZN(new_n1936_));
  NAND2_X1   g01744(.A1(new_n1932_), .A2(new_n1936_), .ZN(new_n1937_));
  NAND2_X1   g01745(.A1(new_n1937_), .A2(new_n1929_), .ZN(new_n1938_));
  AOI22_X1   g01746(.A1(new_n1924_), .A2(\asqrt[56] ), .B1(new_n1919_), .B2(new_n1912_), .ZN(new_n1939_));
  OAI22_X1   g01747(.A1(new_n1939_), .A2(new_n587_), .B1(new_n1928_), .B2(new_n1920_), .ZN(new_n1940_));
  NOR4_X1    g01748(.A1(new_n1854_), .A2(\asqrt[58] ), .A3(new_n1694_), .A4(new_n1699_), .ZN(new_n1941_));
  XOR2_X1    g01749(.A1(new_n1941_), .A2(new_n1721_), .Z(new_n1942_));
  NAND2_X1   g01750(.A1(new_n1942_), .A2(new_n376_), .ZN(new_n1943_));
  AOI21_X1   g01751(.A1(new_n1940_), .A2(\asqrt[58] ), .B(new_n1943_), .ZN(new_n1944_));
  NOR2_X1    g01752(.A1(new_n1944_), .A2(new_n1938_), .ZN(new_n1945_));
  AOI22_X1   g01753(.A1(new_n1940_), .A2(\asqrt[58] ), .B1(new_n1937_), .B2(new_n1929_), .ZN(new_n1946_));
  NOR4_X1    g01754(.A1(new_n1854_), .A2(\asqrt[59] ), .A3(new_n1702_), .A4(new_n1801_), .ZN(new_n1947_));
  XOR2_X1    g01755(.A1(new_n1947_), .A2(new_n1779_), .Z(new_n1948_));
  NAND2_X1   g01756(.A1(new_n1948_), .A2(new_n275_), .ZN(new_n1949_));
  INV_X1     g01757(.I(new_n1949_), .ZN(new_n1950_));
  OAI21_X1   g01758(.A1(new_n1946_), .A2(new_n376_), .B(new_n1950_), .ZN(new_n1951_));
  NAND2_X1   g01759(.A1(new_n1951_), .A2(new_n1945_), .ZN(new_n1952_));
  OAI22_X1   g01760(.A1(new_n1946_), .A2(new_n376_), .B1(new_n1944_), .B2(new_n1938_), .ZN(new_n1953_));
  NOR4_X1    g01761(.A1(new_n1854_), .A2(\asqrt[60] ), .A3(new_n1708_), .A4(new_n1713_), .ZN(new_n1954_));
  XOR2_X1    g01762(.A1(new_n1954_), .A2(new_n1723_), .Z(new_n1955_));
  NAND2_X1   g01763(.A1(new_n1955_), .A2(new_n229_), .ZN(new_n1956_));
  AOI21_X1   g01764(.A1(new_n1953_), .A2(\asqrt[60] ), .B(new_n1956_), .ZN(new_n1957_));
  NOR2_X1    g01765(.A1(new_n1957_), .A2(new_n1952_), .ZN(new_n1958_));
  AOI22_X1   g01766(.A1(new_n1953_), .A2(\asqrt[60] ), .B1(new_n1951_), .B2(new_n1945_), .ZN(new_n1959_));
  INV_X1     g01767(.I(new_n1826_), .ZN(new_n1960_));
  NOR2_X1    g01768(.A1(new_n1960_), .A2(\asqrt[62] ), .ZN(new_n1961_));
  NOR3_X1    g01769(.A1(new_n1959_), .A2(new_n229_), .A3(new_n1961_), .ZN(new_n1962_));
  AOI21_X1   g01770(.A1(new_n1962_), .A2(new_n1958_), .B(new_n1827_), .ZN(new_n1963_));
  NAND3_X1   g01771(.A1(new_n1854_), .A2(new_n1733_), .A3(new_n1808_), .ZN(new_n1964_));
  AOI21_X1   g01772(.A1(new_n1964_), .A2(new_n1817_), .B(\asqrt[63] ), .ZN(new_n1965_));
  AOI21_X1   g01773(.A1(new_n1963_), .A2(new_n1965_), .B(new_n1823_), .ZN(new_n1966_));
  INV_X1     g01774(.I(new_n1823_), .ZN(new_n1967_));
  AOI22_X1   g01775(.A1(new_n1900_), .A2(new_n1897_), .B1(\asqrt[51] ), .B2(new_n1891_), .ZN(new_n1968_));
  INV_X1     g01776(.I(new_n1877_), .ZN(new_n1969_));
  OAI21_X1   g01777(.A1(new_n1968_), .A2(new_n1260_), .B(new_n1969_), .ZN(new_n1970_));
  OAI22_X1   g01778(.A1(new_n1968_), .A2(new_n1260_), .B1(new_n1901_), .B2(new_n1895_), .ZN(new_n1971_));
  AOI22_X1   g01779(.A1(new_n1971_), .A2(\asqrt[53] ), .B1(new_n1970_), .B2(new_n1896_), .ZN(new_n1972_));
  OAI21_X1   g01780(.A1(new_n1972_), .A2(new_n970_), .B(new_n1911_), .ZN(new_n1973_));
  AOI21_X1   g01781(.A1(new_n1971_), .A2(\asqrt[53] ), .B(new_n1884_), .ZN(new_n1974_));
  OAI22_X1   g01782(.A1(new_n1972_), .A2(new_n970_), .B1(new_n1974_), .B2(new_n1904_), .ZN(new_n1975_));
  AOI22_X1   g01783(.A1(new_n1975_), .A2(\asqrt[55] ), .B1(new_n1973_), .B2(new_n1921_), .ZN(new_n1976_));
  INV_X1     g01784(.I(new_n1927_), .ZN(new_n1977_));
  OAI21_X1   g01785(.A1(new_n1976_), .A2(new_n724_), .B(new_n1977_), .ZN(new_n1978_));
  NAND2_X1   g01786(.A1(new_n1978_), .A2(new_n1930_), .ZN(new_n1979_));
  AOI21_X1   g01787(.A1(new_n1975_), .A2(\asqrt[55] ), .B(new_n1917_), .ZN(new_n1980_));
  OAI22_X1   g01788(.A1(new_n1976_), .A2(new_n724_), .B1(new_n1980_), .B2(new_n1922_), .ZN(new_n1981_));
  AOI21_X1   g01789(.A1(new_n1981_), .A2(\asqrt[57] ), .B(new_n1935_), .ZN(new_n1982_));
  NOR2_X1    g01790(.A1(new_n1982_), .A2(new_n1979_), .ZN(new_n1983_));
  AOI22_X1   g01791(.A1(new_n1981_), .A2(\asqrt[57] ), .B1(new_n1978_), .B2(new_n1930_), .ZN(new_n1984_));
  INV_X1     g01792(.I(new_n1943_), .ZN(new_n1985_));
  OAI21_X1   g01793(.A1(new_n1984_), .A2(new_n504_), .B(new_n1985_), .ZN(new_n1986_));
  NAND2_X1   g01794(.A1(new_n1986_), .A2(new_n1983_), .ZN(new_n1987_));
  OAI22_X1   g01795(.A1(new_n1984_), .A2(new_n504_), .B1(new_n1982_), .B2(new_n1979_), .ZN(new_n1988_));
  AOI21_X1   g01796(.A1(new_n1988_), .A2(\asqrt[59] ), .B(new_n1949_), .ZN(new_n1989_));
  NOR2_X1    g01797(.A1(new_n1989_), .A2(new_n1987_), .ZN(new_n1990_));
  AOI22_X1   g01798(.A1(new_n1988_), .A2(\asqrt[59] ), .B1(new_n1986_), .B2(new_n1983_), .ZN(new_n1991_));
  INV_X1     g01799(.I(new_n1956_), .ZN(new_n1992_));
  OAI21_X1   g01800(.A1(new_n1991_), .A2(new_n275_), .B(new_n1992_), .ZN(new_n1993_));
  OAI22_X1   g01801(.A1(new_n1991_), .A2(new_n275_), .B1(new_n1989_), .B2(new_n1987_), .ZN(new_n1994_));
  AOI22_X1   g01802(.A1(new_n1994_), .A2(\asqrt[61] ), .B1(new_n1993_), .B2(new_n1990_), .ZN(new_n1995_));
  NAND4_X1   g01803(.A1(new_n1995_), .A2(new_n196_), .A3(new_n1967_), .A4(new_n1960_), .ZN(new_n1996_));
  NAND2_X1   g01804(.A1(new_n1833_), .A2(new_n1733_), .ZN(new_n1997_));
  XOR2_X1    g01805(.A1(new_n1833_), .A2(\asqrt[63] ), .Z(new_n1998_));
  AOI21_X1   g01806(.A1(\asqrt[49] ), .A2(new_n1997_), .B(new_n1998_), .ZN(new_n1999_));
  INV_X1     g01807(.I(new_n1999_), .ZN(new_n2000_));
  NOR2_X1    g01808(.A1(new_n1996_), .A2(new_n2000_), .ZN(new_n2001_));
  NAND4_X1   g01809(.A1(new_n2001_), .A2(new_n1966_), .A3(\a[97] ), .A4(new_n1811_), .ZN(new_n2002_));
  INV_X1     g01810(.I(\a[97] ), .ZN(new_n2003_));
  NOR2_X1    g01811(.A1(new_n2003_), .A2(\a[96] ), .ZN(new_n2004_));
  INV_X1     g01812(.I(new_n2004_), .ZN(new_n2005_));
  AOI21_X1   g01813(.A1(new_n2002_), .A2(new_n2005_), .B(new_n1751_), .ZN(new_n2006_));
  INV_X1     g01814(.I(new_n1827_), .ZN(new_n2007_));
  NAND2_X1   g01815(.A1(new_n1993_), .A2(new_n1990_), .ZN(new_n2008_));
  INV_X1     g01816(.I(new_n1961_), .ZN(new_n2009_));
  NAND3_X1   g01817(.A1(new_n1994_), .A2(\asqrt[61] ), .A3(new_n2009_), .ZN(new_n2010_));
  OAI21_X1   g01818(.A1(new_n2010_), .A2(new_n2008_), .B(new_n2007_), .ZN(new_n2011_));
  INV_X1     g01819(.I(new_n1965_), .ZN(new_n2012_));
  OAI21_X1   g01820(.A1(new_n2011_), .A2(new_n2012_), .B(new_n1967_), .ZN(new_n2013_));
  OAI22_X1   g01821(.A1(new_n1959_), .A2(new_n229_), .B1(new_n1957_), .B2(new_n1952_), .ZN(new_n2014_));
  NOR4_X1    g01822(.A1(new_n2014_), .A2(\asqrt[62] ), .A3(new_n1823_), .A4(new_n1826_), .ZN(new_n2015_));
  NAND2_X1   g01823(.A1(new_n2015_), .A2(new_n1999_), .ZN(new_n2016_));
  NOR4_X1    g01824(.A1(new_n2016_), .A2(new_n2003_), .A3(new_n1810_), .A4(new_n2013_), .ZN(new_n2017_));
  NOR3_X1    g01825(.A1(new_n2017_), .A2(new_n1738_), .A3(new_n1750_), .ZN(new_n2018_));
  NOR2_X1    g01826(.A1(new_n2018_), .A2(new_n2006_), .ZN(new_n2019_));
  AOI21_X1   g01827(.A1(new_n1979_), .A2(new_n1932_), .B(new_n504_), .ZN(new_n2020_));
  OAI21_X1   g01828(.A1(new_n1983_), .A2(new_n2020_), .B(\asqrt[59] ), .ZN(new_n2021_));
  AOI21_X1   g01829(.A1(new_n1987_), .A2(new_n2021_), .B(new_n275_), .ZN(new_n2022_));
  OAI21_X1   g01830(.A1(new_n1990_), .A2(new_n2022_), .B(\asqrt[61] ), .ZN(new_n2023_));
  NOR3_X1    g01831(.A1(new_n2008_), .A2(new_n2023_), .A3(new_n1961_), .ZN(new_n2024_));
  NOR3_X1    g01832(.A1(new_n2024_), .A2(new_n1827_), .A3(new_n2012_), .ZN(new_n2025_));
  NOR4_X1    g01833(.A1(new_n2025_), .A2(new_n1823_), .A3(new_n1996_), .A4(new_n2000_), .ZN(new_n2026_));
  NOR4_X1    g01834(.A1(new_n1819_), .A2(new_n1733_), .A3(new_n1784_), .A4(new_n1743_), .ZN(new_n2027_));
  NAND2_X1   g01835(.A1(\asqrt[49] ), .A2(\a[96] ), .ZN(new_n2028_));
  XOR2_X1    g01836(.A1(new_n2028_), .A2(new_n2027_), .Z(new_n2029_));
  NOR2_X1    g01837(.A1(new_n2029_), .A2(new_n1747_), .ZN(new_n2030_));
  NOR3_X1    g01838(.A1(new_n2016_), .A2(new_n1810_), .A3(new_n2013_), .ZN(\asqrt[48] ));
  INV_X1     g01839(.I(new_n1931_), .ZN(new_n2032_));
  AOI21_X1   g01840(.A1(new_n2032_), .A2(new_n1920_), .B(new_n587_), .ZN(new_n2033_));
  OAI21_X1   g01841(.A1(new_n2033_), .A2(new_n1929_), .B(\asqrt[58] ), .ZN(new_n2034_));
  AOI21_X1   g01842(.A1(new_n1938_), .A2(new_n2034_), .B(new_n376_), .ZN(new_n2035_));
  OAI21_X1   g01843(.A1(new_n1945_), .A2(new_n2035_), .B(\asqrt[60] ), .ZN(new_n2036_));
  AOI21_X1   g01844(.A1(new_n1952_), .A2(new_n2036_), .B(new_n229_), .ZN(new_n2037_));
  NAND3_X1   g01845(.A1(new_n1958_), .A2(new_n2037_), .A3(new_n2009_), .ZN(new_n2038_));
  NAND3_X1   g01846(.A1(new_n2038_), .A2(new_n2007_), .A3(new_n1965_), .ZN(new_n2039_));
  AOI21_X1   g01847(.A1(new_n2039_), .A2(new_n1967_), .B(new_n2015_), .ZN(new_n2040_));
  NOR2_X1    g01848(.A1(new_n1811_), .A2(new_n1999_), .ZN(new_n2041_));
  NAND2_X1   g01849(.A1(new_n2041_), .A2(\asqrt[49] ), .ZN(new_n2042_));
  INV_X1     g01850(.I(new_n2042_), .ZN(new_n2043_));
  AOI21_X1   g01851(.A1(new_n2040_), .A2(new_n2043_), .B(\a[98] ), .ZN(new_n2044_));
  NOR3_X1    g01852(.A1(new_n2044_), .A2(new_n1845_), .A3(\asqrt[48] ), .ZN(new_n2045_));
  NAND3_X1   g01853(.A1(new_n2001_), .A2(new_n1966_), .A3(new_n1811_), .ZN(new_n2046_));
  OAI21_X1   g01854(.A1(new_n2025_), .A2(new_n1823_), .B(new_n1996_), .ZN(new_n2047_));
  OAI21_X1   g01855(.A1(new_n2047_), .A2(new_n2042_), .B(new_n1840_), .ZN(new_n2048_));
  AOI21_X1   g01856(.A1(new_n2048_), .A2(new_n1828_), .B(new_n2046_), .ZN(new_n2049_));
  NOR4_X1    g01857(.A1(new_n2045_), .A2(new_n2049_), .A3(\asqrt[50] ), .A4(new_n2030_), .ZN(new_n2050_));
  OAI21_X1   g01858(.A1(new_n2017_), .A2(new_n2004_), .B(new_n1750_), .ZN(new_n2051_));
  NAND3_X1   g01859(.A1(new_n2002_), .A2(\a[96] ), .A3(new_n1751_), .ZN(new_n2052_));
  INV_X1     g01860(.I(new_n2030_), .ZN(new_n2053_));
  NAND3_X1   g01861(.A1(new_n2051_), .A2(new_n2052_), .A3(new_n2053_), .ZN(new_n2054_));
  AOI21_X1   g01862(.A1(\asqrt[49] ), .A2(new_n1840_), .B(\a[99] ), .ZN(new_n2055_));
  NOR2_X1    g01863(.A1(new_n1836_), .A2(\a[98] ), .ZN(new_n2056_));
  AOI21_X1   g01864(.A1(\asqrt[49] ), .A2(\a[98] ), .B(new_n1829_), .ZN(new_n2057_));
  OAI21_X1   g01865(.A1(new_n2055_), .A2(new_n2056_), .B(new_n2057_), .ZN(new_n2058_));
  INV_X1     g01866(.I(new_n2058_), .ZN(new_n2059_));
  NAND4_X1   g01867(.A1(new_n2026_), .A2(new_n1811_), .A3(new_n1890_), .A4(new_n2059_), .ZN(new_n2060_));
  OAI21_X1   g01868(.A1(new_n2046_), .A2(new_n2058_), .B(new_n1849_), .ZN(new_n2061_));
  NAND3_X1   g01869(.A1(new_n2061_), .A2(new_n1436_), .A3(new_n2060_), .ZN(new_n2062_));
  AOI21_X1   g01870(.A1(new_n2054_), .A2(\asqrt[50] ), .B(new_n2062_), .ZN(new_n2063_));
  NOR3_X1    g01871(.A1(new_n2063_), .A2(new_n2019_), .A3(new_n2050_), .ZN(new_n2064_));
  NAND2_X1   g01872(.A1(new_n2051_), .A2(new_n2052_), .ZN(new_n2065_));
  NAND3_X1   g01873(.A1(new_n2048_), .A2(new_n1828_), .A3(new_n2046_), .ZN(new_n2066_));
  OAI21_X1   g01874(.A1(new_n2044_), .A2(new_n1845_), .B(\asqrt[48] ), .ZN(new_n2067_));
  NAND4_X1   g01875(.A1(new_n2067_), .A2(new_n2066_), .A3(new_n1595_), .A4(new_n2053_), .ZN(new_n2068_));
  NAND2_X1   g01876(.A1(new_n2068_), .A2(new_n2065_), .ZN(new_n2069_));
  NAND2_X1   g01877(.A1(new_n2054_), .A2(\asqrt[50] ), .ZN(new_n2070_));
  AOI21_X1   g01878(.A1(new_n2069_), .A2(new_n2070_), .B(new_n1436_), .ZN(new_n2071_));
  AOI21_X1   g01879(.A1(new_n1899_), .A2(new_n1898_), .B(\asqrt[51] ), .ZN(new_n2072_));
  AND4_X2    g01880(.A1(new_n1860_), .A2(\asqrt[48] ), .A3(new_n1902_), .A4(new_n2072_), .Z(new_n2073_));
  NOR2_X1    g01881(.A1(new_n1860_), .A2(new_n1436_), .ZN(new_n2074_));
  NOR3_X1    g01882(.A1(new_n2073_), .A2(new_n2074_), .A3(\asqrt[52] ), .ZN(new_n2075_));
  INV_X1     g01883(.I(new_n2075_), .ZN(new_n2076_));
  OAI21_X1   g01884(.A1(new_n2071_), .A2(new_n2076_), .B(new_n2064_), .ZN(new_n2077_));
  OAI21_X1   g01885(.A1(new_n2071_), .A2(new_n2064_), .B(\asqrt[52] ), .ZN(new_n2078_));
  NAND2_X1   g01886(.A1(new_n1893_), .A2(new_n1892_), .ZN(new_n2079_));
  NAND4_X1   g01887(.A1(\asqrt[48] ), .A2(new_n1260_), .A3(new_n2079_), .A4(new_n1968_), .ZN(new_n2080_));
  XOR2_X1    g01888(.A1(new_n2080_), .A2(new_n1903_), .Z(new_n2081_));
  NAND2_X1   g01889(.A1(new_n2081_), .A2(new_n1096_), .ZN(new_n2082_));
  INV_X1     g01890(.I(new_n2082_), .ZN(new_n2083_));
  AOI21_X1   g01891(.A1(new_n2078_), .A2(new_n2083_), .B(new_n2077_), .ZN(new_n2084_));
  AOI21_X1   g01892(.A1(new_n2077_), .A2(new_n2078_), .B(new_n1096_), .ZN(new_n2085_));
  NOR4_X1    g01893(.A1(new_n2046_), .A2(\asqrt[53] ), .A3(new_n1876_), .A4(new_n1971_), .ZN(new_n2086_));
  XOR2_X1    g01894(.A1(new_n2086_), .A2(new_n1905_), .Z(new_n2087_));
  NAND2_X1   g01895(.A1(new_n2087_), .A2(new_n970_), .ZN(new_n2088_));
  OAI21_X1   g01896(.A1(new_n2085_), .A2(new_n2088_), .B(new_n2084_), .ZN(new_n2089_));
  OAI21_X1   g01897(.A1(new_n2084_), .A2(new_n2085_), .B(\asqrt[54] ), .ZN(new_n2090_));
  NOR4_X1    g01898(.A1(new_n2046_), .A2(\asqrt[54] ), .A3(new_n1883_), .A4(new_n1913_), .ZN(new_n2091_));
  XOR2_X1    g01899(.A1(new_n2091_), .A2(new_n1907_), .Z(new_n2092_));
  NAND2_X1   g01900(.A1(new_n2092_), .A2(new_n825_), .ZN(new_n2093_));
  INV_X1     g01901(.I(new_n2093_), .ZN(new_n2094_));
  AOI21_X1   g01902(.A1(new_n2090_), .A2(new_n2094_), .B(new_n2089_), .ZN(new_n2095_));
  AOI21_X1   g01903(.A1(new_n2089_), .A2(new_n2090_), .B(new_n825_), .ZN(new_n2096_));
  NOR4_X1    g01904(.A1(new_n2046_), .A2(\asqrt[55] ), .A3(new_n1909_), .A4(new_n1975_), .ZN(new_n2097_));
  XOR2_X1    g01905(.A1(new_n2097_), .A2(new_n1923_), .Z(new_n2098_));
  NAND2_X1   g01906(.A1(new_n2098_), .A2(new_n724_), .ZN(new_n2099_));
  OAI21_X1   g01907(.A1(new_n2096_), .A2(new_n2099_), .B(new_n2095_), .ZN(new_n2100_));
  OAI21_X1   g01908(.A1(new_n2095_), .A2(new_n2096_), .B(\asqrt[56] ), .ZN(new_n2101_));
  NOR4_X1    g01909(.A1(new_n2046_), .A2(\asqrt[56] ), .A3(new_n1916_), .A4(new_n1924_), .ZN(new_n2102_));
  XOR2_X1    g01910(.A1(new_n2102_), .A2(new_n2032_), .Z(new_n2103_));
  NAND2_X1   g01911(.A1(new_n2103_), .A2(new_n587_), .ZN(new_n2104_));
  INV_X1     g01912(.I(new_n2104_), .ZN(new_n2105_));
  AOI21_X1   g01913(.A1(new_n2101_), .A2(new_n2105_), .B(new_n2100_), .ZN(new_n2106_));
  AOI22_X1   g01914(.A1(new_n2068_), .A2(new_n2065_), .B1(\asqrt[50] ), .B2(new_n2054_), .ZN(new_n2107_));
  OAI21_X1   g01915(.A1(new_n2107_), .A2(new_n1436_), .B(new_n2075_), .ZN(new_n2108_));
  OAI22_X1   g01916(.A1(new_n2107_), .A2(new_n1436_), .B1(new_n2069_), .B2(new_n2063_), .ZN(new_n2109_));
  AOI22_X1   g01917(.A1(new_n2109_), .A2(\asqrt[52] ), .B1(new_n2108_), .B2(new_n2064_), .ZN(new_n2110_));
  INV_X1     g01918(.I(new_n2088_), .ZN(new_n2111_));
  OAI21_X1   g01919(.A1(new_n2110_), .A2(new_n1096_), .B(new_n2111_), .ZN(new_n2112_));
  AOI21_X1   g01920(.A1(new_n2109_), .A2(\asqrt[52] ), .B(new_n2082_), .ZN(new_n2113_));
  OAI22_X1   g01921(.A1(new_n2110_), .A2(new_n1096_), .B1(new_n2113_), .B2(new_n2077_), .ZN(new_n2114_));
  AOI22_X1   g01922(.A1(new_n2114_), .A2(\asqrt[54] ), .B1(new_n2112_), .B2(new_n2084_), .ZN(new_n2115_));
  INV_X1     g01923(.I(new_n2099_), .ZN(new_n2116_));
  OAI21_X1   g01924(.A1(new_n2115_), .A2(new_n825_), .B(new_n2116_), .ZN(new_n2117_));
  AOI21_X1   g01925(.A1(new_n2114_), .A2(\asqrt[54] ), .B(new_n2093_), .ZN(new_n2118_));
  OAI22_X1   g01926(.A1(new_n2115_), .A2(new_n825_), .B1(new_n2118_), .B2(new_n2089_), .ZN(new_n2119_));
  AOI22_X1   g01927(.A1(new_n2119_), .A2(\asqrt[56] ), .B1(new_n2117_), .B2(new_n2095_), .ZN(new_n2120_));
  NOR4_X1    g01928(.A1(new_n2046_), .A2(\asqrt[57] ), .A3(new_n1926_), .A4(new_n1981_), .ZN(new_n2121_));
  XOR2_X1    g01929(.A1(new_n2121_), .A2(new_n1932_), .Z(new_n2122_));
  NAND2_X1   g01930(.A1(new_n2122_), .A2(new_n504_), .ZN(new_n2123_));
  INV_X1     g01931(.I(new_n2123_), .ZN(new_n2124_));
  OAI21_X1   g01932(.A1(new_n2120_), .A2(new_n587_), .B(new_n2124_), .ZN(new_n2125_));
  NAND2_X1   g01933(.A1(new_n2125_), .A2(new_n2106_), .ZN(new_n2126_));
  AOI21_X1   g01934(.A1(new_n2119_), .A2(\asqrt[56] ), .B(new_n2104_), .ZN(new_n2127_));
  OAI22_X1   g01935(.A1(new_n2120_), .A2(new_n587_), .B1(new_n2127_), .B2(new_n2100_), .ZN(new_n2128_));
  NOR4_X1    g01936(.A1(new_n2046_), .A2(\asqrt[58] ), .A3(new_n1934_), .A4(new_n1940_), .ZN(new_n2129_));
  XOR2_X1    g01937(.A1(new_n2129_), .A2(new_n2034_), .Z(new_n2130_));
  NAND2_X1   g01938(.A1(new_n2130_), .A2(new_n376_), .ZN(new_n2131_));
  AOI21_X1   g01939(.A1(new_n2128_), .A2(\asqrt[58] ), .B(new_n2131_), .ZN(new_n2132_));
  NOR2_X1    g01940(.A1(new_n2132_), .A2(new_n2126_), .ZN(new_n2133_));
  AOI22_X1   g01941(.A1(new_n2128_), .A2(\asqrt[58] ), .B1(new_n2125_), .B2(new_n2106_), .ZN(new_n2134_));
  NOR4_X1    g01942(.A1(new_n2046_), .A2(\asqrt[59] ), .A3(new_n1942_), .A4(new_n1988_), .ZN(new_n2135_));
  XOR2_X1    g01943(.A1(new_n2135_), .A2(new_n2021_), .Z(new_n2136_));
  NAND2_X1   g01944(.A1(new_n2136_), .A2(new_n275_), .ZN(new_n2137_));
  INV_X1     g01945(.I(new_n2137_), .ZN(new_n2138_));
  OAI21_X1   g01946(.A1(new_n2134_), .A2(new_n376_), .B(new_n2138_), .ZN(new_n2139_));
  NAND2_X1   g01947(.A1(new_n2139_), .A2(new_n2133_), .ZN(new_n2140_));
  AOI21_X1   g01948(.A1(new_n2100_), .A2(new_n2101_), .B(new_n587_), .ZN(new_n2141_));
  OAI21_X1   g01949(.A1(new_n2106_), .A2(new_n2141_), .B(\asqrt[58] ), .ZN(new_n2142_));
  AOI21_X1   g01950(.A1(new_n2126_), .A2(new_n2142_), .B(new_n376_), .ZN(new_n2143_));
  OAI21_X1   g01951(.A1(new_n2133_), .A2(new_n2143_), .B(\asqrt[60] ), .ZN(new_n2144_));
  AOI21_X1   g01952(.A1(new_n2140_), .A2(new_n2144_), .B(new_n229_), .ZN(new_n2145_));
  NAND2_X1   g01953(.A1(new_n2014_), .A2(\asqrt[62] ), .ZN(new_n2146_));
  NOR2_X1    g01954(.A1(new_n2014_), .A2(\asqrt[62] ), .ZN(new_n2147_));
  NAND2_X1   g01955(.A1(new_n2147_), .A2(new_n1960_), .ZN(new_n2148_));
  NOR3_X1    g01956(.A1(new_n2046_), .A2(new_n2146_), .A3(new_n2148_), .ZN(new_n2149_));
  NOR2_X1    g01957(.A1(new_n2147_), .A2(new_n1960_), .ZN(new_n2150_));
  AOI21_X1   g01958(.A1(new_n2046_), .A2(new_n2150_), .B(new_n2146_), .ZN(new_n2151_));
  NOR2_X1    g01959(.A1(new_n2149_), .A2(new_n2151_), .ZN(new_n2152_));
  NOR3_X1    g01960(.A1(new_n1994_), .A2(\asqrt[61] ), .A3(new_n1955_), .ZN(new_n2153_));
  NAND2_X1   g01961(.A1(\asqrt[48] ), .A2(new_n2153_), .ZN(new_n2154_));
  XOR2_X1    g01962(.A1(new_n2154_), .A2(new_n2037_), .Z(new_n2155_));
  NOR2_X1    g01963(.A1(new_n2155_), .A2(new_n196_), .ZN(new_n2156_));
  INV_X1     g01964(.I(new_n2156_), .ZN(new_n2157_));
  NOR2_X1    g01965(.A1(new_n2050_), .A2(new_n2019_), .ZN(new_n2158_));
  NOR3_X1    g01966(.A1(new_n2018_), .A2(new_n2006_), .A3(new_n2030_), .ZN(new_n2159_));
  NAND4_X1   g01967(.A1(new_n2039_), .A2(new_n2015_), .A3(new_n1967_), .A4(new_n1999_), .ZN(new_n2160_));
  NOR4_X1    g01968(.A1(new_n2160_), .A2(new_n1810_), .A3(new_n1849_), .A4(new_n2058_), .ZN(new_n2161_));
  AOI21_X1   g01969(.A1(\asqrt[48] ), .A2(new_n2059_), .B(new_n1890_), .ZN(new_n2162_));
  NOR3_X1    g01970(.A1(new_n2162_), .A2(\asqrt[51] ), .A3(new_n2161_), .ZN(new_n2163_));
  OAI21_X1   g01971(.A1(new_n2159_), .A2(new_n1595_), .B(new_n2163_), .ZN(new_n2164_));
  NAND2_X1   g01972(.A1(new_n2158_), .A2(new_n2164_), .ZN(new_n2165_));
  NOR2_X1    g01973(.A1(new_n2159_), .A2(new_n1595_), .ZN(new_n2166_));
  OAI21_X1   g01974(.A1(new_n2158_), .A2(new_n2166_), .B(\asqrt[51] ), .ZN(new_n2167_));
  AOI21_X1   g01975(.A1(new_n2167_), .A2(new_n2075_), .B(new_n2165_), .ZN(new_n2168_));
  AOI21_X1   g01976(.A1(new_n2167_), .A2(new_n2165_), .B(new_n1260_), .ZN(new_n2169_));
  OAI21_X1   g01977(.A1(new_n2169_), .A2(new_n2082_), .B(new_n2168_), .ZN(new_n2170_));
  OAI21_X1   g01978(.A1(new_n2168_), .A2(new_n2169_), .B(\asqrt[53] ), .ZN(new_n2171_));
  AOI21_X1   g01979(.A1(new_n2171_), .A2(new_n2111_), .B(new_n2170_), .ZN(new_n2172_));
  AOI21_X1   g01980(.A1(new_n2170_), .A2(new_n2171_), .B(new_n970_), .ZN(new_n2173_));
  OAI21_X1   g01981(.A1(new_n2173_), .A2(new_n2093_), .B(new_n2172_), .ZN(new_n2174_));
  OAI21_X1   g01982(.A1(new_n2172_), .A2(new_n2173_), .B(\asqrt[55] ), .ZN(new_n2175_));
  AOI21_X1   g01983(.A1(new_n2175_), .A2(new_n2116_), .B(new_n2174_), .ZN(new_n2176_));
  AOI21_X1   g01984(.A1(new_n2174_), .A2(new_n2175_), .B(new_n724_), .ZN(new_n2177_));
  OAI21_X1   g01985(.A1(new_n2177_), .A2(new_n2104_), .B(new_n2176_), .ZN(new_n2178_));
  OAI21_X1   g01986(.A1(new_n2176_), .A2(new_n2177_), .B(\asqrt[57] ), .ZN(new_n2179_));
  AOI21_X1   g01987(.A1(new_n2179_), .A2(new_n2124_), .B(new_n2178_), .ZN(new_n2180_));
  AOI21_X1   g01988(.A1(new_n2178_), .A2(new_n2179_), .B(new_n504_), .ZN(new_n2181_));
  OAI21_X1   g01989(.A1(new_n2181_), .A2(new_n2131_), .B(new_n2180_), .ZN(new_n2182_));
  OAI21_X1   g01990(.A1(new_n2180_), .A2(new_n2181_), .B(\asqrt[59] ), .ZN(new_n2183_));
  AOI21_X1   g01991(.A1(new_n2183_), .A2(new_n2138_), .B(new_n2182_), .ZN(new_n2184_));
  INV_X1     g01992(.I(new_n2131_), .ZN(new_n2185_));
  NAND2_X1   g01993(.A1(new_n2142_), .A2(new_n2185_), .ZN(new_n2186_));
  NAND2_X1   g01994(.A1(new_n2126_), .A2(new_n2142_), .ZN(new_n2187_));
  AOI22_X1   g01995(.A1(new_n2187_), .A2(\asqrt[59] ), .B1(new_n2186_), .B2(new_n2180_), .ZN(new_n2188_));
  NOR4_X1    g01996(.A1(new_n2046_), .A2(\asqrt[60] ), .A3(new_n1948_), .A4(new_n1953_), .ZN(new_n2189_));
  XOR2_X1    g01997(.A1(new_n2189_), .A2(new_n2036_), .Z(new_n2190_));
  NAND2_X1   g01998(.A1(new_n2190_), .A2(new_n229_), .ZN(new_n2191_));
  INV_X1     g01999(.I(new_n2191_), .ZN(new_n2192_));
  OAI21_X1   g02000(.A1(new_n2188_), .A2(new_n275_), .B(new_n2192_), .ZN(new_n2193_));
  NAND2_X1   g02001(.A1(new_n2193_), .A2(new_n2184_), .ZN(new_n2194_));
  INV_X1     g02002(.I(new_n2155_), .ZN(new_n2195_));
  NOR2_X1    g02003(.A1(new_n2195_), .A2(\asqrt[62] ), .ZN(new_n2196_));
  INV_X1     g02004(.I(new_n2196_), .ZN(new_n2197_));
  NAND2_X1   g02005(.A1(new_n2145_), .A2(new_n2197_), .ZN(new_n2198_));
  OAI21_X1   g02006(.A1(new_n2198_), .A2(new_n2194_), .B(new_n2157_), .ZN(new_n2199_));
  NAND2_X1   g02007(.A1(new_n1996_), .A2(new_n1823_), .ZN(new_n2200_));
  OAI21_X1   g02008(.A1(\asqrt[48] ), .A2(new_n2200_), .B(new_n2011_), .ZN(new_n2201_));
  NAND2_X1   g02009(.A1(new_n2201_), .A2(new_n231_), .ZN(new_n2202_));
  OAI21_X1   g02010(.A1(new_n2199_), .A2(new_n2202_), .B(new_n2152_), .ZN(new_n2203_));
  OAI21_X1   g02011(.A1(new_n1967_), .A2(new_n2011_), .B(\asqrt[48] ), .ZN(new_n2204_));
  XOR2_X1    g02012(.A1(new_n2011_), .A2(\asqrt[63] ), .Z(new_n2205_));
  NAND2_X1   g02013(.A1(new_n2204_), .A2(new_n2205_), .ZN(new_n2206_));
  INV_X1     g02014(.I(new_n2206_), .ZN(new_n2207_));
  INV_X1     g02015(.I(new_n2152_), .ZN(new_n2208_));
  OAI22_X1   g02016(.A1(new_n2134_), .A2(new_n376_), .B1(new_n2132_), .B2(new_n2126_), .ZN(new_n2209_));
  AOI21_X1   g02017(.A1(new_n2209_), .A2(\asqrt[60] ), .B(new_n2191_), .ZN(new_n2210_));
  AOI22_X1   g02018(.A1(new_n2209_), .A2(\asqrt[60] ), .B1(new_n2139_), .B2(new_n2133_), .ZN(new_n2211_));
  OAI22_X1   g02019(.A1(new_n2211_), .A2(new_n229_), .B1(new_n2210_), .B2(new_n2140_), .ZN(new_n2212_));
  NOR4_X1    g02020(.A1(new_n2212_), .A2(\asqrt[62] ), .A3(new_n2208_), .A4(new_n2155_), .ZN(new_n2213_));
  NAND2_X1   g02021(.A1(new_n2213_), .A2(new_n2207_), .ZN(new_n2214_));
  NOR2_X1    g02022(.A1(new_n1823_), .A2(new_n1811_), .ZN(new_n2215_));
  NAND2_X1   g02023(.A1(new_n2026_), .A2(new_n2215_), .ZN(new_n2216_));
  NOR3_X1    g02024(.A1(new_n2214_), .A2(new_n2203_), .A3(new_n2216_), .ZN(\asqrt[47] ));
  NAND2_X1   g02025(.A1(new_n2140_), .A2(new_n2144_), .ZN(new_n2218_));
  NOR3_X1    g02026(.A1(new_n2218_), .A2(\asqrt[61] ), .A3(new_n2190_), .ZN(new_n2219_));
  NAND2_X1   g02027(.A1(\asqrt[47] ), .A2(new_n2219_), .ZN(new_n2220_));
  XOR2_X1    g02028(.A1(new_n2220_), .A2(new_n2145_), .Z(new_n2221_));
  INV_X1     g02029(.I(new_n2221_), .ZN(new_n2222_));
  INV_X1     g02030(.I(\a[95] ), .ZN(new_n2223_));
  INV_X1     g02031(.I(\a[94] ), .ZN(new_n2224_));
  NOR2_X1    g02032(.A1(\a[92] ), .A2(\a[93] ), .ZN(new_n2225_));
  INV_X1     g02033(.I(new_n2225_), .ZN(new_n2226_));
  NOR4_X1    g02034(.A1(new_n2047_), .A2(new_n2224_), .A3(new_n2041_), .A4(new_n2226_), .ZN(new_n2227_));
  XOR2_X1    g02035(.A1(new_n2227_), .A2(new_n2223_), .Z(new_n2228_));
  NOR4_X1    g02036(.A1(new_n2214_), .A2(new_n2203_), .A3(new_n2223_), .A4(new_n2216_), .ZN(new_n2229_));
  NOR2_X1    g02037(.A1(new_n2223_), .A2(\a[94] ), .ZN(new_n2230_));
  OAI21_X1   g02038(.A1(new_n2229_), .A2(new_n2230_), .B(new_n2228_), .ZN(new_n2231_));
  INV_X1     g02039(.I(new_n2228_), .ZN(new_n2232_));
  NOR2_X1    g02040(.A1(new_n2210_), .A2(new_n2140_), .ZN(new_n2233_));
  NOR3_X1    g02041(.A1(new_n2211_), .A2(new_n229_), .A3(new_n2196_), .ZN(new_n2234_));
  AOI21_X1   g02042(.A1(new_n2234_), .A2(new_n2233_), .B(new_n2156_), .ZN(new_n2235_));
  INV_X1     g02043(.I(new_n2202_), .ZN(new_n2236_));
  AOI21_X1   g02044(.A1(new_n2235_), .A2(new_n2236_), .B(new_n2208_), .ZN(new_n2237_));
  AOI21_X1   g02045(.A1(new_n2212_), .A2(\asqrt[62] ), .B(new_n2152_), .ZN(new_n2238_));
  AOI21_X1   g02046(.A1(new_n2182_), .A2(new_n2183_), .B(new_n275_), .ZN(new_n2239_));
  OAI21_X1   g02047(.A1(new_n2184_), .A2(new_n2239_), .B(\asqrt[61] ), .ZN(new_n2240_));
  NAND4_X1   g02048(.A1(new_n2194_), .A2(new_n196_), .A3(new_n2240_), .A4(new_n2195_), .ZN(new_n2241_));
  NOR3_X1    g02049(.A1(new_n2238_), .A2(new_n2206_), .A3(new_n2241_), .ZN(new_n2242_));
  INV_X1     g02050(.I(new_n2216_), .ZN(new_n2243_));
  NAND4_X1   g02051(.A1(new_n2242_), .A2(\a[95] ), .A3(new_n2237_), .A4(new_n2243_), .ZN(new_n2244_));
  NAND3_X1   g02052(.A1(new_n2244_), .A2(\a[94] ), .A3(new_n2232_), .ZN(new_n2245_));
  NAND2_X1   g02053(.A1(new_n2231_), .A2(new_n2245_), .ZN(new_n2246_));
  NOR2_X1    g02054(.A1(new_n2214_), .A2(new_n2203_), .ZN(new_n2247_));
  NOR4_X1    g02055(.A1(new_n2016_), .A2(new_n1810_), .A3(new_n1823_), .A4(new_n2025_), .ZN(new_n2248_));
  NAND2_X1   g02056(.A1(\asqrt[48] ), .A2(\a[94] ), .ZN(new_n2249_));
  XOR2_X1    g02057(.A1(new_n2249_), .A2(new_n2248_), .Z(new_n2250_));
  NOR2_X1    g02058(.A1(new_n2250_), .A2(new_n2226_), .ZN(new_n2251_));
  INV_X1     g02059(.I(new_n2251_), .ZN(new_n2252_));
  NAND3_X1   g02060(.A1(new_n2242_), .A2(new_n2237_), .A3(new_n2243_), .ZN(new_n2253_));
  NOR4_X1    g02061(.A1(new_n2240_), .A2(new_n2140_), .A3(new_n2210_), .A4(new_n2196_), .ZN(new_n2254_));
  NOR3_X1    g02062(.A1(new_n2254_), .A2(new_n2156_), .A3(new_n2202_), .ZN(new_n2255_));
  AOI22_X1   g02063(.A1(new_n2218_), .A2(\asqrt[61] ), .B1(new_n2193_), .B2(new_n2184_), .ZN(new_n2256_));
  NAND4_X1   g02064(.A1(new_n2256_), .A2(new_n196_), .A3(new_n2152_), .A4(new_n2195_), .ZN(new_n2257_));
  OAI21_X1   g02065(.A1(new_n2255_), .A2(new_n2208_), .B(new_n2257_), .ZN(new_n2258_));
  NOR2_X1    g02066(.A1(new_n2207_), .A2(new_n2243_), .ZN(new_n2259_));
  NAND2_X1   g02067(.A1(new_n2259_), .A2(\asqrt[48] ), .ZN(new_n2260_));
  OAI21_X1   g02068(.A1(new_n2258_), .A2(new_n2260_), .B(new_n1738_), .ZN(new_n2261_));
  NAND3_X1   g02069(.A1(new_n2261_), .A2(new_n1746_), .A3(new_n2253_), .ZN(new_n2262_));
  NAND4_X1   g02070(.A1(new_n2145_), .A2(new_n2184_), .A3(new_n2193_), .A4(new_n2197_), .ZN(new_n2263_));
  NAND3_X1   g02071(.A1(new_n2263_), .A2(new_n2157_), .A3(new_n2236_), .ZN(new_n2264_));
  AOI21_X1   g02072(.A1(new_n2152_), .A2(new_n2264_), .B(new_n2213_), .ZN(new_n2265_));
  INV_X1     g02073(.I(new_n2260_), .ZN(new_n2266_));
  AOI21_X1   g02074(.A1(new_n2265_), .A2(new_n2266_), .B(\a[96] ), .ZN(new_n2267_));
  OAI21_X1   g02075(.A1(new_n2267_), .A2(new_n1747_), .B(\asqrt[47] ), .ZN(new_n2268_));
  NAND4_X1   g02076(.A1(new_n2262_), .A2(new_n2268_), .A3(new_n1854_), .A4(new_n2252_), .ZN(new_n2269_));
  NAND2_X1   g02077(.A1(new_n2269_), .A2(new_n2246_), .ZN(new_n2270_));
  NAND3_X1   g02078(.A1(new_n2231_), .A2(new_n2245_), .A3(new_n2252_), .ZN(new_n2271_));
  AOI21_X1   g02079(.A1(\asqrt[48] ), .A2(new_n1738_), .B(\a[97] ), .ZN(new_n2272_));
  NOR2_X1    g02080(.A1(new_n2002_), .A2(\a[96] ), .ZN(new_n2273_));
  AOI21_X1   g02081(.A1(\asqrt[48] ), .A2(\a[96] ), .B(new_n1749_), .ZN(new_n2274_));
  OAI21_X1   g02082(.A1(new_n2272_), .A2(new_n2273_), .B(new_n2274_), .ZN(new_n2275_));
  INV_X1     g02083(.I(new_n2275_), .ZN(new_n2276_));
  NAND3_X1   g02084(.A1(\asqrt[47] ), .A2(new_n2053_), .A3(new_n2276_), .ZN(new_n2277_));
  OAI21_X1   g02085(.A1(new_n2253_), .A2(new_n2275_), .B(new_n2030_), .ZN(new_n2278_));
  NAND3_X1   g02086(.A1(new_n2277_), .A2(new_n2278_), .A3(new_n1595_), .ZN(new_n2279_));
  AOI21_X1   g02087(.A1(new_n2271_), .A2(\asqrt[49] ), .B(new_n2279_), .ZN(new_n2280_));
  NOR2_X1    g02088(.A1(new_n2270_), .A2(new_n2280_), .ZN(new_n2281_));
  AOI22_X1   g02089(.A1(new_n2269_), .A2(new_n2246_), .B1(\asqrt[49] ), .B2(new_n2271_), .ZN(new_n2282_));
  AOI21_X1   g02090(.A1(new_n2067_), .A2(new_n2066_), .B(\asqrt[50] ), .ZN(new_n2283_));
  NAND2_X1   g02091(.A1(new_n2283_), .A2(new_n2159_), .ZN(new_n2284_));
  NOR3_X1    g02092(.A1(new_n2253_), .A2(new_n2166_), .A3(new_n2284_), .ZN(new_n2285_));
  NOR2_X1    g02093(.A1(new_n2159_), .A2(new_n1595_), .ZN(new_n2286_));
  NOR2_X1    g02094(.A1(new_n2285_), .A2(new_n2286_), .ZN(new_n2287_));
  NAND2_X1   g02095(.A1(new_n2287_), .A2(new_n1436_), .ZN(new_n2288_));
  INV_X1     g02096(.I(new_n2288_), .ZN(new_n2289_));
  OAI21_X1   g02097(.A1(new_n2282_), .A2(new_n1595_), .B(new_n2289_), .ZN(new_n2290_));
  NAND2_X1   g02098(.A1(new_n2290_), .A2(new_n2281_), .ZN(new_n2291_));
  OAI22_X1   g02099(.A1(new_n2282_), .A2(new_n1595_), .B1(new_n2270_), .B2(new_n2280_), .ZN(new_n2292_));
  NAND2_X1   g02100(.A1(new_n2061_), .A2(new_n2060_), .ZN(new_n2293_));
  NAND4_X1   g02101(.A1(\asqrt[47] ), .A2(new_n1436_), .A3(new_n2293_), .A4(new_n2107_), .ZN(new_n2294_));
  XOR2_X1    g02102(.A1(new_n2294_), .A2(new_n2071_), .Z(new_n2295_));
  NAND2_X1   g02103(.A1(new_n2295_), .A2(new_n1260_), .ZN(new_n2296_));
  AOI21_X1   g02104(.A1(new_n2292_), .A2(\asqrt[51] ), .B(new_n2296_), .ZN(new_n2297_));
  NOR2_X1    g02105(.A1(new_n2297_), .A2(new_n2291_), .ZN(new_n2298_));
  AOI22_X1   g02106(.A1(new_n2292_), .A2(\asqrt[51] ), .B1(new_n2290_), .B2(new_n2281_), .ZN(new_n2299_));
  NOR2_X1    g02107(.A1(new_n2073_), .A2(new_n2074_), .ZN(new_n2300_));
  NOR4_X1    g02108(.A1(new_n2253_), .A2(\asqrt[52] ), .A3(new_n2300_), .A4(new_n2109_), .ZN(new_n2301_));
  XOR2_X1    g02109(.A1(new_n2301_), .A2(new_n2078_), .Z(new_n2302_));
  NAND2_X1   g02110(.A1(new_n2302_), .A2(new_n1096_), .ZN(new_n2303_));
  INV_X1     g02111(.I(new_n2303_), .ZN(new_n2304_));
  OAI21_X1   g02112(.A1(new_n2299_), .A2(new_n1260_), .B(new_n2304_), .ZN(new_n2305_));
  NAND2_X1   g02113(.A1(new_n2305_), .A2(new_n2298_), .ZN(new_n2306_));
  OAI22_X1   g02114(.A1(new_n2299_), .A2(new_n1260_), .B1(new_n2297_), .B2(new_n2291_), .ZN(new_n2307_));
  INV_X1     g02115(.I(new_n2110_), .ZN(new_n2308_));
  NOR4_X1    g02116(.A1(new_n2253_), .A2(\asqrt[53] ), .A3(new_n2081_), .A4(new_n2308_), .ZN(new_n2309_));
  XOR2_X1    g02117(.A1(new_n2309_), .A2(new_n2171_), .Z(new_n2310_));
  NAND2_X1   g02118(.A1(new_n2310_), .A2(new_n970_), .ZN(new_n2311_));
  AOI21_X1   g02119(.A1(new_n2307_), .A2(\asqrt[53] ), .B(new_n2311_), .ZN(new_n2312_));
  NOR2_X1    g02120(.A1(new_n2312_), .A2(new_n2306_), .ZN(new_n2313_));
  AOI22_X1   g02121(.A1(new_n2307_), .A2(\asqrt[53] ), .B1(new_n2305_), .B2(new_n2298_), .ZN(new_n2314_));
  NOR4_X1    g02122(.A1(new_n2253_), .A2(\asqrt[54] ), .A3(new_n2087_), .A4(new_n2114_), .ZN(new_n2315_));
  XOR2_X1    g02123(.A1(new_n2315_), .A2(new_n2090_), .Z(new_n2316_));
  NAND2_X1   g02124(.A1(new_n2316_), .A2(new_n825_), .ZN(new_n2317_));
  INV_X1     g02125(.I(new_n2317_), .ZN(new_n2318_));
  OAI21_X1   g02126(.A1(new_n2314_), .A2(new_n970_), .B(new_n2318_), .ZN(new_n2319_));
  NAND2_X1   g02127(.A1(new_n2319_), .A2(new_n2313_), .ZN(new_n2320_));
  OAI22_X1   g02128(.A1(new_n2314_), .A2(new_n970_), .B1(new_n2312_), .B2(new_n2306_), .ZN(new_n2321_));
  INV_X1     g02129(.I(new_n2115_), .ZN(new_n2322_));
  NOR4_X1    g02130(.A1(new_n2253_), .A2(\asqrt[55] ), .A3(new_n2092_), .A4(new_n2322_), .ZN(new_n2323_));
  XOR2_X1    g02131(.A1(new_n2323_), .A2(new_n2175_), .Z(new_n2324_));
  NAND2_X1   g02132(.A1(new_n2324_), .A2(new_n724_), .ZN(new_n2325_));
  AOI21_X1   g02133(.A1(new_n2321_), .A2(\asqrt[55] ), .B(new_n2325_), .ZN(new_n2326_));
  NOR2_X1    g02134(.A1(new_n2326_), .A2(new_n2320_), .ZN(new_n2327_));
  AOI22_X1   g02135(.A1(new_n2321_), .A2(\asqrt[55] ), .B1(new_n2319_), .B2(new_n2313_), .ZN(new_n2328_));
  NOR4_X1    g02136(.A1(new_n2253_), .A2(\asqrt[56] ), .A3(new_n2098_), .A4(new_n2119_), .ZN(new_n2329_));
  XOR2_X1    g02137(.A1(new_n2329_), .A2(new_n2101_), .Z(new_n2330_));
  NAND2_X1   g02138(.A1(new_n2330_), .A2(new_n587_), .ZN(new_n2331_));
  INV_X1     g02139(.I(new_n2331_), .ZN(new_n2332_));
  OAI21_X1   g02140(.A1(new_n2328_), .A2(new_n724_), .B(new_n2332_), .ZN(new_n2333_));
  NAND2_X1   g02141(.A1(new_n2333_), .A2(new_n2327_), .ZN(new_n2334_));
  OAI22_X1   g02142(.A1(new_n2328_), .A2(new_n724_), .B1(new_n2326_), .B2(new_n2320_), .ZN(new_n2335_));
  INV_X1     g02143(.I(new_n2120_), .ZN(new_n2336_));
  NOR4_X1    g02144(.A1(new_n2253_), .A2(\asqrt[57] ), .A3(new_n2103_), .A4(new_n2336_), .ZN(new_n2337_));
  XOR2_X1    g02145(.A1(new_n2337_), .A2(new_n2179_), .Z(new_n2338_));
  NAND2_X1   g02146(.A1(new_n2338_), .A2(new_n504_), .ZN(new_n2339_));
  AOI21_X1   g02147(.A1(new_n2335_), .A2(\asqrt[57] ), .B(new_n2339_), .ZN(new_n2340_));
  NOR2_X1    g02148(.A1(new_n2340_), .A2(new_n2334_), .ZN(new_n2341_));
  AOI22_X1   g02149(.A1(new_n2335_), .A2(\asqrt[57] ), .B1(new_n2333_), .B2(new_n2327_), .ZN(new_n2342_));
  NOR4_X1    g02150(.A1(new_n2253_), .A2(\asqrt[58] ), .A3(new_n2122_), .A4(new_n2128_), .ZN(new_n2343_));
  XOR2_X1    g02151(.A1(new_n2343_), .A2(new_n2142_), .Z(new_n2344_));
  NAND2_X1   g02152(.A1(new_n2344_), .A2(new_n376_), .ZN(new_n2345_));
  INV_X1     g02153(.I(new_n2345_), .ZN(new_n2346_));
  OAI21_X1   g02154(.A1(new_n2342_), .A2(new_n504_), .B(new_n2346_), .ZN(new_n2347_));
  NAND2_X1   g02155(.A1(new_n2347_), .A2(new_n2341_), .ZN(new_n2348_));
  OAI22_X1   g02156(.A1(new_n2342_), .A2(new_n504_), .B1(new_n2340_), .B2(new_n2334_), .ZN(new_n2349_));
  NOR4_X1    g02157(.A1(new_n2253_), .A2(\asqrt[59] ), .A3(new_n2130_), .A4(new_n2187_), .ZN(new_n2350_));
  XOR2_X1    g02158(.A1(new_n2350_), .A2(new_n2183_), .Z(new_n2351_));
  NAND2_X1   g02159(.A1(new_n2351_), .A2(new_n275_), .ZN(new_n2352_));
  AOI21_X1   g02160(.A1(new_n2349_), .A2(\asqrt[59] ), .B(new_n2352_), .ZN(new_n2353_));
  NOR2_X1    g02161(.A1(new_n2353_), .A2(new_n2348_), .ZN(new_n2354_));
  AOI22_X1   g02162(.A1(new_n2349_), .A2(\asqrt[59] ), .B1(new_n2347_), .B2(new_n2341_), .ZN(new_n2355_));
  OAI22_X1   g02163(.A1(new_n2355_), .A2(new_n275_), .B1(new_n2353_), .B2(new_n2348_), .ZN(new_n2356_));
  NOR4_X1    g02164(.A1(new_n2253_), .A2(\asqrt[60] ), .A3(new_n2136_), .A4(new_n2209_), .ZN(new_n2357_));
  XOR2_X1    g02165(.A1(new_n2357_), .A2(new_n2144_), .Z(new_n2358_));
  NAND2_X1   g02166(.A1(new_n2358_), .A2(new_n229_), .ZN(new_n2359_));
  INV_X1     g02167(.I(new_n2359_), .ZN(new_n2360_));
  OAI21_X1   g02168(.A1(new_n2355_), .A2(new_n275_), .B(new_n2360_), .ZN(new_n2361_));
  AOI22_X1   g02169(.A1(new_n2356_), .A2(\asqrt[61] ), .B1(new_n2361_), .B2(new_n2354_), .ZN(new_n2362_));
  NOR2_X1    g02170(.A1(new_n2362_), .A2(new_n196_), .ZN(new_n2363_));
  INV_X1     g02171(.I(new_n2230_), .ZN(new_n2364_));
  AOI21_X1   g02172(.A1(new_n2244_), .A2(new_n2364_), .B(new_n2232_), .ZN(new_n2365_));
  NOR3_X1    g02173(.A1(new_n2229_), .A2(new_n2224_), .A3(new_n2228_), .ZN(new_n2366_));
  NOR2_X1    g02174(.A1(new_n2366_), .A2(new_n2365_), .ZN(new_n2367_));
  NOR3_X1    g02175(.A1(new_n2267_), .A2(new_n1747_), .A3(\asqrt[47] ), .ZN(new_n2368_));
  AOI21_X1   g02176(.A1(new_n2261_), .A2(new_n1746_), .B(new_n2253_), .ZN(new_n2369_));
  NOR4_X1    g02177(.A1(new_n2369_), .A2(new_n2368_), .A3(\asqrt[49] ), .A4(new_n2251_), .ZN(new_n2370_));
  NOR2_X1    g02178(.A1(new_n2370_), .A2(new_n2367_), .ZN(new_n2371_));
  NOR3_X1    g02179(.A1(new_n2366_), .A2(new_n2365_), .A3(new_n2251_), .ZN(new_n2372_));
  NOR3_X1    g02180(.A1(new_n2253_), .A2(new_n2030_), .A3(new_n2275_), .ZN(new_n2373_));
  AOI21_X1   g02181(.A1(\asqrt[47] ), .A2(new_n2276_), .B(new_n2053_), .ZN(new_n2374_));
  NOR3_X1    g02182(.A1(new_n2374_), .A2(new_n2373_), .A3(\asqrt[50] ), .ZN(new_n2375_));
  OAI21_X1   g02183(.A1(new_n2372_), .A2(new_n1854_), .B(new_n2375_), .ZN(new_n2376_));
  NAND2_X1   g02184(.A1(new_n2371_), .A2(new_n2376_), .ZN(new_n2377_));
  OAI22_X1   g02185(.A1(new_n2370_), .A2(new_n2367_), .B1(new_n1854_), .B2(new_n2372_), .ZN(new_n2378_));
  AOI21_X1   g02186(.A1(new_n2378_), .A2(\asqrt[50] ), .B(new_n2288_), .ZN(new_n2379_));
  NOR2_X1    g02187(.A1(new_n2379_), .A2(new_n2377_), .ZN(new_n2380_));
  AOI22_X1   g02188(.A1(new_n2378_), .A2(\asqrt[50] ), .B1(new_n2371_), .B2(new_n2376_), .ZN(new_n2381_));
  INV_X1     g02189(.I(new_n2296_), .ZN(new_n2382_));
  OAI21_X1   g02190(.A1(new_n2381_), .A2(new_n1436_), .B(new_n2382_), .ZN(new_n2383_));
  NAND2_X1   g02191(.A1(new_n2383_), .A2(new_n2380_), .ZN(new_n2384_));
  OAI22_X1   g02192(.A1(new_n2381_), .A2(new_n1436_), .B1(new_n2379_), .B2(new_n2377_), .ZN(new_n2385_));
  AOI21_X1   g02193(.A1(new_n2385_), .A2(\asqrt[52] ), .B(new_n2303_), .ZN(new_n2386_));
  NOR2_X1    g02194(.A1(new_n2386_), .A2(new_n2384_), .ZN(new_n2387_));
  AOI22_X1   g02195(.A1(new_n2385_), .A2(\asqrt[52] ), .B1(new_n2383_), .B2(new_n2380_), .ZN(new_n2388_));
  INV_X1     g02196(.I(new_n2311_), .ZN(new_n2389_));
  OAI21_X1   g02197(.A1(new_n2388_), .A2(new_n1096_), .B(new_n2389_), .ZN(new_n2390_));
  NAND2_X1   g02198(.A1(new_n2390_), .A2(new_n2387_), .ZN(new_n2391_));
  OAI22_X1   g02199(.A1(new_n2388_), .A2(new_n1096_), .B1(new_n2386_), .B2(new_n2384_), .ZN(new_n2392_));
  AOI21_X1   g02200(.A1(new_n2392_), .A2(\asqrt[54] ), .B(new_n2317_), .ZN(new_n2393_));
  NOR2_X1    g02201(.A1(new_n2393_), .A2(new_n2391_), .ZN(new_n2394_));
  AOI22_X1   g02202(.A1(new_n2392_), .A2(\asqrt[54] ), .B1(new_n2390_), .B2(new_n2387_), .ZN(new_n2395_));
  INV_X1     g02203(.I(new_n2325_), .ZN(new_n2396_));
  OAI21_X1   g02204(.A1(new_n2395_), .A2(new_n825_), .B(new_n2396_), .ZN(new_n2397_));
  NAND2_X1   g02205(.A1(new_n2397_), .A2(new_n2394_), .ZN(new_n2398_));
  OAI22_X1   g02206(.A1(new_n2395_), .A2(new_n825_), .B1(new_n2393_), .B2(new_n2391_), .ZN(new_n2399_));
  AOI21_X1   g02207(.A1(new_n2399_), .A2(\asqrt[56] ), .B(new_n2331_), .ZN(new_n2400_));
  NOR2_X1    g02208(.A1(new_n2400_), .A2(new_n2398_), .ZN(new_n2401_));
  AOI22_X1   g02209(.A1(new_n2399_), .A2(\asqrt[56] ), .B1(new_n2397_), .B2(new_n2394_), .ZN(new_n2402_));
  INV_X1     g02210(.I(new_n2339_), .ZN(new_n2403_));
  OAI21_X1   g02211(.A1(new_n2402_), .A2(new_n587_), .B(new_n2403_), .ZN(new_n2404_));
  NAND2_X1   g02212(.A1(new_n2404_), .A2(new_n2401_), .ZN(new_n2405_));
  OAI22_X1   g02213(.A1(new_n2402_), .A2(new_n587_), .B1(new_n2400_), .B2(new_n2398_), .ZN(new_n2406_));
  AOI21_X1   g02214(.A1(new_n2406_), .A2(\asqrt[58] ), .B(new_n2345_), .ZN(new_n2407_));
  NOR2_X1    g02215(.A1(new_n2407_), .A2(new_n2405_), .ZN(new_n2408_));
  AOI22_X1   g02216(.A1(new_n2406_), .A2(\asqrt[58] ), .B1(new_n2404_), .B2(new_n2401_), .ZN(new_n2409_));
  INV_X1     g02217(.I(new_n2352_), .ZN(new_n2410_));
  OAI21_X1   g02218(.A1(new_n2409_), .A2(new_n376_), .B(new_n2410_), .ZN(new_n2411_));
  NAND2_X1   g02219(.A1(new_n2411_), .A2(new_n2408_), .ZN(new_n2412_));
  OAI22_X1   g02220(.A1(new_n2409_), .A2(new_n376_), .B1(new_n2407_), .B2(new_n2405_), .ZN(new_n2413_));
  AOI22_X1   g02221(.A1(new_n2413_), .A2(\asqrt[60] ), .B1(new_n2411_), .B2(new_n2408_), .ZN(new_n2414_));
  AOI21_X1   g02222(.A1(new_n2413_), .A2(\asqrt[60] ), .B(new_n2359_), .ZN(new_n2415_));
  OAI22_X1   g02223(.A1(new_n2414_), .A2(new_n229_), .B1(new_n2415_), .B2(new_n2412_), .ZN(new_n2416_));
  NOR2_X1    g02224(.A1(new_n2416_), .A2(\asqrt[62] ), .ZN(new_n2417_));
  NAND3_X1   g02225(.A1(new_n2247_), .A2(new_n2152_), .A3(new_n2216_), .ZN(new_n2418_));
  NOR2_X1    g02226(.A1(new_n2256_), .A2(new_n196_), .ZN(new_n2419_));
  INV_X1     g02227(.I(new_n2241_), .ZN(new_n2420_));
  NAND3_X1   g02228(.A1(\asqrt[47] ), .A2(new_n2419_), .A3(new_n2420_), .ZN(new_n2421_));
  OAI21_X1   g02229(.A1(new_n2212_), .A2(\asqrt[62] ), .B(new_n2155_), .ZN(new_n2422_));
  OAI21_X1   g02230(.A1(\asqrt[47] ), .A2(new_n2422_), .B(new_n2419_), .ZN(new_n2423_));
  NAND2_X1   g02231(.A1(new_n2423_), .A2(new_n2421_), .ZN(new_n2424_));
  INV_X1     g02232(.I(new_n2424_), .ZN(new_n2425_));
  NOR2_X1    g02233(.A1(new_n2221_), .A2(new_n196_), .ZN(new_n2426_));
  INV_X1     g02234(.I(new_n2426_), .ZN(new_n2427_));
  NAND2_X1   g02235(.A1(new_n2335_), .A2(\asqrt[57] ), .ZN(new_n2428_));
  AOI21_X1   g02236(.A1(new_n2428_), .A2(new_n2334_), .B(new_n504_), .ZN(new_n2429_));
  OAI21_X1   g02237(.A1(new_n2341_), .A2(new_n2429_), .B(\asqrt[59] ), .ZN(new_n2430_));
  AOI21_X1   g02238(.A1(new_n2348_), .A2(new_n2430_), .B(new_n275_), .ZN(new_n2431_));
  OAI21_X1   g02239(.A1(new_n2354_), .A2(new_n2431_), .B(\asqrt[61] ), .ZN(new_n2432_));
  NOR2_X1    g02240(.A1(new_n2222_), .A2(\asqrt[62] ), .ZN(new_n2433_));
  INV_X1     g02241(.I(new_n2433_), .ZN(new_n2434_));
  NAND3_X1   g02242(.A1(new_n2361_), .A2(new_n2354_), .A3(new_n2434_), .ZN(new_n2435_));
  OAI21_X1   g02243(.A1(new_n2435_), .A2(new_n2432_), .B(new_n2427_), .ZN(new_n2436_));
  NAND3_X1   g02244(.A1(new_n2253_), .A2(new_n2208_), .A3(new_n2257_), .ZN(new_n2437_));
  AOI21_X1   g02245(.A1(new_n2437_), .A2(new_n2199_), .B(\asqrt[63] ), .ZN(new_n2438_));
  INV_X1     g02246(.I(new_n2438_), .ZN(new_n2439_));
  OAI21_X1   g02247(.A1(new_n2436_), .A2(new_n2439_), .B(new_n2425_), .ZN(new_n2440_));
  NOR4_X1    g02248(.A1(new_n2416_), .A2(\asqrt[62] ), .A3(new_n2424_), .A4(new_n2221_), .ZN(new_n2441_));
  AOI21_X1   g02249(.A1(new_n2208_), .A2(new_n2235_), .B(new_n2253_), .ZN(new_n2442_));
  XOR2_X1    g02250(.A1(new_n2235_), .A2(\asqrt[63] ), .Z(new_n2443_));
  NOR2_X1    g02251(.A1(new_n2442_), .A2(new_n2443_), .ZN(new_n2444_));
  NAND2_X1   g02252(.A1(new_n2441_), .A2(new_n2444_), .ZN(new_n2445_));
  NOR3_X1    g02253(.A1(new_n2445_), .A2(new_n2418_), .A3(new_n2440_), .ZN(\asqrt[46] ));
  NAND4_X1   g02254(.A1(\asqrt[46] ), .A2(new_n2222_), .A3(new_n2363_), .A4(new_n2417_), .ZN(new_n2447_));
  OAI21_X1   g02255(.A1(new_n2416_), .A2(\asqrt[62] ), .B(new_n2221_), .ZN(new_n2448_));
  OAI21_X1   g02256(.A1(\asqrt[46] ), .A2(new_n2448_), .B(new_n2363_), .ZN(new_n2449_));
  NAND2_X1   g02257(.A1(new_n2447_), .A2(new_n2449_), .ZN(new_n2450_));
  INV_X1     g02258(.I(new_n2450_), .ZN(new_n2451_));
  NAND2_X1   g02259(.A1(new_n2406_), .A2(\asqrt[58] ), .ZN(new_n2452_));
  AOI21_X1   g02260(.A1(new_n2452_), .A2(new_n2405_), .B(new_n376_), .ZN(new_n2453_));
  OAI21_X1   g02261(.A1(new_n2408_), .A2(new_n2453_), .B(\asqrt[60] ), .ZN(new_n2454_));
  AOI21_X1   g02262(.A1(new_n2412_), .A2(new_n2454_), .B(new_n229_), .ZN(new_n2455_));
  NOR3_X1    g02263(.A1(new_n2356_), .A2(\asqrt[61] ), .A3(new_n2358_), .ZN(new_n2456_));
  NAND2_X1   g02264(.A1(\asqrt[46] ), .A2(new_n2456_), .ZN(new_n2457_));
  XOR2_X1    g02265(.A1(new_n2457_), .A2(new_n2455_), .Z(new_n2458_));
  NOR2_X1    g02266(.A1(new_n2458_), .A2(new_n196_), .ZN(new_n2459_));
  INV_X1     g02267(.I(new_n2459_), .ZN(new_n2460_));
  INV_X1     g02268(.I(\a[92] ), .ZN(new_n2461_));
  NOR2_X1    g02269(.A1(\a[90] ), .A2(\a[91] ), .ZN(new_n2462_));
  INV_X1     g02270(.I(new_n2462_), .ZN(new_n2463_));
  NOR3_X1    g02271(.A1(new_n2259_), .A2(new_n2461_), .A3(new_n2463_), .ZN(new_n2464_));
  NAND2_X1   g02272(.A1(new_n2265_), .A2(new_n2464_), .ZN(new_n2465_));
  XOR2_X1    g02273(.A1(new_n2465_), .A2(\a[93] ), .Z(new_n2466_));
  INV_X1     g02274(.I(\a[93] ), .ZN(new_n2467_));
  NOR4_X1    g02275(.A1(new_n2445_), .A2(new_n2467_), .A3(new_n2418_), .A4(new_n2440_), .ZN(new_n2468_));
  NOR2_X1    g02276(.A1(new_n2467_), .A2(\a[92] ), .ZN(new_n2469_));
  OAI21_X1   g02277(.A1(new_n2468_), .A2(new_n2469_), .B(new_n2466_), .ZN(new_n2470_));
  INV_X1     g02278(.I(new_n2466_), .ZN(new_n2471_));
  INV_X1     g02279(.I(new_n2418_), .ZN(new_n2472_));
  NOR3_X1    g02280(.A1(new_n2415_), .A2(new_n2412_), .A3(new_n2433_), .ZN(new_n2473_));
  AOI21_X1   g02281(.A1(new_n2473_), .A2(new_n2455_), .B(new_n2426_), .ZN(new_n2474_));
  AOI21_X1   g02282(.A1(new_n2474_), .A2(new_n2438_), .B(new_n2424_), .ZN(new_n2475_));
  NAND4_X1   g02283(.A1(new_n2362_), .A2(new_n196_), .A3(new_n2425_), .A4(new_n2222_), .ZN(new_n2476_));
  INV_X1     g02284(.I(new_n2444_), .ZN(new_n2477_));
  NOR2_X1    g02285(.A1(new_n2476_), .A2(new_n2477_), .ZN(new_n2478_));
  NAND4_X1   g02286(.A1(new_n2478_), .A2(\a[93] ), .A3(new_n2475_), .A4(new_n2472_), .ZN(new_n2479_));
  NAND3_X1   g02287(.A1(new_n2479_), .A2(\a[92] ), .A3(new_n2471_), .ZN(new_n2480_));
  NAND2_X1   g02288(.A1(new_n2470_), .A2(new_n2480_), .ZN(new_n2481_));
  NOR2_X1    g02289(.A1(new_n2445_), .A2(new_n2440_), .ZN(new_n2482_));
  NOR4_X1    g02290(.A1(new_n2214_), .A2(new_n2208_), .A3(new_n2255_), .A4(new_n2216_), .ZN(new_n2483_));
  NAND2_X1   g02291(.A1(\asqrt[47] ), .A2(\a[92] ), .ZN(new_n2484_));
  XOR2_X1    g02292(.A1(new_n2484_), .A2(new_n2483_), .Z(new_n2485_));
  NOR2_X1    g02293(.A1(new_n2485_), .A2(new_n2463_), .ZN(new_n2486_));
  INV_X1     g02294(.I(new_n2486_), .ZN(new_n2487_));
  NAND3_X1   g02295(.A1(new_n2478_), .A2(new_n2472_), .A3(new_n2475_), .ZN(new_n2488_));
  NOR2_X1    g02296(.A1(new_n2444_), .A2(new_n2472_), .ZN(new_n2489_));
  NAND2_X1   g02297(.A1(new_n2489_), .A2(\asqrt[47] ), .ZN(new_n2490_));
  INV_X1     g02298(.I(new_n2490_), .ZN(new_n2491_));
  NAND3_X1   g02299(.A1(new_n2440_), .A2(new_n2476_), .A3(new_n2491_), .ZN(new_n2492_));
  NAND2_X1   g02300(.A1(new_n2492_), .A2(new_n2224_), .ZN(new_n2493_));
  NAND3_X1   g02301(.A1(new_n2493_), .A2(new_n2225_), .A3(new_n2488_), .ZN(new_n2494_));
  NOR3_X1    g02302(.A1(new_n2475_), .A2(new_n2441_), .A3(new_n2490_), .ZN(new_n2495_));
  OAI21_X1   g02303(.A1(new_n2495_), .A2(\a[94] ), .B(new_n2225_), .ZN(new_n2496_));
  NAND2_X1   g02304(.A1(new_n2496_), .A2(\asqrt[46] ), .ZN(new_n2497_));
  NAND4_X1   g02305(.A1(new_n2497_), .A2(new_n2046_), .A3(new_n2494_), .A4(new_n2487_), .ZN(new_n2498_));
  NAND2_X1   g02306(.A1(new_n2498_), .A2(new_n2481_), .ZN(new_n2499_));
  NAND3_X1   g02307(.A1(new_n2470_), .A2(new_n2480_), .A3(new_n2487_), .ZN(new_n2500_));
  NAND2_X1   g02308(.A1(\asqrt[47] ), .A2(new_n2224_), .ZN(new_n2501_));
  AOI22_X1   g02309(.A1(new_n2501_), .A2(new_n2223_), .B1(new_n2224_), .B2(new_n2229_), .ZN(new_n2502_));
  OAI21_X1   g02310(.A1(new_n2253_), .A2(new_n2224_), .B(new_n2227_), .ZN(new_n2503_));
  NOR2_X1    g02311(.A1(new_n2502_), .A2(new_n2503_), .ZN(new_n2504_));
  NAND3_X1   g02312(.A1(\asqrt[46] ), .A2(new_n2252_), .A3(new_n2504_), .ZN(new_n2505_));
  INV_X1     g02313(.I(new_n2504_), .ZN(new_n2506_));
  OAI21_X1   g02314(.A1(new_n2488_), .A2(new_n2506_), .B(new_n2251_), .ZN(new_n2507_));
  NAND3_X1   g02315(.A1(new_n2505_), .A2(new_n2507_), .A3(new_n1854_), .ZN(new_n2508_));
  AOI21_X1   g02316(.A1(new_n2500_), .A2(\asqrt[48] ), .B(new_n2508_), .ZN(new_n2509_));
  NOR2_X1    g02317(.A1(new_n2499_), .A2(new_n2509_), .ZN(new_n2510_));
  NAND2_X1   g02318(.A1(new_n2500_), .A2(\asqrt[48] ), .ZN(new_n2511_));
  AOI21_X1   g02319(.A1(new_n2499_), .A2(new_n2511_), .B(new_n1854_), .ZN(new_n2512_));
  NOR2_X1    g02320(.A1(new_n2369_), .A2(new_n2368_), .ZN(new_n2513_));
  NOR4_X1    g02321(.A1(new_n2488_), .A2(\asqrt[49] ), .A3(new_n2513_), .A4(new_n2271_), .ZN(new_n2514_));
  AOI21_X1   g02322(.A1(new_n2367_), .A2(new_n2252_), .B(new_n1854_), .ZN(new_n2515_));
  NOR2_X1    g02323(.A1(new_n2514_), .A2(new_n2515_), .ZN(new_n2516_));
  NAND2_X1   g02324(.A1(new_n2516_), .A2(new_n1595_), .ZN(new_n2517_));
  OAI21_X1   g02325(.A1(new_n2512_), .A2(new_n2517_), .B(new_n2510_), .ZN(new_n2518_));
  AOI22_X1   g02326(.A1(new_n2498_), .A2(new_n2481_), .B1(\asqrt[48] ), .B2(new_n2500_), .ZN(new_n2519_));
  OAI22_X1   g02327(.A1(new_n2519_), .A2(new_n1854_), .B1(new_n2499_), .B2(new_n2509_), .ZN(new_n2520_));
  NOR2_X1    g02328(.A1(new_n2282_), .A2(new_n1595_), .ZN(new_n2521_));
  NAND2_X1   g02329(.A1(new_n2277_), .A2(new_n2278_), .ZN(new_n2522_));
  NAND4_X1   g02330(.A1(\asqrt[46] ), .A2(new_n1595_), .A3(new_n2522_), .A4(new_n2282_), .ZN(new_n2523_));
  XOR2_X1    g02331(.A1(new_n2523_), .A2(new_n2521_), .Z(new_n2524_));
  NAND2_X1   g02332(.A1(new_n2524_), .A2(new_n1436_), .ZN(new_n2525_));
  AOI21_X1   g02333(.A1(new_n2520_), .A2(\asqrt[50] ), .B(new_n2525_), .ZN(new_n2526_));
  OAI21_X1   g02334(.A1(new_n2512_), .A2(new_n2510_), .B(\asqrt[50] ), .ZN(new_n2527_));
  AOI21_X1   g02335(.A1(new_n2518_), .A2(new_n2527_), .B(new_n1436_), .ZN(new_n2528_));
  NAND2_X1   g02336(.A1(new_n2292_), .A2(\asqrt[51] ), .ZN(new_n2529_));
  NOR4_X1    g02337(.A1(new_n2488_), .A2(\asqrt[51] ), .A3(new_n2287_), .A4(new_n2292_), .ZN(new_n2530_));
  XOR2_X1    g02338(.A1(new_n2530_), .A2(new_n2529_), .Z(new_n2531_));
  NAND2_X1   g02339(.A1(new_n2531_), .A2(new_n1260_), .ZN(new_n2532_));
  NOR2_X1    g02340(.A1(new_n2528_), .A2(new_n2532_), .ZN(new_n2533_));
  NOR3_X1    g02341(.A1(new_n2533_), .A2(new_n2518_), .A3(new_n2526_), .ZN(new_n2534_));
  INV_X1     g02342(.I(new_n2525_), .ZN(new_n2535_));
  AOI21_X1   g02343(.A1(new_n2527_), .A2(new_n2535_), .B(new_n2518_), .ZN(new_n2536_));
  OAI21_X1   g02344(.A1(new_n2536_), .A2(new_n2528_), .B(\asqrt[52] ), .ZN(new_n2537_));
  NAND2_X1   g02345(.A1(new_n2385_), .A2(\asqrt[52] ), .ZN(new_n2538_));
  NOR4_X1    g02346(.A1(new_n2488_), .A2(\asqrt[52] ), .A3(new_n2295_), .A4(new_n2385_), .ZN(new_n2539_));
  XOR2_X1    g02347(.A1(new_n2539_), .A2(new_n2538_), .Z(new_n2540_));
  NAND2_X1   g02348(.A1(new_n2540_), .A2(new_n1096_), .ZN(new_n2541_));
  INV_X1     g02349(.I(new_n2541_), .ZN(new_n2542_));
  NAND2_X1   g02350(.A1(new_n2537_), .A2(new_n2542_), .ZN(new_n2543_));
  NAND2_X1   g02351(.A1(new_n2543_), .A2(new_n2534_), .ZN(new_n2544_));
  OAI21_X1   g02352(.A1(new_n2528_), .A2(new_n2532_), .B(new_n2536_), .ZN(new_n2545_));
  NAND2_X1   g02353(.A1(new_n2545_), .A2(new_n2537_), .ZN(new_n2546_));
  NAND2_X1   g02354(.A1(new_n2307_), .A2(\asqrt[53] ), .ZN(new_n2547_));
  NOR4_X1    g02355(.A1(new_n2488_), .A2(\asqrt[53] ), .A3(new_n2302_), .A4(new_n2307_), .ZN(new_n2548_));
  XOR2_X1    g02356(.A1(new_n2548_), .A2(new_n2547_), .Z(new_n2549_));
  NAND2_X1   g02357(.A1(new_n2549_), .A2(new_n970_), .ZN(new_n2550_));
  AOI21_X1   g02358(.A1(new_n2546_), .A2(\asqrt[53] ), .B(new_n2550_), .ZN(new_n2551_));
  NOR2_X1    g02359(.A1(new_n2551_), .A2(new_n2544_), .ZN(new_n2552_));
  AOI22_X1   g02360(.A1(new_n2546_), .A2(\asqrt[53] ), .B1(new_n2543_), .B2(new_n2534_), .ZN(new_n2553_));
  NAND2_X1   g02361(.A1(new_n2392_), .A2(\asqrt[54] ), .ZN(new_n2554_));
  NOR4_X1    g02362(.A1(new_n2488_), .A2(\asqrt[54] ), .A3(new_n2310_), .A4(new_n2392_), .ZN(new_n2555_));
  XOR2_X1    g02363(.A1(new_n2555_), .A2(new_n2554_), .Z(new_n2556_));
  NAND2_X1   g02364(.A1(new_n2556_), .A2(new_n825_), .ZN(new_n2557_));
  INV_X1     g02365(.I(new_n2557_), .ZN(new_n2558_));
  OAI21_X1   g02366(.A1(new_n2553_), .A2(new_n970_), .B(new_n2558_), .ZN(new_n2559_));
  NAND2_X1   g02367(.A1(new_n2559_), .A2(new_n2552_), .ZN(new_n2560_));
  OAI22_X1   g02368(.A1(new_n2553_), .A2(new_n970_), .B1(new_n2551_), .B2(new_n2544_), .ZN(new_n2561_));
  NAND2_X1   g02369(.A1(new_n2321_), .A2(\asqrt[55] ), .ZN(new_n2562_));
  NOR4_X1    g02370(.A1(new_n2488_), .A2(\asqrt[55] ), .A3(new_n2316_), .A4(new_n2321_), .ZN(new_n2563_));
  XOR2_X1    g02371(.A1(new_n2563_), .A2(new_n2562_), .Z(new_n2564_));
  NAND2_X1   g02372(.A1(new_n2564_), .A2(new_n724_), .ZN(new_n2565_));
  AOI21_X1   g02373(.A1(new_n2561_), .A2(\asqrt[55] ), .B(new_n2565_), .ZN(new_n2566_));
  NOR2_X1    g02374(.A1(new_n2566_), .A2(new_n2560_), .ZN(new_n2567_));
  AOI22_X1   g02375(.A1(new_n2561_), .A2(\asqrt[55] ), .B1(new_n2559_), .B2(new_n2552_), .ZN(new_n2568_));
  NAND2_X1   g02376(.A1(new_n2399_), .A2(\asqrt[56] ), .ZN(new_n2569_));
  NOR4_X1    g02377(.A1(new_n2488_), .A2(\asqrt[56] ), .A3(new_n2324_), .A4(new_n2399_), .ZN(new_n2570_));
  XOR2_X1    g02378(.A1(new_n2570_), .A2(new_n2569_), .Z(new_n2571_));
  NAND2_X1   g02379(.A1(new_n2571_), .A2(new_n587_), .ZN(new_n2572_));
  INV_X1     g02380(.I(new_n2572_), .ZN(new_n2573_));
  OAI21_X1   g02381(.A1(new_n2568_), .A2(new_n724_), .B(new_n2573_), .ZN(new_n2574_));
  NAND2_X1   g02382(.A1(new_n2574_), .A2(new_n2567_), .ZN(new_n2575_));
  AOI21_X1   g02383(.A1(new_n2545_), .A2(new_n2537_), .B(new_n1096_), .ZN(new_n2576_));
  INV_X1     g02384(.I(new_n2576_), .ZN(new_n2577_));
  AOI21_X1   g02385(.A1(new_n2577_), .A2(new_n2544_), .B(new_n970_), .ZN(new_n2578_));
  OAI21_X1   g02386(.A1(new_n2578_), .A2(new_n2552_), .B(\asqrt[55] ), .ZN(new_n2579_));
  AOI21_X1   g02387(.A1(new_n2560_), .A2(new_n2579_), .B(new_n724_), .ZN(new_n2580_));
  OAI21_X1   g02388(.A1(new_n2567_), .A2(new_n2580_), .B(\asqrt[57] ), .ZN(new_n2581_));
  NOR4_X1    g02389(.A1(new_n2488_), .A2(\asqrt[57] ), .A3(new_n2330_), .A4(new_n2335_), .ZN(new_n2582_));
  XOR2_X1    g02390(.A1(new_n2582_), .A2(new_n2428_), .Z(new_n2583_));
  AND2_X2    g02391(.A1(new_n2583_), .A2(new_n504_), .Z(new_n2584_));
  AOI21_X1   g02392(.A1(new_n2581_), .A2(new_n2584_), .B(new_n2575_), .ZN(new_n2585_));
  OAI22_X1   g02393(.A1(new_n2568_), .A2(new_n724_), .B1(new_n2566_), .B2(new_n2560_), .ZN(new_n2586_));
  AOI22_X1   g02394(.A1(new_n2586_), .A2(\asqrt[57] ), .B1(new_n2574_), .B2(new_n2567_), .ZN(new_n2587_));
  NOR4_X1    g02395(.A1(new_n2488_), .A2(\asqrt[58] ), .A3(new_n2338_), .A4(new_n2406_), .ZN(new_n2588_));
  XOR2_X1    g02396(.A1(new_n2588_), .A2(new_n2452_), .Z(new_n2589_));
  NAND2_X1   g02397(.A1(new_n2589_), .A2(new_n376_), .ZN(new_n2590_));
  INV_X1     g02398(.I(new_n2590_), .ZN(new_n2591_));
  OAI21_X1   g02399(.A1(new_n2587_), .A2(new_n504_), .B(new_n2591_), .ZN(new_n2592_));
  NAND2_X1   g02400(.A1(new_n2592_), .A2(new_n2585_), .ZN(new_n2593_));
  AOI21_X1   g02401(.A1(new_n2575_), .A2(new_n2581_), .B(new_n504_), .ZN(new_n2594_));
  OAI21_X1   g02402(.A1(new_n2585_), .A2(new_n2594_), .B(\asqrt[59] ), .ZN(new_n2595_));
  NOR4_X1    g02403(.A1(new_n2488_), .A2(\asqrt[59] ), .A3(new_n2344_), .A4(new_n2349_), .ZN(new_n2596_));
  XOR2_X1    g02404(.A1(new_n2596_), .A2(new_n2430_), .Z(new_n2597_));
  AND2_X2    g02405(.A1(new_n2597_), .A2(new_n275_), .Z(new_n2598_));
  AOI21_X1   g02406(.A1(new_n2595_), .A2(new_n2598_), .B(new_n2593_), .ZN(new_n2599_));
  INV_X1     g02407(.I(new_n2517_), .ZN(new_n2600_));
  OAI21_X1   g02408(.A1(new_n2519_), .A2(new_n1854_), .B(new_n2600_), .ZN(new_n2601_));
  AOI22_X1   g02409(.A1(new_n2520_), .A2(\asqrt[50] ), .B1(new_n2601_), .B2(new_n2510_), .ZN(new_n2602_));
  OAI22_X1   g02410(.A1(new_n2602_), .A2(new_n1436_), .B1(new_n2526_), .B2(new_n2518_), .ZN(new_n2603_));
  AOI21_X1   g02411(.A1(new_n2603_), .A2(\asqrt[52] ), .B(new_n2541_), .ZN(new_n2604_));
  NOR2_X1    g02412(.A1(new_n2604_), .A2(new_n2545_), .ZN(new_n2605_));
  INV_X1     g02413(.I(new_n2532_), .ZN(new_n2606_));
  OAI21_X1   g02414(.A1(new_n2602_), .A2(new_n1436_), .B(new_n2606_), .ZN(new_n2607_));
  AOI22_X1   g02415(.A1(new_n2603_), .A2(\asqrt[52] ), .B1(new_n2607_), .B2(new_n2536_), .ZN(new_n2608_));
  INV_X1     g02416(.I(new_n2550_), .ZN(new_n2609_));
  OAI21_X1   g02417(.A1(new_n2608_), .A2(new_n1096_), .B(new_n2609_), .ZN(new_n2610_));
  NAND2_X1   g02418(.A1(new_n2610_), .A2(new_n2605_), .ZN(new_n2611_));
  OAI22_X1   g02419(.A1(new_n2608_), .A2(new_n1096_), .B1(new_n2604_), .B2(new_n2545_), .ZN(new_n2612_));
  AOI21_X1   g02420(.A1(new_n2612_), .A2(\asqrt[54] ), .B(new_n2557_), .ZN(new_n2613_));
  NOR2_X1    g02421(.A1(new_n2613_), .A2(new_n2611_), .ZN(new_n2614_));
  AOI22_X1   g02422(.A1(new_n2612_), .A2(\asqrt[54] ), .B1(new_n2610_), .B2(new_n2605_), .ZN(new_n2615_));
  INV_X1     g02423(.I(new_n2565_), .ZN(new_n2616_));
  OAI21_X1   g02424(.A1(new_n2615_), .A2(new_n825_), .B(new_n2616_), .ZN(new_n2617_));
  NAND2_X1   g02425(.A1(new_n2617_), .A2(new_n2614_), .ZN(new_n2618_));
  OAI22_X1   g02426(.A1(new_n2615_), .A2(new_n825_), .B1(new_n2613_), .B2(new_n2611_), .ZN(new_n2619_));
  AOI21_X1   g02427(.A1(new_n2619_), .A2(\asqrt[56] ), .B(new_n2572_), .ZN(new_n2620_));
  NOR2_X1    g02428(.A1(new_n2620_), .A2(new_n2618_), .ZN(new_n2621_));
  AOI22_X1   g02429(.A1(new_n2619_), .A2(\asqrt[56] ), .B1(new_n2617_), .B2(new_n2614_), .ZN(new_n2622_));
  OAI21_X1   g02430(.A1(new_n2622_), .A2(new_n587_), .B(new_n2584_), .ZN(new_n2623_));
  NAND2_X1   g02431(.A1(new_n2623_), .A2(new_n2621_), .ZN(new_n2624_));
  OAI21_X1   g02432(.A1(new_n2605_), .A2(new_n2576_), .B(\asqrt[54] ), .ZN(new_n2625_));
  AOI21_X1   g02433(.A1(new_n2611_), .A2(new_n2625_), .B(new_n825_), .ZN(new_n2626_));
  OAI21_X1   g02434(.A1(new_n2614_), .A2(new_n2626_), .B(\asqrt[56] ), .ZN(new_n2627_));
  AOI21_X1   g02435(.A1(new_n2618_), .A2(new_n2627_), .B(new_n587_), .ZN(new_n2628_));
  OAI21_X1   g02436(.A1(new_n2621_), .A2(new_n2628_), .B(\asqrt[58] ), .ZN(new_n2629_));
  NAND2_X1   g02437(.A1(new_n2624_), .A2(new_n2629_), .ZN(new_n2630_));
  AOI22_X1   g02438(.A1(new_n2630_), .A2(\asqrt[59] ), .B1(new_n2592_), .B2(new_n2585_), .ZN(new_n2631_));
  NOR3_X1    g02439(.A1(new_n2413_), .A2(\asqrt[60] ), .A3(new_n2351_), .ZN(new_n2632_));
  NAND2_X1   g02440(.A1(\asqrt[46] ), .A2(new_n2632_), .ZN(new_n2633_));
  XOR2_X1    g02441(.A1(new_n2633_), .A2(new_n2431_), .Z(new_n2634_));
  NAND2_X1   g02442(.A1(new_n2634_), .A2(new_n229_), .ZN(new_n2635_));
  INV_X1     g02443(.I(new_n2635_), .ZN(new_n2636_));
  OAI21_X1   g02444(.A1(new_n2631_), .A2(new_n275_), .B(new_n2636_), .ZN(new_n2637_));
  OAI22_X1   g02445(.A1(new_n2622_), .A2(new_n587_), .B1(new_n2620_), .B2(new_n2618_), .ZN(new_n2638_));
  AOI21_X1   g02446(.A1(new_n2638_), .A2(\asqrt[58] ), .B(new_n2590_), .ZN(new_n2639_));
  NOR2_X1    g02447(.A1(new_n2639_), .A2(new_n2624_), .ZN(new_n2640_));
  AOI22_X1   g02448(.A1(new_n2638_), .A2(\asqrt[58] ), .B1(new_n2623_), .B2(new_n2621_), .ZN(new_n2641_));
  OAI21_X1   g02449(.A1(new_n2641_), .A2(new_n376_), .B(new_n2598_), .ZN(new_n2642_));
  NAND2_X1   g02450(.A1(new_n2642_), .A2(new_n2640_), .ZN(new_n2643_));
  AOI21_X1   g02451(.A1(new_n2624_), .A2(new_n2629_), .B(new_n376_), .ZN(new_n2644_));
  OAI21_X1   g02452(.A1(new_n2640_), .A2(new_n2644_), .B(\asqrt[60] ), .ZN(new_n2645_));
  AOI21_X1   g02453(.A1(new_n2643_), .A2(new_n2645_), .B(new_n229_), .ZN(new_n2646_));
  INV_X1     g02454(.I(new_n2458_), .ZN(new_n2647_));
  NOR2_X1    g02455(.A1(new_n2647_), .A2(\asqrt[62] ), .ZN(new_n2648_));
  INV_X1     g02456(.I(new_n2648_), .ZN(new_n2649_));
  NAND4_X1   g02457(.A1(new_n2646_), .A2(new_n2599_), .A3(new_n2637_), .A4(new_n2649_), .ZN(new_n2650_));
  NAND2_X1   g02458(.A1(new_n2476_), .A2(new_n2424_), .ZN(new_n2651_));
  OAI21_X1   g02459(.A1(\asqrt[46] ), .A2(new_n2651_), .B(new_n2436_), .ZN(new_n2652_));
  NAND2_X1   g02460(.A1(new_n2652_), .A2(new_n231_), .ZN(new_n2653_));
  INV_X1     g02461(.I(new_n2653_), .ZN(new_n2654_));
  NAND3_X1   g02462(.A1(new_n2650_), .A2(new_n2460_), .A3(new_n2654_), .ZN(new_n2655_));
  OAI22_X1   g02463(.A1(new_n2641_), .A2(new_n376_), .B1(new_n2639_), .B2(new_n2624_), .ZN(new_n2656_));
  AOI21_X1   g02464(.A1(new_n2656_), .A2(\asqrt[60] ), .B(new_n2635_), .ZN(new_n2657_));
  AOI22_X1   g02465(.A1(new_n2656_), .A2(\asqrt[60] ), .B1(new_n2642_), .B2(new_n2640_), .ZN(new_n2658_));
  OAI22_X1   g02466(.A1(new_n2658_), .A2(new_n229_), .B1(new_n2657_), .B2(new_n2643_), .ZN(new_n2659_));
  NOR4_X1    g02467(.A1(new_n2659_), .A2(\asqrt[62] ), .A3(new_n2450_), .A4(new_n2458_), .ZN(new_n2660_));
  AOI21_X1   g02468(.A1(new_n2451_), .A2(new_n2655_), .B(new_n2660_), .ZN(new_n2661_));
  INV_X1     g02469(.I(\a[88] ), .ZN(new_n2662_));
  OAI21_X1   g02470(.A1(new_n2425_), .A2(new_n2436_), .B(\asqrt[46] ), .ZN(new_n2663_));
  XOR2_X1    g02471(.A1(new_n2436_), .A2(\asqrt[63] ), .Z(new_n2664_));
  NAND2_X1   g02472(.A1(new_n2663_), .A2(new_n2664_), .ZN(new_n2665_));
  INV_X1     g02473(.I(new_n2665_), .ZN(new_n2666_));
  NAND3_X1   g02474(.A1(new_n2482_), .A2(new_n2418_), .A3(new_n2425_), .ZN(new_n2667_));
  INV_X1     g02475(.I(new_n2667_), .ZN(new_n2668_));
  NOR2_X1    g02476(.A1(new_n2666_), .A2(new_n2668_), .ZN(new_n2669_));
  NOR2_X1    g02477(.A1(\a[86] ), .A2(\a[87] ), .ZN(new_n2670_));
  INV_X1     g02478(.I(new_n2670_), .ZN(new_n2671_));
  NOR3_X1    g02479(.A1(new_n2669_), .A2(new_n2662_), .A3(new_n2671_), .ZN(new_n2672_));
  NAND2_X1   g02480(.A1(new_n2661_), .A2(new_n2672_), .ZN(new_n2673_));
  XOR2_X1    g02481(.A1(new_n2673_), .A2(\a[89] ), .Z(new_n2674_));
  INV_X1     g02482(.I(\a[89] ), .ZN(new_n2675_));
  NAND2_X1   g02483(.A1(new_n2637_), .A2(new_n2599_), .ZN(new_n2676_));
  NAND2_X1   g02484(.A1(new_n2646_), .A2(new_n2649_), .ZN(new_n2677_));
  OAI21_X1   g02485(.A1(new_n2677_), .A2(new_n2676_), .B(new_n2460_), .ZN(new_n2678_));
  OAI21_X1   g02486(.A1(new_n2678_), .A2(new_n2653_), .B(new_n2451_), .ZN(new_n2679_));
  NAND2_X1   g02487(.A1(new_n2660_), .A2(new_n2666_), .ZN(new_n2680_));
  NOR2_X1    g02488(.A1(new_n2680_), .A2(new_n2679_), .ZN(new_n2681_));
  NAND3_X1   g02489(.A1(new_n2681_), .A2(new_n2451_), .A3(new_n2667_), .ZN(new_n2682_));
  NAND2_X1   g02490(.A1(new_n2643_), .A2(new_n2645_), .ZN(new_n2683_));
  AOI22_X1   g02491(.A1(new_n2683_), .A2(\asqrt[61] ), .B1(new_n2637_), .B2(new_n2599_), .ZN(new_n2684_));
  NOR2_X1    g02492(.A1(new_n2684_), .A2(new_n196_), .ZN(new_n2685_));
  AOI21_X1   g02493(.A1(new_n2593_), .A2(new_n2595_), .B(new_n275_), .ZN(new_n2686_));
  OAI21_X1   g02494(.A1(new_n2599_), .A2(new_n2686_), .B(\asqrt[61] ), .ZN(new_n2687_));
  NAND4_X1   g02495(.A1(new_n2676_), .A2(new_n196_), .A3(new_n2687_), .A4(new_n2647_), .ZN(new_n2688_));
  INV_X1     g02496(.I(new_n2688_), .ZN(new_n2689_));
  NOR3_X1    g02497(.A1(new_n2680_), .A2(new_n2679_), .A3(new_n2667_), .ZN(\asqrt[45] ));
  NAND3_X1   g02498(.A1(\asqrt[45] ), .A2(new_n2685_), .A3(new_n2689_), .ZN(new_n2691_));
  OAI21_X1   g02499(.A1(new_n2659_), .A2(\asqrt[62] ), .B(new_n2458_), .ZN(new_n2692_));
  OAI21_X1   g02500(.A1(\asqrt[45] ), .A2(new_n2692_), .B(new_n2685_), .ZN(new_n2693_));
  NAND2_X1   g02501(.A1(new_n2693_), .A2(new_n2691_), .ZN(new_n2694_));
  INV_X1     g02502(.I(new_n2694_), .ZN(new_n2695_));
  INV_X1     g02503(.I(new_n2634_), .ZN(new_n2696_));
  NAND4_X1   g02504(.A1(\asqrt[45] ), .A2(new_n229_), .A3(new_n2696_), .A4(new_n2658_), .ZN(new_n2697_));
  XOR2_X1    g02505(.A1(new_n2697_), .A2(new_n2646_), .Z(new_n2698_));
  NOR2_X1    g02506(.A1(new_n2698_), .A2(new_n196_), .ZN(new_n2699_));
  INV_X1     g02507(.I(new_n2699_), .ZN(new_n2700_));
  INV_X1     g02508(.I(\a[91] ), .ZN(new_n2701_));
  INV_X1     g02509(.I(\a[90] ), .ZN(new_n2702_));
  NOR2_X1    g02510(.A1(new_n2475_), .A2(new_n2441_), .ZN(new_n2703_));
  INV_X1     g02511(.I(new_n2703_), .ZN(new_n2704_));
  NOR2_X1    g02512(.A1(\a[88] ), .A2(\a[89] ), .ZN(new_n2705_));
  INV_X1     g02513(.I(new_n2705_), .ZN(new_n2706_));
  NOR4_X1    g02514(.A1(new_n2704_), .A2(new_n2702_), .A3(new_n2489_), .A4(new_n2706_), .ZN(new_n2707_));
  XOR2_X1    g02515(.A1(new_n2707_), .A2(new_n2701_), .Z(new_n2708_));
  NOR4_X1    g02516(.A1(new_n2680_), .A2(new_n2679_), .A3(new_n2701_), .A4(new_n2667_), .ZN(new_n2709_));
  NOR2_X1    g02517(.A1(new_n2701_), .A2(\a[90] ), .ZN(new_n2710_));
  OAI21_X1   g02518(.A1(new_n2709_), .A2(new_n2710_), .B(new_n2708_), .ZN(new_n2711_));
  INV_X1     g02519(.I(new_n2708_), .ZN(new_n2712_));
  NOR2_X1    g02520(.A1(new_n2657_), .A2(new_n2643_), .ZN(new_n2713_));
  NOR3_X1    g02521(.A1(new_n2658_), .A2(new_n229_), .A3(new_n2648_), .ZN(new_n2714_));
  AOI21_X1   g02522(.A1(new_n2714_), .A2(new_n2713_), .B(new_n2459_), .ZN(new_n2715_));
  AOI21_X1   g02523(.A1(new_n2715_), .A2(new_n2654_), .B(new_n2450_), .ZN(new_n2716_));
  AOI21_X1   g02524(.A1(new_n2659_), .A2(\asqrt[62] ), .B(new_n2451_), .ZN(new_n2717_));
  NOR3_X1    g02525(.A1(new_n2717_), .A2(new_n2688_), .A3(new_n2665_), .ZN(new_n2718_));
  NAND4_X1   g02526(.A1(new_n2718_), .A2(\a[91] ), .A3(new_n2716_), .A4(new_n2668_), .ZN(new_n2719_));
  NAND3_X1   g02527(.A1(new_n2719_), .A2(\a[90] ), .A3(new_n2712_), .ZN(new_n2720_));
  NAND2_X1   g02528(.A1(new_n2711_), .A2(new_n2720_), .ZN(new_n2721_));
  NOR2_X1    g02529(.A1(new_n2436_), .A2(new_n2439_), .ZN(new_n2722_));
  NOR4_X1    g02530(.A1(new_n2445_), .A2(new_n2418_), .A3(new_n2424_), .A4(new_n2722_), .ZN(new_n2723_));
  NOR2_X1    g02531(.A1(new_n2488_), .A2(new_n2702_), .ZN(new_n2724_));
  XNOR2_X1   g02532(.A1(new_n2724_), .A2(new_n2723_), .ZN(new_n2725_));
  NOR2_X1    g02533(.A1(new_n2725_), .A2(new_n2706_), .ZN(new_n2726_));
  INV_X1     g02534(.I(new_n2726_), .ZN(new_n2727_));
  NAND3_X1   g02535(.A1(new_n2718_), .A2(new_n2716_), .A3(new_n2668_), .ZN(new_n2728_));
  NOR4_X1    g02536(.A1(new_n2687_), .A2(new_n2643_), .A3(new_n2657_), .A4(new_n2648_), .ZN(new_n2729_));
  NOR3_X1    g02537(.A1(new_n2729_), .A2(new_n2459_), .A3(new_n2653_), .ZN(new_n2730_));
  NAND4_X1   g02538(.A1(new_n2684_), .A2(new_n196_), .A3(new_n2451_), .A4(new_n2647_), .ZN(new_n2731_));
  OAI21_X1   g02539(.A1(new_n2730_), .A2(new_n2450_), .B(new_n2731_), .ZN(new_n2732_));
  NAND2_X1   g02540(.A1(new_n2669_), .A2(\asqrt[46] ), .ZN(new_n2733_));
  OAI21_X1   g02541(.A1(new_n2732_), .A2(new_n2733_), .B(new_n2461_), .ZN(new_n2734_));
  NAND3_X1   g02542(.A1(new_n2734_), .A2(new_n2462_), .A3(new_n2728_), .ZN(new_n2735_));
  INV_X1     g02543(.I(new_n2733_), .ZN(new_n2736_));
  AOI21_X1   g02544(.A1(new_n2661_), .A2(new_n2736_), .B(\a[92] ), .ZN(new_n2737_));
  OAI21_X1   g02545(.A1(new_n2737_), .A2(new_n2463_), .B(\asqrt[45] ), .ZN(new_n2738_));
  NAND4_X1   g02546(.A1(new_n2735_), .A2(new_n2738_), .A3(new_n2253_), .A4(new_n2727_), .ZN(new_n2739_));
  NAND2_X1   g02547(.A1(new_n2739_), .A2(new_n2721_), .ZN(new_n2740_));
  NAND3_X1   g02548(.A1(new_n2711_), .A2(new_n2720_), .A3(new_n2727_), .ZN(new_n2741_));
  AOI21_X1   g02549(.A1(\asqrt[46] ), .A2(new_n2461_), .B(\a[93] ), .ZN(new_n2742_));
  NOR2_X1    g02550(.A1(new_n2479_), .A2(\a[92] ), .ZN(new_n2743_));
  AOI21_X1   g02551(.A1(\asqrt[46] ), .A2(\a[92] ), .B(new_n2465_), .ZN(new_n2744_));
  OAI21_X1   g02552(.A1(new_n2742_), .A2(new_n2743_), .B(new_n2744_), .ZN(new_n2745_));
  INV_X1     g02553(.I(new_n2745_), .ZN(new_n2746_));
  NAND3_X1   g02554(.A1(\asqrt[45] ), .A2(new_n2487_), .A3(new_n2746_), .ZN(new_n2747_));
  OAI21_X1   g02555(.A1(new_n2728_), .A2(new_n2745_), .B(new_n2486_), .ZN(new_n2748_));
  NAND3_X1   g02556(.A1(new_n2747_), .A2(new_n2748_), .A3(new_n2046_), .ZN(new_n2749_));
  AOI21_X1   g02557(.A1(new_n2741_), .A2(\asqrt[47] ), .B(new_n2749_), .ZN(new_n2750_));
  NOR2_X1    g02558(.A1(new_n2740_), .A2(new_n2750_), .ZN(new_n2751_));
  AOI22_X1   g02559(.A1(new_n2739_), .A2(new_n2721_), .B1(\asqrt[47] ), .B2(new_n2741_), .ZN(new_n2752_));
  INV_X1     g02560(.I(new_n2469_), .ZN(new_n2753_));
  AOI21_X1   g02561(.A1(new_n2479_), .A2(new_n2753_), .B(new_n2471_), .ZN(new_n2754_));
  INV_X1     g02562(.I(new_n2480_), .ZN(new_n2755_));
  NOR3_X1    g02563(.A1(new_n2755_), .A2(new_n2754_), .A3(new_n2486_), .ZN(new_n2756_));
  AOI21_X1   g02564(.A1(new_n2497_), .A2(new_n2494_), .B(\asqrt[48] ), .ZN(new_n2757_));
  AND4_X2    g02565(.A1(new_n2756_), .A2(\asqrt[45] ), .A3(new_n2511_), .A4(new_n2757_), .Z(new_n2758_));
  NOR2_X1    g02566(.A1(new_n2756_), .A2(new_n2046_), .ZN(new_n2759_));
  NOR3_X1    g02567(.A1(new_n2758_), .A2(\asqrt[49] ), .A3(new_n2759_), .ZN(new_n2760_));
  OAI21_X1   g02568(.A1(new_n2752_), .A2(new_n2046_), .B(new_n2760_), .ZN(new_n2761_));
  NAND2_X1   g02569(.A1(new_n2761_), .A2(new_n2751_), .ZN(new_n2762_));
  OAI22_X1   g02570(.A1(new_n2752_), .A2(new_n2046_), .B1(new_n2740_), .B2(new_n2750_), .ZN(new_n2763_));
  NAND2_X1   g02571(.A1(new_n2505_), .A2(new_n2507_), .ZN(new_n2764_));
  NAND4_X1   g02572(.A1(\asqrt[45] ), .A2(new_n1854_), .A3(new_n2764_), .A4(new_n2519_), .ZN(new_n2765_));
  XOR2_X1    g02573(.A1(new_n2765_), .A2(new_n2512_), .Z(new_n2766_));
  NAND2_X1   g02574(.A1(new_n2766_), .A2(new_n1595_), .ZN(new_n2767_));
  AOI21_X1   g02575(.A1(new_n2763_), .A2(\asqrt[49] ), .B(new_n2767_), .ZN(new_n2768_));
  NOR2_X1    g02576(.A1(new_n2768_), .A2(new_n2762_), .ZN(new_n2769_));
  AOI22_X1   g02577(.A1(new_n2763_), .A2(\asqrt[49] ), .B1(new_n2761_), .B2(new_n2751_), .ZN(new_n2770_));
  NOR4_X1    g02578(.A1(new_n2728_), .A2(\asqrt[50] ), .A3(new_n2516_), .A4(new_n2520_), .ZN(new_n2771_));
  XOR2_X1    g02579(.A1(new_n2771_), .A2(new_n2527_), .Z(new_n2772_));
  NAND2_X1   g02580(.A1(new_n2772_), .A2(new_n1436_), .ZN(new_n2773_));
  INV_X1     g02581(.I(new_n2773_), .ZN(new_n2774_));
  OAI21_X1   g02582(.A1(new_n2770_), .A2(new_n1595_), .B(new_n2774_), .ZN(new_n2775_));
  NAND2_X1   g02583(.A1(new_n2775_), .A2(new_n2769_), .ZN(new_n2776_));
  OAI22_X1   g02584(.A1(new_n2770_), .A2(new_n1595_), .B1(new_n2768_), .B2(new_n2762_), .ZN(new_n2777_));
  NOR2_X1    g02585(.A1(new_n2524_), .A2(\asqrt[51] ), .ZN(new_n2778_));
  NAND3_X1   g02586(.A1(\asqrt[45] ), .A2(new_n2602_), .A3(new_n2778_), .ZN(new_n2779_));
  XOR2_X1    g02587(.A1(new_n2779_), .A2(new_n2528_), .Z(new_n2780_));
  NAND2_X1   g02588(.A1(new_n2780_), .A2(new_n1260_), .ZN(new_n2781_));
  AOI21_X1   g02589(.A1(new_n2777_), .A2(\asqrt[51] ), .B(new_n2781_), .ZN(new_n2782_));
  NOR2_X1    g02590(.A1(new_n2782_), .A2(new_n2776_), .ZN(new_n2783_));
  AOI22_X1   g02591(.A1(new_n2777_), .A2(\asqrt[51] ), .B1(new_n2775_), .B2(new_n2769_), .ZN(new_n2784_));
  NOR4_X1    g02592(.A1(new_n2728_), .A2(\asqrt[52] ), .A3(new_n2531_), .A4(new_n2603_), .ZN(new_n2785_));
  XOR2_X1    g02593(.A1(new_n2785_), .A2(new_n2537_), .Z(new_n2786_));
  NAND2_X1   g02594(.A1(new_n2786_), .A2(new_n1096_), .ZN(new_n2787_));
  INV_X1     g02595(.I(new_n2787_), .ZN(new_n2788_));
  OAI21_X1   g02596(.A1(new_n2784_), .A2(new_n1260_), .B(new_n2788_), .ZN(new_n2789_));
  NAND2_X1   g02597(.A1(new_n2789_), .A2(new_n2783_), .ZN(new_n2790_));
  OAI22_X1   g02598(.A1(new_n2784_), .A2(new_n1260_), .B1(new_n2782_), .B2(new_n2776_), .ZN(new_n2791_));
  NOR4_X1    g02599(.A1(new_n2728_), .A2(\asqrt[53] ), .A3(new_n2540_), .A4(new_n2546_), .ZN(new_n2792_));
  XOR2_X1    g02600(.A1(new_n2792_), .A2(new_n2577_), .Z(new_n2793_));
  NAND2_X1   g02601(.A1(new_n2793_), .A2(new_n970_), .ZN(new_n2794_));
  AOI21_X1   g02602(.A1(new_n2791_), .A2(\asqrt[53] ), .B(new_n2794_), .ZN(new_n2795_));
  NOR2_X1    g02603(.A1(new_n2795_), .A2(new_n2790_), .ZN(new_n2796_));
  AOI22_X1   g02604(.A1(new_n2791_), .A2(\asqrt[53] ), .B1(new_n2789_), .B2(new_n2783_), .ZN(new_n2797_));
  NOR4_X1    g02605(.A1(new_n2728_), .A2(\asqrt[54] ), .A3(new_n2549_), .A4(new_n2612_), .ZN(new_n2798_));
  XOR2_X1    g02606(.A1(new_n2798_), .A2(new_n2625_), .Z(new_n2799_));
  NAND2_X1   g02607(.A1(new_n2799_), .A2(new_n825_), .ZN(new_n2800_));
  INV_X1     g02608(.I(new_n2800_), .ZN(new_n2801_));
  OAI21_X1   g02609(.A1(new_n2797_), .A2(new_n970_), .B(new_n2801_), .ZN(new_n2802_));
  NAND2_X1   g02610(.A1(new_n2802_), .A2(new_n2796_), .ZN(new_n2803_));
  OAI22_X1   g02611(.A1(new_n2797_), .A2(new_n970_), .B1(new_n2795_), .B2(new_n2790_), .ZN(new_n2804_));
  NOR4_X1    g02612(.A1(new_n2728_), .A2(\asqrt[55] ), .A3(new_n2556_), .A4(new_n2561_), .ZN(new_n2805_));
  XOR2_X1    g02613(.A1(new_n2805_), .A2(new_n2579_), .Z(new_n2806_));
  NAND2_X1   g02614(.A1(new_n2806_), .A2(new_n724_), .ZN(new_n2807_));
  AOI21_X1   g02615(.A1(new_n2804_), .A2(\asqrt[55] ), .B(new_n2807_), .ZN(new_n2808_));
  NOR2_X1    g02616(.A1(new_n2808_), .A2(new_n2803_), .ZN(new_n2809_));
  AOI22_X1   g02617(.A1(new_n2804_), .A2(\asqrt[55] ), .B1(new_n2802_), .B2(new_n2796_), .ZN(new_n2810_));
  NOR4_X1    g02618(.A1(new_n2728_), .A2(\asqrt[56] ), .A3(new_n2564_), .A4(new_n2619_), .ZN(new_n2811_));
  XOR2_X1    g02619(.A1(new_n2811_), .A2(new_n2627_), .Z(new_n2812_));
  NAND2_X1   g02620(.A1(new_n2812_), .A2(new_n587_), .ZN(new_n2813_));
  INV_X1     g02621(.I(new_n2813_), .ZN(new_n2814_));
  OAI21_X1   g02622(.A1(new_n2810_), .A2(new_n724_), .B(new_n2814_), .ZN(new_n2815_));
  NAND2_X1   g02623(.A1(new_n2815_), .A2(new_n2809_), .ZN(new_n2816_));
  OAI22_X1   g02624(.A1(new_n2810_), .A2(new_n724_), .B1(new_n2808_), .B2(new_n2803_), .ZN(new_n2817_));
  NOR4_X1    g02625(.A1(new_n2728_), .A2(\asqrt[57] ), .A3(new_n2571_), .A4(new_n2586_), .ZN(new_n2818_));
  XOR2_X1    g02626(.A1(new_n2818_), .A2(new_n2581_), .Z(new_n2819_));
  NAND2_X1   g02627(.A1(new_n2819_), .A2(new_n504_), .ZN(new_n2820_));
  AOI21_X1   g02628(.A1(new_n2817_), .A2(\asqrt[57] ), .B(new_n2820_), .ZN(new_n2821_));
  NOR2_X1    g02629(.A1(new_n2821_), .A2(new_n2816_), .ZN(new_n2822_));
  AOI22_X1   g02630(.A1(new_n2817_), .A2(\asqrt[57] ), .B1(new_n2815_), .B2(new_n2809_), .ZN(new_n2823_));
  NOR4_X1    g02631(.A1(new_n2728_), .A2(\asqrt[58] ), .A3(new_n2583_), .A4(new_n2638_), .ZN(new_n2824_));
  XOR2_X1    g02632(.A1(new_n2824_), .A2(new_n2629_), .Z(new_n2825_));
  NAND2_X1   g02633(.A1(new_n2825_), .A2(new_n376_), .ZN(new_n2826_));
  INV_X1     g02634(.I(new_n2826_), .ZN(new_n2827_));
  OAI21_X1   g02635(.A1(new_n2823_), .A2(new_n504_), .B(new_n2827_), .ZN(new_n2828_));
  NAND2_X1   g02636(.A1(new_n2828_), .A2(new_n2822_), .ZN(new_n2829_));
  OAI22_X1   g02637(.A1(new_n2823_), .A2(new_n504_), .B1(new_n2821_), .B2(new_n2816_), .ZN(new_n2830_));
  NOR4_X1    g02638(.A1(new_n2728_), .A2(\asqrt[59] ), .A3(new_n2589_), .A4(new_n2630_), .ZN(new_n2831_));
  XOR2_X1    g02639(.A1(new_n2831_), .A2(new_n2595_), .Z(new_n2832_));
  NAND2_X1   g02640(.A1(new_n2832_), .A2(new_n275_), .ZN(new_n2833_));
  AOI21_X1   g02641(.A1(new_n2830_), .A2(\asqrt[59] ), .B(new_n2833_), .ZN(new_n2834_));
  NOR2_X1    g02642(.A1(new_n2834_), .A2(new_n2829_), .ZN(new_n2835_));
  AOI22_X1   g02643(.A1(new_n2830_), .A2(\asqrt[59] ), .B1(new_n2828_), .B2(new_n2822_), .ZN(new_n2836_));
  NOR4_X1    g02644(.A1(new_n2728_), .A2(\asqrt[60] ), .A3(new_n2597_), .A4(new_n2656_), .ZN(new_n2837_));
  XOR2_X1    g02645(.A1(new_n2837_), .A2(new_n2645_), .Z(new_n2838_));
  NAND2_X1   g02646(.A1(new_n2838_), .A2(new_n229_), .ZN(new_n2839_));
  INV_X1     g02647(.I(new_n2839_), .ZN(new_n2840_));
  OAI21_X1   g02648(.A1(new_n2836_), .A2(new_n275_), .B(new_n2840_), .ZN(new_n2841_));
  NAND2_X1   g02649(.A1(new_n2841_), .A2(new_n2835_), .ZN(new_n2842_));
  OAI22_X1   g02650(.A1(new_n2836_), .A2(new_n275_), .B1(new_n2834_), .B2(new_n2829_), .ZN(new_n2843_));
  INV_X1     g02651(.I(new_n2698_), .ZN(new_n2844_));
  NOR2_X1    g02652(.A1(new_n2844_), .A2(\asqrt[62] ), .ZN(new_n2845_));
  INV_X1     g02653(.I(new_n2845_), .ZN(new_n2846_));
  NAND3_X1   g02654(.A1(new_n2843_), .A2(\asqrt[61] ), .A3(new_n2846_), .ZN(new_n2847_));
  OAI21_X1   g02655(.A1(new_n2847_), .A2(new_n2842_), .B(new_n2700_), .ZN(new_n2848_));
  NAND3_X1   g02656(.A1(new_n2728_), .A2(new_n2450_), .A3(new_n2731_), .ZN(new_n2849_));
  AOI21_X1   g02657(.A1(new_n2849_), .A2(new_n2678_), .B(\asqrt[63] ), .ZN(new_n2850_));
  INV_X1     g02658(.I(new_n2850_), .ZN(new_n2851_));
  OAI21_X1   g02659(.A1(new_n2848_), .A2(new_n2851_), .B(new_n2695_), .ZN(new_n2852_));
  INV_X1     g02660(.I(new_n2710_), .ZN(new_n2853_));
  AOI21_X1   g02661(.A1(new_n2719_), .A2(new_n2853_), .B(new_n2712_), .ZN(new_n2854_));
  NOR3_X1    g02662(.A1(new_n2709_), .A2(new_n2702_), .A3(new_n2708_), .ZN(new_n2855_));
  NOR2_X1    g02663(.A1(new_n2855_), .A2(new_n2854_), .ZN(new_n2856_));
  NOR3_X1    g02664(.A1(new_n2737_), .A2(new_n2463_), .A3(\asqrt[45] ), .ZN(new_n2857_));
  AOI21_X1   g02665(.A1(new_n2734_), .A2(new_n2462_), .B(new_n2728_), .ZN(new_n2858_));
  NOR4_X1    g02666(.A1(new_n2858_), .A2(new_n2857_), .A3(\asqrt[47] ), .A4(new_n2726_), .ZN(new_n2859_));
  NOR2_X1    g02667(.A1(new_n2859_), .A2(new_n2856_), .ZN(new_n2860_));
  NOR3_X1    g02668(.A1(new_n2855_), .A2(new_n2854_), .A3(new_n2726_), .ZN(new_n2861_));
  NOR3_X1    g02669(.A1(new_n2728_), .A2(new_n2486_), .A3(new_n2745_), .ZN(new_n2862_));
  AOI21_X1   g02670(.A1(\asqrt[45] ), .A2(new_n2746_), .B(new_n2487_), .ZN(new_n2863_));
  NOR3_X1    g02671(.A1(new_n2863_), .A2(new_n2862_), .A3(\asqrt[48] ), .ZN(new_n2864_));
  OAI21_X1   g02672(.A1(new_n2861_), .A2(new_n2253_), .B(new_n2864_), .ZN(new_n2865_));
  NAND2_X1   g02673(.A1(new_n2860_), .A2(new_n2865_), .ZN(new_n2866_));
  OAI22_X1   g02674(.A1(new_n2859_), .A2(new_n2856_), .B1(new_n2253_), .B2(new_n2861_), .ZN(new_n2867_));
  INV_X1     g02675(.I(new_n2760_), .ZN(new_n2868_));
  AOI21_X1   g02676(.A1(new_n2867_), .A2(\asqrt[48] ), .B(new_n2868_), .ZN(new_n2869_));
  NOR2_X1    g02677(.A1(new_n2869_), .A2(new_n2866_), .ZN(new_n2870_));
  AOI22_X1   g02678(.A1(new_n2867_), .A2(\asqrt[48] ), .B1(new_n2860_), .B2(new_n2865_), .ZN(new_n2871_));
  INV_X1     g02679(.I(new_n2767_), .ZN(new_n2872_));
  OAI21_X1   g02680(.A1(new_n2871_), .A2(new_n1854_), .B(new_n2872_), .ZN(new_n2873_));
  NAND2_X1   g02681(.A1(new_n2873_), .A2(new_n2870_), .ZN(new_n2874_));
  OAI22_X1   g02682(.A1(new_n2871_), .A2(new_n1854_), .B1(new_n2869_), .B2(new_n2866_), .ZN(new_n2875_));
  AOI21_X1   g02683(.A1(new_n2875_), .A2(\asqrt[50] ), .B(new_n2773_), .ZN(new_n2876_));
  NOR2_X1    g02684(.A1(new_n2876_), .A2(new_n2874_), .ZN(new_n2877_));
  AOI22_X1   g02685(.A1(new_n2875_), .A2(\asqrt[50] ), .B1(new_n2873_), .B2(new_n2870_), .ZN(new_n2878_));
  INV_X1     g02686(.I(new_n2781_), .ZN(new_n2879_));
  OAI21_X1   g02687(.A1(new_n2878_), .A2(new_n1436_), .B(new_n2879_), .ZN(new_n2880_));
  NAND2_X1   g02688(.A1(new_n2880_), .A2(new_n2877_), .ZN(new_n2881_));
  OAI22_X1   g02689(.A1(new_n2878_), .A2(new_n1436_), .B1(new_n2876_), .B2(new_n2874_), .ZN(new_n2882_));
  AOI21_X1   g02690(.A1(new_n2882_), .A2(\asqrt[52] ), .B(new_n2787_), .ZN(new_n2883_));
  NOR2_X1    g02691(.A1(new_n2883_), .A2(new_n2881_), .ZN(new_n2884_));
  AOI22_X1   g02692(.A1(new_n2882_), .A2(\asqrt[52] ), .B1(new_n2880_), .B2(new_n2877_), .ZN(new_n2885_));
  INV_X1     g02693(.I(new_n2794_), .ZN(new_n2886_));
  OAI21_X1   g02694(.A1(new_n2885_), .A2(new_n1096_), .B(new_n2886_), .ZN(new_n2887_));
  NAND2_X1   g02695(.A1(new_n2887_), .A2(new_n2884_), .ZN(new_n2888_));
  OAI22_X1   g02696(.A1(new_n2885_), .A2(new_n1096_), .B1(new_n2883_), .B2(new_n2881_), .ZN(new_n2889_));
  AOI21_X1   g02697(.A1(new_n2889_), .A2(\asqrt[54] ), .B(new_n2800_), .ZN(new_n2890_));
  NOR2_X1    g02698(.A1(new_n2890_), .A2(new_n2888_), .ZN(new_n2891_));
  AOI22_X1   g02699(.A1(new_n2889_), .A2(\asqrt[54] ), .B1(new_n2887_), .B2(new_n2884_), .ZN(new_n2892_));
  INV_X1     g02700(.I(new_n2807_), .ZN(new_n2893_));
  OAI21_X1   g02701(.A1(new_n2892_), .A2(new_n825_), .B(new_n2893_), .ZN(new_n2894_));
  NAND2_X1   g02702(.A1(new_n2894_), .A2(new_n2891_), .ZN(new_n2895_));
  OAI22_X1   g02703(.A1(new_n2892_), .A2(new_n825_), .B1(new_n2890_), .B2(new_n2888_), .ZN(new_n2896_));
  AOI21_X1   g02704(.A1(new_n2896_), .A2(\asqrt[56] ), .B(new_n2813_), .ZN(new_n2897_));
  NOR2_X1    g02705(.A1(new_n2897_), .A2(new_n2895_), .ZN(new_n2898_));
  AOI22_X1   g02706(.A1(new_n2896_), .A2(\asqrt[56] ), .B1(new_n2894_), .B2(new_n2891_), .ZN(new_n2899_));
  INV_X1     g02707(.I(new_n2820_), .ZN(new_n2900_));
  OAI21_X1   g02708(.A1(new_n2899_), .A2(new_n587_), .B(new_n2900_), .ZN(new_n2901_));
  NAND2_X1   g02709(.A1(new_n2901_), .A2(new_n2898_), .ZN(new_n2902_));
  OAI22_X1   g02710(.A1(new_n2899_), .A2(new_n587_), .B1(new_n2897_), .B2(new_n2895_), .ZN(new_n2903_));
  AOI21_X1   g02711(.A1(new_n2903_), .A2(\asqrt[58] ), .B(new_n2826_), .ZN(new_n2904_));
  NOR2_X1    g02712(.A1(new_n2904_), .A2(new_n2902_), .ZN(new_n2905_));
  AOI22_X1   g02713(.A1(new_n2903_), .A2(\asqrt[58] ), .B1(new_n2901_), .B2(new_n2898_), .ZN(new_n2906_));
  INV_X1     g02714(.I(new_n2833_), .ZN(new_n2907_));
  OAI21_X1   g02715(.A1(new_n2906_), .A2(new_n376_), .B(new_n2907_), .ZN(new_n2908_));
  NAND2_X1   g02716(.A1(new_n2908_), .A2(new_n2905_), .ZN(new_n2909_));
  OAI22_X1   g02717(.A1(new_n2906_), .A2(new_n376_), .B1(new_n2904_), .B2(new_n2902_), .ZN(new_n2910_));
  AOI21_X1   g02718(.A1(new_n2910_), .A2(\asqrt[60] ), .B(new_n2839_), .ZN(new_n2911_));
  AOI22_X1   g02719(.A1(new_n2910_), .A2(\asqrt[60] ), .B1(new_n2908_), .B2(new_n2905_), .ZN(new_n2912_));
  OAI22_X1   g02720(.A1(new_n2912_), .A2(new_n229_), .B1(new_n2911_), .B2(new_n2909_), .ZN(new_n2913_));
  NOR4_X1    g02721(.A1(new_n2913_), .A2(\asqrt[62] ), .A3(new_n2694_), .A4(new_n2698_), .ZN(new_n2914_));
  AOI21_X1   g02722(.A1(new_n2450_), .A2(new_n2715_), .B(new_n2728_), .ZN(new_n2915_));
  XOR2_X1    g02723(.A1(new_n2715_), .A2(\asqrt[63] ), .Z(new_n2916_));
  NOR2_X1    g02724(.A1(new_n2915_), .A2(new_n2916_), .ZN(new_n2917_));
  NAND2_X1   g02725(.A1(new_n2914_), .A2(new_n2917_), .ZN(new_n2918_));
  NOR4_X1    g02726(.A1(new_n2918_), .A2(new_n2675_), .A3(new_n2682_), .A4(new_n2852_), .ZN(new_n2919_));
  NOR2_X1    g02727(.A1(new_n2675_), .A2(\a[88] ), .ZN(new_n2920_));
  OAI21_X1   g02728(.A1(new_n2919_), .A2(new_n2920_), .B(new_n2674_), .ZN(new_n2921_));
  INV_X1     g02729(.I(new_n2674_), .ZN(new_n2922_));
  INV_X1     g02730(.I(new_n2682_), .ZN(new_n2923_));
  NOR2_X1    g02731(.A1(new_n2911_), .A2(new_n2909_), .ZN(new_n2924_));
  NOR3_X1    g02732(.A1(new_n2912_), .A2(new_n229_), .A3(new_n2845_), .ZN(new_n2925_));
  AOI21_X1   g02733(.A1(new_n2925_), .A2(new_n2924_), .B(new_n2699_), .ZN(new_n2926_));
  AOI21_X1   g02734(.A1(new_n2926_), .A2(new_n2850_), .B(new_n2694_), .ZN(new_n2927_));
  AOI22_X1   g02735(.A1(new_n2843_), .A2(\asqrt[61] ), .B1(new_n2841_), .B2(new_n2835_), .ZN(new_n2928_));
  NAND4_X1   g02736(.A1(new_n2928_), .A2(new_n196_), .A3(new_n2695_), .A4(new_n2844_), .ZN(new_n2929_));
  INV_X1     g02737(.I(new_n2917_), .ZN(new_n2930_));
  NOR2_X1    g02738(.A1(new_n2929_), .A2(new_n2930_), .ZN(new_n2931_));
  NAND4_X1   g02739(.A1(new_n2931_), .A2(new_n2927_), .A3(\a[89] ), .A4(new_n2923_), .ZN(new_n2932_));
  NAND3_X1   g02740(.A1(new_n2932_), .A2(\a[88] ), .A3(new_n2922_), .ZN(new_n2933_));
  NAND2_X1   g02741(.A1(new_n2921_), .A2(new_n2933_), .ZN(new_n2934_));
  NOR2_X1    g02742(.A1(new_n2918_), .A2(new_n2852_), .ZN(new_n2935_));
  NOR4_X1    g02743(.A1(new_n2680_), .A2(new_n2450_), .A3(new_n2730_), .A4(new_n2667_), .ZN(new_n2936_));
  NAND2_X1   g02744(.A1(\asqrt[45] ), .A2(\a[88] ), .ZN(new_n2937_));
  XOR2_X1    g02745(.A1(new_n2937_), .A2(new_n2936_), .Z(new_n2938_));
  NOR2_X1    g02746(.A1(new_n2938_), .A2(new_n2671_), .ZN(new_n2939_));
  INV_X1     g02747(.I(new_n2939_), .ZN(new_n2940_));
  NAND3_X1   g02748(.A1(new_n2931_), .A2(new_n2927_), .A3(new_n2923_), .ZN(new_n2941_));
  NAND2_X1   g02749(.A1(new_n2804_), .A2(\asqrt[55] ), .ZN(new_n2942_));
  AOI21_X1   g02750(.A1(new_n2942_), .A2(new_n2803_), .B(new_n724_), .ZN(new_n2943_));
  OAI21_X1   g02751(.A1(new_n2809_), .A2(new_n2943_), .B(\asqrt[57] ), .ZN(new_n2944_));
  AOI21_X1   g02752(.A1(new_n2816_), .A2(new_n2944_), .B(new_n504_), .ZN(new_n2945_));
  OAI21_X1   g02753(.A1(new_n2822_), .A2(new_n2945_), .B(\asqrt[59] ), .ZN(new_n2946_));
  AOI21_X1   g02754(.A1(new_n2829_), .A2(new_n2946_), .B(new_n275_), .ZN(new_n2947_));
  OAI21_X1   g02755(.A1(new_n2835_), .A2(new_n2947_), .B(\asqrt[61] ), .ZN(new_n2948_));
  NOR3_X1    g02756(.A1(new_n2842_), .A2(new_n2948_), .A3(new_n2845_), .ZN(new_n2949_));
  NOR3_X1    g02757(.A1(new_n2949_), .A2(new_n2699_), .A3(new_n2851_), .ZN(new_n2950_));
  OAI21_X1   g02758(.A1(new_n2950_), .A2(new_n2694_), .B(new_n2929_), .ZN(new_n2951_));
  NOR2_X1    g02759(.A1(new_n2917_), .A2(new_n2923_), .ZN(new_n2952_));
  NAND2_X1   g02760(.A1(new_n2952_), .A2(\asqrt[45] ), .ZN(new_n2953_));
  OAI21_X1   g02761(.A1(new_n2951_), .A2(new_n2953_), .B(new_n2702_), .ZN(new_n2954_));
  NAND3_X1   g02762(.A1(new_n2954_), .A2(new_n2705_), .A3(new_n2941_), .ZN(new_n2955_));
  NOR3_X1    g02763(.A1(new_n2918_), .A2(new_n2682_), .A3(new_n2852_), .ZN(\asqrt[44] ));
  NAND2_X1   g02764(.A1(new_n2889_), .A2(\asqrt[54] ), .ZN(new_n2957_));
  AOI21_X1   g02765(.A1(new_n2957_), .A2(new_n2888_), .B(new_n825_), .ZN(new_n2958_));
  OAI21_X1   g02766(.A1(new_n2891_), .A2(new_n2958_), .B(\asqrt[56] ), .ZN(new_n2959_));
  AOI21_X1   g02767(.A1(new_n2895_), .A2(new_n2959_), .B(new_n587_), .ZN(new_n2960_));
  OAI21_X1   g02768(.A1(new_n2898_), .A2(new_n2960_), .B(\asqrt[58] ), .ZN(new_n2961_));
  AOI21_X1   g02769(.A1(new_n2902_), .A2(new_n2961_), .B(new_n376_), .ZN(new_n2962_));
  OAI21_X1   g02770(.A1(new_n2905_), .A2(new_n2962_), .B(\asqrt[60] ), .ZN(new_n2963_));
  AOI21_X1   g02771(.A1(new_n2909_), .A2(new_n2963_), .B(new_n229_), .ZN(new_n2964_));
  NAND4_X1   g02772(.A1(new_n2964_), .A2(new_n2835_), .A3(new_n2841_), .A4(new_n2846_), .ZN(new_n2965_));
  NAND3_X1   g02773(.A1(new_n2965_), .A2(new_n2700_), .A3(new_n2850_), .ZN(new_n2966_));
  AOI21_X1   g02774(.A1(new_n2695_), .A2(new_n2966_), .B(new_n2914_), .ZN(new_n2967_));
  INV_X1     g02775(.I(new_n2953_), .ZN(new_n2968_));
  AOI21_X1   g02776(.A1(new_n2967_), .A2(new_n2968_), .B(\a[90] ), .ZN(new_n2969_));
  OAI21_X1   g02777(.A1(new_n2969_), .A2(new_n2706_), .B(\asqrt[44] ), .ZN(new_n2970_));
  NAND4_X1   g02778(.A1(new_n2970_), .A2(new_n2955_), .A3(new_n2488_), .A4(new_n2940_), .ZN(new_n2971_));
  NAND2_X1   g02779(.A1(new_n2971_), .A2(new_n2934_), .ZN(new_n2972_));
  NAND3_X1   g02780(.A1(new_n2921_), .A2(new_n2933_), .A3(new_n2940_), .ZN(new_n2973_));
  NAND2_X1   g02781(.A1(\asqrt[45] ), .A2(new_n2702_), .ZN(new_n2974_));
  AOI22_X1   g02782(.A1(new_n2974_), .A2(new_n2701_), .B1(new_n2702_), .B2(new_n2709_), .ZN(new_n2975_));
  OAI21_X1   g02783(.A1(new_n2728_), .A2(new_n2702_), .B(new_n2707_), .ZN(new_n2976_));
  NOR2_X1    g02784(.A1(new_n2975_), .A2(new_n2976_), .ZN(new_n2977_));
  NAND3_X1   g02785(.A1(\asqrt[44] ), .A2(new_n2727_), .A3(new_n2977_), .ZN(new_n2978_));
  INV_X1     g02786(.I(new_n2977_), .ZN(new_n2979_));
  OAI21_X1   g02787(.A1(new_n2941_), .A2(new_n2979_), .B(new_n2726_), .ZN(new_n2980_));
  NAND3_X1   g02788(.A1(new_n2978_), .A2(new_n2980_), .A3(new_n2253_), .ZN(new_n2981_));
  AOI21_X1   g02789(.A1(new_n2973_), .A2(\asqrt[46] ), .B(new_n2981_), .ZN(new_n2982_));
  NOR2_X1    g02790(.A1(new_n2972_), .A2(new_n2982_), .ZN(new_n2983_));
  NAND2_X1   g02791(.A1(new_n2973_), .A2(\asqrt[46] ), .ZN(new_n2984_));
  AOI21_X1   g02792(.A1(new_n2972_), .A2(new_n2984_), .B(new_n2253_), .ZN(new_n2985_));
  NOR2_X1    g02793(.A1(new_n2858_), .A2(new_n2857_), .ZN(new_n2986_));
  NOR4_X1    g02794(.A1(new_n2941_), .A2(\asqrt[47] ), .A3(new_n2986_), .A4(new_n2741_), .ZN(new_n2987_));
  AOI21_X1   g02795(.A1(new_n2856_), .A2(new_n2727_), .B(new_n2253_), .ZN(new_n2988_));
  NOR2_X1    g02796(.A1(new_n2987_), .A2(new_n2988_), .ZN(new_n2989_));
  NAND2_X1   g02797(.A1(new_n2989_), .A2(new_n2046_), .ZN(new_n2990_));
  OAI21_X1   g02798(.A1(new_n2985_), .A2(new_n2990_), .B(new_n2983_), .ZN(new_n2991_));
  OAI21_X1   g02799(.A1(new_n2985_), .A2(new_n2983_), .B(\asqrt[48] ), .ZN(new_n2992_));
  NOR2_X1    g02800(.A1(new_n2752_), .A2(new_n2046_), .ZN(new_n2993_));
  NAND2_X1   g02801(.A1(new_n2747_), .A2(new_n2748_), .ZN(new_n2994_));
  NAND4_X1   g02802(.A1(\asqrt[44] ), .A2(new_n2046_), .A3(new_n2994_), .A4(new_n2752_), .ZN(new_n2995_));
  XOR2_X1    g02803(.A1(new_n2995_), .A2(new_n2993_), .Z(new_n2996_));
  NAND2_X1   g02804(.A1(new_n2996_), .A2(new_n1854_), .ZN(new_n2997_));
  INV_X1     g02805(.I(new_n2997_), .ZN(new_n2998_));
  AOI21_X1   g02806(.A1(new_n2992_), .A2(new_n2998_), .B(new_n2991_), .ZN(new_n2999_));
  AOI21_X1   g02807(.A1(new_n2991_), .A2(new_n2992_), .B(new_n1854_), .ZN(new_n3000_));
  NAND2_X1   g02808(.A1(new_n2763_), .A2(\asqrt[49] ), .ZN(new_n3001_));
  NOR2_X1    g02809(.A1(new_n2758_), .A2(new_n2759_), .ZN(new_n3002_));
  NOR4_X1    g02810(.A1(new_n2941_), .A2(\asqrt[49] ), .A3(new_n3002_), .A4(new_n2763_), .ZN(new_n3003_));
  XOR2_X1    g02811(.A1(new_n3003_), .A2(new_n3001_), .Z(new_n3004_));
  NAND2_X1   g02812(.A1(new_n3004_), .A2(new_n1595_), .ZN(new_n3005_));
  OAI21_X1   g02813(.A1(new_n3000_), .A2(new_n3005_), .B(new_n2999_), .ZN(new_n3006_));
  AOI22_X1   g02814(.A1(new_n2971_), .A2(new_n2934_), .B1(\asqrt[46] ), .B2(new_n2973_), .ZN(new_n3007_));
  OAI22_X1   g02815(.A1(new_n3007_), .A2(new_n2253_), .B1(new_n2972_), .B2(new_n2982_), .ZN(new_n3008_));
  AOI21_X1   g02816(.A1(new_n3008_), .A2(\asqrt[48] ), .B(new_n2997_), .ZN(new_n3009_));
  INV_X1     g02817(.I(new_n2990_), .ZN(new_n3010_));
  OAI21_X1   g02818(.A1(new_n3007_), .A2(new_n2253_), .B(new_n3010_), .ZN(new_n3011_));
  AOI22_X1   g02819(.A1(new_n3008_), .A2(\asqrt[48] ), .B1(new_n3011_), .B2(new_n2983_), .ZN(new_n3012_));
  OAI22_X1   g02820(.A1(new_n3012_), .A2(new_n1854_), .B1(new_n3009_), .B2(new_n2991_), .ZN(new_n3013_));
  NOR4_X1    g02821(.A1(new_n2941_), .A2(\asqrt[50] ), .A3(new_n2766_), .A4(new_n2875_), .ZN(new_n3014_));
  AOI21_X1   g02822(.A1(new_n3001_), .A2(new_n2762_), .B(new_n1595_), .ZN(new_n3015_));
  NOR2_X1    g02823(.A1(new_n3014_), .A2(new_n3015_), .ZN(new_n3016_));
  NAND2_X1   g02824(.A1(new_n3016_), .A2(new_n1436_), .ZN(new_n3017_));
  AOI21_X1   g02825(.A1(new_n3013_), .A2(\asqrt[50] ), .B(new_n3017_), .ZN(new_n3018_));
  NOR2_X1    g02826(.A1(new_n3018_), .A2(new_n3006_), .ZN(new_n3019_));
  INV_X1     g02827(.I(new_n3005_), .ZN(new_n3020_));
  OAI21_X1   g02828(.A1(new_n3012_), .A2(new_n1854_), .B(new_n3020_), .ZN(new_n3021_));
  AOI22_X1   g02829(.A1(new_n3013_), .A2(\asqrt[50] ), .B1(new_n3021_), .B2(new_n2999_), .ZN(new_n3022_));
  NAND2_X1   g02830(.A1(new_n2777_), .A2(\asqrt[51] ), .ZN(new_n3023_));
  NOR4_X1    g02831(.A1(new_n2941_), .A2(\asqrt[51] ), .A3(new_n2772_), .A4(new_n2777_), .ZN(new_n3024_));
  XOR2_X1    g02832(.A1(new_n3024_), .A2(new_n3023_), .Z(new_n3025_));
  NAND2_X1   g02833(.A1(new_n3025_), .A2(new_n1260_), .ZN(new_n3026_));
  INV_X1     g02834(.I(new_n3026_), .ZN(new_n3027_));
  OAI21_X1   g02835(.A1(new_n3022_), .A2(new_n1436_), .B(new_n3027_), .ZN(new_n3028_));
  NAND2_X1   g02836(.A1(new_n3028_), .A2(new_n3019_), .ZN(new_n3029_));
  OAI22_X1   g02837(.A1(new_n3022_), .A2(new_n1436_), .B1(new_n3018_), .B2(new_n3006_), .ZN(new_n3030_));
  NOR4_X1    g02838(.A1(new_n2941_), .A2(\asqrt[52] ), .A3(new_n2780_), .A4(new_n2882_), .ZN(new_n3031_));
  AOI21_X1   g02839(.A1(new_n3023_), .A2(new_n2776_), .B(new_n1260_), .ZN(new_n3032_));
  NOR2_X1    g02840(.A1(new_n3031_), .A2(new_n3032_), .ZN(new_n3033_));
  NAND2_X1   g02841(.A1(new_n3033_), .A2(new_n1096_), .ZN(new_n3034_));
  AOI21_X1   g02842(.A1(new_n3030_), .A2(\asqrt[52] ), .B(new_n3034_), .ZN(new_n3035_));
  NOR2_X1    g02843(.A1(new_n3035_), .A2(new_n3029_), .ZN(new_n3036_));
  AOI22_X1   g02844(.A1(new_n3030_), .A2(\asqrt[52] ), .B1(new_n3028_), .B2(new_n3019_), .ZN(new_n3037_));
  NOR2_X1    g02845(.A1(new_n2885_), .A2(new_n1096_), .ZN(new_n3038_));
  NOR4_X1    g02846(.A1(new_n2941_), .A2(\asqrt[53] ), .A3(new_n2786_), .A4(new_n2791_), .ZN(new_n3039_));
  XNOR2_X1   g02847(.A1(new_n3039_), .A2(new_n3038_), .ZN(new_n3040_));
  NAND2_X1   g02848(.A1(new_n3040_), .A2(new_n970_), .ZN(new_n3041_));
  INV_X1     g02849(.I(new_n3041_), .ZN(new_n3042_));
  OAI21_X1   g02850(.A1(new_n3037_), .A2(new_n1096_), .B(new_n3042_), .ZN(new_n3043_));
  NAND2_X1   g02851(.A1(new_n3043_), .A2(new_n3036_), .ZN(new_n3044_));
  OAI22_X1   g02852(.A1(new_n3037_), .A2(new_n1096_), .B1(new_n3035_), .B2(new_n3029_), .ZN(new_n3045_));
  NOR4_X1    g02853(.A1(new_n2941_), .A2(\asqrt[54] ), .A3(new_n2793_), .A4(new_n2889_), .ZN(new_n3046_));
  XOR2_X1    g02854(.A1(new_n3046_), .A2(new_n2957_), .Z(new_n3047_));
  NAND2_X1   g02855(.A1(new_n3047_), .A2(new_n825_), .ZN(new_n3048_));
  AOI21_X1   g02856(.A1(new_n3045_), .A2(\asqrt[54] ), .B(new_n3048_), .ZN(new_n3049_));
  NOR2_X1    g02857(.A1(new_n3049_), .A2(new_n3044_), .ZN(new_n3050_));
  AOI22_X1   g02858(.A1(new_n3045_), .A2(\asqrt[54] ), .B1(new_n3043_), .B2(new_n3036_), .ZN(new_n3051_));
  NOR4_X1    g02859(.A1(new_n2941_), .A2(\asqrt[55] ), .A3(new_n2799_), .A4(new_n2804_), .ZN(new_n3052_));
  XOR2_X1    g02860(.A1(new_n3052_), .A2(new_n2942_), .Z(new_n3053_));
  NAND2_X1   g02861(.A1(new_n3053_), .A2(new_n724_), .ZN(new_n3054_));
  INV_X1     g02862(.I(new_n3054_), .ZN(new_n3055_));
  OAI21_X1   g02863(.A1(new_n3051_), .A2(new_n825_), .B(new_n3055_), .ZN(new_n3056_));
  NAND2_X1   g02864(.A1(new_n3056_), .A2(new_n3050_), .ZN(new_n3057_));
  OAI22_X1   g02865(.A1(new_n3051_), .A2(new_n825_), .B1(new_n3049_), .B2(new_n3044_), .ZN(new_n3058_));
  NOR4_X1    g02866(.A1(new_n2941_), .A2(\asqrt[56] ), .A3(new_n2806_), .A4(new_n2896_), .ZN(new_n3059_));
  XOR2_X1    g02867(.A1(new_n3059_), .A2(new_n2959_), .Z(new_n3060_));
  NAND2_X1   g02868(.A1(new_n3060_), .A2(new_n587_), .ZN(new_n3061_));
  AOI21_X1   g02869(.A1(new_n3058_), .A2(\asqrt[56] ), .B(new_n3061_), .ZN(new_n3062_));
  NOR2_X1    g02870(.A1(new_n3062_), .A2(new_n3057_), .ZN(new_n3063_));
  AOI22_X1   g02871(.A1(new_n3058_), .A2(\asqrt[56] ), .B1(new_n3056_), .B2(new_n3050_), .ZN(new_n3064_));
  NOR4_X1    g02872(.A1(new_n2941_), .A2(\asqrt[57] ), .A3(new_n2812_), .A4(new_n2817_), .ZN(new_n3065_));
  XOR2_X1    g02873(.A1(new_n3065_), .A2(new_n2944_), .Z(new_n3066_));
  NAND2_X1   g02874(.A1(new_n3066_), .A2(new_n504_), .ZN(new_n3067_));
  INV_X1     g02875(.I(new_n3067_), .ZN(new_n3068_));
  OAI21_X1   g02876(.A1(new_n3064_), .A2(new_n587_), .B(new_n3068_), .ZN(new_n3069_));
  NAND2_X1   g02877(.A1(new_n3069_), .A2(new_n3063_), .ZN(new_n3070_));
  OAI22_X1   g02878(.A1(new_n3064_), .A2(new_n587_), .B1(new_n3062_), .B2(new_n3057_), .ZN(new_n3071_));
  NOR4_X1    g02879(.A1(new_n2941_), .A2(\asqrt[58] ), .A3(new_n2819_), .A4(new_n2903_), .ZN(new_n3072_));
  XOR2_X1    g02880(.A1(new_n3072_), .A2(new_n2961_), .Z(new_n3073_));
  NAND2_X1   g02881(.A1(new_n3073_), .A2(new_n376_), .ZN(new_n3074_));
  AOI21_X1   g02882(.A1(new_n3071_), .A2(\asqrt[58] ), .B(new_n3074_), .ZN(new_n3075_));
  NOR2_X1    g02883(.A1(new_n3075_), .A2(new_n3070_), .ZN(new_n3076_));
  AOI22_X1   g02884(.A1(new_n3071_), .A2(\asqrt[58] ), .B1(new_n3069_), .B2(new_n3063_), .ZN(new_n3077_));
  NOR4_X1    g02885(.A1(new_n2941_), .A2(\asqrt[59] ), .A3(new_n2825_), .A4(new_n2830_), .ZN(new_n3078_));
  XOR2_X1    g02886(.A1(new_n3078_), .A2(new_n2946_), .Z(new_n3079_));
  AND2_X2    g02887(.A1(new_n3079_), .A2(new_n275_), .Z(new_n3080_));
  OAI21_X1   g02888(.A1(new_n3077_), .A2(new_n376_), .B(new_n3080_), .ZN(new_n3081_));
  NAND2_X1   g02889(.A1(new_n3081_), .A2(new_n3076_), .ZN(new_n3082_));
  NAND2_X1   g02890(.A1(new_n3045_), .A2(\asqrt[54] ), .ZN(new_n3083_));
  AOI21_X1   g02891(.A1(new_n3083_), .A2(new_n3044_), .B(new_n825_), .ZN(new_n3084_));
  OAI21_X1   g02892(.A1(new_n3050_), .A2(new_n3084_), .B(\asqrt[56] ), .ZN(new_n3085_));
  AOI21_X1   g02893(.A1(new_n3057_), .A2(new_n3085_), .B(new_n587_), .ZN(new_n3086_));
  OAI21_X1   g02894(.A1(new_n3063_), .A2(new_n3086_), .B(\asqrt[58] ), .ZN(new_n3087_));
  AOI21_X1   g02895(.A1(new_n3070_), .A2(new_n3087_), .B(new_n376_), .ZN(new_n3088_));
  OAI21_X1   g02896(.A1(new_n3076_), .A2(new_n3088_), .B(\asqrt[60] ), .ZN(new_n3089_));
  AOI21_X1   g02897(.A1(new_n3082_), .A2(new_n3089_), .B(new_n229_), .ZN(new_n3090_));
  NOR2_X1    g02898(.A1(new_n2928_), .A2(new_n196_), .ZN(new_n3091_));
  NOR2_X1    g02899(.A1(new_n2913_), .A2(\asqrt[62] ), .ZN(new_n3092_));
  NAND3_X1   g02900(.A1(new_n3092_), .A2(new_n3091_), .A3(new_n2844_), .ZN(new_n3093_));
  NOR2_X1    g02901(.A1(new_n2941_), .A2(new_n3093_), .ZN(new_n3094_));
  OR3_X2     g02902(.A1(\asqrt[44] ), .A2(new_n2844_), .A3(new_n3092_), .Z(new_n3095_));
  AOI21_X1   g02903(.A1(new_n3095_), .A2(new_n3091_), .B(new_n3094_), .ZN(new_n3096_));
  NOR3_X1    g02904(.A1(new_n2843_), .A2(\asqrt[61] ), .A3(new_n2838_), .ZN(new_n3097_));
  NAND2_X1   g02905(.A1(\asqrt[44] ), .A2(new_n3097_), .ZN(new_n3098_));
  XOR2_X1    g02906(.A1(new_n3098_), .A2(new_n2964_), .Z(new_n3099_));
  NOR2_X1    g02907(.A1(new_n3099_), .A2(new_n196_), .ZN(new_n3100_));
  INV_X1     g02908(.I(new_n3100_), .ZN(new_n3101_));
  NOR2_X1    g02909(.A1(new_n3000_), .A2(new_n3005_), .ZN(new_n3102_));
  NOR3_X1    g02910(.A1(new_n3102_), .A2(new_n2991_), .A3(new_n3009_), .ZN(new_n3103_));
  OAI21_X1   g02911(.A1(new_n2999_), .A2(new_n3000_), .B(\asqrt[50] ), .ZN(new_n3104_));
  INV_X1     g02912(.I(new_n3017_), .ZN(new_n3105_));
  NAND2_X1   g02913(.A1(new_n3104_), .A2(new_n3105_), .ZN(new_n3106_));
  NAND2_X1   g02914(.A1(new_n3106_), .A2(new_n3103_), .ZN(new_n3107_));
  NAND2_X1   g02915(.A1(new_n3006_), .A2(new_n3104_), .ZN(new_n3108_));
  AOI21_X1   g02916(.A1(new_n3108_), .A2(\asqrt[51] ), .B(new_n3026_), .ZN(new_n3109_));
  NOR2_X1    g02917(.A1(new_n3109_), .A2(new_n3107_), .ZN(new_n3110_));
  AOI22_X1   g02918(.A1(new_n3108_), .A2(\asqrt[51] ), .B1(new_n3106_), .B2(new_n3103_), .ZN(new_n3111_));
  INV_X1     g02919(.I(new_n3034_), .ZN(new_n3112_));
  OAI21_X1   g02920(.A1(new_n3111_), .A2(new_n1260_), .B(new_n3112_), .ZN(new_n3113_));
  NAND2_X1   g02921(.A1(new_n3113_), .A2(new_n3110_), .ZN(new_n3114_));
  OAI22_X1   g02922(.A1(new_n3111_), .A2(new_n1260_), .B1(new_n3109_), .B2(new_n3107_), .ZN(new_n3115_));
  AOI21_X1   g02923(.A1(new_n3115_), .A2(\asqrt[53] ), .B(new_n3041_), .ZN(new_n3116_));
  NOR2_X1    g02924(.A1(new_n3116_), .A2(new_n3114_), .ZN(new_n3117_));
  AOI22_X1   g02925(.A1(new_n3115_), .A2(\asqrt[53] ), .B1(new_n3113_), .B2(new_n3110_), .ZN(new_n3118_));
  INV_X1     g02926(.I(new_n3048_), .ZN(new_n3119_));
  OAI21_X1   g02927(.A1(new_n3118_), .A2(new_n970_), .B(new_n3119_), .ZN(new_n3120_));
  NAND2_X1   g02928(.A1(new_n3120_), .A2(new_n3117_), .ZN(new_n3121_));
  OAI22_X1   g02929(.A1(new_n3118_), .A2(new_n970_), .B1(new_n3116_), .B2(new_n3114_), .ZN(new_n3122_));
  AOI21_X1   g02930(.A1(new_n3122_), .A2(\asqrt[55] ), .B(new_n3054_), .ZN(new_n3123_));
  NOR2_X1    g02931(.A1(new_n3123_), .A2(new_n3121_), .ZN(new_n3124_));
  AOI22_X1   g02932(.A1(new_n3122_), .A2(\asqrt[55] ), .B1(new_n3120_), .B2(new_n3117_), .ZN(new_n3125_));
  INV_X1     g02933(.I(new_n3061_), .ZN(new_n3126_));
  OAI21_X1   g02934(.A1(new_n3125_), .A2(new_n724_), .B(new_n3126_), .ZN(new_n3127_));
  NAND2_X1   g02935(.A1(new_n3127_), .A2(new_n3124_), .ZN(new_n3128_));
  NAND2_X1   g02936(.A1(new_n3115_), .A2(\asqrt[53] ), .ZN(new_n3129_));
  AOI21_X1   g02937(.A1(new_n3129_), .A2(new_n3114_), .B(new_n970_), .ZN(new_n3130_));
  OAI21_X1   g02938(.A1(new_n3117_), .A2(new_n3130_), .B(\asqrt[55] ), .ZN(new_n3131_));
  AOI21_X1   g02939(.A1(new_n3121_), .A2(new_n3131_), .B(new_n724_), .ZN(new_n3132_));
  OAI21_X1   g02940(.A1(new_n3124_), .A2(new_n3132_), .B(\asqrt[57] ), .ZN(new_n3133_));
  AOI21_X1   g02941(.A1(new_n3133_), .A2(new_n3068_), .B(new_n3128_), .ZN(new_n3134_));
  OAI22_X1   g02942(.A1(new_n3125_), .A2(new_n724_), .B1(new_n3123_), .B2(new_n3121_), .ZN(new_n3135_));
  AOI22_X1   g02943(.A1(new_n3135_), .A2(\asqrt[57] ), .B1(new_n3127_), .B2(new_n3124_), .ZN(new_n3136_));
  INV_X1     g02944(.I(new_n3074_), .ZN(new_n3137_));
  OAI21_X1   g02945(.A1(new_n3136_), .A2(new_n504_), .B(new_n3137_), .ZN(new_n3138_));
  NAND2_X1   g02946(.A1(new_n3138_), .A2(new_n3134_), .ZN(new_n3139_));
  AOI21_X1   g02947(.A1(new_n3128_), .A2(new_n3133_), .B(new_n504_), .ZN(new_n3140_));
  OAI21_X1   g02948(.A1(new_n3134_), .A2(new_n3140_), .B(\asqrt[59] ), .ZN(new_n3141_));
  AOI21_X1   g02949(.A1(new_n3141_), .A2(new_n3080_), .B(new_n3139_), .ZN(new_n3142_));
  NAND2_X1   g02950(.A1(new_n3070_), .A2(new_n3087_), .ZN(new_n3143_));
  AOI22_X1   g02951(.A1(new_n3143_), .A2(\asqrt[59] ), .B1(new_n3138_), .B2(new_n3134_), .ZN(new_n3144_));
  NOR4_X1    g02952(.A1(new_n2941_), .A2(\asqrt[60] ), .A3(new_n2832_), .A4(new_n2910_), .ZN(new_n3145_));
  XOR2_X1    g02953(.A1(new_n3145_), .A2(new_n2963_), .Z(new_n3146_));
  NAND2_X1   g02954(.A1(new_n3146_), .A2(new_n229_), .ZN(new_n3147_));
  INV_X1     g02955(.I(new_n3147_), .ZN(new_n3148_));
  OAI21_X1   g02956(.A1(new_n3144_), .A2(new_n275_), .B(new_n3148_), .ZN(new_n3149_));
  NAND2_X1   g02957(.A1(new_n3149_), .A2(new_n3142_), .ZN(new_n3150_));
  INV_X1     g02958(.I(new_n3099_), .ZN(new_n3151_));
  NOR2_X1    g02959(.A1(new_n3151_), .A2(\asqrt[62] ), .ZN(new_n3152_));
  INV_X1     g02960(.I(new_n3152_), .ZN(new_n3153_));
  NAND2_X1   g02961(.A1(new_n3090_), .A2(new_n3153_), .ZN(new_n3154_));
  OAI21_X1   g02962(.A1(new_n3154_), .A2(new_n3150_), .B(new_n3101_), .ZN(new_n3155_));
  NAND2_X1   g02963(.A1(new_n2929_), .A2(new_n2694_), .ZN(new_n3156_));
  OAI21_X1   g02964(.A1(\asqrt[44] ), .A2(new_n3156_), .B(new_n2848_), .ZN(new_n3157_));
  NAND2_X1   g02965(.A1(new_n3157_), .A2(new_n231_), .ZN(new_n3158_));
  OAI21_X1   g02966(.A1(new_n3155_), .A2(new_n3158_), .B(new_n3096_), .ZN(new_n3159_));
  OAI21_X1   g02967(.A1(new_n2695_), .A2(new_n2848_), .B(\asqrt[44] ), .ZN(new_n3160_));
  XOR2_X1    g02968(.A1(new_n2848_), .A2(\asqrt[63] ), .Z(new_n3161_));
  NAND2_X1   g02969(.A1(new_n3160_), .A2(new_n3161_), .ZN(new_n3162_));
  INV_X1     g02970(.I(new_n3162_), .ZN(new_n3163_));
  INV_X1     g02971(.I(new_n3096_), .ZN(new_n3164_));
  OAI22_X1   g02972(.A1(new_n3077_), .A2(new_n376_), .B1(new_n3075_), .B2(new_n3070_), .ZN(new_n3165_));
  AOI21_X1   g02973(.A1(new_n3165_), .A2(\asqrt[60] ), .B(new_n3147_), .ZN(new_n3166_));
  AOI22_X1   g02974(.A1(new_n3165_), .A2(\asqrt[60] ), .B1(new_n3081_), .B2(new_n3076_), .ZN(new_n3167_));
  OAI22_X1   g02975(.A1(new_n3167_), .A2(new_n229_), .B1(new_n3166_), .B2(new_n3082_), .ZN(new_n3168_));
  NOR4_X1    g02976(.A1(new_n3168_), .A2(\asqrt[62] ), .A3(new_n3164_), .A4(new_n3099_), .ZN(new_n3169_));
  NAND2_X1   g02977(.A1(new_n3169_), .A2(new_n3163_), .ZN(new_n3170_));
  NAND3_X1   g02978(.A1(new_n2935_), .A2(new_n2682_), .A3(new_n2695_), .ZN(new_n3171_));
  NOR3_X1    g02979(.A1(new_n3170_), .A2(new_n3159_), .A3(new_n3171_), .ZN(\asqrt[43] ));
  NAND2_X1   g02980(.A1(new_n3082_), .A2(new_n3089_), .ZN(new_n3173_));
  NOR3_X1    g02981(.A1(new_n3173_), .A2(\asqrt[61] ), .A3(new_n3146_), .ZN(new_n3174_));
  NAND2_X1   g02982(.A1(\asqrt[43] ), .A2(new_n3174_), .ZN(new_n3175_));
  XOR2_X1    g02983(.A1(new_n3175_), .A2(new_n3090_), .Z(new_n3176_));
  INV_X1     g02984(.I(new_n3176_), .ZN(new_n3177_));
  INV_X1     g02985(.I(\a[87] ), .ZN(new_n3178_));
  INV_X1     g02986(.I(\a[86] ), .ZN(new_n3179_));
  NOR2_X1    g02987(.A1(\a[84] ), .A2(\a[85] ), .ZN(new_n3180_));
  INV_X1     g02988(.I(new_n3180_), .ZN(new_n3181_));
  NOR4_X1    g02989(.A1(new_n2951_), .A2(new_n3179_), .A3(new_n2952_), .A4(new_n3181_), .ZN(new_n3182_));
  XOR2_X1    g02990(.A1(new_n3182_), .A2(new_n3178_), .Z(new_n3183_));
  NOR4_X1    g02991(.A1(new_n3170_), .A2(new_n3159_), .A3(new_n3178_), .A4(new_n3171_), .ZN(new_n3184_));
  NOR2_X1    g02992(.A1(new_n3178_), .A2(\a[86] ), .ZN(new_n3185_));
  OAI21_X1   g02993(.A1(new_n3184_), .A2(new_n3185_), .B(new_n3183_), .ZN(new_n3186_));
  INV_X1     g02994(.I(new_n3183_), .ZN(new_n3187_));
  NOR2_X1    g02995(.A1(new_n3166_), .A2(new_n3082_), .ZN(new_n3188_));
  NOR3_X1    g02996(.A1(new_n3167_), .A2(new_n229_), .A3(new_n3152_), .ZN(new_n3189_));
  AOI21_X1   g02997(.A1(new_n3189_), .A2(new_n3188_), .B(new_n3100_), .ZN(new_n3190_));
  INV_X1     g02998(.I(new_n3158_), .ZN(new_n3191_));
  AOI21_X1   g02999(.A1(new_n3190_), .A2(new_n3191_), .B(new_n3164_), .ZN(new_n3192_));
  AOI21_X1   g03000(.A1(new_n3168_), .A2(\asqrt[62] ), .B(new_n3096_), .ZN(new_n3193_));
  AOI21_X1   g03001(.A1(new_n3139_), .A2(new_n3141_), .B(new_n275_), .ZN(new_n3194_));
  OAI21_X1   g03002(.A1(new_n3142_), .A2(new_n3194_), .B(\asqrt[61] ), .ZN(new_n3195_));
  NAND4_X1   g03003(.A1(new_n3150_), .A2(new_n196_), .A3(new_n3195_), .A4(new_n3151_), .ZN(new_n3196_));
  NOR3_X1    g03004(.A1(new_n3193_), .A2(new_n3162_), .A3(new_n3196_), .ZN(new_n3197_));
  INV_X1     g03005(.I(new_n3171_), .ZN(new_n3198_));
  NAND4_X1   g03006(.A1(new_n3197_), .A2(\a[87] ), .A3(new_n3192_), .A4(new_n3198_), .ZN(new_n3199_));
  NAND3_X1   g03007(.A1(new_n3199_), .A2(\a[86] ), .A3(new_n3187_), .ZN(new_n3200_));
  NAND2_X1   g03008(.A1(new_n3186_), .A2(new_n3200_), .ZN(new_n3201_));
  NOR2_X1    g03009(.A1(new_n3170_), .A2(new_n3159_), .ZN(new_n3202_));
  NOR4_X1    g03010(.A1(new_n2918_), .A2(new_n2682_), .A3(new_n2694_), .A4(new_n2950_), .ZN(new_n3203_));
  NAND2_X1   g03011(.A1(\asqrt[44] ), .A2(\a[86] ), .ZN(new_n3204_));
  XOR2_X1    g03012(.A1(new_n3204_), .A2(new_n3203_), .Z(new_n3205_));
  NOR2_X1    g03013(.A1(new_n3205_), .A2(new_n3181_), .ZN(new_n3206_));
  INV_X1     g03014(.I(new_n3206_), .ZN(new_n3207_));
  NAND3_X1   g03015(.A1(new_n3197_), .A2(new_n3192_), .A3(new_n3198_), .ZN(new_n3208_));
  NOR4_X1    g03016(.A1(new_n3195_), .A2(new_n3082_), .A3(new_n3166_), .A4(new_n3152_), .ZN(new_n3209_));
  NOR3_X1    g03017(.A1(new_n3209_), .A2(new_n3100_), .A3(new_n3158_), .ZN(new_n3210_));
  AOI22_X1   g03018(.A1(new_n3173_), .A2(\asqrt[61] ), .B1(new_n3149_), .B2(new_n3142_), .ZN(new_n3211_));
  NAND4_X1   g03019(.A1(new_n3211_), .A2(new_n196_), .A3(new_n3096_), .A4(new_n3151_), .ZN(new_n3212_));
  OAI21_X1   g03020(.A1(new_n3210_), .A2(new_n3164_), .B(new_n3212_), .ZN(new_n3213_));
  NOR2_X1    g03021(.A1(new_n3163_), .A2(new_n3198_), .ZN(new_n3214_));
  NAND2_X1   g03022(.A1(new_n3214_), .A2(\asqrt[44] ), .ZN(new_n3215_));
  OAI21_X1   g03023(.A1(new_n3213_), .A2(new_n3215_), .B(new_n2662_), .ZN(new_n3216_));
  NAND3_X1   g03024(.A1(new_n3216_), .A2(new_n2670_), .A3(new_n3208_), .ZN(new_n3217_));
  NAND4_X1   g03025(.A1(new_n3090_), .A2(new_n3142_), .A3(new_n3149_), .A4(new_n3153_), .ZN(new_n3218_));
  NAND3_X1   g03026(.A1(new_n3218_), .A2(new_n3101_), .A3(new_n3191_), .ZN(new_n3219_));
  AOI21_X1   g03027(.A1(new_n3096_), .A2(new_n3219_), .B(new_n3169_), .ZN(new_n3220_));
  INV_X1     g03028(.I(new_n3215_), .ZN(new_n3221_));
  AOI21_X1   g03029(.A1(new_n3220_), .A2(new_n3221_), .B(\a[88] ), .ZN(new_n3222_));
  OAI21_X1   g03030(.A1(new_n3222_), .A2(new_n2671_), .B(\asqrt[43] ), .ZN(new_n3223_));
  NAND4_X1   g03031(.A1(new_n3217_), .A2(new_n3223_), .A3(new_n2728_), .A4(new_n3207_), .ZN(new_n3224_));
  NAND2_X1   g03032(.A1(new_n3224_), .A2(new_n3201_), .ZN(new_n3225_));
  NAND3_X1   g03033(.A1(new_n3186_), .A2(new_n3200_), .A3(new_n3207_), .ZN(new_n3226_));
  AOI21_X1   g03034(.A1(\asqrt[44] ), .A2(new_n2662_), .B(\a[89] ), .ZN(new_n3227_));
  NOR2_X1    g03035(.A1(new_n2932_), .A2(\a[88] ), .ZN(new_n3228_));
  AOI21_X1   g03036(.A1(\asqrt[44] ), .A2(\a[88] ), .B(new_n2673_), .ZN(new_n3229_));
  OAI21_X1   g03037(.A1(new_n3227_), .A2(new_n3228_), .B(new_n3229_), .ZN(new_n3230_));
  INV_X1     g03038(.I(new_n3230_), .ZN(new_n3231_));
  NAND3_X1   g03039(.A1(\asqrt[43] ), .A2(new_n2940_), .A3(new_n3231_), .ZN(new_n3232_));
  OAI21_X1   g03040(.A1(new_n3208_), .A2(new_n3230_), .B(new_n2939_), .ZN(new_n3233_));
  NAND3_X1   g03041(.A1(new_n3232_), .A2(new_n3233_), .A3(new_n2488_), .ZN(new_n3234_));
  AOI21_X1   g03042(.A1(new_n3226_), .A2(\asqrt[45] ), .B(new_n3234_), .ZN(new_n3235_));
  NOR2_X1    g03043(.A1(new_n3225_), .A2(new_n3235_), .ZN(new_n3236_));
  AOI22_X1   g03044(.A1(new_n3224_), .A2(new_n3201_), .B1(\asqrt[45] ), .B2(new_n3226_), .ZN(new_n3237_));
  INV_X1     g03045(.I(new_n2973_), .ZN(new_n3238_));
  AOI21_X1   g03046(.A1(new_n2970_), .A2(new_n2955_), .B(\asqrt[46] ), .ZN(new_n3239_));
  AND4_X2    g03047(.A1(new_n3238_), .A2(\asqrt[43] ), .A3(new_n2984_), .A4(new_n3239_), .Z(new_n3240_));
  NOR2_X1    g03048(.A1(new_n3238_), .A2(new_n2488_), .ZN(new_n3241_));
  NOR3_X1    g03049(.A1(new_n3240_), .A2(\asqrt[47] ), .A3(new_n3241_), .ZN(new_n3242_));
  OAI21_X1   g03050(.A1(new_n3237_), .A2(new_n2488_), .B(new_n3242_), .ZN(new_n3243_));
  NAND2_X1   g03051(.A1(new_n3243_), .A2(new_n3236_), .ZN(new_n3244_));
  OAI22_X1   g03052(.A1(new_n3237_), .A2(new_n2488_), .B1(new_n3225_), .B2(new_n3235_), .ZN(new_n3245_));
  NAND2_X1   g03053(.A1(new_n2978_), .A2(new_n2980_), .ZN(new_n3246_));
  NAND4_X1   g03054(.A1(\asqrt[43] ), .A2(new_n2253_), .A3(new_n3246_), .A4(new_n3007_), .ZN(new_n3247_));
  XOR2_X1    g03055(.A1(new_n3247_), .A2(new_n2985_), .Z(new_n3248_));
  NAND2_X1   g03056(.A1(new_n3248_), .A2(new_n2046_), .ZN(new_n3249_));
  AOI21_X1   g03057(.A1(new_n3245_), .A2(\asqrt[47] ), .B(new_n3249_), .ZN(new_n3250_));
  NOR2_X1    g03058(.A1(new_n3250_), .A2(new_n3244_), .ZN(new_n3251_));
  AOI22_X1   g03059(.A1(new_n3245_), .A2(\asqrt[47] ), .B1(new_n3243_), .B2(new_n3236_), .ZN(new_n3252_));
  NOR4_X1    g03060(.A1(new_n3208_), .A2(\asqrt[48] ), .A3(new_n2989_), .A4(new_n3008_), .ZN(new_n3253_));
  XOR2_X1    g03061(.A1(new_n3253_), .A2(new_n2992_), .Z(new_n3254_));
  NAND2_X1   g03062(.A1(new_n3254_), .A2(new_n1854_), .ZN(new_n3255_));
  INV_X1     g03063(.I(new_n3255_), .ZN(new_n3256_));
  OAI21_X1   g03064(.A1(new_n3252_), .A2(new_n2046_), .B(new_n3256_), .ZN(new_n3257_));
  NAND2_X1   g03065(.A1(new_n3257_), .A2(new_n3251_), .ZN(new_n3258_));
  OAI22_X1   g03066(.A1(new_n3252_), .A2(new_n2046_), .B1(new_n3250_), .B2(new_n3244_), .ZN(new_n3259_));
  NOR2_X1    g03067(.A1(new_n2996_), .A2(\asqrt[49] ), .ZN(new_n3260_));
  NAND3_X1   g03068(.A1(\asqrt[43] ), .A2(new_n3012_), .A3(new_n3260_), .ZN(new_n3261_));
  XOR2_X1    g03069(.A1(new_n3261_), .A2(new_n3000_), .Z(new_n3262_));
  NAND2_X1   g03070(.A1(new_n3262_), .A2(new_n1595_), .ZN(new_n3263_));
  AOI21_X1   g03071(.A1(new_n3259_), .A2(\asqrt[49] ), .B(new_n3263_), .ZN(new_n3264_));
  NOR2_X1    g03072(.A1(new_n3264_), .A2(new_n3258_), .ZN(new_n3265_));
  AOI22_X1   g03073(.A1(new_n3259_), .A2(\asqrt[49] ), .B1(new_n3257_), .B2(new_n3251_), .ZN(new_n3266_));
  NOR4_X1    g03074(.A1(new_n3208_), .A2(\asqrt[50] ), .A3(new_n3004_), .A4(new_n3013_), .ZN(new_n3267_));
  XOR2_X1    g03075(.A1(new_n3267_), .A2(new_n3104_), .Z(new_n3268_));
  NAND2_X1   g03076(.A1(new_n3268_), .A2(new_n1436_), .ZN(new_n3269_));
  INV_X1     g03077(.I(new_n3269_), .ZN(new_n3270_));
  OAI21_X1   g03078(.A1(new_n3266_), .A2(new_n1595_), .B(new_n3270_), .ZN(new_n3271_));
  NAND2_X1   g03079(.A1(new_n3271_), .A2(new_n3265_), .ZN(new_n3272_));
  OAI22_X1   g03080(.A1(new_n3266_), .A2(new_n1595_), .B1(new_n3264_), .B2(new_n3258_), .ZN(new_n3273_));
  NAND2_X1   g03081(.A1(new_n3108_), .A2(\asqrt[51] ), .ZN(new_n3274_));
  NOR4_X1    g03082(.A1(new_n3208_), .A2(\asqrt[51] ), .A3(new_n3016_), .A4(new_n3108_), .ZN(new_n3275_));
  XOR2_X1    g03083(.A1(new_n3275_), .A2(new_n3274_), .Z(new_n3276_));
  NAND2_X1   g03084(.A1(new_n3276_), .A2(new_n1260_), .ZN(new_n3277_));
  AOI21_X1   g03085(.A1(new_n3273_), .A2(\asqrt[51] ), .B(new_n3277_), .ZN(new_n3278_));
  NOR2_X1    g03086(.A1(new_n3278_), .A2(new_n3272_), .ZN(new_n3279_));
  AOI22_X1   g03087(.A1(new_n3273_), .A2(\asqrt[51] ), .B1(new_n3271_), .B2(new_n3265_), .ZN(new_n3280_));
  NOR4_X1    g03088(.A1(new_n3208_), .A2(\asqrt[52] ), .A3(new_n3025_), .A4(new_n3030_), .ZN(new_n3281_));
  AOI21_X1   g03089(.A1(new_n3274_), .A2(new_n3107_), .B(new_n1260_), .ZN(new_n3282_));
  NOR2_X1    g03090(.A1(new_n3281_), .A2(new_n3282_), .ZN(new_n3283_));
  NAND2_X1   g03091(.A1(new_n3283_), .A2(new_n1096_), .ZN(new_n3284_));
  INV_X1     g03092(.I(new_n3284_), .ZN(new_n3285_));
  OAI21_X1   g03093(.A1(new_n3280_), .A2(new_n1260_), .B(new_n3285_), .ZN(new_n3286_));
  NAND2_X1   g03094(.A1(new_n3286_), .A2(new_n3279_), .ZN(new_n3287_));
  OAI22_X1   g03095(.A1(new_n3280_), .A2(new_n1260_), .B1(new_n3278_), .B2(new_n3272_), .ZN(new_n3288_));
  NOR4_X1    g03096(.A1(new_n3208_), .A2(\asqrt[53] ), .A3(new_n3033_), .A4(new_n3115_), .ZN(new_n3289_));
  XOR2_X1    g03097(.A1(new_n3289_), .A2(new_n3129_), .Z(new_n3290_));
  NAND2_X1   g03098(.A1(new_n3290_), .A2(new_n970_), .ZN(new_n3291_));
  AOI21_X1   g03099(.A1(new_n3288_), .A2(\asqrt[53] ), .B(new_n3291_), .ZN(new_n3292_));
  NOR2_X1    g03100(.A1(new_n3292_), .A2(new_n3287_), .ZN(new_n3293_));
  AOI22_X1   g03101(.A1(new_n3288_), .A2(\asqrt[53] ), .B1(new_n3286_), .B2(new_n3279_), .ZN(new_n3294_));
  NOR4_X1    g03102(.A1(new_n3208_), .A2(\asqrt[54] ), .A3(new_n3040_), .A4(new_n3045_), .ZN(new_n3295_));
  XOR2_X1    g03103(.A1(new_n3295_), .A2(new_n3083_), .Z(new_n3296_));
  NAND2_X1   g03104(.A1(new_n3296_), .A2(new_n825_), .ZN(new_n3297_));
  INV_X1     g03105(.I(new_n3297_), .ZN(new_n3298_));
  OAI21_X1   g03106(.A1(new_n3294_), .A2(new_n970_), .B(new_n3298_), .ZN(new_n3299_));
  NAND2_X1   g03107(.A1(new_n3299_), .A2(new_n3293_), .ZN(new_n3300_));
  OAI22_X1   g03108(.A1(new_n3294_), .A2(new_n970_), .B1(new_n3292_), .B2(new_n3287_), .ZN(new_n3301_));
  NOR4_X1    g03109(.A1(new_n3208_), .A2(\asqrt[55] ), .A3(new_n3047_), .A4(new_n3122_), .ZN(new_n3302_));
  XOR2_X1    g03110(.A1(new_n3302_), .A2(new_n3131_), .Z(new_n3303_));
  NAND2_X1   g03111(.A1(new_n3303_), .A2(new_n724_), .ZN(new_n3304_));
  AOI21_X1   g03112(.A1(new_n3301_), .A2(\asqrt[55] ), .B(new_n3304_), .ZN(new_n3305_));
  NOR2_X1    g03113(.A1(new_n3305_), .A2(new_n3300_), .ZN(new_n3306_));
  AOI22_X1   g03114(.A1(new_n3301_), .A2(\asqrt[55] ), .B1(new_n3299_), .B2(new_n3293_), .ZN(new_n3307_));
  NOR4_X1    g03115(.A1(new_n3208_), .A2(\asqrt[56] ), .A3(new_n3053_), .A4(new_n3058_), .ZN(new_n3308_));
  XOR2_X1    g03116(.A1(new_n3308_), .A2(new_n3085_), .Z(new_n3309_));
  NAND2_X1   g03117(.A1(new_n3309_), .A2(new_n587_), .ZN(new_n3310_));
  INV_X1     g03118(.I(new_n3310_), .ZN(new_n3311_));
  OAI21_X1   g03119(.A1(new_n3307_), .A2(new_n724_), .B(new_n3311_), .ZN(new_n3312_));
  NAND2_X1   g03120(.A1(new_n3312_), .A2(new_n3306_), .ZN(new_n3313_));
  OAI22_X1   g03121(.A1(new_n3307_), .A2(new_n724_), .B1(new_n3305_), .B2(new_n3300_), .ZN(new_n3314_));
  NOR4_X1    g03122(.A1(new_n3208_), .A2(\asqrt[57] ), .A3(new_n3060_), .A4(new_n3135_), .ZN(new_n3315_));
  XOR2_X1    g03123(.A1(new_n3315_), .A2(new_n3133_), .Z(new_n3316_));
  NAND2_X1   g03124(.A1(new_n3316_), .A2(new_n504_), .ZN(new_n3317_));
  AOI21_X1   g03125(.A1(new_n3314_), .A2(\asqrt[57] ), .B(new_n3317_), .ZN(new_n3318_));
  NOR2_X1    g03126(.A1(new_n3318_), .A2(new_n3313_), .ZN(new_n3319_));
  AOI22_X1   g03127(.A1(new_n3314_), .A2(\asqrt[57] ), .B1(new_n3312_), .B2(new_n3306_), .ZN(new_n3320_));
  NOR4_X1    g03128(.A1(new_n3208_), .A2(\asqrt[58] ), .A3(new_n3066_), .A4(new_n3071_), .ZN(new_n3321_));
  XOR2_X1    g03129(.A1(new_n3321_), .A2(new_n3087_), .Z(new_n3322_));
  NAND2_X1   g03130(.A1(new_n3322_), .A2(new_n376_), .ZN(new_n3323_));
  INV_X1     g03131(.I(new_n3323_), .ZN(new_n3324_));
  OAI21_X1   g03132(.A1(new_n3320_), .A2(new_n504_), .B(new_n3324_), .ZN(new_n3325_));
  NAND2_X1   g03133(.A1(new_n3325_), .A2(new_n3319_), .ZN(new_n3326_));
  OAI22_X1   g03134(.A1(new_n3320_), .A2(new_n504_), .B1(new_n3318_), .B2(new_n3313_), .ZN(new_n3327_));
  NOR4_X1    g03135(.A1(new_n3208_), .A2(\asqrt[59] ), .A3(new_n3073_), .A4(new_n3143_), .ZN(new_n3328_));
  XOR2_X1    g03136(.A1(new_n3328_), .A2(new_n3141_), .Z(new_n3329_));
  NAND2_X1   g03137(.A1(new_n3329_), .A2(new_n275_), .ZN(new_n3330_));
  AOI21_X1   g03138(.A1(new_n3327_), .A2(\asqrt[59] ), .B(new_n3330_), .ZN(new_n3331_));
  NOR2_X1    g03139(.A1(new_n3331_), .A2(new_n3326_), .ZN(new_n3332_));
  AOI22_X1   g03140(.A1(new_n3327_), .A2(\asqrt[59] ), .B1(new_n3325_), .B2(new_n3319_), .ZN(new_n3333_));
  OAI22_X1   g03141(.A1(new_n3333_), .A2(new_n275_), .B1(new_n3331_), .B2(new_n3326_), .ZN(new_n3334_));
  NOR4_X1    g03142(.A1(new_n3208_), .A2(\asqrt[60] ), .A3(new_n3079_), .A4(new_n3165_), .ZN(new_n3335_));
  XOR2_X1    g03143(.A1(new_n3335_), .A2(new_n3089_), .Z(new_n3336_));
  NAND2_X1   g03144(.A1(new_n3336_), .A2(new_n229_), .ZN(new_n3337_));
  INV_X1     g03145(.I(new_n3337_), .ZN(new_n3338_));
  OAI21_X1   g03146(.A1(new_n3333_), .A2(new_n275_), .B(new_n3338_), .ZN(new_n3339_));
  AOI22_X1   g03147(.A1(new_n3334_), .A2(\asqrt[61] ), .B1(new_n3339_), .B2(new_n3332_), .ZN(new_n3340_));
  NOR2_X1    g03148(.A1(new_n3340_), .A2(new_n196_), .ZN(new_n3341_));
  INV_X1     g03149(.I(new_n3185_), .ZN(new_n3342_));
  AOI21_X1   g03150(.A1(new_n3199_), .A2(new_n3342_), .B(new_n3187_), .ZN(new_n3343_));
  NOR3_X1    g03151(.A1(new_n3184_), .A2(new_n3179_), .A3(new_n3183_), .ZN(new_n3344_));
  NOR2_X1    g03152(.A1(new_n3344_), .A2(new_n3343_), .ZN(new_n3345_));
  NOR3_X1    g03153(.A1(new_n3222_), .A2(new_n2671_), .A3(\asqrt[43] ), .ZN(new_n3346_));
  AOI21_X1   g03154(.A1(new_n3216_), .A2(new_n2670_), .B(new_n3208_), .ZN(new_n3347_));
  NOR4_X1    g03155(.A1(new_n3347_), .A2(new_n3346_), .A3(\asqrt[45] ), .A4(new_n3206_), .ZN(new_n3348_));
  NOR2_X1    g03156(.A1(new_n3348_), .A2(new_n3345_), .ZN(new_n3349_));
  NOR3_X1    g03157(.A1(new_n3344_), .A2(new_n3343_), .A3(new_n3206_), .ZN(new_n3350_));
  NOR3_X1    g03158(.A1(new_n3208_), .A2(new_n2939_), .A3(new_n3230_), .ZN(new_n3351_));
  AOI21_X1   g03159(.A1(\asqrt[43] ), .A2(new_n3231_), .B(new_n2940_), .ZN(new_n3352_));
  NOR3_X1    g03160(.A1(new_n3352_), .A2(new_n3351_), .A3(\asqrt[46] ), .ZN(new_n3353_));
  OAI21_X1   g03161(.A1(new_n3350_), .A2(new_n2728_), .B(new_n3353_), .ZN(new_n3354_));
  NAND2_X1   g03162(.A1(new_n3349_), .A2(new_n3354_), .ZN(new_n3355_));
  OAI22_X1   g03163(.A1(new_n3348_), .A2(new_n3345_), .B1(new_n2728_), .B2(new_n3350_), .ZN(new_n3356_));
  INV_X1     g03164(.I(new_n3242_), .ZN(new_n3357_));
  AOI21_X1   g03165(.A1(new_n3356_), .A2(\asqrt[46] ), .B(new_n3357_), .ZN(new_n3358_));
  NOR2_X1    g03166(.A1(new_n3358_), .A2(new_n3355_), .ZN(new_n3359_));
  AOI22_X1   g03167(.A1(new_n3356_), .A2(\asqrt[46] ), .B1(new_n3349_), .B2(new_n3354_), .ZN(new_n3360_));
  INV_X1     g03168(.I(new_n3249_), .ZN(new_n3361_));
  OAI21_X1   g03169(.A1(new_n3360_), .A2(new_n2253_), .B(new_n3361_), .ZN(new_n3362_));
  NAND2_X1   g03170(.A1(new_n3362_), .A2(new_n3359_), .ZN(new_n3363_));
  OAI22_X1   g03171(.A1(new_n3360_), .A2(new_n2253_), .B1(new_n3358_), .B2(new_n3355_), .ZN(new_n3364_));
  AOI21_X1   g03172(.A1(new_n3364_), .A2(\asqrt[48] ), .B(new_n3255_), .ZN(new_n3365_));
  NOR2_X1    g03173(.A1(new_n3365_), .A2(new_n3363_), .ZN(new_n3366_));
  AOI22_X1   g03174(.A1(new_n3364_), .A2(\asqrt[48] ), .B1(new_n3362_), .B2(new_n3359_), .ZN(new_n3367_));
  INV_X1     g03175(.I(new_n3263_), .ZN(new_n3368_));
  OAI21_X1   g03176(.A1(new_n3367_), .A2(new_n1854_), .B(new_n3368_), .ZN(new_n3369_));
  NAND2_X1   g03177(.A1(new_n3369_), .A2(new_n3366_), .ZN(new_n3370_));
  OAI22_X1   g03178(.A1(new_n3367_), .A2(new_n1854_), .B1(new_n3365_), .B2(new_n3363_), .ZN(new_n3371_));
  AOI21_X1   g03179(.A1(new_n3371_), .A2(\asqrt[50] ), .B(new_n3269_), .ZN(new_n3372_));
  NOR2_X1    g03180(.A1(new_n3372_), .A2(new_n3370_), .ZN(new_n3373_));
  AOI22_X1   g03181(.A1(new_n3371_), .A2(\asqrt[50] ), .B1(new_n3369_), .B2(new_n3366_), .ZN(new_n3374_));
  INV_X1     g03182(.I(new_n3277_), .ZN(new_n3375_));
  OAI21_X1   g03183(.A1(new_n3374_), .A2(new_n1436_), .B(new_n3375_), .ZN(new_n3376_));
  NAND2_X1   g03184(.A1(new_n3376_), .A2(new_n3373_), .ZN(new_n3377_));
  OAI22_X1   g03185(.A1(new_n3374_), .A2(new_n1436_), .B1(new_n3372_), .B2(new_n3370_), .ZN(new_n3378_));
  AOI21_X1   g03186(.A1(new_n3378_), .A2(\asqrt[52] ), .B(new_n3284_), .ZN(new_n3379_));
  NOR2_X1    g03187(.A1(new_n3379_), .A2(new_n3377_), .ZN(new_n3380_));
  AOI22_X1   g03188(.A1(new_n3378_), .A2(\asqrt[52] ), .B1(new_n3376_), .B2(new_n3373_), .ZN(new_n3381_));
  INV_X1     g03189(.I(new_n3291_), .ZN(new_n3382_));
  OAI21_X1   g03190(.A1(new_n3381_), .A2(new_n1096_), .B(new_n3382_), .ZN(new_n3383_));
  NAND2_X1   g03191(.A1(new_n3383_), .A2(new_n3380_), .ZN(new_n3384_));
  OAI22_X1   g03192(.A1(new_n3381_), .A2(new_n1096_), .B1(new_n3379_), .B2(new_n3377_), .ZN(new_n3385_));
  AOI21_X1   g03193(.A1(new_n3385_), .A2(\asqrt[54] ), .B(new_n3297_), .ZN(new_n3386_));
  NOR2_X1    g03194(.A1(new_n3386_), .A2(new_n3384_), .ZN(new_n3387_));
  AOI22_X1   g03195(.A1(new_n3385_), .A2(\asqrt[54] ), .B1(new_n3383_), .B2(new_n3380_), .ZN(new_n3388_));
  INV_X1     g03196(.I(new_n3304_), .ZN(new_n3389_));
  OAI21_X1   g03197(.A1(new_n3388_), .A2(new_n825_), .B(new_n3389_), .ZN(new_n3390_));
  NAND2_X1   g03198(.A1(new_n3390_), .A2(new_n3387_), .ZN(new_n3391_));
  OAI22_X1   g03199(.A1(new_n3388_), .A2(new_n825_), .B1(new_n3386_), .B2(new_n3384_), .ZN(new_n3392_));
  AOI21_X1   g03200(.A1(new_n3392_), .A2(\asqrt[56] ), .B(new_n3310_), .ZN(new_n3393_));
  NOR2_X1    g03201(.A1(new_n3393_), .A2(new_n3391_), .ZN(new_n3394_));
  AOI22_X1   g03202(.A1(new_n3392_), .A2(\asqrt[56] ), .B1(new_n3390_), .B2(new_n3387_), .ZN(new_n3395_));
  INV_X1     g03203(.I(new_n3317_), .ZN(new_n3396_));
  OAI21_X1   g03204(.A1(new_n3395_), .A2(new_n587_), .B(new_n3396_), .ZN(new_n3397_));
  NAND2_X1   g03205(.A1(new_n3397_), .A2(new_n3394_), .ZN(new_n3398_));
  OAI22_X1   g03206(.A1(new_n3395_), .A2(new_n587_), .B1(new_n3393_), .B2(new_n3391_), .ZN(new_n3399_));
  AOI21_X1   g03207(.A1(new_n3399_), .A2(\asqrt[58] ), .B(new_n3323_), .ZN(new_n3400_));
  NOR2_X1    g03208(.A1(new_n3400_), .A2(new_n3398_), .ZN(new_n3401_));
  AOI22_X1   g03209(.A1(new_n3399_), .A2(\asqrt[58] ), .B1(new_n3397_), .B2(new_n3394_), .ZN(new_n3402_));
  INV_X1     g03210(.I(new_n3330_), .ZN(new_n3403_));
  OAI21_X1   g03211(.A1(new_n3402_), .A2(new_n376_), .B(new_n3403_), .ZN(new_n3404_));
  NAND2_X1   g03212(.A1(new_n3404_), .A2(new_n3401_), .ZN(new_n3405_));
  OAI22_X1   g03213(.A1(new_n3402_), .A2(new_n376_), .B1(new_n3400_), .B2(new_n3398_), .ZN(new_n3406_));
  AOI22_X1   g03214(.A1(new_n3406_), .A2(\asqrt[60] ), .B1(new_n3404_), .B2(new_n3401_), .ZN(new_n3407_));
  AOI21_X1   g03215(.A1(new_n3406_), .A2(\asqrt[60] ), .B(new_n3337_), .ZN(new_n3408_));
  OAI22_X1   g03216(.A1(new_n3407_), .A2(new_n229_), .B1(new_n3408_), .B2(new_n3405_), .ZN(new_n3409_));
  NOR2_X1    g03217(.A1(new_n3409_), .A2(\asqrt[62] ), .ZN(new_n3410_));
  NAND3_X1   g03218(.A1(new_n3202_), .A2(new_n3096_), .A3(new_n3171_), .ZN(new_n3411_));
  NOR2_X1    g03219(.A1(new_n3211_), .A2(new_n196_), .ZN(new_n3412_));
  INV_X1     g03220(.I(new_n3196_), .ZN(new_n3413_));
  NAND3_X1   g03221(.A1(\asqrt[43] ), .A2(new_n3412_), .A3(new_n3413_), .ZN(new_n3414_));
  OAI21_X1   g03222(.A1(new_n3168_), .A2(\asqrt[62] ), .B(new_n3099_), .ZN(new_n3415_));
  OAI21_X1   g03223(.A1(\asqrt[43] ), .A2(new_n3415_), .B(new_n3412_), .ZN(new_n3416_));
  NAND2_X1   g03224(.A1(new_n3416_), .A2(new_n3414_), .ZN(new_n3417_));
  INV_X1     g03225(.I(new_n3417_), .ZN(new_n3418_));
  NOR2_X1    g03226(.A1(new_n3176_), .A2(new_n196_), .ZN(new_n3419_));
  INV_X1     g03227(.I(new_n3419_), .ZN(new_n3420_));
  NAND2_X1   g03228(.A1(new_n3314_), .A2(\asqrt[57] ), .ZN(new_n3421_));
  AOI21_X1   g03229(.A1(new_n3421_), .A2(new_n3313_), .B(new_n504_), .ZN(new_n3422_));
  OAI21_X1   g03230(.A1(new_n3319_), .A2(new_n3422_), .B(\asqrt[59] ), .ZN(new_n3423_));
  AOI21_X1   g03231(.A1(new_n3326_), .A2(new_n3423_), .B(new_n275_), .ZN(new_n3424_));
  OAI21_X1   g03232(.A1(new_n3332_), .A2(new_n3424_), .B(\asqrt[61] ), .ZN(new_n3425_));
  NOR2_X1    g03233(.A1(new_n3177_), .A2(\asqrt[62] ), .ZN(new_n3426_));
  INV_X1     g03234(.I(new_n3426_), .ZN(new_n3427_));
  NAND3_X1   g03235(.A1(new_n3339_), .A2(new_n3332_), .A3(new_n3427_), .ZN(new_n3428_));
  OAI21_X1   g03236(.A1(new_n3428_), .A2(new_n3425_), .B(new_n3420_), .ZN(new_n3429_));
  NAND3_X1   g03237(.A1(new_n3208_), .A2(new_n3164_), .A3(new_n3212_), .ZN(new_n3430_));
  AOI21_X1   g03238(.A1(new_n3430_), .A2(new_n3155_), .B(\asqrt[63] ), .ZN(new_n3431_));
  INV_X1     g03239(.I(new_n3431_), .ZN(new_n3432_));
  OAI21_X1   g03240(.A1(new_n3429_), .A2(new_n3432_), .B(new_n3418_), .ZN(new_n3433_));
  NOR4_X1    g03241(.A1(new_n3409_), .A2(\asqrt[62] ), .A3(new_n3417_), .A4(new_n3176_), .ZN(new_n3434_));
  AOI21_X1   g03242(.A1(new_n3164_), .A2(new_n3190_), .B(new_n3208_), .ZN(new_n3435_));
  XOR2_X1    g03243(.A1(new_n3190_), .A2(\asqrt[63] ), .Z(new_n3436_));
  NOR2_X1    g03244(.A1(new_n3435_), .A2(new_n3436_), .ZN(new_n3437_));
  NAND2_X1   g03245(.A1(new_n3434_), .A2(new_n3437_), .ZN(new_n3438_));
  NOR3_X1    g03246(.A1(new_n3438_), .A2(new_n3411_), .A3(new_n3433_), .ZN(\asqrt[42] ));
  NAND4_X1   g03247(.A1(\asqrt[42] ), .A2(new_n3177_), .A3(new_n3341_), .A4(new_n3410_), .ZN(new_n3440_));
  OAI21_X1   g03248(.A1(new_n3409_), .A2(\asqrt[62] ), .B(new_n3176_), .ZN(new_n3441_));
  OAI21_X1   g03249(.A1(\asqrt[42] ), .A2(new_n3441_), .B(new_n3341_), .ZN(new_n3442_));
  NAND2_X1   g03250(.A1(new_n3440_), .A2(new_n3442_), .ZN(new_n3443_));
  INV_X1     g03251(.I(new_n3443_), .ZN(new_n3444_));
  NAND2_X1   g03252(.A1(new_n3399_), .A2(\asqrt[58] ), .ZN(new_n3445_));
  AOI21_X1   g03253(.A1(new_n3445_), .A2(new_n3398_), .B(new_n376_), .ZN(new_n3446_));
  OAI21_X1   g03254(.A1(new_n3401_), .A2(new_n3446_), .B(\asqrt[60] ), .ZN(new_n3447_));
  AOI21_X1   g03255(.A1(new_n3405_), .A2(new_n3447_), .B(new_n229_), .ZN(new_n3448_));
  NOR3_X1    g03256(.A1(new_n3334_), .A2(\asqrt[61] ), .A3(new_n3336_), .ZN(new_n3449_));
  NAND2_X1   g03257(.A1(\asqrt[42] ), .A2(new_n3449_), .ZN(new_n3450_));
  XOR2_X1    g03258(.A1(new_n3450_), .A2(new_n3448_), .Z(new_n3451_));
  NOR2_X1    g03259(.A1(new_n3451_), .A2(new_n196_), .ZN(new_n3452_));
  INV_X1     g03260(.I(new_n3452_), .ZN(new_n3453_));
  INV_X1     g03261(.I(\a[84] ), .ZN(new_n3454_));
  NOR2_X1    g03262(.A1(\a[82] ), .A2(\a[83] ), .ZN(new_n3455_));
  INV_X1     g03263(.I(new_n3455_), .ZN(new_n3456_));
  NOR3_X1    g03264(.A1(new_n3214_), .A2(new_n3454_), .A3(new_n3456_), .ZN(new_n3457_));
  NAND2_X1   g03265(.A1(new_n3220_), .A2(new_n3457_), .ZN(new_n3458_));
  XOR2_X1    g03266(.A1(new_n3458_), .A2(\a[85] ), .Z(new_n3459_));
  INV_X1     g03267(.I(\a[85] ), .ZN(new_n3460_));
  NOR4_X1    g03268(.A1(new_n3438_), .A2(new_n3460_), .A3(new_n3411_), .A4(new_n3433_), .ZN(new_n3461_));
  NOR2_X1    g03269(.A1(new_n3460_), .A2(\a[84] ), .ZN(new_n3462_));
  OAI21_X1   g03270(.A1(new_n3461_), .A2(new_n3462_), .B(new_n3459_), .ZN(new_n3463_));
  INV_X1     g03271(.I(new_n3459_), .ZN(new_n3464_));
  INV_X1     g03272(.I(new_n3411_), .ZN(new_n3465_));
  NOR3_X1    g03273(.A1(new_n3408_), .A2(new_n3405_), .A3(new_n3426_), .ZN(new_n3466_));
  AOI21_X1   g03274(.A1(new_n3466_), .A2(new_n3448_), .B(new_n3419_), .ZN(new_n3467_));
  AOI21_X1   g03275(.A1(new_n3467_), .A2(new_n3431_), .B(new_n3417_), .ZN(new_n3468_));
  NAND4_X1   g03276(.A1(new_n3340_), .A2(new_n196_), .A3(new_n3418_), .A4(new_n3177_), .ZN(new_n3469_));
  INV_X1     g03277(.I(new_n3437_), .ZN(new_n3470_));
  NOR2_X1    g03278(.A1(new_n3469_), .A2(new_n3470_), .ZN(new_n3471_));
  NAND4_X1   g03279(.A1(new_n3471_), .A2(\a[85] ), .A3(new_n3468_), .A4(new_n3465_), .ZN(new_n3472_));
  NAND3_X1   g03280(.A1(new_n3472_), .A2(\a[84] ), .A3(new_n3464_), .ZN(new_n3473_));
  NAND2_X1   g03281(.A1(new_n3463_), .A2(new_n3473_), .ZN(new_n3474_));
  NOR2_X1    g03282(.A1(new_n3438_), .A2(new_n3433_), .ZN(new_n3475_));
  NOR4_X1    g03283(.A1(new_n3170_), .A2(new_n3164_), .A3(new_n3210_), .A4(new_n3171_), .ZN(new_n3476_));
  NAND2_X1   g03284(.A1(\asqrt[43] ), .A2(\a[84] ), .ZN(new_n3477_));
  XOR2_X1    g03285(.A1(new_n3477_), .A2(new_n3476_), .Z(new_n3478_));
  NOR2_X1    g03286(.A1(new_n3478_), .A2(new_n3456_), .ZN(new_n3479_));
  INV_X1     g03287(.I(new_n3479_), .ZN(new_n3480_));
  NAND3_X1   g03288(.A1(new_n3471_), .A2(new_n3465_), .A3(new_n3468_), .ZN(new_n3481_));
  NOR2_X1    g03289(.A1(new_n3437_), .A2(new_n3465_), .ZN(new_n3482_));
  NAND2_X1   g03290(.A1(new_n3482_), .A2(\asqrt[43] ), .ZN(new_n3483_));
  INV_X1     g03291(.I(new_n3483_), .ZN(new_n3484_));
  NAND3_X1   g03292(.A1(new_n3433_), .A2(new_n3469_), .A3(new_n3484_), .ZN(new_n3485_));
  NAND2_X1   g03293(.A1(new_n3485_), .A2(new_n3179_), .ZN(new_n3486_));
  NAND3_X1   g03294(.A1(new_n3486_), .A2(new_n3180_), .A3(new_n3481_), .ZN(new_n3487_));
  NOR3_X1    g03295(.A1(new_n3468_), .A2(new_n3434_), .A3(new_n3483_), .ZN(new_n3488_));
  OAI21_X1   g03296(.A1(new_n3488_), .A2(\a[86] ), .B(new_n3180_), .ZN(new_n3489_));
  NAND2_X1   g03297(.A1(new_n3489_), .A2(\asqrt[42] ), .ZN(new_n3490_));
  NAND4_X1   g03298(.A1(new_n3490_), .A2(new_n2941_), .A3(new_n3487_), .A4(new_n3480_), .ZN(new_n3491_));
  NAND2_X1   g03299(.A1(new_n3491_), .A2(new_n3474_), .ZN(new_n3492_));
  NAND3_X1   g03300(.A1(new_n3463_), .A2(new_n3473_), .A3(new_n3480_), .ZN(new_n3493_));
  NAND2_X1   g03301(.A1(\asqrt[43] ), .A2(new_n3179_), .ZN(new_n3494_));
  AOI22_X1   g03302(.A1(new_n3494_), .A2(new_n3178_), .B1(new_n3179_), .B2(new_n3184_), .ZN(new_n3495_));
  OAI21_X1   g03303(.A1(new_n3208_), .A2(new_n3179_), .B(new_n3182_), .ZN(new_n3496_));
  NOR2_X1    g03304(.A1(new_n3495_), .A2(new_n3496_), .ZN(new_n3497_));
  NAND3_X1   g03305(.A1(\asqrt[42] ), .A2(new_n3207_), .A3(new_n3497_), .ZN(new_n3498_));
  INV_X1     g03306(.I(new_n3497_), .ZN(new_n3499_));
  OAI21_X1   g03307(.A1(new_n3481_), .A2(new_n3499_), .B(new_n3206_), .ZN(new_n3500_));
  NAND3_X1   g03308(.A1(new_n3498_), .A2(new_n3500_), .A3(new_n2728_), .ZN(new_n3501_));
  AOI21_X1   g03309(.A1(new_n3493_), .A2(\asqrt[44] ), .B(new_n3501_), .ZN(new_n3502_));
  NOR2_X1    g03310(.A1(new_n3492_), .A2(new_n3502_), .ZN(new_n3503_));
  NAND2_X1   g03311(.A1(new_n3493_), .A2(\asqrt[44] ), .ZN(new_n3504_));
  AOI21_X1   g03312(.A1(new_n3492_), .A2(new_n3504_), .B(new_n2728_), .ZN(new_n3505_));
  NOR2_X1    g03313(.A1(new_n3347_), .A2(new_n3346_), .ZN(new_n3506_));
  NOR4_X1    g03314(.A1(new_n3481_), .A2(\asqrt[45] ), .A3(new_n3506_), .A4(new_n3226_), .ZN(new_n3507_));
  AOI21_X1   g03315(.A1(new_n3345_), .A2(new_n3207_), .B(new_n2728_), .ZN(new_n3508_));
  NOR2_X1    g03316(.A1(new_n3507_), .A2(new_n3508_), .ZN(new_n3509_));
  NAND2_X1   g03317(.A1(new_n3509_), .A2(new_n2488_), .ZN(new_n3510_));
  OAI21_X1   g03318(.A1(new_n3505_), .A2(new_n3510_), .B(new_n3503_), .ZN(new_n3511_));
  AOI22_X1   g03319(.A1(new_n3491_), .A2(new_n3474_), .B1(\asqrt[44] ), .B2(new_n3493_), .ZN(new_n3512_));
  OAI22_X1   g03320(.A1(new_n3512_), .A2(new_n2728_), .B1(new_n3492_), .B2(new_n3502_), .ZN(new_n3513_));
  NOR2_X1    g03321(.A1(new_n3237_), .A2(new_n2488_), .ZN(new_n3514_));
  NAND2_X1   g03322(.A1(new_n3232_), .A2(new_n3233_), .ZN(new_n3515_));
  NAND4_X1   g03323(.A1(\asqrt[42] ), .A2(new_n2488_), .A3(new_n3515_), .A4(new_n3237_), .ZN(new_n3516_));
  XOR2_X1    g03324(.A1(new_n3516_), .A2(new_n3514_), .Z(new_n3517_));
  NAND2_X1   g03325(.A1(new_n3517_), .A2(new_n2253_), .ZN(new_n3518_));
  AOI21_X1   g03326(.A1(new_n3513_), .A2(\asqrt[46] ), .B(new_n3518_), .ZN(new_n3519_));
  OAI21_X1   g03327(.A1(new_n3505_), .A2(new_n3503_), .B(\asqrt[46] ), .ZN(new_n3520_));
  AOI21_X1   g03328(.A1(new_n3511_), .A2(new_n3520_), .B(new_n2253_), .ZN(new_n3521_));
  NAND2_X1   g03329(.A1(new_n3245_), .A2(\asqrt[47] ), .ZN(new_n3522_));
  OAI21_X1   g03330(.A1(new_n3240_), .A2(new_n3241_), .B(new_n2253_), .ZN(new_n3523_));
  NOR3_X1    g03331(.A1(new_n3481_), .A2(new_n3245_), .A3(new_n3523_), .ZN(new_n3524_));
  XOR2_X1    g03332(.A1(new_n3524_), .A2(new_n3522_), .Z(new_n3525_));
  NAND2_X1   g03333(.A1(new_n3525_), .A2(new_n2046_), .ZN(new_n3526_));
  NOR2_X1    g03334(.A1(new_n3521_), .A2(new_n3526_), .ZN(new_n3527_));
  NOR3_X1    g03335(.A1(new_n3527_), .A2(new_n3511_), .A3(new_n3519_), .ZN(new_n3528_));
  INV_X1     g03336(.I(new_n3518_), .ZN(new_n3529_));
  AOI21_X1   g03337(.A1(new_n3520_), .A2(new_n3529_), .B(new_n3511_), .ZN(new_n3530_));
  OAI21_X1   g03338(.A1(new_n3530_), .A2(new_n3521_), .B(\asqrt[48] ), .ZN(new_n3531_));
  NAND2_X1   g03339(.A1(new_n3364_), .A2(\asqrt[48] ), .ZN(new_n3532_));
  NOR4_X1    g03340(.A1(new_n3481_), .A2(\asqrt[48] ), .A3(new_n3248_), .A4(new_n3364_), .ZN(new_n3533_));
  XOR2_X1    g03341(.A1(new_n3533_), .A2(new_n3532_), .Z(new_n3534_));
  NAND2_X1   g03342(.A1(new_n3534_), .A2(new_n1854_), .ZN(new_n3535_));
  INV_X1     g03343(.I(new_n3535_), .ZN(new_n3536_));
  NAND2_X1   g03344(.A1(new_n3531_), .A2(new_n3536_), .ZN(new_n3537_));
  NAND2_X1   g03345(.A1(new_n3537_), .A2(new_n3528_), .ZN(new_n3538_));
  OAI21_X1   g03346(.A1(new_n3521_), .A2(new_n3526_), .B(new_n3530_), .ZN(new_n3539_));
  NAND2_X1   g03347(.A1(new_n3539_), .A2(new_n3531_), .ZN(new_n3540_));
  NAND2_X1   g03348(.A1(new_n3259_), .A2(\asqrt[49] ), .ZN(new_n3541_));
  NOR4_X1    g03349(.A1(new_n3481_), .A2(\asqrt[49] ), .A3(new_n3254_), .A4(new_n3259_), .ZN(new_n3542_));
  XOR2_X1    g03350(.A1(new_n3542_), .A2(new_n3541_), .Z(new_n3543_));
  NAND2_X1   g03351(.A1(new_n3543_), .A2(new_n1595_), .ZN(new_n3544_));
  AOI21_X1   g03352(.A1(new_n3540_), .A2(\asqrt[49] ), .B(new_n3544_), .ZN(new_n3545_));
  NOR2_X1    g03353(.A1(new_n3545_), .A2(new_n3538_), .ZN(new_n3546_));
  AOI22_X1   g03354(.A1(new_n3540_), .A2(\asqrt[49] ), .B1(new_n3537_), .B2(new_n3528_), .ZN(new_n3547_));
  NAND2_X1   g03355(.A1(new_n3371_), .A2(\asqrt[50] ), .ZN(new_n3548_));
  NOR4_X1    g03356(.A1(new_n3481_), .A2(\asqrt[50] ), .A3(new_n3262_), .A4(new_n3371_), .ZN(new_n3549_));
  XOR2_X1    g03357(.A1(new_n3549_), .A2(new_n3548_), .Z(new_n3550_));
  NAND2_X1   g03358(.A1(new_n3550_), .A2(new_n1436_), .ZN(new_n3551_));
  INV_X1     g03359(.I(new_n3551_), .ZN(new_n3552_));
  OAI21_X1   g03360(.A1(new_n3547_), .A2(new_n1595_), .B(new_n3552_), .ZN(new_n3553_));
  NAND2_X1   g03361(.A1(new_n3553_), .A2(new_n3546_), .ZN(new_n3554_));
  OAI22_X1   g03362(.A1(new_n3547_), .A2(new_n1595_), .B1(new_n3545_), .B2(new_n3538_), .ZN(new_n3555_));
  NAND2_X1   g03363(.A1(new_n3273_), .A2(\asqrt[51] ), .ZN(new_n3556_));
  NOR4_X1    g03364(.A1(new_n3481_), .A2(\asqrt[51] ), .A3(new_n3268_), .A4(new_n3273_), .ZN(new_n3557_));
  XOR2_X1    g03365(.A1(new_n3557_), .A2(new_n3556_), .Z(new_n3558_));
  NAND2_X1   g03366(.A1(new_n3558_), .A2(new_n1260_), .ZN(new_n3559_));
  AOI21_X1   g03367(.A1(new_n3555_), .A2(\asqrt[51] ), .B(new_n3559_), .ZN(new_n3560_));
  NOR2_X1    g03368(.A1(new_n3560_), .A2(new_n3554_), .ZN(new_n3561_));
  AOI22_X1   g03369(.A1(new_n3555_), .A2(\asqrt[51] ), .B1(new_n3553_), .B2(new_n3546_), .ZN(new_n3562_));
  NAND2_X1   g03370(.A1(new_n3378_), .A2(\asqrt[52] ), .ZN(new_n3563_));
  NOR4_X1    g03371(.A1(new_n3481_), .A2(\asqrt[52] ), .A3(new_n3276_), .A4(new_n3378_), .ZN(new_n3564_));
  XOR2_X1    g03372(.A1(new_n3564_), .A2(new_n3563_), .Z(new_n3565_));
  NAND2_X1   g03373(.A1(new_n3565_), .A2(new_n1096_), .ZN(new_n3566_));
  INV_X1     g03374(.I(new_n3566_), .ZN(new_n3567_));
  OAI21_X1   g03375(.A1(new_n3562_), .A2(new_n1260_), .B(new_n3567_), .ZN(new_n3568_));
  NAND2_X1   g03376(.A1(new_n3568_), .A2(new_n3561_), .ZN(new_n3569_));
  OAI22_X1   g03377(.A1(new_n3562_), .A2(new_n1260_), .B1(new_n3560_), .B2(new_n3554_), .ZN(new_n3570_));
  NAND2_X1   g03378(.A1(new_n3288_), .A2(\asqrt[53] ), .ZN(new_n3571_));
  NOR4_X1    g03379(.A1(new_n3481_), .A2(\asqrt[53] ), .A3(new_n3283_), .A4(new_n3288_), .ZN(new_n3572_));
  XOR2_X1    g03380(.A1(new_n3572_), .A2(new_n3571_), .Z(new_n3573_));
  NAND2_X1   g03381(.A1(new_n3573_), .A2(new_n970_), .ZN(new_n3574_));
  AOI21_X1   g03382(.A1(new_n3570_), .A2(\asqrt[53] ), .B(new_n3574_), .ZN(new_n3575_));
  NOR2_X1    g03383(.A1(new_n3575_), .A2(new_n3569_), .ZN(new_n3576_));
  AOI22_X1   g03384(.A1(new_n3570_), .A2(\asqrt[53] ), .B1(new_n3568_), .B2(new_n3561_), .ZN(new_n3577_));
  NAND2_X1   g03385(.A1(new_n3385_), .A2(\asqrt[54] ), .ZN(new_n3578_));
  NOR4_X1    g03386(.A1(new_n3481_), .A2(\asqrt[54] ), .A3(new_n3290_), .A4(new_n3385_), .ZN(new_n3579_));
  XOR2_X1    g03387(.A1(new_n3579_), .A2(new_n3578_), .Z(new_n3580_));
  NAND2_X1   g03388(.A1(new_n3580_), .A2(new_n825_), .ZN(new_n3581_));
  INV_X1     g03389(.I(new_n3581_), .ZN(new_n3582_));
  OAI21_X1   g03390(.A1(new_n3577_), .A2(new_n970_), .B(new_n3582_), .ZN(new_n3583_));
  NAND2_X1   g03391(.A1(new_n3583_), .A2(new_n3576_), .ZN(new_n3584_));
  OAI22_X1   g03392(.A1(new_n3577_), .A2(new_n970_), .B1(new_n3575_), .B2(new_n3569_), .ZN(new_n3585_));
  NAND2_X1   g03393(.A1(new_n3301_), .A2(\asqrt[55] ), .ZN(new_n3586_));
  NOR4_X1    g03394(.A1(new_n3481_), .A2(\asqrt[55] ), .A3(new_n3296_), .A4(new_n3301_), .ZN(new_n3587_));
  XOR2_X1    g03395(.A1(new_n3587_), .A2(new_n3586_), .Z(new_n3588_));
  NAND2_X1   g03396(.A1(new_n3588_), .A2(new_n724_), .ZN(new_n3589_));
  AOI21_X1   g03397(.A1(new_n3585_), .A2(\asqrt[55] ), .B(new_n3589_), .ZN(new_n3590_));
  NOR2_X1    g03398(.A1(new_n3590_), .A2(new_n3584_), .ZN(new_n3591_));
  AOI22_X1   g03399(.A1(new_n3585_), .A2(\asqrt[55] ), .B1(new_n3583_), .B2(new_n3576_), .ZN(new_n3592_));
  NAND2_X1   g03400(.A1(new_n3392_), .A2(\asqrt[56] ), .ZN(new_n3593_));
  NOR4_X1    g03401(.A1(new_n3481_), .A2(\asqrt[56] ), .A3(new_n3303_), .A4(new_n3392_), .ZN(new_n3594_));
  XOR2_X1    g03402(.A1(new_n3594_), .A2(new_n3593_), .Z(new_n3595_));
  NAND2_X1   g03403(.A1(new_n3595_), .A2(new_n587_), .ZN(new_n3596_));
  INV_X1     g03404(.I(new_n3596_), .ZN(new_n3597_));
  OAI21_X1   g03405(.A1(new_n3592_), .A2(new_n724_), .B(new_n3597_), .ZN(new_n3598_));
  NAND2_X1   g03406(.A1(new_n3598_), .A2(new_n3591_), .ZN(new_n3599_));
  NOR2_X1    g03407(.A1(new_n3592_), .A2(new_n724_), .ZN(new_n3600_));
  OAI21_X1   g03408(.A1(new_n3600_), .A2(new_n3591_), .B(\asqrt[57] ), .ZN(new_n3601_));
  NOR4_X1    g03409(.A1(new_n3481_), .A2(\asqrt[57] ), .A3(new_n3309_), .A4(new_n3314_), .ZN(new_n3602_));
  XOR2_X1    g03410(.A1(new_n3602_), .A2(new_n3421_), .Z(new_n3603_));
  NAND2_X1   g03411(.A1(new_n3603_), .A2(new_n504_), .ZN(new_n3604_));
  INV_X1     g03412(.I(new_n3604_), .ZN(new_n3605_));
  AOI21_X1   g03413(.A1(new_n3601_), .A2(new_n3605_), .B(new_n3599_), .ZN(new_n3606_));
  OAI22_X1   g03414(.A1(new_n3592_), .A2(new_n724_), .B1(new_n3590_), .B2(new_n3584_), .ZN(new_n3607_));
  AOI22_X1   g03415(.A1(new_n3607_), .A2(\asqrt[57] ), .B1(new_n3598_), .B2(new_n3591_), .ZN(new_n3608_));
  NOR4_X1    g03416(.A1(new_n3481_), .A2(\asqrt[58] ), .A3(new_n3316_), .A4(new_n3399_), .ZN(new_n3609_));
  XOR2_X1    g03417(.A1(new_n3609_), .A2(new_n3445_), .Z(new_n3610_));
  NAND2_X1   g03418(.A1(new_n3610_), .A2(new_n376_), .ZN(new_n3611_));
  INV_X1     g03419(.I(new_n3611_), .ZN(new_n3612_));
  OAI21_X1   g03420(.A1(new_n3608_), .A2(new_n504_), .B(new_n3612_), .ZN(new_n3613_));
  NAND2_X1   g03421(.A1(new_n3613_), .A2(new_n3606_), .ZN(new_n3614_));
  AOI21_X1   g03422(.A1(new_n3601_), .A2(new_n3599_), .B(new_n504_), .ZN(new_n3615_));
  OAI21_X1   g03423(.A1(new_n3606_), .A2(new_n3615_), .B(\asqrt[59] ), .ZN(new_n3616_));
  NOR4_X1    g03424(.A1(new_n3481_), .A2(\asqrt[59] ), .A3(new_n3322_), .A4(new_n3327_), .ZN(new_n3617_));
  XOR2_X1    g03425(.A1(new_n3617_), .A2(new_n3423_), .Z(new_n3618_));
  AND2_X2    g03426(.A1(new_n3618_), .A2(new_n275_), .Z(new_n3619_));
  AOI21_X1   g03427(.A1(new_n3616_), .A2(new_n3619_), .B(new_n3614_), .ZN(new_n3620_));
  INV_X1     g03428(.I(new_n3510_), .ZN(new_n3621_));
  OAI21_X1   g03429(.A1(new_n3512_), .A2(new_n2728_), .B(new_n3621_), .ZN(new_n3622_));
  AOI22_X1   g03430(.A1(new_n3513_), .A2(\asqrt[46] ), .B1(new_n3622_), .B2(new_n3503_), .ZN(new_n3623_));
  OAI22_X1   g03431(.A1(new_n3623_), .A2(new_n2253_), .B1(new_n3519_), .B2(new_n3511_), .ZN(new_n3624_));
  AOI21_X1   g03432(.A1(new_n3624_), .A2(\asqrt[48] ), .B(new_n3535_), .ZN(new_n3625_));
  NOR2_X1    g03433(.A1(new_n3625_), .A2(new_n3539_), .ZN(new_n3626_));
  INV_X1     g03434(.I(new_n3526_), .ZN(new_n3627_));
  OAI21_X1   g03435(.A1(new_n3623_), .A2(new_n2253_), .B(new_n3627_), .ZN(new_n3628_));
  AOI22_X1   g03436(.A1(new_n3624_), .A2(\asqrt[48] ), .B1(new_n3628_), .B2(new_n3530_), .ZN(new_n3629_));
  INV_X1     g03437(.I(new_n3544_), .ZN(new_n3630_));
  OAI21_X1   g03438(.A1(new_n3629_), .A2(new_n1854_), .B(new_n3630_), .ZN(new_n3631_));
  NAND2_X1   g03439(.A1(new_n3631_), .A2(new_n3626_), .ZN(new_n3632_));
  OAI22_X1   g03440(.A1(new_n3629_), .A2(new_n1854_), .B1(new_n3625_), .B2(new_n3539_), .ZN(new_n3633_));
  AOI21_X1   g03441(.A1(new_n3633_), .A2(\asqrt[50] ), .B(new_n3551_), .ZN(new_n3634_));
  NOR2_X1    g03442(.A1(new_n3634_), .A2(new_n3632_), .ZN(new_n3635_));
  AOI22_X1   g03443(.A1(new_n3633_), .A2(\asqrt[50] ), .B1(new_n3631_), .B2(new_n3626_), .ZN(new_n3636_));
  INV_X1     g03444(.I(new_n3559_), .ZN(new_n3637_));
  OAI21_X1   g03445(.A1(new_n3636_), .A2(new_n1436_), .B(new_n3637_), .ZN(new_n3638_));
  NAND2_X1   g03446(.A1(new_n3638_), .A2(new_n3635_), .ZN(new_n3639_));
  OAI22_X1   g03447(.A1(new_n3636_), .A2(new_n1436_), .B1(new_n3634_), .B2(new_n3632_), .ZN(new_n3640_));
  AOI21_X1   g03448(.A1(new_n3640_), .A2(\asqrt[52] ), .B(new_n3566_), .ZN(new_n3641_));
  NOR2_X1    g03449(.A1(new_n3641_), .A2(new_n3639_), .ZN(new_n3642_));
  AOI22_X1   g03450(.A1(new_n3640_), .A2(\asqrt[52] ), .B1(new_n3638_), .B2(new_n3635_), .ZN(new_n3643_));
  INV_X1     g03451(.I(new_n3574_), .ZN(new_n3644_));
  OAI21_X1   g03452(.A1(new_n3643_), .A2(new_n1096_), .B(new_n3644_), .ZN(new_n3645_));
  NAND2_X1   g03453(.A1(new_n3645_), .A2(new_n3642_), .ZN(new_n3646_));
  OAI22_X1   g03454(.A1(new_n3643_), .A2(new_n1096_), .B1(new_n3641_), .B2(new_n3639_), .ZN(new_n3647_));
  AOI21_X1   g03455(.A1(new_n3647_), .A2(\asqrt[54] ), .B(new_n3581_), .ZN(new_n3648_));
  NOR2_X1    g03456(.A1(new_n3648_), .A2(new_n3646_), .ZN(new_n3649_));
  AOI22_X1   g03457(.A1(new_n3647_), .A2(\asqrt[54] ), .B1(new_n3645_), .B2(new_n3642_), .ZN(new_n3650_));
  INV_X1     g03458(.I(new_n3589_), .ZN(new_n3651_));
  OAI21_X1   g03459(.A1(new_n3650_), .A2(new_n825_), .B(new_n3651_), .ZN(new_n3652_));
  NAND2_X1   g03460(.A1(new_n3652_), .A2(new_n3649_), .ZN(new_n3653_));
  OAI22_X1   g03461(.A1(new_n3650_), .A2(new_n825_), .B1(new_n3648_), .B2(new_n3646_), .ZN(new_n3654_));
  AOI21_X1   g03462(.A1(new_n3654_), .A2(\asqrt[56] ), .B(new_n3596_), .ZN(new_n3655_));
  NOR2_X1    g03463(.A1(new_n3655_), .A2(new_n3653_), .ZN(new_n3656_));
  AOI22_X1   g03464(.A1(new_n3654_), .A2(\asqrt[56] ), .B1(new_n3652_), .B2(new_n3649_), .ZN(new_n3657_));
  OAI21_X1   g03465(.A1(new_n3657_), .A2(new_n587_), .B(new_n3605_), .ZN(new_n3658_));
  NAND2_X1   g03466(.A1(new_n3658_), .A2(new_n3656_), .ZN(new_n3659_));
  NAND2_X1   g03467(.A1(new_n3647_), .A2(\asqrt[54] ), .ZN(new_n3660_));
  AOI21_X1   g03468(.A1(new_n3660_), .A2(new_n3646_), .B(new_n825_), .ZN(new_n3661_));
  OAI21_X1   g03469(.A1(new_n3649_), .A2(new_n3661_), .B(\asqrt[56] ), .ZN(new_n3662_));
  AOI21_X1   g03470(.A1(new_n3653_), .A2(new_n3662_), .B(new_n587_), .ZN(new_n3663_));
  OAI21_X1   g03471(.A1(new_n3656_), .A2(new_n3663_), .B(\asqrt[58] ), .ZN(new_n3664_));
  NAND2_X1   g03472(.A1(new_n3659_), .A2(new_n3664_), .ZN(new_n3665_));
  AOI22_X1   g03473(.A1(new_n3665_), .A2(\asqrt[59] ), .B1(new_n3613_), .B2(new_n3606_), .ZN(new_n3666_));
  NOR4_X1    g03474(.A1(new_n3481_), .A2(\asqrt[60] ), .A3(new_n3329_), .A4(new_n3406_), .ZN(new_n3667_));
  XOR2_X1    g03475(.A1(new_n3667_), .A2(new_n3447_), .Z(new_n3668_));
  NAND2_X1   g03476(.A1(new_n3668_), .A2(new_n229_), .ZN(new_n3669_));
  INV_X1     g03477(.I(new_n3669_), .ZN(new_n3670_));
  OAI21_X1   g03478(.A1(new_n3666_), .A2(new_n275_), .B(new_n3670_), .ZN(new_n3671_));
  OAI22_X1   g03479(.A1(new_n3657_), .A2(new_n587_), .B1(new_n3655_), .B2(new_n3653_), .ZN(new_n3672_));
  AOI21_X1   g03480(.A1(new_n3672_), .A2(\asqrt[58] ), .B(new_n3611_), .ZN(new_n3673_));
  NOR2_X1    g03481(.A1(new_n3673_), .A2(new_n3659_), .ZN(new_n3674_));
  AOI22_X1   g03482(.A1(new_n3672_), .A2(\asqrt[58] ), .B1(new_n3658_), .B2(new_n3656_), .ZN(new_n3675_));
  OAI21_X1   g03483(.A1(new_n3675_), .A2(new_n376_), .B(new_n3619_), .ZN(new_n3676_));
  NAND2_X1   g03484(.A1(new_n3676_), .A2(new_n3674_), .ZN(new_n3677_));
  AOI21_X1   g03485(.A1(new_n3659_), .A2(new_n3664_), .B(new_n376_), .ZN(new_n3678_));
  OAI21_X1   g03486(.A1(new_n3674_), .A2(new_n3678_), .B(\asqrt[60] ), .ZN(new_n3679_));
  AOI21_X1   g03487(.A1(new_n3677_), .A2(new_n3679_), .B(new_n229_), .ZN(new_n3680_));
  INV_X1     g03488(.I(new_n3451_), .ZN(new_n3681_));
  NOR2_X1    g03489(.A1(new_n3681_), .A2(\asqrt[62] ), .ZN(new_n3682_));
  INV_X1     g03490(.I(new_n3682_), .ZN(new_n3683_));
  NAND4_X1   g03491(.A1(new_n3680_), .A2(new_n3620_), .A3(new_n3671_), .A4(new_n3683_), .ZN(new_n3684_));
  NAND3_X1   g03492(.A1(new_n3481_), .A2(new_n3417_), .A3(new_n3469_), .ZN(new_n3685_));
  AOI21_X1   g03493(.A1(new_n3685_), .A2(new_n3429_), .B(\asqrt[63] ), .ZN(new_n3686_));
  NAND3_X1   g03494(.A1(new_n3684_), .A2(new_n3453_), .A3(new_n3686_), .ZN(new_n3687_));
  OAI22_X1   g03495(.A1(new_n3675_), .A2(new_n376_), .B1(new_n3673_), .B2(new_n3659_), .ZN(new_n3688_));
  AOI21_X1   g03496(.A1(new_n3688_), .A2(\asqrt[60] ), .B(new_n3669_), .ZN(new_n3689_));
  AOI22_X1   g03497(.A1(new_n3688_), .A2(\asqrt[60] ), .B1(new_n3676_), .B2(new_n3674_), .ZN(new_n3690_));
  OAI22_X1   g03498(.A1(new_n3690_), .A2(new_n229_), .B1(new_n3689_), .B2(new_n3677_), .ZN(new_n3691_));
  NOR4_X1    g03499(.A1(new_n3691_), .A2(\asqrt[62] ), .A3(new_n3443_), .A4(new_n3451_), .ZN(new_n3692_));
  AOI21_X1   g03500(.A1(new_n3444_), .A2(new_n3687_), .B(new_n3692_), .ZN(new_n3693_));
  INV_X1     g03501(.I(\a[80] ), .ZN(new_n3694_));
  OAI21_X1   g03502(.A1(new_n3418_), .A2(new_n3429_), .B(\asqrt[42] ), .ZN(new_n3695_));
  XOR2_X1    g03503(.A1(new_n3429_), .A2(\asqrt[63] ), .Z(new_n3696_));
  NAND2_X1   g03504(.A1(new_n3695_), .A2(new_n3696_), .ZN(new_n3697_));
  INV_X1     g03505(.I(new_n3697_), .ZN(new_n3698_));
  NAND3_X1   g03506(.A1(new_n3475_), .A2(new_n3411_), .A3(new_n3418_), .ZN(new_n3699_));
  INV_X1     g03507(.I(new_n3699_), .ZN(new_n3700_));
  NOR2_X1    g03508(.A1(new_n3698_), .A2(new_n3700_), .ZN(new_n3701_));
  NOR2_X1    g03509(.A1(\a[78] ), .A2(\a[79] ), .ZN(new_n3702_));
  INV_X1     g03510(.I(new_n3702_), .ZN(new_n3703_));
  NOR3_X1    g03511(.A1(new_n3701_), .A2(new_n3694_), .A3(new_n3703_), .ZN(new_n3704_));
  NAND2_X1   g03512(.A1(new_n3693_), .A2(new_n3704_), .ZN(new_n3705_));
  XOR2_X1    g03513(.A1(new_n3705_), .A2(\a[81] ), .Z(new_n3706_));
  INV_X1     g03514(.I(\a[81] ), .ZN(new_n3707_));
  NAND2_X1   g03515(.A1(new_n3671_), .A2(new_n3620_), .ZN(new_n3708_));
  NAND2_X1   g03516(.A1(new_n3680_), .A2(new_n3683_), .ZN(new_n3709_));
  OAI21_X1   g03517(.A1(new_n3709_), .A2(new_n3708_), .B(new_n3453_), .ZN(new_n3710_));
  INV_X1     g03518(.I(new_n3686_), .ZN(new_n3711_));
  OAI21_X1   g03519(.A1(new_n3710_), .A2(new_n3711_), .B(new_n3444_), .ZN(new_n3712_));
  NAND2_X1   g03520(.A1(new_n3692_), .A2(new_n3698_), .ZN(new_n3713_));
  NOR2_X1    g03521(.A1(new_n3713_), .A2(new_n3712_), .ZN(new_n3714_));
  NAND3_X1   g03522(.A1(new_n3714_), .A2(new_n3444_), .A3(new_n3699_), .ZN(new_n3715_));
  NAND2_X1   g03523(.A1(new_n3677_), .A2(new_n3679_), .ZN(new_n3716_));
  AOI22_X1   g03524(.A1(new_n3716_), .A2(\asqrt[61] ), .B1(new_n3671_), .B2(new_n3620_), .ZN(new_n3717_));
  NOR2_X1    g03525(.A1(new_n3717_), .A2(new_n196_), .ZN(new_n3718_));
  AOI21_X1   g03526(.A1(new_n3614_), .A2(new_n3616_), .B(new_n275_), .ZN(new_n3719_));
  OAI21_X1   g03527(.A1(new_n3620_), .A2(new_n3719_), .B(\asqrt[61] ), .ZN(new_n3720_));
  NAND4_X1   g03528(.A1(new_n3708_), .A2(new_n196_), .A3(new_n3720_), .A4(new_n3681_), .ZN(new_n3721_));
  INV_X1     g03529(.I(new_n3721_), .ZN(new_n3722_));
  NOR3_X1    g03530(.A1(new_n3713_), .A2(new_n3712_), .A3(new_n3699_), .ZN(\asqrt[41] ));
  NAND3_X1   g03531(.A1(\asqrt[41] ), .A2(new_n3718_), .A3(new_n3722_), .ZN(new_n3724_));
  OAI21_X1   g03532(.A1(new_n3691_), .A2(\asqrt[62] ), .B(new_n3451_), .ZN(new_n3725_));
  OAI21_X1   g03533(.A1(\asqrt[41] ), .A2(new_n3725_), .B(new_n3718_), .ZN(new_n3726_));
  NAND2_X1   g03534(.A1(new_n3726_), .A2(new_n3724_), .ZN(new_n3727_));
  INV_X1     g03535(.I(new_n3727_), .ZN(new_n3728_));
  NOR3_X1    g03536(.A1(new_n3716_), .A2(\asqrt[61] ), .A3(new_n3668_), .ZN(new_n3729_));
  NAND2_X1   g03537(.A1(\asqrt[41] ), .A2(new_n3729_), .ZN(new_n3730_));
  XOR2_X1    g03538(.A1(new_n3730_), .A2(new_n3680_), .Z(new_n3731_));
  NOR2_X1    g03539(.A1(new_n3731_), .A2(new_n196_), .ZN(new_n3732_));
  INV_X1     g03540(.I(new_n3732_), .ZN(new_n3733_));
  INV_X1     g03541(.I(\a[82] ), .ZN(new_n3734_));
  NOR2_X1    g03542(.A1(\a[80] ), .A2(\a[81] ), .ZN(new_n3735_));
  INV_X1     g03543(.I(new_n3735_), .ZN(new_n3736_));
  NOR3_X1    g03544(.A1(new_n3482_), .A2(new_n3734_), .A3(new_n3736_), .ZN(new_n3737_));
  NAND3_X1   g03545(.A1(new_n3433_), .A2(new_n3469_), .A3(new_n3737_), .ZN(new_n3738_));
  XOR2_X1    g03546(.A1(new_n3738_), .A2(\a[83] ), .Z(new_n3739_));
  INV_X1     g03547(.I(\a[83] ), .ZN(new_n3740_));
  NOR4_X1    g03548(.A1(new_n3713_), .A2(new_n3712_), .A3(new_n3740_), .A4(new_n3699_), .ZN(new_n3741_));
  NOR2_X1    g03549(.A1(new_n3739_), .A2(\a[82] ), .ZN(new_n3742_));
  OAI21_X1   g03550(.A1(new_n3741_), .A2(new_n3742_), .B(new_n3739_), .ZN(new_n3743_));
  INV_X1     g03551(.I(new_n3739_), .ZN(new_n3744_));
  NOR2_X1    g03552(.A1(new_n3689_), .A2(new_n3677_), .ZN(new_n3745_));
  NOR3_X1    g03553(.A1(new_n3690_), .A2(new_n229_), .A3(new_n3682_), .ZN(new_n3746_));
  AOI21_X1   g03554(.A1(new_n3746_), .A2(new_n3745_), .B(new_n3452_), .ZN(new_n3747_));
  AOI21_X1   g03555(.A1(new_n3747_), .A2(new_n3686_), .B(new_n3443_), .ZN(new_n3748_));
  AOI21_X1   g03556(.A1(new_n3691_), .A2(\asqrt[62] ), .B(new_n3444_), .ZN(new_n3749_));
  NOR3_X1    g03557(.A1(new_n3749_), .A2(new_n3721_), .A3(new_n3697_), .ZN(new_n3750_));
  NAND4_X1   g03558(.A1(new_n3750_), .A2(\a[83] ), .A3(new_n3748_), .A4(new_n3700_), .ZN(new_n3751_));
  NAND3_X1   g03559(.A1(new_n3751_), .A2(\a[82] ), .A3(new_n3744_), .ZN(new_n3752_));
  NAND2_X1   g03560(.A1(new_n3743_), .A2(new_n3752_), .ZN(new_n3753_));
  NAND2_X1   g03561(.A1(new_n3467_), .A2(new_n3431_), .ZN(new_n3754_));
  NAND4_X1   g03562(.A1(new_n3471_), .A2(new_n3465_), .A3(new_n3418_), .A4(new_n3754_), .ZN(new_n3755_));
  NOR2_X1    g03563(.A1(new_n3481_), .A2(new_n3734_), .ZN(new_n3756_));
  XOR2_X1    g03564(.A1(new_n3756_), .A2(new_n3755_), .Z(new_n3757_));
  NOR2_X1    g03565(.A1(new_n3757_), .A2(new_n3736_), .ZN(new_n3758_));
  INV_X1     g03566(.I(new_n3758_), .ZN(new_n3759_));
  NAND3_X1   g03567(.A1(new_n3750_), .A2(new_n3748_), .A3(new_n3700_), .ZN(new_n3760_));
  NOR4_X1    g03568(.A1(new_n3720_), .A2(new_n3677_), .A3(new_n3689_), .A4(new_n3682_), .ZN(new_n3761_));
  NOR3_X1    g03569(.A1(new_n3761_), .A2(new_n3452_), .A3(new_n3711_), .ZN(new_n3762_));
  NAND4_X1   g03570(.A1(new_n3717_), .A2(new_n196_), .A3(new_n3444_), .A4(new_n3681_), .ZN(new_n3763_));
  OAI21_X1   g03571(.A1(new_n3762_), .A2(new_n3443_), .B(new_n3763_), .ZN(new_n3764_));
  NAND2_X1   g03572(.A1(new_n3701_), .A2(\asqrt[42] ), .ZN(new_n3765_));
  OAI21_X1   g03573(.A1(new_n3764_), .A2(new_n3765_), .B(new_n3454_), .ZN(new_n3766_));
  NAND3_X1   g03574(.A1(new_n3766_), .A2(new_n3455_), .A3(new_n3760_), .ZN(new_n3767_));
  INV_X1     g03575(.I(new_n3765_), .ZN(new_n3768_));
  AOI21_X1   g03576(.A1(new_n3693_), .A2(new_n3768_), .B(\a[84] ), .ZN(new_n3769_));
  OAI21_X1   g03577(.A1(new_n3769_), .A2(new_n3456_), .B(\asqrt[41] ), .ZN(new_n3770_));
  NAND4_X1   g03578(.A1(new_n3767_), .A2(new_n3770_), .A3(new_n3208_), .A4(new_n3759_), .ZN(new_n3771_));
  NAND2_X1   g03579(.A1(new_n3771_), .A2(new_n3753_), .ZN(new_n3772_));
  NAND3_X1   g03580(.A1(new_n3743_), .A2(new_n3752_), .A3(new_n3759_), .ZN(new_n3773_));
  AOI21_X1   g03581(.A1(\asqrt[42] ), .A2(new_n3454_), .B(\a[85] ), .ZN(new_n3774_));
  NOR2_X1    g03582(.A1(new_n3472_), .A2(\a[84] ), .ZN(new_n3775_));
  AOI21_X1   g03583(.A1(\asqrt[42] ), .A2(\a[84] ), .B(new_n3458_), .ZN(new_n3776_));
  OAI21_X1   g03584(.A1(new_n3774_), .A2(new_n3775_), .B(new_n3776_), .ZN(new_n3777_));
  INV_X1     g03585(.I(new_n3777_), .ZN(new_n3778_));
  NAND3_X1   g03586(.A1(\asqrt[41] ), .A2(new_n3480_), .A3(new_n3778_), .ZN(new_n3779_));
  OAI21_X1   g03587(.A1(new_n3760_), .A2(new_n3777_), .B(new_n3479_), .ZN(new_n3780_));
  NAND3_X1   g03588(.A1(new_n3779_), .A2(new_n3780_), .A3(new_n2941_), .ZN(new_n3781_));
  AOI21_X1   g03589(.A1(new_n3773_), .A2(\asqrt[43] ), .B(new_n3781_), .ZN(new_n3782_));
  NOR2_X1    g03590(.A1(new_n3772_), .A2(new_n3782_), .ZN(new_n3783_));
  AOI22_X1   g03591(.A1(new_n3771_), .A2(new_n3753_), .B1(\asqrt[43] ), .B2(new_n3773_), .ZN(new_n3784_));
  INV_X1     g03592(.I(new_n3462_), .ZN(new_n3785_));
  AOI21_X1   g03593(.A1(new_n3472_), .A2(new_n3785_), .B(new_n3464_), .ZN(new_n3786_));
  INV_X1     g03594(.I(new_n3473_), .ZN(new_n3787_));
  NOR3_X1    g03595(.A1(new_n3787_), .A2(new_n3786_), .A3(new_n3479_), .ZN(new_n3788_));
  AOI21_X1   g03596(.A1(new_n3490_), .A2(new_n3487_), .B(\asqrt[44] ), .ZN(new_n3789_));
  AND4_X2    g03597(.A1(new_n3788_), .A2(\asqrt[41] ), .A3(new_n3504_), .A4(new_n3789_), .Z(new_n3790_));
  NOR2_X1    g03598(.A1(new_n3788_), .A2(new_n2941_), .ZN(new_n3791_));
  NOR3_X1    g03599(.A1(new_n3790_), .A2(\asqrt[45] ), .A3(new_n3791_), .ZN(new_n3792_));
  OAI21_X1   g03600(.A1(new_n3784_), .A2(new_n2941_), .B(new_n3792_), .ZN(new_n3793_));
  NAND2_X1   g03601(.A1(new_n3793_), .A2(new_n3783_), .ZN(new_n3794_));
  OAI22_X1   g03602(.A1(new_n3784_), .A2(new_n2941_), .B1(new_n3772_), .B2(new_n3782_), .ZN(new_n3795_));
  NAND2_X1   g03603(.A1(new_n3498_), .A2(new_n3500_), .ZN(new_n3796_));
  NAND4_X1   g03604(.A1(\asqrt[41] ), .A2(new_n2728_), .A3(new_n3796_), .A4(new_n3512_), .ZN(new_n3797_));
  XOR2_X1    g03605(.A1(new_n3797_), .A2(new_n3505_), .Z(new_n3798_));
  NAND2_X1   g03606(.A1(new_n3798_), .A2(new_n2488_), .ZN(new_n3799_));
  AOI21_X1   g03607(.A1(new_n3795_), .A2(\asqrt[45] ), .B(new_n3799_), .ZN(new_n3800_));
  NOR2_X1    g03608(.A1(new_n3800_), .A2(new_n3794_), .ZN(new_n3801_));
  AOI22_X1   g03609(.A1(new_n3795_), .A2(\asqrt[45] ), .B1(new_n3793_), .B2(new_n3783_), .ZN(new_n3802_));
  NOR4_X1    g03610(.A1(new_n3760_), .A2(\asqrt[46] ), .A3(new_n3509_), .A4(new_n3513_), .ZN(new_n3803_));
  XOR2_X1    g03611(.A1(new_n3803_), .A2(new_n3520_), .Z(new_n3804_));
  NAND2_X1   g03612(.A1(new_n3804_), .A2(new_n2253_), .ZN(new_n3805_));
  INV_X1     g03613(.I(new_n3805_), .ZN(new_n3806_));
  OAI21_X1   g03614(.A1(new_n3802_), .A2(new_n2488_), .B(new_n3806_), .ZN(new_n3807_));
  NAND2_X1   g03615(.A1(new_n3807_), .A2(new_n3801_), .ZN(new_n3808_));
  OAI22_X1   g03616(.A1(new_n3802_), .A2(new_n2488_), .B1(new_n3800_), .B2(new_n3794_), .ZN(new_n3809_));
  NAND2_X1   g03617(.A1(new_n3511_), .A2(new_n3520_), .ZN(new_n3810_));
  NOR4_X1    g03618(.A1(new_n3760_), .A2(\asqrt[47] ), .A3(new_n3517_), .A4(new_n3810_), .ZN(new_n3811_));
  XNOR2_X1   g03619(.A1(new_n3811_), .A2(new_n3521_), .ZN(new_n3812_));
  NAND2_X1   g03620(.A1(new_n3812_), .A2(new_n2046_), .ZN(new_n3813_));
  AOI21_X1   g03621(.A1(new_n3809_), .A2(\asqrt[47] ), .B(new_n3813_), .ZN(new_n3814_));
  NOR2_X1    g03622(.A1(new_n3814_), .A2(new_n3808_), .ZN(new_n3815_));
  AOI22_X1   g03623(.A1(new_n3809_), .A2(\asqrt[47] ), .B1(new_n3807_), .B2(new_n3801_), .ZN(new_n3816_));
  NOR4_X1    g03624(.A1(new_n3760_), .A2(\asqrt[48] ), .A3(new_n3525_), .A4(new_n3624_), .ZN(new_n3817_));
  XOR2_X1    g03625(.A1(new_n3817_), .A2(new_n3531_), .Z(new_n3818_));
  NAND2_X1   g03626(.A1(new_n3818_), .A2(new_n1854_), .ZN(new_n3819_));
  INV_X1     g03627(.I(new_n3819_), .ZN(new_n3820_));
  OAI21_X1   g03628(.A1(new_n3816_), .A2(new_n2046_), .B(new_n3820_), .ZN(new_n3821_));
  NAND2_X1   g03629(.A1(new_n3821_), .A2(new_n3815_), .ZN(new_n3822_));
  OAI22_X1   g03630(.A1(new_n3816_), .A2(new_n2046_), .B1(new_n3814_), .B2(new_n3808_), .ZN(new_n3823_));
  NOR2_X1    g03631(.A1(new_n3629_), .A2(new_n1854_), .ZN(new_n3824_));
  NOR4_X1    g03632(.A1(new_n3760_), .A2(\asqrt[49] ), .A3(new_n3534_), .A4(new_n3540_), .ZN(new_n3825_));
  XNOR2_X1   g03633(.A1(new_n3825_), .A2(new_n3824_), .ZN(new_n3826_));
  NAND2_X1   g03634(.A1(new_n3826_), .A2(new_n1595_), .ZN(new_n3827_));
  AOI21_X1   g03635(.A1(new_n3823_), .A2(\asqrt[49] ), .B(new_n3827_), .ZN(new_n3828_));
  NOR2_X1    g03636(.A1(new_n3828_), .A2(new_n3822_), .ZN(new_n3829_));
  AOI22_X1   g03637(.A1(new_n3823_), .A2(\asqrt[49] ), .B1(new_n3821_), .B2(new_n3815_), .ZN(new_n3830_));
  NAND2_X1   g03638(.A1(new_n3633_), .A2(\asqrt[50] ), .ZN(new_n3831_));
  NOR4_X1    g03639(.A1(new_n3760_), .A2(\asqrt[50] ), .A3(new_n3543_), .A4(new_n3633_), .ZN(new_n3832_));
  XOR2_X1    g03640(.A1(new_n3832_), .A2(new_n3831_), .Z(new_n3833_));
  NAND2_X1   g03641(.A1(new_n3833_), .A2(new_n1436_), .ZN(new_n3834_));
  INV_X1     g03642(.I(new_n3834_), .ZN(new_n3835_));
  OAI21_X1   g03643(.A1(new_n3830_), .A2(new_n1595_), .B(new_n3835_), .ZN(new_n3836_));
  NAND2_X1   g03644(.A1(new_n3836_), .A2(new_n3829_), .ZN(new_n3837_));
  OAI22_X1   g03645(.A1(new_n3830_), .A2(new_n1595_), .B1(new_n3828_), .B2(new_n3822_), .ZN(new_n3838_));
  NAND2_X1   g03646(.A1(new_n3555_), .A2(\asqrt[51] ), .ZN(new_n3839_));
  NOR4_X1    g03647(.A1(new_n3760_), .A2(\asqrt[51] ), .A3(new_n3550_), .A4(new_n3555_), .ZN(new_n3840_));
  XOR2_X1    g03648(.A1(new_n3840_), .A2(new_n3839_), .Z(new_n3841_));
  NAND2_X1   g03649(.A1(new_n3841_), .A2(new_n1260_), .ZN(new_n3842_));
  AOI21_X1   g03650(.A1(new_n3838_), .A2(\asqrt[51] ), .B(new_n3842_), .ZN(new_n3843_));
  NOR2_X1    g03651(.A1(new_n3843_), .A2(new_n3837_), .ZN(new_n3844_));
  AOI22_X1   g03652(.A1(new_n3838_), .A2(\asqrt[51] ), .B1(new_n3836_), .B2(new_n3829_), .ZN(new_n3845_));
  NAND2_X1   g03653(.A1(new_n3640_), .A2(\asqrt[52] ), .ZN(new_n3846_));
  NOR4_X1    g03654(.A1(new_n3760_), .A2(\asqrt[52] ), .A3(new_n3558_), .A4(new_n3640_), .ZN(new_n3847_));
  XOR2_X1    g03655(.A1(new_n3847_), .A2(new_n3846_), .Z(new_n3848_));
  NAND2_X1   g03656(.A1(new_n3848_), .A2(new_n1096_), .ZN(new_n3849_));
  INV_X1     g03657(.I(new_n3849_), .ZN(new_n3850_));
  OAI21_X1   g03658(.A1(new_n3845_), .A2(new_n1260_), .B(new_n3850_), .ZN(new_n3851_));
  NAND2_X1   g03659(.A1(new_n3851_), .A2(new_n3844_), .ZN(new_n3852_));
  OAI22_X1   g03660(.A1(new_n3845_), .A2(new_n1260_), .B1(new_n3843_), .B2(new_n3837_), .ZN(new_n3853_));
  NOR2_X1    g03661(.A1(new_n3643_), .A2(new_n1096_), .ZN(new_n3854_));
  NOR4_X1    g03662(.A1(new_n3760_), .A2(\asqrt[53] ), .A3(new_n3565_), .A4(new_n3570_), .ZN(new_n3855_));
  XNOR2_X1   g03663(.A1(new_n3855_), .A2(new_n3854_), .ZN(new_n3856_));
  NAND2_X1   g03664(.A1(new_n3856_), .A2(new_n970_), .ZN(new_n3857_));
  AOI21_X1   g03665(.A1(new_n3853_), .A2(\asqrt[53] ), .B(new_n3857_), .ZN(new_n3858_));
  NOR2_X1    g03666(.A1(new_n3858_), .A2(new_n3852_), .ZN(new_n3859_));
  AOI22_X1   g03667(.A1(new_n3853_), .A2(\asqrt[53] ), .B1(new_n3851_), .B2(new_n3844_), .ZN(new_n3860_));
  NOR4_X1    g03668(.A1(new_n3760_), .A2(\asqrt[54] ), .A3(new_n3573_), .A4(new_n3647_), .ZN(new_n3861_));
  XOR2_X1    g03669(.A1(new_n3861_), .A2(new_n3660_), .Z(new_n3862_));
  NAND2_X1   g03670(.A1(new_n3862_), .A2(new_n825_), .ZN(new_n3863_));
  INV_X1     g03671(.I(new_n3863_), .ZN(new_n3864_));
  OAI21_X1   g03672(.A1(new_n3860_), .A2(new_n970_), .B(new_n3864_), .ZN(new_n3865_));
  NAND2_X1   g03673(.A1(new_n3865_), .A2(new_n3859_), .ZN(new_n3866_));
  OAI22_X1   g03674(.A1(new_n3860_), .A2(new_n970_), .B1(new_n3858_), .B2(new_n3852_), .ZN(new_n3867_));
  NOR4_X1    g03675(.A1(new_n3760_), .A2(\asqrt[55] ), .A3(new_n3580_), .A4(new_n3585_), .ZN(new_n3868_));
  XNOR2_X1   g03676(.A1(new_n3868_), .A2(new_n3661_), .ZN(new_n3869_));
  NAND2_X1   g03677(.A1(new_n3869_), .A2(new_n724_), .ZN(new_n3870_));
  AOI21_X1   g03678(.A1(new_n3867_), .A2(\asqrt[55] ), .B(new_n3870_), .ZN(new_n3871_));
  NOR2_X1    g03679(.A1(new_n3871_), .A2(new_n3866_), .ZN(new_n3872_));
  AOI22_X1   g03680(.A1(new_n3867_), .A2(\asqrt[55] ), .B1(new_n3865_), .B2(new_n3859_), .ZN(new_n3873_));
  NOR4_X1    g03681(.A1(new_n3760_), .A2(\asqrt[56] ), .A3(new_n3588_), .A4(new_n3654_), .ZN(new_n3874_));
  XOR2_X1    g03682(.A1(new_n3874_), .A2(new_n3662_), .Z(new_n3875_));
  NAND2_X1   g03683(.A1(new_n3875_), .A2(new_n587_), .ZN(new_n3876_));
  INV_X1     g03684(.I(new_n3876_), .ZN(new_n3877_));
  OAI21_X1   g03685(.A1(new_n3873_), .A2(new_n724_), .B(new_n3877_), .ZN(new_n3878_));
  NAND2_X1   g03686(.A1(new_n3878_), .A2(new_n3872_), .ZN(new_n3879_));
  OAI22_X1   g03687(.A1(new_n3873_), .A2(new_n724_), .B1(new_n3871_), .B2(new_n3866_), .ZN(new_n3880_));
  NOR4_X1    g03688(.A1(new_n3760_), .A2(\asqrt[57] ), .A3(new_n3595_), .A4(new_n3607_), .ZN(new_n3881_));
  XOR2_X1    g03689(.A1(new_n3881_), .A2(new_n3601_), .Z(new_n3882_));
  NAND2_X1   g03690(.A1(new_n3882_), .A2(new_n504_), .ZN(new_n3883_));
  AOI21_X1   g03691(.A1(new_n3880_), .A2(\asqrt[57] ), .B(new_n3883_), .ZN(new_n3884_));
  NOR2_X1    g03692(.A1(new_n3884_), .A2(new_n3879_), .ZN(new_n3885_));
  AOI22_X1   g03693(.A1(new_n3880_), .A2(\asqrt[57] ), .B1(new_n3878_), .B2(new_n3872_), .ZN(new_n3886_));
  NOR4_X1    g03694(.A1(new_n3760_), .A2(\asqrt[58] ), .A3(new_n3603_), .A4(new_n3672_), .ZN(new_n3887_));
  XOR2_X1    g03695(.A1(new_n3887_), .A2(new_n3664_), .Z(new_n3888_));
  NAND2_X1   g03696(.A1(new_n3888_), .A2(new_n376_), .ZN(new_n3889_));
  INV_X1     g03697(.I(new_n3889_), .ZN(new_n3890_));
  OAI21_X1   g03698(.A1(new_n3886_), .A2(new_n504_), .B(new_n3890_), .ZN(new_n3891_));
  NAND2_X1   g03699(.A1(new_n3891_), .A2(new_n3885_), .ZN(new_n3892_));
  OAI22_X1   g03700(.A1(new_n3886_), .A2(new_n504_), .B1(new_n3884_), .B2(new_n3879_), .ZN(new_n3893_));
  NOR4_X1    g03701(.A1(new_n3760_), .A2(\asqrt[59] ), .A3(new_n3610_), .A4(new_n3665_), .ZN(new_n3894_));
  XOR2_X1    g03702(.A1(new_n3894_), .A2(new_n3616_), .Z(new_n3895_));
  NAND2_X1   g03703(.A1(new_n3895_), .A2(new_n275_), .ZN(new_n3896_));
  AOI21_X1   g03704(.A1(new_n3893_), .A2(\asqrt[59] ), .B(new_n3896_), .ZN(new_n3897_));
  NOR2_X1    g03705(.A1(new_n3897_), .A2(new_n3892_), .ZN(new_n3898_));
  AOI22_X1   g03706(.A1(new_n3893_), .A2(\asqrt[59] ), .B1(new_n3891_), .B2(new_n3885_), .ZN(new_n3899_));
  NOR4_X1    g03707(.A1(new_n3760_), .A2(\asqrt[60] ), .A3(new_n3618_), .A4(new_n3688_), .ZN(new_n3900_));
  XOR2_X1    g03708(.A1(new_n3900_), .A2(new_n3679_), .Z(new_n3901_));
  NAND2_X1   g03709(.A1(new_n3901_), .A2(new_n229_), .ZN(new_n3902_));
  INV_X1     g03710(.I(new_n3902_), .ZN(new_n3903_));
  OAI21_X1   g03711(.A1(new_n3899_), .A2(new_n275_), .B(new_n3903_), .ZN(new_n3904_));
  NAND2_X1   g03712(.A1(new_n3904_), .A2(new_n3898_), .ZN(new_n3905_));
  OAI22_X1   g03713(.A1(new_n3899_), .A2(new_n275_), .B1(new_n3897_), .B2(new_n3892_), .ZN(new_n3906_));
  INV_X1     g03714(.I(new_n3731_), .ZN(new_n3907_));
  NOR2_X1    g03715(.A1(new_n3907_), .A2(\asqrt[62] ), .ZN(new_n3908_));
  INV_X1     g03716(.I(new_n3908_), .ZN(new_n3909_));
  NAND3_X1   g03717(.A1(new_n3906_), .A2(\asqrt[61] ), .A3(new_n3909_), .ZN(new_n3910_));
  OAI21_X1   g03718(.A1(new_n3910_), .A2(new_n3905_), .B(new_n3733_), .ZN(new_n3911_));
  NAND3_X1   g03719(.A1(new_n3760_), .A2(new_n3443_), .A3(new_n3763_), .ZN(new_n3912_));
  AOI21_X1   g03720(.A1(new_n3912_), .A2(new_n3710_), .B(\asqrt[63] ), .ZN(new_n3913_));
  INV_X1     g03721(.I(new_n3913_), .ZN(new_n3914_));
  OAI21_X1   g03722(.A1(new_n3911_), .A2(new_n3914_), .B(new_n3728_), .ZN(new_n3915_));
  INV_X1     g03723(.I(new_n3742_), .ZN(new_n3916_));
  AOI21_X1   g03724(.A1(new_n3751_), .A2(new_n3916_), .B(new_n3744_), .ZN(new_n3917_));
  NOR3_X1    g03725(.A1(new_n3741_), .A2(new_n3734_), .A3(new_n3739_), .ZN(new_n3918_));
  NOR2_X1    g03726(.A1(new_n3918_), .A2(new_n3917_), .ZN(new_n3919_));
  NOR3_X1    g03727(.A1(new_n3769_), .A2(new_n3456_), .A3(\asqrt[41] ), .ZN(new_n3920_));
  AOI21_X1   g03728(.A1(new_n3766_), .A2(new_n3455_), .B(new_n3760_), .ZN(new_n3921_));
  NOR4_X1    g03729(.A1(new_n3921_), .A2(new_n3920_), .A3(\asqrt[43] ), .A4(new_n3758_), .ZN(new_n3922_));
  NOR2_X1    g03730(.A1(new_n3922_), .A2(new_n3919_), .ZN(new_n3923_));
  NOR3_X1    g03731(.A1(new_n3918_), .A2(new_n3917_), .A3(new_n3758_), .ZN(new_n3924_));
  NOR3_X1    g03732(.A1(new_n3760_), .A2(new_n3479_), .A3(new_n3777_), .ZN(new_n3925_));
  AOI21_X1   g03733(.A1(\asqrt[41] ), .A2(new_n3778_), .B(new_n3480_), .ZN(new_n3926_));
  NOR3_X1    g03734(.A1(new_n3926_), .A2(new_n3925_), .A3(\asqrt[44] ), .ZN(new_n3927_));
  OAI21_X1   g03735(.A1(new_n3924_), .A2(new_n3208_), .B(new_n3927_), .ZN(new_n3928_));
  NAND2_X1   g03736(.A1(new_n3923_), .A2(new_n3928_), .ZN(new_n3929_));
  OAI22_X1   g03737(.A1(new_n3922_), .A2(new_n3919_), .B1(new_n3208_), .B2(new_n3924_), .ZN(new_n3930_));
  INV_X1     g03738(.I(new_n3792_), .ZN(new_n3931_));
  AOI21_X1   g03739(.A1(new_n3930_), .A2(\asqrt[44] ), .B(new_n3931_), .ZN(new_n3932_));
  NOR2_X1    g03740(.A1(new_n3932_), .A2(new_n3929_), .ZN(new_n3933_));
  AOI22_X1   g03741(.A1(new_n3930_), .A2(\asqrt[44] ), .B1(new_n3923_), .B2(new_n3928_), .ZN(new_n3934_));
  INV_X1     g03742(.I(new_n3799_), .ZN(new_n3935_));
  OAI21_X1   g03743(.A1(new_n3934_), .A2(new_n2728_), .B(new_n3935_), .ZN(new_n3936_));
  NAND2_X1   g03744(.A1(new_n3936_), .A2(new_n3933_), .ZN(new_n3937_));
  OAI22_X1   g03745(.A1(new_n3934_), .A2(new_n2728_), .B1(new_n3932_), .B2(new_n3929_), .ZN(new_n3938_));
  AOI21_X1   g03746(.A1(new_n3938_), .A2(\asqrt[46] ), .B(new_n3805_), .ZN(new_n3939_));
  NOR2_X1    g03747(.A1(new_n3939_), .A2(new_n3937_), .ZN(new_n3940_));
  AOI22_X1   g03748(.A1(new_n3938_), .A2(\asqrt[46] ), .B1(new_n3936_), .B2(new_n3933_), .ZN(new_n3941_));
  INV_X1     g03749(.I(new_n3813_), .ZN(new_n3942_));
  OAI21_X1   g03750(.A1(new_n3941_), .A2(new_n2253_), .B(new_n3942_), .ZN(new_n3943_));
  NAND2_X1   g03751(.A1(new_n3943_), .A2(new_n3940_), .ZN(new_n3944_));
  OAI22_X1   g03752(.A1(new_n3941_), .A2(new_n2253_), .B1(new_n3939_), .B2(new_n3937_), .ZN(new_n3945_));
  AOI21_X1   g03753(.A1(new_n3945_), .A2(\asqrt[48] ), .B(new_n3819_), .ZN(new_n3946_));
  NOR2_X1    g03754(.A1(new_n3946_), .A2(new_n3944_), .ZN(new_n3947_));
  AOI22_X1   g03755(.A1(new_n3945_), .A2(\asqrt[48] ), .B1(new_n3943_), .B2(new_n3940_), .ZN(new_n3948_));
  INV_X1     g03756(.I(new_n3827_), .ZN(new_n3949_));
  OAI21_X1   g03757(.A1(new_n3948_), .A2(new_n1854_), .B(new_n3949_), .ZN(new_n3950_));
  NAND2_X1   g03758(.A1(new_n3950_), .A2(new_n3947_), .ZN(new_n3951_));
  OAI22_X1   g03759(.A1(new_n3948_), .A2(new_n1854_), .B1(new_n3946_), .B2(new_n3944_), .ZN(new_n3952_));
  AOI21_X1   g03760(.A1(new_n3952_), .A2(\asqrt[50] ), .B(new_n3834_), .ZN(new_n3953_));
  NOR2_X1    g03761(.A1(new_n3953_), .A2(new_n3951_), .ZN(new_n3954_));
  AOI22_X1   g03762(.A1(new_n3952_), .A2(\asqrt[50] ), .B1(new_n3950_), .B2(new_n3947_), .ZN(new_n3955_));
  INV_X1     g03763(.I(new_n3842_), .ZN(new_n3956_));
  OAI21_X1   g03764(.A1(new_n3955_), .A2(new_n1436_), .B(new_n3956_), .ZN(new_n3957_));
  NAND2_X1   g03765(.A1(new_n3957_), .A2(new_n3954_), .ZN(new_n3958_));
  OAI22_X1   g03766(.A1(new_n3955_), .A2(new_n1436_), .B1(new_n3953_), .B2(new_n3951_), .ZN(new_n3959_));
  AOI21_X1   g03767(.A1(new_n3959_), .A2(\asqrt[52] ), .B(new_n3849_), .ZN(new_n3960_));
  NOR2_X1    g03768(.A1(new_n3960_), .A2(new_n3958_), .ZN(new_n3961_));
  AOI22_X1   g03769(.A1(new_n3959_), .A2(\asqrt[52] ), .B1(new_n3957_), .B2(new_n3954_), .ZN(new_n3962_));
  INV_X1     g03770(.I(new_n3857_), .ZN(new_n3963_));
  OAI21_X1   g03771(.A1(new_n3962_), .A2(new_n1096_), .B(new_n3963_), .ZN(new_n3964_));
  NAND2_X1   g03772(.A1(new_n3964_), .A2(new_n3961_), .ZN(new_n3965_));
  OAI22_X1   g03773(.A1(new_n3962_), .A2(new_n1096_), .B1(new_n3960_), .B2(new_n3958_), .ZN(new_n3966_));
  AOI21_X1   g03774(.A1(new_n3966_), .A2(\asqrt[54] ), .B(new_n3863_), .ZN(new_n3967_));
  NOR2_X1    g03775(.A1(new_n3967_), .A2(new_n3965_), .ZN(new_n3968_));
  AOI22_X1   g03776(.A1(new_n3966_), .A2(\asqrt[54] ), .B1(new_n3964_), .B2(new_n3961_), .ZN(new_n3969_));
  INV_X1     g03777(.I(new_n3870_), .ZN(new_n3970_));
  OAI21_X1   g03778(.A1(new_n3969_), .A2(new_n825_), .B(new_n3970_), .ZN(new_n3971_));
  NAND2_X1   g03779(.A1(new_n3971_), .A2(new_n3968_), .ZN(new_n3972_));
  OAI22_X1   g03780(.A1(new_n3969_), .A2(new_n825_), .B1(new_n3967_), .B2(new_n3965_), .ZN(new_n3973_));
  AOI21_X1   g03781(.A1(new_n3973_), .A2(\asqrt[56] ), .B(new_n3876_), .ZN(new_n3974_));
  NOR2_X1    g03782(.A1(new_n3974_), .A2(new_n3972_), .ZN(new_n3975_));
  AOI22_X1   g03783(.A1(new_n3973_), .A2(\asqrt[56] ), .B1(new_n3971_), .B2(new_n3968_), .ZN(new_n3976_));
  INV_X1     g03784(.I(new_n3883_), .ZN(new_n3977_));
  OAI21_X1   g03785(.A1(new_n3976_), .A2(new_n587_), .B(new_n3977_), .ZN(new_n3978_));
  NAND2_X1   g03786(.A1(new_n3978_), .A2(new_n3975_), .ZN(new_n3979_));
  OAI22_X1   g03787(.A1(new_n3976_), .A2(new_n587_), .B1(new_n3974_), .B2(new_n3972_), .ZN(new_n3980_));
  AOI21_X1   g03788(.A1(new_n3980_), .A2(\asqrt[58] ), .B(new_n3889_), .ZN(new_n3981_));
  NOR2_X1    g03789(.A1(new_n3981_), .A2(new_n3979_), .ZN(new_n3982_));
  AOI22_X1   g03790(.A1(new_n3980_), .A2(\asqrt[58] ), .B1(new_n3978_), .B2(new_n3975_), .ZN(new_n3983_));
  INV_X1     g03791(.I(new_n3896_), .ZN(new_n3984_));
  OAI21_X1   g03792(.A1(new_n3983_), .A2(new_n376_), .B(new_n3984_), .ZN(new_n3985_));
  NAND2_X1   g03793(.A1(new_n3985_), .A2(new_n3982_), .ZN(new_n3986_));
  OAI22_X1   g03794(.A1(new_n3983_), .A2(new_n376_), .B1(new_n3981_), .B2(new_n3979_), .ZN(new_n3987_));
  AOI21_X1   g03795(.A1(new_n3987_), .A2(\asqrt[60] ), .B(new_n3902_), .ZN(new_n3988_));
  AOI22_X1   g03796(.A1(new_n3987_), .A2(\asqrt[60] ), .B1(new_n3985_), .B2(new_n3982_), .ZN(new_n3989_));
  OAI22_X1   g03797(.A1(new_n3989_), .A2(new_n229_), .B1(new_n3988_), .B2(new_n3986_), .ZN(new_n3990_));
  NOR4_X1    g03798(.A1(new_n3990_), .A2(\asqrt[62] ), .A3(new_n3727_), .A4(new_n3731_), .ZN(new_n3991_));
  NAND2_X1   g03799(.A1(new_n3747_), .A2(new_n3443_), .ZN(new_n3992_));
  XOR2_X1    g03800(.A1(new_n3747_), .A2(\asqrt[63] ), .Z(new_n3993_));
  AOI21_X1   g03801(.A1(\asqrt[41] ), .A2(new_n3992_), .B(new_n3993_), .ZN(new_n3994_));
  NAND2_X1   g03802(.A1(new_n3991_), .A2(new_n3994_), .ZN(new_n3995_));
  NOR4_X1    g03803(.A1(new_n3995_), .A2(new_n3707_), .A3(new_n3715_), .A4(new_n3915_), .ZN(new_n3996_));
  NOR2_X1    g03804(.A1(new_n3707_), .A2(\a[80] ), .ZN(new_n3997_));
  OAI21_X1   g03805(.A1(new_n3996_), .A2(new_n3997_), .B(new_n3706_), .ZN(new_n3998_));
  INV_X1     g03806(.I(new_n3706_), .ZN(new_n3999_));
  INV_X1     g03807(.I(new_n3715_), .ZN(new_n4000_));
  NOR2_X1    g03808(.A1(new_n3988_), .A2(new_n3986_), .ZN(new_n4001_));
  NOR3_X1    g03809(.A1(new_n3989_), .A2(new_n229_), .A3(new_n3908_), .ZN(new_n4002_));
  AOI21_X1   g03810(.A1(new_n4002_), .A2(new_n4001_), .B(new_n3732_), .ZN(new_n4003_));
  AOI21_X1   g03811(.A1(new_n4003_), .A2(new_n3913_), .B(new_n3727_), .ZN(new_n4004_));
  AOI22_X1   g03812(.A1(new_n3906_), .A2(\asqrt[61] ), .B1(new_n3904_), .B2(new_n3898_), .ZN(new_n4005_));
  NAND4_X1   g03813(.A1(new_n4005_), .A2(new_n196_), .A3(new_n3728_), .A4(new_n3907_), .ZN(new_n4006_));
  INV_X1     g03814(.I(new_n3994_), .ZN(new_n4007_));
  NOR2_X1    g03815(.A1(new_n4006_), .A2(new_n4007_), .ZN(new_n4008_));
  NAND4_X1   g03816(.A1(new_n4008_), .A2(new_n4004_), .A3(\a[81] ), .A4(new_n4000_), .ZN(new_n4009_));
  NAND3_X1   g03817(.A1(new_n4009_), .A2(\a[80] ), .A3(new_n3999_), .ZN(new_n4010_));
  NAND2_X1   g03818(.A1(new_n3998_), .A2(new_n4010_), .ZN(new_n4011_));
  NOR2_X1    g03819(.A1(new_n3995_), .A2(new_n3915_), .ZN(new_n4012_));
  NOR4_X1    g03820(.A1(new_n3713_), .A2(new_n3443_), .A3(new_n3762_), .A4(new_n3699_), .ZN(new_n4013_));
  NAND2_X1   g03821(.A1(\asqrt[41] ), .A2(\a[80] ), .ZN(new_n4014_));
  XOR2_X1    g03822(.A1(new_n4014_), .A2(new_n4013_), .Z(new_n4015_));
  NOR2_X1    g03823(.A1(new_n4015_), .A2(new_n3703_), .ZN(new_n4016_));
  INV_X1     g03824(.I(new_n4016_), .ZN(new_n4017_));
  NAND3_X1   g03825(.A1(new_n4008_), .A2(new_n4004_), .A3(new_n4000_), .ZN(new_n4018_));
  NAND2_X1   g03826(.A1(new_n3867_), .A2(\asqrt[55] ), .ZN(new_n4019_));
  AOI21_X1   g03827(.A1(new_n4019_), .A2(new_n3866_), .B(new_n724_), .ZN(new_n4020_));
  OAI21_X1   g03828(.A1(new_n3872_), .A2(new_n4020_), .B(\asqrt[57] ), .ZN(new_n4021_));
  AOI21_X1   g03829(.A1(new_n3879_), .A2(new_n4021_), .B(new_n504_), .ZN(new_n4022_));
  OAI21_X1   g03830(.A1(new_n3885_), .A2(new_n4022_), .B(\asqrt[59] ), .ZN(new_n4023_));
  AOI21_X1   g03831(.A1(new_n3892_), .A2(new_n4023_), .B(new_n275_), .ZN(new_n4024_));
  OAI21_X1   g03832(.A1(new_n3898_), .A2(new_n4024_), .B(\asqrt[61] ), .ZN(new_n4025_));
  NOR3_X1    g03833(.A1(new_n3905_), .A2(new_n4025_), .A3(new_n3908_), .ZN(new_n4026_));
  NOR3_X1    g03834(.A1(new_n4026_), .A2(new_n3732_), .A3(new_n3914_), .ZN(new_n4027_));
  OAI21_X1   g03835(.A1(new_n4027_), .A2(new_n3727_), .B(new_n4006_), .ZN(new_n4028_));
  NOR2_X1    g03836(.A1(new_n4000_), .A2(new_n3994_), .ZN(new_n4029_));
  NAND2_X1   g03837(.A1(new_n4029_), .A2(\asqrt[41] ), .ZN(new_n4030_));
  OAI21_X1   g03838(.A1(new_n4028_), .A2(new_n4030_), .B(new_n3734_), .ZN(new_n4031_));
  NAND3_X1   g03839(.A1(new_n4031_), .A2(new_n3735_), .A3(new_n4018_), .ZN(new_n4032_));
  NOR4_X1    g03840(.A1(new_n3915_), .A2(new_n3715_), .A3(new_n4006_), .A4(new_n4007_), .ZN(\asqrt[40] ));
  NAND2_X1   g03841(.A1(new_n3973_), .A2(\asqrt[56] ), .ZN(new_n4034_));
  AOI21_X1   g03842(.A1(new_n4034_), .A2(new_n3972_), .B(new_n587_), .ZN(new_n4035_));
  OAI21_X1   g03843(.A1(new_n3975_), .A2(new_n4035_), .B(\asqrt[58] ), .ZN(new_n4036_));
  AOI21_X1   g03844(.A1(new_n3979_), .A2(new_n4036_), .B(new_n376_), .ZN(new_n4037_));
  OAI21_X1   g03845(.A1(new_n3982_), .A2(new_n4037_), .B(\asqrt[60] ), .ZN(new_n4038_));
  AOI21_X1   g03846(.A1(new_n3986_), .A2(new_n4038_), .B(new_n229_), .ZN(new_n4039_));
  NAND4_X1   g03847(.A1(new_n4039_), .A2(new_n3898_), .A3(new_n3904_), .A4(new_n3909_), .ZN(new_n4040_));
  NAND3_X1   g03848(.A1(new_n4040_), .A2(new_n3733_), .A3(new_n3913_), .ZN(new_n4041_));
  AOI21_X1   g03849(.A1(new_n3728_), .A2(new_n4041_), .B(new_n3991_), .ZN(new_n4042_));
  INV_X1     g03850(.I(new_n4030_), .ZN(new_n4043_));
  AOI21_X1   g03851(.A1(new_n4042_), .A2(new_n4043_), .B(\a[82] ), .ZN(new_n4044_));
  OAI21_X1   g03852(.A1(new_n4044_), .A2(new_n3736_), .B(\asqrt[40] ), .ZN(new_n4045_));
  NAND4_X1   g03853(.A1(new_n4045_), .A2(new_n4032_), .A3(new_n3481_), .A4(new_n4017_), .ZN(new_n4046_));
  NAND2_X1   g03854(.A1(new_n4046_), .A2(new_n4011_), .ZN(new_n4047_));
  NAND3_X1   g03855(.A1(new_n3998_), .A2(new_n4010_), .A3(new_n4017_), .ZN(new_n4048_));
  AOI21_X1   g03856(.A1(\asqrt[41] ), .A2(new_n3734_), .B(\a[83] ), .ZN(new_n4049_));
  NOR2_X1    g03857(.A1(new_n3751_), .A2(\a[82] ), .ZN(new_n4050_));
  AOI21_X1   g03858(.A1(\asqrt[41] ), .A2(\a[82] ), .B(new_n3738_), .ZN(new_n4051_));
  OAI21_X1   g03859(.A1(new_n4050_), .A2(new_n4049_), .B(new_n4051_), .ZN(new_n4052_));
  INV_X1     g03860(.I(new_n4052_), .ZN(new_n4053_));
  NAND3_X1   g03861(.A1(\asqrt[40] ), .A2(new_n3759_), .A3(new_n4053_), .ZN(new_n4054_));
  OAI21_X1   g03862(.A1(new_n4018_), .A2(new_n4052_), .B(new_n3758_), .ZN(new_n4055_));
  NAND3_X1   g03863(.A1(new_n4055_), .A2(new_n4054_), .A3(new_n3208_), .ZN(new_n4056_));
  AOI21_X1   g03864(.A1(new_n4048_), .A2(\asqrt[42] ), .B(new_n4056_), .ZN(new_n4057_));
  NOR2_X1    g03865(.A1(new_n4047_), .A2(new_n4057_), .ZN(new_n4058_));
  NAND2_X1   g03866(.A1(new_n4048_), .A2(\asqrt[42] ), .ZN(new_n4059_));
  AOI21_X1   g03867(.A1(new_n4047_), .A2(new_n4059_), .B(new_n3208_), .ZN(new_n4060_));
  NOR2_X1    g03868(.A1(new_n3921_), .A2(new_n3920_), .ZN(new_n4061_));
  NOR4_X1    g03869(.A1(new_n4018_), .A2(\asqrt[43] ), .A3(new_n4061_), .A4(new_n3773_), .ZN(new_n4062_));
  AOI21_X1   g03870(.A1(new_n3919_), .A2(new_n3759_), .B(new_n3208_), .ZN(new_n4063_));
  NOR2_X1    g03871(.A1(new_n4062_), .A2(new_n4063_), .ZN(new_n4064_));
  NAND2_X1   g03872(.A1(new_n4064_), .A2(new_n2941_), .ZN(new_n4065_));
  OAI21_X1   g03873(.A1(new_n4060_), .A2(new_n4065_), .B(new_n4058_), .ZN(new_n4066_));
  OAI21_X1   g03874(.A1(new_n4060_), .A2(new_n4058_), .B(\asqrt[44] ), .ZN(new_n4067_));
  NAND2_X1   g03875(.A1(new_n3930_), .A2(\asqrt[44] ), .ZN(new_n4068_));
  NOR2_X1    g03876(.A1(new_n3926_), .A2(new_n3925_), .ZN(new_n4069_));
  NOR4_X1    g03877(.A1(new_n4018_), .A2(\asqrt[44] ), .A3(new_n4069_), .A4(new_n3930_), .ZN(new_n4070_));
  XOR2_X1    g03878(.A1(new_n4070_), .A2(new_n4068_), .Z(new_n4071_));
  NAND2_X1   g03879(.A1(new_n4071_), .A2(new_n2728_), .ZN(new_n4072_));
  INV_X1     g03880(.I(new_n4072_), .ZN(new_n4073_));
  AOI21_X1   g03881(.A1(new_n4067_), .A2(new_n4073_), .B(new_n4066_), .ZN(new_n4074_));
  AOI21_X1   g03882(.A1(new_n4066_), .A2(new_n4067_), .B(new_n2728_), .ZN(new_n4075_));
  NAND2_X1   g03883(.A1(new_n3795_), .A2(\asqrt[45] ), .ZN(new_n4076_));
  NOR2_X1    g03884(.A1(new_n3790_), .A2(new_n3791_), .ZN(new_n4077_));
  NOR4_X1    g03885(.A1(new_n4018_), .A2(\asqrt[45] ), .A3(new_n4077_), .A4(new_n3795_), .ZN(new_n4078_));
  XOR2_X1    g03886(.A1(new_n4078_), .A2(new_n4076_), .Z(new_n4079_));
  NAND2_X1   g03887(.A1(new_n4079_), .A2(new_n2488_), .ZN(new_n4080_));
  OAI21_X1   g03888(.A1(new_n4075_), .A2(new_n4080_), .B(new_n4074_), .ZN(new_n4081_));
  OAI21_X1   g03889(.A1(new_n4074_), .A2(new_n4075_), .B(\asqrt[46] ), .ZN(new_n4082_));
  NOR4_X1    g03890(.A1(new_n4018_), .A2(\asqrt[46] ), .A3(new_n3798_), .A4(new_n3938_), .ZN(new_n4083_));
  AOI21_X1   g03891(.A1(new_n4076_), .A2(new_n3794_), .B(new_n2488_), .ZN(new_n4084_));
  NOR2_X1    g03892(.A1(new_n4083_), .A2(new_n4084_), .ZN(new_n4085_));
  NAND2_X1   g03893(.A1(new_n4085_), .A2(new_n2253_), .ZN(new_n4086_));
  INV_X1     g03894(.I(new_n4086_), .ZN(new_n4087_));
  AOI21_X1   g03895(.A1(new_n4082_), .A2(new_n4087_), .B(new_n4081_), .ZN(new_n4088_));
  AOI22_X1   g03896(.A1(new_n4046_), .A2(new_n4011_), .B1(\asqrt[42] ), .B2(new_n4048_), .ZN(new_n4089_));
  INV_X1     g03897(.I(new_n4065_), .ZN(new_n4090_));
  OAI21_X1   g03898(.A1(new_n4089_), .A2(new_n3208_), .B(new_n4090_), .ZN(new_n4091_));
  OAI22_X1   g03899(.A1(new_n4089_), .A2(new_n3208_), .B1(new_n4047_), .B2(new_n4057_), .ZN(new_n4092_));
  AOI22_X1   g03900(.A1(new_n4092_), .A2(\asqrt[44] ), .B1(new_n4091_), .B2(new_n4058_), .ZN(new_n4093_));
  INV_X1     g03901(.I(new_n4080_), .ZN(new_n4094_));
  OAI21_X1   g03902(.A1(new_n4093_), .A2(new_n2728_), .B(new_n4094_), .ZN(new_n4095_));
  AOI21_X1   g03903(.A1(new_n4092_), .A2(\asqrt[44] ), .B(new_n4072_), .ZN(new_n4096_));
  OAI22_X1   g03904(.A1(new_n4093_), .A2(new_n2728_), .B1(new_n4096_), .B2(new_n4066_), .ZN(new_n4097_));
  AOI22_X1   g03905(.A1(new_n4097_), .A2(\asqrt[46] ), .B1(new_n4095_), .B2(new_n4074_), .ZN(new_n4098_));
  NAND2_X1   g03906(.A1(new_n3809_), .A2(\asqrt[47] ), .ZN(new_n4099_));
  NOR4_X1    g03907(.A1(new_n4018_), .A2(\asqrt[47] ), .A3(new_n3804_), .A4(new_n3809_), .ZN(new_n4100_));
  XOR2_X1    g03908(.A1(new_n4100_), .A2(new_n4099_), .Z(new_n4101_));
  NAND2_X1   g03909(.A1(new_n4101_), .A2(new_n2046_), .ZN(new_n4102_));
  INV_X1     g03910(.I(new_n4102_), .ZN(new_n4103_));
  OAI21_X1   g03911(.A1(new_n4098_), .A2(new_n2253_), .B(new_n4103_), .ZN(new_n4104_));
  NAND2_X1   g03912(.A1(new_n4104_), .A2(new_n4088_), .ZN(new_n4105_));
  AOI21_X1   g03913(.A1(new_n4097_), .A2(\asqrt[46] ), .B(new_n4086_), .ZN(new_n4106_));
  OAI22_X1   g03914(.A1(new_n4098_), .A2(new_n2253_), .B1(new_n4106_), .B2(new_n4081_), .ZN(new_n4107_));
  NOR4_X1    g03915(.A1(new_n4018_), .A2(\asqrt[48] ), .A3(new_n3812_), .A4(new_n3945_), .ZN(new_n4108_));
  AOI21_X1   g03916(.A1(new_n4099_), .A2(new_n3808_), .B(new_n2046_), .ZN(new_n4109_));
  NOR2_X1    g03917(.A1(new_n4108_), .A2(new_n4109_), .ZN(new_n4110_));
  NAND2_X1   g03918(.A1(new_n4110_), .A2(new_n1854_), .ZN(new_n4111_));
  AOI21_X1   g03919(.A1(new_n4107_), .A2(\asqrt[48] ), .B(new_n4111_), .ZN(new_n4112_));
  NOR2_X1    g03920(.A1(new_n4112_), .A2(new_n4105_), .ZN(new_n4113_));
  AOI22_X1   g03921(.A1(new_n4107_), .A2(\asqrt[48] ), .B1(new_n4104_), .B2(new_n4088_), .ZN(new_n4114_));
  NAND2_X1   g03922(.A1(new_n3823_), .A2(\asqrt[49] ), .ZN(new_n4115_));
  NOR4_X1    g03923(.A1(new_n4018_), .A2(\asqrt[49] ), .A3(new_n3818_), .A4(new_n3823_), .ZN(new_n4116_));
  XOR2_X1    g03924(.A1(new_n4116_), .A2(new_n4115_), .Z(new_n4117_));
  NAND2_X1   g03925(.A1(new_n4117_), .A2(new_n1595_), .ZN(new_n4118_));
  INV_X1     g03926(.I(new_n4118_), .ZN(new_n4119_));
  OAI21_X1   g03927(.A1(new_n4114_), .A2(new_n1854_), .B(new_n4119_), .ZN(new_n4120_));
  NAND2_X1   g03928(.A1(new_n4120_), .A2(new_n4113_), .ZN(new_n4121_));
  OAI22_X1   g03929(.A1(new_n4114_), .A2(new_n1854_), .B1(new_n4112_), .B2(new_n4105_), .ZN(new_n4122_));
  NOR4_X1    g03930(.A1(new_n4018_), .A2(\asqrt[50] ), .A3(new_n3826_), .A4(new_n3952_), .ZN(new_n4123_));
  AOI21_X1   g03931(.A1(new_n4115_), .A2(new_n3822_), .B(new_n1595_), .ZN(new_n4124_));
  NOR2_X1    g03932(.A1(new_n4123_), .A2(new_n4124_), .ZN(new_n4125_));
  NAND2_X1   g03933(.A1(new_n4125_), .A2(new_n1436_), .ZN(new_n4126_));
  AOI21_X1   g03934(.A1(new_n4122_), .A2(\asqrt[50] ), .B(new_n4126_), .ZN(new_n4127_));
  NOR2_X1    g03935(.A1(new_n4127_), .A2(new_n4121_), .ZN(new_n4128_));
  AOI22_X1   g03936(.A1(new_n4122_), .A2(\asqrt[50] ), .B1(new_n4120_), .B2(new_n4113_), .ZN(new_n4129_));
  NAND2_X1   g03937(.A1(new_n3838_), .A2(\asqrt[51] ), .ZN(new_n4130_));
  NOR4_X1    g03938(.A1(new_n4018_), .A2(\asqrt[51] ), .A3(new_n3833_), .A4(new_n3838_), .ZN(new_n4131_));
  XOR2_X1    g03939(.A1(new_n4131_), .A2(new_n4130_), .Z(new_n4132_));
  NAND2_X1   g03940(.A1(new_n4132_), .A2(new_n1260_), .ZN(new_n4133_));
  INV_X1     g03941(.I(new_n4133_), .ZN(new_n4134_));
  OAI21_X1   g03942(.A1(new_n4129_), .A2(new_n1436_), .B(new_n4134_), .ZN(new_n4135_));
  NAND2_X1   g03943(.A1(new_n4135_), .A2(new_n4128_), .ZN(new_n4136_));
  OAI22_X1   g03944(.A1(new_n4129_), .A2(new_n1436_), .B1(new_n4127_), .B2(new_n4121_), .ZN(new_n4137_));
  NAND2_X1   g03945(.A1(new_n3959_), .A2(\asqrt[52] ), .ZN(new_n4138_));
  NOR4_X1    g03946(.A1(new_n4018_), .A2(\asqrt[52] ), .A3(new_n3841_), .A4(new_n3959_), .ZN(new_n4139_));
  XOR2_X1    g03947(.A1(new_n4139_), .A2(new_n4138_), .Z(new_n4140_));
  NAND2_X1   g03948(.A1(new_n4140_), .A2(new_n1096_), .ZN(new_n4141_));
  AOI21_X1   g03949(.A1(new_n4137_), .A2(\asqrt[52] ), .B(new_n4141_), .ZN(new_n4142_));
  NOR2_X1    g03950(.A1(new_n4142_), .A2(new_n4136_), .ZN(new_n4143_));
  AOI22_X1   g03951(.A1(new_n4137_), .A2(\asqrt[52] ), .B1(new_n4135_), .B2(new_n4128_), .ZN(new_n4144_));
  NOR4_X1    g03952(.A1(new_n4018_), .A2(\asqrt[53] ), .A3(new_n3848_), .A4(new_n3853_), .ZN(new_n4145_));
  AOI21_X1   g03953(.A1(new_n4138_), .A2(new_n3958_), .B(new_n1096_), .ZN(new_n4146_));
  NOR2_X1    g03954(.A1(new_n4145_), .A2(new_n4146_), .ZN(new_n4147_));
  NAND2_X1   g03955(.A1(new_n4147_), .A2(new_n970_), .ZN(new_n4148_));
  INV_X1     g03956(.I(new_n4148_), .ZN(new_n4149_));
  OAI21_X1   g03957(.A1(new_n4144_), .A2(new_n1096_), .B(new_n4149_), .ZN(new_n4150_));
  NAND2_X1   g03958(.A1(new_n4150_), .A2(new_n4143_), .ZN(new_n4151_));
  OAI22_X1   g03959(.A1(new_n4144_), .A2(new_n1096_), .B1(new_n4142_), .B2(new_n4136_), .ZN(new_n4152_));
  NAND2_X1   g03960(.A1(new_n3966_), .A2(\asqrt[54] ), .ZN(new_n4153_));
  NOR4_X1    g03961(.A1(new_n4018_), .A2(\asqrt[54] ), .A3(new_n3856_), .A4(new_n3966_), .ZN(new_n4154_));
  XOR2_X1    g03962(.A1(new_n4154_), .A2(new_n4153_), .Z(new_n4155_));
  NAND2_X1   g03963(.A1(new_n4155_), .A2(new_n825_), .ZN(new_n4156_));
  AOI21_X1   g03964(.A1(new_n4152_), .A2(\asqrt[54] ), .B(new_n4156_), .ZN(new_n4157_));
  NOR2_X1    g03965(.A1(new_n4157_), .A2(new_n4151_), .ZN(new_n4158_));
  AOI22_X1   g03966(.A1(new_n4152_), .A2(\asqrt[54] ), .B1(new_n4150_), .B2(new_n4143_), .ZN(new_n4159_));
  NOR4_X1    g03967(.A1(new_n4018_), .A2(\asqrt[55] ), .A3(new_n3862_), .A4(new_n3867_), .ZN(new_n4160_));
  XOR2_X1    g03968(.A1(new_n4160_), .A2(new_n4019_), .Z(new_n4161_));
  NAND2_X1   g03969(.A1(new_n4161_), .A2(new_n724_), .ZN(new_n4162_));
  INV_X1     g03970(.I(new_n4162_), .ZN(new_n4163_));
  OAI21_X1   g03971(.A1(new_n4159_), .A2(new_n825_), .B(new_n4163_), .ZN(new_n4164_));
  NAND2_X1   g03972(.A1(new_n4164_), .A2(new_n4158_), .ZN(new_n4165_));
  OAI22_X1   g03973(.A1(new_n4159_), .A2(new_n825_), .B1(new_n4157_), .B2(new_n4151_), .ZN(new_n4166_));
  NOR4_X1    g03974(.A1(new_n4018_), .A2(\asqrt[56] ), .A3(new_n3869_), .A4(new_n3973_), .ZN(new_n4167_));
  XOR2_X1    g03975(.A1(new_n4167_), .A2(new_n4034_), .Z(new_n4168_));
  NAND2_X1   g03976(.A1(new_n4168_), .A2(new_n587_), .ZN(new_n4169_));
  AOI21_X1   g03977(.A1(new_n4166_), .A2(\asqrt[56] ), .B(new_n4169_), .ZN(new_n4170_));
  NOR2_X1    g03978(.A1(new_n4170_), .A2(new_n4165_), .ZN(new_n4171_));
  AOI22_X1   g03979(.A1(new_n4166_), .A2(\asqrt[56] ), .B1(new_n4164_), .B2(new_n4158_), .ZN(new_n4172_));
  NOR4_X1    g03980(.A1(new_n4018_), .A2(\asqrt[57] ), .A3(new_n3875_), .A4(new_n3880_), .ZN(new_n4173_));
  XOR2_X1    g03981(.A1(new_n4173_), .A2(new_n4021_), .Z(new_n4174_));
  AND2_X2    g03982(.A1(new_n4174_), .A2(new_n504_), .Z(new_n4175_));
  OAI21_X1   g03983(.A1(new_n4172_), .A2(new_n587_), .B(new_n4175_), .ZN(new_n4176_));
  NAND2_X1   g03984(.A1(new_n4176_), .A2(new_n4171_), .ZN(new_n4177_));
  OAI22_X1   g03985(.A1(new_n4172_), .A2(new_n587_), .B1(new_n4170_), .B2(new_n4165_), .ZN(new_n4178_));
  NOR4_X1    g03986(.A1(new_n4018_), .A2(\asqrt[58] ), .A3(new_n3882_), .A4(new_n3980_), .ZN(new_n4179_));
  XOR2_X1    g03987(.A1(new_n4179_), .A2(new_n4036_), .Z(new_n4180_));
  NAND2_X1   g03988(.A1(new_n4180_), .A2(new_n376_), .ZN(new_n4181_));
  AOI21_X1   g03989(.A1(new_n4178_), .A2(\asqrt[58] ), .B(new_n4181_), .ZN(new_n4182_));
  NOR2_X1    g03990(.A1(new_n4182_), .A2(new_n4177_), .ZN(new_n4183_));
  AOI22_X1   g03991(.A1(new_n4178_), .A2(\asqrt[58] ), .B1(new_n4176_), .B2(new_n4171_), .ZN(new_n4184_));
  NOR4_X1    g03992(.A1(new_n4018_), .A2(\asqrt[59] ), .A3(new_n3888_), .A4(new_n3893_), .ZN(new_n4185_));
  XOR2_X1    g03993(.A1(new_n4185_), .A2(new_n4023_), .Z(new_n4186_));
  AND2_X2    g03994(.A1(new_n4186_), .A2(new_n275_), .Z(new_n4187_));
  OAI21_X1   g03995(.A1(new_n4184_), .A2(new_n376_), .B(new_n4187_), .ZN(new_n4188_));
  NAND2_X1   g03996(.A1(new_n4188_), .A2(new_n4183_), .ZN(new_n4189_));
  NAND2_X1   g03997(.A1(new_n4137_), .A2(\asqrt[52] ), .ZN(new_n4190_));
  AOI21_X1   g03998(.A1(new_n4190_), .A2(new_n4136_), .B(new_n1096_), .ZN(new_n4191_));
  OAI21_X1   g03999(.A1(new_n4143_), .A2(new_n4191_), .B(\asqrt[54] ), .ZN(new_n4192_));
  AOI21_X1   g04000(.A1(new_n4151_), .A2(new_n4192_), .B(new_n825_), .ZN(new_n4193_));
  OAI21_X1   g04001(.A1(new_n4158_), .A2(new_n4193_), .B(\asqrt[56] ), .ZN(new_n4194_));
  AOI21_X1   g04002(.A1(new_n4165_), .A2(new_n4194_), .B(new_n587_), .ZN(new_n4195_));
  OAI21_X1   g04003(.A1(new_n4171_), .A2(new_n4195_), .B(\asqrt[58] ), .ZN(new_n4196_));
  AOI21_X1   g04004(.A1(new_n4177_), .A2(new_n4196_), .B(new_n376_), .ZN(new_n4197_));
  OAI21_X1   g04005(.A1(new_n4183_), .A2(new_n4197_), .B(\asqrt[60] ), .ZN(new_n4198_));
  AOI21_X1   g04006(.A1(new_n4189_), .A2(new_n4198_), .B(new_n229_), .ZN(new_n4199_));
  NOR2_X1    g04007(.A1(new_n4005_), .A2(new_n196_), .ZN(new_n4200_));
  NOR2_X1    g04008(.A1(new_n3990_), .A2(\asqrt[62] ), .ZN(new_n4201_));
  NAND3_X1   g04009(.A1(new_n4201_), .A2(new_n4200_), .A3(new_n3907_), .ZN(new_n4202_));
  NOR2_X1    g04010(.A1(new_n4018_), .A2(new_n4202_), .ZN(new_n4203_));
  OR3_X2     g04011(.A1(\asqrt[40] ), .A2(new_n3907_), .A3(new_n4201_), .Z(new_n4204_));
  AOI21_X1   g04012(.A1(new_n4204_), .A2(new_n4200_), .B(new_n4203_), .ZN(new_n4205_));
  NOR4_X1    g04013(.A1(new_n4018_), .A2(\asqrt[61] ), .A3(new_n3901_), .A4(new_n3906_), .ZN(new_n4206_));
  XOR2_X1    g04014(.A1(new_n4206_), .A2(new_n4025_), .Z(new_n4207_));
  NOR2_X1    g04015(.A1(new_n4207_), .A2(new_n196_), .ZN(new_n4208_));
  INV_X1     g04016(.I(new_n4208_), .ZN(new_n4209_));
  NOR2_X1    g04017(.A1(new_n4075_), .A2(new_n4080_), .ZN(new_n4210_));
  NOR3_X1    g04018(.A1(new_n4210_), .A2(new_n4066_), .A3(new_n4096_), .ZN(new_n4211_));
  NAND2_X1   g04019(.A1(new_n4082_), .A2(new_n4087_), .ZN(new_n4212_));
  NAND2_X1   g04020(.A1(new_n4212_), .A2(new_n4211_), .ZN(new_n4213_));
  NAND2_X1   g04021(.A1(new_n4081_), .A2(new_n4082_), .ZN(new_n4214_));
  AOI21_X1   g04022(.A1(new_n4214_), .A2(\asqrt[47] ), .B(new_n4102_), .ZN(new_n4215_));
  NOR2_X1    g04023(.A1(new_n4215_), .A2(new_n4213_), .ZN(new_n4216_));
  AOI21_X1   g04024(.A1(new_n4081_), .A2(new_n4082_), .B(new_n2253_), .ZN(new_n4217_));
  OAI21_X1   g04025(.A1(new_n4088_), .A2(new_n4217_), .B(\asqrt[48] ), .ZN(new_n4218_));
  INV_X1     g04026(.I(new_n4111_), .ZN(new_n4219_));
  NAND2_X1   g04027(.A1(new_n4218_), .A2(new_n4219_), .ZN(new_n4220_));
  NAND2_X1   g04028(.A1(new_n4220_), .A2(new_n4216_), .ZN(new_n4221_));
  AOI22_X1   g04029(.A1(new_n4214_), .A2(\asqrt[47] ), .B1(new_n4212_), .B2(new_n4211_), .ZN(new_n4222_));
  OAI22_X1   g04030(.A1(new_n4222_), .A2(new_n2046_), .B1(new_n4215_), .B2(new_n4213_), .ZN(new_n4223_));
  AOI21_X1   g04031(.A1(new_n4223_), .A2(\asqrt[49] ), .B(new_n4118_), .ZN(new_n4224_));
  NOR2_X1    g04032(.A1(new_n4224_), .A2(new_n4221_), .ZN(new_n4225_));
  AOI22_X1   g04033(.A1(new_n4223_), .A2(\asqrt[49] ), .B1(new_n4220_), .B2(new_n4216_), .ZN(new_n4226_));
  INV_X1     g04034(.I(new_n4126_), .ZN(new_n4227_));
  OAI21_X1   g04035(.A1(new_n4226_), .A2(new_n1595_), .B(new_n4227_), .ZN(new_n4228_));
  NAND2_X1   g04036(.A1(new_n4228_), .A2(new_n4225_), .ZN(new_n4229_));
  OAI22_X1   g04037(.A1(new_n4226_), .A2(new_n1595_), .B1(new_n4224_), .B2(new_n4221_), .ZN(new_n4230_));
  AOI21_X1   g04038(.A1(new_n4230_), .A2(\asqrt[51] ), .B(new_n4133_), .ZN(new_n4231_));
  NOR2_X1    g04039(.A1(new_n4231_), .A2(new_n4229_), .ZN(new_n4232_));
  AOI22_X1   g04040(.A1(new_n4230_), .A2(\asqrt[51] ), .B1(new_n4228_), .B2(new_n4225_), .ZN(new_n4233_));
  INV_X1     g04041(.I(new_n4141_), .ZN(new_n4234_));
  OAI21_X1   g04042(.A1(new_n4233_), .A2(new_n1260_), .B(new_n4234_), .ZN(new_n4235_));
  NAND2_X1   g04043(.A1(new_n4235_), .A2(new_n4232_), .ZN(new_n4236_));
  OAI22_X1   g04044(.A1(new_n4233_), .A2(new_n1260_), .B1(new_n4231_), .B2(new_n4229_), .ZN(new_n4237_));
  AOI21_X1   g04045(.A1(new_n4237_), .A2(\asqrt[53] ), .B(new_n4148_), .ZN(new_n4238_));
  NOR2_X1    g04046(.A1(new_n4238_), .A2(new_n4236_), .ZN(new_n4239_));
  AOI22_X1   g04047(.A1(new_n4237_), .A2(\asqrt[53] ), .B1(new_n4235_), .B2(new_n4232_), .ZN(new_n4240_));
  INV_X1     g04048(.I(new_n4156_), .ZN(new_n4241_));
  OAI21_X1   g04049(.A1(new_n4240_), .A2(new_n970_), .B(new_n4241_), .ZN(new_n4242_));
  NAND2_X1   g04050(.A1(new_n4242_), .A2(new_n4239_), .ZN(new_n4243_));
  OAI22_X1   g04051(.A1(new_n4240_), .A2(new_n970_), .B1(new_n4238_), .B2(new_n4236_), .ZN(new_n4244_));
  AOI21_X1   g04052(.A1(new_n4244_), .A2(\asqrt[55] ), .B(new_n4162_), .ZN(new_n4245_));
  NOR2_X1    g04053(.A1(new_n4245_), .A2(new_n4243_), .ZN(new_n4246_));
  AOI22_X1   g04054(.A1(new_n4244_), .A2(\asqrt[55] ), .B1(new_n4242_), .B2(new_n4239_), .ZN(new_n4247_));
  INV_X1     g04055(.I(new_n4169_), .ZN(new_n4248_));
  OAI21_X1   g04056(.A1(new_n4247_), .A2(new_n724_), .B(new_n4248_), .ZN(new_n4249_));
  NAND2_X1   g04057(.A1(new_n4249_), .A2(new_n4246_), .ZN(new_n4250_));
  NAND2_X1   g04058(.A1(new_n4237_), .A2(\asqrt[53] ), .ZN(new_n4251_));
  AOI21_X1   g04059(.A1(new_n4251_), .A2(new_n4236_), .B(new_n970_), .ZN(new_n4252_));
  OAI21_X1   g04060(.A1(new_n4239_), .A2(new_n4252_), .B(\asqrt[55] ), .ZN(new_n4253_));
  AOI21_X1   g04061(.A1(new_n4243_), .A2(new_n4253_), .B(new_n724_), .ZN(new_n4254_));
  OAI21_X1   g04062(.A1(new_n4246_), .A2(new_n4254_), .B(\asqrt[57] ), .ZN(new_n4255_));
  AOI21_X1   g04063(.A1(new_n4255_), .A2(new_n4175_), .B(new_n4250_), .ZN(new_n4256_));
  OAI22_X1   g04064(.A1(new_n4247_), .A2(new_n724_), .B1(new_n4245_), .B2(new_n4243_), .ZN(new_n4257_));
  AOI22_X1   g04065(.A1(new_n4257_), .A2(\asqrt[57] ), .B1(new_n4249_), .B2(new_n4246_), .ZN(new_n4258_));
  INV_X1     g04066(.I(new_n4181_), .ZN(new_n4259_));
  OAI21_X1   g04067(.A1(new_n4258_), .A2(new_n504_), .B(new_n4259_), .ZN(new_n4260_));
  NAND2_X1   g04068(.A1(new_n4260_), .A2(new_n4256_), .ZN(new_n4261_));
  AOI21_X1   g04069(.A1(new_n4250_), .A2(new_n4255_), .B(new_n504_), .ZN(new_n4262_));
  OAI21_X1   g04070(.A1(new_n4256_), .A2(new_n4262_), .B(\asqrt[59] ), .ZN(new_n4263_));
  AOI21_X1   g04071(.A1(new_n4263_), .A2(new_n4187_), .B(new_n4261_), .ZN(new_n4264_));
  NAND2_X1   g04072(.A1(new_n4177_), .A2(new_n4196_), .ZN(new_n4265_));
  AOI22_X1   g04073(.A1(new_n4265_), .A2(\asqrt[59] ), .B1(new_n4260_), .B2(new_n4256_), .ZN(new_n4266_));
  NOR4_X1    g04074(.A1(new_n4018_), .A2(\asqrt[60] ), .A3(new_n3895_), .A4(new_n3987_), .ZN(new_n4267_));
  XOR2_X1    g04075(.A1(new_n4267_), .A2(new_n4038_), .Z(new_n4268_));
  NAND2_X1   g04076(.A1(new_n4268_), .A2(new_n229_), .ZN(new_n4269_));
  INV_X1     g04077(.I(new_n4269_), .ZN(new_n4270_));
  OAI21_X1   g04078(.A1(new_n4266_), .A2(new_n275_), .B(new_n4270_), .ZN(new_n4271_));
  NAND2_X1   g04079(.A1(new_n4271_), .A2(new_n4264_), .ZN(new_n4272_));
  INV_X1     g04080(.I(new_n4207_), .ZN(new_n4273_));
  NOR2_X1    g04081(.A1(new_n4273_), .A2(\asqrt[62] ), .ZN(new_n4274_));
  INV_X1     g04082(.I(new_n4274_), .ZN(new_n4275_));
  NAND2_X1   g04083(.A1(new_n4199_), .A2(new_n4275_), .ZN(new_n4276_));
  OAI21_X1   g04084(.A1(new_n4276_), .A2(new_n4272_), .B(new_n4209_), .ZN(new_n4277_));
  NAND2_X1   g04085(.A1(new_n4006_), .A2(new_n3727_), .ZN(new_n4278_));
  OAI21_X1   g04086(.A1(\asqrt[40] ), .A2(new_n4278_), .B(new_n3911_), .ZN(new_n4279_));
  NAND2_X1   g04087(.A1(new_n4279_), .A2(new_n231_), .ZN(new_n4280_));
  OAI21_X1   g04088(.A1(new_n4277_), .A2(new_n4280_), .B(new_n4205_), .ZN(new_n4281_));
  OAI21_X1   g04089(.A1(new_n3728_), .A2(new_n3911_), .B(\asqrt[40] ), .ZN(new_n4282_));
  XOR2_X1    g04090(.A1(new_n3911_), .A2(\asqrt[63] ), .Z(new_n4283_));
  NAND2_X1   g04091(.A1(new_n4282_), .A2(new_n4283_), .ZN(new_n4284_));
  INV_X1     g04092(.I(new_n4284_), .ZN(new_n4285_));
  INV_X1     g04093(.I(new_n4205_), .ZN(new_n4286_));
  OAI22_X1   g04094(.A1(new_n4184_), .A2(new_n376_), .B1(new_n4182_), .B2(new_n4177_), .ZN(new_n4287_));
  AOI21_X1   g04095(.A1(new_n4287_), .A2(\asqrt[60] ), .B(new_n4269_), .ZN(new_n4288_));
  AOI22_X1   g04096(.A1(new_n4287_), .A2(\asqrt[60] ), .B1(new_n4188_), .B2(new_n4183_), .ZN(new_n4289_));
  OAI22_X1   g04097(.A1(new_n4289_), .A2(new_n229_), .B1(new_n4288_), .B2(new_n4189_), .ZN(new_n4290_));
  NOR4_X1    g04098(.A1(new_n4290_), .A2(\asqrt[62] ), .A3(new_n4286_), .A4(new_n4207_), .ZN(new_n4291_));
  NAND2_X1   g04099(.A1(new_n4291_), .A2(new_n4285_), .ZN(new_n4292_));
  NAND3_X1   g04100(.A1(new_n4012_), .A2(new_n3715_), .A3(new_n3728_), .ZN(new_n4293_));
  NOR3_X1    g04101(.A1(new_n4292_), .A2(new_n4281_), .A3(new_n4293_), .ZN(\asqrt[39] ));
  NAND2_X1   g04102(.A1(new_n4189_), .A2(new_n4198_), .ZN(new_n4295_));
  NOR3_X1    g04103(.A1(new_n4295_), .A2(\asqrt[61] ), .A3(new_n4268_), .ZN(new_n4296_));
  NAND2_X1   g04104(.A1(\asqrt[39] ), .A2(new_n4296_), .ZN(new_n4297_));
  XOR2_X1    g04105(.A1(new_n4297_), .A2(new_n4199_), .Z(new_n4298_));
  INV_X1     g04106(.I(new_n4298_), .ZN(new_n4299_));
  INV_X1     g04107(.I(\a[79] ), .ZN(new_n4300_));
  INV_X1     g04108(.I(\a[78] ), .ZN(new_n4301_));
  NOR2_X1    g04109(.A1(\a[76] ), .A2(\a[77] ), .ZN(new_n4302_));
  INV_X1     g04110(.I(new_n4302_), .ZN(new_n4303_));
  NOR4_X1    g04111(.A1(new_n4028_), .A2(new_n4301_), .A3(new_n4029_), .A4(new_n4303_), .ZN(new_n4304_));
  XOR2_X1    g04112(.A1(new_n4304_), .A2(new_n4300_), .Z(new_n4305_));
  NOR4_X1    g04113(.A1(new_n4292_), .A2(new_n4281_), .A3(new_n4300_), .A4(new_n4293_), .ZN(new_n4306_));
  NOR2_X1    g04114(.A1(new_n4300_), .A2(\a[78] ), .ZN(new_n4307_));
  OAI21_X1   g04115(.A1(new_n4306_), .A2(new_n4307_), .B(new_n4305_), .ZN(new_n4308_));
  INV_X1     g04116(.I(new_n4305_), .ZN(new_n4309_));
  NOR2_X1    g04117(.A1(new_n4288_), .A2(new_n4189_), .ZN(new_n4310_));
  NOR3_X1    g04118(.A1(new_n4289_), .A2(new_n229_), .A3(new_n4274_), .ZN(new_n4311_));
  AOI21_X1   g04119(.A1(new_n4311_), .A2(new_n4310_), .B(new_n4208_), .ZN(new_n4312_));
  INV_X1     g04120(.I(new_n4280_), .ZN(new_n4313_));
  AOI21_X1   g04121(.A1(new_n4312_), .A2(new_n4313_), .B(new_n4286_), .ZN(new_n4314_));
  AOI21_X1   g04122(.A1(new_n4290_), .A2(\asqrt[62] ), .B(new_n4205_), .ZN(new_n4315_));
  AOI21_X1   g04123(.A1(new_n4261_), .A2(new_n4263_), .B(new_n275_), .ZN(new_n4316_));
  OAI21_X1   g04124(.A1(new_n4264_), .A2(new_n4316_), .B(\asqrt[61] ), .ZN(new_n4317_));
  NAND4_X1   g04125(.A1(new_n4272_), .A2(new_n196_), .A3(new_n4317_), .A4(new_n4273_), .ZN(new_n4318_));
  NOR3_X1    g04126(.A1(new_n4315_), .A2(new_n4284_), .A3(new_n4318_), .ZN(new_n4319_));
  INV_X1     g04127(.I(new_n4293_), .ZN(new_n4320_));
  NAND4_X1   g04128(.A1(new_n4319_), .A2(\a[79] ), .A3(new_n4314_), .A4(new_n4320_), .ZN(new_n4321_));
  NAND3_X1   g04129(.A1(new_n4321_), .A2(\a[78] ), .A3(new_n4309_), .ZN(new_n4322_));
  NAND2_X1   g04130(.A1(new_n4308_), .A2(new_n4322_), .ZN(new_n4323_));
  NOR2_X1    g04131(.A1(new_n4292_), .A2(new_n4281_), .ZN(new_n4324_));
  NOR4_X1    g04132(.A1(new_n3995_), .A2(new_n3715_), .A3(new_n3727_), .A4(new_n4027_), .ZN(new_n4325_));
  NAND2_X1   g04133(.A1(\asqrt[40] ), .A2(\a[78] ), .ZN(new_n4326_));
  XOR2_X1    g04134(.A1(new_n4326_), .A2(new_n4325_), .Z(new_n4327_));
  NOR2_X1    g04135(.A1(new_n4327_), .A2(new_n4303_), .ZN(new_n4328_));
  INV_X1     g04136(.I(new_n4328_), .ZN(new_n4329_));
  NAND3_X1   g04137(.A1(new_n4319_), .A2(new_n4314_), .A3(new_n4320_), .ZN(new_n4330_));
  NOR4_X1    g04138(.A1(new_n4317_), .A2(new_n4189_), .A3(new_n4288_), .A4(new_n4274_), .ZN(new_n4331_));
  NOR3_X1    g04139(.A1(new_n4331_), .A2(new_n4208_), .A3(new_n4280_), .ZN(new_n4332_));
  AOI22_X1   g04140(.A1(new_n4295_), .A2(\asqrt[61] ), .B1(new_n4271_), .B2(new_n4264_), .ZN(new_n4333_));
  NAND4_X1   g04141(.A1(new_n4333_), .A2(new_n196_), .A3(new_n4205_), .A4(new_n4273_), .ZN(new_n4334_));
  OAI21_X1   g04142(.A1(new_n4332_), .A2(new_n4286_), .B(new_n4334_), .ZN(new_n4335_));
  NOR2_X1    g04143(.A1(new_n4285_), .A2(new_n4320_), .ZN(new_n4336_));
  NAND2_X1   g04144(.A1(new_n4336_), .A2(\asqrt[40] ), .ZN(new_n4337_));
  OAI21_X1   g04145(.A1(new_n4335_), .A2(new_n4337_), .B(new_n3694_), .ZN(new_n4338_));
  NAND3_X1   g04146(.A1(new_n4338_), .A2(new_n3702_), .A3(new_n4330_), .ZN(new_n4339_));
  NAND4_X1   g04147(.A1(new_n4199_), .A2(new_n4264_), .A3(new_n4271_), .A4(new_n4275_), .ZN(new_n4340_));
  NAND3_X1   g04148(.A1(new_n4340_), .A2(new_n4209_), .A3(new_n4313_), .ZN(new_n4341_));
  AOI21_X1   g04149(.A1(new_n4205_), .A2(new_n4341_), .B(new_n4291_), .ZN(new_n4342_));
  INV_X1     g04150(.I(new_n4337_), .ZN(new_n4343_));
  AOI21_X1   g04151(.A1(new_n4342_), .A2(new_n4343_), .B(\a[80] ), .ZN(new_n4344_));
  OAI21_X1   g04152(.A1(new_n4344_), .A2(new_n3703_), .B(\asqrt[39] ), .ZN(new_n4345_));
  NAND4_X1   g04153(.A1(new_n4339_), .A2(new_n4345_), .A3(new_n3760_), .A4(new_n4329_), .ZN(new_n4346_));
  NAND2_X1   g04154(.A1(new_n4346_), .A2(new_n4323_), .ZN(new_n4347_));
  NAND3_X1   g04155(.A1(new_n4308_), .A2(new_n4322_), .A3(new_n4329_), .ZN(new_n4348_));
  AOI21_X1   g04156(.A1(\asqrt[40] ), .A2(new_n3694_), .B(\a[81] ), .ZN(new_n4349_));
  NOR2_X1    g04157(.A1(new_n4009_), .A2(\a[80] ), .ZN(new_n4350_));
  AOI21_X1   g04158(.A1(\asqrt[40] ), .A2(\a[80] ), .B(new_n3705_), .ZN(new_n4351_));
  OAI21_X1   g04159(.A1(new_n4349_), .A2(new_n4350_), .B(new_n4351_), .ZN(new_n4352_));
  INV_X1     g04160(.I(new_n4352_), .ZN(new_n4353_));
  NAND3_X1   g04161(.A1(\asqrt[39] ), .A2(new_n4017_), .A3(new_n4353_), .ZN(new_n4354_));
  OAI21_X1   g04162(.A1(new_n4330_), .A2(new_n4352_), .B(new_n4016_), .ZN(new_n4355_));
  NAND3_X1   g04163(.A1(new_n4354_), .A2(new_n4355_), .A3(new_n3481_), .ZN(new_n4356_));
  AOI21_X1   g04164(.A1(new_n4348_), .A2(\asqrt[41] ), .B(new_n4356_), .ZN(new_n4357_));
  NOR2_X1    g04165(.A1(new_n4347_), .A2(new_n4357_), .ZN(new_n4358_));
  AOI22_X1   g04166(.A1(new_n4346_), .A2(new_n4323_), .B1(\asqrt[41] ), .B2(new_n4348_), .ZN(new_n4359_));
  INV_X1     g04167(.I(new_n3997_), .ZN(new_n4360_));
  AOI21_X1   g04168(.A1(new_n4009_), .A2(new_n4360_), .B(new_n3999_), .ZN(new_n4361_));
  INV_X1     g04169(.I(new_n4010_), .ZN(new_n4362_));
  NOR3_X1    g04170(.A1(new_n4362_), .A2(new_n4361_), .A3(new_n4016_), .ZN(new_n4363_));
  AOI21_X1   g04171(.A1(new_n4045_), .A2(new_n4032_), .B(\asqrt[42] ), .ZN(new_n4364_));
  AND4_X2    g04172(.A1(new_n4363_), .A2(\asqrt[39] ), .A3(new_n4059_), .A4(new_n4364_), .Z(new_n4365_));
  NOR2_X1    g04173(.A1(new_n4363_), .A2(new_n3481_), .ZN(new_n4366_));
  NOR3_X1    g04174(.A1(new_n4365_), .A2(\asqrt[43] ), .A3(new_n4366_), .ZN(new_n4367_));
  OAI21_X1   g04175(.A1(new_n4359_), .A2(new_n3481_), .B(new_n4367_), .ZN(new_n4368_));
  NAND2_X1   g04176(.A1(new_n4368_), .A2(new_n4358_), .ZN(new_n4369_));
  OAI22_X1   g04177(.A1(new_n4359_), .A2(new_n3481_), .B1(new_n4347_), .B2(new_n4357_), .ZN(new_n4370_));
  NAND2_X1   g04178(.A1(new_n4055_), .A2(new_n4054_), .ZN(new_n4371_));
  NAND4_X1   g04179(.A1(\asqrt[39] ), .A2(new_n3208_), .A3(new_n4371_), .A4(new_n4089_), .ZN(new_n4372_));
  XOR2_X1    g04180(.A1(new_n4372_), .A2(new_n4060_), .Z(new_n4373_));
  NAND2_X1   g04181(.A1(new_n4373_), .A2(new_n2941_), .ZN(new_n4374_));
  AOI21_X1   g04182(.A1(new_n4370_), .A2(\asqrt[43] ), .B(new_n4374_), .ZN(new_n4375_));
  NOR2_X1    g04183(.A1(new_n4375_), .A2(new_n4369_), .ZN(new_n4376_));
  AOI22_X1   g04184(.A1(new_n4370_), .A2(\asqrt[43] ), .B1(new_n4368_), .B2(new_n4358_), .ZN(new_n4377_));
  NOR4_X1    g04185(.A1(new_n4330_), .A2(\asqrt[44] ), .A3(new_n4064_), .A4(new_n4092_), .ZN(new_n4378_));
  XOR2_X1    g04186(.A1(new_n4378_), .A2(new_n4067_), .Z(new_n4379_));
  NAND2_X1   g04187(.A1(new_n4379_), .A2(new_n2728_), .ZN(new_n4380_));
  INV_X1     g04188(.I(new_n4380_), .ZN(new_n4381_));
  OAI21_X1   g04189(.A1(new_n4377_), .A2(new_n2941_), .B(new_n4381_), .ZN(new_n4382_));
  NAND2_X1   g04190(.A1(new_n4382_), .A2(new_n4376_), .ZN(new_n4383_));
  OAI22_X1   g04191(.A1(new_n4377_), .A2(new_n2941_), .B1(new_n4375_), .B2(new_n4369_), .ZN(new_n4384_));
  NAND2_X1   g04192(.A1(new_n4066_), .A2(new_n4067_), .ZN(new_n4385_));
  NOR4_X1    g04193(.A1(new_n4330_), .A2(\asqrt[45] ), .A3(new_n4071_), .A4(new_n4385_), .ZN(new_n4386_));
  XNOR2_X1   g04194(.A1(new_n4386_), .A2(new_n4075_), .ZN(new_n4387_));
  NAND2_X1   g04195(.A1(new_n4387_), .A2(new_n2488_), .ZN(new_n4388_));
  AOI21_X1   g04196(.A1(new_n4384_), .A2(\asqrt[45] ), .B(new_n4388_), .ZN(new_n4389_));
  NOR2_X1    g04197(.A1(new_n4389_), .A2(new_n4383_), .ZN(new_n4390_));
  AOI22_X1   g04198(.A1(new_n4384_), .A2(\asqrt[45] ), .B1(new_n4382_), .B2(new_n4376_), .ZN(new_n4391_));
  NOR4_X1    g04199(.A1(new_n4330_), .A2(\asqrt[46] ), .A3(new_n4079_), .A4(new_n4097_), .ZN(new_n4392_));
  XOR2_X1    g04200(.A1(new_n4392_), .A2(new_n4082_), .Z(new_n4393_));
  NAND2_X1   g04201(.A1(new_n4393_), .A2(new_n2253_), .ZN(new_n4394_));
  INV_X1     g04202(.I(new_n4394_), .ZN(new_n4395_));
  OAI21_X1   g04203(.A1(new_n4391_), .A2(new_n2488_), .B(new_n4395_), .ZN(new_n4396_));
  NAND2_X1   g04204(.A1(new_n4396_), .A2(new_n4390_), .ZN(new_n4397_));
  OAI22_X1   g04205(.A1(new_n4391_), .A2(new_n2488_), .B1(new_n4389_), .B2(new_n4383_), .ZN(new_n4398_));
  NOR4_X1    g04206(.A1(new_n4330_), .A2(\asqrt[47] ), .A3(new_n4085_), .A4(new_n4214_), .ZN(new_n4399_));
  XNOR2_X1   g04207(.A1(new_n4399_), .A2(new_n4217_), .ZN(new_n4400_));
  NAND2_X1   g04208(.A1(new_n4400_), .A2(new_n2046_), .ZN(new_n4401_));
  AOI21_X1   g04209(.A1(new_n4398_), .A2(\asqrt[47] ), .B(new_n4401_), .ZN(new_n4402_));
  NOR2_X1    g04210(.A1(new_n4402_), .A2(new_n4397_), .ZN(new_n4403_));
  AOI22_X1   g04211(.A1(new_n4398_), .A2(\asqrt[47] ), .B1(new_n4396_), .B2(new_n4390_), .ZN(new_n4404_));
  NOR4_X1    g04212(.A1(new_n4330_), .A2(\asqrt[48] ), .A3(new_n4101_), .A4(new_n4107_), .ZN(new_n4405_));
  XOR2_X1    g04213(.A1(new_n4405_), .A2(new_n4218_), .Z(new_n4406_));
  NAND2_X1   g04214(.A1(new_n4406_), .A2(new_n1854_), .ZN(new_n4407_));
  INV_X1     g04215(.I(new_n4407_), .ZN(new_n4408_));
  OAI21_X1   g04216(.A1(new_n4404_), .A2(new_n2046_), .B(new_n4408_), .ZN(new_n4409_));
  NAND2_X1   g04217(.A1(new_n4409_), .A2(new_n4403_), .ZN(new_n4410_));
  OAI22_X1   g04218(.A1(new_n4404_), .A2(new_n2046_), .B1(new_n4402_), .B2(new_n4397_), .ZN(new_n4411_));
  NAND2_X1   g04219(.A1(new_n4223_), .A2(\asqrt[49] ), .ZN(new_n4412_));
  NOR4_X1    g04220(.A1(new_n4330_), .A2(\asqrt[49] ), .A3(new_n4110_), .A4(new_n4223_), .ZN(new_n4413_));
  XOR2_X1    g04221(.A1(new_n4413_), .A2(new_n4412_), .Z(new_n4414_));
  NAND2_X1   g04222(.A1(new_n4414_), .A2(new_n1595_), .ZN(new_n4415_));
  AOI21_X1   g04223(.A1(new_n4411_), .A2(\asqrt[49] ), .B(new_n4415_), .ZN(new_n4416_));
  NOR2_X1    g04224(.A1(new_n4416_), .A2(new_n4410_), .ZN(new_n4417_));
  AOI22_X1   g04225(.A1(new_n4411_), .A2(\asqrt[49] ), .B1(new_n4409_), .B2(new_n4403_), .ZN(new_n4418_));
  NOR4_X1    g04226(.A1(new_n4330_), .A2(\asqrt[50] ), .A3(new_n4117_), .A4(new_n4122_), .ZN(new_n4419_));
  AOI21_X1   g04227(.A1(new_n4412_), .A2(new_n4221_), .B(new_n1595_), .ZN(new_n4420_));
  NOR2_X1    g04228(.A1(new_n4419_), .A2(new_n4420_), .ZN(new_n4421_));
  NAND2_X1   g04229(.A1(new_n4421_), .A2(new_n1436_), .ZN(new_n4422_));
  INV_X1     g04230(.I(new_n4422_), .ZN(new_n4423_));
  OAI21_X1   g04231(.A1(new_n4418_), .A2(new_n1595_), .B(new_n4423_), .ZN(new_n4424_));
  NAND2_X1   g04232(.A1(new_n4424_), .A2(new_n4417_), .ZN(new_n4425_));
  OAI22_X1   g04233(.A1(new_n4418_), .A2(new_n1595_), .B1(new_n4416_), .B2(new_n4410_), .ZN(new_n4426_));
  NOR2_X1    g04234(.A1(new_n4129_), .A2(new_n1436_), .ZN(new_n4427_));
  NOR4_X1    g04235(.A1(new_n4330_), .A2(\asqrt[51] ), .A3(new_n4125_), .A4(new_n4230_), .ZN(new_n4428_));
  XNOR2_X1   g04236(.A1(new_n4428_), .A2(new_n4427_), .ZN(new_n4429_));
  NAND2_X1   g04237(.A1(new_n4429_), .A2(new_n1260_), .ZN(new_n4430_));
  AOI21_X1   g04238(.A1(new_n4426_), .A2(\asqrt[51] ), .B(new_n4430_), .ZN(new_n4431_));
  NOR2_X1    g04239(.A1(new_n4431_), .A2(new_n4425_), .ZN(new_n4432_));
  AOI22_X1   g04240(.A1(new_n4426_), .A2(\asqrt[51] ), .B1(new_n4424_), .B2(new_n4417_), .ZN(new_n4433_));
  NOR4_X1    g04241(.A1(new_n4330_), .A2(\asqrt[52] ), .A3(new_n4132_), .A4(new_n4137_), .ZN(new_n4434_));
  XOR2_X1    g04242(.A1(new_n4434_), .A2(new_n4190_), .Z(new_n4435_));
  NAND2_X1   g04243(.A1(new_n4435_), .A2(new_n1096_), .ZN(new_n4436_));
  INV_X1     g04244(.I(new_n4436_), .ZN(new_n4437_));
  OAI21_X1   g04245(.A1(new_n4433_), .A2(new_n1260_), .B(new_n4437_), .ZN(new_n4438_));
  NAND2_X1   g04246(.A1(new_n4438_), .A2(new_n4432_), .ZN(new_n4439_));
  OAI22_X1   g04247(.A1(new_n4433_), .A2(new_n1260_), .B1(new_n4431_), .B2(new_n4425_), .ZN(new_n4440_));
  NOR4_X1    g04248(.A1(new_n4330_), .A2(\asqrt[53] ), .A3(new_n4140_), .A4(new_n4237_), .ZN(new_n4441_));
  XOR2_X1    g04249(.A1(new_n4441_), .A2(new_n4251_), .Z(new_n4442_));
  NAND2_X1   g04250(.A1(new_n4442_), .A2(new_n970_), .ZN(new_n4443_));
  AOI21_X1   g04251(.A1(new_n4440_), .A2(\asqrt[53] ), .B(new_n4443_), .ZN(new_n4444_));
  NOR2_X1    g04252(.A1(new_n4444_), .A2(new_n4439_), .ZN(new_n4445_));
  AOI22_X1   g04253(.A1(new_n4440_), .A2(\asqrt[53] ), .B1(new_n4438_), .B2(new_n4432_), .ZN(new_n4446_));
  NOR4_X1    g04254(.A1(new_n4330_), .A2(\asqrt[54] ), .A3(new_n4147_), .A4(new_n4152_), .ZN(new_n4447_));
  XOR2_X1    g04255(.A1(new_n4447_), .A2(new_n4192_), .Z(new_n4448_));
  NAND2_X1   g04256(.A1(new_n4448_), .A2(new_n825_), .ZN(new_n4449_));
  INV_X1     g04257(.I(new_n4449_), .ZN(new_n4450_));
  OAI21_X1   g04258(.A1(new_n4446_), .A2(new_n970_), .B(new_n4450_), .ZN(new_n4451_));
  NAND2_X1   g04259(.A1(new_n4451_), .A2(new_n4445_), .ZN(new_n4452_));
  OAI22_X1   g04260(.A1(new_n4446_), .A2(new_n970_), .B1(new_n4444_), .B2(new_n4439_), .ZN(new_n4453_));
  NOR4_X1    g04261(.A1(new_n4330_), .A2(\asqrt[55] ), .A3(new_n4155_), .A4(new_n4244_), .ZN(new_n4454_));
  XOR2_X1    g04262(.A1(new_n4454_), .A2(new_n4253_), .Z(new_n4455_));
  NAND2_X1   g04263(.A1(new_n4455_), .A2(new_n724_), .ZN(new_n4456_));
  AOI21_X1   g04264(.A1(new_n4453_), .A2(\asqrt[55] ), .B(new_n4456_), .ZN(new_n4457_));
  NOR2_X1    g04265(.A1(new_n4457_), .A2(new_n4452_), .ZN(new_n4458_));
  AOI22_X1   g04266(.A1(new_n4453_), .A2(\asqrt[55] ), .B1(new_n4451_), .B2(new_n4445_), .ZN(new_n4459_));
  NOR4_X1    g04267(.A1(new_n4330_), .A2(\asqrt[56] ), .A3(new_n4161_), .A4(new_n4166_), .ZN(new_n4460_));
  XOR2_X1    g04268(.A1(new_n4460_), .A2(new_n4194_), .Z(new_n4461_));
  NAND2_X1   g04269(.A1(new_n4461_), .A2(new_n587_), .ZN(new_n4462_));
  INV_X1     g04270(.I(new_n4462_), .ZN(new_n4463_));
  OAI21_X1   g04271(.A1(new_n4459_), .A2(new_n724_), .B(new_n4463_), .ZN(new_n4464_));
  NAND2_X1   g04272(.A1(new_n4464_), .A2(new_n4458_), .ZN(new_n4465_));
  OAI22_X1   g04273(.A1(new_n4459_), .A2(new_n724_), .B1(new_n4457_), .B2(new_n4452_), .ZN(new_n4466_));
  NOR4_X1    g04274(.A1(new_n4330_), .A2(\asqrt[57] ), .A3(new_n4168_), .A4(new_n4257_), .ZN(new_n4467_));
  XOR2_X1    g04275(.A1(new_n4467_), .A2(new_n4255_), .Z(new_n4468_));
  NAND2_X1   g04276(.A1(new_n4468_), .A2(new_n504_), .ZN(new_n4469_));
  AOI21_X1   g04277(.A1(new_n4466_), .A2(\asqrt[57] ), .B(new_n4469_), .ZN(new_n4470_));
  NOR2_X1    g04278(.A1(new_n4470_), .A2(new_n4465_), .ZN(new_n4471_));
  AOI22_X1   g04279(.A1(new_n4466_), .A2(\asqrt[57] ), .B1(new_n4464_), .B2(new_n4458_), .ZN(new_n4472_));
  NOR4_X1    g04280(.A1(new_n4330_), .A2(\asqrt[58] ), .A3(new_n4174_), .A4(new_n4178_), .ZN(new_n4473_));
  XOR2_X1    g04281(.A1(new_n4473_), .A2(new_n4196_), .Z(new_n4474_));
  NAND2_X1   g04282(.A1(new_n4474_), .A2(new_n376_), .ZN(new_n4475_));
  INV_X1     g04283(.I(new_n4475_), .ZN(new_n4476_));
  OAI21_X1   g04284(.A1(new_n4472_), .A2(new_n504_), .B(new_n4476_), .ZN(new_n4477_));
  NAND2_X1   g04285(.A1(new_n4477_), .A2(new_n4471_), .ZN(new_n4478_));
  OAI22_X1   g04286(.A1(new_n4472_), .A2(new_n504_), .B1(new_n4470_), .B2(new_n4465_), .ZN(new_n4479_));
  NOR4_X1    g04287(.A1(new_n4330_), .A2(\asqrt[59] ), .A3(new_n4180_), .A4(new_n4265_), .ZN(new_n4480_));
  XOR2_X1    g04288(.A1(new_n4480_), .A2(new_n4263_), .Z(new_n4481_));
  NAND2_X1   g04289(.A1(new_n4481_), .A2(new_n275_), .ZN(new_n4482_));
  AOI21_X1   g04290(.A1(new_n4479_), .A2(\asqrt[59] ), .B(new_n4482_), .ZN(new_n4483_));
  NOR2_X1    g04291(.A1(new_n4483_), .A2(new_n4478_), .ZN(new_n4484_));
  AOI22_X1   g04292(.A1(new_n4479_), .A2(\asqrt[59] ), .B1(new_n4477_), .B2(new_n4471_), .ZN(new_n4485_));
  OAI22_X1   g04293(.A1(new_n4485_), .A2(new_n275_), .B1(new_n4483_), .B2(new_n4478_), .ZN(new_n4486_));
  NOR4_X1    g04294(.A1(new_n4330_), .A2(\asqrt[60] ), .A3(new_n4186_), .A4(new_n4287_), .ZN(new_n4487_));
  XOR2_X1    g04295(.A1(new_n4487_), .A2(new_n4198_), .Z(new_n4488_));
  NAND2_X1   g04296(.A1(new_n4488_), .A2(new_n229_), .ZN(new_n4489_));
  INV_X1     g04297(.I(new_n4489_), .ZN(new_n4490_));
  OAI21_X1   g04298(.A1(new_n4485_), .A2(new_n275_), .B(new_n4490_), .ZN(new_n4491_));
  AOI22_X1   g04299(.A1(new_n4486_), .A2(\asqrt[61] ), .B1(new_n4491_), .B2(new_n4484_), .ZN(new_n4492_));
  NOR2_X1    g04300(.A1(new_n4492_), .A2(new_n196_), .ZN(new_n4493_));
  INV_X1     g04301(.I(new_n4307_), .ZN(new_n4494_));
  AOI21_X1   g04302(.A1(new_n4321_), .A2(new_n4494_), .B(new_n4309_), .ZN(new_n4495_));
  NOR3_X1    g04303(.A1(new_n4306_), .A2(new_n4301_), .A3(new_n4305_), .ZN(new_n4496_));
  NOR2_X1    g04304(.A1(new_n4496_), .A2(new_n4495_), .ZN(new_n4497_));
  NOR3_X1    g04305(.A1(new_n4344_), .A2(new_n3703_), .A3(\asqrt[39] ), .ZN(new_n4498_));
  AOI21_X1   g04306(.A1(new_n4338_), .A2(new_n3702_), .B(new_n4330_), .ZN(new_n4499_));
  NOR4_X1    g04307(.A1(new_n4499_), .A2(new_n4498_), .A3(\asqrt[41] ), .A4(new_n4328_), .ZN(new_n4500_));
  NOR2_X1    g04308(.A1(new_n4500_), .A2(new_n4497_), .ZN(new_n4501_));
  NOR3_X1    g04309(.A1(new_n4496_), .A2(new_n4495_), .A3(new_n4328_), .ZN(new_n4502_));
  NOR3_X1    g04310(.A1(new_n4330_), .A2(new_n4016_), .A3(new_n4352_), .ZN(new_n4503_));
  AOI21_X1   g04311(.A1(\asqrt[39] ), .A2(new_n4353_), .B(new_n4017_), .ZN(new_n4504_));
  NOR3_X1    g04312(.A1(new_n4504_), .A2(new_n4503_), .A3(\asqrt[42] ), .ZN(new_n4505_));
  OAI21_X1   g04313(.A1(new_n4502_), .A2(new_n3760_), .B(new_n4505_), .ZN(new_n4506_));
  NAND2_X1   g04314(.A1(new_n4501_), .A2(new_n4506_), .ZN(new_n4507_));
  OAI22_X1   g04315(.A1(new_n4500_), .A2(new_n4497_), .B1(new_n3760_), .B2(new_n4502_), .ZN(new_n4508_));
  INV_X1     g04316(.I(new_n4367_), .ZN(new_n4509_));
  AOI21_X1   g04317(.A1(new_n4508_), .A2(\asqrt[42] ), .B(new_n4509_), .ZN(new_n4510_));
  NOR2_X1    g04318(.A1(new_n4510_), .A2(new_n4507_), .ZN(new_n4511_));
  AOI22_X1   g04319(.A1(new_n4508_), .A2(\asqrt[42] ), .B1(new_n4501_), .B2(new_n4506_), .ZN(new_n4512_));
  INV_X1     g04320(.I(new_n4374_), .ZN(new_n4513_));
  OAI21_X1   g04321(.A1(new_n4512_), .A2(new_n3208_), .B(new_n4513_), .ZN(new_n4514_));
  NAND2_X1   g04322(.A1(new_n4514_), .A2(new_n4511_), .ZN(new_n4515_));
  OAI22_X1   g04323(.A1(new_n4512_), .A2(new_n3208_), .B1(new_n4510_), .B2(new_n4507_), .ZN(new_n4516_));
  AOI21_X1   g04324(.A1(new_n4516_), .A2(\asqrt[44] ), .B(new_n4380_), .ZN(new_n4517_));
  NOR2_X1    g04325(.A1(new_n4517_), .A2(new_n4515_), .ZN(new_n4518_));
  AOI22_X1   g04326(.A1(new_n4516_), .A2(\asqrt[44] ), .B1(new_n4514_), .B2(new_n4511_), .ZN(new_n4519_));
  INV_X1     g04327(.I(new_n4388_), .ZN(new_n4520_));
  OAI21_X1   g04328(.A1(new_n4519_), .A2(new_n2728_), .B(new_n4520_), .ZN(new_n4521_));
  NAND2_X1   g04329(.A1(new_n4521_), .A2(new_n4518_), .ZN(new_n4522_));
  OAI22_X1   g04330(.A1(new_n4519_), .A2(new_n2728_), .B1(new_n4517_), .B2(new_n4515_), .ZN(new_n4523_));
  AOI21_X1   g04331(.A1(new_n4523_), .A2(\asqrt[46] ), .B(new_n4394_), .ZN(new_n4524_));
  NOR2_X1    g04332(.A1(new_n4524_), .A2(new_n4522_), .ZN(new_n4525_));
  AOI22_X1   g04333(.A1(new_n4523_), .A2(\asqrt[46] ), .B1(new_n4521_), .B2(new_n4518_), .ZN(new_n4526_));
  INV_X1     g04334(.I(new_n4401_), .ZN(new_n4527_));
  OAI21_X1   g04335(.A1(new_n4526_), .A2(new_n2253_), .B(new_n4527_), .ZN(new_n4528_));
  NAND2_X1   g04336(.A1(new_n4528_), .A2(new_n4525_), .ZN(new_n4529_));
  OAI22_X1   g04337(.A1(new_n4526_), .A2(new_n2253_), .B1(new_n4524_), .B2(new_n4522_), .ZN(new_n4530_));
  AOI21_X1   g04338(.A1(new_n4530_), .A2(\asqrt[48] ), .B(new_n4407_), .ZN(new_n4531_));
  NOR2_X1    g04339(.A1(new_n4531_), .A2(new_n4529_), .ZN(new_n4532_));
  AOI22_X1   g04340(.A1(new_n4530_), .A2(\asqrt[48] ), .B1(new_n4528_), .B2(new_n4525_), .ZN(new_n4533_));
  INV_X1     g04341(.I(new_n4415_), .ZN(new_n4534_));
  OAI21_X1   g04342(.A1(new_n4533_), .A2(new_n1854_), .B(new_n4534_), .ZN(new_n4535_));
  NAND2_X1   g04343(.A1(new_n4535_), .A2(new_n4532_), .ZN(new_n4536_));
  OAI22_X1   g04344(.A1(new_n4533_), .A2(new_n1854_), .B1(new_n4531_), .B2(new_n4529_), .ZN(new_n4537_));
  AOI21_X1   g04345(.A1(new_n4537_), .A2(\asqrt[50] ), .B(new_n4422_), .ZN(new_n4538_));
  NOR2_X1    g04346(.A1(new_n4538_), .A2(new_n4536_), .ZN(new_n4539_));
  AOI22_X1   g04347(.A1(new_n4537_), .A2(\asqrt[50] ), .B1(new_n4535_), .B2(new_n4532_), .ZN(new_n4540_));
  INV_X1     g04348(.I(new_n4430_), .ZN(new_n4541_));
  OAI21_X1   g04349(.A1(new_n4540_), .A2(new_n1436_), .B(new_n4541_), .ZN(new_n4542_));
  NAND2_X1   g04350(.A1(new_n4542_), .A2(new_n4539_), .ZN(new_n4543_));
  OAI22_X1   g04351(.A1(new_n4540_), .A2(new_n1436_), .B1(new_n4538_), .B2(new_n4536_), .ZN(new_n4544_));
  AOI21_X1   g04352(.A1(new_n4544_), .A2(\asqrt[52] ), .B(new_n4436_), .ZN(new_n4545_));
  NOR2_X1    g04353(.A1(new_n4545_), .A2(new_n4543_), .ZN(new_n4546_));
  AOI22_X1   g04354(.A1(new_n4544_), .A2(\asqrt[52] ), .B1(new_n4542_), .B2(new_n4539_), .ZN(new_n4547_));
  INV_X1     g04355(.I(new_n4443_), .ZN(new_n4548_));
  OAI21_X1   g04356(.A1(new_n4547_), .A2(new_n1096_), .B(new_n4548_), .ZN(new_n4549_));
  NAND2_X1   g04357(.A1(new_n4549_), .A2(new_n4546_), .ZN(new_n4550_));
  OAI22_X1   g04358(.A1(new_n4547_), .A2(new_n1096_), .B1(new_n4545_), .B2(new_n4543_), .ZN(new_n4551_));
  AOI21_X1   g04359(.A1(new_n4551_), .A2(\asqrt[54] ), .B(new_n4449_), .ZN(new_n4552_));
  NOR2_X1    g04360(.A1(new_n4552_), .A2(new_n4550_), .ZN(new_n4553_));
  AOI22_X1   g04361(.A1(new_n4551_), .A2(\asqrt[54] ), .B1(new_n4549_), .B2(new_n4546_), .ZN(new_n4554_));
  INV_X1     g04362(.I(new_n4456_), .ZN(new_n4555_));
  OAI21_X1   g04363(.A1(new_n4554_), .A2(new_n825_), .B(new_n4555_), .ZN(new_n4556_));
  NAND2_X1   g04364(.A1(new_n4556_), .A2(new_n4553_), .ZN(new_n4557_));
  OAI22_X1   g04365(.A1(new_n4554_), .A2(new_n825_), .B1(new_n4552_), .B2(new_n4550_), .ZN(new_n4558_));
  AOI21_X1   g04366(.A1(new_n4558_), .A2(\asqrt[56] ), .B(new_n4462_), .ZN(new_n4559_));
  NOR2_X1    g04367(.A1(new_n4559_), .A2(new_n4557_), .ZN(new_n4560_));
  AOI22_X1   g04368(.A1(new_n4558_), .A2(\asqrt[56] ), .B1(new_n4556_), .B2(new_n4553_), .ZN(new_n4561_));
  INV_X1     g04369(.I(new_n4469_), .ZN(new_n4562_));
  OAI21_X1   g04370(.A1(new_n4561_), .A2(new_n587_), .B(new_n4562_), .ZN(new_n4563_));
  NAND2_X1   g04371(.A1(new_n4563_), .A2(new_n4560_), .ZN(new_n4564_));
  OAI22_X1   g04372(.A1(new_n4561_), .A2(new_n587_), .B1(new_n4559_), .B2(new_n4557_), .ZN(new_n4565_));
  AOI21_X1   g04373(.A1(new_n4565_), .A2(\asqrt[58] ), .B(new_n4475_), .ZN(new_n4566_));
  NOR2_X1    g04374(.A1(new_n4566_), .A2(new_n4564_), .ZN(new_n4567_));
  AOI22_X1   g04375(.A1(new_n4565_), .A2(\asqrt[58] ), .B1(new_n4563_), .B2(new_n4560_), .ZN(new_n4568_));
  INV_X1     g04376(.I(new_n4482_), .ZN(new_n4569_));
  OAI21_X1   g04377(.A1(new_n4568_), .A2(new_n376_), .B(new_n4569_), .ZN(new_n4570_));
  NAND2_X1   g04378(.A1(new_n4570_), .A2(new_n4567_), .ZN(new_n4571_));
  OAI22_X1   g04379(.A1(new_n4568_), .A2(new_n376_), .B1(new_n4566_), .B2(new_n4564_), .ZN(new_n4572_));
  AOI22_X1   g04380(.A1(new_n4572_), .A2(\asqrt[60] ), .B1(new_n4570_), .B2(new_n4567_), .ZN(new_n4573_));
  AOI21_X1   g04381(.A1(new_n4572_), .A2(\asqrt[60] ), .B(new_n4489_), .ZN(new_n4574_));
  OAI22_X1   g04382(.A1(new_n4573_), .A2(new_n229_), .B1(new_n4574_), .B2(new_n4571_), .ZN(new_n4575_));
  NOR2_X1    g04383(.A1(new_n4575_), .A2(\asqrt[62] ), .ZN(new_n4576_));
  NAND3_X1   g04384(.A1(new_n4324_), .A2(new_n4205_), .A3(new_n4293_), .ZN(new_n4577_));
  NOR2_X1    g04385(.A1(new_n4333_), .A2(new_n196_), .ZN(new_n4578_));
  INV_X1     g04386(.I(new_n4318_), .ZN(new_n4579_));
  NAND3_X1   g04387(.A1(\asqrt[39] ), .A2(new_n4578_), .A3(new_n4579_), .ZN(new_n4580_));
  OAI21_X1   g04388(.A1(new_n4290_), .A2(\asqrt[62] ), .B(new_n4207_), .ZN(new_n4581_));
  OAI21_X1   g04389(.A1(\asqrt[39] ), .A2(new_n4581_), .B(new_n4578_), .ZN(new_n4582_));
  NAND2_X1   g04390(.A1(new_n4582_), .A2(new_n4580_), .ZN(new_n4583_));
  INV_X1     g04391(.I(new_n4583_), .ZN(new_n4584_));
  NOR2_X1    g04392(.A1(new_n4298_), .A2(new_n196_), .ZN(new_n4585_));
  INV_X1     g04393(.I(new_n4585_), .ZN(new_n4586_));
  NAND2_X1   g04394(.A1(new_n4479_), .A2(\asqrt[59] ), .ZN(new_n4587_));
  AOI21_X1   g04395(.A1(new_n4587_), .A2(new_n4478_), .B(new_n275_), .ZN(new_n4588_));
  OAI21_X1   g04396(.A1(new_n4484_), .A2(new_n4588_), .B(\asqrt[61] ), .ZN(new_n4589_));
  NOR2_X1    g04397(.A1(new_n4299_), .A2(\asqrt[62] ), .ZN(new_n4590_));
  INV_X1     g04398(.I(new_n4590_), .ZN(new_n4591_));
  NAND3_X1   g04399(.A1(new_n4491_), .A2(new_n4484_), .A3(new_n4591_), .ZN(new_n4592_));
  OAI21_X1   g04400(.A1(new_n4592_), .A2(new_n4589_), .B(new_n4586_), .ZN(new_n4593_));
  NAND3_X1   g04401(.A1(new_n4330_), .A2(new_n4286_), .A3(new_n4334_), .ZN(new_n4594_));
  AOI21_X1   g04402(.A1(new_n4594_), .A2(new_n4277_), .B(\asqrt[63] ), .ZN(new_n4595_));
  INV_X1     g04403(.I(new_n4595_), .ZN(new_n4596_));
  OAI21_X1   g04404(.A1(new_n4593_), .A2(new_n4596_), .B(new_n4584_), .ZN(new_n4597_));
  NOR4_X1    g04405(.A1(new_n4575_), .A2(\asqrt[62] ), .A3(new_n4583_), .A4(new_n4298_), .ZN(new_n4598_));
  NAND2_X1   g04406(.A1(new_n4312_), .A2(new_n4286_), .ZN(new_n4599_));
  XOR2_X1    g04407(.A1(new_n4312_), .A2(\asqrt[63] ), .Z(new_n4600_));
  AOI21_X1   g04408(.A1(\asqrt[39] ), .A2(new_n4599_), .B(new_n4600_), .ZN(new_n4601_));
  NAND2_X1   g04409(.A1(new_n4598_), .A2(new_n4601_), .ZN(new_n4602_));
  NOR3_X1    g04410(.A1(new_n4602_), .A2(new_n4577_), .A3(new_n4597_), .ZN(\asqrt[38] ));
  NAND4_X1   g04411(.A1(\asqrt[38] ), .A2(new_n4299_), .A3(new_n4493_), .A4(new_n4576_), .ZN(new_n4604_));
  OAI21_X1   g04412(.A1(new_n4575_), .A2(\asqrt[62] ), .B(new_n4298_), .ZN(new_n4605_));
  OAI21_X1   g04413(.A1(\asqrt[38] ), .A2(new_n4605_), .B(new_n4493_), .ZN(new_n4606_));
  NAND2_X1   g04414(.A1(new_n4604_), .A2(new_n4606_), .ZN(new_n4607_));
  INV_X1     g04415(.I(new_n4607_), .ZN(new_n4608_));
  NAND2_X1   g04416(.A1(new_n4565_), .A2(\asqrt[58] ), .ZN(new_n4609_));
  AOI21_X1   g04417(.A1(new_n4609_), .A2(new_n4564_), .B(new_n376_), .ZN(new_n4610_));
  OAI21_X1   g04418(.A1(new_n4567_), .A2(new_n4610_), .B(\asqrt[60] ), .ZN(new_n4611_));
  AOI21_X1   g04419(.A1(new_n4571_), .A2(new_n4611_), .B(new_n229_), .ZN(new_n4612_));
  NOR3_X1    g04420(.A1(new_n4486_), .A2(\asqrt[61] ), .A3(new_n4488_), .ZN(new_n4613_));
  NAND2_X1   g04421(.A1(\asqrt[38] ), .A2(new_n4613_), .ZN(new_n4614_));
  XOR2_X1    g04422(.A1(new_n4614_), .A2(new_n4612_), .Z(new_n4615_));
  NOR2_X1    g04423(.A1(new_n4615_), .A2(new_n196_), .ZN(new_n4616_));
  INV_X1     g04424(.I(new_n4616_), .ZN(new_n4617_));
  INV_X1     g04425(.I(\a[76] ), .ZN(new_n4618_));
  NOR2_X1    g04426(.A1(\a[74] ), .A2(\a[75] ), .ZN(new_n4619_));
  INV_X1     g04427(.I(new_n4619_), .ZN(new_n4620_));
  NOR3_X1    g04428(.A1(new_n4336_), .A2(new_n4618_), .A3(new_n4620_), .ZN(new_n4621_));
  NAND2_X1   g04429(.A1(new_n4342_), .A2(new_n4621_), .ZN(new_n4622_));
  XOR2_X1    g04430(.A1(new_n4622_), .A2(\a[77] ), .Z(new_n4623_));
  INV_X1     g04431(.I(\a[77] ), .ZN(new_n4624_));
  NOR4_X1    g04432(.A1(new_n4602_), .A2(new_n4624_), .A3(new_n4577_), .A4(new_n4597_), .ZN(new_n4625_));
  NOR2_X1    g04433(.A1(new_n4624_), .A2(\a[76] ), .ZN(new_n4626_));
  OAI21_X1   g04434(.A1(new_n4625_), .A2(new_n4626_), .B(new_n4623_), .ZN(new_n4627_));
  INV_X1     g04435(.I(new_n4623_), .ZN(new_n4628_));
  INV_X1     g04436(.I(new_n4577_), .ZN(new_n4629_));
  NOR3_X1    g04437(.A1(new_n4574_), .A2(new_n4571_), .A3(new_n4590_), .ZN(new_n4630_));
  AOI21_X1   g04438(.A1(new_n4630_), .A2(new_n4612_), .B(new_n4585_), .ZN(new_n4631_));
  AOI21_X1   g04439(.A1(new_n4631_), .A2(new_n4595_), .B(new_n4583_), .ZN(new_n4632_));
  NAND4_X1   g04440(.A1(new_n4492_), .A2(new_n196_), .A3(new_n4584_), .A4(new_n4299_), .ZN(new_n4633_));
  INV_X1     g04441(.I(new_n4601_), .ZN(new_n4634_));
  NOR2_X1    g04442(.A1(new_n4633_), .A2(new_n4634_), .ZN(new_n4635_));
  NAND4_X1   g04443(.A1(new_n4635_), .A2(\a[77] ), .A3(new_n4632_), .A4(new_n4629_), .ZN(new_n4636_));
  NAND3_X1   g04444(.A1(new_n4636_), .A2(\a[76] ), .A3(new_n4628_), .ZN(new_n4637_));
  NAND2_X1   g04445(.A1(new_n4627_), .A2(new_n4637_), .ZN(new_n4638_));
  NOR2_X1    g04446(.A1(new_n4602_), .A2(new_n4597_), .ZN(new_n4639_));
  NOR4_X1    g04447(.A1(new_n4292_), .A2(new_n4286_), .A3(new_n4332_), .A4(new_n4293_), .ZN(new_n4640_));
  NAND2_X1   g04448(.A1(\asqrt[39] ), .A2(\a[76] ), .ZN(new_n4641_));
  XOR2_X1    g04449(.A1(new_n4641_), .A2(new_n4640_), .Z(new_n4642_));
  NOR2_X1    g04450(.A1(new_n4642_), .A2(new_n4620_), .ZN(new_n4643_));
  INV_X1     g04451(.I(new_n4643_), .ZN(new_n4644_));
  NAND3_X1   g04452(.A1(new_n4635_), .A2(new_n4629_), .A3(new_n4632_), .ZN(new_n4645_));
  NOR2_X1    g04453(.A1(new_n4629_), .A2(new_n4601_), .ZN(new_n4646_));
  NAND2_X1   g04454(.A1(new_n4646_), .A2(\asqrt[39] ), .ZN(new_n4647_));
  INV_X1     g04455(.I(new_n4647_), .ZN(new_n4648_));
  NAND3_X1   g04456(.A1(new_n4597_), .A2(new_n4633_), .A3(new_n4648_), .ZN(new_n4649_));
  NAND2_X1   g04457(.A1(new_n4649_), .A2(new_n4301_), .ZN(new_n4650_));
  NAND3_X1   g04458(.A1(new_n4650_), .A2(new_n4302_), .A3(new_n4645_), .ZN(new_n4651_));
  NOR3_X1    g04459(.A1(new_n4632_), .A2(new_n4598_), .A3(new_n4647_), .ZN(new_n4652_));
  OAI21_X1   g04460(.A1(new_n4652_), .A2(\a[78] ), .B(new_n4302_), .ZN(new_n4653_));
  NAND2_X1   g04461(.A1(new_n4653_), .A2(\asqrt[38] ), .ZN(new_n4654_));
  NAND4_X1   g04462(.A1(new_n4654_), .A2(new_n4018_), .A3(new_n4651_), .A4(new_n4644_), .ZN(new_n4655_));
  NAND2_X1   g04463(.A1(new_n4655_), .A2(new_n4638_), .ZN(new_n4656_));
  NAND3_X1   g04464(.A1(new_n4627_), .A2(new_n4637_), .A3(new_n4644_), .ZN(new_n4657_));
  NAND2_X1   g04465(.A1(\asqrt[39] ), .A2(new_n4301_), .ZN(new_n4658_));
  AOI22_X1   g04466(.A1(new_n4658_), .A2(new_n4300_), .B1(new_n4301_), .B2(new_n4306_), .ZN(new_n4659_));
  OAI21_X1   g04467(.A1(new_n4330_), .A2(new_n4301_), .B(new_n4304_), .ZN(new_n4660_));
  NOR2_X1    g04468(.A1(new_n4659_), .A2(new_n4660_), .ZN(new_n4661_));
  NAND3_X1   g04469(.A1(\asqrt[38] ), .A2(new_n4329_), .A3(new_n4661_), .ZN(new_n4662_));
  INV_X1     g04470(.I(new_n4661_), .ZN(new_n4663_));
  OAI21_X1   g04471(.A1(new_n4645_), .A2(new_n4663_), .B(new_n4328_), .ZN(new_n4664_));
  NAND3_X1   g04472(.A1(new_n4662_), .A2(new_n4664_), .A3(new_n3760_), .ZN(new_n4665_));
  AOI21_X1   g04473(.A1(new_n4657_), .A2(\asqrt[40] ), .B(new_n4665_), .ZN(new_n4666_));
  NOR2_X1    g04474(.A1(new_n4656_), .A2(new_n4666_), .ZN(new_n4667_));
  NAND2_X1   g04475(.A1(new_n4657_), .A2(\asqrt[40] ), .ZN(new_n4668_));
  AOI21_X1   g04476(.A1(new_n4656_), .A2(new_n4668_), .B(new_n3760_), .ZN(new_n4669_));
  NOR2_X1    g04477(.A1(new_n4499_), .A2(new_n4498_), .ZN(new_n4670_));
  NOR4_X1    g04478(.A1(new_n4645_), .A2(\asqrt[41] ), .A3(new_n4670_), .A4(new_n4348_), .ZN(new_n4671_));
  AOI21_X1   g04479(.A1(new_n4497_), .A2(new_n4329_), .B(new_n3760_), .ZN(new_n4672_));
  NOR2_X1    g04480(.A1(new_n4671_), .A2(new_n4672_), .ZN(new_n4673_));
  NAND2_X1   g04481(.A1(new_n4673_), .A2(new_n3481_), .ZN(new_n4674_));
  OAI21_X1   g04482(.A1(new_n4669_), .A2(new_n4674_), .B(new_n4667_), .ZN(new_n4675_));
  AOI22_X1   g04483(.A1(new_n4655_), .A2(new_n4638_), .B1(\asqrt[40] ), .B2(new_n4657_), .ZN(new_n4676_));
  OAI22_X1   g04484(.A1(new_n4676_), .A2(new_n3760_), .B1(new_n4656_), .B2(new_n4666_), .ZN(new_n4677_));
  NOR2_X1    g04485(.A1(new_n4359_), .A2(new_n3481_), .ZN(new_n4678_));
  NAND2_X1   g04486(.A1(new_n4354_), .A2(new_n4355_), .ZN(new_n4679_));
  NAND4_X1   g04487(.A1(\asqrt[38] ), .A2(new_n3481_), .A3(new_n4679_), .A4(new_n4359_), .ZN(new_n4680_));
  XOR2_X1    g04488(.A1(new_n4680_), .A2(new_n4678_), .Z(new_n4681_));
  NAND2_X1   g04489(.A1(new_n4681_), .A2(new_n3208_), .ZN(new_n4682_));
  AOI21_X1   g04490(.A1(new_n4677_), .A2(\asqrt[42] ), .B(new_n4682_), .ZN(new_n4683_));
  OAI21_X1   g04491(.A1(new_n4669_), .A2(new_n4667_), .B(\asqrt[42] ), .ZN(new_n4684_));
  AOI21_X1   g04492(.A1(new_n4675_), .A2(new_n4684_), .B(new_n3208_), .ZN(new_n4685_));
  NAND2_X1   g04493(.A1(new_n4370_), .A2(\asqrt[43] ), .ZN(new_n4686_));
  OAI21_X1   g04494(.A1(new_n4365_), .A2(new_n4366_), .B(new_n3208_), .ZN(new_n4687_));
  NOR3_X1    g04495(.A1(new_n4645_), .A2(new_n4370_), .A3(new_n4687_), .ZN(new_n4688_));
  XOR2_X1    g04496(.A1(new_n4688_), .A2(new_n4686_), .Z(new_n4689_));
  NAND2_X1   g04497(.A1(new_n4689_), .A2(new_n2941_), .ZN(new_n4690_));
  NOR2_X1    g04498(.A1(new_n4685_), .A2(new_n4690_), .ZN(new_n4691_));
  NOR3_X1    g04499(.A1(new_n4691_), .A2(new_n4675_), .A3(new_n4683_), .ZN(new_n4692_));
  INV_X1     g04500(.I(new_n4682_), .ZN(new_n4693_));
  AOI21_X1   g04501(.A1(new_n4684_), .A2(new_n4693_), .B(new_n4675_), .ZN(new_n4694_));
  OAI21_X1   g04502(.A1(new_n4694_), .A2(new_n4685_), .B(\asqrt[44] ), .ZN(new_n4695_));
  NAND2_X1   g04503(.A1(new_n4516_), .A2(\asqrt[44] ), .ZN(new_n4696_));
  NOR4_X1    g04504(.A1(new_n4645_), .A2(\asqrt[44] ), .A3(new_n4373_), .A4(new_n4516_), .ZN(new_n4697_));
  XOR2_X1    g04505(.A1(new_n4697_), .A2(new_n4696_), .Z(new_n4698_));
  NAND2_X1   g04506(.A1(new_n4698_), .A2(new_n2728_), .ZN(new_n4699_));
  INV_X1     g04507(.I(new_n4699_), .ZN(new_n4700_));
  NAND2_X1   g04508(.A1(new_n4695_), .A2(new_n4700_), .ZN(new_n4701_));
  NAND2_X1   g04509(.A1(new_n4701_), .A2(new_n4692_), .ZN(new_n4702_));
  OAI21_X1   g04510(.A1(new_n4685_), .A2(new_n4690_), .B(new_n4694_), .ZN(new_n4703_));
  NAND2_X1   g04511(.A1(new_n4703_), .A2(new_n4695_), .ZN(new_n4704_));
  NAND2_X1   g04512(.A1(new_n4384_), .A2(\asqrt[45] ), .ZN(new_n4705_));
  NOR4_X1    g04513(.A1(new_n4645_), .A2(\asqrt[45] ), .A3(new_n4379_), .A4(new_n4384_), .ZN(new_n4706_));
  XOR2_X1    g04514(.A1(new_n4706_), .A2(new_n4705_), .Z(new_n4707_));
  NAND2_X1   g04515(.A1(new_n4707_), .A2(new_n2488_), .ZN(new_n4708_));
  AOI21_X1   g04516(.A1(new_n4704_), .A2(\asqrt[45] ), .B(new_n4708_), .ZN(new_n4709_));
  NOR2_X1    g04517(.A1(new_n4709_), .A2(new_n4702_), .ZN(new_n4710_));
  AOI21_X1   g04518(.A1(new_n4695_), .A2(new_n4700_), .B(new_n4703_), .ZN(new_n4711_));
  AOI21_X1   g04519(.A1(new_n4703_), .A2(new_n4695_), .B(new_n2728_), .ZN(new_n4712_));
  OAI21_X1   g04520(.A1(new_n4711_), .A2(new_n4712_), .B(\asqrt[46] ), .ZN(new_n4713_));
  NAND2_X1   g04521(.A1(new_n4523_), .A2(\asqrt[46] ), .ZN(new_n4714_));
  NOR4_X1    g04522(.A1(new_n4645_), .A2(\asqrt[46] ), .A3(new_n4387_), .A4(new_n4523_), .ZN(new_n4715_));
  XOR2_X1    g04523(.A1(new_n4715_), .A2(new_n4714_), .Z(new_n4716_));
  NAND2_X1   g04524(.A1(new_n4716_), .A2(new_n2253_), .ZN(new_n4717_));
  INV_X1     g04525(.I(new_n4717_), .ZN(new_n4718_));
  NAND2_X1   g04526(.A1(new_n4713_), .A2(new_n4718_), .ZN(new_n4719_));
  NAND2_X1   g04527(.A1(new_n4719_), .A2(new_n4710_), .ZN(new_n4720_));
  AOI22_X1   g04528(.A1(new_n4704_), .A2(\asqrt[45] ), .B1(new_n4701_), .B2(new_n4692_), .ZN(new_n4721_));
  OAI22_X1   g04529(.A1(new_n4721_), .A2(new_n2488_), .B1(new_n4709_), .B2(new_n4702_), .ZN(new_n4722_));
  NAND2_X1   g04530(.A1(new_n4398_), .A2(\asqrt[47] ), .ZN(new_n4723_));
  NOR4_X1    g04531(.A1(new_n4645_), .A2(\asqrt[47] ), .A3(new_n4393_), .A4(new_n4398_), .ZN(new_n4724_));
  XOR2_X1    g04532(.A1(new_n4724_), .A2(new_n4723_), .Z(new_n4725_));
  NAND2_X1   g04533(.A1(new_n4725_), .A2(new_n2046_), .ZN(new_n4726_));
  AOI21_X1   g04534(.A1(new_n4722_), .A2(\asqrt[47] ), .B(new_n4726_), .ZN(new_n4727_));
  NOR2_X1    g04535(.A1(new_n4727_), .A2(new_n4720_), .ZN(new_n4728_));
  AOI22_X1   g04536(.A1(new_n4722_), .A2(\asqrt[47] ), .B1(new_n4719_), .B2(new_n4710_), .ZN(new_n4729_));
  NAND2_X1   g04537(.A1(new_n4530_), .A2(\asqrt[48] ), .ZN(new_n4730_));
  NOR4_X1    g04538(.A1(new_n4645_), .A2(\asqrt[48] ), .A3(new_n4400_), .A4(new_n4530_), .ZN(new_n4731_));
  XOR2_X1    g04539(.A1(new_n4731_), .A2(new_n4730_), .Z(new_n4732_));
  NAND2_X1   g04540(.A1(new_n4732_), .A2(new_n1854_), .ZN(new_n4733_));
  INV_X1     g04541(.I(new_n4733_), .ZN(new_n4734_));
  OAI21_X1   g04542(.A1(new_n4729_), .A2(new_n2046_), .B(new_n4734_), .ZN(new_n4735_));
  NAND2_X1   g04543(.A1(new_n4735_), .A2(new_n4728_), .ZN(new_n4736_));
  OAI22_X1   g04544(.A1(new_n4729_), .A2(new_n2046_), .B1(new_n4727_), .B2(new_n4720_), .ZN(new_n4737_));
  NAND2_X1   g04545(.A1(new_n4411_), .A2(\asqrt[49] ), .ZN(new_n4738_));
  NOR4_X1    g04546(.A1(new_n4645_), .A2(\asqrt[49] ), .A3(new_n4406_), .A4(new_n4411_), .ZN(new_n4739_));
  XOR2_X1    g04547(.A1(new_n4739_), .A2(new_n4738_), .Z(new_n4740_));
  NAND2_X1   g04548(.A1(new_n4740_), .A2(new_n1595_), .ZN(new_n4741_));
  AOI21_X1   g04549(.A1(new_n4737_), .A2(\asqrt[49] ), .B(new_n4741_), .ZN(new_n4742_));
  NOR2_X1    g04550(.A1(new_n4742_), .A2(new_n4736_), .ZN(new_n4743_));
  AOI22_X1   g04551(.A1(new_n4737_), .A2(\asqrt[49] ), .B1(new_n4735_), .B2(new_n4728_), .ZN(new_n4744_));
  NAND2_X1   g04552(.A1(new_n4537_), .A2(\asqrt[50] ), .ZN(new_n4745_));
  NOR4_X1    g04553(.A1(new_n4645_), .A2(\asqrt[50] ), .A3(new_n4414_), .A4(new_n4537_), .ZN(new_n4746_));
  XOR2_X1    g04554(.A1(new_n4746_), .A2(new_n4745_), .Z(new_n4747_));
  NAND2_X1   g04555(.A1(new_n4747_), .A2(new_n1436_), .ZN(new_n4748_));
  INV_X1     g04556(.I(new_n4748_), .ZN(new_n4749_));
  OAI21_X1   g04557(.A1(new_n4744_), .A2(new_n1595_), .B(new_n4749_), .ZN(new_n4750_));
  NAND2_X1   g04558(.A1(new_n4750_), .A2(new_n4743_), .ZN(new_n4751_));
  OAI22_X1   g04559(.A1(new_n4744_), .A2(new_n1595_), .B1(new_n4742_), .B2(new_n4736_), .ZN(new_n4752_));
  NAND2_X1   g04560(.A1(new_n4426_), .A2(\asqrt[51] ), .ZN(new_n4753_));
  NOR4_X1    g04561(.A1(new_n4645_), .A2(\asqrt[51] ), .A3(new_n4421_), .A4(new_n4426_), .ZN(new_n4754_));
  XOR2_X1    g04562(.A1(new_n4754_), .A2(new_n4753_), .Z(new_n4755_));
  NAND2_X1   g04563(.A1(new_n4755_), .A2(new_n1260_), .ZN(new_n4756_));
  AOI21_X1   g04564(.A1(new_n4752_), .A2(\asqrt[51] ), .B(new_n4756_), .ZN(new_n4757_));
  NOR2_X1    g04565(.A1(new_n4757_), .A2(new_n4751_), .ZN(new_n4758_));
  AOI22_X1   g04566(.A1(new_n4752_), .A2(\asqrt[51] ), .B1(new_n4750_), .B2(new_n4743_), .ZN(new_n4759_));
  NAND2_X1   g04567(.A1(new_n4544_), .A2(\asqrt[52] ), .ZN(new_n4760_));
  NOR4_X1    g04568(.A1(new_n4645_), .A2(\asqrt[52] ), .A3(new_n4429_), .A4(new_n4544_), .ZN(new_n4761_));
  XOR2_X1    g04569(.A1(new_n4761_), .A2(new_n4760_), .Z(new_n4762_));
  NAND2_X1   g04570(.A1(new_n4762_), .A2(new_n1096_), .ZN(new_n4763_));
  INV_X1     g04571(.I(new_n4763_), .ZN(new_n4764_));
  OAI21_X1   g04572(.A1(new_n4759_), .A2(new_n1260_), .B(new_n4764_), .ZN(new_n4765_));
  NAND2_X1   g04573(.A1(new_n4765_), .A2(new_n4758_), .ZN(new_n4766_));
  OAI22_X1   g04574(.A1(new_n4759_), .A2(new_n1260_), .B1(new_n4757_), .B2(new_n4751_), .ZN(new_n4767_));
  NAND2_X1   g04575(.A1(new_n4440_), .A2(\asqrt[53] ), .ZN(new_n4768_));
  NOR4_X1    g04576(.A1(new_n4645_), .A2(\asqrt[53] ), .A3(new_n4435_), .A4(new_n4440_), .ZN(new_n4769_));
  XOR2_X1    g04577(.A1(new_n4769_), .A2(new_n4768_), .Z(new_n4770_));
  NAND2_X1   g04578(.A1(new_n4770_), .A2(new_n970_), .ZN(new_n4771_));
  AOI21_X1   g04579(.A1(new_n4767_), .A2(\asqrt[53] ), .B(new_n4771_), .ZN(new_n4772_));
  NOR2_X1    g04580(.A1(new_n4772_), .A2(new_n4766_), .ZN(new_n4773_));
  AOI22_X1   g04581(.A1(new_n4767_), .A2(\asqrt[53] ), .B1(new_n4765_), .B2(new_n4758_), .ZN(new_n4774_));
  NAND2_X1   g04582(.A1(new_n4551_), .A2(\asqrt[54] ), .ZN(new_n4775_));
  NOR4_X1    g04583(.A1(new_n4645_), .A2(\asqrt[54] ), .A3(new_n4442_), .A4(new_n4551_), .ZN(new_n4776_));
  XOR2_X1    g04584(.A1(new_n4776_), .A2(new_n4775_), .Z(new_n4777_));
  NAND2_X1   g04585(.A1(new_n4777_), .A2(new_n825_), .ZN(new_n4778_));
  INV_X1     g04586(.I(new_n4778_), .ZN(new_n4779_));
  OAI21_X1   g04587(.A1(new_n4774_), .A2(new_n970_), .B(new_n4779_), .ZN(new_n4780_));
  NAND2_X1   g04588(.A1(new_n4780_), .A2(new_n4773_), .ZN(new_n4781_));
  OAI22_X1   g04589(.A1(new_n4774_), .A2(new_n970_), .B1(new_n4772_), .B2(new_n4766_), .ZN(new_n4782_));
  NAND2_X1   g04590(.A1(new_n4453_), .A2(\asqrt[55] ), .ZN(new_n4783_));
  NOR4_X1    g04591(.A1(new_n4645_), .A2(\asqrt[55] ), .A3(new_n4448_), .A4(new_n4453_), .ZN(new_n4784_));
  XOR2_X1    g04592(.A1(new_n4784_), .A2(new_n4783_), .Z(new_n4785_));
  NAND2_X1   g04593(.A1(new_n4785_), .A2(new_n724_), .ZN(new_n4786_));
  AOI21_X1   g04594(.A1(new_n4782_), .A2(\asqrt[55] ), .B(new_n4786_), .ZN(new_n4787_));
  NOR2_X1    g04595(.A1(new_n4787_), .A2(new_n4781_), .ZN(new_n4788_));
  AOI22_X1   g04596(.A1(new_n4782_), .A2(\asqrt[55] ), .B1(new_n4780_), .B2(new_n4773_), .ZN(new_n4789_));
  NAND2_X1   g04597(.A1(new_n4558_), .A2(\asqrt[56] ), .ZN(new_n4790_));
  NOR4_X1    g04598(.A1(new_n4645_), .A2(\asqrt[56] ), .A3(new_n4455_), .A4(new_n4558_), .ZN(new_n4791_));
  XOR2_X1    g04599(.A1(new_n4791_), .A2(new_n4790_), .Z(new_n4792_));
  NAND2_X1   g04600(.A1(new_n4792_), .A2(new_n587_), .ZN(new_n4793_));
  INV_X1     g04601(.I(new_n4793_), .ZN(new_n4794_));
  OAI21_X1   g04602(.A1(new_n4789_), .A2(new_n724_), .B(new_n4794_), .ZN(new_n4795_));
  NAND2_X1   g04603(.A1(new_n4795_), .A2(new_n4788_), .ZN(new_n4796_));
  NAND2_X1   g04604(.A1(new_n4782_), .A2(\asqrt[55] ), .ZN(new_n4797_));
  AOI21_X1   g04605(.A1(new_n4797_), .A2(new_n4781_), .B(new_n724_), .ZN(new_n4798_));
  OAI21_X1   g04606(.A1(new_n4788_), .A2(new_n4798_), .B(\asqrt[57] ), .ZN(new_n4799_));
  NOR2_X1    g04607(.A1(new_n4561_), .A2(new_n587_), .ZN(new_n4800_));
  NOR4_X1    g04608(.A1(new_n4645_), .A2(\asqrt[57] ), .A3(new_n4461_), .A4(new_n4466_), .ZN(new_n4801_));
  XNOR2_X1   g04609(.A1(new_n4801_), .A2(new_n4800_), .ZN(new_n4802_));
  NAND2_X1   g04610(.A1(new_n4802_), .A2(new_n504_), .ZN(new_n4803_));
  INV_X1     g04611(.I(new_n4803_), .ZN(new_n4804_));
  AOI21_X1   g04612(.A1(new_n4799_), .A2(new_n4804_), .B(new_n4796_), .ZN(new_n4805_));
  OAI22_X1   g04613(.A1(new_n4789_), .A2(new_n724_), .B1(new_n4787_), .B2(new_n4781_), .ZN(new_n4806_));
  AOI22_X1   g04614(.A1(new_n4806_), .A2(\asqrt[57] ), .B1(new_n4795_), .B2(new_n4788_), .ZN(new_n4807_));
  NOR4_X1    g04615(.A1(new_n4645_), .A2(\asqrt[58] ), .A3(new_n4468_), .A4(new_n4565_), .ZN(new_n4808_));
  XOR2_X1    g04616(.A1(new_n4808_), .A2(new_n4609_), .Z(new_n4809_));
  NAND2_X1   g04617(.A1(new_n4809_), .A2(new_n376_), .ZN(new_n4810_));
  INV_X1     g04618(.I(new_n4810_), .ZN(new_n4811_));
  OAI21_X1   g04619(.A1(new_n4807_), .A2(new_n504_), .B(new_n4811_), .ZN(new_n4812_));
  NAND2_X1   g04620(.A1(new_n4812_), .A2(new_n4805_), .ZN(new_n4813_));
  AOI21_X1   g04621(.A1(new_n4796_), .A2(new_n4799_), .B(new_n504_), .ZN(new_n4814_));
  OAI21_X1   g04622(.A1(new_n4805_), .A2(new_n4814_), .B(\asqrt[59] ), .ZN(new_n4815_));
  NOR4_X1    g04623(.A1(new_n4645_), .A2(\asqrt[59] ), .A3(new_n4474_), .A4(new_n4479_), .ZN(new_n4816_));
  XOR2_X1    g04624(.A1(new_n4816_), .A2(new_n4587_), .Z(new_n4817_));
  AND2_X2    g04625(.A1(new_n4817_), .A2(new_n275_), .Z(new_n4818_));
  AOI21_X1   g04626(.A1(new_n4815_), .A2(new_n4818_), .B(new_n4813_), .ZN(new_n4819_));
  INV_X1     g04627(.I(new_n4674_), .ZN(new_n4820_));
  OAI21_X1   g04628(.A1(new_n4676_), .A2(new_n3760_), .B(new_n4820_), .ZN(new_n4821_));
  AOI22_X1   g04629(.A1(new_n4677_), .A2(\asqrt[42] ), .B1(new_n4821_), .B2(new_n4667_), .ZN(new_n4822_));
  INV_X1     g04630(.I(new_n4690_), .ZN(new_n4823_));
  OAI21_X1   g04631(.A1(new_n4822_), .A2(new_n3208_), .B(new_n4823_), .ZN(new_n4824_));
  OAI22_X1   g04632(.A1(new_n4822_), .A2(new_n3208_), .B1(new_n4683_), .B2(new_n4675_), .ZN(new_n4825_));
  AOI22_X1   g04633(.A1(new_n4825_), .A2(\asqrt[44] ), .B1(new_n4824_), .B2(new_n4694_), .ZN(new_n4826_));
  INV_X1     g04634(.I(new_n4708_), .ZN(new_n4827_));
  OAI21_X1   g04635(.A1(new_n4826_), .A2(new_n2728_), .B(new_n4827_), .ZN(new_n4828_));
  NAND2_X1   g04636(.A1(new_n4828_), .A2(new_n4711_), .ZN(new_n4829_));
  AOI21_X1   g04637(.A1(new_n4825_), .A2(\asqrt[44] ), .B(new_n4699_), .ZN(new_n4830_));
  OAI22_X1   g04638(.A1(new_n4826_), .A2(new_n2728_), .B1(new_n4830_), .B2(new_n4703_), .ZN(new_n4831_));
  AOI21_X1   g04639(.A1(new_n4831_), .A2(\asqrt[46] ), .B(new_n4717_), .ZN(new_n4832_));
  NOR2_X1    g04640(.A1(new_n4832_), .A2(new_n4829_), .ZN(new_n4833_));
  AOI22_X1   g04641(.A1(new_n4831_), .A2(\asqrt[46] ), .B1(new_n4828_), .B2(new_n4711_), .ZN(new_n4834_));
  INV_X1     g04642(.I(new_n4726_), .ZN(new_n4835_));
  OAI21_X1   g04643(.A1(new_n4834_), .A2(new_n2253_), .B(new_n4835_), .ZN(new_n4836_));
  NAND2_X1   g04644(.A1(new_n4836_), .A2(new_n4833_), .ZN(new_n4837_));
  OAI22_X1   g04645(.A1(new_n4834_), .A2(new_n2253_), .B1(new_n4832_), .B2(new_n4829_), .ZN(new_n4838_));
  AOI21_X1   g04646(.A1(new_n4838_), .A2(\asqrt[48] ), .B(new_n4733_), .ZN(new_n4839_));
  NOR2_X1    g04647(.A1(new_n4839_), .A2(new_n4837_), .ZN(new_n4840_));
  AOI22_X1   g04648(.A1(new_n4838_), .A2(\asqrt[48] ), .B1(new_n4836_), .B2(new_n4833_), .ZN(new_n4841_));
  INV_X1     g04649(.I(new_n4741_), .ZN(new_n4842_));
  OAI21_X1   g04650(.A1(new_n4841_), .A2(new_n1854_), .B(new_n4842_), .ZN(new_n4843_));
  NAND2_X1   g04651(.A1(new_n4843_), .A2(new_n4840_), .ZN(new_n4844_));
  OAI22_X1   g04652(.A1(new_n4841_), .A2(new_n1854_), .B1(new_n4839_), .B2(new_n4837_), .ZN(new_n4845_));
  AOI21_X1   g04653(.A1(new_n4845_), .A2(\asqrt[50] ), .B(new_n4748_), .ZN(new_n4846_));
  NOR2_X1    g04654(.A1(new_n4846_), .A2(new_n4844_), .ZN(new_n4847_));
  AOI22_X1   g04655(.A1(new_n4845_), .A2(\asqrt[50] ), .B1(new_n4843_), .B2(new_n4840_), .ZN(new_n4848_));
  INV_X1     g04656(.I(new_n4756_), .ZN(new_n4849_));
  OAI21_X1   g04657(.A1(new_n4848_), .A2(new_n1436_), .B(new_n4849_), .ZN(new_n4850_));
  NAND2_X1   g04658(.A1(new_n4850_), .A2(new_n4847_), .ZN(new_n4851_));
  OAI22_X1   g04659(.A1(new_n4848_), .A2(new_n1436_), .B1(new_n4846_), .B2(new_n4844_), .ZN(new_n4852_));
  AOI21_X1   g04660(.A1(new_n4852_), .A2(\asqrt[52] ), .B(new_n4763_), .ZN(new_n4853_));
  NOR2_X1    g04661(.A1(new_n4853_), .A2(new_n4851_), .ZN(new_n4854_));
  AOI22_X1   g04662(.A1(new_n4852_), .A2(\asqrt[52] ), .B1(new_n4850_), .B2(new_n4847_), .ZN(new_n4855_));
  INV_X1     g04663(.I(new_n4771_), .ZN(new_n4856_));
  OAI21_X1   g04664(.A1(new_n4855_), .A2(new_n1096_), .B(new_n4856_), .ZN(new_n4857_));
  NAND2_X1   g04665(.A1(new_n4857_), .A2(new_n4854_), .ZN(new_n4858_));
  OAI22_X1   g04666(.A1(new_n4855_), .A2(new_n1096_), .B1(new_n4853_), .B2(new_n4851_), .ZN(new_n4859_));
  AOI21_X1   g04667(.A1(new_n4859_), .A2(\asqrt[54] ), .B(new_n4778_), .ZN(new_n4860_));
  NOR2_X1    g04668(.A1(new_n4860_), .A2(new_n4858_), .ZN(new_n4861_));
  AOI22_X1   g04669(.A1(new_n4859_), .A2(\asqrt[54] ), .B1(new_n4857_), .B2(new_n4854_), .ZN(new_n4862_));
  INV_X1     g04670(.I(new_n4786_), .ZN(new_n4863_));
  OAI21_X1   g04671(.A1(new_n4862_), .A2(new_n825_), .B(new_n4863_), .ZN(new_n4864_));
  NAND2_X1   g04672(.A1(new_n4864_), .A2(new_n4861_), .ZN(new_n4865_));
  OAI22_X1   g04673(.A1(new_n4862_), .A2(new_n825_), .B1(new_n4860_), .B2(new_n4858_), .ZN(new_n4866_));
  AOI21_X1   g04674(.A1(new_n4866_), .A2(\asqrt[56] ), .B(new_n4793_), .ZN(new_n4867_));
  NOR2_X1    g04675(.A1(new_n4867_), .A2(new_n4865_), .ZN(new_n4868_));
  AOI22_X1   g04676(.A1(new_n4866_), .A2(\asqrt[56] ), .B1(new_n4864_), .B2(new_n4861_), .ZN(new_n4869_));
  OAI21_X1   g04677(.A1(new_n4869_), .A2(new_n587_), .B(new_n4804_), .ZN(new_n4870_));
  NAND2_X1   g04678(.A1(new_n4870_), .A2(new_n4868_), .ZN(new_n4871_));
  NAND2_X1   g04679(.A1(new_n4859_), .A2(\asqrt[54] ), .ZN(new_n4872_));
  AOI21_X1   g04680(.A1(new_n4872_), .A2(new_n4858_), .B(new_n825_), .ZN(new_n4873_));
  OAI21_X1   g04681(.A1(new_n4861_), .A2(new_n4873_), .B(\asqrt[56] ), .ZN(new_n4874_));
  AOI21_X1   g04682(.A1(new_n4865_), .A2(new_n4874_), .B(new_n587_), .ZN(new_n4875_));
  OAI21_X1   g04683(.A1(new_n4868_), .A2(new_n4875_), .B(\asqrt[58] ), .ZN(new_n4876_));
  NAND2_X1   g04684(.A1(new_n4871_), .A2(new_n4876_), .ZN(new_n4877_));
  AOI22_X1   g04685(.A1(new_n4877_), .A2(\asqrt[59] ), .B1(new_n4812_), .B2(new_n4805_), .ZN(new_n4878_));
  NOR4_X1    g04686(.A1(new_n4645_), .A2(\asqrt[60] ), .A3(new_n4481_), .A4(new_n4572_), .ZN(new_n4879_));
  XOR2_X1    g04687(.A1(new_n4879_), .A2(new_n4611_), .Z(new_n4880_));
  NAND2_X1   g04688(.A1(new_n4880_), .A2(new_n229_), .ZN(new_n4881_));
  INV_X1     g04689(.I(new_n4881_), .ZN(new_n4882_));
  OAI21_X1   g04690(.A1(new_n4878_), .A2(new_n275_), .B(new_n4882_), .ZN(new_n4883_));
  OAI22_X1   g04691(.A1(new_n4869_), .A2(new_n587_), .B1(new_n4867_), .B2(new_n4865_), .ZN(new_n4884_));
  AOI21_X1   g04692(.A1(new_n4884_), .A2(\asqrt[58] ), .B(new_n4810_), .ZN(new_n4885_));
  NOR2_X1    g04693(.A1(new_n4885_), .A2(new_n4871_), .ZN(new_n4886_));
  AOI22_X1   g04694(.A1(new_n4884_), .A2(\asqrt[58] ), .B1(new_n4870_), .B2(new_n4868_), .ZN(new_n4887_));
  OAI21_X1   g04695(.A1(new_n4887_), .A2(new_n376_), .B(new_n4818_), .ZN(new_n4888_));
  NAND2_X1   g04696(.A1(new_n4888_), .A2(new_n4886_), .ZN(new_n4889_));
  AOI21_X1   g04697(.A1(new_n4871_), .A2(new_n4876_), .B(new_n376_), .ZN(new_n4890_));
  OAI21_X1   g04698(.A1(new_n4886_), .A2(new_n4890_), .B(\asqrt[60] ), .ZN(new_n4891_));
  AOI21_X1   g04699(.A1(new_n4889_), .A2(new_n4891_), .B(new_n229_), .ZN(new_n4892_));
  INV_X1     g04700(.I(new_n4615_), .ZN(new_n4893_));
  NOR2_X1    g04701(.A1(new_n4893_), .A2(\asqrt[62] ), .ZN(new_n4894_));
  INV_X1     g04702(.I(new_n4894_), .ZN(new_n4895_));
  NAND4_X1   g04703(.A1(new_n4892_), .A2(new_n4819_), .A3(new_n4883_), .A4(new_n4895_), .ZN(new_n4896_));
  NAND2_X1   g04704(.A1(new_n4633_), .A2(new_n4583_), .ZN(new_n4897_));
  OAI21_X1   g04705(.A1(\asqrt[38] ), .A2(new_n4897_), .B(new_n4593_), .ZN(new_n4898_));
  NAND2_X1   g04706(.A1(new_n4898_), .A2(new_n231_), .ZN(new_n4899_));
  INV_X1     g04707(.I(new_n4899_), .ZN(new_n4900_));
  NAND3_X1   g04708(.A1(new_n4896_), .A2(new_n4617_), .A3(new_n4900_), .ZN(new_n4901_));
  OAI22_X1   g04709(.A1(new_n4887_), .A2(new_n376_), .B1(new_n4885_), .B2(new_n4871_), .ZN(new_n4902_));
  AOI21_X1   g04710(.A1(new_n4902_), .A2(\asqrt[60] ), .B(new_n4881_), .ZN(new_n4903_));
  AOI22_X1   g04711(.A1(new_n4902_), .A2(\asqrt[60] ), .B1(new_n4888_), .B2(new_n4886_), .ZN(new_n4904_));
  OAI22_X1   g04712(.A1(new_n4904_), .A2(new_n229_), .B1(new_n4903_), .B2(new_n4889_), .ZN(new_n4905_));
  NOR4_X1    g04713(.A1(new_n4905_), .A2(\asqrt[62] ), .A3(new_n4607_), .A4(new_n4615_), .ZN(new_n4906_));
  AOI21_X1   g04714(.A1(new_n4608_), .A2(new_n4901_), .B(new_n4906_), .ZN(new_n4907_));
  INV_X1     g04715(.I(\a[72] ), .ZN(new_n4908_));
  OAI21_X1   g04716(.A1(new_n4584_), .A2(new_n4593_), .B(\asqrt[38] ), .ZN(new_n4909_));
  XOR2_X1    g04717(.A1(new_n4593_), .A2(\asqrt[63] ), .Z(new_n4910_));
  NAND2_X1   g04718(.A1(new_n4909_), .A2(new_n4910_), .ZN(new_n4911_));
  INV_X1     g04719(.I(new_n4911_), .ZN(new_n4912_));
  NAND3_X1   g04720(.A1(new_n4639_), .A2(new_n4577_), .A3(new_n4584_), .ZN(new_n4913_));
  INV_X1     g04721(.I(new_n4913_), .ZN(new_n4914_));
  NOR2_X1    g04722(.A1(new_n4912_), .A2(new_n4914_), .ZN(new_n4915_));
  NOR2_X1    g04723(.A1(\a[70] ), .A2(\a[71] ), .ZN(new_n4916_));
  INV_X1     g04724(.I(new_n4916_), .ZN(new_n4917_));
  NOR3_X1    g04725(.A1(new_n4915_), .A2(new_n4908_), .A3(new_n4917_), .ZN(new_n4918_));
  NAND2_X1   g04726(.A1(new_n4907_), .A2(new_n4918_), .ZN(new_n4919_));
  XOR2_X1    g04727(.A1(new_n4919_), .A2(\a[73] ), .Z(new_n4920_));
  INV_X1     g04728(.I(\a[73] ), .ZN(new_n4921_));
  NAND2_X1   g04729(.A1(new_n4883_), .A2(new_n4819_), .ZN(new_n4922_));
  NAND2_X1   g04730(.A1(new_n4892_), .A2(new_n4895_), .ZN(new_n4923_));
  OAI21_X1   g04731(.A1(new_n4923_), .A2(new_n4922_), .B(new_n4617_), .ZN(new_n4924_));
  OAI21_X1   g04732(.A1(new_n4924_), .A2(new_n4899_), .B(new_n4608_), .ZN(new_n4925_));
  NAND2_X1   g04733(.A1(new_n4906_), .A2(new_n4912_), .ZN(new_n4926_));
  NOR2_X1    g04734(.A1(new_n4926_), .A2(new_n4925_), .ZN(new_n4927_));
  NAND3_X1   g04735(.A1(new_n4927_), .A2(new_n4608_), .A3(new_n4913_), .ZN(new_n4928_));
  NAND2_X1   g04736(.A1(new_n4889_), .A2(new_n4891_), .ZN(new_n4929_));
  AOI22_X1   g04737(.A1(new_n4929_), .A2(\asqrt[61] ), .B1(new_n4883_), .B2(new_n4819_), .ZN(new_n4930_));
  NOR2_X1    g04738(.A1(new_n4930_), .A2(new_n196_), .ZN(new_n4931_));
  AOI21_X1   g04739(.A1(new_n4813_), .A2(new_n4815_), .B(new_n275_), .ZN(new_n4932_));
  OAI21_X1   g04740(.A1(new_n4819_), .A2(new_n4932_), .B(\asqrt[61] ), .ZN(new_n4933_));
  NAND4_X1   g04741(.A1(new_n4922_), .A2(new_n196_), .A3(new_n4933_), .A4(new_n4893_), .ZN(new_n4934_));
  INV_X1     g04742(.I(new_n4934_), .ZN(new_n4935_));
  NOR3_X1    g04743(.A1(new_n4926_), .A2(new_n4925_), .A3(new_n4913_), .ZN(\asqrt[37] ));
  NAND3_X1   g04744(.A1(\asqrt[37] ), .A2(new_n4931_), .A3(new_n4935_), .ZN(new_n4937_));
  OAI21_X1   g04745(.A1(new_n4905_), .A2(\asqrt[62] ), .B(new_n4615_), .ZN(new_n4938_));
  OAI21_X1   g04746(.A1(\asqrt[37] ), .A2(new_n4938_), .B(new_n4931_), .ZN(new_n4939_));
  NAND2_X1   g04747(.A1(new_n4939_), .A2(new_n4937_), .ZN(new_n4940_));
  INV_X1     g04748(.I(new_n4940_), .ZN(new_n4941_));
  NOR3_X1    g04749(.A1(new_n4929_), .A2(\asqrt[61] ), .A3(new_n4880_), .ZN(new_n4942_));
  NAND2_X1   g04750(.A1(\asqrt[37] ), .A2(new_n4942_), .ZN(new_n4943_));
  XOR2_X1    g04751(.A1(new_n4943_), .A2(new_n4892_), .Z(new_n4944_));
  NOR2_X1    g04752(.A1(new_n4944_), .A2(new_n196_), .ZN(new_n4945_));
  INV_X1     g04753(.I(new_n4945_), .ZN(new_n4946_));
  INV_X1     g04754(.I(\a[74] ), .ZN(new_n4947_));
  NOR2_X1    g04755(.A1(\a[72] ), .A2(\a[73] ), .ZN(new_n4948_));
  INV_X1     g04756(.I(new_n4948_), .ZN(new_n4949_));
  NOR3_X1    g04757(.A1(new_n4646_), .A2(new_n4947_), .A3(new_n4949_), .ZN(new_n4950_));
  NAND3_X1   g04758(.A1(new_n4597_), .A2(new_n4633_), .A3(new_n4950_), .ZN(new_n4951_));
  XOR2_X1    g04759(.A1(new_n4951_), .A2(\a[75] ), .Z(new_n4952_));
  INV_X1     g04760(.I(\a[75] ), .ZN(new_n4953_));
  NOR4_X1    g04761(.A1(new_n4926_), .A2(new_n4925_), .A3(new_n4953_), .A4(new_n4913_), .ZN(new_n4954_));
  NOR2_X1    g04762(.A1(new_n4952_), .A2(\a[74] ), .ZN(new_n4955_));
  OAI21_X1   g04763(.A1(new_n4954_), .A2(new_n4955_), .B(new_n4952_), .ZN(new_n4956_));
  INV_X1     g04764(.I(new_n4952_), .ZN(new_n4957_));
  NOR2_X1    g04765(.A1(new_n4903_), .A2(new_n4889_), .ZN(new_n4958_));
  NOR3_X1    g04766(.A1(new_n4904_), .A2(new_n229_), .A3(new_n4894_), .ZN(new_n4959_));
  AOI21_X1   g04767(.A1(new_n4959_), .A2(new_n4958_), .B(new_n4616_), .ZN(new_n4960_));
  AOI21_X1   g04768(.A1(new_n4960_), .A2(new_n4900_), .B(new_n4607_), .ZN(new_n4961_));
  AOI21_X1   g04769(.A1(new_n4905_), .A2(\asqrt[62] ), .B(new_n4608_), .ZN(new_n4962_));
  NOR3_X1    g04770(.A1(new_n4962_), .A2(new_n4934_), .A3(new_n4911_), .ZN(new_n4963_));
  NAND4_X1   g04771(.A1(new_n4963_), .A2(\a[75] ), .A3(new_n4961_), .A4(new_n4914_), .ZN(new_n4964_));
  NAND3_X1   g04772(.A1(new_n4964_), .A2(\a[74] ), .A3(new_n4957_), .ZN(new_n4965_));
  NAND2_X1   g04773(.A1(new_n4956_), .A2(new_n4965_), .ZN(new_n4966_));
  NAND2_X1   g04774(.A1(new_n4631_), .A2(new_n4595_), .ZN(new_n4967_));
  NAND4_X1   g04775(.A1(new_n4635_), .A2(new_n4629_), .A3(new_n4584_), .A4(new_n4967_), .ZN(new_n4968_));
  NOR2_X1    g04776(.A1(new_n4645_), .A2(new_n4947_), .ZN(new_n4969_));
  XOR2_X1    g04777(.A1(new_n4969_), .A2(new_n4968_), .Z(new_n4970_));
  NOR2_X1    g04778(.A1(new_n4970_), .A2(new_n4949_), .ZN(new_n4971_));
  INV_X1     g04779(.I(new_n4971_), .ZN(new_n4972_));
  NAND3_X1   g04780(.A1(new_n4963_), .A2(new_n4961_), .A3(new_n4914_), .ZN(new_n4973_));
  NOR4_X1    g04781(.A1(new_n4933_), .A2(new_n4889_), .A3(new_n4903_), .A4(new_n4894_), .ZN(new_n4974_));
  NOR3_X1    g04782(.A1(new_n4974_), .A2(new_n4616_), .A3(new_n4899_), .ZN(new_n4975_));
  NAND4_X1   g04783(.A1(new_n4930_), .A2(new_n196_), .A3(new_n4608_), .A4(new_n4893_), .ZN(new_n4976_));
  OAI21_X1   g04784(.A1(new_n4975_), .A2(new_n4607_), .B(new_n4976_), .ZN(new_n4977_));
  NAND2_X1   g04785(.A1(new_n4915_), .A2(\asqrt[38] ), .ZN(new_n4978_));
  OAI21_X1   g04786(.A1(new_n4977_), .A2(new_n4978_), .B(new_n4618_), .ZN(new_n4979_));
  NAND3_X1   g04787(.A1(new_n4979_), .A2(new_n4619_), .A3(new_n4973_), .ZN(new_n4980_));
  INV_X1     g04788(.I(new_n4978_), .ZN(new_n4981_));
  AOI21_X1   g04789(.A1(new_n4907_), .A2(new_n4981_), .B(\a[76] ), .ZN(new_n4982_));
  OAI21_X1   g04790(.A1(new_n4982_), .A2(new_n4620_), .B(\asqrt[37] ), .ZN(new_n4983_));
  NAND4_X1   g04791(.A1(new_n4980_), .A2(new_n4983_), .A3(new_n4330_), .A4(new_n4972_), .ZN(new_n4984_));
  NAND2_X1   g04792(.A1(new_n4984_), .A2(new_n4966_), .ZN(new_n4985_));
  NAND3_X1   g04793(.A1(new_n4956_), .A2(new_n4965_), .A3(new_n4972_), .ZN(new_n4986_));
  AOI21_X1   g04794(.A1(\asqrt[38] ), .A2(new_n4618_), .B(\a[77] ), .ZN(new_n4987_));
  NOR2_X1    g04795(.A1(new_n4636_), .A2(\a[76] ), .ZN(new_n4988_));
  AOI21_X1   g04796(.A1(\asqrt[38] ), .A2(\a[76] ), .B(new_n4622_), .ZN(new_n4989_));
  OAI21_X1   g04797(.A1(new_n4987_), .A2(new_n4988_), .B(new_n4989_), .ZN(new_n4990_));
  INV_X1     g04798(.I(new_n4990_), .ZN(new_n4991_));
  NAND3_X1   g04799(.A1(\asqrt[37] ), .A2(new_n4644_), .A3(new_n4991_), .ZN(new_n4992_));
  OAI21_X1   g04800(.A1(new_n4973_), .A2(new_n4990_), .B(new_n4643_), .ZN(new_n4993_));
  NAND3_X1   g04801(.A1(new_n4992_), .A2(new_n4993_), .A3(new_n4018_), .ZN(new_n4994_));
  AOI21_X1   g04802(.A1(new_n4986_), .A2(\asqrt[39] ), .B(new_n4994_), .ZN(new_n4995_));
  NOR2_X1    g04803(.A1(new_n4985_), .A2(new_n4995_), .ZN(new_n4996_));
  AOI22_X1   g04804(.A1(new_n4984_), .A2(new_n4966_), .B1(\asqrt[39] ), .B2(new_n4986_), .ZN(new_n4997_));
  INV_X1     g04805(.I(new_n4626_), .ZN(new_n4998_));
  AOI21_X1   g04806(.A1(new_n4636_), .A2(new_n4998_), .B(new_n4628_), .ZN(new_n4999_));
  INV_X1     g04807(.I(new_n4637_), .ZN(new_n5000_));
  NOR3_X1    g04808(.A1(new_n5000_), .A2(new_n4999_), .A3(new_n4643_), .ZN(new_n5001_));
  AOI21_X1   g04809(.A1(new_n4654_), .A2(new_n4651_), .B(\asqrt[40] ), .ZN(new_n5002_));
  AND4_X2    g04810(.A1(new_n5001_), .A2(\asqrt[37] ), .A3(new_n4668_), .A4(new_n5002_), .Z(new_n5003_));
  NOR2_X1    g04811(.A1(new_n5001_), .A2(new_n4018_), .ZN(new_n5004_));
  NOR3_X1    g04812(.A1(new_n5003_), .A2(\asqrt[41] ), .A3(new_n5004_), .ZN(new_n5005_));
  OAI21_X1   g04813(.A1(new_n4997_), .A2(new_n4018_), .B(new_n5005_), .ZN(new_n5006_));
  NAND2_X1   g04814(.A1(new_n5006_), .A2(new_n4996_), .ZN(new_n5007_));
  OAI22_X1   g04815(.A1(new_n4997_), .A2(new_n4018_), .B1(new_n4985_), .B2(new_n4995_), .ZN(new_n5008_));
  NAND2_X1   g04816(.A1(new_n4662_), .A2(new_n4664_), .ZN(new_n5009_));
  NAND4_X1   g04817(.A1(\asqrt[37] ), .A2(new_n3760_), .A3(new_n5009_), .A4(new_n4676_), .ZN(new_n5010_));
  XOR2_X1    g04818(.A1(new_n5010_), .A2(new_n4669_), .Z(new_n5011_));
  NAND2_X1   g04819(.A1(new_n5011_), .A2(new_n3481_), .ZN(new_n5012_));
  AOI21_X1   g04820(.A1(new_n5008_), .A2(\asqrt[41] ), .B(new_n5012_), .ZN(new_n5013_));
  NOR2_X1    g04821(.A1(new_n5013_), .A2(new_n5007_), .ZN(new_n5014_));
  AOI22_X1   g04822(.A1(new_n5008_), .A2(\asqrt[41] ), .B1(new_n5006_), .B2(new_n4996_), .ZN(new_n5015_));
  NOR4_X1    g04823(.A1(new_n4973_), .A2(\asqrt[42] ), .A3(new_n4673_), .A4(new_n4677_), .ZN(new_n5016_));
  XOR2_X1    g04824(.A1(new_n5016_), .A2(new_n4684_), .Z(new_n5017_));
  NAND2_X1   g04825(.A1(new_n5017_), .A2(new_n3208_), .ZN(new_n5018_));
  INV_X1     g04826(.I(new_n5018_), .ZN(new_n5019_));
  OAI21_X1   g04827(.A1(new_n5015_), .A2(new_n3481_), .B(new_n5019_), .ZN(new_n5020_));
  NAND2_X1   g04828(.A1(new_n5020_), .A2(new_n5014_), .ZN(new_n5021_));
  OAI22_X1   g04829(.A1(new_n5015_), .A2(new_n3481_), .B1(new_n5013_), .B2(new_n5007_), .ZN(new_n5022_));
  NAND2_X1   g04830(.A1(new_n4675_), .A2(new_n4684_), .ZN(new_n5023_));
  NOR4_X1    g04831(.A1(new_n4973_), .A2(\asqrt[43] ), .A3(new_n4681_), .A4(new_n5023_), .ZN(new_n5024_));
  XNOR2_X1   g04832(.A1(new_n5024_), .A2(new_n4685_), .ZN(new_n5025_));
  NAND2_X1   g04833(.A1(new_n5025_), .A2(new_n2941_), .ZN(new_n5026_));
  AOI21_X1   g04834(.A1(new_n5022_), .A2(\asqrt[43] ), .B(new_n5026_), .ZN(new_n5027_));
  NOR2_X1    g04835(.A1(new_n5027_), .A2(new_n5021_), .ZN(new_n5028_));
  AOI22_X1   g04836(.A1(new_n5022_), .A2(\asqrt[43] ), .B1(new_n5020_), .B2(new_n5014_), .ZN(new_n5029_));
  NOR4_X1    g04837(.A1(new_n4973_), .A2(\asqrt[44] ), .A3(new_n4689_), .A4(new_n4825_), .ZN(new_n5030_));
  XOR2_X1    g04838(.A1(new_n5030_), .A2(new_n4695_), .Z(new_n5031_));
  NAND2_X1   g04839(.A1(new_n5031_), .A2(new_n2728_), .ZN(new_n5032_));
  INV_X1     g04840(.I(new_n5032_), .ZN(new_n5033_));
  OAI21_X1   g04841(.A1(new_n5029_), .A2(new_n2941_), .B(new_n5033_), .ZN(new_n5034_));
  NAND2_X1   g04842(.A1(new_n5034_), .A2(new_n5028_), .ZN(new_n5035_));
  OAI22_X1   g04843(.A1(new_n5029_), .A2(new_n2941_), .B1(new_n5027_), .B2(new_n5021_), .ZN(new_n5036_));
  NOR4_X1    g04844(.A1(new_n4973_), .A2(\asqrt[45] ), .A3(new_n4698_), .A4(new_n4704_), .ZN(new_n5037_));
  XNOR2_X1   g04845(.A1(new_n5037_), .A2(new_n4712_), .ZN(new_n5038_));
  NAND2_X1   g04846(.A1(new_n5038_), .A2(new_n2488_), .ZN(new_n5039_));
  AOI21_X1   g04847(.A1(new_n5036_), .A2(\asqrt[45] ), .B(new_n5039_), .ZN(new_n5040_));
  NOR2_X1    g04848(.A1(new_n5040_), .A2(new_n5035_), .ZN(new_n5041_));
  AOI22_X1   g04849(.A1(new_n5036_), .A2(\asqrt[45] ), .B1(new_n5034_), .B2(new_n5028_), .ZN(new_n5042_));
  NOR4_X1    g04850(.A1(new_n4973_), .A2(\asqrt[46] ), .A3(new_n4707_), .A4(new_n4831_), .ZN(new_n5043_));
  XOR2_X1    g04851(.A1(new_n5043_), .A2(new_n4713_), .Z(new_n5044_));
  NAND2_X1   g04852(.A1(new_n5044_), .A2(new_n2253_), .ZN(new_n5045_));
  INV_X1     g04853(.I(new_n5045_), .ZN(new_n5046_));
  OAI21_X1   g04854(.A1(new_n5042_), .A2(new_n2488_), .B(new_n5046_), .ZN(new_n5047_));
  NAND2_X1   g04855(.A1(new_n5047_), .A2(new_n5041_), .ZN(new_n5048_));
  OAI22_X1   g04856(.A1(new_n5042_), .A2(new_n2488_), .B1(new_n5040_), .B2(new_n5035_), .ZN(new_n5049_));
  NAND2_X1   g04857(.A1(new_n4722_), .A2(\asqrt[47] ), .ZN(new_n5050_));
  NOR4_X1    g04858(.A1(new_n4973_), .A2(\asqrt[47] ), .A3(new_n4716_), .A4(new_n4722_), .ZN(new_n5051_));
  XOR2_X1    g04859(.A1(new_n5051_), .A2(new_n5050_), .Z(new_n5052_));
  NAND2_X1   g04860(.A1(new_n5052_), .A2(new_n2046_), .ZN(new_n5053_));
  AOI21_X1   g04861(.A1(new_n5049_), .A2(\asqrt[47] ), .B(new_n5053_), .ZN(new_n5054_));
  NOR2_X1    g04862(.A1(new_n5054_), .A2(new_n5048_), .ZN(new_n5055_));
  AOI22_X1   g04863(.A1(new_n5049_), .A2(\asqrt[47] ), .B1(new_n5047_), .B2(new_n5041_), .ZN(new_n5056_));
  NAND2_X1   g04864(.A1(new_n4838_), .A2(\asqrt[48] ), .ZN(new_n5057_));
  NOR4_X1    g04865(.A1(new_n4973_), .A2(\asqrt[48] ), .A3(new_n4725_), .A4(new_n4838_), .ZN(new_n5058_));
  XOR2_X1    g04866(.A1(new_n5058_), .A2(new_n5057_), .Z(new_n5059_));
  NAND2_X1   g04867(.A1(new_n5059_), .A2(new_n1854_), .ZN(new_n5060_));
  INV_X1     g04868(.I(new_n5060_), .ZN(new_n5061_));
  OAI21_X1   g04869(.A1(new_n5056_), .A2(new_n2046_), .B(new_n5061_), .ZN(new_n5062_));
  NAND2_X1   g04870(.A1(new_n5062_), .A2(new_n5055_), .ZN(new_n5063_));
  OAI22_X1   g04871(.A1(new_n5056_), .A2(new_n2046_), .B1(new_n5054_), .B2(new_n5048_), .ZN(new_n5064_));
  NAND2_X1   g04872(.A1(new_n4737_), .A2(\asqrt[49] ), .ZN(new_n5065_));
  NOR4_X1    g04873(.A1(new_n4973_), .A2(\asqrt[49] ), .A3(new_n4732_), .A4(new_n4737_), .ZN(new_n5066_));
  XOR2_X1    g04874(.A1(new_n5066_), .A2(new_n5065_), .Z(new_n5067_));
  NAND2_X1   g04875(.A1(new_n5067_), .A2(new_n1595_), .ZN(new_n5068_));
  AOI21_X1   g04876(.A1(new_n5064_), .A2(\asqrt[49] ), .B(new_n5068_), .ZN(new_n5069_));
  NOR2_X1    g04877(.A1(new_n5069_), .A2(new_n5063_), .ZN(new_n5070_));
  AOI22_X1   g04878(.A1(new_n5064_), .A2(\asqrt[49] ), .B1(new_n5062_), .B2(new_n5055_), .ZN(new_n5071_));
  NAND2_X1   g04879(.A1(new_n4845_), .A2(\asqrt[50] ), .ZN(new_n5072_));
  NOR4_X1    g04880(.A1(new_n4973_), .A2(\asqrt[50] ), .A3(new_n4740_), .A4(new_n4845_), .ZN(new_n5073_));
  XOR2_X1    g04881(.A1(new_n5073_), .A2(new_n5072_), .Z(new_n5074_));
  NAND2_X1   g04882(.A1(new_n5074_), .A2(new_n1436_), .ZN(new_n5075_));
  INV_X1     g04883(.I(new_n5075_), .ZN(new_n5076_));
  OAI21_X1   g04884(.A1(new_n5071_), .A2(new_n1595_), .B(new_n5076_), .ZN(new_n5077_));
  NAND2_X1   g04885(.A1(new_n5077_), .A2(new_n5070_), .ZN(new_n5078_));
  OAI22_X1   g04886(.A1(new_n5071_), .A2(new_n1595_), .B1(new_n5069_), .B2(new_n5063_), .ZN(new_n5079_));
  NAND2_X1   g04887(.A1(new_n4752_), .A2(\asqrt[51] ), .ZN(new_n5080_));
  NOR4_X1    g04888(.A1(new_n4973_), .A2(\asqrt[51] ), .A3(new_n4747_), .A4(new_n4752_), .ZN(new_n5081_));
  XOR2_X1    g04889(.A1(new_n5081_), .A2(new_n5080_), .Z(new_n5082_));
  NAND2_X1   g04890(.A1(new_n5082_), .A2(new_n1260_), .ZN(new_n5083_));
  AOI21_X1   g04891(.A1(new_n5079_), .A2(\asqrt[51] ), .B(new_n5083_), .ZN(new_n5084_));
  NOR2_X1    g04892(.A1(new_n5084_), .A2(new_n5078_), .ZN(new_n5085_));
  AOI22_X1   g04893(.A1(new_n5079_), .A2(\asqrt[51] ), .B1(new_n5077_), .B2(new_n5070_), .ZN(new_n5086_));
  NAND2_X1   g04894(.A1(new_n4852_), .A2(\asqrt[52] ), .ZN(new_n5087_));
  NOR4_X1    g04895(.A1(new_n4973_), .A2(\asqrt[52] ), .A3(new_n4755_), .A4(new_n4852_), .ZN(new_n5088_));
  XOR2_X1    g04896(.A1(new_n5088_), .A2(new_n5087_), .Z(new_n5089_));
  NAND2_X1   g04897(.A1(new_n5089_), .A2(new_n1096_), .ZN(new_n5090_));
  INV_X1     g04898(.I(new_n5090_), .ZN(new_n5091_));
  OAI21_X1   g04899(.A1(new_n5086_), .A2(new_n1260_), .B(new_n5091_), .ZN(new_n5092_));
  NAND2_X1   g04900(.A1(new_n5092_), .A2(new_n5085_), .ZN(new_n5093_));
  OAI22_X1   g04901(.A1(new_n5086_), .A2(new_n1260_), .B1(new_n5084_), .B2(new_n5078_), .ZN(new_n5094_));
  NOR2_X1    g04902(.A1(new_n4855_), .A2(new_n1096_), .ZN(new_n5095_));
  NOR4_X1    g04903(.A1(new_n4973_), .A2(\asqrt[53] ), .A3(new_n4762_), .A4(new_n4767_), .ZN(new_n5096_));
  XNOR2_X1   g04904(.A1(new_n5096_), .A2(new_n5095_), .ZN(new_n5097_));
  NAND2_X1   g04905(.A1(new_n5097_), .A2(new_n970_), .ZN(new_n5098_));
  AOI21_X1   g04906(.A1(new_n5094_), .A2(\asqrt[53] ), .B(new_n5098_), .ZN(new_n5099_));
  NOR2_X1    g04907(.A1(new_n5099_), .A2(new_n5093_), .ZN(new_n5100_));
  AOI22_X1   g04908(.A1(new_n5094_), .A2(\asqrt[53] ), .B1(new_n5092_), .B2(new_n5085_), .ZN(new_n5101_));
  NOR4_X1    g04909(.A1(new_n4973_), .A2(\asqrt[54] ), .A3(new_n4770_), .A4(new_n4859_), .ZN(new_n5102_));
  XOR2_X1    g04910(.A1(new_n5102_), .A2(new_n4872_), .Z(new_n5103_));
  NAND2_X1   g04911(.A1(new_n5103_), .A2(new_n825_), .ZN(new_n5104_));
  INV_X1     g04912(.I(new_n5104_), .ZN(new_n5105_));
  OAI21_X1   g04913(.A1(new_n5101_), .A2(new_n970_), .B(new_n5105_), .ZN(new_n5106_));
  NAND2_X1   g04914(.A1(new_n5106_), .A2(new_n5100_), .ZN(new_n5107_));
  OAI22_X1   g04915(.A1(new_n5101_), .A2(new_n970_), .B1(new_n5099_), .B2(new_n5093_), .ZN(new_n5108_));
  NOR4_X1    g04916(.A1(new_n4973_), .A2(\asqrt[55] ), .A3(new_n4777_), .A4(new_n4782_), .ZN(new_n5109_));
  XOR2_X1    g04917(.A1(new_n5109_), .A2(new_n4797_), .Z(new_n5110_));
  NAND2_X1   g04918(.A1(new_n5110_), .A2(new_n724_), .ZN(new_n5111_));
  AOI21_X1   g04919(.A1(new_n5108_), .A2(\asqrt[55] ), .B(new_n5111_), .ZN(new_n5112_));
  NOR2_X1    g04920(.A1(new_n5112_), .A2(new_n5107_), .ZN(new_n5113_));
  AOI22_X1   g04921(.A1(new_n5108_), .A2(\asqrt[55] ), .B1(new_n5106_), .B2(new_n5100_), .ZN(new_n5114_));
  NOR4_X1    g04922(.A1(new_n4973_), .A2(\asqrt[56] ), .A3(new_n4785_), .A4(new_n4866_), .ZN(new_n5115_));
  XOR2_X1    g04923(.A1(new_n5115_), .A2(new_n4874_), .Z(new_n5116_));
  NAND2_X1   g04924(.A1(new_n5116_), .A2(new_n587_), .ZN(new_n5117_));
  INV_X1     g04925(.I(new_n5117_), .ZN(new_n5118_));
  OAI21_X1   g04926(.A1(new_n5114_), .A2(new_n724_), .B(new_n5118_), .ZN(new_n5119_));
  NAND2_X1   g04927(.A1(new_n5119_), .A2(new_n5113_), .ZN(new_n5120_));
  OAI22_X1   g04928(.A1(new_n5114_), .A2(new_n724_), .B1(new_n5112_), .B2(new_n5107_), .ZN(new_n5121_));
  NOR4_X1    g04929(.A1(new_n4973_), .A2(\asqrt[57] ), .A3(new_n4792_), .A4(new_n4806_), .ZN(new_n5122_));
  XOR2_X1    g04930(.A1(new_n5122_), .A2(new_n4799_), .Z(new_n5123_));
  NAND2_X1   g04931(.A1(new_n5123_), .A2(new_n504_), .ZN(new_n5124_));
  AOI21_X1   g04932(.A1(new_n5121_), .A2(\asqrt[57] ), .B(new_n5124_), .ZN(new_n5125_));
  NOR2_X1    g04933(.A1(new_n5125_), .A2(new_n5120_), .ZN(new_n5126_));
  AOI22_X1   g04934(.A1(new_n5121_), .A2(\asqrt[57] ), .B1(new_n5119_), .B2(new_n5113_), .ZN(new_n5127_));
  NOR4_X1    g04935(.A1(new_n4973_), .A2(\asqrt[58] ), .A3(new_n4802_), .A4(new_n4884_), .ZN(new_n5128_));
  XOR2_X1    g04936(.A1(new_n5128_), .A2(new_n4876_), .Z(new_n5129_));
  NAND2_X1   g04937(.A1(new_n5129_), .A2(new_n376_), .ZN(new_n5130_));
  INV_X1     g04938(.I(new_n5130_), .ZN(new_n5131_));
  OAI21_X1   g04939(.A1(new_n5127_), .A2(new_n504_), .B(new_n5131_), .ZN(new_n5132_));
  NAND2_X1   g04940(.A1(new_n5132_), .A2(new_n5126_), .ZN(new_n5133_));
  OAI22_X1   g04941(.A1(new_n5127_), .A2(new_n504_), .B1(new_n5125_), .B2(new_n5120_), .ZN(new_n5134_));
  NOR4_X1    g04942(.A1(new_n4973_), .A2(\asqrt[59] ), .A3(new_n4809_), .A4(new_n4877_), .ZN(new_n5135_));
  XOR2_X1    g04943(.A1(new_n5135_), .A2(new_n4815_), .Z(new_n5136_));
  NAND2_X1   g04944(.A1(new_n5136_), .A2(new_n275_), .ZN(new_n5137_));
  AOI21_X1   g04945(.A1(new_n5134_), .A2(\asqrt[59] ), .B(new_n5137_), .ZN(new_n5138_));
  NOR2_X1    g04946(.A1(new_n5138_), .A2(new_n5133_), .ZN(new_n5139_));
  AOI22_X1   g04947(.A1(new_n5134_), .A2(\asqrt[59] ), .B1(new_n5132_), .B2(new_n5126_), .ZN(new_n5140_));
  NOR4_X1    g04948(.A1(new_n4973_), .A2(\asqrt[60] ), .A3(new_n4817_), .A4(new_n4902_), .ZN(new_n5141_));
  XOR2_X1    g04949(.A1(new_n5141_), .A2(new_n4891_), .Z(new_n5142_));
  NAND2_X1   g04950(.A1(new_n5142_), .A2(new_n229_), .ZN(new_n5143_));
  INV_X1     g04951(.I(new_n5143_), .ZN(new_n5144_));
  OAI21_X1   g04952(.A1(new_n5140_), .A2(new_n275_), .B(new_n5144_), .ZN(new_n5145_));
  NAND2_X1   g04953(.A1(new_n5145_), .A2(new_n5139_), .ZN(new_n5146_));
  OAI22_X1   g04954(.A1(new_n5140_), .A2(new_n275_), .B1(new_n5138_), .B2(new_n5133_), .ZN(new_n5147_));
  INV_X1     g04955(.I(new_n4944_), .ZN(new_n5148_));
  NOR2_X1    g04956(.A1(new_n5148_), .A2(\asqrt[62] ), .ZN(new_n5149_));
  INV_X1     g04957(.I(new_n5149_), .ZN(new_n5150_));
  NAND3_X1   g04958(.A1(new_n5147_), .A2(\asqrt[61] ), .A3(new_n5150_), .ZN(new_n5151_));
  OAI21_X1   g04959(.A1(new_n5151_), .A2(new_n5146_), .B(new_n4946_), .ZN(new_n5152_));
  NAND3_X1   g04960(.A1(new_n4973_), .A2(new_n4607_), .A3(new_n4976_), .ZN(new_n5153_));
  AOI21_X1   g04961(.A1(new_n5153_), .A2(new_n4924_), .B(\asqrt[63] ), .ZN(new_n5154_));
  INV_X1     g04962(.I(new_n5154_), .ZN(new_n5155_));
  OAI21_X1   g04963(.A1(new_n5152_), .A2(new_n5155_), .B(new_n4941_), .ZN(new_n5156_));
  INV_X1     g04964(.I(new_n4955_), .ZN(new_n5157_));
  AOI21_X1   g04965(.A1(new_n4964_), .A2(new_n5157_), .B(new_n4957_), .ZN(new_n5158_));
  NOR3_X1    g04966(.A1(new_n4954_), .A2(new_n4947_), .A3(new_n4952_), .ZN(new_n5159_));
  NOR2_X1    g04967(.A1(new_n5159_), .A2(new_n5158_), .ZN(new_n5160_));
  NOR3_X1    g04968(.A1(new_n4982_), .A2(new_n4620_), .A3(\asqrt[37] ), .ZN(new_n5161_));
  AOI21_X1   g04969(.A1(new_n4979_), .A2(new_n4619_), .B(new_n4973_), .ZN(new_n5162_));
  NOR4_X1    g04970(.A1(new_n5162_), .A2(new_n5161_), .A3(\asqrt[39] ), .A4(new_n4971_), .ZN(new_n5163_));
  NOR2_X1    g04971(.A1(new_n5163_), .A2(new_n5160_), .ZN(new_n5164_));
  NOR3_X1    g04972(.A1(new_n5159_), .A2(new_n5158_), .A3(new_n4971_), .ZN(new_n5165_));
  NOR3_X1    g04973(.A1(new_n4973_), .A2(new_n4643_), .A3(new_n4990_), .ZN(new_n5166_));
  AOI21_X1   g04974(.A1(\asqrt[37] ), .A2(new_n4991_), .B(new_n4644_), .ZN(new_n5167_));
  NOR3_X1    g04975(.A1(new_n5167_), .A2(new_n5166_), .A3(\asqrt[40] ), .ZN(new_n5168_));
  OAI21_X1   g04976(.A1(new_n5165_), .A2(new_n4330_), .B(new_n5168_), .ZN(new_n5169_));
  NAND2_X1   g04977(.A1(new_n5164_), .A2(new_n5169_), .ZN(new_n5170_));
  OAI22_X1   g04978(.A1(new_n5163_), .A2(new_n5160_), .B1(new_n4330_), .B2(new_n5165_), .ZN(new_n5171_));
  INV_X1     g04979(.I(new_n5005_), .ZN(new_n5172_));
  AOI21_X1   g04980(.A1(new_n5171_), .A2(\asqrt[40] ), .B(new_n5172_), .ZN(new_n5173_));
  NOR2_X1    g04981(.A1(new_n5173_), .A2(new_n5170_), .ZN(new_n5174_));
  AOI22_X1   g04982(.A1(new_n5171_), .A2(\asqrt[40] ), .B1(new_n5164_), .B2(new_n5169_), .ZN(new_n5175_));
  INV_X1     g04983(.I(new_n5012_), .ZN(new_n5176_));
  OAI21_X1   g04984(.A1(new_n5175_), .A2(new_n3760_), .B(new_n5176_), .ZN(new_n5177_));
  NAND2_X1   g04985(.A1(new_n5177_), .A2(new_n5174_), .ZN(new_n5178_));
  OAI22_X1   g04986(.A1(new_n5175_), .A2(new_n3760_), .B1(new_n5173_), .B2(new_n5170_), .ZN(new_n5179_));
  AOI21_X1   g04987(.A1(new_n5179_), .A2(\asqrt[42] ), .B(new_n5018_), .ZN(new_n5180_));
  NOR2_X1    g04988(.A1(new_n5180_), .A2(new_n5178_), .ZN(new_n5181_));
  AOI22_X1   g04989(.A1(new_n5179_), .A2(\asqrt[42] ), .B1(new_n5177_), .B2(new_n5174_), .ZN(new_n5182_));
  INV_X1     g04990(.I(new_n5026_), .ZN(new_n5183_));
  OAI21_X1   g04991(.A1(new_n5182_), .A2(new_n3208_), .B(new_n5183_), .ZN(new_n5184_));
  NAND2_X1   g04992(.A1(new_n5184_), .A2(new_n5181_), .ZN(new_n5185_));
  OAI22_X1   g04993(.A1(new_n5182_), .A2(new_n3208_), .B1(new_n5180_), .B2(new_n5178_), .ZN(new_n5186_));
  AOI21_X1   g04994(.A1(new_n5186_), .A2(\asqrt[44] ), .B(new_n5032_), .ZN(new_n5187_));
  NOR2_X1    g04995(.A1(new_n5187_), .A2(new_n5185_), .ZN(new_n5188_));
  AOI22_X1   g04996(.A1(new_n5186_), .A2(\asqrt[44] ), .B1(new_n5184_), .B2(new_n5181_), .ZN(new_n5189_));
  INV_X1     g04997(.I(new_n5039_), .ZN(new_n5190_));
  OAI21_X1   g04998(.A1(new_n5189_), .A2(new_n2728_), .B(new_n5190_), .ZN(new_n5191_));
  NAND2_X1   g04999(.A1(new_n5191_), .A2(new_n5188_), .ZN(new_n5192_));
  OAI22_X1   g05000(.A1(new_n5189_), .A2(new_n2728_), .B1(new_n5187_), .B2(new_n5185_), .ZN(new_n5193_));
  AOI21_X1   g05001(.A1(new_n5193_), .A2(\asqrt[46] ), .B(new_n5045_), .ZN(new_n5194_));
  NOR2_X1    g05002(.A1(new_n5194_), .A2(new_n5192_), .ZN(new_n5195_));
  AOI22_X1   g05003(.A1(new_n5193_), .A2(\asqrt[46] ), .B1(new_n5191_), .B2(new_n5188_), .ZN(new_n5196_));
  INV_X1     g05004(.I(new_n5053_), .ZN(new_n5197_));
  OAI21_X1   g05005(.A1(new_n5196_), .A2(new_n2253_), .B(new_n5197_), .ZN(new_n5198_));
  NAND2_X1   g05006(.A1(new_n5198_), .A2(new_n5195_), .ZN(new_n5199_));
  OAI22_X1   g05007(.A1(new_n5196_), .A2(new_n2253_), .B1(new_n5194_), .B2(new_n5192_), .ZN(new_n5200_));
  AOI21_X1   g05008(.A1(new_n5200_), .A2(\asqrt[48] ), .B(new_n5060_), .ZN(new_n5201_));
  NOR2_X1    g05009(.A1(new_n5201_), .A2(new_n5199_), .ZN(new_n5202_));
  AOI22_X1   g05010(.A1(new_n5200_), .A2(\asqrt[48] ), .B1(new_n5198_), .B2(new_n5195_), .ZN(new_n5203_));
  INV_X1     g05011(.I(new_n5068_), .ZN(new_n5204_));
  OAI21_X1   g05012(.A1(new_n5203_), .A2(new_n1854_), .B(new_n5204_), .ZN(new_n5205_));
  NAND2_X1   g05013(.A1(new_n5205_), .A2(new_n5202_), .ZN(new_n5206_));
  OAI22_X1   g05014(.A1(new_n5203_), .A2(new_n1854_), .B1(new_n5201_), .B2(new_n5199_), .ZN(new_n5207_));
  AOI21_X1   g05015(.A1(new_n5207_), .A2(\asqrt[50] ), .B(new_n5075_), .ZN(new_n5208_));
  NOR2_X1    g05016(.A1(new_n5208_), .A2(new_n5206_), .ZN(new_n5209_));
  AOI22_X1   g05017(.A1(new_n5207_), .A2(\asqrt[50] ), .B1(new_n5205_), .B2(new_n5202_), .ZN(new_n5210_));
  INV_X1     g05018(.I(new_n5083_), .ZN(new_n5211_));
  OAI21_X1   g05019(.A1(new_n5210_), .A2(new_n1436_), .B(new_n5211_), .ZN(new_n5212_));
  NAND2_X1   g05020(.A1(new_n5212_), .A2(new_n5209_), .ZN(new_n5213_));
  OAI22_X1   g05021(.A1(new_n5210_), .A2(new_n1436_), .B1(new_n5208_), .B2(new_n5206_), .ZN(new_n5214_));
  AOI21_X1   g05022(.A1(new_n5214_), .A2(\asqrt[52] ), .B(new_n5090_), .ZN(new_n5215_));
  NOR2_X1    g05023(.A1(new_n5215_), .A2(new_n5213_), .ZN(new_n5216_));
  AOI22_X1   g05024(.A1(new_n5214_), .A2(\asqrt[52] ), .B1(new_n5212_), .B2(new_n5209_), .ZN(new_n5217_));
  INV_X1     g05025(.I(new_n5098_), .ZN(new_n5218_));
  OAI21_X1   g05026(.A1(new_n5217_), .A2(new_n1096_), .B(new_n5218_), .ZN(new_n5219_));
  NAND2_X1   g05027(.A1(new_n5219_), .A2(new_n5216_), .ZN(new_n5220_));
  OAI22_X1   g05028(.A1(new_n5217_), .A2(new_n1096_), .B1(new_n5215_), .B2(new_n5213_), .ZN(new_n5221_));
  AOI21_X1   g05029(.A1(new_n5221_), .A2(\asqrt[54] ), .B(new_n5104_), .ZN(new_n5222_));
  NOR2_X1    g05030(.A1(new_n5222_), .A2(new_n5220_), .ZN(new_n5223_));
  AOI22_X1   g05031(.A1(new_n5221_), .A2(\asqrt[54] ), .B1(new_n5219_), .B2(new_n5216_), .ZN(new_n5224_));
  INV_X1     g05032(.I(new_n5111_), .ZN(new_n5225_));
  OAI21_X1   g05033(.A1(new_n5224_), .A2(new_n825_), .B(new_n5225_), .ZN(new_n5226_));
  NAND2_X1   g05034(.A1(new_n5226_), .A2(new_n5223_), .ZN(new_n5227_));
  OAI22_X1   g05035(.A1(new_n5224_), .A2(new_n825_), .B1(new_n5222_), .B2(new_n5220_), .ZN(new_n5228_));
  AOI21_X1   g05036(.A1(new_n5228_), .A2(\asqrt[56] ), .B(new_n5117_), .ZN(new_n5229_));
  NOR2_X1    g05037(.A1(new_n5229_), .A2(new_n5227_), .ZN(new_n5230_));
  AOI22_X1   g05038(.A1(new_n5228_), .A2(\asqrt[56] ), .B1(new_n5226_), .B2(new_n5223_), .ZN(new_n5231_));
  INV_X1     g05039(.I(new_n5124_), .ZN(new_n5232_));
  OAI21_X1   g05040(.A1(new_n5231_), .A2(new_n587_), .B(new_n5232_), .ZN(new_n5233_));
  NAND2_X1   g05041(.A1(new_n5233_), .A2(new_n5230_), .ZN(new_n5234_));
  OAI22_X1   g05042(.A1(new_n5231_), .A2(new_n587_), .B1(new_n5229_), .B2(new_n5227_), .ZN(new_n5235_));
  AOI21_X1   g05043(.A1(new_n5235_), .A2(\asqrt[58] ), .B(new_n5130_), .ZN(new_n5236_));
  NOR2_X1    g05044(.A1(new_n5236_), .A2(new_n5234_), .ZN(new_n5237_));
  AOI22_X1   g05045(.A1(new_n5235_), .A2(\asqrt[58] ), .B1(new_n5233_), .B2(new_n5230_), .ZN(new_n5238_));
  INV_X1     g05046(.I(new_n5137_), .ZN(new_n5239_));
  OAI21_X1   g05047(.A1(new_n5238_), .A2(new_n376_), .B(new_n5239_), .ZN(new_n5240_));
  NAND2_X1   g05048(.A1(new_n5240_), .A2(new_n5237_), .ZN(new_n5241_));
  OAI22_X1   g05049(.A1(new_n5238_), .A2(new_n376_), .B1(new_n5236_), .B2(new_n5234_), .ZN(new_n5242_));
  AOI21_X1   g05050(.A1(new_n5242_), .A2(\asqrt[60] ), .B(new_n5143_), .ZN(new_n5243_));
  AOI22_X1   g05051(.A1(new_n5242_), .A2(\asqrt[60] ), .B1(new_n5240_), .B2(new_n5237_), .ZN(new_n5244_));
  OAI22_X1   g05052(.A1(new_n5244_), .A2(new_n229_), .B1(new_n5243_), .B2(new_n5241_), .ZN(new_n5245_));
  NOR4_X1    g05053(.A1(new_n5245_), .A2(\asqrt[62] ), .A3(new_n4940_), .A4(new_n4944_), .ZN(new_n5246_));
  NAND2_X1   g05054(.A1(new_n4960_), .A2(new_n4607_), .ZN(new_n5247_));
  XOR2_X1    g05055(.A1(new_n4960_), .A2(\asqrt[63] ), .Z(new_n5248_));
  AOI21_X1   g05056(.A1(\asqrt[37] ), .A2(new_n5247_), .B(new_n5248_), .ZN(new_n5249_));
  NAND2_X1   g05057(.A1(new_n5246_), .A2(new_n5249_), .ZN(new_n5250_));
  NOR4_X1    g05058(.A1(new_n5250_), .A2(new_n4921_), .A3(new_n4928_), .A4(new_n5156_), .ZN(new_n5251_));
  NOR2_X1    g05059(.A1(new_n4921_), .A2(\a[72] ), .ZN(new_n5252_));
  OAI21_X1   g05060(.A1(new_n5251_), .A2(new_n5252_), .B(new_n4920_), .ZN(new_n5253_));
  INV_X1     g05061(.I(new_n4920_), .ZN(new_n5254_));
  INV_X1     g05062(.I(new_n4928_), .ZN(new_n5255_));
  NOR2_X1    g05063(.A1(new_n5243_), .A2(new_n5241_), .ZN(new_n5256_));
  NOR3_X1    g05064(.A1(new_n5244_), .A2(new_n229_), .A3(new_n5149_), .ZN(new_n5257_));
  AOI21_X1   g05065(.A1(new_n5257_), .A2(new_n5256_), .B(new_n4945_), .ZN(new_n5258_));
  AOI21_X1   g05066(.A1(new_n5258_), .A2(new_n5154_), .B(new_n4940_), .ZN(new_n5259_));
  AOI22_X1   g05067(.A1(new_n5147_), .A2(\asqrt[61] ), .B1(new_n5145_), .B2(new_n5139_), .ZN(new_n5260_));
  NAND4_X1   g05068(.A1(new_n5260_), .A2(new_n196_), .A3(new_n4941_), .A4(new_n5148_), .ZN(new_n5261_));
  INV_X1     g05069(.I(new_n5249_), .ZN(new_n5262_));
  NOR2_X1    g05070(.A1(new_n5261_), .A2(new_n5262_), .ZN(new_n5263_));
  NAND4_X1   g05071(.A1(new_n5263_), .A2(new_n5259_), .A3(\a[73] ), .A4(new_n5255_), .ZN(new_n5264_));
  NAND3_X1   g05072(.A1(new_n5264_), .A2(\a[72] ), .A3(new_n5254_), .ZN(new_n5265_));
  NAND2_X1   g05073(.A1(new_n5253_), .A2(new_n5265_), .ZN(new_n5266_));
  NOR2_X1    g05074(.A1(new_n5250_), .A2(new_n5156_), .ZN(new_n5267_));
  NOR4_X1    g05075(.A1(new_n4926_), .A2(new_n4607_), .A3(new_n4975_), .A4(new_n4913_), .ZN(new_n5268_));
  NAND2_X1   g05076(.A1(\asqrt[37] ), .A2(\a[72] ), .ZN(new_n5269_));
  XOR2_X1    g05077(.A1(new_n5269_), .A2(new_n5268_), .Z(new_n5270_));
  NOR2_X1    g05078(.A1(new_n5270_), .A2(new_n4917_), .ZN(new_n5271_));
  INV_X1     g05079(.I(new_n5271_), .ZN(new_n5272_));
  NAND3_X1   g05080(.A1(new_n5263_), .A2(new_n5259_), .A3(new_n5255_), .ZN(new_n5273_));
  NAND2_X1   g05081(.A1(new_n5121_), .A2(\asqrt[57] ), .ZN(new_n5274_));
  AOI21_X1   g05082(.A1(new_n5274_), .A2(new_n5120_), .B(new_n504_), .ZN(new_n5275_));
  OAI21_X1   g05083(.A1(new_n5126_), .A2(new_n5275_), .B(\asqrt[59] ), .ZN(new_n5276_));
  AOI21_X1   g05084(.A1(new_n5133_), .A2(new_n5276_), .B(new_n275_), .ZN(new_n5277_));
  OAI21_X1   g05085(.A1(new_n5139_), .A2(new_n5277_), .B(\asqrt[61] ), .ZN(new_n5278_));
  NOR3_X1    g05086(.A1(new_n5146_), .A2(new_n5278_), .A3(new_n5149_), .ZN(new_n5279_));
  NOR3_X1    g05087(.A1(new_n5279_), .A2(new_n4945_), .A3(new_n5155_), .ZN(new_n5280_));
  OAI21_X1   g05088(.A1(new_n5280_), .A2(new_n4940_), .B(new_n5261_), .ZN(new_n5281_));
  NOR2_X1    g05089(.A1(new_n5255_), .A2(new_n5249_), .ZN(new_n5282_));
  NAND2_X1   g05090(.A1(new_n5282_), .A2(\asqrt[37] ), .ZN(new_n5283_));
  OAI21_X1   g05091(.A1(new_n5281_), .A2(new_n5283_), .B(new_n4947_), .ZN(new_n5284_));
  NAND3_X1   g05092(.A1(new_n5284_), .A2(new_n4948_), .A3(new_n5273_), .ZN(new_n5285_));
  NOR4_X1    g05093(.A1(new_n5156_), .A2(new_n4928_), .A3(new_n5261_), .A4(new_n5262_), .ZN(\asqrt[36] ));
  NAND2_X1   g05094(.A1(new_n5221_), .A2(\asqrt[54] ), .ZN(new_n5287_));
  AOI21_X1   g05095(.A1(new_n5287_), .A2(new_n5220_), .B(new_n825_), .ZN(new_n5288_));
  OAI21_X1   g05096(.A1(new_n5223_), .A2(new_n5288_), .B(\asqrt[56] ), .ZN(new_n5289_));
  AOI21_X1   g05097(.A1(new_n5227_), .A2(new_n5289_), .B(new_n587_), .ZN(new_n5290_));
  OAI21_X1   g05098(.A1(new_n5230_), .A2(new_n5290_), .B(\asqrt[58] ), .ZN(new_n5291_));
  AOI21_X1   g05099(.A1(new_n5234_), .A2(new_n5291_), .B(new_n376_), .ZN(new_n5292_));
  OAI21_X1   g05100(.A1(new_n5237_), .A2(new_n5292_), .B(\asqrt[60] ), .ZN(new_n5293_));
  AOI21_X1   g05101(.A1(new_n5241_), .A2(new_n5293_), .B(new_n229_), .ZN(new_n5294_));
  NAND4_X1   g05102(.A1(new_n5294_), .A2(new_n5139_), .A3(new_n5145_), .A4(new_n5150_), .ZN(new_n5295_));
  NAND3_X1   g05103(.A1(new_n5295_), .A2(new_n4946_), .A3(new_n5154_), .ZN(new_n5296_));
  AOI21_X1   g05104(.A1(new_n4941_), .A2(new_n5296_), .B(new_n5246_), .ZN(new_n5297_));
  INV_X1     g05105(.I(new_n5283_), .ZN(new_n5298_));
  AOI21_X1   g05106(.A1(new_n5297_), .A2(new_n5298_), .B(\a[74] ), .ZN(new_n5299_));
  OAI21_X1   g05107(.A1(new_n5299_), .A2(new_n4949_), .B(\asqrt[36] ), .ZN(new_n5300_));
  NAND4_X1   g05108(.A1(new_n5300_), .A2(new_n5285_), .A3(new_n4645_), .A4(new_n5272_), .ZN(new_n5301_));
  NAND2_X1   g05109(.A1(new_n5301_), .A2(new_n5266_), .ZN(new_n5302_));
  NAND3_X1   g05110(.A1(new_n5253_), .A2(new_n5265_), .A3(new_n5272_), .ZN(new_n5303_));
  AOI21_X1   g05111(.A1(\asqrt[37] ), .A2(new_n4947_), .B(\a[75] ), .ZN(new_n5304_));
  NOR2_X1    g05112(.A1(new_n4964_), .A2(\a[74] ), .ZN(new_n5305_));
  AOI21_X1   g05113(.A1(\asqrt[37] ), .A2(\a[74] ), .B(new_n4951_), .ZN(new_n5306_));
  OAI21_X1   g05114(.A1(new_n5305_), .A2(new_n5304_), .B(new_n5306_), .ZN(new_n5307_));
  INV_X1     g05115(.I(new_n5307_), .ZN(new_n5308_));
  NAND3_X1   g05116(.A1(\asqrt[36] ), .A2(new_n4972_), .A3(new_n5308_), .ZN(new_n5309_));
  OAI21_X1   g05117(.A1(new_n5273_), .A2(new_n5307_), .B(new_n4971_), .ZN(new_n5310_));
  NAND3_X1   g05118(.A1(new_n5310_), .A2(new_n5309_), .A3(new_n4330_), .ZN(new_n5311_));
  AOI21_X1   g05119(.A1(new_n5303_), .A2(\asqrt[38] ), .B(new_n5311_), .ZN(new_n5312_));
  NOR2_X1    g05120(.A1(new_n5302_), .A2(new_n5312_), .ZN(new_n5313_));
  NAND2_X1   g05121(.A1(new_n5303_), .A2(\asqrt[38] ), .ZN(new_n5314_));
  AOI21_X1   g05122(.A1(new_n5302_), .A2(new_n5314_), .B(new_n4330_), .ZN(new_n5315_));
  NAND2_X1   g05123(.A1(new_n4986_), .A2(\asqrt[39] ), .ZN(new_n5316_));
  NAND2_X1   g05124(.A1(new_n4980_), .A2(new_n4983_), .ZN(new_n5317_));
  NAND3_X1   g05125(.A1(new_n5317_), .A2(new_n5165_), .A3(new_n4330_), .ZN(new_n5318_));
  NOR2_X1    g05126(.A1(new_n5273_), .A2(new_n5318_), .ZN(new_n5319_));
  AND2_X2    g05127(.A1(new_n5319_), .A2(new_n5316_), .Z(new_n5320_));
  NOR2_X1    g05128(.A1(new_n5319_), .A2(new_n5316_), .ZN(new_n5321_));
  NOR3_X1    g05129(.A1(new_n5320_), .A2(\asqrt[40] ), .A3(new_n5321_), .ZN(new_n5322_));
  INV_X1     g05130(.I(new_n5322_), .ZN(new_n5323_));
  OAI21_X1   g05131(.A1(new_n5315_), .A2(new_n5323_), .B(new_n5313_), .ZN(new_n5324_));
  OAI21_X1   g05132(.A1(new_n5315_), .A2(new_n5313_), .B(\asqrt[40] ), .ZN(new_n5325_));
  NOR2_X1    g05133(.A1(new_n5167_), .A2(new_n5166_), .ZN(new_n5326_));
  NOR4_X1    g05134(.A1(new_n5273_), .A2(\asqrt[40] ), .A3(new_n5326_), .A4(new_n5171_), .ZN(new_n5327_));
  AOI21_X1   g05135(.A1(new_n4985_), .A2(new_n5316_), .B(new_n4018_), .ZN(new_n5328_));
  NOR2_X1    g05136(.A1(new_n5327_), .A2(new_n5328_), .ZN(new_n5329_));
  NAND2_X1   g05137(.A1(new_n5329_), .A2(new_n3760_), .ZN(new_n5330_));
  INV_X1     g05138(.I(new_n5330_), .ZN(new_n5331_));
  AOI21_X1   g05139(.A1(new_n5325_), .A2(new_n5331_), .B(new_n5324_), .ZN(new_n5332_));
  AOI21_X1   g05140(.A1(new_n5324_), .A2(new_n5325_), .B(new_n3760_), .ZN(new_n5333_));
  NAND2_X1   g05141(.A1(new_n5008_), .A2(\asqrt[41] ), .ZN(new_n5334_));
  NOR2_X1    g05142(.A1(new_n5003_), .A2(new_n5004_), .ZN(new_n5335_));
  NOR4_X1    g05143(.A1(new_n5273_), .A2(\asqrt[41] ), .A3(new_n5335_), .A4(new_n5008_), .ZN(new_n5336_));
  XOR2_X1    g05144(.A1(new_n5336_), .A2(new_n5334_), .Z(new_n5337_));
  NAND2_X1   g05145(.A1(new_n5337_), .A2(new_n3481_), .ZN(new_n5338_));
  OAI21_X1   g05146(.A1(new_n5333_), .A2(new_n5338_), .B(new_n5332_), .ZN(new_n5339_));
  OAI21_X1   g05147(.A1(new_n5332_), .A2(new_n5333_), .B(\asqrt[42] ), .ZN(new_n5340_));
  NOR4_X1    g05148(.A1(new_n5273_), .A2(\asqrt[42] ), .A3(new_n5011_), .A4(new_n5179_), .ZN(new_n5341_));
  AOI21_X1   g05149(.A1(new_n5334_), .A2(new_n5007_), .B(new_n3481_), .ZN(new_n5342_));
  NOR2_X1    g05150(.A1(new_n5341_), .A2(new_n5342_), .ZN(new_n5343_));
  NAND2_X1   g05151(.A1(new_n5343_), .A2(new_n3208_), .ZN(new_n5344_));
  INV_X1     g05152(.I(new_n5344_), .ZN(new_n5345_));
  AOI21_X1   g05153(.A1(new_n5340_), .A2(new_n5345_), .B(new_n5339_), .ZN(new_n5346_));
  AOI22_X1   g05154(.A1(new_n5301_), .A2(new_n5266_), .B1(\asqrt[38] ), .B2(new_n5303_), .ZN(new_n5347_));
  OAI21_X1   g05155(.A1(new_n5347_), .A2(new_n4330_), .B(new_n5322_), .ZN(new_n5348_));
  OAI22_X1   g05156(.A1(new_n5347_), .A2(new_n4330_), .B1(new_n5302_), .B2(new_n5312_), .ZN(new_n5349_));
  AOI22_X1   g05157(.A1(new_n5349_), .A2(\asqrt[40] ), .B1(new_n5348_), .B2(new_n5313_), .ZN(new_n5350_));
  INV_X1     g05158(.I(new_n5338_), .ZN(new_n5351_));
  OAI21_X1   g05159(.A1(new_n5350_), .A2(new_n3760_), .B(new_n5351_), .ZN(new_n5352_));
  AOI21_X1   g05160(.A1(new_n5349_), .A2(\asqrt[40] ), .B(new_n5330_), .ZN(new_n5353_));
  OAI22_X1   g05161(.A1(new_n5350_), .A2(new_n3760_), .B1(new_n5353_), .B2(new_n5324_), .ZN(new_n5354_));
  AOI22_X1   g05162(.A1(new_n5354_), .A2(\asqrt[42] ), .B1(new_n5352_), .B2(new_n5332_), .ZN(new_n5355_));
  NAND2_X1   g05163(.A1(new_n5022_), .A2(\asqrt[43] ), .ZN(new_n5356_));
  NOR4_X1    g05164(.A1(new_n5273_), .A2(\asqrt[43] ), .A3(new_n5017_), .A4(new_n5022_), .ZN(new_n5357_));
  XOR2_X1    g05165(.A1(new_n5357_), .A2(new_n5356_), .Z(new_n5358_));
  NAND2_X1   g05166(.A1(new_n5358_), .A2(new_n2941_), .ZN(new_n5359_));
  INV_X1     g05167(.I(new_n5359_), .ZN(new_n5360_));
  OAI21_X1   g05168(.A1(new_n5355_), .A2(new_n3208_), .B(new_n5360_), .ZN(new_n5361_));
  NAND2_X1   g05169(.A1(new_n5361_), .A2(new_n5346_), .ZN(new_n5362_));
  AOI21_X1   g05170(.A1(new_n5354_), .A2(\asqrt[42] ), .B(new_n5344_), .ZN(new_n5363_));
  OAI22_X1   g05171(.A1(new_n5355_), .A2(new_n3208_), .B1(new_n5363_), .B2(new_n5339_), .ZN(new_n5364_));
  NOR4_X1    g05172(.A1(new_n5273_), .A2(\asqrt[44] ), .A3(new_n5025_), .A4(new_n5186_), .ZN(new_n5365_));
  AOI21_X1   g05173(.A1(new_n5356_), .A2(new_n5021_), .B(new_n2941_), .ZN(new_n5366_));
  NOR2_X1    g05174(.A1(new_n5365_), .A2(new_n5366_), .ZN(new_n5367_));
  NAND2_X1   g05175(.A1(new_n5367_), .A2(new_n2728_), .ZN(new_n5368_));
  AOI21_X1   g05176(.A1(new_n5364_), .A2(\asqrt[44] ), .B(new_n5368_), .ZN(new_n5369_));
  NOR2_X1    g05177(.A1(new_n5369_), .A2(new_n5362_), .ZN(new_n5370_));
  AOI22_X1   g05178(.A1(new_n5364_), .A2(\asqrt[44] ), .B1(new_n5361_), .B2(new_n5346_), .ZN(new_n5371_));
  NAND2_X1   g05179(.A1(new_n5036_), .A2(\asqrt[45] ), .ZN(new_n5372_));
  NOR4_X1    g05180(.A1(new_n5273_), .A2(\asqrt[45] ), .A3(new_n5031_), .A4(new_n5036_), .ZN(new_n5373_));
  XOR2_X1    g05181(.A1(new_n5373_), .A2(new_n5372_), .Z(new_n5374_));
  NAND2_X1   g05182(.A1(new_n5374_), .A2(new_n2488_), .ZN(new_n5375_));
  INV_X1     g05183(.I(new_n5375_), .ZN(new_n5376_));
  OAI21_X1   g05184(.A1(new_n5371_), .A2(new_n2728_), .B(new_n5376_), .ZN(new_n5377_));
  NAND2_X1   g05185(.A1(new_n5377_), .A2(new_n5370_), .ZN(new_n5378_));
  OAI22_X1   g05186(.A1(new_n5371_), .A2(new_n2728_), .B1(new_n5369_), .B2(new_n5362_), .ZN(new_n5379_));
  NOR4_X1    g05187(.A1(new_n5273_), .A2(\asqrt[46] ), .A3(new_n5038_), .A4(new_n5193_), .ZN(new_n5380_));
  AOI21_X1   g05188(.A1(new_n5372_), .A2(new_n5035_), .B(new_n2488_), .ZN(new_n5381_));
  NOR2_X1    g05189(.A1(new_n5380_), .A2(new_n5381_), .ZN(new_n5382_));
  NAND2_X1   g05190(.A1(new_n5382_), .A2(new_n2253_), .ZN(new_n5383_));
  AOI21_X1   g05191(.A1(new_n5379_), .A2(\asqrt[46] ), .B(new_n5383_), .ZN(new_n5384_));
  NOR2_X1    g05192(.A1(new_n5384_), .A2(new_n5378_), .ZN(new_n5385_));
  AOI22_X1   g05193(.A1(new_n5379_), .A2(\asqrt[46] ), .B1(new_n5377_), .B2(new_n5370_), .ZN(new_n5386_));
  NAND2_X1   g05194(.A1(new_n5049_), .A2(\asqrt[47] ), .ZN(new_n5387_));
  NOR4_X1    g05195(.A1(new_n5273_), .A2(\asqrt[47] ), .A3(new_n5044_), .A4(new_n5049_), .ZN(new_n5388_));
  XOR2_X1    g05196(.A1(new_n5388_), .A2(new_n5387_), .Z(new_n5389_));
  NAND2_X1   g05197(.A1(new_n5389_), .A2(new_n2046_), .ZN(new_n5390_));
  INV_X1     g05198(.I(new_n5390_), .ZN(new_n5391_));
  OAI21_X1   g05199(.A1(new_n5386_), .A2(new_n2253_), .B(new_n5391_), .ZN(new_n5392_));
  NAND2_X1   g05200(.A1(new_n5392_), .A2(new_n5385_), .ZN(new_n5393_));
  OAI22_X1   g05201(.A1(new_n5386_), .A2(new_n2253_), .B1(new_n5384_), .B2(new_n5378_), .ZN(new_n5394_));
  NAND2_X1   g05202(.A1(new_n5200_), .A2(\asqrt[48] ), .ZN(new_n5395_));
  NOR4_X1    g05203(.A1(new_n5273_), .A2(\asqrt[48] ), .A3(new_n5052_), .A4(new_n5200_), .ZN(new_n5396_));
  XOR2_X1    g05204(.A1(new_n5396_), .A2(new_n5395_), .Z(new_n5397_));
  NAND2_X1   g05205(.A1(new_n5397_), .A2(new_n1854_), .ZN(new_n5398_));
  AOI21_X1   g05206(.A1(new_n5394_), .A2(\asqrt[48] ), .B(new_n5398_), .ZN(new_n5399_));
  NOR2_X1    g05207(.A1(new_n5399_), .A2(new_n5393_), .ZN(new_n5400_));
  AOI22_X1   g05208(.A1(new_n5394_), .A2(\asqrt[48] ), .B1(new_n5392_), .B2(new_n5385_), .ZN(new_n5401_));
  NOR4_X1    g05209(.A1(new_n5273_), .A2(\asqrt[49] ), .A3(new_n5059_), .A4(new_n5064_), .ZN(new_n5402_));
  AOI21_X1   g05210(.A1(new_n5395_), .A2(new_n5199_), .B(new_n1854_), .ZN(new_n5403_));
  NOR2_X1    g05211(.A1(new_n5402_), .A2(new_n5403_), .ZN(new_n5404_));
  NAND2_X1   g05212(.A1(new_n5404_), .A2(new_n1595_), .ZN(new_n5405_));
  INV_X1     g05213(.I(new_n5405_), .ZN(new_n5406_));
  OAI21_X1   g05214(.A1(new_n5401_), .A2(new_n1854_), .B(new_n5406_), .ZN(new_n5407_));
  NAND2_X1   g05215(.A1(new_n5407_), .A2(new_n5400_), .ZN(new_n5408_));
  OAI22_X1   g05216(.A1(new_n5401_), .A2(new_n1854_), .B1(new_n5399_), .B2(new_n5393_), .ZN(new_n5409_));
  NAND2_X1   g05217(.A1(new_n5207_), .A2(\asqrt[50] ), .ZN(new_n5410_));
  NOR4_X1    g05218(.A1(new_n5273_), .A2(\asqrt[50] ), .A3(new_n5067_), .A4(new_n5207_), .ZN(new_n5411_));
  XOR2_X1    g05219(.A1(new_n5411_), .A2(new_n5410_), .Z(new_n5412_));
  NAND2_X1   g05220(.A1(new_n5412_), .A2(new_n1436_), .ZN(new_n5413_));
  AOI21_X1   g05221(.A1(new_n5409_), .A2(\asqrt[50] ), .B(new_n5413_), .ZN(new_n5414_));
  NOR2_X1    g05222(.A1(new_n5414_), .A2(new_n5408_), .ZN(new_n5415_));
  AOI22_X1   g05223(.A1(new_n5409_), .A2(\asqrt[50] ), .B1(new_n5407_), .B2(new_n5400_), .ZN(new_n5416_));
  NOR4_X1    g05224(.A1(new_n5273_), .A2(\asqrt[51] ), .A3(new_n5074_), .A4(new_n5079_), .ZN(new_n5417_));
  AOI21_X1   g05225(.A1(new_n5410_), .A2(new_n5206_), .B(new_n1436_), .ZN(new_n5418_));
  NOR2_X1    g05226(.A1(new_n5417_), .A2(new_n5418_), .ZN(new_n5419_));
  NAND2_X1   g05227(.A1(new_n5419_), .A2(new_n1260_), .ZN(new_n5420_));
  INV_X1     g05228(.I(new_n5420_), .ZN(new_n5421_));
  OAI21_X1   g05229(.A1(new_n5416_), .A2(new_n1436_), .B(new_n5421_), .ZN(new_n5422_));
  NAND2_X1   g05230(.A1(new_n5422_), .A2(new_n5415_), .ZN(new_n5423_));
  OAI22_X1   g05231(.A1(new_n5416_), .A2(new_n1436_), .B1(new_n5414_), .B2(new_n5408_), .ZN(new_n5424_));
  NAND2_X1   g05232(.A1(new_n5214_), .A2(\asqrt[52] ), .ZN(new_n5425_));
  NOR4_X1    g05233(.A1(new_n5273_), .A2(\asqrt[52] ), .A3(new_n5082_), .A4(new_n5214_), .ZN(new_n5426_));
  XOR2_X1    g05234(.A1(new_n5426_), .A2(new_n5425_), .Z(new_n5427_));
  NAND2_X1   g05235(.A1(new_n5427_), .A2(new_n1096_), .ZN(new_n5428_));
  AOI21_X1   g05236(.A1(new_n5424_), .A2(\asqrt[52] ), .B(new_n5428_), .ZN(new_n5429_));
  NOR2_X1    g05237(.A1(new_n5429_), .A2(new_n5423_), .ZN(new_n5430_));
  AOI22_X1   g05238(.A1(new_n5424_), .A2(\asqrt[52] ), .B1(new_n5422_), .B2(new_n5415_), .ZN(new_n5431_));
  NOR4_X1    g05239(.A1(new_n5273_), .A2(\asqrt[53] ), .A3(new_n5089_), .A4(new_n5094_), .ZN(new_n5432_));
  AOI21_X1   g05240(.A1(new_n5425_), .A2(new_n5213_), .B(new_n1096_), .ZN(new_n5433_));
  NOR2_X1    g05241(.A1(new_n5432_), .A2(new_n5433_), .ZN(new_n5434_));
  NAND2_X1   g05242(.A1(new_n5434_), .A2(new_n970_), .ZN(new_n5435_));
  INV_X1     g05243(.I(new_n5435_), .ZN(new_n5436_));
  OAI21_X1   g05244(.A1(new_n5431_), .A2(new_n1096_), .B(new_n5436_), .ZN(new_n5437_));
  NAND2_X1   g05245(.A1(new_n5437_), .A2(new_n5430_), .ZN(new_n5438_));
  OAI22_X1   g05246(.A1(new_n5431_), .A2(new_n1096_), .B1(new_n5429_), .B2(new_n5423_), .ZN(new_n5439_));
  NOR4_X1    g05247(.A1(new_n5273_), .A2(\asqrt[54] ), .A3(new_n5097_), .A4(new_n5221_), .ZN(new_n5440_));
  XOR2_X1    g05248(.A1(new_n5440_), .A2(new_n5287_), .Z(new_n5441_));
  NAND2_X1   g05249(.A1(new_n5441_), .A2(new_n825_), .ZN(new_n5442_));
  AOI21_X1   g05250(.A1(new_n5439_), .A2(\asqrt[54] ), .B(new_n5442_), .ZN(new_n5443_));
  NOR2_X1    g05251(.A1(new_n5443_), .A2(new_n5438_), .ZN(new_n5444_));
  AOI22_X1   g05252(.A1(new_n5439_), .A2(\asqrt[54] ), .B1(new_n5437_), .B2(new_n5430_), .ZN(new_n5445_));
  NOR4_X1    g05253(.A1(new_n5273_), .A2(\asqrt[55] ), .A3(new_n5103_), .A4(new_n5108_), .ZN(new_n5446_));
  XNOR2_X1   g05254(.A1(new_n5446_), .A2(new_n5288_), .ZN(new_n5447_));
  NAND2_X1   g05255(.A1(new_n5447_), .A2(new_n724_), .ZN(new_n5448_));
  INV_X1     g05256(.I(new_n5448_), .ZN(new_n5449_));
  OAI21_X1   g05257(.A1(new_n5445_), .A2(new_n825_), .B(new_n5449_), .ZN(new_n5450_));
  NAND2_X1   g05258(.A1(new_n5450_), .A2(new_n5444_), .ZN(new_n5451_));
  OAI22_X1   g05259(.A1(new_n5445_), .A2(new_n825_), .B1(new_n5443_), .B2(new_n5438_), .ZN(new_n5452_));
  NOR4_X1    g05260(.A1(new_n5273_), .A2(\asqrt[56] ), .A3(new_n5110_), .A4(new_n5228_), .ZN(new_n5453_));
  XOR2_X1    g05261(.A1(new_n5453_), .A2(new_n5289_), .Z(new_n5454_));
  NAND2_X1   g05262(.A1(new_n5454_), .A2(new_n587_), .ZN(new_n5455_));
  AOI21_X1   g05263(.A1(new_n5452_), .A2(\asqrt[56] ), .B(new_n5455_), .ZN(new_n5456_));
  NOR2_X1    g05264(.A1(new_n5456_), .A2(new_n5451_), .ZN(new_n5457_));
  AOI22_X1   g05265(.A1(new_n5452_), .A2(\asqrt[56] ), .B1(new_n5450_), .B2(new_n5444_), .ZN(new_n5458_));
  NOR4_X1    g05266(.A1(new_n5273_), .A2(\asqrt[57] ), .A3(new_n5116_), .A4(new_n5121_), .ZN(new_n5459_));
  XOR2_X1    g05267(.A1(new_n5459_), .A2(new_n5274_), .Z(new_n5460_));
  NAND2_X1   g05268(.A1(new_n5460_), .A2(new_n504_), .ZN(new_n5461_));
  INV_X1     g05269(.I(new_n5461_), .ZN(new_n5462_));
  OAI21_X1   g05270(.A1(new_n5458_), .A2(new_n587_), .B(new_n5462_), .ZN(new_n5463_));
  NAND2_X1   g05271(.A1(new_n5463_), .A2(new_n5457_), .ZN(new_n5464_));
  OAI22_X1   g05272(.A1(new_n5458_), .A2(new_n587_), .B1(new_n5456_), .B2(new_n5451_), .ZN(new_n5465_));
  NOR4_X1    g05273(.A1(new_n5273_), .A2(\asqrt[58] ), .A3(new_n5123_), .A4(new_n5235_), .ZN(new_n5466_));
  XOR2_X1    g05274(.A1(new_n5466_), .A2(new_n5291_), .Z(new_n5467_));
  NAND2_X1   g05275(.A1(new_n5467_), .A2(new_n376_), .ZN(new_n5468_));
  AOI21_X1   g05276(.A1(new_n5465_), .A2(\asqrt[58] ), .B(new_n5468_), .ZN(new_n5469_));
  NOR2_X1    g05277(.A1(new_n5469_), .A2(new_n5464_), .ZN(new_n5470_));
  AOI22_X1   g05278(.A1(new_n5465_), .A2(\asqrt[58] ), .B1(new_n5463_), .B2(new_n5457_), .ZN(new_n5471_));
  NOR4_X1    g05279(.A1(new_n5273_), .A2(\asqrt[59] ), .A3(new_n5129_), .A4(new_n5134_), .ZN(new_n5472_));
  XOR2_X1    g05280(.A1(new_n5472_), .A2(new_n5276_), .Z(new_n5473_));
  AND2_X2    g05281(.A1(new_n5473_), .A2(new_n275_), .Z(new_n5474_));
  OAI21_X1   g05282(.A1(new_n5471_), .A2(new_n376_), .B(new_n5474_), .ZN(new_n5475_));
  NAND2_X1   g05283(.A1(new_n5475_), .A2(new_n5470_), .ZN(new_n5476_));
  NAND2_X1   g05284(.A1(new_n5452_), .A2(\asqrt[56] ), .ZN(new_n5477_));
  AOI21_X1   g05285(.A1(new_n5477_), .A2(new_n5451_), .B(new_n587_), .ZN(new_n5478_));
  OAI21_X1   g05286(.A1(new_n5457_), .A2(new_n5478_), .B(\asqrt[58] ), .ZN(new_n5479_));
  AOI21_X1   g05287(.A1(new_n5464_), .A2(new_n5479_), .B(new_n376_), .ZN(new_n5480_));
  OAI21_X1   g05288(.A1(new_n5470_), .A2(new_n5480_), .B(\asqrt[60] ), .ZN(new_n5481_));
  AOI21_X1   g05289(.A1(new_n5476_), .A2(new_n5481_), .B(new_n229_), .ZN(new_n5482_));
  NOR2_X1    g05290(.A1(new_n5260_), .A2(new_n196_), .ZN(new_n5483_));
  NOR2_X1    g05291(.A1(new_n5245_), .A2(\asqrt[62] ), .ZN(new_n5484_));
  NAND3_X1   g05292(.A1(new_n5484_), .A2(new_n5483_), .A3(new_n5148_), .ZN(new_n5485_));
  NOR2_X1    g05293(.A1(new_n5273_), .A2(new_n5485_), .ZN(new_n5486_));
  OR3_X2     g05294(.A1(\asqrt[36] ), .A2(new_n5148_), .A3(new_n5484_), .Z(new_n5487_));
  AOI21_X1   g05295(.A1(new_n5487_), .A2(new_n5483_), .B(new_n5486_), .ZN(new_n5488_));
  NOR4_X1    g05296(.A1(new_n5273_), .A2(\asqrt[61] ), .A3(new_n5142_), .A4(new_n5147_), .ZN(new_n5489_));
  XOR2_X1    g05297(.A1(new_n5489_), .A2(new_n5278_), .Z(new_n5490_));
  NOR2_X1    g05298(.A1(new_n5490_), .A2(new_n196_), .ZN(new_n5491_));
  INV_X1     g05299(.I(new_n5491_), .ZN(new_n5492_));
  NOR2_X1    g05300(.A1(new_n5333_), .A2(new_n5338_), .ZN(new_n5493_));
  NOR3_X1    g05301(.A1(new_n5493_), .A2(new_n5324_), .A3(new_n5353_), .ZN(new_n5494_));
  NAND2_X1   g05302(.A1(new_n5340_), .A2(new_n5345_), .ZN(new_n5495_));
  NAND2_X1   g05303(.A1(new_n5495_), .A2(new_n5494_), .ZN(new_n5496_));
  NAND2_X1   g05304(.A1(new_n5339_), .A2(new_n5340_), .ZN(new_n5497_));
  AOI21_X1   g05305(.A1(new_n5497_), .A2(\asqrt[43] ), .B(new_n5359_), .ZN(new_n5498_));
  NOR2_X1    g05306(.A1(new_n5498_), .A2(new_n5496_), .ZN(new_n5499_));
  AOI21_X1   g05307(.A1(new_n5339_), .A2(new_n5340_), .B(new_n3208_), .ZN(new_n5500_));
  OAI21_X1   g05308(.A1(new_n5346_), .A2(new_n5500_), .B(\asqrt[44] ), .ZN(new_n5501_));
  INV_X1     g05309(.I(new_n5368_), .ZN(new_n5502_));
  NAND2_X1   g05310(.A1(new_n5501_), .A2(new_n5502_), .ZN(new_n5503_));
  NAND2_X1   g05311(.A1(new_n5503_), .A2(new_n5499_), .ZN(new_n5504_));
  AOI22_X1   g05312(.A1(new_n5497_), .A2(\asqrt[43] ), .B1(new_n5495_), .B2(new_n5494_), .ZN(new_n5505_));
  OAI22_X1   g05313(.A1(new_n5505_), .A2(new_n2941_), .B1(new_n5498_), .B2(new_n5496_), .ZN(new_n5506_));
  AOI21_X1   g05314(.A1(new_n5506_), .A2(\asqrt[45] ), .B(new_n5375_), .ZN(new_n5507_));
  NOR2_X1    g05315(.A1(new_n5507_), .A2(new_n5504_), .ZN(new_n5508_));
  AOI22_X1   g05316(.A1(new_n5506_), .A2(\asqrt[45] ), .B1(new_n5503_), .B2(new_n5499_), .ZN(new_n5509_));
  INV_X1     g05317(.I(new_n5383_), .ZN(new_n5510_));
  OAI21_X1   g05318(.A1(new_n5509_), .A2(new_n2488_), .B(new_n5510_), .ZN(new_n5511_));
  NAND2_X1   g05319(.A1(new_n5511_), .A2(new_n5508_), .ZN(new_n5512_));
  OAI22_X1   g05320(.A1(new_n5509_), .A2(new_n2488_), .B1(new_n5507_), .B2(new_n5504_), .ZN(new_n5513_));
  AOI21_X1   g05321(.A1(new_n5513_), .A2(\asqrt[47] ), .B(new_n5390_), .ZN(new_n5514_));
  NOR2_X1    g05322(.A1(new_n5514_), .A2(new_n5512_), .ZN(new_n5515_));
  AOI22_X1   g05323(.A1(new_n5513_), .A2(\asqrt[47] ), .B1(new_n5511_), .B2(new_n5508_), .ZN(new_n5516_));
  INV_X1     g05324(.I(new_n5398_), .ZN(new_n5517_));
  OAI21_X1   g05325(.A1(new_n5516_), .A2(new_n2046_), .B(new_n5517_), .ZN(new_n5518_));
  NAND2_X1   g05326(.A1(new_n5518_), .A2(new_n5515_), .ZN(new_n5519_));
  OAI22_X1   g05327(.A1(new_n5516_), .A2(new_n2046_), .B1(new_n5514_), .B2(new_n5512_), .ZN(new_n5520_));
  AOI21_X1   g05328(.A1(new_n5520_), .A2(\asqrt[49] ), .B(new_n5405_), .ZN(new_n5521_));
  NOR2_X1    g05329(.A1(new_n5521_), .A2(new_n5519_), .ZN(new_n5522_));
  AOI22_X1   g05330(.A1(new_n5520_), .A2(\asqrt[49] ), .B1(new_n5518_), .B2(new_n5515_), .ZN(new_n5523_));
  INV_X1     g05331(.I(new_n5413_), .ZN(new_n5524_));
  OAI21_X1   g05332(.A1(new_n5523_), .A2(new_n1595_), .B(new_n5524_), .ZN(new_n5525_));
  NAND2_X1   g05333(.A1(new_n5525_), .A2(new_n5522_), .ZN(new_n5526_));
  OAI22_X1   g05334(.A1(new_n5523_), .A2(new_n1595_), .B1(new_n5521_), .B2(new_n5519_), .ZN(new_n5527_));
  AOI21_X1   g05335(.A1(new_n5527_), .A2(\asqrt[51] ), .B(new_n5420_), .ZN(new_n5528_));
  NOR2_X1    g05336(.A1(new_n5528_), .A2(new_n5526_), .ZN(new_n5529_));
  AOI22_X1   g05337(.A1(new_n5527_), .A2(\asqrt[51] ), .B1(new_n5525_), .B2(new_n5522_), .ZN(new_n5530_));
  INV_X1     g05338(.I(new_n5428_), .ZN(new_n5531_));
  OAI21_X1   g05339(.A1(new_n5530_), .A2(new_n1260_), .B(new_n5531_), .ZN(new_n5532_));
  NAND2_X1   g05340(.A1(new_n5532_), .A2(new_n5529_), .ZN(new_n5533_));
  OAI22_X1   g05341(.A1(new_n5530_), .A2(new_n1260_), .B1(new_n5528_), .B2(new_n5526_), .ZN(new_n5534_));
  AOI21_X1   g05342(.A1(new_n5534_), .A2(\asqrt[53] ), .B(new_n5435_), .ZN(new_n5535_));
  NOR2_X1    g05343(.A1(new_n5535_), .A2(new_n5533_), .ZN(new_n5536_));
  AOI22_X1   g05344(.A1(new_n5534_), .A2(\asqrt[53] ), .B1(new_n5532_), .B2(new_n5529_), .ZN(new_n5537_));
  INV_X1     g05345(.I(new_n5442_), .ZN(new_n5538_));
  OAI21_X1   g05346(.A1(new_n5537_), .A2(new_n970_), .B(new_n5538_), .ZN(new_n5539_));
  NAND2_X1   g05347(.A1(new_n5539_), .A2(new_n5536_), .ZN(new_n5540_));
  OAI22_X1   g05348(.A1(new_n5537_), .A2(new_n970_), .B1(new_n5535_), .B2(new_n5533_), .ZN(new_n5541_));
  AOI21_X1   g05349(.A1(new_n5541_), .A2(\asqrt[55] ), .B(new_n5448_), .ZN(new_n5542_));
  NOR2_X1    g05350(.A1(new_n5542_), .A2(new_n5540_), .ZN(new_n5543_));
  AOI22_X1   g05351(.A1(new_n5541_), .A2(\asqrt[55] ), .B1(new_n5539_), .B2(new_n5536_), .ZN(new_n5544_));
  INV_X1     g05352(.I(new_n5455_), .ZN(new_n5545_));
  OAI21_X1   g05353(.A1(new_n5544_), .A2(new_n724_), .B(new_n5545_), .ZN(new_n5546_));
  NAND2_X1   g05354(.A1(new_n5546_), .A2(new_n5543_), .ZN(new_n5547_));
  OAI22_X1   g05355(.A1(new_n5544_), .A2(new_n724_), .B1(new_n5542_), .B2(new_n5540_), .ZN(new_n5548_));
  AOI21_X1   g05356(.A1(new_n5548_), .A2(\asqrt[57] ), .B(new_n5461_), .ZN(new_n5549_));
  NOR2_X1    g05357(.A1(new_n5549_), .A2(new_n5547_), .ZN(new_n5550_));
  AOI22_X1   g05358(.A1(new_n5548_), .A2(\asqrt[57] ), .B1(new_n5546_), .B2(new_n5543_), .ZN(new_n5551_));
  INV_X1     g05359(.I(new_n5468_), .ZN(new_n5552_));
  OAI21_X1   g05360(.A1(new_n5551_), .A2(new_n504_), .B(new_n5552_), .ZN(new_n5553_));
  NAND2_X1   g05361(.A1(new_n5553_), .A2(new_n5550_), .ZN(new_n5554_));
  NAND2_X1   g05362(.A1(new_n5541_), .A2(\asqrt[55] ), .ZN(new_n5555_));
  AOI21_X1   g05363(.A1(new_n5555_), .A2(new_n5540_), .B(new_n724_), .ZN(new_n5556_));
  OAI21_X1   g05364(.A1(new_n5543_), .A2(new_n5556_), .B(\asqrt[57] ), .ZN(new_n5557_));
  AOI21_X1   g05365(.A1(new_n5547_), .A2(new_n5557_), .B(new_n504_), .ZN(new_n5558_));
  OAI21_X1   g05366(.A1(new_n5550_), .A2(new_n5558_), .B(\asqrt[59] ), .ZN(new_n5559_));
  AOI21_X1   g05367(.A1(new_n5559_), .A2(new_n5474_), .B(new_n5554_), .ZN(new_n5560_));
  OAI22_X1   g05368(.A1(new_n5551_), .A2(new_n504_), .B1(new_n5549_), .B2(new_n5547_), .ZN(new_n5561_));
  AOI22_X1   g05369(.A1(new_n5561_), .A2(\asqrt[59] ), .B1(new_n5553_), .B2(new_n5550_), .ZN(new_n5562_));
  NOR4_X1    g05370(.A1(new_n5273_), .A2(\asqrt[60] ), .A3(new_n5136_), .A4(new_n5242_), .ZN(new_n5563_));
  XOR2_X1    g05371(.A1(new_n5563_), .A2(new_n5293_), .Z(new_n5564_));
  NAND2_X1   g05372(.A1(new_n5564_), .A2(new_n229_), .ZN(new_n5565_));
  INV_X1     g05373(.I(new_n5565_), .ZN(new_n5566_));
  OAI21_X1   g05374(.A1(new_n5562_), .A2(new_n275_), .B(new_n5566_), .ZN(new_n5567_));
  NAND2_X1   g05375(.A1(new_n5567_), .A2(new_n5560_), .ZN(new_n5568_));
  INV_X1     g05376(.I(new_n5490_), .ZN(new_n5569_));
  NOR2_X1    g05377(.A1(new_n5569_), .A2(\asqrt[62] ), .ZN(new_n5570_));
  INV_X1     g05378(.I(new_n5570_), .ZN(new_n5571_));
  NAND2_X1   g05379(.A1(new_n5482_), .A2(new_n5571_), .ZN(new_n5572_));
  OAI21_X1   g05380(.A1(new_n5572_), .A2(new_n5568_), .B(new_n5492_), .ZN(new_n5573_));
  NOR3_X1    g05381(.A1(\asqrt[36] ), .A2(new_n4941_), .A3(new_n5246_), .ZN(new_n5574_));
  OAI21_X1   g05382(.A1(new_n5574_), .A2(new_n5258_), .B(new_n231_), .ZN(new_n5575_));
  OAI21_X1   g05383(.A1(new_n5573_), .A2(new_n5575_), .B(new_n5488_), .ZN(new_n5576_));
  OAI21_X1   g05384(.A1(new_n4941_), .A2(new_n5152_), .B(\asqrt[36] ), .ZN(new_n5577_));
  XOR2_X1    g05385(.A1(new_n5152_), .A2(\asqrt[63] ), .Z(new_n5578_));
  NAND2_X1   g05386(.A1(new_n5577_), .A2(new_n5578_), .ZN(new_n5579_));
  INV_X1     g05387(.I(new_n5579_), .ZN(new_n5580_));
  INV_X1     g05388(.I(new_n5488_), .ZN(new_n5581_));
  OAI22_X1   g05389(.A1(new_n5471_), .A2(new_n376_), .B1(new_n5469_), .B2(new_n5464_), .ZN(new_n5582_));
  AOI21_X1   g05390(.A1(new_n5582_), .A2(\asqrt[60] ), .B(new_n5565_), .ZN(new_n5583_));
  AOI22_X1   g05391(.A1(new_n5582_), .A2(\asqrt[60] ), .B1(new_n5475_), .B2(new_n5470_), .ZN(new_n5584_));
  OAI22_X1   g05392(.A1(new_n5584_), .A2(new_n229_), .B1(new_n5583_), .B2(new_n5476_), .ZN(new_n5585_));
  NOR4_X1    g05393(.A1(new_n5585_), .A2(\asqrt[62] ), .A3(new_n5581_), .A4(new_n5490_), .ZN(new_n5586_));
  NAND2_X1   g05394(.A1(new_n5586_), .A2(new_n5580_), .ZN(new_n5587_));
  NAND3_X1   g05395(.A1(new_n5267_), .A2(new_n4928_), .A3(new_n4941_), .ZN(new_n5588_));
  NOR3_X1    g05396(.A1(new_n5587_), .A2(new_n5576_), .A3(new_n5588_), .ZN(\asqrt[35] ));
  NAND2_X1   g05397(.A1(new_n5476_), .A2(new_n5481_), .ZN(new_n5590_));
  NOR3_X1    g05398(.A1(new_n5590_), .A2(\asqrt[61] ), .A3(new_n5564_), .ZN(new_n5591_));
  NAND2_X1   g05399(.A1(\asqrt[35] ), .A2(new_n5591_), .ZN(new_n5592_));
  XOR2_X1    g05400(.A1(new_n5592_), .A2(new_n5482_), .Z(new_n5593_));
  INV_X1     g05401(.I(new_n5593_), .ZN(new_n5594_));
  INV_X1     g05402(.I(\a[70] ), .ZN(new_n5595_));
  NOR2_X1    g05403(.A1(\a[68] ), .A2(\a[69] ), .ZN(new_n5596_));
  INV_X1     g05404(.I(new_n5596_), .ZN(new_n5597_));
  NOR3_X1    g05405(.A1(new_n5282_), .A2(new_n5595_), .A3(new_n5597_), .ZN(new_n5598_));
  NAND2_X1   g05406(.A1(new_n5297_), .A2(new_n5598_), .ZN(new_n5599_));
  XOR2_X1    g05407(.A1(new_n5599_), .A2(\a[71] ), .Z(new_n5600_));
  INV_X1     g05408(.I(\a[71] ), .ZN(new_n5601_));
  NOR4_X1    g05409(.A1(new_n5587_), .A2(new_n5576_), .A3(new_n5601_), .A4(new_n5588_), .ZN(new_n5602_));
  NOR2_X1    g05410(.A1(new_n5601_), .A2(\a[70] ), .ZN(new_n5603_));
  OAI21_X1   g05411(.A1(new_n5602_), .A2(new_n5603_), .B(new_n5600_), .ZN(new_n5604_));
  INV_X1     g05412(.I(new_n5600_), .ZN(new_n5605_));
  NOR2_X1    g05413(.A1(new_n5583_), .A2(new_n5476_), .ZN(new_n5606_));
  NOR3_X1    g05414(.A1(new_n5584_), .A2(new_n229_), .A3(new_n5570_), .ZN(new_n5607_));
  AOI21_X1   g05415(.A1(new_n5607_), .A2(new_n5606_), .B(new_n5491_), .ZN(new_n5608_));
  INV_X1     g05416(.I(new_n5575_), .ZN(new_n5609_));
  AOI21_X1   g05417(.A1(new_n5608_), .A2(new_n5609_), .B(new_n5581_), .ZN(new_n5610_));
  AOI21_X1   g05418(.A1(new_n5585_), .A2(\asqrt[62] ), .B(new_n5488_), .ZN(new_n5611_));
  AOI21_X1   g05419(.A1(new_n5554_), .A2(new_n5559_), .B(new_n275_), .ZN(new_n5612_));
  OAI21_X1   g05420(.A1(new_n5560_), .A2(new_n5612_), .B(\asqrt[61] ), .ZN(new_n5613_));
  NAND4_X1   g05421(.A1(new_n5568_), .A2(new_n5613_), .A3(new_n196_), .A4(new_n5569_), .ZN(new_n5614_));
  NOR3_X1    g05422(.A1(new_n5611_), .A2(new_n5579_), .A3(new_n5614_), .ZN(new_n5615_));
  INV_X1     g05423(.I(new_n5588_), .ZN(new_n5616_));
  NAND4_X1   g05424(.A1(new_n5615_), .A2(\a[71] ), .A3(new_n5610_), .A4(new_n5616_), .ZN(new_n5617_));
  NAND3_X1   g05425(.A1(new_n5617_), .A2(\a[70] ), .A3(new_n5605_), .ZN(new_n5618_));
  NAND2_X1   g05426(.A1(new_n5604_), .A2(new_n5618_), .ZN(new_n5619_));
  NOR2_X1    g05427(.A1(new_n5587_), .A2(new_n5576_), .ZN(new_n5620_));
  NAND4_X1   g05428(.A1(new_n5263_), .A2(new_n5255_), .A3(new_n4941_), .A4(new_n5296_), .ZN(new_n5621_));
  NOR2_X1    g05429(.A1(new_n5273_), .A2(new_n5595_), .ZN(new_n5622_));
  XOR2_X1    g05430(.A1(new_n5622_), .A2(new_n5621_), .Z(new_n5623_));
  NOR2_X1    g05431(.A1(new_n5623_), .A2(new_n5597_), .ZN(new_n5624_));
  INV_X1     g05432(.I(new_n5624_), .ZN(new_n5625_));
  NAND3_X1   g05433(.A1(new_n5615_), .A2(new_n5610_), .A3(new_n5616_), .ZN(new_n5626_));
  NOR4_X1    g05434(.A1(new_n5613_), .A2(new_n5476_), .A3(new_n5583_), .A4(new_n5570_), .ZN(new_n5627_));
  NOR3_X1    g05435(.A1(new_n5627_), .A2(new_n5491_), .A3(new_n5575_), .ZN(new_n5628_));
  AOI22_X1   g05436(.A1(new_n5590_), .A2(\asqrt[61] ), .B1(new_n5567_), .B2(new_n5560_), .ZN(new_n5629_));
  NAND4_X1   g05437(.A1(new_n5629_), .A2(new_n196_), .A3(new_n5488_), .A4(new_n5569_), .ZN(new_n5630_));
  OAI21_X1   g05438(.A1(new_n5628_), .A2(new_n5581_), .B(new_n5630_), .ZN(new_n5631_));
  NOR2_X1    g05439(.A1(new_n5580_), .A2(new_n5616_), .ZN(new_n5632_));
  NAND2_X1   g05440(.A1(new_n5632_), .A2(\asqrt[36] ), .ZN(new_n5633_));
  OAI21_X1   g05441(.A1(new_n5631_), .A2(new_n5633_), .B(new_n4908_), .ZN(new_n5634_));
  NAND3_X1   g05442(.A1(new_n5634_), .A2(new_n4916_), .A3(new_n5626_), .ZN(new_n5635_));
  NAND4_X1   g05443(.A1(new_n5482_), .A2(new_n5560_), .A3(new_n5567_), .A4(new_n5571_), .ZN(new_n5636_));
  NAND3_X1   g05444(.A1(new_n5636_), .A2(new_n5492_), .A3(new_n5609_), .ZN(new_n5637_));
  AOI21_X1   g05445(.A1(new_n5488_), .A2(new_n5637_), .B(new_n5586_), .ZN(new_n5638_));
  INV_X1     g05446(.I(new_n5633_), .ZN(new_n5639_));
  AOI21_X1   g05447(.A1(new_n5638_), .A2(new_n5639_), .B(\a[72] ), .ZN(new_n5640_));
  OAI21_X1   g05448(.A1(new_n5640_), .A2(new_n4917_), .B(\asqrt[35] ), .ZN(new_n5641_));
  NAND4_X1   g05449(.A1(new_n5635_), .A2(new_n5641_), .A3(new_n4973_), .A4(new_n5625_), .ZN(new_n5642_));
  NAND2_X1   g05450(.A1(new_n5642_), .A2(new_n5619_), .ZN(new_n5643_));
  NAND3_X1   g05451(.A1(new_n5604_), .A2(new_n5618_), .A3(new_n5625_), .ZN(new_n5644_));
  AOI21_X1   g05452(.A1(\asqrt[36] ), .A2(new_n4908_), .B(\a[73] ), .ZN(new_n5645_));
  NOR2_X1    g05453(.A1(new_n5264_), .A2(\a[72] ), .ZN(new_n5646_));
  AOI21_X1   g05454(.A1(\asqrt[36] ), .A2(\a[72] ), .B(new_n4919_), .ZN(new_n5647_));
  OAI21_X1   g05455(.A1(new_n5645_), .A2(new_n5646_), .B(new_n5647_), .ZN(new_n5648_));
  INV_X1     g05456(.I(new_n5648_), .ZN(new_n5649_));
  NAND3_X1   g05457(.A1(\asqrt[35] ), .A2(new_n5272_), .A3(new_n5649_), .ZN(new_n5650_));
  OAI21_X1   g05458(.A1(new_n5626_), .A2(new_n5648_), .B(new_n5271_), .ZN(new_n5651_));
  NAND3_X1   g05459(.A1(new_n5650_), .A2(new_n5651_), .A3(new_n4645_), .ZN(new_n5652_));
  AOI21_X1   g05460(.A1(new_n5644_), .A2(\asqrt[37] ), .B(new_n5652_), .ZN(new_n5653_));
  NOR2_X1    g05461(.A1(new_n5643_), .A2(new_n5653_), .ZN(new_n5654_));
  AOI22_X1   g05462(.A1(new_n5642_), .A2(new_n5619_), .B1(\asqrt[37] ), .B2(new_n5644_), .ZN(new_n5655_));
  INV_X1     g05463(.I(new_n5252_), .ZN(new_n5656_));
  AOI21_X1   g05464(.A1(new_n5264_), .A2(new_n5656_), .B(new_n5254_), .ZN(new_n5657_));
  INV_X1     g05465(.I(new_n5265_), .ZN(new_n5658_));
  NOR3_X1    g05466(.A1(new_n5658_), .A2(new_n5657_), .A3(new_n5271_), .ZN(new_n5659_));
  AOI21_X1   g05467(.A1(new_n5300_), .A2(new_n5285_), .B(\asqrt[38] ), .ZN(new_n5660_));
  AND4_X2    g05468(.A1(new_n5659_), .A2(\asqrt[35] ), .A3(new_n5314_), .A4(new_n5660_), .Z(new_n5661_));
  NOR2_X1    g05469(.A1(new_n5659_), .A2(new_n4645_), .ZN(new_n5662_));
  NOR3_X1    g05470(.A1(new_n5661_), .A2(\asqrt[39] ), .A3(new_n5662_), .ZN(new_n5663_));
  OAI21_X1   g05471(.A1(new_n5655_), .A2(new_n4645_), .B(new_n5663_), .ZN(new_n5664_));
  NAND2_X1   g05472(.A1(new_n5664_), .A2(new_n5654_), .ZN(new_n5665_));
  OAI22_X1   g05473(.A1(new_n5655_), .A2(new_n4645_), .B1(new_n5643_), .B2(new_n5653_), .ZN(new_n5666_));
  NAND2_X1   g05474(.A1(new_n5310_), .A2(new_n5309_), .ZN(new_n5667_));
  NAND4_X1   g05475(.A1(\asqrt[35] ), .A2(new_n4330_), .A3(new_n5667_), .A4(new_n5347_), .ZN(new_n5668_));
  XOR2_X1    g05476(.A1(new_n5668_), .A2(new_n5315_), .Z(new_n5669_));
  NAND2_X1   g05477(.A1(new_n5669_), .A2(new_n4018_), .ZN(new_n5670_));
  AOI21_X1   g05478(.A1(new_n5666_), .A2(\asqrt[39] ), .B(new_n5670_), .ZN(new_n5671_));
  NOR2_X1    g05479(.A1(new_n5671_), .A2(new_n5665_), .ZN(new_n5672_));
  AOI22_X1   g05480(.A1(new_n5666_), .A2(\asqrt[39] ), .B1(new_n5664_), .B2(new_n5654_), .ZN(new_n5673_));
  NOR2_X1    g05481(.A1(new_n5320_), .A2(new_n5321_), .ZN(new_n5674_));
  NOR4_X1    g05482(.A1(new_n5626_), .A2(\asqrt[40] ), .A3(new_n5674_), .A4(new_n5349_), .ZN(new_n5675_));
  XOR2_X1    g05483(.A1(new_n5675_), .A2(new_n5325_), .Z(new_n5676_));
  NAND2_X1   g05484(.A1(new_n5676_), .A2(new_n3760_), .ZN(new_n5677_));
  INV_X1     g05485(.I(new_n5677_), .ZN(new_n5678_));
  OAI21_X1   g05486(.A1(new_n5673_), .A2(new_n4018_), .B(new_n5678_), .ZN(new_n5679_));
  NAND2_X1   g05487(.A1(new_n5679_), .A2(new_n5672_), .ZN(new_n5680_));
  OAI22_X1   g05488(.A1(new_n5673_), .A2(new_n4018_), .B1(new_n5671_), .B2(new_n5665_), .ZN(new_n5681_));
  NOR2_X1    g05489(.A1(new_n5329_), .A2(\asqrt[41] ), .ZN(new_n5682_));
  NAND3_X1   g05490(.A1(\asqrt[35] ), .A2(new_n5350_), .A3(new_n5682_), .ZN(new_n5683_));
  XOR2_X1    g05491(.A1(new_n5683_), .A2(new_n5333_), .Z(new_n5684_));
  NAND2_X1   g05492(.A1(new_n5684_), .A2(new_n3481_), .ZN(new_n5685_));
  AOI21_X1   g05493(.A1(new_n5681_), .A2(\asqrt[41] ), .B(new_n5685_), .ZN(new_n5686_));
  NOR2_X1    g05494(.A1(new_n5686_), .A2(new_n5680_), .ZN(new_n5687_));
  AOI22_X1   g05495(.A1(new_n5681_), .A2(\asqrt[41] ), .B1(new_n5679_), .B2(new_n5672_), .ZN(new_n5688_));
  NOR4_X1    g05496(.A1(new_n5626_), .A2(\asqrt[42] ), .A3(new_n5337_), .A4(new_n5354_), .ZN(new_n5689_));
  XOR2_X1    g05497(.A1(new_n5689_), .A2(new_n5340_), .Z(new_n5690_));
  NAND2_X1   g05498(.A1(new_n5690_), .A2(new_n3208_), .ZN(new_n5691_));
  INV_X1     g05499(.I(new_n5691_), .ZN(new_n5692_));
  OAI21_X1   g05500(.A1(new_n5688_), .A2(new_n3481_), .B(new_n5692_), .ZN(new_n5693_));
  NAND2_X1   g05501(.A1(new_n5693_), .A2(new_n5687_), .ZN(new_n5694_));
  OAI22_X1   g05502(.A1(new_n5688_), .A2(new_n3481_), .B1(new_n5686_), .B2(new_n5680_), .ZN(new_n5695_));
  NOR4_X1    g05503(.A1(new_n5626_), .A2(\asqrt[43] ), .A3(new_n5343_), .A4(new_n5497_), .ZN(new_n5696_));
  XNOR2_X1   g05504(.A1(new_n5696_), .A2(new_n5500_), .ZN(new_n5697_));
  NAND2_X1   g05505(.A1(new_n5697_), .A2(new_n2941_), .ZN(new_n5698_));
  AOI21_X1   g05506(.A1(new_n5695_), .A2(\asqrt[43] ), .B(new_n5698_), .ZN(new_n5699_));
  NOR2_X1    g05507(.A1(new_n5699_), .A2(new_n5694_), .ZN(new_n5700_));
  AOI22_X1   g05508(.A1(new_n5695_), .A2(\asqrt[43] ), .B1(new_n5693_), .B2(new_n5687_), .ZN(new_n5701_));
  NOR4_X1    g05509(.A1(new_n5626_), .A2(\asqrt[44] ), .A3(new_n5358_), .A4(new_n5364_), .ZN(new_n5702_));
  XOR2_X1    g05510(.A1(new_n5702_), .A2(new_n5501_), .Z(new_n5703_));
  NAND2_X1   g05511(.A1(new_n5703_), .A2(new_n2728_), .ZN(new_n5704_));
  INV_X1     g05512(.I(new_n5704_), .ZN(new_n5705_));
  OAI21_X1   g05513(.A1(new_n5701_), .A2(new_n2941_), .B(new_n5705_), .ZN(new_n5706_));
  NAND2_X1   g05514(.A1(new_n5706_), .A2(new_n5700_), .ZN(new_n5707_));
  OAI22_X1   g05515(.A1(new_n5701_), .A2(new_n2941_), .B1(new_n5699_), .B2(new_n5694_), .ZN(new_n5708_));
  NAND2_X1   g05516(.A1(new_n5506_), .A2(\asqrt[45] ), .ZN(new_n5709_));
  NOR4_X1    g05517(.A1(new_n5626_), .A2(\asqrt[45] ), .A3(new_n5367_), .A4(new_n5506_), .ZN(new_n5710_));
  XOR2_X1    g05518(.A1(new_n5710_), .A2(new_n5709_), .Z(new_n5711_));
  NAND2_X1   g05519(.A1(new_n5711_), .A2(new_n2488_), .ZN(new_n5712_));
  AOI21_X1   g05520(.A1(new_n5708_), .A2(\asqrt[45] ), .B(new_n5712_), .ZN(new_n5713_));
  NOR2_X1    g05521(.A1(new_n5713_), .A2(new_n5707_), .ZN(new_n5714_));
  AOI22_X1   g05522(.A1(new_n5708_), .A2(\asqrt[45] ), .B1(new_n5706_), .B2(new_n5700_), .ZN(new_n5715_));
  NOR4_X1    g05523(.A1(new_n5626_), .A2(\asqrt[46] ), .A3(new_n5374_), .A4(new_n5379_), .ZN(new_n5716_));
  AOI21_X1   g05524(.A1(new_n5709_), .A2(new_n5504_), .B(new_n2488_), .ZN(new_n5717_));
  NOR2_X1    g05525(.A1(new_n5716_), .A2(new_n5717_), .ZN(new_n5718_));
  NAND2_X1   g05526(.A1(new_n5718_), .A2(new_n2253_), .ZN(new_n5719_));
  INV_X1     g05527(.I(new_n5719_), .ZN(new_n5720_));
  OAI21_X1   g05528(.A1(new_n5715_), .A2(new_n2488_), .B(new_n5720_), .ZN(new_n5721_));
  NAND2_X1   g05529(.A1(new_n5721_), .A2(new_n5714_), .ZN(new_n5722_));
  OAI22_X1   g05530(.A1(new_n5715_), .A2(new_n2488_), .B1(new_n5713_), .B2(new_n5707_), .ZN(new_n5723_));
  NAND2_X1   g05531(.A1(new_n5513_), .A2(\asqrt[47] ), .ZN(new_n5724_));
  NOR4_X1    g05532(.A1(new_n5626_), .A2(\asqrt[47] ), .A3(new_n5382_), .A4(new_n5513_), .ZN(new_n5725_));
  XOR2_X1    g05533(.A1(new_n5725_), .A2(new_n5724_), .Z(new_n5726_));
  NAND2_X1   g05534(.A1(new_n5726_), .A2(new_n2046_), .ZN(new_n5727_));
  AOI21_X1   g05535(.A1(new_n5723_), .A2(\asqrt[47] ), .B(new_n5727_), .ZN(new_n5728_));
  NOR2_X1    g05536(.A1(new_n5728_), .A2(new_n5722_), .ZN(new_n5729_));
  AOI22_X1   g05537(.A1(new_n5723_), .A2(\asqrt[47] ), .B1(new_n5721_), .B2(new_n5714_), .ZN(new_n5730_));
  NOR4_X1    g05538(.A1(new_n5626_), .A2(\asqrt[48] ), .A3(new_n5389_), .A4(new_n5394_), .ZN(new_n5731_));
  AOI21_X1   g05539(.A1(new_n5724_), .A2(new_n5512_), .B(new_n2046_), .ZN(new_n5732_));
  NOR2_X1    g05540(.A1(new_n5731_), .A2(new_n5732_), .ZN(new_n5733_));
  NAND2_X1   g05541(.A1(new_n5733_), .A2(new_n1854_), .ZN(new_n5734_));
  INV_X1     g05542(.I(new_n5734_), .ZN(new_n5735_));
  OAI21_X1   g05543(.A1(new_n5730_), .A2(new_n2046_), .B(new_n5735_), .ZN(new_n5736_));
  NAND2_X1   g05544(.A1(new_n5736_), .A2(new_n5729_), .ZN(new_n5737_));
  OAI22_X1   g05545(.A1(new_n5730_), .A2(new_n2046_), .B1(new_n5728_), .B2(new_n5722_), .ZN(new_n5738_));
  NAND2_X1   g05546(.A1(new_n5520_), .A2(\asqrt[49] ), .ZN(new_n5739_));
  NOR4_X1    g05547(.A1(new_n5626_), .A2(\asqrt[49] ), .A3(new_n5397_), .A4(new_n5520_), .ZN(new_n5740_));
  XOR2_X1    g05548(.A1(new_n5740_), .A2(new_n5739_), .Z(new_n5741_));
  NAND2_X1   g05549(.A1(new_n5741_), .A2(new_n1595_), .ZN(new_n5742_));
  AOI21_X1   g05550(.A1(new_n5738_), .A2(\asqrt[49] ), .B(new_n5742_), .ZN(new_n5743_));
  NOR2_X1    g05551(.A1(new_n5743_), .A2(new_n5737_), .ZN(new_n5744_));
  AOI22_X1   g05552(.A1(new_n5738_), .A2(\asqrt[49] ), .B1(new_n5736_), .B2(new_n5729_), .ZN(new_n5745_));
  NOR4_X1    g05553(.A1(new_n5626_), .A2(\asqrt[50] ), .A3(new_n5404_), .A4(new_n5409_), .ZN(new_n5746_));
  AOI21_X1   g05554(.A1(new_n5739_), .A2(new_n5519_), .B(new_n1595_), .ZN(new_n5747_));
  NOR2_X1    g05555(.A1(new_n5746_), .A2(new_n5747_), .ZN(new_n5748_));
  NAND2_X1   g05556(.A1(new_n5748_), .A2(new_n1436_), .ZN(new_n5749_));
  INV_X1     g05557(.I(new_n5749_), .ZN(new_n5750_));
  OAI21_X1   g05558(.A1(new_n5745_), .A2(new_n1595_), .B(new_n5750_), .ZN(new_n5751_));
  NAND2_X1   g05559(.A1(new_n5751_), .A2(new_n5744_), .ZN(new_n5752_));
  OAI22_X1   g05560(.A1(new_n5745_), .A2(new_n1595_), .B1(new_n5743_), .B2(new_n5737_), .ZN(new_n5753_));
  NAND2_X1   g05561(.A1(new_n5527_), .A2(\asqrt[51] ), .ZN(new_n5754_));
  NOR4_X1    g05562(.A1(new_n5626_), .A2(\asqrt[51] ), .A3(new_n5412_), .A4(new_n5527_), .ZN(new_n5755_));
  XOR2_X1    g05563(.A1(new_n5755_), .A2(new_n5754_), .Z(new_n5756_));
  NAND2_X1   g05564(.A1(new_n5756_), .A2(new_n1260_), .ZN(new_n5757_));
  AOI21_X1   g05565(.A1(new_n5753_), .A2(\asqrt[51] ), .B(new_n5757_), .ZN(new_n5758_));
  NOR2_X1    g05566(.A1(new_n5758_), .A2(new_n5752_), .ZN(new_n5759_));
  AOI22_X1   g05567(.A1(new_n5753_), .A2(\asqrt[51] ), .B1(new_n5751_), .B2(new_n5744_), .ZN(new_n5760_));
  NOR4_X1    g05568(.A1(new_n5626_), .A2(\asqrt[52] ), .A3(new_n5419_), .A4(new_n5424_), .ZN(new_n5761_));
  AOI21_X1   g05569(.A1(new_n5754_), .A2(new_n5526_), .B(new_n1260_), .ZN(new_n5762_));
  NOR2_X1    g05570(.A1(new_n5761_), .A2(new_n5762_), .ZN(new_n5763_));
  NAND2_X1   g05571(.A1(new_n5763_), .A2(new_n1096_), .ZN(new_n5764_));
  INV_X1     g05572(.I(new_n5764_), .ZN(new_n5765_));
  OAI21_X1   g05573(.A1(new_n5760_), .A2(new_n1260_), .B(new_n5765_), .ZN(new_n5766_));
  NAND2_X1   g05574(.A1(new_n5766_), .A2(new_n5759_), .ZN(new_n5767_));
  OAI22_X1   g05575(.A1(new_n5760_), .A2(new_n1260_), .B1(new_n5758_), .B2(new_n5752_), .ZN(new_n5768_));
  NAND2_X1   g05576(.A1(new_n5534_), .A2(\asqrt[53] ), .ZN(new_n5769_));
  NOR4_X1    g05577(.A1(new_n5626_), .A2(\asqrt[53] ), .A3(new_n5427_), .A4(new_n5534_), .ZN(new_n5770_));
  XOR2_X1    g05578(.A1(new_n5770_), .A2(new_n5769_), .Z(new_n5771_));
  NAND2_X1   g05579(.A1(new_n5771_), .A2(new_n970_), .ZN(new_n5772_));
  AOI21_X1   g05580(.A1(new_n5768_), .A2(\asqrt[53] ), .B(new_n5772_), .ZN(new_n5773_));
  NOR2_X1    g05581(.A1(new_n5773_), .A2(new_n5767_), .ZN(new_n5774_));
  AOI22_X1   g05582(.A1(new_n5768_), .A2(\asqrt[53] ), .B1(new_n5766_), .B2(new_n5759_), .ZN(new_n5775_));
  NOR4_X1    g05583(.A1(new_n5626_), .A2(\asqrt[54] ), .A3(new_n5434_), .A4(new_n5439_), .ZN(new_n5776_));
  AOI21_X1   g05584(.A1(new_n5769_), .A2(new_n5533_), .B(new_n970_), .ZN(new_n5777_));
  NOR2_X1    g05585(.A1(new_n5776_), .A2(new_n5777_), .ZN(new_n5778_));
  NAND2_X1   g05586(.A1(new_n5778_), .A2(new_n825_), .ZN(new_n5779_));
  INV_X1     g05587(.I(new_n5779_), .ZN(new_n5780_));
  OAI21_X1   g05588(.A1(new_n5775_), .A2(new_n970_), .B(new_n5780_), .ZN(new_n5781_));
  NAND2_X1   g05589(.A1(new_n5781_), .A2(new_n5774_), .ZN(new_n5782_));
  OAI22_X1   g05590(.A1(new_n5775_), .A2(new_n970_), .B1(new_n5773_), .B2(new_n5767_), .ZN(new_n5783_));
  NOR4_X1    g05591(.A1(new_n5626_), .A2(\asqrt[55] ), .A3(new_n5441_), .A4(new_n5541_), .ZN(new_n5784_));
  XOR2_X1    g05592(.A1(new_n5784_), .A2(new_n5555_), .Z(new_n5785_));
  NAND2_X1   g05593(.A1(new_n5785_), .A2(new_n724_), .ZN(new_n5786_));
  AOI21_X1   g05594(.A1(new_n5783_), .A2(\asqrt[55] ), .B(new_n5786_), .ZN(new_n5787_));
  NOR2_X1    g05595(.A1(new_n5787_), .A2(new_n5782_), .ZN(new_n5788_));
  AOI22_X1   g05596(.A1(new_n5783_), .A2(\asqrt[55] ), .B1(new_n5781_), .B2(new_n5774_), .ZN(new_n5789_));
  NOR4_X1    g05597(.A1(new_n5626_), .A2(\asqrt[56] ), .A3(new_n5447_), .A4(new_n5452_), .ZN(new_n5790_));
  XOR2_X1    g05598(.A1(new_n5790_), .A2(new_n5477_), .Z(new_n5791_));
  NAND2_X1   g05599(.A1(new_n5791_), .A2(new_n587_), .ZN(new_n5792_));
  INV_X1     g05600(.I(new_n5792_), .ZN(new_n5793_));
  OAI21_X1   g05601(.A1(new_n5789_), .A2(new_n724_), .B(new_n5793_), .ZN(new_n5794_));
  NAND2_X1   g05602(.A1(new_n5794_), .A2(new_n5788_), .ZN(new_n5795_));
  OAI22_X1   g05603(.A1(new_n5789_), .A2(new_n724_), .B1(new_n5787_), .B2(new_n5782_), .ZN(new_n5796_));
  NOR4_X1    g05604(.A1(new_n5626_), .A2(\asqrt[57] ), .A3(new_n5454_), .A4(new_n5548_), .ZN(new_n5797_));
  XOR2_X1    g05605(.A1(new_n5797_), .A2(new_n5557_), .Z(new_n5798_));
  NAND2_X1   g05606(.A1(new_n5798_), .A2(new_n504_), .ZN(new_n5799_));
  AOI21_X1   g05607(.A1(new_n5796_), .A2(\asqrt[57] ), .B(new_n5799_), .ZN(new_n5800_));
  NOR2_X1    g05608(.A1(new_n5800_), .A2(new_n5795_), .ZN(new_n5801_));
  AOI22_X1   g05609(.A1(new_n5796_), .A2(\asqrt[57] ), .B1(new_n5794_), .B2(new_n5788_), .ZN(new_n5802_));
  NOR4_X1    g05610(.A1(new_n5626_), .A2(\asqrt[58] ), .A3(new_n5460_), .A4(new_n5465_), .ZN(new_n5803_));
  XOR2_X1    g05611(.A1(new_n5803_), .A2(new_n5479_), .Z(new_n5804_));
  NAND2_X1   g05612(.A1(new_n5804_), .A2(new_n376_), .ZN(new_n5805_));
  INV_X1     g05613(.I(new_n5805_), .ZN(new_n5806_));
  OAI21_X1   g05614(.A1(new_n5802_), .A2(new_n504_), .B(new_n5806_), .ZN(new_n5807_));
  NAND2_X1   g05615(.A1(new_n5807_), .A2(new_n5801_), .ZN(new_n5808_));
  OAI22_X1   g05616(.A1(new_n5802_), .A2(new_n504_), .B1(new_n5800_), .B2(new_n5795_), .ZN(new_n5809_));
  NOR4_X1    g05617(.A1(new_n5626_), .A2(\asqrt[59] ), .A3(new_n5467_), .A4(new_n5561_), .ZN(new_n5810_));
  XOR2_X1    g05618(.A1(new_n5810_), .A2(new_n5559_), .Z(new_n5811_));
  NAND2_X1   g05619(.A1(new_n5811_), .A2(new_n275_), .ZN(new_n5812_));
  AOI21_X1   g05620(.A1(new_n5809_), .A2(\asqrt[59] ), .B(new_n5812_), .ZN(new_n5813_));
  NOR2_X1    g05621(.A1(new_n5813_), .A2(new_n5808_), .ZN(new_n5814_));
  AOI22_X1   g05622(.A1(new_n5809_), .A2(\asqrt[59] ), .B1(new_n5807_), .B2(new_n5801_), .ZN(new_n5815_));
  OAI22_X1   g05623(.A1(new_n5815_), .A2(new_n275_), .B1(new_n5813_), .B2(new_n5808_), .ZN(new_n5816_));
  NOR4_X1    g05624(.A1(new_n5626_), .A2(\asqrt[60] ), .A3(new_n5473_), .A4(new_n5582_), .ZN(new_n5817_));
  XOR2_X1    g05625(.A1(new_n5817_), .A2(new_n5481_), .Z(new_n5818_));
  NAND2_X1   g05626(.A1(new_n5818_), .A2(new_n229_), .ZN(new_n5819_));
  INV_X1     g05627(.I(new_n5819_), .ZN(new_n5820_));
  OAI21_X1   g05628(.A1(new_n5815_), .A2(new_n275_), .B(new_n5820_), .ZN(new_n5821_));
  AOI22_X1   g05629(.A1(new_n5816_), .A2(\asqrt[61] ), .B1(new_n5821_), .B2(new_n5814_), .ZN(new_n5822_));
  NOR2_X1    g05630(.A1(new_n5822_), .A2(new_n196_), .ZN(new_n5823_));
  INV_X1     g05631(.I(new_n5603_), .ZN(new_n5824_));
  AOI21_X1   g05632(.A1(new_n5617_), .A2(new_n5824_), .B(new_n5605_), .ZN(new_n5825_));
  NOR3_X1    g05633(.A1(new_n5602_), .A2(new_n5595_), .A3(new_n5600_), .ZN(new_n5826_));
  NOR2_X1    g05634(.A1(new_n5826_), .A2(new_n5825_), .ZN(new_n5827_));
  NOR3_X1    g05635(.A1(new_n5640_), .A2(new_n4917_), .A3(\asqrt[35] ), .ZN(new_n5828_));
  AOI21_X1   g05636(.A1(new_n5634_), .A2(new_n4916_), .B(new_n5626_), .ZN(new_n5829_));
  NOR4_X1    g05637(.A1(new_n5829_), .A2(new_n5828_), .A3(\asqrt[37] ), .A4(new_n5624_), .ZN(new_n5830_));
  NOR2_X1    g05638(.A1(new_n5830_), .A2(new_n5827_), .ZN(new_n5831_));
  NOR3_X1    g05639(.A1(new_n5826_), .A2(new_n5825_), .A3(new_n5624_), .ZN(new_n5832_));
  NOR3_X1    g05640(.A1(new_n5626_), .A2(new_n5271_), .A3(new_n5648_), .ZN(new_n5833_));
  AOI21_X1   g05641(.A1(\asqrt[35] ), .A2(new_n5649_), .B(new_n5272_), .ZN(new_n5834_));
  NOR3_X1    g05642(.A1(new_n5834_), .A2(new_n5833_), .A3(\asqrt[38] ), .ZN(new_n5835_));
  OAI21_X1   g05643(.A1(new_n5832_), .A2(new_n4973_), .B(new_n5835_), .ZN(new_n5836_));
  NAND2_X1   g05644(.A1(new_n5831_), .A2(new_n5836_), .ZN(new_n5837_));
  OAI22_X1   g05645(.A1(new_n5830_), .A2(new_n5827_), .B1(new_n4973_), .B2(new_n5832_), .ZN(new_n5838_));
  INV_X1     g05646(.I(new_n5663_), .ZN(new_n5839_));
  AOI21_X1   g05647(.A1(new_n5838_), .A2(\asqrt[38] ), .B(new_n5839_), .ZN(new_n5840_));
  NOR2_X1    g05648(.A1(new_n5840_), .A2(new_n5837_), .ZN(new_n5841_));
  AOI22_X1   g05649(.A1(new_n5838_), .A2(\asqrt[38] ), .B1(new_n5831_), .B2(new_n5836_), .ZN(new_n5842_));
  INV_X1     g05650(.I(new_n5670_), .ZN(new_n5843_));
  OAI21_X1   g05651(.A1(new_n5842_), .A2(new_n4330_), .B(new_n5843_), .ZN(new_n5844_));
  NAND2_X1   g05652(.A1(new_n5844_), .A2(new_n5841_), .ZN(new_n5845_));
  OAI22_X1   g05653(.A1(new_n5842_), .A2(new_n4330_), .B1(new_n5840_), .B2(new_n5837_), .ZN(new_n5846_));
  AOI21_X1   g05654(.A1(new_n5846_), .A2(\asqrt[40] ), .B(new_n5677_), .ZN(new_n5847_));
  NOR2_X1    g05655(.A1(new_n5847_), .A2(new_n5845_), .ZN(new_n5848_));
  AOI22_X1   g05656(.A1(new_n5846_), .A2(\asqrt[40] ), .B1(new_n5844_), .B2(new_n5841_), .ZN(new_n5849_));
  INV_X1     g05657(.I(new_n5685_), .ZN(new_n5850_));
  OAI21_X1   g05658(.A1(new_n5849_), .A2(new_n3760_), .B(new_n5850_), .ZN(new_n5851_));
  NAND2_X1   g05659(.A1(new_n5851_), .A2(new_n5848_), .ZN(new_n5852_));
  OAI22_X1   g05660(.A1(new_n5849_), .A2(new_n3760_), .B1(new_n5847_), .B2(new_n5845_), .ZN(new_n5853_));
  AOI21_X1   g05661(.A1(new_n5853_), .A2(\asqrt[42] ), .B(new_n5691_), .ZN(new_n5854_));
  NOR2_X1    g05662(.A1(new_n5854_), .A2(new_n5852_), .ZN(new_n5855_));
  AOI22_X1   g05663(.A1(new_n5853_), .A2(\asqrt[42] ), .B1(new_n5851_), .B2(new_n5848_), .ZN(new_n5856_));
  INV_X1     g05664(.I(new_n5698_), .ZN(new_n5857_));
  OAI21_X1   g05665(.A1(new_n5856_), .A2(new_n3208_), .B(new_n5857_), .ZN(new_n5858_));
  NAND2_X1   g05666(.A1(new_n5858_), .A2(new_n5855_), .ZN(new_n5859_));
  OAI22_X1   g05667(.A1(new_n5856_), .A2(new_n3208_), .B1(new_n5854_), .B2(new_n5852_), .ZN(new_n5860_));
  AOI21_X1   g05668(.A1(new_n5860_), .A2(\asqrt[44] ), .B(new_n5704_), .ZN(new_n5861_));
  NOR2_X1    g05669(.A1(new_n5861_), .A2(new_n5859_), .ZN(new_n5862_));
  AOI22_X1   g05670(.A1(new_n5860_), .A2(\asqrt[44] ), .B1(new_n5858_), .B2(new_n5855_), .ZN(new_n5863_));
  INV_X1     g05671(.I(new_n5712_), .ZN(new_n5864_));
  OAI21_X1   g05672(.A1(new_n5863_), .A2(new_n2728_), .B(new_n5864_), .ZN(new_n5865_));
  NAND2_X1   g05673(.A1(new_n5865_), .A2(new_n5862_), .ZN(new_n5866_));
  OAI22_X1   g05674(.A1(new_n5863_), .A2(new_n2728_), .B1(new_n5861_), .B2(new_n5859_), .ZN(new_n5867_));
  AOI21_X1   g05675(.A1(new_n5867_), .A2(\asqrt[46] ), .B(new_n5719_), .ZN(new_n5868_));
  NOR2_X1    g05676(.A1(new_n5868_), .A2(new_n5866_), .ZN(new_n5869_));
  AOI22_X1   g05677(.A1(new_n5867_), .A2(\asqrt[46] ), .B1(new_n5865_), .B2(new_n5862_), .ZN(new_n5870_));
  INV_X1     g05678(.I(new_n5727_), .ZN(new_n5871_));
  OAI21_X1   g05679(.A1(new_n5870_), .A2(new_n2253_), .B(new_n5871_), .ZN(new_n5872_));
  NAND2_X1   g05680(.A1(new_n5872_), .A2(new_n5869_), .ZN(new_n5873_));
  OAI22_X1   g05681(.A1(new_n5870_), .A2(new_n2253_), .B1(new_n5868_), .B2(new_n5866_), .ZN(new_n5874_));
  AOI21_X1   g05682(.A1(new_n5874_), .A2(\asqrt[48] ), .B(new_n5734_), .ZN(new_n5875_));
  NOR2_X1    g05683(.A1(new_n5875_), .A2(new_n5873_), .ZN(new_n5876_));
  AOI22_X1   g05684(.A1(new_n5874_), .A2(\asqrt[48] ), .B1(new_n5872_), .B2(new_n5869_), .ZN(new_n5877_));
  INV_X1     g05685(.I(new_n5742_), .ZN(new_n5878_));
  OAI21_X1   g05686(.A1(new_n5877_), .A2(new_n1854_), .B(new_n5878_), .ZN(new_n5879_));
  NAND2_X1   g05687(.A1(new_n5879_), .A2(new_n5876_), .ZN(new_n5880_));
  OAI22_X1   g05688(.A1(new_n5877_), .A2(new_n1854_), .B1(new_n5875_), .B2(new_n5873_), .ZN(new_n5881_));
  AOI21_X1   g05689(.A1(new_n5881_), .A2(\asqrt[50] ), .B(new_n5749_), .ZN(new_n5882_));
  NOR2_X1    g05690(.A1(new_n5882_), .A2(new_n5880_), .ZN(new_n5883_));
  AOI22_X1   g05691(.A1(new_n5881_), .A2(\asqrt[50] ), .B1(new_n5879_), .B2(new_n5876_), .ZN(new_n5884_));
  INV_X1     g05692(.I(new_n5757_), .ZN(new_n5885_));
  OAI21_X1   g05693(.A1(new_n5884_), .A2(new_n1436_), .B(new_n5885_), .ZN(new_n5886_));
  NAND2_X1   g05694(.A1(new_n5886_), .A2(new_n5883_), .ZN(new_n5887_));
  OAI22_X1   g05695(.A1(new_n5884_), .A2(new_n1436_), .B1(new_n5882_), .B2(new_n5880_), .ZN(new_n5888_));
  AOI21_X1   g05696(.A1(new_n5888_), .A2(\asqrt[52] ), .B(new_n5764_), .ZN(new_n5889_));
  NOR2_X1    g05697(.A1(new_n5889_), .A2(new_n5887_), .ZN(new_n5890_));
  AOI22_X1   g05698(.A1(new_n5888_), .A2(\asqrt[52] ), .B1(new_n5886_), .B2(new_n5883_), .ZN(new_n5891_));
  INV_X1     g05699(.I(new_n5772_), .ZN(new_n5892_));
  OAI21_X1   g05700(.A1(new_n5891_), .A2(new_n1096_), .B(new_n5892_), .ZN(new_n5893_));
  NAND2_X1   g05701(.A1(new_n5893_), .A2(new_n5890_), .ZN(new_n5894_));
  OAI22_X1   g05702(.A1(new_n5891_), .A2(new_n1096_), .B1(new_n5889_), .B2(new_n5887_), .ZN(new_n5895_));
  AOI21_X1   g05703(.A1(new_n5895_), .A2(\asqrt[54] ), .B(new_n5779_), .ZN(new_n5896_));
  NOR2_X1    g05704(.A1(new_n5896_), .A2(new_n5894_), .ZN(new_n5897_));
  AOI22_X1   g05705(.A1(new_n5895_), .A2(\asqrt[54] ), .B1(new_n5893_), .B2(new_n5890_), .ZN(new_n5898_));
  INV_X1     g05706(.I(new_n5786_), .ZN(new_n5899_));
  OAI21_X1   g05707(.A1(new_n5898_), .A2(new_n825_), .B(new_n5899_), .ZN(new_n5900_));
  NAND2_X1   g05708(.A1(new_n5900_), .A2(new_n5897_), .ZN(new_n5901_));
  OAI22_X1   g05709(.A1(new_n5898_), .A2(new_n825_), .B1(new_n5896_), .B2(new_n5894_), .ZN(new_n5902_));
  AOI21_X1   g05710(.A1(new_n5902_), .A2(\asqrt[56] ), .B(new_n5792_), .ZN(new_n5903_));
  NOR2_X1    g05711(.A1(new_n5903_), .A2(new_n5901_), .ZN(new_n5904_));
  AOI22_X1   g05712(.A1(new_n5902_), .A2(\asqrt[56] ), .B1(new_n5900_), .B2(new_n5897_), .ZN(new_n5905_));
  INV_X1     g05713(.I(new_n5799_), .ZN(new_n5906_));
  OAI21_X1   g05714(.A1(new_n5905_), .A2(new_n587_), .B(new_n5906_), .ZN(new_n5907_));
  NAND2_X1   g05715(.A1(new_n5907_), .A2(new_n5904_), .ZN(new_n5908_));
  OAI22_X1   g05716(.A1(new_n5905_), .A2(new_n587_), .B1(new_n5903_), .B2(new_n5901_), .ZN(new_n5909_));
  AOI21_X1   g05717(.A1(new_n5909_), .A2(\asqrt[58] ), .B(new_n5805_), .ZN(new_n5910_));
  NOR2_X1    g05718(.A1(new_n5910_), .A2(new_n5908_), .ZN(new_n5911_));
  AOI22_X1   g05719(.A1(new_n5909_), .A2(\asqrt[58] ), .B1(new_n5907_), .B2(new_n5904_), .ZN(new_n5912_));
  INV_X1     g05720(.I(new_n5812_), .ZN(new_n5913_));
  OAI21_X1   g05721(.A1(new_n5912_), .A2(new_n376_), .B(new_n5913_), .ZN(new_n5914_));
  NAND2_X1   g05722(.A1(new_n5914_), .A2(new_n5911_), .ZN(new_n5915_));
  OAI22_X1   g05723(.A1(new_n5912_), .A2(new_n376_), .B1(new_n5910_), .B2(new_n5908_), .ZN(new_n5916_));
  AOI22_X1   g05724(.A1(new_n5916_), .A2(\asqrt[60] ), .B1(new_n5914_), .B2(new_n5911_), .ZN(new_n5917_));
  AOI21_X1   g05725(.A1(new_n5916_), .A2(\asqrt[60] ), .B(new_n5819_), .ZN(new_n5918_));
  OAI22_X1   g05726(.A1(new_n5917_), .A2(new_n229_), .B1(new_n5918_), .B2(new_n5915_), .ZN(new_n5919_));
  NOR2_X1    g05727(.A1(new_n5919_), .A2(\asqrt[62] ), .ZN(new_n5920_));
  NAND3_X1   g05728(.A1(new_n5620_), .A2(new_n5488_), .A3(new_n5588_), .ZN(new_n5921_));
  NOR2_X1    g05729(.A1(new_n5629_), .A2(new_n196_), .ZN(new_n5922_));
  INV_X1     g05730(.I(new_n5614_), .ZN(new_n5923_));
  NAND3_X1   g05731(.A1(\asqrt[35] ), .A2(new_n5922_), .A3(new_n5923_), .ZN(new_n5924_));
  OAI21_X1   g05732(.A1(new_n5585_), .A2(\asqrt[62] ), .B(new_n5490_), .ZN(new_n5925_));
  OAI21_X1   g05733(.A1(\asqrt[35] ), .A2(new_n5925_), .B(new_n5922_), .ZN(new_n5926_));
  NAND2_X1   g05734(.A1(new_n5926_), .A2(new_n5924_), .ZN(new_n5927_));
  INV_X1     g05735(.I(new_n5927_), .ZN(new_n5928_));
  NOR2_X1    g05736(.A1(new_n5593_), .A2(new_n196_), .ZN(new_n5929_));
  INV_X1     g05737(.I(new_n5929_), .ZN(new_n5930_));
  NAND2_X1   g05738(.A1(new_n5796_), .A2(\asqrt[57] ), .ZN(new_n5931_));
  AOI21_X1   g05739(.A1(new_n5931_), .A2(new_n5795_), .B(new_n504_), .ZN(new_n5932_));
  OAI21_X1   g05740(.A1(new_n5801_), .A2(new_n5932_), .B(\asqrt[59] ), .ZN(new_n5933_));
  AOI21_X1   g05741(.A1(new_n5808_), .A2(new_n5933_), .B(new_n275_), .ZN(new_n5934_));
  OAI21_X1   g05742(.A1(new_n5814_), .A2(new_n5934_), .B(\asqrt[61] ), .ZN(new_n5935_));
  NOR2_X1    g05743(.A1(new_n5594_), .A2(\asqrt[62] ), .ZN(new_n5936_));
  INV_X1     g05744(.I(new_n5936_), .ZN(new_n5937_));
  NAND3_X1   g05745(.A1(new_n5821_), .A2(new_n5814_), .A3(new_n5937_), .ZN(new_n5938_));
  OAI21_X1   g05746(.A1(new_n5938_), .A2(new_n5935_), .B(new_n5930_), .ZN(new_n5939_));
  NAND3_X1   g05747(.A1(new_n5626_), .A2(new_n5581_), .A3(new_n5630_), .ZN(new_n5940_));
  AOI21_X1   g05748(.A1(new_n5940_), .A2(new_n5573_), .B(\asqrt[63] ), .ZN(new_n5941_));
  INV_X1     g05749(.I(new_n5941_), .ZN(new_n5942_));
  OAI21_X1   g05750(.A1(new_n5939_), .A2(new_n5942_), .B(new_n5928_), .ZN(new_n5943_));
  NOR4_X1    g05751(.A1(new_n5919_), .A2(\asqrt[62] ), .A3(new_n5927_), .A4(new_n5593_), .ZN(new_n5944_));
  NAND2_X1   g05752(.A1(new_n5608_), .A2(new_n5581_), .ZN(new_n5945_));
  XOR2_X1    g05753(.A1(new_n5608_), .A2(\asqrt[63] ), .Z(new_n5946_));
  AOI21_X1   g05754(.A1(\asqrt[35] ), .A2(new_n5945_), .B(new_n5946_), .ZN(new_n5947_));
  NAND2_X1   g05755(.A1(new_n5944_), .A2(new_n5947_), .ZN(new_n5948_));
  NOR3_X1    g05756(.A1(new_n5948_), .A2(new_n5921_), .A3(new_n5943_), .ZN(\asqrt[34] ));
  NAND4_X1   g05757(.A1(\asqrt[34] ), .A2(new_n5594_), .A3(new_n5823_), .A4(new_n5920_), .ZN(new_n5950_));
  OAI21_X1   g05758(.A1(new_n5919_), .A2(\asqrt[62] ), .B(new_n5593_), .ZN(new_n5951_));
  OAI21_X1   g05759(.A1(\asqrt[34] ), .A2(new_n5951_), .B(new_n5823_), .ZN(new_n5952_));
  NAND2_X1   g05760(.A1(new_n5950_), .A2(new_n5952_), .ZN(new_n5953_));
  INV_X1     g05761(.I(new_n5953_), .ZN(new_n5954_));
  NAND2_X1   g05762(.A1(new_n5909_), .A2(\asqrt[58] ), .ZN(new_n5955_));
  AOI21_X1   g05763(.A1(new_n5955_), .A2(new_n5908_), .B(new_n376_), .ZN(new_n5956_));
  OAI21_X1   g05764(.A1(new_n5911_), .A2(new_n5956_), .B(\asqrt[60] ), .ZN(new_n5957_));
  AOI21_X1   g05765(.A1(new_n5915_), .A2(new_n5957_), .B(new_n229_), .ZN(new_n5958_));
  NOR3_X1    g05766(.A1(new_n5816_), .A2(\asqrt[61] ), .A3(new_n5818_), .ZN(new_n5959_));
  NAND2_X1   g05767(.A1(\asqrt[34] ), .A2(new_n5959_), .ZN(new_n5960_));
  XOR2_X1    g05768(.A1(new_n5960_), .A2(new_n5958_), .Z(new_n5961_));
  NOR2_X1    g05769(.A1(new_n5961_), .A2(new_n196_), .ZN(new_n5962_));
  INV_X1     g05770(.I(new_n5962_), .ZN(new_n5963_));
  INV_X1     g05771(.I(\a[68] ), .ZN(new_n5964_));
  NOR2_X1    g05772(.A1(\a[66] ), .A2(\a[67] ), .ZN(new_n5965_));
  INV_X1     g05773(.I(new_n5965_), .ZN(new_n5966_));
  NOR3_X1    g05774(.A1(new_n5632_), .A2(new_n5964_), .A3(new_n5966_), .ZN(new_n5967_));
  NAND2_X1   g05775(.A1(new_n5638_), .A2(new_n5967_), .ZN(new_n5968_));
  XOR2_X1    g05776(.A1(new_n5968_), .A2(\a[69] ), .Z(new_n5969_));
  INV_X1     g05777(.I(\a[69] ), .ZN(new_n5970_));
  NOR4_X1    g05778(.A1(new_n5948_), .A2(new_n5970_), .A3(new_n5921_), .A4(new_n5943_), .ZN(new_n5971_));
  NOR2_X1    g05779(.A1(new_n5970_), .A2(\a[68] ), .ZN(new_n5972_));
  OAI21_X1   g05780(.A1(new_n5971_), .A2(new_n5972_), .B(new_n5969_), .ZN(new_n5973_));
  INV_X1     g05781(.I(new_n5969_), .ZN(new_n5974_));
  INV_X1     g05782(.I(new_n5921_), .ZN(new_n5975_));
  NOR3_X1    g05783(.A1(new_n5918_), .A2(new_n5915_), .A3(new_n5936_), .ZN(new_n5976_));
  AOI21_X1   g05784(.A1(new_n5976_), .A2(new_n5958_), .B(new_n5929_), .ZN(new_n5977_));
  AOI21_X1   g05785(.A1(new_n5977_), .A2(new_n5941_), .B(new_n5927_), .ZN(new_n5978_));
  NAND4_X1   g05786(.A1(new_n5822_), .A2(new_n196_), .A3(new_n5928_), .A4(new_n5594_), .ZN(new_n5979_));
  INV_X1     g05787(.I(new_n5947_), .ZN(new_n5980_));
  NOR2_X1    g05788(.A1(new_n5979_), .A2(new_n5980_), .ZN(new_n5981_));
  NAND4_X1   g05789(.A1(new_n5981_), .A2(\a[69] ), .A3(new_n5978_), .A4(new_n5975_), .ZN(new_n5982_));
  NAND3_X1   g05790(.A1(new_n5982_), .A2(\a[68] ), .A3(new_n5974_), .ZN(new_n5983_));
  NAND2_X1   g05791(.A1(new_n5973_), .A2(new_n5983_), .ZN(new_n5984_));
  NOR2_X1    g05792(.A1(new_n5948_), .A2(new_n5943_), .ZN(new_n5985_));
  NOR4_X1    g05793(.A1(new_n5587_), .A2(new_n5581_), .A3(new_n5628_), .A4(new_n5588_), .ZN(new_n5986_));
  NAND2_X1   g05794(.A1(\asqrt[35] ), .A2(\a[68] ), .ZN(new_n5987_));
  XOR2_X1    g05795(.A1(new_n5987_), .A2(new_n5986_), .Z(new_n5988_));
  NOR2_X1    g05796(.A1(new_n5988_), .A2(new_n5966_), .ZN(new_n5989_));
  INV_X1     g05797(.I(new_n5989_), .ZN(new_n5990_));
  NAND3_X1   g05798(.A1(new_n5981_), .A2(new_n5975_), .A3(new_n5978_), .ZN(new_n5991_));
  NOR2_X1    g05799(.A1(new_n5975_), .A2(new_n5947_), .ZN(new_n5992_));
  NAND2_X1   g05800(.A1(new_n5992_), .A2(\asqrt[35] ), .ZN(new_n5993_));
  INV_X1     g05801(.I(new_n5993_), .ZN(new_n5994_));
  NAND3_X1   g05802(.A1(new_n5943_), .A2(new_n5979_), .A3(new_n5994_), .ZN(new_n5995_));
  NAND2_X1   g05803(.A1(new_n5995_), .A2(new_n5595_), .ZN(new_n5996_));
  NAND3_X1   g05804(.A1(new_n5996_), .A2(new_n5596_), .A3(new_n5991_), .ZN(new_n5997_));
  NOR3_X1    g05805(.A1(new_n5978_), .A2(new_n5944_), .A3(new_n5993_), .ZN(new_n5998_));
  OAI21_X1   g05806(.A1(new_n5998_), .A2(\a[70] ), .B(new_n5596_), .ZN(new_n5999_));
  NAND2_X1   g05807(.A1(new_n5999_), .A2(\asqrt[34] ), .ZN(new_n6000_));
  NAND4_X1   g05808(.A1(new_n6000_), .A2(new_n5273_), .A3(new_n5997_), .A4(new_n5990_), .ZN(new_n6001_));
  NAND2_X1   g05809(.A1(new_n6001_), .A2(new_n5984_), .ZN(new_n6002_));
  NAND3_X1   g05810(.A1(new_n5973_), .A2(new_n5983_), .A3(new_n5990_), .ZN(new_n6003_));
  AOI21_X1   g05811(.A1(\asqrt[35] ), .A2(new_n5595_), .B(\a[71] ), .ZN(new_n6004_));
  NOR2_X1    g05812(.A1(new_n5617_), .A2(\a[70] ), .ZN(new_n6005_));
  AOI21_X1   g05813(.A1(\asqrt[35] ), .A2(\a[70] ), .B(new_n5599_), .ZN(new_n6006_));
  OAI21_X1   g05814(.A1(new_n6005_), .A2(new_n6004_), .B(new_n6006_), .ZN(new_n6007_));
  INV_X1     g05815(.I(new_n6007_), .ZN(new_n6008_));
  NAND3_X1   g05816(.A1(\asqrt[34] ), .A2(new_n5625_), .A3(new_n6008_), .ZN(new_n6009_));
  OAI21_X1   g05817(.A1(new_n5991_), .A2(new_n6007_), .B(new_n5624_), .ZN(new_n6010_));
  NAND3_X1   g05818(.A1(new_n6009_), .A2(new_n6010_), .A3(new_n4973_), .ZN(new_n6011_));
  AOI21_X1   g05819(.A1(new_n6003_), .A2(\asqrt[36] ), .B(new_n6011_), .ZN(new_n6012_));
  NOR2_X1    g05820(.A1(new_n6002_), .A2(new_n6012_), .ZN(new_n6013_));
  NAND2_X1   g05821(.A1(new_n6003_), .A2(\asqrt[36] ), .ZN(new_n6014_));
  AOI21_X1   g05822(.A1(new_n6002_), .A2(new_n6014_), .B(new_n4973_), .ZN(new_n6015_));
  NOR2_X1    g05823(.A1(new_n5829_), .A2(new_n5828_), .ZN(new_n6016_));
  NOR4_X1    g05824(.A1(new_n5991_), .A2(\asqrt[37] ), .A3(new_n6016_), .A4(new_n5644_), .ZN(new_n6017_));
  AOI21_X1   g05825(.A1(new_n5827_), .A2(new_n5625_), .B(new_n4973_), .ZN(new_n6018_));
  NOR2_X1    g05826(.A1(new_n6017_), .A2(new_n6018_), .ZN(new_n6019_));
  NAND2_X1   g05827(.A1(new_n6019_), .A2(new_n4645_), .ZN(new_n6020_));
  OAI21_X1   g05828(.A1(new_n6015_), .A2(new_n6020_), .B(new_n6013_), .ZN(new_n6021_));
  AOI22_X1   g05829(.A1(new_n6001_), .A2(new_n5984_), .B1(\asqrt[36] ), .B2(new_n6003_), .ZN(new_n6022_));
  OAI22_X1   g05830(.A1(new_n6022_), .A2(new_n4973_), .B1(new_n6002_), .B2(new_n6012_), .ZN(new_n6023_));
  NOR2_X1    g05831(.A1(new_n5655_), .A2(new_n4645_), .ZN(new_n6024_));
  NAND2_X1   g05832(.A1(new_n5650_), .A2(new_n5651_), .ZN(new_n6025_));
  NAND4_X1   g05833(.A1(\asqrt[34] ), .A2(new_n4645_), .A3(new_n6025_), .A4(new_n5655_), .ZN(new_n6026_));
  XOR2_X1    g05834(.A1(new_n6026_), .A2(new_n6024_), .Z(new_n6027_));
  NAND2_X1   g05835(.A1(new_n6027_), .A2(new_n4330_), .ZN(new_n6028_));
  AOI21_X1   g05836(.A1(new_n6023_), .A2(\asqrt[38] ), .B(new_n6028_), .ZN(new_n6029_));
  OAI21_X1   g05837(.A1(new_n6015_), .A2(new_n6013_), .B(\asqrt[38] ), .ZN(new_n6030_));
  AOI21_X1   g05838(.A1(new_n6021_), .A2(new_n6030_), .B(new_n4330_), .ZN(new_n6031_));
  NAND2_X1   g05839(.A1(new_n5666_), .A2(\asqrt[39] ), .ZN(new_n6032_));
  OAI21_X1   g05840(.A1(new_n5661_), .A2(new_n5662_), .B(new_n4330_), .ZN(new_n6033_));
  NOR2_X1    g05841(.A1(new_n5666_), .A2(new_n6033_), .ZN(new_n6034_));
  NAND2_X1   g05842(.A1(\asqrt[34] ), .A2(new_n6034_), .ZN(new_n6035_));
  XNOR2_X1   g05843(.A1(new_n6035_), .A2(new_n6032_), .ZN(new_n6036_));
  NAND2_X1   g05844(.A1(new_n6036_), .A2(new_n4018_), .ZN(new_n6037_));
  NOR2_X1    g05845(.A1(new_n6031_), .A2(new_n6037_), .ZN(new_n6038_));
  NOR3_X1    g05846(.A1(new_n6038_), .A2(new_n6021_), .A3(new_n6029_), .ZN(new_n6039_));
  INV_X1     g05847(.I(new_n6028_), .ZN(new_n6040_));
  AOI21_X1   g05848(.A1(new_n6030_), .A2(new_n6040_), .B(new_n6021_), .ZN(new_n6041_));
  OAI21_X1   g05849(.A1(new_n6041_), .A2(new_n6031_), .B(\asqrt[40] ), .ZN(new_n6042_));
  NAND2_X1   g05850(.A1(new_n5846_), .A2(\asqrt[40] ), .ZN(new_n6043_));
  NOR4_X1    g05851(.A1(new_n5991_), .A2(\asqrt[40] ), .A3(new_n5669_), .A4(new_n5846_), .ZN(new_n6044_));
  XOR2_X1    g05852(.A1(new_n6044_), .A2(new_n6043_), .Z(new_n6045_));
  NAND2_X1   g05853(.A1(new_n6045_), .A2(new_n3760_), .ZN(new_n6046_));
  INV_X1     g05854(.I(new_n6046_), .ZN(new_n6047_));
  NAND2_X1   g05855(.A1(new_n6042_), .A2(new_n6047_), .ZN(new_n6048_));
  NAND2_X1   g05856(.A1(new_n6048_), .A2(new_n6039_), .ZN(new_n6049_));
  OAI21_X1   g05857(.A1(new_n6031_), .A2(new_n6037_), .B(new_n6041_), .ZN(new_n6050_));
  NAND2_X1   g05858(.A1(new_n6050_), .A2(new_n6042_), .ZN(new_n6051_));
  NAND2_X1   g05859(.A1(new_n5681_), .A2(\asqrt[41] ), .ZN(new_n6052_));
  NOR4_X1    g05860(.A1(new_n5991_), .A2(\asqrt[41] ), .A3(new_n5676_), .A4(new_n5681_), .ZN(new_n6053_));
  XOR2_X1    g05861(.A1(new_n6053_), .A2(new_n6052_), .Z(new_n6054_));
  NAND2_X1   g05862(.A1(new_n6054_), .A2(new_n3481_), .ZN(new_n6055_));
  AOI21_X1   g05863(.A1(new_n6051_), .A2(\asqrt[41] ), .B(new_n6055_), .ZN(new_n6056_));
  NOR2_X1    g05864(.A1(new_n6056_), .A2(new_n6049_), .ZN(new_n6057_));
  AOI21_X1   g05865(.A1(new_n6042_), .A2(new_n6047_), .B(new_n6050_), .ZN(new_n6058_));
  AOI21_X1   g05866(.A1(new_n6050_), .A2(new_n6042_), .B(new_n3760_), .ZN(new_n6059_));
  OAI21_X1   g05867(.A1(new_n6058_), .A2(new_n6059_), .B(\asqrt[42] ), .ZN(new_n6060_));
  NAND2_X1   g05868(.A1(new_n5853_), .A2(\asqrt[42] ), .ZN(new_n6061_));
  NOR4_X1    g05869(.A1(new_n5991_), .A2(\asqrt[42] ), .A3(new_n5684_), .A4(new_n5853_), .ZN(new_n6062_));
  XOR2_X1    g05870(.A1(new_n6062_), .A2(new_n6061_), .Z(new_n6063_));
  NAND2_X1   g05871(.A1(new_n6063_), .A2(new_n3208_), .ZN(new_n6064_));
  INV_X1     g05872(.I(new_n6064_), .ZN(new_n6065_));
  NAND2_X1   g05873(.A1(new_n6060_), .A2(new_n6065_), .ZN(new_n6066_));
  NAND2_X1   g05874(.A1(new_n6066_), .A2(new_n6057_), .ZN(new_n6067_));
  AOI22_X1   g05875(.A1(new_n6051_), .A2(\asqrt[41] ), .B1(new_n6048_), .B2(new_n6039_), .ZN(new_n6068_));
  OAI22_X1   g05876(.A1(new_n6068_), .A2(new_n3481_), .B1(new_n6056_), .B2(new_n6049_), .ZN(new_n6069_));
  NAND2_X1   g05877(.A1(new_n5695_), .A2(\asqrt[43] ), .ZN(new_n6070_));
  NOR4_X1    g05878(.A1(new_n5991_), .A2(\asqrt[43] ), .A3(new_n5690_), .A4(new_n5695_), .ZN(new_n6071_));
  XOR2_X1    g05879(.A1(new_n6071_), .A2(new_n6070_), .Z(new_n6072_));
  NAND2_X1   g05880(.A1(new_n6072_), .A2(new_n2941_), .ZN(new_n6073_));
  AOI21_X1   g05881(.A1(new_n6069_), .A2(\asqrt[43] ), .B(new_n6073_), .ZN(new_n6074_));
  NOR2_X1    g05882(.A1(new_n6074_), .A2(new_n6067_), .ZN(new_n6075_));
  AOI22_X1   g05883(.A1(new_n6069_), .A2(\asqrt[43] ), .B1(new_n6066_), .B2(new_n6057_), .ZN(new_n6076_));
  NAND2_X1   g05884(.A1(new_n5860_), .A2(\asqrt[44] ), .ZN(new_n6077_));
  NOR4_X1    g05885(.A1(new_n5991_), .A2(\asqrt[44] ), .A3(new_n5697_), .A4(new_n5860_), .ZN(new_n6078_));
  XOR2_X1    g05886(.A1(new_n6078_), .A2(new_n6077_), .Z(new_n6079_));
  NAND2_X1   g05887(.A1(new_n6079_), .A2(new_n2728_), .ZN(new_n6080_));
  INV_X1     g05888(.I(new_n6080_), .ZN(new_n6081_));
  OAI21_X1   g05889(.A1(new_n6076_), .A2(new_n2941_), .B(new_n6081_), .ZN(new_n6082_));
  NAND2_X1   g05890(.A1(new_n6082_), .A2(new_n6075_), .ZN(new_n6083_));
  OAI22_X1   g05891(.A1(new_n6076_), .A2(new_n2941_), .B1(new_n6074_), .B2(new_n6067_), .ZN(new_n6084_));
  NAND2_X1   g05892(.A1(new_n5708_), .A2(\asqrt[45] ), .ZN(new_n6085_));
  NOR4_X1    g05893(.A1(new_n5991_), .A2(\asqrt[45] ), .A3(new_n5703_), .A4(new_n5708_), .ZN(new_n6086_));
  XOR2_X1    g05894(.A1(new_n6086_), .A2(new_n6085_), .Z(new_n6087_));
  NAND2_X1   g05895(.A1(new_n6087_), .A2(new_n2488_), .ZN(new_n6088_));
  AOI21_X1   g05896(.A1(new_n6084_), .A2(\asqrt[45] ), .B(new_n6088_), .ZN(new_n6089_));
  NOR2_X1    g05897(.A1(new_n6089_), .A2(new_n6083_), .ZN(new_n6090_));
  AOI22_X1   g05898(.A1(new_n6084_), .A2(\asqrt[45] ), .B1(new_n6082_), .B2(new_n6075_), .ZN(new_n6091_));
  NAND2_X1   g05899(.A1(new_n5867_), .A2(\asqrt[46] ), .ZN(new_n6092_));
  NOR4_X1    g05900(.A1(new_n5991_), .A2(\asqrt[46] ), .A3(new_n5711_), .A4(new_n5867_), .ZN(new_n6093_));
  XOR2_X1    g05901(.A1(new_n6093_), .A2(new_n6092_), .Z(new_n6094_));
  NAND2_X1   g05902(.A1(new_n6094_), .A2(new_n2253_), .ZN(new_n6095_));
  INV_X1     g05903(.I(new_n6095_), .ZN(new_n6096_));
  OAI21_X1   g05904(.A1(new_n6091_), .A2(new_n2488_), .B(new_n6096_), .ZN(new_n6097_));
  NAND2_X1   g05905(.A1(new_n6097_), .A2(new_n6090_), .ZN(new_n6098_));
  OAI22_X1   g05906(.A1(new_n6091_), .A2(new_n2488_), .B1(new_n6089_), .B2(new_n6083_), .ZN(new_n6099_));
  NAND2_X1   g05907(.A1(new_n5723_), .A2(\asqrt[47] ), .ZN(new_n6100_));
  NOR4_X1    g05908(.A1(new_n5991_), .A2(\asqrt[47] ), .A3(new_n5718_), .A4(new_n5723_), .ZN(new_n6101_));
  XOR2_X1    g05909(.A1(new_n6101_), .A2(new_n6100_), .Z(new_n6102_));
  NAND2_X1   g05910(.A1(new_n6102_), .A2(new_n2046_), .ZN(new_n6103_));
  AOI21_X1   g05911(.A1(new_n6099_), .A2(\asqrt[47] ), .B(new_n6103_), .ZN(new_n6104_));
  NOR2_X1    g05912(.A1(new_n6104_), .A2(new_n6098_), .ZN(new_n6105_));
  AOI22_X1   g05913(.A1(new_n6099_), .A2(\asqrt[47] ), .B1(new_n6097_), .B2(new_n6090_), .ZN(new_n6106_));
  NAND2_X1   g05914(.A1(new_n5874_), .A2(\asqrt[48] ), .ZN(new_n6107_));
  NOR4_X1    g05915(.A1(new_n5991_), .A2(\asqrt[48] ), .A3(new_n5726_), .A4(new_n5874_), .ZN(new_n6108_));
  XOR2_X1    g05916(.A1(new_n6108_), .A2(new_n6107_), .Z(new_n6109_));
  NAND2_X1   g05917(.A1(new_n6109_), .A2(new_n1854_), .ZN(new_n6110_));
  INV_X1     g05918(.I(new_n6110_), .ZN(new_n6111_));
  OAI21_X1   g05919(.A1(new_n6106_), .A2(new_n2046_), .B(new_n6111_), .ZN(new_n6112_));
  NAND2_X1   g05920(.A1(new_n6112_), .A2(new_n6105_), .ZN(new_n6113_));
  OAI22_X1   g05921(.A1(new_n6106_), .A2(new_n2046_), .B1(new_n6104_), .B2(new_n6098_), .ZN(new_n6114_));
  NAND2_X1   g05922(.A1(new_n5738_), .A2(\asqrt[49] ), .ZN(new_n6115_));
  NOR4_X1    g05923(.A1(new_n5991_), .A2(\asqrt[49] ), .A3(new_n5733_), .A4(new_n5738_), .ZN(new_n6116_));
  XOR2_X1    g05924(.A1(new_n6116_), .A2(new_n6115_), .Z(new_n6117_));
  NAND2_X1   g05925(.A1(new_n6117_), .A2(new_n1595_), .ZN(new_n6118_));
  AOI21_X1   g05926(.A1(new_n6114_), .A2(\asqrt[49] ), .B(new_n6118_), .ZN(new_n6119_));
  NOR2_X1    g05927(.A1(new_n6119_), .A2(new_n6113_), .ZN(new_n6120_));
  AOI22_X1   g05928(.A1(new_n6114_), .A2(\asqrt[49] ), .B1(new_n6112_), .B2(new_n6105_), .ZN(new_n6121_));
  NAND2_X1   g05929(.A1(new_n5881_), .A2(\asqrt[50] ), .ZN(new_n6122_));
  NOR4_X1    g05930(.A1(new_n5991_), .A2(\asqrt[50] ), .A3(new_n5741_), .A4(new_n5881_), .ZN(new_n6123_));
  XOR2_X1    g05931(.A1(new_n6123_), .A2(new_n6122_), .Z(new_n6124_));
  NAND2_X1   g05932(.A1(new_n6124_), .A2(new_n1436_), .ZN(new_n6125_));
  INV_X1     g05933(.I(new_n6125_), .ZN(new_n6126_));
  OAI21_X1   g05934(.A1(new_n6121_), .A2(new_n1595_), .B(new_n6126_), .ZN(new_n6127_));
  NAND2_X1   g05935(.A1(new_n6127_), .A2(new_n6120_), .ZN(new_n6128_));
  OAI22_X1   g05936(.A1(new_n6121_), .A2(new_n1595_), .B1(new_n6119_), .B2(new_n6113_), .ZN(new_n6129_));
  NAND2_X1   g05937(.A1(new_n5753_), .A2(\asqrt[51] ), .ZN(new_n6130_));
  NOR4_X1    g05938(.A1(new_n5991_), .A2(\asqrt[51] ), .A3(new_n5748_), .A4(new_n5753_), .ZN(new_n6131_));
  XOR2_X1    g05939(.A1(new_n6131_), .A2(new_n6130_), .Z(new_n6132_));
  NAND2_X1   g05940(.A1(new_n6132_), .A2(new_n1260_), .ZN(new_n6133_));
  AOI21_X1   g05941(.A1(new_n6129_), .A2(\asqrt[51] ), .B(new_n6133_), .ZN(new_n6134_));
  NOR2_X1    g05942(.A1(new_n6134_), .A2(new_n6128_), .ZN(new_n6135_));
  AOI22_X1   g05943(.A1(new_n6129_), .A2(\asqrt[51] ), .B1(new_n6127_), .B2(new_n6120_), .ZN(new_n6136_));
  NAND2_X1   g05944(.A1(new_n5888_), .A2(\asqrt[52] ), .ZN(new_n6137_));
  NOR4_X1    g05945(.A1(new_n5991_), .A2(\asqrt[52] ), .A3(new_n5756_), .A4(new_n5888_), .ZN(new_n6138_));
  XOR2_X1    g05946(.A1(new_n6138_), .A2(new_n6137_), .Z(new_n6139_));
  NAND2_X1   g05947(.A1(new_n6139_), .A2(new_n1096_), .ZN(new_n6140_));
  INV_X1     g05948(.I(new_n6140_), .ZN(new_n6141_));
  OAI21_X1   g05949(.A1(new_n6136_), .A2(new_n1260_), .B(new_n6141_), .ZN(new_n6142_));
  NAND2_X1   g05950(.A1(new_n6142_), .A2(new_n6135_), .ZN(new_n6143_));
  OAI22_X1   g05951(.A1(new_n6136_), .A2(new_n1260_), .B1(new_n6134_), .B2(new_n6128_), .ZN(new_n6144_));
  NAND2_X1   g05952(.A1(new_n5768_), .A2(\asqrt[53] ), .ZN(new_n6145_));
  NOR4_X1    g05953(.A1(new_n5991_), .A2(\asqrt[53] ), .A3(new_n5763_), .A4(new_n5768_), .ZN(new_n6146_));
  XOR2_X1    g05954(.A1(new_n6146_), .A2(new_n6145_), .Z(new_n6147_));
  NAND2_X1   g05955(.A1(new_n6147_), .A2(new_n970_), .ZN(new_n6148_));
  AOI21_X1   g05956(.A1(new_n6144_), .A2(\asqrt[53] ), .B(new_n6148_), .ZN(new_n6149_));
  NOR2_X1    g05957(.A1(new_n6149_), .A2(new_n6143_), .ZN(new_n6150_));
  AOI22_X1   g05958(.A1(new_n6144_), .A2(\asqrt[53] ), .B1(new_n6142_), .B2(new_n6135_), .ZN(new_n6151_));
  NAND2_X1   g05959(.A1(new_n5895_), .A2(\asqrt[54] ), .ZN(new_n6152_));
  NOR4_X1    g05960(.A1(new_n5991_), .A2(\asqrt[54] ), .A3(new_n5771_), .A4(new_n5895_), .ZN(new_n6153_));
  XOR2_X1    g05961(.A1(new_n6153_), .A2(new_n6152_), .Z(new_n6154_));
  NAND2_X1   g05962(.A1(new_n6154_), .A2(new_n825_), .ZN(new_n6155_));
  INV_X1     g05963(.I(new_n6155_), .ZN(new_n6156_));
  OAI21_X1   g05964(.A1(new_n6151_), .A2(new_n970_), .B(new_n6156_), .ZN(new_n6157_));
  NAND2_X1   g05965(.A1(new_n6157_), .A2(new_n6150_), .ZN(new_n6158_));
  OAI22_X1   g05966(.A1(new_n6151_), .A2(new_n970_), .B1(new_n6149_), .B2(new_n6143_), .ZN(new_n6159_));
  NAND2_X1   g05967(.A1(new_n5783_), .A2(\asqrt[55] ), .ZN(new_n6160_));
  NOR4_X1    g05968(.A1(new_n5991_), .A2(\asqrt[55] ), .A3(new_n5778_), .A4(new_n5783_), .ZN(new_n6161_));
  XOR2_X1    g05969(.A1(new_n6161_), .A2(new_n6160_), .Z(new_n6162_));
  NAND2_X1   g05970(.A1(new_n6162_), .A2(new_n724_), .ZN(new_n6163_));
  AOI21_X1   g05971(.A1(new_n6159_), .A2(\asqrt[55] ), .B(new_n6163_), .ZN(new_n6164_));
  NOR2_X1    g05972(.A1(new_n6164_), .A2(new_n6158_), .ZN(new_n6165_));
  AOI22_X1   g05973(.A1(new_n6159_), .A2(\asqrt[55] ), .B1(new_n6157_), .B2(new_n6150_), .ZN(new_n6166_));
  NAND2_X1   g05974(.A1(new_n5902_), .A2(\asqrt[56] ), .ZN(new_n6167_));
  NOR4_X1    g05975(.A1(new_n5991_), .A2(\asqrt[56] ), .A3(new_n5785_), .A4(new_n5902_), .ZN(new_n6168_));
  XOR2_X1    g05976(.A1(new_n6168_), .A2(new_n6167_), .Z(new_n6169_));
  NAND2_X1   g05977(.A1(new_n6169_), .A2(new_n587_), .ZN(new_n6170_));
  INV_X1     g05978(.I(new_n6170_), .ZN(new_n6171_));
  OAI21_X1   g05979(.A1(new_n6166_), .A2(new_n724_), .B(new_n6171_), .ZN(new_n6172_));
  NAND2_X1   g05980(.A1(new_n6172_), .A2(new_n6165_), .ZN(new_n6173_));
  NAND2_X1   g05981(.A1(new_n6144_), .A2(\asqrt[53] ), .ZN(new_n6174_));
  AOI21_X1   g05982(.A1(new_n6174_), .A2(new_n6143_), .B(new_n970_), .ZN(new_n6175_));
  OAI21_X1   g05983(.A1(new_n6150_), .A2(new_n6175_), .B(\asqrt[55] ), .ZN(new_n6176_));
  AOI21_X1   g05984(.A1(new_n6158_), .A2(new_n6176_), .B(new_n724_), .ZN(new_n6177_));
  OAI21_X1   g05985(.A1(new_n6165_), .A2(new_n6177_), .B(\asqrt[57] ), .ZN(new_n6178_));
  NOR4_X1    g05986(.A1(new_n5991_), .A2(\asqrt[57] ), .A3(new_n5791_), .A4(new_n5796_), .ZN(new_n6179_));
  XOR2_X1    g05987(.A1(new_n6179_), .A2(new_n5931_), .Z(new_n6180_));
  NAND2_X1   g05988(.A1(new_n6180_), .A2(new_n504_), .ZN(new_n6181_));
  INV_X1     g05989(.I(new_n6181_), .ZN(new_n6182_));
  AOI21_X1   g05990(.A1(new_n6178_), .A2(new_n6182_), .B(new_n6173_), .ZN(new_n6183_));
  OAI22_X1   g05991(.A1(new_n6166_), .A2(new_n724_), .B1(new_n6164_), .B2(new_n6158_), .ZN(new_n6184_));
  AOI22_X1   g05992(.A1(new_n6184_), .A2(\asqrt[57] ), .B1(new_n6172_), .B2(new_n6165_), .ZN(new_n6185_));
  NOR4_X1    g05993(.A1(new_n5991_), .A2(\asqrt[58] ), .A3(new_n5798_), .A4(new_n5909_), .ZN(new_n6186_));
  XOR2_X1    g05994(.A1(new_n6186_), .A2(new_n5955_), .Z(new_n6187_));
  NAND2_X1   g05995(.A1(new_n6187_), .A2(new_n376_), .ZN(new_n6188_));
  INV_X1     g05996(.I(new_n6188_), .ZN(new_n6189_));
  OAI21_X1   g05997(.A1(new_n6185_), .A2(new_n504_), .B(new_n6189_), .ZN(new_n6190_));
  NAND2_X1   g05998(.A1(new_n6190_), .A2(new_n6183_), .ZN(new_n6191_));
  AOI21_X1   g05999(.A1(new_n6173_), .A2(new_n6178_), .B(new_n504_), .ZN(new_n6192_));
  OAI21_X1   g06000(.A1(new_n6183_), .A2(new_n6192_), .B(\asqrt[59] ), .ZN(new_n6193_));
  NOR4_X1    g06001(.A1(new_n5991_), .A2(\asqrt[59] ), .A3(new_n5804_), .A4(new_n5809_), .ZN(new_n6194_));
  XOR2_X1    g06002(.A1(new_n6194_), .A2(new_n5933_), .Z(new_n6195_));
  AND2_X2    g06003(.A1(new_n6195_), .A2(new_n275_), .Z(new_n6196_));
  AOI21_X1   g06004(.A1(new_n6193_), .A2(new_n6196_), .B(new_n6191_), .ZN(new_n6197_));
  INV_X1     g06005(.I(new_n6020_), .ZN(new_n6198_));
  OAI21_X1   g06006(.A1(new_n6022_), .A2(new_n4973_), .B(new_n6198_), .ZN(new_n6199_));
  AOI22_X1   g06007(.A1(new_n6023_), .A2(\asqrt[38] ), .B1(new_n6199_), .B2(new_n6013_), .ZN(new_n6200_));
  INV_X1     g06008(.I(new_n6037_), .ZN(new_n6201_));
  OAI21_X1   g06009(.A1(new_n6200_), .A2(new_n4330_), .B(new_n6201_), .ZN(new_n6202_));
  OAI22_X1   g06010(.A1(new_n6200_), .A2(new_n4330_), .B1(new_n6029_), .B2(new_n6021_), .ZN(new_n6203_));
  AOI22_X1   g06011(.A1(new_n6203_), .A2(\asqrt[40] ), .B1(new_n6202_), .B2(new_n6041_), .ZN(new_n6204_));
  INV_X1     g06012(.I(new_n6055_), .ZN(new_n6205_));
  OAI21_X1   g06013(.A1(new_n6204_), .A2(new_n3760_), .B(new_n6205_), .ZN(new_n6206_));
  NAND2_X1   g06014(.A1(new_n6206_), .A2(new_n6058_), .ZN(new_n6207_));
  AOI21_X1   g06015(.A1(new_n6203_), .A2(\asqrt[40] ), .B(new_n6046_), .ZN(new_n6208_));
  OAI22_X1   g06016(.A1(new_n6204_), .A2(new_n3760_), .B1(new_n6208_), .B2(new_n6050_), .ZN(new_n6209_));
  AOI21_X1   g06017(.A1(new_n6209_), .A2(\asqrt[42] ), .B(new_n6064_), .ZN(new_n6210_));
  NOR2_X1    g06018(.A1(new_n6210_), .A2(new_n6207_), .ZN(new_n6211_));
  AOI22_X1   g06019(.A1(new_n6209_), .A2(\asqrt[42] ), .B1(new_n6206_), .B2(new_n6058_), .ZN(new_n6212_));
  INV_X1     g06020(.I(new_n6073_), .ZN(new_n6213_));
  OAI21_X1   g06021(.A1(new_n6212_), .A2(new_n3208_), .B(new_n6213_), .ZN(new_n6214_));
  NAND2_X1   g06022(.A1(new_n6214_), .A2(new_n6211_), .ZN(new_n6215_));
  OAI22_X1   g06023(.A1(new_n6212_), .A2(new_n3208_), .B1(new_n6210_), .B2(new_n6207_), .ZN(new_n6216_));
  AOI21_X1   g06024(.A1(new_n6216_), .A2(\asqrt[44] ), .B(new_n6080_), .ZN(new_n6217_));
  NOR2_X1    g06025(.A1(new_n6217_), .A2(new_n6215_), .ZN(new_n6218_));
  AOI22_X1   g06026(.A1(new_n6216_), .A2(\asqrt[44] ), .B1(new_n6214_), .B2(new_n6211_), .ZN(new_n6219_));
  INV_X1     g06027(.I(new_n6088_), .ZN(new_n6220_));
  OAI21_X1   g06028(.A1(new_n6219_), .A2(new_n2728_), .B(new_n6220_), .ZN(new_n6221_));
  NAND2_X1   g06029(.A1(new_n6221_), .A2(new_n6218_), .ZN(new_n6222_));
  OAI22_X1   g06030(.A1(new_n6219_), .A2(new_n2728_), .B1(new_n6217_), .B2(new_n6215_), .ZN(new_n6223_));
  AOI21_X1   g06031(.A1(new_n6223_), .A2(\asqrt[46] ), .B(new_n6095_), .ZN(new_n6224_));
  NOR2_X1    g06032(.A1(new_n6224_), .A2(new_n6222_), .ZN(new_n6225_));
  AOI22_X1   g06033(.A1(new_n6223_), .A2(\asqrt[46] ), .B1(new_n6221_), .B2(new_n6218_), .ZN(new_n6226_));
  INV_X1     g06034(.I(new_n6103_), .ZN(new_n6227_));
  OAI21_X1   g06035(.A1(new_n6226_), .A2(new_n2253_), .B(new_n6227_), .ZN(new_n6228_));
  NAND2_X1   g06036(.A1(new_n6228_), .A2(new_n6225_), .ZN(new_n6229_));
  OAI22_X1   g06037(.A1(new_n6226_), .A2(new_n2253_), .B1(new_n6224_), .B2(new_n6222_), .ZN(new_n6230_));
  AOI21_X1   g06038(.A1(new_n6230_), .A2(\asqrt[48] ), .B(new_n6110_), .ZN(new_n6231_));
  NOR2_X1    g06039(.A1(new_n6231_), .A2(new_n6229_), .ZN(new_n6232_));
  AOI22_X1   g06040(.A1(new_n6230_), .A2(\asqrt[48] ), .B1(new_n6228_), .B2(new_n6225_), .ZN(new_n6233_));
  INV_X1     g06041(.I(new_n6118_), .ZN(new_n6234_));
  OAI21_X1   g06042(.A1(new_n6233_), .A2(new_n1854_), .B(new_n6234_), .ZN(new_n6235_));
  NAND2_X1   g06043(.A1(new_n6235_), .A2(new_n6232_), .ZN(new_n6236_));
  OAI22_X1   g06044(.A1(new_n6233_), .A2(new_n1854_), .B1(new_n6231_), .B2(new_n6229_), .ZN(new_n6237_));
  AOI21_X1   g06045(.A1(new_n6237_), .A2(\asqrt[50] ), .B(new_n6125_), .ZN(new_n6238_));
  NOR2_X1    g06046(.A1(new_n6238_), .A2(new_n6236_), .ZN(new_n6239_));
  AOI22_X1   g06047(.A1(new_n6237_), .A2(\asqrt[50] ), .B1(new_n6235_), .B2(new_n6232_), .ZN(new_n6240_));
  INV_X1     g06048(.I(new_n6133_), .ZN(new_n6241_));
  OAI21_X1   g06049(.A1(new_n6240_), .A2(new_n1436_), .B(new_n6241_), .ZN(new_n6242_));
  NAND2_X1   g06050(.A1(new_n6242_), .A2(new_n6239_), .ZN(new_n6243_));
  OAI22_X1   g06051(.A1(new_n6240_), .A2(new_n1436_), .B1(new_n6238_), .B2(new_n6236_), .ZN(new_n6244_));
  AOI21_X1   g06052(.A1(new_n6244_), .A2(\asqrt[52] ), .B(new_n6140_), .ZN(new_n6245_));
  NOR2_X1    g06053(.A1(new_n6245_), .A2(new_n6243_), .ZN(new_n6246_));
  AOI22_X1   g06054(.A1(new_n6244_), .A2(\asqrt[52] ), .B1(new_n6242_), .B2(new_n6239_), .ZN(new_n6247_));
  INV_X1     g06055(.I(new_n6148_), .ZN(new_n6248_));
  OAI21_X1   g06056(.A1(new_n6247_), .A2(new_n1096_), .B(new_n6248_), .ZN(new_n6249_));
  NAND2_X1   g06057(.A1(new_n6249_), .A2(new_n6246_), .ZN(new_n6250_));
  OAI22_X1   g06058(.A1(new_n6247_), .A2(new_n1096_), .B1(new_n6245_), .B2(new_n6243_), .ZN(new_n6251_));
  AOI21_X1   g06059(.A1(new_n6251_), .A2(\asqrt[54] ), .B(new_n6155_), .ZN(new_n6252_));
  NOR2_X1    g06060(.A1(new_n6252_), .A2(new_n6250_), .ZN(new_n6253_));
  AOI22_X1   g06061(.A1(new_n6251_), .A2(\asqrt[54] ), .B1(new_n6249_), .B2(new_n6246_), .ZN(new_n6254_));
  INV_X1     g06062(.I(new_n6163_), .ZN(new_n6255_));
  OAI21_X1   g06063(.A1(new_n6254_), .A2(new_n825_), .B(new_n6255_), .ZN(new_n6256_));
  NAND2_X1   g06064(.A1(new_n6256_), .A2(new_n6253_), .ZN(new_n6257_));
  OAI22_X1   g06065(.A1(new_n6254_), .A2(new_n825_), .B1(new_n6252_), .B2(new_n6250_), .ZN(new_n6258_));
  AOI21_X1   g06066(.A1(new_n6258_), .A2(\asqrt[56] ), .B(new_n6170_), .ZN(new_n6259_));
  NOR2_X1    g06067(.A1(new_n6259_), .A2(new_n6257_), .ZN(new_n6260_));
  AOI22_X1   g06068(.A1(new_n6258_), .A2(\asqrt[56] ), .B1(new_n6256_), .B2(new_n6253_), .ZN(new_n6261_));
  OAI21_X1   g06069(.A1(new_n6261_), .A2(new_n587_), .B(new_n6182_), .ZN(new_n6262_));
  NAND2_X1   g06070(.A1(new_n6262_), .A2(new_n6260_), .ZN(new_n6263_));
  NAND2_X1   g06071(.A1(new_n6251_), .A2(\asqrt[54] ), .ZN(new_n6264_));
  AOI21_X1   g06072(.A1(new_n6264_), .A2(new_n6250_), .B(new_n825_), .ZN(new_n6265_));
  OAI21_X1   g06073(.A1(new_n6253_), .A2(new_n6265_), .B(\asqrt[56] ), .ZN(new_n6266_));
  AOI21_X1   g06074(.A1(new_n6257_), .A2(new_n6266_), .B(new_n587_), .ZN(new_n6267_));
  OAI21_X1   g06075(.A1(new_n6260_), .A2(new_n6267_), .B(\asqrt[58] ), .ZN(new_n6268_));
  NAND2_X1   g06076(.A1(new_n6263_), .A2(new_n6268_), .ZN(new_n6269_));
  AOI22_X1   g06077(.A1(new_n6269_), .A2(\asqrt[59] ), .B1(new_n6190_), .B2(new_n6183_), .ZN(new_n6270_));
  NOR4_X1    g06078(.A1(new_n5991_), .A2(\asqrt[60] ), .A3(new_n5811_), .A4(new_n5916_), .ZN(new_n6271_));
  XOR2_X1    g06079(.A1(new_n6271_), .A2(new_n5957_), .Z(new_n6272_));
  NAND2_X1   g06080(.A1(new_n6272_), .A2(new_n229_), .ZN(new_n6273_));
  INV_X1     g06081(.I(new_n6273_), .ZN(new_n6274_));
  OAI21_X1   g06082(.A1(new_n6270_), .A2(new_n275_), .B(new_n6274_), .ZN(new_n6275_));
  OAI22_X1   g06083(.A1(new_n6261_), .A2(new_n587_), .B1(new_n6259_), .B2(new_n6257_), .ZN(new_n6276_));
  AOI21_X1   g06084(.A1(new_n6276_), .A2(\asqrt[58] ), .B(new_n6188_), .ZN(new_n6277_));
  NOR2_X1    g06085(.A1(new_n6277_), .A2(new_n6263_), .ZN(new_n6278_));
  AOI22_X1   g06086(.A1(new_n6276_), .A2(\asqrt[58] ), .B1(new_n6262_), .B2(new_n6260_), .ZN(new_n6279_));
  OAI21_X1   g06087(.A1(new_n6279_), .A2(new_n376_), .B(new_n6196_), .ZN(new_n6280_));
  NAND2_X1   g06088(.A1(new_n6280_), .A2(new_n6278_), .ZN(new_n6281_));
  AOI21_X1   g06089(.A1(new_n6263_), .A2(new_n6268_), .B(new_n376_), .ZN(new_n6282_));
  OAI21_X1   g06090(.A1(new_n6278_), .A2(new_n6282_), .B(\asqrt[60] ), .ZN(new_n6283_));
  AOI21_X1   g06091(.A1(new_n6281_), .A2(new_n6283_), .B(new_n229_), .ZN(new_n6284_));
  INV_X1     g06092(.I(new_n5961_), .ZN(new_n6285_));
  NOR2_X1    g06093(.A1(new_n6285_), .A2(\asqrt[62] ), .ZN(new_n6286_));
  INV_X1     g06094(.I(new_n6286_), .ZN(new_n6287_));
  NAND4_X1   g06095(.A1(new_n6284_), .A2(new_n6197_), .A3(new_n6275_), .A4(new_n6287_), .ZN(new_n6288_));
  NAND2_X1   g06096(.A1(new_n5979_), .A2(new_n5927_), .ZN(new_n6289_));
  OAI21_X1   g06097(.A1(\asqrt[34] ), .A2(new_n6289_), .B(new_n5939_), .ZN(new_n6290_));
  NAND2_X1   g06098(.A1(new_n6290_), .A2(new_n231_), .ZN(new_n6291_));
  INV_X1     g06099(.I(new_n6291_), .ZN(new_n6292_));
  NAND3_X1   g06100(.A1(new_n6288_), .A2(new_n5963_), .A3(new_n6292_), .ZN(new_n6293_));
  OAI22_X1   g06101(.A1(new_n6279_), .A2(new_n376_), .B1(new_n6277_), .B2(new_n6263_), .ZN(new_n6294_));
  AOI21_X1   g06102(.A1(new_n6294_), .A2(\asqrt[60] ), .B(new_n6273_), .ZN(new_n6295_));
  AOI22_X1   g06103(.A1(new_n6294_), .A2(\asqrt[60] ), .B1(new_n6280_), .B2(new_n6278_), .ZN(new_n6296_));
  OAI22_X1   g06104(.A1(new_n6296_), .A2(new_n229_), .B1(new_n6295_), .B2(new_n6281_), .ZN(new_n6297_));
  NOR4_X1    g06105(.A1(new_n6297_), .A2(\asqrt[62] ), .A3(new_n5953_), .A4(new_n5961_), .ZN(new_n6298_));
  AOI21_X1   g06106(.A1(new_n5954_), .A2(new_n6293_), .B(new_n6298_), .ZN(new_n6299_));
  INV_X1     g06107(.I(\a[64] ), .ZN(new_n6300_));
  OAI21_X1   g06108(.A1(new_n5928_), .A2(new_n5939_), .B(\asqrt[34] ), .ZN(new_n6301_));
  XOR2_X1    g06109(.A1(new_n5939_), .A2(\asqrt[63] ), .Z(new_n6302_));
  NAND2_X1   g06110(.A1(new_n6301_), .A2(new_n6302_), .ZN(new_n6303_));
  INV_X1     g06111(.I(new_n6303_), .ZN(new_n6304_));
  NAND3_X1   g06112(.A1(new_n5985_), .A2(new_n5921_), .A3(new_n5928_), .ZN(new_n6305_));
  INV_X1     g06113(.I(new_n6305_), .ZN(new_n6306_));
  NOR2_X1    g06114(.A1(new_n6304_), .A2(new_n6306_), .ZN(new_n6307_));
  NOR2_X1    g06115(.A1(\a[62] ), .A2(\a[63] ), .ZN(new_n6308_));
  INV_X1     g06116(.I(new_n6308_), .ZN(new_n6309_));
  NOR3_X1    g06117(.A1(new_n6307_), .A2(new_n6300_), .A3(new_n6309_), .ZN(new_n6310_));
  NAND2_X1   g06118(.A1(new_n6299_), .A2(new_n6310_), .ZN(new_n6311_));
  XOR2_X1    g06119(.A1(new_n6311_), .A2(\a[65] ), .Z(new_n6312_));
  INV_X1     g06120(.I(\a[65] ), .ZN(new_n6313_));
  NAND2_X1   g06121(.A1(new_n6275_), .A2(new_n6197_), .ZN(new_n6314_));
  NAND2_X1   g06122(.A1(new_n6284_), .A2(new_n6287_), .ZN(new_n6315_));
  OAI21_X1   g06123(.A1(new_n6315_), .A2(new_n6314_), .B(new_n5963_), .ZN(new_n6316_));
  OAI21_X1   g06124(.A1(new_n6316_), .A2(new_n6291_), .B(new_n5954_), .ZN(new_n6317_));
  NAND2_X1   g06125(.A1(new_n6298_), .A2(new_n6304_), .ZN(new_n6318_));
  NOR2_X1    g06126(.A1(new_n6318_), .A2(new_n6317_), .ZN(new_n6319_));
  NAND3_X1   g06127(.A1(new_n6319_), .A2(new_n5954_), .A3(new_n6305_), .ZN(new_n6320_));
  NAND2_X1   g06128(.A1(new_n6281_), .A2(new_n6283_), .ZN(new_n6321_));
  AOI22_X1   g06129(.A1(new_n6321_), .A2(\asqrt[61] ), .B1(new_n6275_), .B2(new_n6197_), .ZN(new_n6322_));
  NOR2_X1    g06130(.A1(new_n6322_), .A2(new_n196_), .ZN(new_n6323_));
  AOI21_X1   g06131(.A1(new_n6191_), .A2(new_n6193_), .B(new_n275_), .ZN(new_n6324_));
  OAI21_X1   g06132(.A1(new_n6197_), .A2(new_n6324_), .B(\asqrt[61] ), .ZN(new_n6325_));
  NAND4_X1   g06133(.A1(new_n6314_), .A2(new_n196_), .A3(new_n6325_), .A4(new_n6285_), .ZN(new_n6326_));
  INV_X1     g06134(.I(new_n6326_), .ZN(new_n6327_));
  NOR3_X1    g06135(.A1(new_n6318_), .A2(new_n6317_), .A3(new_n6305_), .ZN(\asqrt[33] ));
  NAND3_X1   g06136(.A1(\asqrt[33] ), .A2(new_n6323_), .A3(new_n6327_), .ZN(new_n6329_));
  OAI21_X1   g06137(.A1(new_n6297_), .A2(\asqrt[62] ), .B(new_n5961_), .ZN(new_n6330_));
  OAI21_X1   g06138(.A1(\asqrt[33] ), .A2(new_n6330_), .B(new_n6323_), .ZN(new_n6331_));
  NAND2_X1   g06139(.A1(new_n6331_), .A2(new_n6329_), .ZN(new_n6332_));
  INV_X1     g06140(.I(new_n6332_), .ZN(new_n6333_));
  NOR3_X1    g06141(.A1(new_n6321_), .A2(\asqrt[61] ), .A3(new_n6272_), .ZN(new_n6334_));
  NAND2_X1   g06142(.A1(\asqrt[33] ), .A2(new_n6334_), .ZN(new_n6335_));
  XOR2_X1    g06143(.A1(new_n6335_), .A2(new_n6284_), .Z(new_n6336_));
  NOR2_X1    g06144(.A1(new_n6336_), .A2(new_n196_), .ZN(new_n6337_));
  INV_X1     g06145(.I(new_n6337_), .ZN(new_n6338_));
  INV_X1     g06146(.I(\a[66] ), .ZN(new_n6339_));
  NOR2_X1    g06147(.A1(\a[64] ), .A2(\a[65] ), .ZN(new_n6340_));
  INV_X1     g06148(.I(new_n6340_), .ZN(new_n6341_));
  NOR3_X1    g06149(.A1(new_n5992_), .A2(new_n6339_), .A3(new_n6341_), .ZN(new_n6342_));
  NAND3_X1   g06150(.A1(new_n5943_), .A2(new_n5979_), .A3(new_n6342_), .ZN(new_n6343_));
  XOR2_X1    g06151(.A1(new_n6343_), .A2(\a[67] ), .Z(new_n6344_));
  INV_X1     g06152(.I(\a[67] ), .ZN(new_n6345_));
  NOR4_X1    g06153(.A1(new_n6318_), .A2(new_n6317_), .A3(new_n6345_), .A4(new_n6305_), .ZN(new_n6346_));
  NOR2_X1    g06154(.A1(new_n6344_), .A2(\a[66] ), .ZN(new_n6347_));
  OAI21_X1   g06155(.A1(new_n6346_), .A2(new_n6347_), .B(new_n6344_), .ZN(new_n6348_));
  INV_X1     g06156(.I(new_n6344_), .ZN(new_n6349_));
  NOR2_X1    g06157(.A1(new_n6295_), .A2(new_n6281_), .ZN(new_n6350_));
  NOR3_X1    g06158(.A1(new_n6296_), .A2(new_n229_), .A3(new_n6286_), .ZN(new_n6351_));
  AOI21_X1   g06159(.A1(new_n6351_), .A2(new_n6350_), .B(new_n5962_), .ZN(new_n6352_));
  AOI21_X1   g06160(.A1(new_n6352_), .A2(new_n6292_), .B(new_n5953_), .ZN(new_n6353_));
  AOI21_X1   g06161(.A1(new_n6297_), .A2(\asqrt[62] ), .B(new_n5954_), .ZN(new_n6354_));
  NOR3_X1    g06162(.A1(new_n6354_), .A2(new_n6326_), .A3(new_n6303_), .ZN(new_n6355_));
  NAND4_X1   g06163(.A1(new_n6355_), .A2(\a[67] ), .A3(new_n6353_), .A4(new_n6306_), .ZN(new_n6356_));
  NAND3_X1   g06164(.A1(new_n6356_), .A2(\a[66] ), .A3(new_n6349_), .ZN(new_n6357_));
  NAND2_X1   g06165(.A1(new_n6348_), .A2(new_n6357_), .ZN(new_n6358_));
  NAND2_X1   g06166(.A1(new_n5977_), .A2(new_n5941_), .ZN(new_n6359_));
  NAND4_X1   g06167(.A1(new_n5981_), .A2(new_n5975_), .A3(new_n5928_), .A4(new_n6359_), .ZN(new_n6360_));
  NOR2_X1    g06168(.A1(new_n5991_), .A2(new_n6339_), .ZN(new_n6361_));
  XOR2_X1    g06169(.A1(new_n6361_), .A2(new_n6360_), .Z(new_n6362_));
  NOR2_X1    g06170(.A1(new_n6362_), .A2(new_n6341_), .ZN(new_n6363_));
  INV_X1     g06171(.I(new_n6363_), .ZN(new_n6364_));
  NAND3_X1   g06172(.A1(new_n6355_), .A2(new_n6353_), .A3(new_n6306_), .ZN(new_n6365_));
  NOR4_X1    g06173(.A1(new_n6325_), .A2(new_n6281_), .A3(new_n6295_), .A4(new_n6286_), .ZN(new_n6366_));
  NOR3_X1    g06174(.A1(new_n6366_), .A2(new_n5962_), .A3(new_n6291_), .ZN(new_n6367_));
  NAND4_X1   g06175(.A1(new_n6322_), .A2(new_n196_), .A3(new_n5954_), .A4(new_n6285_), .ZN(new_n6368_));
  OAI21_X1   g06176(.A1(new_n6367_), .A2(new_n5953_), .B(new_n6368_), .ZN(new_n6369_));
  NAND2_X1   g06177(.A1(new_n6307_), .A2(\asqrt[34] ), .ZN(new_n6370_));
  OAI21_X1   g06178(.A1(new_n6369_), .A2(new_n6370_), .B(new_n5964_), .ZN(new_n6371_));
  NAND3_X1   g06179(.A1(new_n6371_), .A2(new_n5965_), .A3(new_n6365_), .ZN(new_n6372_));
  INV_X1     g06180(.I(new_n6370_), .ZN(new_n6373_));
  AOI21_X1   g06181(.A1(new_n6299_), .A2(new_n6373_), .B(\a[68] ), .ZN(new_n6374_));
  OAI21_X1   g06182(.A1(new_n6374_), .A2(new_n5966_), .B(\asqrt[33] ), .ZN(new_n6375_));
  NAND4_X1   g06183(.A1(new_n6372_), .A2(new_n6375_), .A3(new_n5626_), .A4(new_n6364_), .ZN(new_n6376_));
  NAND2_X1   g06184(.A1(new_n6376_), .A2(new_n6358_), .ZN(new_n6377_));
  NAND3_X1   g06185(.A1(new_n6348_), .A2(new_n6357_), .A3(new_n6364_), .ZN(new_n6378_));
  AOI21_X1   g06186(.A1(\asqrt[34] ), .A2(new_n5964_), .B(\a[69] ), .ZN(new_n6379_));
  NOR2_X1    g06187(.A1(new_n5982_), .A2(\a[68] ), .ZN(new_n6380_));
  AOI21_X1   g06188(.A1(\asqrt[34] ), .A2(\a[68] ), .B(new_n5968_), .ZN(new_n6381_));
  OAI21_X1   g06189(.A1(new_n6379_), .A2(new_n6380_), .B(new_n6381_), .ZN(new_n6382_));
  INV_X1     g06190(.I(new_n6382_), .ZN(new_n6383_));
  NAND3_X1   g06191(.A1(\asqrt[33] ), .A2(new_n5990_), .A3(new_n6383_), .ZN(new_n6384_));
  OAI21_X1   g06192(.A1(new_n6365_), .A2(new_n6382_), .B(new_n5989_), .ZN(new_n6385_));
  NAND3_X1   g06193(.A1(new_n6384_), .A2(new_n6385_), .A3(new_n5273_), .ZN(new_n6386_));
  AOI21_X1   g06194(.A1(new_n6378_), .A2(\asqrt[35] ), .B(new_n6386_), .ZN(new_n6387_));
  NOR2_X1    g06195(.A1(new_n6377_), .A2(new_n6387_), .ZN(new_n6388_));
  AOI22_X1   g06196(.A1(new_n6376_), .A2(new_n6358_), .B1(\asqrt[35] ), .B2(new_n6378_), .ZN(new_n6389_));
  INV_X1     g06197(.I(new_n5972_), .ZN(new_n6390_));
  AOI21_X1   g06198(.A1(new_n5982_), .A2(new_n6390_), .B(new_n5974_), .ZN(new_n6391_));
  INV_X1     g06199(.I(new_n5983_), .ZN(new_n6392_));
  NOR3_X1    g06200(.A1(new_n6392_), .A2(new_n6391_), .A3(new_n5989_), .ZN(new_n6393_));
  AOI21_X1   g06201(.A1(new_n6000_), .A2(new_n5997_), .B(\asqrt[36] ), .ZN(new_n6394_));
  AND4_X2    g06202(.A1(new_n6393_), .A2(\asqrt[33] ), .A3(new_n6014_), .A4(new_n6394_), .Z(new_n6395_));
  NOR2_X1    g06203(.A1(new_n6393_), .A2(new_n5273_), .ZN(new_n6396_));
  NOR3_X1    g06204(.A1(new_n6395_), .A2(\asqrt[37] ), .A3(new_n6396_), .ZN(new_n6397_));
  OAI21_X1   g06205(.A1(new_n6389_), .A2(new_n5273_), .B(new_n6397_), .ZN(new_n6398_));
  NAND2_X1   g06206(.A1(new_n6398_), .A2(new_n6388_), .ZN(new_n6399_));
  OAI22_X1   g06207(.A1(new_n6389_), .A2(new_n5273_), .B1(new_n6377_), .B2(new_n6387_), .ZN(new_n6400_));
  NAND2_X1   g06208(.A1(new_n6009_), .A2(new_n6010_), .ZN(new_n6401_));
  NAND4_X1   g06209(.A1(\asqrt[33] ), .A2(new_n4973_), .A3(new_n6401_), .A4(new_n6022_), .ZN(new_n6402_));
  XOR2_X1    g06210(.A1(new_n6402_), .A2(new_n6015_), .Z(new_n6403_));
  NAND2_X1   g06211(.A1(new_n6403_), .A2(new_n4645_), .ZN(new_n6404_));
  AOI21_X1   g06212(.A1(new_n6400_), .A2(\asqrt[37] ), .B(new_n6404_), .ZN(new_n6405_));
  NOR2_X1    g06213(.A1(new_n6405_), .A2(new_n6399_), .ZN(new_n6406_));
  AOI22_X1   g06214(.A1(new_n6400_), .A2(\asqrt[37] ), .B1(new_n6398_), .B2(new_n6388_), .ZN(new_n6407_));
  NOR4_X1    g06215(.A1(new_n6365_), .A2(\asqrt[38] ), .A3(new_n6019_), .A4(new_n6023_), .ZN(new_n6408_));
  XOR2_X1    g06216(.A1(new_n6408_), .A2(new_n6030_), .Z(new_n6409_));
  NAND2_X1   g06217(.A1(new_n6409_), .A2(new_n4330_), .ZN(new_n6410_));
  INV_X1     g06218(.I(new_n6410_), .ZN(new_n6411_));
  OAI21_X1   g06219(.A1(new_n6407_), .A2(new_n4645_), .B(new_n6411_), .ZN(new_n6412_));
  NAND2_X1   g06220(.A1(new_n6412_), .A2(new_n6406_), .ZN(new_n6413_));
  OAI22_X1   g06221(.A1(new_n6407_), .A2(new_n4645_), .B1(new_n6405_), .B2(new_n6399_), .ZN(new_n6414_));
  NOR2_X1    g06222(.A1(new_n6027_), .A2(\asqrt[39] ), .ZN(new_n6415_));
  NAND3_X1   g06223(.A1(\asqrt[33] ), .A2(new_n6200_), .A3(new_n6415_), .ZN(new_n6416_));
  XOR2_X1    g06224(.A1(new_n6416_), .A2(new_n6031_), .Z(new_n6417_));
  NAND2_X1   g06225(.A1(new_n6417_), .A2(new_n4018_), .ZN(new_n6418_));
  AOI21_X1   g06226(.A1(new_n6414_), .A2(\asqrt[39] ), .B(new_n6418_), .ZN(new_n6419_));
  NOR2_X1    g06227(.A1(new_n6419_), .A2(new_n6413_), .ZN(new_n6420_));
  AOI22_X1   g06228(.A1(new_n6414_), .A2(\asqrt[39] ), .B1(new_n6412_), .B2(new_n6406_), .ZN(new_n6421_));
  NOR4_X1    g06229(.A1(new_n6365_), .A2(\asqrt[40] ), .A3(new_n6036_), .A4(new_n6203_), .ZN(new_n6422_));
  XOR2_X1    g06230(.A1(new_n6422_), .A2(new_n6042_), .Z(new_n6423_));
  NAND2_X1   g06231(.A1(new_n6423_), .A2(new_n3760_), .ZN(new_n6424_));
  INV_X1     g06232(.I(new_n6424_), .ZN(new_n6425_));
  OAI21_X1   g06233(.A1(new_n6421_), .A2(new_n4018_), .B(new_n6425_), .ZN(new_n6426_));
  NAND2_X1   g06234(.A1(new_n6426_), .A2(new_n6420_), .ZN(new_n6427_));
  OAI22_X1   g06235(.A1(new_n6421_), .A2(new_n4018_), .B1(new_n6419_), .B2(new_n6413_), .ZN(new_n6428_));
  NOR4_X1    g06236(.A1(new_n6365_), .A2(\asqrt[41] ), .A3(new_n6045_), .A4(new_n6051_), .ZN(new_n6429_));
  XNOR2_X1   g06237(.A1(new_n6429_), .A2(new_n6059_), .ZN(new_n6430_));
  NAND2_X1   g06238(.A1(new_n6430_), .A2(new_n3481_), .ZN(new_n6431_));
  AOI21_X1   g06239(.A1(new_n6428_), .A2(\asqrt[41] ), .B(new_n6431_), .ZN(new_n6432_));
  NOR2_X1    g06240(.A1(new_n6432_), .A2(new_n6427_), .ZN(new_n6433_));
  AOI22_X1   g06241(.A1(new_n6428_), .A2(\asqrt[41] ), .B1(new_n6426_), .B2(new_n6420_), .ZN(new_n6434_));
  NOR4_X1    g06242(.A1(new_n6365_), .A2(\asqrt[42] ), .A3(new_n6054_), .A4(new_n6209_), .ZN(new_n6435_));
  XOR2_X1    g06243(.A1(new_n6435_), .A2(new_n6060_), .Z(new_n6436_));
  NAND2_X1   g06244(.A1(new_n6436_), .A2(new_n3208_), .ZN(new_n6437_));
  INV_X1     g06245(.I(new_n6437_), .ZN(new_n6438_));
  OAI21_X1   g06246(.A1(new_n6434_), .A2(new_n3481_), .B(new_n6438_), .ZN(new_n6439_));
  NAND2_X1   g06247(.A1(new_n6439_), .A2(new_n6433_), .ZN(new_n6440_));
  OAI22_X1   g06248(.A1(new_n6434_), .A2(new_n3481_), .B1(new_n6432_), .B2(new_n6427_), .ZN(new_n6441_));
  NAND2_X1   g06249(.A1(new_n6069_), .A2(\asqrt[43] ), .ZN(new_n6442_));
  NOR4_X1    g06250(.A1(new_n6365_), .A2(\asqrt[43] ), .A3(new_n6063_), .A4(new_n6069_), .ZN(new_n6443_));
  XOR2_X1    g06251(.A1(new_n6443_), .A2(new_n6442_), .Z(new_n6444_));
  NAND2_X1   g06252(.A1(new_n6444_), .A2(new_n2941_), .ZN(new_n6445_));
  AOI21_X1   g06253(.A1(new_n6441_), .A2(\asqrt[43] ), .B(new_n6445_), .ZN(new_n6446_));
  NOR2_X1    g06254(.A1(new_n6446_), .A2(new_n6440_), .ZN(new_n6447_));
  AOI22_X1   g06255(.A1(new_n6441_), .A2(\asqrt[43] ), .B1(new_n6439_), .B2(new_n6433_), .ZN(new_n6448_));
  NAND2_X1   g06256(.A1(new_n6216_), .A2(\asqrt[44] ), .ZN(new_n6449_));
  NOR4_X1    g06257(.A1(new_n6365_), .A2(\asqrt[44] ), .A3(new_n6072_), .A4(new_n6216_), .ZN(new_n6450_));
  XOR2_X1    g06258(.A1(new_n6450_), .A2(new_n6449_), .Z(new_n6451_));
  NAND2_X1   g06259(.A1(new_n6451_), .A2(new_n2728_), .ZN(new_n6452_));
  INV_X1     g06260(.I(new_n6452_), .ZN(new_n6453_));
  OAI21_X1   g06261(.A1(new_n6448_), .A2(new_n2941_), .B(new_n6453_), .ZN(new_n6454_));
  NAND2_X1   g06262(.A1(new_n6454_), .A2(new_n6447_), .ZN(new_n6455_));
  OAI22_X1   g06263(.A1(new_n6448_), .A2(new_n2941_), .B1(new_n6446_), .B2(new_n6440_), .ZN(new_n6456_));
  NAND2_X1   g06264(.A1(new_n6084_), .A2(\asqrt[45] ), .ZN(new_n6457_));
  NOR4_X1    g06265(.A1(new_n6365_), .A2(\asqrt[45] ), .A3(new_n6079_), .A4(new_n6084_), .ZN(new_n6458_));
  XOR2_X1    g06266(.A1(new_n6458_), .A2(new_n6457_), .Z(new_n6459_));
  NAND2_X1   g06267(.A1(new_n6459_), .A2(new_n2488_), .ZN(new_n6460_));
  AOI21_X1   g06268(.A1(new_n6456_), .A2(\asqrt[45] ), .B(new_n6460_), .ZN(new_n6461_));
  NOR2_X1    g06269(.A1(new_n6461_), .A2(new_n6455_), .ZN(new_n6462_));
  AOI22_X1   g06270(.A1(new_n6456_), .A2(\asqrt[45] ), .B1(new_n6454_), .B2(new_n6447_), .ZN(new_n6463_));
  NAND2_X1   g06271(.A1(new_n6223_), .A2(\asqrt[46] ), .ZN(new_n6464_));
  NOR4_X1    g06272(.A1(new_n6365_), .A2(\asqrt[46] ), .A3(new_n6087_), .A4(new_n6223_), .ZN(new_n6465_));
  XOR2_X1    g06273(.A1(new_n6465_), .A2(new_n6464_), .Z(new_n6466_));
  NAND2_X1   g06274(.A1(new_n6466_), .A2(new_n2253_), .ZN(new_n6467_));
  INV_X1     g06275(.I(new_n6467_), .ZN(new_n6468_));
  OAI21_X1   g06276(.A1(new_n6463_), .A2(new_n2488_), .B(new_n6468_), .ZN(new_n6469_));
  NAND2_X1   g06277(.A1(new_n6469_), .A2(new_n6462_), .ZN(new_n6470_));
  OAI22_X1   g06278(.A1(new_n6463_), .A2(new_n2488_), .B1(new_n6461_), .B2(new_n6455_), .ZN(new_n6471_));
  NAND2_X1   g06279(.A1(new_n6099_), .A2(\asqrt[47] ), .ZN(new_n6472_));
  NOR4_X1    g06280(.A1(new_n6365_), .A2(\asqrt[47] ), .A3(new_n6094_), .A4(new_n6099_), .ZN(new_n6473_));
  XOR2_X1    g06281(.A1(new_n6473_), .A2(new_n6472_), .Z(new_n6474_));
  NAND2_X1   g06282(.A1(new_n6474_), .A2(new_n2046_), .ZN(new_n6475_));
  AOI21_X1   g06283(.A1(new_n6471_), .A2(\asqrt[47] ), .B(new_n6475_), .ZN(new_n6476_));
  NOR2_X1    g06284(.A1(new_n6476_), .A2(new_n6470_), .ZN(new_n6477_));
  AOI22_X1   g06285(.A1(new_n6471_), .A2(\asqrt[47] ), .B1(new_n6469_), .B2(new_n6462_), .ZN(new_n6478_));
  NAND2_X1   g06286(.A1(new_n6230_), .A2(\asqrt[48] ), .ZN(new_n6479_));
  NOR4_X1    g06287(.A1(new_n6365_), .A2(\asqrt[48] ), .A3(new_n6102_), .A4(new_n6230_), .ZN(new_n6480_));
  XOR2_X1    g06288(.A1(new_n6480_), .A2(new_n6479_), .Z(new_n6481_));
  NAND2_X1   g06289(.A1(new_n6481_), .A2(new_n1854_), .ZN(new_n6482_));
  INV_X1     g06290(.I(new_n6482_), .ZN(new_n6483_));
  OAI21_X1   g06291(.A1(new_n6478_), .A2(new_n2046_), .B(new_n6483_), .ZN(new_n6484_));
  NAND2_X1   g06292(.A1(new_n6484_), .A2(new_n6477_), .ZN(new_n6485_));
  OAI22_X1   g06293(.A1(new_n6478_), .A2(new_n2046_), .B1(new_n6476_), .B2(new_n6470_), .ZN(new_n6486_));
  NAND2_X1   g06294(.A1(new_n6114_), .A2(\asqrt[49] ), .ZN(new_n6487_));
  NOR4_X1    g06295(.A1(new_n6365_), .A2(\asqrt[49] ), .A3(new_n6109_), .A4(new_n6114_), .ZN(new_n6488_));
  XOR2_X1    g06296(.A1(new_n6488_), .A2(new_n6487_), .Z(new_n6489_));
  NAND2_X1   g06297(.A1(new_n6489_), .A2(new_n1595_), .ZN(new_n6490_));
  AOI21_X1   g06298(.A1(new_n6486_), .A2(\asqrt[49] ), .B(new_n6490_), .ZN(new_n6491_));
  NOR2_X1    g06299(.A1(new_n6491_), .A2(new_n6485_), .ZN(new_n6492_));
  AOI22_X1   g06300(.A1(new_n6486_), .A2(\asqrt[49] ), .B1(new_n6484_), .B2(new_n6477_), .ZN(new_n6493_));
  NAND2_X1   g06301(.A1(new_n6237_), .A2(\asqrt[50] ), .ZN(new_n6494_));
  NOR4_X1    g06302(.A1(new_n6365_), .A2(\asqrt[50] ), .A3(new_n6117_), .A4(new_n6237_), .ZN(new_n6495_));
  XOR2_X1    g06303(.A1(new_n6495_), .A2(new_n6494_), .Z(new_n6496_));
  NAND2_X1   g06304(.A1(new_n6496_), .A2(new_n1436_), .ZN(new_n6497_));
  INV_X1     g06305(.I(new_n6497_), .ZN(new_n6498_));
  OAI21_X1   g06306(.A1(new_n6493_), .A2(new_n1595_), .B(new_n6498_), .ZN(new_n6499_));
  NAND2_X1   g06307(.A1(new_n6499_), .A2(new_n6492_), .ZN(new_n6500_));
  OAI22_X1   g06308(.A1(new_n6493_), .A2(new_n1595_), .B1(new_n6491_), .B2(new_n6485_), .ZN(new_n6501_));
  NAND2_X1   g06309(.A1(new_n6129_), .A2(\asqrt[51] ), .ZN(new_n6502_));
  NOR4_X1    g06310(.A1(new_n6365_), .A2(\asqrt[51] ), .A3(new_n6124_), .A4(new_n6129_), .ZN(new_n6503_));
  XOR2_X1    g06311(.A1(new_n6503_), .A2(new_n6502_), .Z(new_n6504_));
  NAND2_X1   g06312(.A1(new_n6504_), .A2(new_n1260_), .ZN(new_n6505_));
  AOI21_X1   g06313(.A1(new_n6501_), .A2(\asqrt[51] ), .B(new_n6505_), .ZN(new_n6506_));
  NOR2_X1    g06314(.A1(new_n6506_), .A2(new_n6500_), .ZN(new_n6507_));
  AOI22_X1   g06315(.A1(new_n6501_), .A2(\asqrt[51] ), .B1(new_n6499_), .B2(new_n6492_), .ZN(new_n6508_));
  NAND2_X1   g06316(.A1(new_n6244_), .A2(\asqrt[52] ), .ZN(new_n6509_));
  NOR4_X1    g06317(.A1(new_n6365_), .A2(\asqrt[52] ), .A3(new_n6132_), .A4(new_n6244_), .ZN(new_n6510_));
  XOR2_X1    g06318(.A1(new_n6510_), .A2(new_n6509_), .Z(new_n6511_));
  NAND2_X1   g06319(.A1(new_n6511_), .A2(new_n1096_), .ZN(new_n6512_));
  INV_X1     g06320(.I(new_n6512_), .ZN(new_n6513_));
  OAI21_X1   g06321(.A1(new_n6508_), .A2(new_n1260_), .B(new_n6513_), .ZN(new_n6514_));
  NAND2_X1   g06322(.A1(new_n6514_), .A2(new_n6507_), .ZN(new_n6515_));
  OAI22_X1   g06323(.A1(new_n6508_), .A2(new_n1260_), .B1(new_n6506_), .B2(new_n6500_), .ZN(new_n6516_));
  NOR4_X1    g06324(.A1(new_n6365_), .A2(\asqrt[53] ), .A3(new_n6139_), .A4(new_n6144_), .ZN(new_n6517_));
  XOR2_X1    g06325(.A1(new_n6517_), .A2(new_n6174_), .Z(new_n6518_));
  NAND2_X1   g06326(.A1(new_n6518_), .A2(new_n970_), .ZN(new_n6519_));
  AOI21_X1   g06327(.A1(new_n6516_), .A2(\asqrt[53] ), .B(new_n6519_), .ZN(new_n6520_));
  NOR2_X1    g06328(.A1(new_n6520_), .A2(new_n6515_), .ZN(new_n6521_));
  AOI22_X1   g06329(.A1(new_n6516_), .A2(\asqrt[53] ), .B1(new_n6514_), .B2(new_n6507_), .ZN(new_n6522_));
  NOR4_X1    g06330(.A1(new_n6365_), .A2(\asqrt[54] ), .A3(new_n6147_), .A4(new_n6251_), .ZN(new_n6523_));
  XOR2_X1    g06331(.A1(new_n6523_), .A2(new_n6264_), .Z(new_n6524_));
  NAND2_X1   g06332(.A1(new_n6524_), .A2(new_n825_), .ZN(new_n6525_));
  INV_X1     g06333(.I(new_n6525_), .ZN(new_n6526_));
  OAI21_X1   g06334(.A1(new_n6522_), .A2(new_n970_), .B(new_n6526_), .ZN(new_n6527_));
  NAND2_X1   g06335(.A1(new_n6527_), .A2(new_n6521_), .ZN(new_n6528_));
  OAI22_X1   g06336(.A1(new_n6522_), .A2(new_n970_), .B1(new_n6520_), .B2(new_n6515_), .ZN(new_n6529_));
  NOR4_X1    g06337(.A1(new_n6365_), .A2(\asqrt[55] ), .A3(new_n6154_), .A4(new_n6159_), .ZN(new_n6530_));
  XOR2_X1    g06338(.A1(new_n6530_), .A2(new_n6176_), .Z(new_n6531_));
  NAND2_X1   g06339(.A1(new_n6531_), .A2(new_n724_), .ZN(new_n6532_));
  AOI21_X1   g06340(.A1(new_n6529_), .A2(\asqrt[55] ), .B(new_n6532_), .ZN(new_n6533_));
  NOR2_X1    g06341(.A1(new_n6533_), .A2(new_n6528_), .ZN(new_n6534_));
  AOI22_X1   g06342(.A1(new_n6529_), .A2(\asqrt[55] ), .B1(new_n6527_), .B2(new_n6521_), .ZN(new_n6535_));
  NOR4_X1    g06343(.A1(new_n6365_), .A2(\asqrt[56] ), .A3(new_n6162_), .A4(new_n6258_), .ZN(new_n6536_));
  XOR2_X1    g06344(.A1(new_n6536_), .A2(new_n6266_), .Z(new_n6537_));
  NAND2_X1   g06345(.A1(new_n6537_), .A2(new_n587_), .ZN(new_n6538_));
  INV_X1     g06346(.I(new_n6538_), .ZN(new_n6539_));
  OAI21_X1   g06347(.A1(new_n6535_), .A2(new_n724_), .B(new_n6539_), .ZN(new_n6540_));
  NAND2_X1   g06348(.A1(new_n6540_), .A2(new_n6534_), .ZN(new_n6541_));
  OAI22_X1   g06349(.A1(new_n6535_), .A2(new_n724_), .B1(new_n6533_), .B2(new_n6528_), .ZN(new_n6542_));
  NOR4_X1    g06350(.A1(new_n6365_), .A2(\asqrt[57] ), .A3(new_n6169_), .A4(new_n6184_), .ZN(new_n6543_));
  XOR2_X1    g06351(.A1(new_n6543_), .A2(new_n6178_), .Z(new_n6544_));
  NAND2_X1   g06352(.A1(new_n6544_), .A2(new_n504_), .ZN(new_n6545_));
  AOI21_X1   g06353(.A1(new_n6542_), .A2(\asqrt[57] ), .B(new_n6545_), .ZN(new_n6546_));
  NOR2_X1    g06354(.A1(new_n6546_), .A2(new_n6541_), .ZN(new_n6547_));
  AOI22_X1   g06355(.A1(new_n6542_), .A2(\asqrt[57] ), .B1(new_n6540_), .B2(new_n6534_), .ZN(new_n6548_));
  NOR4_X1    g06356(.A1(new_n6365_), .A2(\asqrt[58] ), .A3(new_n6180_), .A4(new_n6276_), .ZN(new_n6549_));
  XOR2_X1    g06357(.A1(new_n6549_), .A2(new_n6268_), .Z(new_n6550_));
  NAND2_X1   g06358(.A1(new_n6550_), .A2(new_n376_), .ZN(new_n6551_));
  INV_X1     g06359(.I(new_n6551_), .ZN(new_n6552_));
  OAI21_X1   g06360(.A1(new_n6548_), .A2(new_n504_), .B(new_n6552_), .ZN(new_n6553_));
  NAND2_X1   g06361(.A1(new_n6553_), .A2(new_n6547_), .ZN(new_n6554_));
  OAI22_X1   g06362(.A1(new_n6548_), .A2(new_n504_), .B1(new_n6546_), .B2(new_n6541_), .ZN(new_n6555_));
  NOR4_X1    g06363(.A1(new_n6365_), .A2(\asqrt[59] ), .A3(new_n6187_), .A4(new_n6269_), .ZN(new_n6556_));
  XOR2_X1    g06364(.A1(new_n6556_), .A2(new_n6193_), .Z(new_n6557_));
  NAND2_X1   g06365(.A1(new_n6557_), .A2(new_n275_), .ZN(new_n6558_));
  AOI21_X1   g06366(.A1(new_n6555_), .A2(\asqrt[59] ), .B(new_n6558_), .ZN(new_n6559_));
  NOR2_X1    g06367(.A1(new_n6559_), .A2(new_n6554_), .ZN(new_n6560_));
  AOI22_X1   g06368(.A1(new_n6555_), .A2(\asqrt[59] ), .B1(new_n6553_), .B2(new_n6547_), .ZN(new_n6561_));
  NOR4_X1    g06369(.A1(new_n6365_), .A2(\asqrt[60] ), .A3(new_n6195_), .A4(new_n6294_), .ZN(new_n6562_));
  XOR2_X1    g06370(.A1(new_n6562_), .A2(new_n6283_), .Z(new_n6563_));
  NAND2_X1   g06371(.A1(new_n6563_), .A2(new_n229_), .ZN(new_n6564_));
  INV_X1     g06372(.I(new_n6564_), .ZN(new_n6565_));
  OAI21_X1   g06373(.A1(new_n6561_), .A2(new_n275_), .B(new_n6565_), .ZN(new_n6566_));
  NAND2_X1   g06374(.A1(new_n6566_), .A2(new_n6560_), .ZN(new_n6567_));
  OAI22_X1   g06375(.A1(new_n6561_), .A2(new_n275_), .B1(new_n6559_), .B2(new_n6554_), .ZN(new_n6568_));
  INV_X1     g06376(.I(new_n6336_), .ZN(new_n6569_));
  NOR2_X1    g06377(.A1(new_n6569_), .A2(\asqrt[62] ), .ZN(new_n6570_));
  INV_X1     g06378(.I(new_n6570_), .ZN(new_n6571_));
  NAND3_X1   g06379(.A1(new_n6568_), .A2(\asqrt[61] ), .A3(new_n6571_), .ZN(new_n6572_));
  OAI21_X1   g06380(.A1(new_n6572_), .A2(new_n6567_), .B(new_n6338_), .ZN(new_n6573_));
  NAND3_X1   g06381(.A1(new_n6365_), .A2(new_n5953_), .A3(new_n6368_), .ZN(new_n6574_));
  AOI21_X1   g06382(.A1(new_n6574_), .A2(new_n6316_), .B(\asqrt[63] ), .ZN(new_n6575_));
  INV_X1     g06383(.I(new_n6575_), .ZN(new_n6576_));
  OAI21_X1   g06384(.A1(new_n6573_), .A2(new_n6576_), .B(new_n6333_), .ZN(new_n6577_));
  INV_X1     g06385(.I(new_n6347_), .ZN(new_n6578_));
  AOI21_X1   g06386(.A1(new_n6356_), .A2(new_n6578_), .B(new_n6349_), .ZN(new_n6579_));
  NOR3_X1    g06387(.A1(new_n6346_), .A2(new_n6339_), .A3(new_n6344_), .ZN(new_n6580_));
  NOR2_X1    g06388(.A1(new_n6580_), .A2(new_n6579_), .ZN(new_n6581_));
  NOR3_X1    g06389(.A1(new_n6374_), .A2(new_n5966_), .A3(\asqrt[33] ), .ZN(new_n6582_));
  AOI21_X1   g06390(.A1(new_n6371_), .A2(new_n5965_), .B(new_n6365_), .ZN(new_n6583_));
  NOR4_X1    g06391(.A1(new_n6583_), .A2(new_n6582_), .A3(\asqrt[35] ), .A4(new_n6363_), .ZN(new_n6584_));
  NOR2_X1    g06392(.A1(new_n6584_), .A2(new_n6581_), .ZN(new_n6585_));
  NOR3_X1    g06393(.A1(new_n6580_), .A2(new_n6579_), .A3(new_n6363_), .ZN(new_n6586_));
  NOR3_X1    g06394(.A1(new_n6365_), .A2(new_n5989_), .A3(new_n6382_), .ZN(new_n6587_));
  AOI21_X1   g06395(.A1(\asqrt[33] ), .A2(new_n6383_), .B(new_n5990_), .ZN(new_n6588_));
  NOR3_X1    g06396(.A1(new_n6588_), .A2(new_n6587_), .A3(\asqrt[36] ), .ZN(new_n6589_));
  OAI21_X1   g06397(.A1(new_n6586_), .A2(new_n5626_), .B(new_n6589_), .ZN(new_n6590_));
  NAND2_X1   g06398(.A1(new_n6585_), .A2(new_n6590_), .ZN(new_n6591_));
  OAI22_X1   g06399(.A1(new_n6584_), .A2(new_n6581_), .B1(new_n5626_), .B2(new_n6586_), .ZN(new_n6592_));
  INV_X1     g06400(.I(new_n6397_), .ZN(new_n6593_));
  AOI21_X1   g06401(.A1(new_n6592_), .A2(\asqrt[36] ), .B(new_n6593_), .ZN(new_n6594_));
  NOR2_X1    g06402(.A1(new_n6594_), .A2(new_n6591_), .ZN(new_n6595_));
  AOI22_X1   g06403(.A1(new_n6592_), .A2(\asqrt[36] ), .B1(new_n6585_), .B2(new_n6590_), .ZN(new_n6596_));
  INV_X1     g06404(.I(new_n6404_), .ZN(new_n6597_));
  OAI21_X1   g06405(.A1(new_n6596_), .A2(new_n4973_), .B(new_n6597_), .ZN(new_n6598_));
  NAND2_X1   g06406(.A1(new_n6598_), .A2(new_n6595_), .ZN(new_n6599_));
  OAI22_X1   g06407(.A1(new_n6596_), .A2(new_n4973_), .B1(new_n6594_), .B2(new_n6591_), .ZN(new_n6600_));
  AOI21_X1   g06408(.A1(new_n6600_), .A2(\asqrt[38] ), .B(new_n6410_), .ZN(new_n6601_));
  NOR2_X1    g06409(.A1(new_n6601_), .A2(new_n6599_), .ZN(new_n6602_));
  AOI22_X1   g06410(.A1(new_n6600_), .A2(\asqrt[38] ), .B1(new_n6598_), .B2(new_n6595_), .ZN(new_n6603_));
  INV_X1     g06411(.I(new_n6418_), .ZN(new_n6604_));
  OAI21_X1   g06412(.A1(new_n6603_), .A2(new_n4330_), .B(new_n6604_), .ZN(new_n6605_));
  NAND2_X1   g06413(.A1(new_n6605_), .A2(new_n6602_), .ZN(new_n6606_));
  OAI22_X1   g06414(.A1(new_n6603_), .A2(new_n4330_), .B1(new_n6601_), .B2(new_n6599_), .ZN(new_n6607_));
  AOI21_X1   g06415(.A1(new_n6607_), .A2(\asqrt[40] ), .B(new_n6424_), .ZN(new_n6608_));
  NOR2_X1    g06416(.A1(new_n6608_), .A2(new_n6606_), .ZN(new_n6609_));
  AOI22_X1   g06417(.A1(new_n6607_), .A2(\asqrt[40] ), .B1(new_n6605_), .B2(new_n6602_), .ZN(new_n6610_));
  INV_X1     g06418(.I(new_n6431_), .ZN(new_n6611_));
  OAI21_X1   g06419(.A1(new_n6610_), .A2(new_n3760_), .B(new_n6611_), .ZN(new_n6612_));
  NAND2_X1   g06420(.A1(new_n6612_), .A2(new_n6609_), .ZN(new_n6613_));
  OAI22_X1   g06421(.A1(new_n6610_), .A2(new_n3760_), .B1(new_n6608_), .B2(new_n6606_), .ZN(new_n6614_));
  AOI21_X1   g06422(.A1(new_n6614_), .A2(\asqrt[42] ), .B(new_n6437_), .ZN(new_n6615_));
  NOR2_X1    g06423(.A1(new_n6615_), .A2(new_n6613_), .ZN(new_n6616_));
  AOI22_X1   g06424(.A1(new_n6614_), .A2(\asqrt[42] ), .B1(new_n6612_), .B2(new_n6609_), .ZN(new_n6617_));
  INV_X1     g06425(.I(new_n6445_), .ZN(new_n6618_));
  OAI21_X1   g06426(.A1(new_n6617_), .A2(new_n3208_), .B(new_n6618_), .ZN(new_n6619_));
  NAND2_X1   g06427(.A1(new_n6619_), .A2(new_n6616_), .ZN(new_n6620_));
  OAI22_X1   g06428(.A1(new_n6617_), .A2(new_n3208_), .B1(new_n6615_), .B2(new_n6613_), .ZN(new_n6621_));
  AOI21_X1   g06429(.A1(new_n6621_), .A2(\asqrt[44] ), .B(new_n6452_), .ZN(new_n6622_));
  NOR2_X1    g06430(.A1(new_n6622_), .A2(new_n6620_), .ZN(new_n6623_));
  AOI22_X1   g06431(.A1(new_n6621_), .A2(\asqrt[44] ), .B1(new_n6619_), .B2(new_n6616_), .ZN(new_n6624_));
  INV_X1     g06432(.I(new_n6460_), .ZN(new_n6625_));
  OAI21_X1   g06433(.A1(new_n6624_), .A2(new_n2728_), .B(new_n6625_), .ZN(new_n6626_));
  NAND2_X1   g06434(.A1(new_n6626_), .A2(new_n6623_), .ZN(new_n6627_));
  OAI22_X1   g06435(.A1(new_n6624_), .A2(new_n2728_), .B1(new_n6622_), .B2(new_n6620_), .ZN(new_n6628_));
  AOI21_X1   g06436(.A1(new_n6628_), .A2(\asqrt[46] ), .B(new_n6467_), .ZN(new_n6629_));
  NOR2_X1    g06437(.A1(new_n6629_), .A2(new_n6627_), .ZN(new_n6630_));
  AOI22_X1   g06438(.A1(new_n6628_), .A2(\asqrt[46] ), .B1(new_n6626_), .B2(new_n6623_), .ZN(new_n6631_));
  INV_X1     g06439(.I(new_n6475_), .ZN(new_n6632_));
  OAI21_X1   g06440(.A1(new_n6631_), .A2(new_n2253_), .B(new_n6632_), .ZN(new_n6633_));
  NAND2_X1   g06441(.A1(new_n6633_), .A2(new_n6630_), .ZN(new_n6634_));
  OAI22_X1   g06442(.A1(new_n6631_), .A2(new_n2253_), .B1(new_n6629_), .B2(new_n6627_), .ZN(new_n6635_));
  AOI21_X1   g06443(.A1(new_n6635_), .A2(\asqrt[48] ), .B(new_n6482_), .ZN(new_n6636_));
  NOR2_X1    g06444(.A1(new_n6636_), .A2(new_n6634_), .ZN(new_n6637_));
  AOI22_X1   g06445(.A1(new_n6635_), .A2(\asqrt[48] ), .B1(new_n6633_), .B2(new_n6630_), .ZN(new_n6638_));
  INV_X1     g06446(.I(new_n6490_), .ZN(new_n6639_));
  OAI21_X1   g06447(.A1(new_n6638_), .A2(new_n1854_), .B(new_n6639_), .ZN(new_n6640_));
  NAND2_X1   g06448(.A1(new_n6640_), .A2(new_n6637_), .ZN(new_n6641_));
  OAI22_X1   g06449(.A1(new_n6638_), .A2(new_n1854_), .B1(new_n6636_), .B2(new_n6634_), .ZN(new_n6642_));
  AOI21_X1   g06450(.A1(new_n6642_), .A2(\asqrt[50] ), .B(new_n6497_), .ZN(new_n6643_));
  NOR2_X1    g06451(.A1(new_n6643_), .A2(new_n6641_), .ZN(new_n6644_));
  AOI22_X1   g06452(.A1(new_n6642_), .A2(\asqrt[50] ), .B1(new_n6640_), .B2(new_n6637_), .ZN(new_n6645_));
  INV_X1     g06453(.I(new_n6505_), .ZN(new_n6646_));
  OAI21_X1   g06454(.A1(new_n6645_), .A2(new_n1436_), .B(new_n6646_), .ZN(new_n6647_));
  NAND2_X1   g06455(.A1(new_n6647_), .A2(new_n6644_), .ZN(new_n6648_));
  OAI22_X1   g06456(.A1(new_n6645_), .A2(new_n1436_), .B1(new_n6643_), .B2(new_n6641_), .ZN(new_n6649_));
  AOI21_X1   g06457(.A1(new_n6649_), .A2(\asqrt[52] ), .B(new_n6512_), .ZN(new_n6650_));
  NOR2_X1    g06458(.A1(new_n6650_), .A2(new_n6648_), .ZN(new_n6651_));
  AOI22_X1   g06459(.A1(new_n6649_), .A2(\asqrt[52] ), .B1(new_n6647_), .B2(new_n6644_), .ZN(new_n6652_));
  INV_X1     g06460(.I(new_n6519_), .ZN(new_n6653_));
  OAI21_X1   g06461(.A1(new_n6652_), .A2(new_n1096_), .B(new_n6653_), .ZN(new_n6654_));
  NAND2_X1   g06462(.A1(new_n6654_), .A2(new_n6651_), .ZN(new_n6655_));
  OAI22_X1   g06463(.A1(new_n6652_), .A2(new_n1096_), .B1(new_n6650_), .B2(new_n6648_), .ZN(new_n6656_));
  AOI21_X1   g06464(.A1(new_n6656_), .A2(\asqrt[54] ), .B(new_n6525_), .ZN(new_n6657_));
  NOR2_X1    g06465(.A1(new_n6657_), .A2(new_n6655_), .ZN(new_n6658_));
  AOI22_X1   g06466(.A1(new_n6656_), .A2(\asqrt[54] ), .B1(new_n6654_), .B2(new_n6651_), .ZN(new_n6659_));
  INV_X1     g06467(.I(new_n6532_), .ZN(new_n6660_));
  OAI21_X1   g06468(.A1(new_n6659_), .A2(new_n825_), .B(new_n6660_), .ZN(new_n6661_));
  NAND2_X1   g06469(.A1(new_n6661_), .A2(new_n6658_), .ZN(new_n6662_));
  OAI22_X1   g06470(.A1(new_n6659_), .A2(new_n825_), .B1(new_n6657_), .B2(new_n6655_), .ZN(new_n6663_));
  AOI21_X1   g06471(.A1(new_n6663_), .A2(\asqrt[56] ), .B(new_n6538_), .ZN(new_n6664_));
  NOR2_X1    g06472(.A1(new_n6664_), .A2(new_n6662_), .ZN(new_n6665_));
  AOI22_X1   g06473(.A1(new_n6663_), .A2(\asqrt[56] ), .B1(new_n6661_), .B2(new_n6658_), .ZN(new_n6666_));
  INV_X1     g06474(.I(new_n6545_), .ZN(new_n6667_));
  OAI21_X1   g06475(.A1(new_n6666_), .A2(new_n587_), .B(new_n6667_), .ZN(new_n6668_));
  NAND2_X1   g06476(.A1(new_n6668_), .A2(new_n6665_), .ZN(new_n6669_));
  OAI22_X1   g06477(.A1(new_n6666_), .A2(new_n587_), .B1(new_n6664_), .B2(new_n6662_), .ZN(new_n6670_));
  AOI21_X1   g06478(.A1(new_n6670_), .A2(\asqrt[58] ), .B(new_n6551_), .ZN(new_n6671_));
  NOR2_X1    g06479(.A1(new_n6671_), .A2(new_n6669_), .ZN(new_n6672_));
  AOI22_X1   g06480(.A1(new_n6670_), .A2(\asqrt[58] ), .B1(new_n6668_), .B2(new_n6665_), .ZN(new_n6673_));
  INV_X1     g06481(.I(new_n6558_), .ZN(new_n6674_));
  OAI21_X1   g06482(.A1(new_n6673_), .A2(new_n376_), .B(new_n6674_), .ZN(new_n6675_));
  NAND2_X1   g06483(.A1(new_n6675_), .A2(new_n6672_), .ZN(new_n6676_));
  OAI22_X1   g06484(.A1(new_n6673_), .A2(new_n376_), .B1(new_n6671_), .B2(new_n6669_), .ZN(new_n6677_));
  AOI21_X1   g06485(.A1(new_n6677_), .A2(\asqrt[60] ), .B(new_n6564_), .ZN(new_n6678_));
  AOI22_X1   g06486(.A1(new_n6677_), .A2(\asqrt[60] ), .B1(new_n6675_), .B2(new_n6672_), .ZN(new_n6679_));
  OAI22_X1   g06487(.A1(new_n6679_), .A2(new_n229_), .B1(new_n6678_), .B2(new_n6676_), .ZN(new_n6680_));
  NOR4_X1    g06488(.A1(new_n6680_), .A2(\asqrt[62] ), .A3(new_n6332_), .A4(new_n6336_), .ZN(new_n6681_));
  NAND2_X1   g06489(.A1(new_n6352_), .A2(new_n5953_), .ZN(new_n6682_));
  XOR2_X1    g06490(.A1(new_n6352_), .A2(\asqrt[63] ), .Z(new_n6683_));
  AOI21_X1   g06491(.A1(\asqrt[33] ), .A2(new_n6682_), .B(new_n6683_), .ZN(new_n6684_));
  NAND2_X1   g06492(.A1(new_n6681_), .A2(new_n6684_), .ZN(new_n6685_));
  NOR4_X1    g06493(.A1(new_n6685_), .A2(new_n6313_), .A3(new_n6320_), .A4(new_n6577_), .ZN(new_n6686_));
  NOR2_X1    g06494(.A1(new_n6313_), .A2(\a[64] ), .ZN(new_n6687_));
  OAI21_X1   g06495(.A1(new_n6686_), .A2(new_n6687_), .B(new_n6312_), .ZN(new_n6688_));
  INV_X1     g06496(.I(new_n6312_), .ZN(new_n6689_));
  INV_X1     g06497(.I(new_n6320_), .ZN(new_n6690_));
  NOR2_X1    g06498(.A1(new_n6678_), .A2(new_n6676_), .ZN(new_n6691_));
  NOR3_X1    g06499(.A1(new_n6679_), .A2(new_n229_), .A3(new_n6570_), .ZN(new_n6692_));
  AOI21_X1   g06500(.A1(new_n6692_), .A2(new_n6691_), .B(new_n6337_), .ZN(new_n6693_));
  AOI21_X1   g06501(.A1(new_n6693_), .A2(new_n6575_), .B(new_n6332_), .ZN(new_n6694_));
  AOI22_X1   g06502(.A1(new_n6568_), .A2(\asqrt[61] ), .B1(new_n6566_), .B2(new_n6560_), .ZN(new_n6695_));
  NAND4_X1   g06503(.A1(new_n6695_), .A2(new_n196_), .A3(new_n6333_), .A4(new_n6569_), .ZN(new_n6696_));
  INV_X1     g06504(.I(new_n6684_), .ZN(new_n6697_));
  NOR2_X1    g06505(.A1(new_n6696_), .A2(new_n6697_), .ZN(new_n6698_));
  NAND4_X1   g06506(.A1(new_n6698_), .A2(new_n6694_), .A3(\a[65] ), .A4(new_n6690_), .ZN(new_n6699_));
  NAND3_X1   g06507(.A1(new_n6699_), .A2(\a[64] ), .A3(new_n6689_), .ZN(new_n6700_));
  NAND2_X1   g06508(.A1(new_n6688_), .A2(new_n6700_), .ZN(new_n6701_));
  NOR2_X1    g06509(.A1(new_n6685_), .A2(new_n6577_), .ZN(new_n6702_));
  NOR4_X1    g06510(.A1(new_n6318_), .A2(new_n5953_), .A3(new_n6367_), .A4(new_n6305_), .ZN(new_n6703_));
  NAND2_X1   g06511(.A1(\asqrt[33] ), .A2(\a[64] ), .ZN(new_n6704_));
  XOR2_X1    g06512(.A1(new_n6704_), .A2(new_n6703_), .Z(new_n6705_));
  NOR2_X1    g06513(.A1(new_n6705_), .A2(new_n6309_), .ZN(new_n6706_));
  INV_X1     g06514(.I(new_n6706_), .ZN(new_n6707_));
  NAND3_X1   g06515(.A1(new_n6698_), .A2(new_n6694_), .A3(new_n6690_), .ZN(new_n6708_));
  NAND2_X1   g06516(.A1(new_n6529_), .A2(\asqrt[55] ), .ZN(new_n6709_));
  AOI21_X1   g06517(.A1(new_n6709_), .A2(new_n6528_), .B(new_n724_), .ZN(new_n6710_));
  OAI21_X1   g06518(.A1(new_n6534_), .A2(new_n6710_), .B(\asqrt[57] ), .ZN(new_n6711_));
  AOI21_X1   g06519(.A1(new_n6541_), .A2(new_n6711_), .B(new_n504_), .ZN(new_n6712_));
  OAI21_X1   g06520(.A1(new_n6547_), .A2(new_n6712_), .B(\asqrt[59] ), .ZN(new_n6713_));
  AOI21_X1   g06521(.A1(new_n6554_), .A2(new_n6713_), .B(new_n275_), .ZN(new_n6714_));
  OAI21_X1   g06522(.A1(new_n6560_), .A2(new_n6714_), .B(\asqrt[61] ), .ZN(new_n6715_));
  NOR3_X1    g06523(.A1(new_n6567_), .A2(new_n6715_), .A3(new_n6570_), .ZN(new_n6716_));
  NOR3_X1    g06524(.A1(new_n6716_), .A2(new_n6337_), .A3(new_n6576_), .ZN(new_n6717_));
  OAI21_X1   g06525(.A1(new_n6717_), .A2(new_n6332_), .B(new_n6696_), .ZN(new_n6718_));
  NOR2_X1    g06526(.A1(new_n6690_), .A2(new_n6684_), .ZN(new_n6719_));
  NAND2_X1   g06527(.A1(new_n6719_), .A2(\asqrt[33] ), .ZN(new_n6720_));
  OAI21_X1   g06528(.A1(new_n6718_), .A2(new_n6720_), .B(new_n6339_), .ZN(new_n6721_));
  NAND3_X1   g06529(.A1(new_n6721_), .A2(new_n6340_), .A3(new_n6708_), .ZN(new_n6722_));
  NOR4_X1    g06530(.A1(new_n6577_), .A2(new_n6320_), .A3(new_n6696_), .A4(new_n6697_), .ZN(\asqrt[32] ));
  NAND2_X1   g06531(.A1(new_n6656_), .A2(\asqrt[54] ), .ZN(new_n6724_));
  AOI21_X1   g06532(.A1(new_n6724_), .A2(new_n6655_), .B(new_n825_), .ZN(new_n6725_));
  OAI21_X1   g06533(.A1(new_n6658_), .A2(new_n6725_), .B(\asqrt[56] ), .ZN(new_n6726_));
  AOI21_X1   g06534(.A1(new_n6662_), .A2(new_n6726_), .B(new_n587_), .ZN(new_n6727_));
  OAI21_X1   g06535(.A1(new_n6665_), .A2(new_n6727_), .B(\asqrt[58] ), .ZN(new_n6728_));
  AOI21_X1   g06536(.A1(new_n6669_), .A2(new_n6728_), .B(new_n376_), .ZN(new_n6729_));
  OAI21_X1   g06537(.A1(new_n6672_), .A2(new_n6729_), .B(\asqrt[60] ), .ZN(new_n6730_));
  AOI21_X1   g06538(.A1(new_n6676_), .A2(new_n6730_), .B(new_n229_), .ZN(new_n6731_));
  NAND4_X1   g06539(.A1(new_n6731_), .A2(new_n6560_), .A3(new_n6566_), .A4(new_n6571_), .ZN(new_n6732_));
  NAND3_X1   g06540(.A1(new_n6732_), .A2(new_n6338_), .A3(new_n6575_), .ZN(new_n6733_));
  AOI21_X1   g06541(.A1(new_n6333_), .A2(new_n6733_), .B(new_n6681_), .ZN(new_n6734_));
  INV_X1     g06542(.I(new_n6720_), .ZN(new_n6735_));
  AOI21_X1   g06543(.A1(new_n6734_), .A2(new_n6735_), .B(\a[66] ), .ZN(new_n6736_));
  OAI21_X1   g06544(.A1(new_n6736_), .A2(new_n6341_), .B(\asqrt[32] ), .ZN(new_n6737_));
  NAND4_X1   g06545(.A1(new_n6737_), .A2(new_n6722_), .A3(new_n5991_), .A4(new_n6707_), .ZN(new_n6738_));
  NAND2_X1   g06546(.A1(new_n6738_), .A2(new_n6701_), .ZN(new_n6739_));
  NAND3_X1   g06547(.A1(new_n6688_), .A2(new_n6700_), .A3(new_n6707_), .ZN(new_n6740_));
  AOI21_X1   g06548(.A1(\asqrt[33] ), .A2(new_n6339_), .B(\a[67] ), .ZN(new_n6741_));
  NOR2_X1    g06549(.A1(new_n6356_), .A2(\a[66] ), .ZN(new_n6742_));
  AOI21_X1   g06550(.A1(\asqrt[33] ), .A2(\a[66] ), .B(new_n6343_), .ZN(new_n6743_));
  OAI21_X1   g06551(.A1(new_n6742_), .A2(new_n6741_), .B(new_n6743_), .ZN(new_n6744_));
  INV_X1     g06552(.I(new_n6744_), .ZN(new_n6745_));
  NAND3_X1   g06553(.A1(\asqrt[32] ), .A2(new_n6364_), .A3(new_n6745_), .ZN(new_n6746_));
  OAI21_X1   g06554(.A1(new_n6708_), .A2(new_n6744_), .B(new_n6363_), .ZN(new_n6747_));
  NAND3_X1   g06555(.A1(new_n6747_), .A2(new_n6746_), .A3(new_n5626_), .ZN(new_n6748_));
  AOI21_X1   g06556(.A1(new_n6740_), .A2(\asqrt[34] ), .B(new_n6748_), .ZN(new_n6749_));
  NOR2_X1    g06557(.A1(new_n6739_), .A2(new_n6749_), .ZN(new_n6750_));
  NAND2_X1   g06558(.A1(new_n6740_), .A2(\asqrt[34] ), .ZN(new_n6751_));
  AOI21_X1   g06559(.A1(new_n6739_), .A2(new_n6751_), .B(new_n5626_), .ZN(new_n6752_));
  NAND2_X1   g06560(.A1(new_n6378_), .A2(\asqrt[35] ), .ZN(new_n6753_));
  NAND2_X1   g06561(.A1(new_n6372_), .A2(new_n6375_), .ZN(new_n6754_));
  NAND3_X1   g06562(.A1(new_n6754_), .A2(new_n6586_), .A3(new_n5626_), .ZN(new_n6755_));
  NOR2_X1    g06563(.A1(new_n6708_), .A2(new_n6755_), .ZN(new_n6756_));
  AND2_X2    g06564(.A1(new_n6756_), .A2(new_n6753_), .Z(new_n6757_));
  NOR2_X1    g06565(.A1(new_n6756_), .A2(new_n6753_), .ZN(new_n6758_));
  NOR3_X1    g06566(.A1(new_n6757_), .A2(\asqrt[36] ), .A3(new_n6758_), .ZN(new_n6759_));
  INV_X1     g06567(.I(new_n6759_), .ZN(new_n6760_));
  OAI21_X1   g06568(.A1(new_n6752_), .A2(new_n6760_), .B(new_n6750_), .ZN(new_n6761_));
  OAI21_X1   g06569(.A1(new_n6752_), .A2(new_n6750_), .B(\asqrt[36] ), .ZN(new_n6762_));
  NAND2_X1   g06570(.A1(new_n6592_), .A2(\asqrt[36] ), .ZN(new_n6763_));
  NOR2_X1    g06571(.A1(new_n6588_), .A2(new_n6587_), .ZN(new_n6764_));
  NOR4_X1    g06572(.A1(new_n6708_), .A2(\asqrt[36] ), .A3(new_n6764_), .A4(new_n6592_), .ZN(new_n6765_));
  XOR2_X1    g06573(.A1(new_n6765_), .A2(new_n6763_), .Z(new_n6766_));
  NAND2_X1   g06574(.A1(new_n6766_), .A2(new_n4973_), .ZN(new_n6767_));
  INV_X1     g06575(.I(new_n6767_), .ZN(new_n6768_));
  AOI21_X1   g06576(.A1(new_n6762_), .A2(new_n6768_), .B(new_n6761_), .ZN(new_n6769_));
  AOI21_X1   g06577(.A1(new_n6761_), .A2(new_n6762_), .B(new_n4973_), .ZN(new_n6770_));
  NAND2_X1   g06578(.A1(new_n6400_), .A2(\asqrt[37] ), .ZN(new_n6771_));
  NOR2_X1    g06579(.A1(new_n6395_), .A2(new_n6396_), .ZN(new_n6772_));
  NOR4_X1    g06580(.A1(new_n6708_), .A2(\asqrt[37] ), .A3(new_n6772_), .A4(new_n6400_), .ZN(new_n6773_));
  XOR2_X1    g06581(.A1(new_n6773_), .A2(new_n6771_), .Z(new_n6774_));
  NAND2_X1   g06582(.A1(new_n6774_), .A2(new_n4645_), .ZN(new_n6775_));
  OAI21_X1   g06583(.A1(new_n6770_), .A2(new_n6775_), .B(new_n6769_), .ZN(new_n6776_));
  OAI21_X1   g06584(.A1(new_n6769_), .A2(new_n6770_), .B(\asqrt[38] ), .ZN(new_n6777_));
  NOR4_X1    g06585(.A1(new_n6708_), .A2(\asqrt[38] ), .A3(new_n6403_), .A4(new_n6600_), .ZN(new_n6778_));
  AOI21_X1   g06586(.A1(new_n6771_), .A2(new_n6399_), .B(new_n4645_), .ZN(new_n6779_));
  NOR2_X1    g06587(.A1(new_n6778_), .A2(new_n6779_), .ZN(new_n6780_));
  NAND2_X1   g06588(.A1(new_n6780_), .A2(new_n4330_), .ZN(new_n6781_));
  INV_X1     g06589(.I(new_n6781_), .ZN(new_n6782_));
  AOI21_X1   g06590(.A1(new_n6777_), .A2(new_n6782_), .B(new_n6776_), .ZN(new_n6783_));
  AOI22_X1   g06591(.A1(new_n6738_), .A2(new_n6701_), .B1(\asqrt[34] ), .B2(new_n6740_), .ZN(new_n6784_));
  OAI21_X1   g06592(.A1(new_n6784_), .A2(new_n5626_), .B(new_n6759_), .ZN(new_n6785_));
  OAI22_X1   g06593(.A1(new_n6784_), .A2(new_n5626_), .B1(new_n6739_), .B2(new_n6749_), .ZN(new_n6786_));
  AOI22_X1   g06594(.A1(new_n6786_), .A2(\asqrt[36] ), .B1(new_n6785_), .B2(new_n6750_), .ZN(new_n6787_));
  INV_X1     g06595(.I(new_n6775_), .ZN(new_n6788_));
  OAI21_X1   g06596(.A1(new_n6787_), .A2(new_n4973_), .B(new_n6788_), .ZN(new_n6789_));
  AOI21_X1   g06597(.A1(new_n6786_), .A2(\asqrt[36] ), .B(new_n6767_), .ZN(new_n6790_));
  OAI22_X1   g06598(.A1(new_n6787_), .A2(new_n4973_), .B1(new_n6790_), .B2(new_n6761_), .ZN(new_n6791_));
  AOI22_X1   g06599(.A1(new_n6791_), .A2(\asqrt[38] ), .B1(new_n6789_), .B2(new_n6769_), .ZN(new_n6792_));
  NAND2_X1   g06600(.A1(new_n6414_), .A2(\asqrt[39] ), .ZN(new_n6793_));
  NOR4_X1    g06601(.A1(new_n6708_), .A2(\asqrt[39] ), .A3(new_n6409_), .A4(new_n6414_), .ZN(new_n6794_));
  XOR2_X1    g06602(.A1(new_n6794_), .A2(new_n6793_), .Z(new_n6795_));
  NAND2_X1   g06603(.A1(new_n6795_), .A2(new_n4018_), .ZN(new_n6796_));
  INV_X1     g06604(.I(new_n6796_), .ZN(new_n6797_));
  OAI21_X1   g06605(.A1(new_n6792_), .A2(new_n4330_), .B(new_n6797_), .ZN(new_n6798_));
  NAND2_X1   g06606(.A1(new_n6798_), .A2(new_n6783_), .ZN(new_n6799_));
  AOI21_X1   g06607(.A1(new_n6791_), .A2(\asqrt[38] ), .B(new_n6781_), .ZN(new_n6800_));
  OAI22_X1   g06608(.A1(new_n6792_), .A2(new_n4330_), .B1(new_n6800_), .B2(new_n6776_), .ZN(new_n6801_));
  NOR4_X1    g06609(.A1(new_n6708_), .A2(\asqrt[40] ), .A3(new_n6417_), .A4(new_n6607_), .ZN(new_n6802_));
  AOI21_X1   g06610(.A1(new_n6793_), .A2(new_n6413_), .B(new_n4018_), .ZN(new_n6803_));
  NOR2_X1    g06611(.A1(new_n6802_), .A2(new_n6803_), .ZN(new_n6804_));
  NAND2_X1   g06612(.A1(new_n6804_), .A2(new_n3760_), .ZN(new_n6805_));
  AOI21_X1   g06613(.A1(new_n6801_), .A2(\asqrt[40] ), .B(new_n6805_), .ZN(new_n6806_));
  NOR2_X1    g06614(.A1(new_n6806_), .A2(new_n6799_), .ZN(new_n6807_));
  AOI22_X1   g06615(.A1(new_n6801_), .A2(\asqrt[40] ), .B1(new_n6798_), .B2(new_n6783_), .ZN(new_n6808_));
  NAND2_X1   g06616(.A1(new_n6428_), .A2(\asqrt[41] ), .ZN(new_n6809_));
  NOR4_X1    g06617(.A1(new_n6708_), .A2(\asqrt[41] ), .A3(new_n6423_), .A4(new_n6428_), .ZN(new_n6810_));
  XOR2_X1    g06618(.A1(new_n6810_), .A2(new_n6809_), .Z(new_n6811_));
  NAND2_X1   g06619(.A1(new_n6811_), .A2(new_n3481_), .ZN(new_n6812_));
  INV_X1     g06620(.I(new_n6812_), .ZN(new_n6813_));
  OAI21_X1   g06621(.A1(new_n6808_), .A2(new_n3760_), .B(new_n6813_), .ZN(new_n6814_));
  NAND2_X1   g06622(.A1(new_n6814_), .A2(new_n6807_), .ZN(new_n6815_));
  OAI22_X1   g06623(.A1(new_n6808_), .A2(new_n3760_), .B1(new_n6806_), .B2(new_n6799_), .ZN(new_n6816_));
  NOR4_X1    g06624(.A1(new_n6708_), .A2(\asqrt[42] ), .A3(new_n6430_), .A4(new_n6614_), .ZN(new_n6817_));
  AOI21_X1   g06625(.A1(new_n6809_), .A2(new_n6427_), .B(new_n3481_), .ZN(new_n6818_));
  NOR2_X1    g06626(.A1(new_n6817_), .A2(new_n6818_), .ZN(new_n6819_));
  NAND2_X1   g06627(.A1(new_n6819_), .A2(new_n3208_), .ZN(new_n6820_));
  AOI21_X1   g06628(.A1(new_n6816_), .A2(\asqrt[42] ), .B(new_n6820_), .ZN(new_n6821_));
  NOR2_X1    g06629(.A1(new_n6821_), .A2(new_n6815_), .ZN(new_n6822_));
  AOI22_X1   g06630(.A1(new_n6816_), .A2(\asqrt[42] ), .B1(new_n6814_), .B2(new_n6807_), .ZN(new_n6823_));
  NAND2_X1   g06631(.A1(new_n6441_), .A2(\asqrt[43] ), .ZN(new_n6824_));
  NOR4_X1    g06632(.A1(new_n6708_), .A2(\asqrt[43] ), .A3(new_n6436_), .A4(new_n6441_), .ZN(new_n6825_));
  XOR2_X1    g06633(.A1(new_n6825_), .A2(new_n6824_), .Z(new_n6826_));
  NAND2_X1   g06634(.A1(new_n6826_), .A2(new_n2941_), .ZN(new_n6827_));
  INV_X1     g06635(.I(new_n6827_), .ZN(new_n6828_));
  OAI21_X1   g06636(.A1(new_n6823_), .A2(new_n3208_), .B(new_n6828_), .ZN(new_n6829_));
  NAND2_X1   g06637(.A1(new_n6829_), .A2(new_n6822_), .ZN(new_n6830_));
  OAI22_X1   g06638(.A1(new_n6823_), .A2(new_n3208_), .B1(new_n6821_), .B2(new_n6815_), .ZN(new_n6831_));
  NAND2_X1   g06639(.A1(new_n6621_), .A2(\asqrt[44] ), .ZN(new_n6832_));
  NOR4_X1    g06640(.A1(new_n6708_), .A2(\asqrt[44] ), .A3(new_n6444_), .A4(new_n6621_), .ZN(new_n6833_));
  XOR2_X1    g06641(.A1(new_n6833_), .A2(new_n6832_), .Z(new_n6834_));
  NAND2_X1   g06642(.A1(new_n6834_), .A2(new_n2728_), .ZN(new_n6835_));
  AOI21_X1   g06643(.A1(new_n6831_), .A2(\asqrt[44] ), .B(new_n6835_), .ZN(new_n6836_));
  NOR2_X1    g06644(.A1(new_n6836_), .A2(new_n6830_), .ZN(new_n6837_));
  AOI22_X1   g06645(.A1(new_n6831_), .A2(\asqrt[44] ), .B1(new_n6829_), .B2(new_n6822_), .ZN(new_n6838_));
  NOR4_X1    g06646(.A1(new_n6708_), .A2(\asqrt[45] ), .A3(new_n6451_), .A4(new_n6456_), .ZN(new_n6839_));
  AOI21_X1   g06647(.A1(new_n6832_), .A2(new_n6620_), .B(new_n2728_), .ZN(new_n6840_));
  NOR2_X1    g06648(.A1(new_n6839_), .A2(new_n6840_), .ZN(new_n6841_));
  NAND2_X1   g06649(.A1(new_n6841_), .A2(new_n2488_), .ZN(new_n6842_));
  INV_X1     g06650(.I(new_n6842_), .ZN(new_n6843_));
  OAI21_X1   g06651(.A1(new_n6838_), .A2(new_n2728_), .B(new_n6843_), .ZN(new_n6844_));
  NAND2_X1   g06652(.A1(new_n6844_), .A2(new_n6837_), .ZN(new_n6845_));
  OAI22_X1   g06653(.A1(new_n6838_), .A2(new_n2728_), .B1(new_n6836_), .B2(new_n6830_), .ZN(new_n6846_));
  NAND2_X1   g06654(.A1(new_n6628_), .A2(\asqrt[46] ), .ZN(new_n6847_));
  NOR4_X1    g06655(.A1(new_n6708_), .A2(\asqrt[46] ), .A3(new_n6459_), .A4(new_n6628_), .ZN(new_n6848_));
  XOR2_X1    g06656(.A1(new_n6848_), .A2(new_n6847_), .Z(new_n6849_));
  NAND2_X1   g06657(.A1(new_n6849_), .A2(new_n2253_), .ZN(new_n6850_));
  AOI21_X1   g06658(.A1(new_n6846_), .A2(\asqrt[46] ), .B(new_n6850_), .ZN(new_n6851_));
  NOR2_X1    g06659(.A1(new_n6851_), .A2(new_n6845_), .ZN(new_n6852_));
  AOI22_X1   g06660(.A1(new_n6846_), .A2(\asqrt[46] ), .B1(new_n6844_), .B2(new_n6837_), .ZN(new_n6853_));
  NOR4_X1    g06661(.A1(new_n6708_), .A2(\asqrt[47] ), .A3(new_n6466_), .A4(new_n6471_), .ZN(new_n6854_));
  AOI21_X1   g06662(.A1(new_n6847_), .A2(new_n6627_), .B(new_n2253_), .ZN(new_n6855_));
  NOR2_X1    g06663(.A1(new_n6854_), .A2(new_n6855_), .ZN(new_n6856_));
  NAND2_X1   g06664(.A1(new_n6856_), .A2(new_n2046_), .ZN(new_n6857_));
  INV_X1     g06665(.I(new_n6857_), .ZN(new_n6858_));
  OAI21_X1   g06666(.A1(new_n6853_), .A2(new_n2253_), .B(new_n6858_), .ZN(new_n6859_));
  NAND2_X1   g06667(.A1(new_n6859_), .A2(new_n6852_), .ZN(new_n6860_));
  OAI22_X1   g06668(.A1(new_n6853_), .A2(new_n2253_), .B1(new_n6851_), .B2(new_n6845_), .ZN(new_n6861_));
  NAND2_X1   g06669(.A1(new_n6635_), .A2(\asqrt[48] ), .ZN(new_n6862_));
  NOR4_X1    g06670(.A1(new_n6708_), .A2(\asqrt[48] ), .A3(new_n6474_), .A4(new_n6635_), .ZN(new_n6863_));
  XOR2_X1    g06671(.A1(new_n6863_), .A2(new_n6862_), .Z(new_n6864_));
  NAND2_X1   g06672(.A1(new_n6864_), .A2(new_n1854_), .ZN(new_n6865_));
  AOI21_X1   g06673(.A1(new_n6861_), .A2(\asqrt[48] ), .B(new_n6865_), .ZN(new_n6866_));
  NOR2_X1    g06674(.A1(new_n6866_), .A2(new_n6860_), .ZN(new_n6867_));
  AOI22_X1   g06675(.A1(new_n6861_), .A2(\asqrt[48] ), .B1(new_n6859_), .B2(new_n6852_), .ZN(new_n6868_));
  NOR4_X1    g06676(.A1(new_n6708_), .A2(\asqrt[49] ), .A3(new_n6481_), .A4(new_n6486_), .ZN(new_n6869_));
  AOI21_X1   g06677(.A1(new_n6862_), .A2(new_n6634_), .B(new_n1854_), .ZN(new_n6870_));
  NOR2_X1    g06678(.A1(new_n6869_), .A2(new_n6870_), .ZN(new_n6871_));
  NAND2_X1   g06679(.A1(new_n6871_), .A2(new_n1595_), .ZN(new_n6872_));
  INV_X1     g06680(.I(new_n6872_), .ZN(new_n6873_));
  OAI21_X1   g06681(.A1(new_n6868_), .A2(new_n1854_), .B(new_n6873_), .ZN(new_n6874_));
  NAND2_X1   g06682(.A1(new_n6874_), .A2(new_n6867_), .ZN(new_n6875_));
  OAI22_X1   g06683(.A1(new_n6868_), .A2(new_n1854_), .B1(new_n6866_), .B2(new_n6860_), .ZN(new_n6876_));
  NAND2_X1   g06684(.A1(new_n6642_), .A2(\asqrt[50] ), .ZN(new_n6877_));
  NOR4_X1    g06685(.A1(new_n6708_), .A2(\asqrt[50] ), .A3(new_n6489_), .A4(new_n6642_), .ZN(new_n6878_));
  XOR2_X1    g06686(.A1(new_n6878_), .A2(new_n6877_), .Z(new_n6879_));
  NAND2_X1   g06687(.A1(new_n6879_), .A2(new_n1436_), .ZN(new_n6880_));
  AOI21_X1   g06688(.A1(new_n6876_), .A2(\asqrt[50] ), .B(new_n6880_), .ZN(new_n6881_));
  NOR2_X1    g06689(.A1(new_n6881_), .A2(new_n6875_), .ZN(new_n6882_));
  AOI22_X1   g06690(.A1(new_n6876_), .A2(\asqrt[50] ), .B1(new_n6874_), .B2(new_n6867_), .ZN(new_n6883_));
  NOR4_X1    g06691(.A1(new_n6708_), .A2(\asqrt[51] ), .A3(new_n6496_), .A4(new_n6501_), .ZN(new_n6884_));
  AOI21_X1   g06692(.A1(new_n6877_), .A2(new_n6641_), .B(new_n1436_), .ZN(new_n6885_));
  NOR2_X1    g06693(.A1(new_n6884_), .A2(new_n6885_), .ZN(new_n6886_));
  NAND2_X1   g06694(.A1(new_n6886_), .A2(new_n1260_), .ZN(new_n6887_));
  INV_X1     g06695(.I(new_n6887_), .ZN(new_n6888_));
  OAI21_X1   g06696(.A1(new_n6883_), .A2(new_n1436_), .B(new_n6888_), .ZN(new_n6889_));
  NAND2_X1   g06697(.A1(new_n6889_), .A2(new_n6882_), .ZN(new_n6890_));
  OAI22_X1   g06698(.A1(new_n6883_), .A2(new_n1436_), .B1(new_n6881_), .B2(new_n6875_), .ZN(new_n6891_));
  NAND2_X1   g06699(.A1(new_n6649_), .A2(\asqrt[52] ), .ZN(new_n6892_));
  NOR4_X1    g06700(.A1(new_n6708_), .A2(\asqrt[52] ), .A3(new_n6504_), .A4(new_n6649_), .ZN(new_n6893_));
  XOR2_X1    g06701(.A1(new_n6893_), .A2(new_n6892_), .Z(new_n6894_));
  NAND2_X1   g06702(.A1(new_n6894_), .A2(new_n1096_), .ZN(new_n6895_));
  AOI21_X1   g06703(.A1(new_n6891_), .A2(\asqrt[52] ), .B(new_n6895_), .ZN(new_n6896_));
  NOR2_X1    g06704(.A1(new_n6896_), .A2(new_n6890_), .ZN(new_n6897_));
  AOI22_X1   g06705(.A1(new_n6891_), .A2(\asqrt[52] ), .B1(new_n6889_), .B2(new_n6882_), .ZN(new_n6898_));
  NOR2_X1    g06706(.A1(new_n6652_), .A2(new_n1096_), .ZN(new_n6899_));
  NOR4_X1    g06707(.A1(new_n6708_), .A2(\asqrt[53] ), .A3(new_n6511_), .A4(new_n6516_), .ZN(new_n6900_));
  XNOR2_X1   g06708(.A1(new_n6900_), .A2(new_n6899_), .ZN(new_n6901_));
  NAND2_X1   g06709(.A1(new_n6901_), .A2(new_n970_), .ZN(new_n6902_));
  INV_X1     g06710(.I(new_n6902_), .ZN(new_n6903_));
  OAI21_X1   g06711(.A1(new_n6898_), .A2(new_n1096_), .B(new_n6903_), .ZN(new_n6904_));
  NAND2_X1   g06712(.A1(new_n6904_), .A2(new_n6897_), .ZN(new_n6905_));
  OAI22_X1   g06713(.A1(new_n6898_), .A2(new_n1096_), .B1(new_n6896_), .B2(new_n6890_), .ZN(new_n6906_));
  NOR4_X1    g06714(.A1(new_n6708_), .A2(\asqrt[54] ), .A3(new_n6518_), .A4(new_n6656_), .ZN(new_n6907_));
  XOR2_X1    g06715(.A1(new_n6907_), .A2(new_n6724_), .Z(new_n6908_));
  NAND2_X1   g06716(.A1(new_n6908_), .A2(new_n825_), .ZN(new_n6909_));
  AOI21_X1   g06717(.A1(new_n6906_), .A2(\asqrt[54] ), .B(new_n6909_), .ZN(new_n6910_));
  NOR2_X1    g06718(.A1(new_n6910_), .A2(new_n6905_), .ZN(new_n6911_));
  AOI22_X1   g06719(.A1(new_n6906_), .A2(\asqrt[54] ), .B1(new_n6904_), .B2(new_n6897_), .ZN(new_n6912_));
  NOR4_X1    g06720(.A1(new_n6708_), .A2(\asqrt[55] ), .A3(new_n6524_), .A4(new_n6529_), .ZN(new_n6913_));
  XOR2_X1    g06721(.A1(new_n6913_), .A2(new_n6709_), .Z(new_n6914_));
  NAND2_X1   g06722(.A1(new_n6914_), .A2(new_n724_), .ZN(new_n6915_));
  INV_X1     g06723(.I(new_n6915_), .ZN(new_n6916_));
  OAI21_X1   g06724(.A1(new_n6912_), .A2(new_n825_), .B(new_n6916_), .ZN(new_n6917_));
  NAND2_X1   g06725(.A1(new_n6917_), .A2(new_n6911_), .ZN(new_n6918_));
  OAI22_X1   g06726(.A1(new_n6912_), .A2(new_n825_), .B1(new_n6910_), .B2(new_n6905_), .ZN(new_n6919_));
  NOR4_X1    g06727(.A1(new_n6708_), .A2(\asqrt[56] ), .A3(new_n6531_), .A4(new_n6663_), .ZN(new_n6920_));
  XOR2_X1    g06728(.A1(new_n6920_), .A2(new_n6726_), .Z(new_n6921_));
  NAND2_X1   g06729(.A1(new_n6921_), .A2(new_n587_), .ZN(new_n6922_));
  AOI21_X1   g06730(.A1(new_n6919_), .A2(\asqrt[56] ), .B(new_n6922_), .ZN(new_n6923_));
  NOR2_X1    g06731(.A1(new_n6923_), .A2(new_n6918_), .ZN(new_n6924_));
  AOI22_X1   g06732(.A1(new_n6919_), .A2(\asqrt[56] ), .B1(new_n6917_), .B2(new_n6911_), .ZN(new_n6925_));
  NOR4_X1    g06733(.A1(new_n6708_), .A2(\asqrt[57] ), .A3(new_n6537_), .A4(new_n6542_), .ZN(new_n6926_));
  XOR2_X1    g06734(.A1(new_n6926_), .A2(new_n6711_), .Z(new_n6927_));
  NAND2_X1   g06735(.A1(new_n6927_), .A2(new_n504_), .ZN(new_n6928_));
  INV_X1     g06736(.I(new_n6928_), .ZN(new_n6929_));
  OAI21_X1   g06737(.A1(new_n6925_), .A2(new_n587_), .B(new_n6929_), .ZN(new_n6930_));
  NAND2_X1   g06738(.A1(new_n6930_), .A2(new_n6924_), .ZN(new_n6931_));
  OAI22_X1   g06739(.A1(new_n6925_), .A2(new_n587_), .B1(new_n6923_), .B2(new_n6918_), .ZN(new_n6932_));
  NOR4_X1    g06740(.A1(new_n6708_), .A2(\asqrt[58] ), .A3(new_n6544_), .A4(new_n6670_), .ZN(new_n6933_));
  XOR2_X1    g06741(.A1(new_n6933_), .A2(new_n6728_), .Z(new_n6934_));
  NAND2_X1   g06742(.A1(new_n6934_), .A2(new_n376_), .ZN(new_n6935_));
  AOI21_X1   g06743(.A1(new_n6932_), .A2(\asqrt[58] ), .B(new_n6935_), .ZN(new_n6936_));
  NOR2_X1    g06744(.A1(new_n6936_), .A2(new_n6931_), .ZN(new_n6937_));
  AOI22_X1   g06745(.A1(new_n6932_), .A2(\asqrt[58] ), .B1(new_n6930_), .B2(new_n6924_), .ZN(new_n6938_));
  NOR4_X1    g06746(.A1(new_n6708_), .A2(\asqrt[59] ), .A3(new_n6550_), .A4(new_n6555_), .ZN(new_n6939_));
  XOR2_X1    g06747(.A1(new_n6939_), .A2(new_n6713_), .Z(new_n6940_));
  AND2_X2    g06748(.A1(new_n6940_), .A2(new_n275_), .Z(new_n6941_));
  OAI21_X1   g06749(.A1(new_n6938_), .A2(new_n376_), .B(new_n6941_), .ZN(new_n6942_));
  NAND2_X1   g06750(.A1(new_n6942_), .A2(new_n6937_), .ZN(new_n6943_));
  NAND2_X1   g06751(.A1(new_n6906_), .A2(\asqrt[54] ), .ZN(new_n6944_));
  AOI21_X1   g06752(.A1(new_n6944_), .A2(new_n6905_), .B(new_n825_), .ZN(new_n6945_));
  OAI21_X1   g06753(.A1(new_n6911_), .A2(new_n6945_), .B(\asqrt[56] ), .ZN(new_n6946_));
  AOI21_X1   g06754(.A1(new_n6918_), .A2(new_n6946_), .B(new_n587_), .ZN(new_n6947_));
  OAI21_X1   g06755(.A1(new_n6924_), .A2(new_n6947_), .B(\asqrt[58] ), .ZN(new_n6948_));
  AOI21_X1   g06756(.A1(new_n6931_), .A2(new_n6948_), .B(new_n376_), .ZN(new_n6949_));
  OAI21_X1   g06757(.A1(new_n6937_), .A2(new_n6949_), .B(\asqrt[60] ), .ZN(new_n6950_));
  AOI21_X1   g06758(.A1(new_n6943_), .A2(new_n6950_), .B(new_n229_), .ZN(new_n6951_));
  NOR2_X1    g06759(.A1(new_n6695_), .A2(new_n196_), .ZN(new_n6952_));
  NOR2_X1    g06760(.A1(new_n6680_), .A2(\asqrt[62] ), .ZN(new_n6953_));
  NAND3_X1   g06761(.A1(new_n6953_), .A2(new_n6952_), .A3(new_n6569_), .ZN(new_n6954_));
  NOR2_X1    g06762(.A1(new_n6708_), .A2(new_n6954_), .ZN(new_n6955_));
  OR3_X2     g06763(.A1(\asqrt[32] ), .A2(new_n6569_), .A3(new_n6953_), .Z(new_n6956_));
  AOI21_X1   g06764(.A1(new_n6956_), .A2(new_n6952_), .B(new_n6955_), .ZN(new_n6957_));
  NOR4_X1    g06765(.A1(new_n6708_), .A2(\asqrt[61] ), .A3(new_n6563_), .A4(new_n6568_), .ZN(new_n6958_));
  XOR2_X1    g06766(.A1(new_n6958_), .A2(new_n6715_), .Z(new_n6959_));
  NOR2_X1    g06767(.A1(new_n6959_), .A2(new_n196_), .ZN(new_n6960_));
  INV_X1     g06768(.I(new_n6960_), .ZN(new_n6961_));
  NOR2_X1    g06769(.A1(new_n6770_), .A2(new_n6775_), .ZN(new_n6962_));
  NOR3_X1    g06770(.A1(new_n6962_), .A2(new_n6761_), .A3(new_n6790_), .ZN(new_n6963_));
  NAND2_X1   g06771(.A1(new_n6777_), .A2(new_n6782_), .ZN(new_n6964_));
  NAND2_X1   g06772(.A1(new_n6964_), .A2(new_n6963_), .ZN(new_n6965_));
  NAND2_X1   g06773(.A1(new_n6776_), .A2(new_n6777_), .ZN(new_n6966_));
  AOI21_X1   g06774(.A1(new_n6966_), .A2(\asqrt[39] ), .B(new_n6796_), .ZN(new_n6967_));
  NOR2_X1    g06775(.A1(new_n6967_), .A2(new_n6965_), .ZN(new_n6968_));
  AOI21_X1   g06776(.A1(new_n6776_), .A2(new_n6777_), .B(new_n4330_), .ZN(new_n6969_));
  OAI21_X1   g06777(.A1(new_n6783_), .A2(new_n6969_), .B(\asqrt[40] ), .ZN(new_n6970_));
  INV_X1     g06778(.I(new_n6805_), .ZN(new_n6971_));
  NAND2_X1   g06779(.A1(new_n6970_), .A2(new_n6971_), .ZN(new_n6972_));
  NAND2_X1   g06780(.A1(new_n6972_), .A2(new_n6968_), .ZN(new_n6973_));
  AOI22_X1   g06781(.A1(new_n6966_), .A2(\asqrt[39] ), .B1(new_n6964_), .B2(new_n6963_), .ZN(new_n6974_));
  OAI22_X1   g06782(.A1(new_n6974_), .A2(new_n4018_), .B1(new_n6967_), .B2(new_n6965_), .ZN(new_n6975_));
  AOI21_X1   g06783(.A1(new_n6975_), .A2(\asqrt[41] ), .B(new_n6812_), .ZN(new_n6976_));
  NOR2_X1    g06784(.A1(new_n6976_), .A2(new_n6973_), .ZN(new_n6977_));
  AOI22_X1   g06785(.A1(new_n6975_), .A2(\asqrt[41] ), .B1(new_n6972_), .B2(new_n6968_), .ZN(new_n6978_));
  INV_X1     g06786(.I(new_n6820_), .ZN(new_n6979_));
  OAI21_X1   g06787(.A1(new_n6978_), .A2(new_n3481_), .B(new_n6979_), .ZN(new_n6980_));
  NAND2_X1   g06788(.A1(new_n6980_), .A2(new_n6977_), .ZN(new_n6981_));
  OAI22_X1   g06789(.A1(new_n6978_), .A2(new_n3481_), .B1(new_n6976_), .B2(new_n6973_), .ZN(new_n6982_));
  AOI21_X1   g06790(.A1(new_n6982_), .A2(\asqrt[43] ), .B(new_n6827_), .ZN(new_n6983_));
  NOR2_X1    g06791(.A1(new_n6983_), .A2(new_n6981_), .ZN(new_n6984_));
  AOI22_X1   g06792(.A1(new_n6982_), .A2(\asqrt[43] ), .B1(new_n6980_), .B2(new_n6977_), .ZN(new_n6985_));
  INV_X1     g06793(.I(new_n6835_), .ZN(new_n6986_));
  OAI21_X1   g06794(.A1(new_n6985_), .A2(new_n2941_), .B(new_n6986_), .ZN(new_n6987_));
  NAND2_X1   g06795(.A1(new_n6987_), .A2(new_n6984_), .ZN(new_n6988_));
  OAI22_X1   g06796(.A1(new_n6985_), .A2(new_n2941_), .B1(new_n6983_), .B2(new_n6981_), .ZN(new_n6989_));
  AOI21_X1   g06797(.A1(new_n6989_), .A2(\asqrt[45] ), .B(new_n6842_), .ZN(new_n6990_));
  NOR2_X1    g06798(.A1(new_n6990_), .A2(new_n6988_), .ZN(new_n6991_));
  AOI22_X1   g06799(.A1(new_n6989_), .A2(\asqrt[45] ), .B1(new_n6987_), .B2(new_n6984_), .ZN(new_n6992_));
  INV_X1     g06800(.I(new_n6850_), .ZN(new_n6993_));
  OAI21_X1   g06801(.A1(new_n6992_), .A2(new_n2488_), .B(new_n6993_), .ZN(new_n6994_));
  NAND2_X1   g06802(.A1(new_n6994_), .A2(new_n6991_), .ZN(new_n6995_));
  OAI22_X1   g06803(.A1(new_n6992_), .A2(new_n2488_), .B1(new_n6990_), .B2(new_n6988_), .ZN(new_n6996_));
  AOI21_X1   g06804(.A1(new_n6996_), .A2(\asqrt[47] ), .B(new_n6857_), .ZN(new_n6997_));
  NOR2_X1    g06805(.A1(new_n6997_), .A2(new_n6995_), .ZN(new_n6998_));
  AOI22_X1   g06806(.A1(new_n6996_), .A2(\asqrt[47] ), .B1(new_n6994_), .B2(new_n6991_), .ZN(new_n6999_));
  INV_X1     g06807(.I(new_n6865_), .ZN(new_n7000_));
  OAI21_X1   g06808(.A1(new_n6999_), .A2(new_n2046_), .B(new_n7000_), .ZN(new_n7001_));
  NAND2_X1   g06809(.A1(new_n7001_), .A2(new_n6998_), .ZN(new_n7002_));
  OAI22_X1   g06810(.A1(new_n6999_), .A2(new_n2046_), .B1(new_n6997_), .B2(new_n6995_), .ZN(new_n7003_));
  AOI21_X1   g06811(.A1(new_n7003_), .A2(\asqrt[49] ), .B(new_n6872_), .ZN(new_n7004_));
  NOR2_X1    g06812(.A1(new_n7004_), .A2(new_n7002_), .ZN(new_n7005_));
  AOI22_X1   g06813(.A1(new_n7003_), .A2(\asqrt[49] ), .B1(new_n7001_), .B2(new_n6998_), .ZN(new_n7006_));
  INV_X1     g06814(.I(new_n6880_), .ZN(new_n7007_));
  OAI21_X1   g06815(.A1(new_n7006_), .A2(new_n1595_), .B(new_n7007_), .ZN(new_n7008_));
  NAND2_X1   g06816(.A1(new_n7008_), .A2(new_n7005_), .ZN(new_n7009_));
  OAI22_X1   g06817(.A1(new_n7006_), .A2(new_n1595_), .B1(new_n7004_), .B2(new_n7002_), .ZN(new_n7010_));
  AOI21_X1   g06818(.A1(new_n7010_), .A2(\asqrt[51] ), .B(new_n6887_), .ZN(new_n7011_));
  NOR2_X1    g06819(.A1(new_n7011_), .A2(new_n7009_), .ZN(new_n7012_));
  AOI22_X1   g06820(.A1(new_n7010_), .A2(\asqrt[51] ), .B1(new_n7008_), .B2(new_n7005_), .ZN(new_n7013_));
  INV_X1     g06821(.I(new_n6895_), .ZN(new_n7014_));
  OAI21_X1   g06822(.A1(new_n7013_), .A2(new_n1260_), .B(new_n7014_), .ZN(new_n7015_));
  NAND2_X1   g06823(.A1(new_n7015_), .A2(new_n7012_), .ZN(new_n7016_));
  OAI22_X1   g06824(.A1(new_n7013_), .A2(new_n1260_), .B1(new_n7011_), .B2(new_n7009_), .ZN(new_n7017_));
  AOI21_X1   g06825(.A1(new_n7017_), .A2(\asqrt[53] ), .B(new_n6902_), .ZN(new_n7018_));
  NOR2_X1    g06826(.A1(new_n7018_), .A2(new_n7016_), .ZN(new_n7019_));
  AOI22_X1   g06827(.A1(new_n7017_), .A2(\asqrt[53] ), .B1(new_n7015_), .B2(new_n7012_), .ZN(new_n7020_));
  INV_X1     g06828(.I(new_n6909_), .ZN(new_n7021_));
  OAI21_X1   g06829(.A1(new_n7020_), .A2(new_n970_), .B(new_n7021_), .ZN(new_n7022_));
  NAND2_X1   g06830(.A1(new_n7022_), .A2(new_n7019_), .ZN(new_n7023_));
  OAI22_X1   g06831(.A1(new_n7020_), .A2(new_n970_), .B1(new_n7018_), .B2(new_n7016_), .ZN(new_n7024_));
  AOI21_X1   g06832(.A1(new_n7024_), .A2(\asqrt[55] ), .B(new_n6915_), .ZN(new_n7025_));
  NOR2_X1    g06833(.A1(new_n7025_), .A2(new_n7023_), .ZN(new_n7026_));
  AOI22_X1   g06834(.A1(new_n7024_), .A2(\asqrt[55] ), .B1(new_n7022_), .B2(new_n7019_), .ZN(new_n7027_));
  INV_X1     g06835(.I(new_n6922_), .ZN(new_n7028_));
  OAI21_X1   g06836(.A1(new_n7027_), .A2(new_n724_), .B(new_n7028_), .ZN(new_n7029_));
  NAND2_X1   g06837(.A1(new_n7029_), .A2(new_n7026_), .ZN(new_n7030_));
  NAND2_X1   g06838(.A1(new_n7017_), .A2(\asqrt[53] ), .ZN(new_n7031_));
  AOI21_X1   g06839(.A1(new_n7031_), .A2(new_n7016_), .B(new_n970_), .ZN(new_n7032_));
  OAI21_X1   g06840(.A1(new_n7019_), .A2(new_n7032_), .B(\asqrt[55] ), .ZN(new_n7033_));
  AOI21_X1   g06841(.A1(new_n7023_), .A2(new_n7033_), .B(new_n724_), .ZN(new_n7034_));
  OAI21_X1   g06842(.A1(new_n7026_), .A2(new_n7034_), .B(\asqrt[57] ), .ZN(new_n7035_));
  AOI21_X1   g06843(.A1(new_n7035_), .A2(new_n6929_), .B(new_n7030_), .ZN(new_n7036_));
  OAI22_X1   g06844(.A1(new_n7027_), .A2(new_n724_), .B1(new_n7025_), .B2(new_n7023_), .ZN(new_n7037_));
  AOI22_X1   g06845(.A1(new_n7037_), .A2(\asqrt[57] ), .B1(new_n7029_), .B2(new_n7026_), .ZN(new_n7038_));
  INV_X1     g06846(.I(new_n6935_), .ZN(new_n7039_));
  OAI21_X1   g06847(.A1(new_n7038_), .A2(new_n504_), .B(new_n7039_), .ZN(new_n7040_));
  NAND2_X1   g06848(.A1(new_n7040_), .A2(new_n7036_), .ZN(new_n7041_));
  AOI21_X1   g06849(.A1(new_n7030_), .A2(new_n7035_), .B(new_n504_), .ZN(new_n7042_));
  OAI21_X1   g06850(.A1(new_n7036_), .A2(new_n7042_), .B(\asqrt[59] ), .ZN(new_n7043_));
  AOI21_X1   g06851(.A1(new_n7043_), .A2(new_n6941_), .B(new_n7041_), .ZN(new_n7044_));
  NAND2_X1   g06852(.A1(new_n6931_), .A2(new_n6948_), .ZN(new_n7045_));
  AOI22_X1   g06853(.A1(new_n7045_), .A2(\asqrt[59] ), .B1(new_n7040_), .B2(new_n7036_), .ZN(new_n7046_));
  NOR4_X1    g06854(.A1(new_n6708_), .A2(\asqrt[60] ), .A3(new_n6557_), .A4(new_n6677_), .ZN(new_n7047_));
  XOR2_X1    g06855(.A1(new_n7047_), .A2(new_n6730_), .Z(new_n7048_));
  NAND2_X1   g06856(.A1(new_n7048_), .A2(new_n229_), .ZN(new_n7049_));
  INV_X1     g06857(.I(new_n7049_), .ZN(new_n7050_));
  OAI21_X1   g06858(.A1(new_n7046_), .A2(new_n275_), .B(new_n7050_), .ZN(new_n7051_));
  NAND2_X1   g06859(.A1(new_n7051_), .A2(new_n7044_), .ZN(new_n7052_));
  INV_X1     g06860(.I(new_n6959_), .ZN(new_n7053_));
  NOR2_X1    g06861(.A1(new_n7053_), .A2(\asqrt[62] ), .ZN(new_n7054_));
  INV_X1     g06862(.I(new_n7054_), .ZN(new_n7055_));
  NAND2_X1   g06863(.A1(new_n6951_), .A2(new_n7055_), .ZN(new_n7056_));
  OAI21_X1   g06864(.A1(new_n7056_), .A2(new_n7052_), .B(new_n6961_), .ZN(new_n7057_));
  NAND2_X1   g06865(.A1(new_n6696_), .A2(new_n6332_), .ZN(new_n7058_));
  OAI21_X1   g06866(.A1(\asqrt[32] ), .A2(new_n7058_), .B(new_n6573_), .ZN(new_n7059_));
  NAND2_X1   g06867(.A1(new_n7059_), .A2(new_n231_), .ZN(new_n7060_));
  OAI21_X1   g06868(.A1(new_n7057_), .A2(new_n7060_), .B(new_n6957_), .ZN(new_n7061_));
  OAI21_X1   g06869(.A1(new_n6333_), .A2(new_n6573_), .B(\asqrt[32] ), .ZN(new_n7062_));
  XOR2_X1    g06870(.A1(new_n6573_), .A2(\asqrt[63] ), .Z(new_n7063_));
  NAND2_X1   g06871(.A1(new_n7062_), .A2(new_n7063_), .ZN(new_n7064_));
  INV_X1     g06872(.I(new_n7064_), .ZN(new_n7065_));
  INV_X1     g06873(.I(new_n6957_), .ZN(new_n7066_));
  OAI22_X1   g06874(.A1(new_n6938_), .A2(new_n376_), .B1(new_n6936_), .B2(new_n6931_), .ZN(new_n7067_));
  AOI21_X1   g06875(.A1(new_n7067_), .A2(\asqrt[60] ), .B(new_n7049_), .ZN(new_n7068_));
  AOI22_X1   g06876(.A1(new_n7067_), .A2(\asqrt[60] ), .B1(new_n6942_), .B2(new_n6937_), .ZN(new_n7069_));
  OAI22_X1   g06877(.A1(new_n7069_), .A2(new_n229_), .B1(new_n7068_), .B2(new_n6943_), .ZN(new_n7070_));
  NOR4_X1    g06878(.A1(new_n7070_), .A2(\asqrt[62] ), .A3(new_n7066_), .A4(new_n6959_), .ZN(new_n7071_));
  NAND2_X1   g06879(.A1(new_n7071_), .A2(new_n7065_), .ZN(new_n7072_));
  NAND3_X1   g06880(.A1(new_n6702_), .A2(new_n6320_), .A3(new_n6333_), .ZN(new_n7073_));
  NOR3_X1    g06881(.A1(new_n7072_), .A2(new_n7061_), .A3(new_n7073_), .ZN(\asqrt[31] ));
  NAND2_X1   g06882(.A1(new_n6943_), .A2(new_n6950_), .ZN(new_n7075_));
  NOR3_X1    g06883(.A1(new_n7075_), .A2(\asqrt[61] ), .A3(new_n7048_), .ZN(new_n7076_));
  NAND2_X1   g06884(.A1(\asqrt[31] ), .A2(new_n7076_), .ZN(new_n7077_));
  XOR2_X1    g06885(.A1(new_n7077_), .A2(new_n6951_), .Z(new_n7078_));
  INV_X1     g06886(.I(new_n7078_), .ZN(new_n7079_));
  INV_X1     g06887(.I(\a[63] ), .ZN(new_n7080_));
  INV_X1     g06888(.I(\a[62] ), .ZN(new_n7081_));
  NOR2_X1    g06889(.A1(\a[60] ), .A2(\a[61] ), .ZN(new_n7082_));
  INV_X1     g06890(.I(new_n7082_), .ZN(new_n7083_));
  NOR4_X1    g06891(.A1(new_n6718_), .A2(new_n7081_), .A3(new_n6719_), .A4(new_n7083_), .ZN(new_n7084_));
  XOR2_X1    g06892(.A1(new_n7084_), .A2(new_n7080_), .Z(new_n7085_));
  NOR4_X1    g06893(.A1(new_n7072_), .A2(new_n7061_), .A3(new_n7080_), .A4(new_n7073_), .ZN(new_n7086_));
  NOR2_X1    g06894(.A1(new_n7080_), .A2(\a[62] ), .ZN(new_n7087_));
  OAI21_X1   g06895(.A1(new_n7086_), .A2(new_n7087_), .B(new_n7085_), .ZN(new_n7088_));
  INV_X1     g06896(.I(new_n7085_), .ZN(new_n7089_));
  NOR2_X1    g06897(.A1(new_n7068_), .A2(new_n6943_), .ZN(new_n7090_));
  NOR3_X1    g06898(.A1(new_n7069_), .A2(new_n229_), .A3(new_n7054_), .ZN(new_n7091_));
  AOI21_X1   g06899(.A1(new_n7091_), .A2(new_n7090_), .B(new_n6960_), .ZN(new_n7092_));
  INV_X1     g06900(.I(new_n7060_), .ZN(new_n7093_));
  AOI21_X1   g06901(.A1(new_n7092_), .A2(new_n7093_), .B(new_n7066_), .ZN(new_n7094_));
  AOI21_X1   g06902(.A1(new_n7070_), .A2(\asqrt[62] ), .B(new_n6957_), .ZN(new_n7095_));
  AOI21_X1   g06903(.A1(new_n7041_), .A2(new_n7043_), .B(new_n275_), .ZN(new_n7096_));
  OAI21_X1   g06904(.A1(new_n7044_), .A2(new_n7096_), .B(\asqrt[61] ), .ZN(new_n7097_));
  NAND4_X1   g06905(.A1(new_n7052_), .A2(new_n196_), .A3(new_n7097_), .A4(new_n7053_), .ZN(new_n7098_));
  NOR3_X1    g06906(.A1(new_n7095_), .A2(new_n7064_), .A3(new_n7098_), .ZN(new_n7099_));
  INV_X1     g06907(.I(new_n7073_), .ZN(new_n7100_));
  NAND4_X1   g06908(.A1(new_n7099_), .A2(\a[63] ), .A3(new_n7094_), .A4(new_n7100_), .ZN(new_n7101_));
  NAND3_X1   g06909(.A1(new_n7101_), .A2(\a[62] ), .A3(new_n7089_), .ZN(new_n7102_));
  NAND2_X1   g06910(.A1(new_n7088_), .A2(new_n7102_), .ZN(new_n7103_));
  NOR2_X1    g06911(.A1(new_n7072_), .A2(new_n7061_), .ZN(new_n7104_));
  NOR4_X1    g06912(.A1(new_n6685_), .A2(new_n6320_), .A3(new_n6332_), .A4(new_n6717_), .ZN(new_n7105_));
  NAND2_X1   g06913(.A1(\asqrt[32] ), .A2(\a[62] ), .ZN(new_n7106_));
  XOR2_X1    g06914(.A1(new_n7106_), .A2(new_n7105_), .Z(new_n7107_));
  NOR2_X1    g06915(.A1(new_n7107_), .A2(new_n7083_), .ZN(new_n7108_));
  INV_X1     g06916(.I(new_n7108_), .ZN(new_n7109_));
  NAND3_X1   g06917(.A1(new_n7099_), .A2(new_n7094_), .A3(new_n7100_), .ZN(new_n7110_));
  NOR4_X1    g06918(.A1(new_n7097_), .A2(new_n6943_), .A3(new_n7068_), .A4(new_n7054_), .ZN(new_n7111_));
  NOR3_X1    g06919(.A1(new_n7111_), .A2(new_n6960_), .A3(new_n7060_), .ZN(new_n7112_));
  AOI22_X1   g06920(.A1(new_n7075_), .A2(\asqrt[61] ), .B1(new_n7051_), .B2(new_n7044_), .ZN(new_n7113_));
  NAND4_X1   g06921(.A1(new_n7113_), .A2(new_n196_), .A3(new_n6957_), .A4(new_n7053_), .ZN(new_n7114_));
  OAI21_X1   g06922(.A1(new_n7112_), .A2(new_n7066_), .B(new_n7114_), .ZN(new_n7115_));
  NOR2_X1    g06923(.A1(new_n7065_), .A2(new_n7100_), .ZN(new_n7116_));
  NAND2_X1   g06924(.A1(new_n7116_), .A2(\asqrt[32] ), .ZN(new_n7117_));
  OAI21_X1   g06925(.A1(new_n7115_), .A2(new_n7117_), .B(new_n6300_), .ZN(new_n7118_));
  NAND3_X1   g06926(.A1(new_n7118_), .A2(new_n6308_), .A3(new_n7110_), .ZN(new_n7119_));
  NAND4_X1   g06927(.A1(new_n6951_), .A2(new_n7044_), .A3(new_n7051_), .A4(new_n7055_), .ZN(new_n7120_));
  NAND3_X1   g06928(.A1(new_n7120_), .A2(new_n6961_), .A3(new_n7093_), .ZN(new_n7121_));
  AOI21_X1   g06929(.A1(new_n6957_), .A2(new_n7121_), .B(new_n7071_), .ZN(new_n7122_));
  INV_X1     g06930(.I(new_n7117_), .ZN(new_n7123_));
  AOI21_X1   g06931(.A1(new_n7122_), .A2(new_n7123_), .B(\a[64] ), .ZN(new_n7124_));
  OAI21_X1   g06932(.A1(new_n7124_), .A2(new_n6309_), .B(\asqrt[31] ), .ZN(new_n7125_));
  NAND4_X1   g06933(.A1(new_n7119_), .A2(new_n7125_), .A3(new_n6365_), .A4(new_n7109_), .ZN(new_n7126_));
  NAND2_X1   g06934(.A1(new_n7126_), .A2(new_n7103_), .ZN(new_n7127_));
  NAND3_X1   g06935(.A1(new_n7088_), .A2(new_n7102_), .A3(new_n7109_), .ZN(new_n7128_));
  NOR2_X1    g06936(.A1(new_n6708_), .A2(\a[64] ), .ZN(new_n7129_));
  OAI22_X1   g06937(.A1(new_n7129_), .A2(\a[65] ), .B1(\a[64] ), .B2(new_n6699_), .ZN(new_n7130_));
  AOI21_X1   g06938(.A1(\asqrt[32] ), .A2(\a[64] ), .B(new_n6311_), .ZN(new_n7131_));
  AND2_X2    g06939(.A1(new_n7130_), .A2(new_n7131_), .Z(new_n7132_));
  NAND3_X1   g06940(.A1(\asqrt[31] ), .A2(new_n6707_), .A3(new_n7132_), .ZN(new_n7133_));
  INV_X1     g06941(.I(new_n7132_), .ZN(new_n7134_));
  OAI21_X1   g06942(.A1(new_n7110_), .A2(new_n7134_), .B(new_n6706_), .ZN(new_n7135_));
  NAND3_X1   g06943(.A1(new_n7133_), .A2(new_n7135_), .A3(new_n5991_), .ZN(new_n7136_));
  AOI21_X1   g06944(.A1(new_n7128_), .A2(\asqrt[33] ), .B(new_n7136_), .ZN(new_n7137_));
  NOR2_X1    g06945(.A1(new_n7127_), .A2(new_n7137_), .ZN(new_n7138_));
  AOI22_X1   g06946(.A1(new_n7126_), .A2(new_n7103_), .B1(\asqrt[33] ), .B2(new_n7128_), .ZN(new_n7139_));
  INV_X1     g06947(.I(new_n6687_), .ZN(new_n7140_));
  AOI21_X1   g06948(.A1(new_n6699_), .A2(new_n7140_), .B(new_n6689_), .ZN(new_n7141_));
  INV_X1     g06949(.I(new_n6700_), .ZN(new_n7142_));
  NOR3_X1    g06950(.A1(new_n7142_), .A2(new_n7141_), .A3(new_n6706_), .ZN(new_n7143_));
  AOI21_X1   g06951(.A1(new_n6737_), .A2(new_n6722_), .B(\asqrt[34] ), .ZN(new_n7144_));
  AND4_X2    g06952(.A1(new_n7143_), .A2(\asqrt[31] ), .A3(new_n6751_), .A4(new_n7144_), .Z(new_n7145_));
  NOR2_X1    g06953(.A1(new_n7143_), .A2(new_n5991_), .ZN(new_n7146_));
  NOR3_X1    g06954(.A1(new_n7145_), .A2(\asqrt[35] ), .A3(new_n7146_), .ZN(new_n7147_));
  OAI21_X1   g06955(.A1(new_n7139_), .A2(new_n5991_), .B(new_n7147_), .ZN(new_n7148_));
  NAND2_X1   g06956(.A1(new_n7148_), .A2(new_n7138_), .ZN(new_n7149_));
  OAI22_X1   g06957(.A1(new_n7139_), .A2(new_n5991_), .B1(new_n7127_), .B2(new_n7137_), .ZN(new_n7150_));
  NAND2_X1   g06958(.A1(new_n6747_), .A2(new_n6746_), .ZN(new_n7151_));
  NAND4_X1   g06959(.A1(\asqrt[31] ), .A2(new_n5626_), .A3(new_n7151_), .A4(new_n6784_), .ZN(new_n7152_));
  XOR2_X1    g06960(.A1(new_n7152_), .A2(new_n6752_), .Z(new_n7153_));
  NAND2_X1   g06961(.A1(new_n7153_), .A2(new_n5273_), .ZN(new_n7154_));
  AOI21_X1   g06962(.A1(new_n7150_), .A2(\asqrt[35] ), .B(new_n7154_), .ZN(new_n7155_));
  NOR2_X1    g06963(.A1(new_n7155_), .A2(new_n7149_), .ZN(new_n7156_));
  AOI22_X1   g06964(.A1(new_n7150_), .A2(\asqrt[35] ), .B1(new_n7148_), .B2(new_n7138_), .ZN(new_n7157_));
  NOR2_X1    g06965(.A1(new_n6757_), .A2(new_n6758_), .ZN(new_n7158_));
  NOR4_X1    g06966(.A1(new_n7110_), .A2(\asqrt[36] ), .A3(new_n7158_), .A4(new_n6786_), .ZN(new_n7159_));
  XOR2_X1    g06967(.A1(new_n7159_), .A2(new_n6762_), .Z(new_n7160_));
  NAND2_X1   g06968(.A1(new_n7160_), .A2(new_n4973_), .ZN(new_n7161_));
  INV_X1     g06969(.I(new_n7161_), .ZN(new_n7162_));
  OAI21_X1   g06970(.A1(new_n7157_), .A2(new_n5273_), .B(new_n7162_), .ZN(new_n7163_));
  NAND2_X1   g06971(.A1(new_n7163_), .A2(new_n7156_), .ZN(new_n7164_));
  OAI22_X1   g06972(.A1(new_n7157_), .A2(new_n5273_), .B1(new_n7155_), .B2(new_n7149_), .ZN(new_n7165_));
  NOR2_X1    g06973(.A1(new_n6766_), .A2(\asqrt[37] ), .ZN(new_n7166_));
  NAND3_X1   g06974(.A1(\asqrt[31] ), .A2(new_n6787_), .A3(new_n7166_), .ZN(new_n7167_));
  XOR2_X1    g06975(.A1(new_n7167_), .A2(new_n6770_), .Z(new_n7168_));
  NAND2_X1   g06976(.A1(new_n7168_), .A2(new_n4645_), .ZN(new_n7169_));
  AOI21_X1   g06977(.A1(new_n7165_), .A2(\asqrt[37] ), .B(new_n7169_), .ZN(new_n7170_));
  NOR2_X1    g06978(.A1(new_n7170_), .A2(new_n7164_), .ZN(new_n7171_));
  AOI22_X1   g06979(.A1(new_n7165_), .A2(\asqrt[37] ), .B1(new_n7163_), .B2(new_n7156_), .ZN(new_n7172_));
  NOR4_X1    g06980(.A1(new_n7110_), .A2(\asqrt[38] ), .A3(new_n6774_), .A4(new_n6791_), .ZN(new_n7173_));
  XOR2_X1    g06981(.A1(new_n7173_), .A2(new_n6777_), .Z(new_n7174_));
  NAND2_X1   g06982(.A1(new_n7174_), .A2(new_n4330_), .ZN(new_n7175_));
  INV_X1     g06983(.I(new_n7175_), .ZN(new_n7176_));
  OAI21_X1   g06984(.A1(new_n7172_), .A2(new_n4645_), .B(new_n7176_), .ZN(new_n7177_));
  NAND2_X1   g06985(.A1(new_n7177_), .A2(new_n7171_), .ZN(new_n7178_));
  OAI22_X1   g06986(.A1(new_n7172_), .A2(new_n4645_), .B1(new_n7170_), .B2(new_n7164_), .ZN(new_n7179_));
  NOR4_X1    g06987(.A1(new_n7110_), .A2(\asqrt[39] ), .A3(new_n6780_), .A4(new_n6966_), .ZN(new_n7180_));
  XNOR2_X1   g06988(.A1(new_n7180_), .A2(new_n6969_), .ZN(new_n7181_));
  NAND2_X1   g06989(.A1(new_n7181_), .A2(new_n4018_), .ZN(new_n7182_));
  AOI21_X1   g06990(.A1(new_n7179_), .A2(\asqrt[39] ), .B(new_n7182_), .ZN(new_n7183_));
  NOR2_X1    g06991(.A1(new_n7183_), .A2(new_n7178_), .ZN(new_n7184_));
  AOI22_X1   g06992(.A1(new_n7179_), .A2(\asqrt[39] ), .B1(new_n7177_), .B2(new_n7171_), .ZN(new_n7185_));
  NOR4_X1    g06993(.A1(new_n7110_), .A2(\asqrt[40] ), .A3(new_n6795_), .A4(new_n6801_), .ZN(new_n7186_));
  XOR2_X1    g06994(.A1(new_n7186_), .A2(new_n6970_), .Z(new_n7187_));
  NAND2_X1   g06995(.A1(new_n7187_), .A2(new_n3760_), .ZN(new_n7188_));
  INV_X1     g06996(.I(new_n7188_), .ZN(new_n7189_));
  OAI21_X1   g06997(.A1(new_n7185_), .A2(new_n4018_), .B(new_n7189_), .ZN(new_n7190_));
  NAND2_X1   g06998(.A1(new_n7190_), .A2(new_n7184_), .ZN(new_n7191_));
  OAI22_X1   g06999(.A1(new_n7185_), .A2(new_n4018_), .B1(new_n7183_), .B2(new_n7178_), .ZN(new_n7192_));
  NAND2_X1   g07000(.A1(new_n6975_), .A2(\asqrt[41] ), .ZN(new_n7193_));
  NOR4_X1    g07001(.A1(new_n7110_), .A2(\asqrt[41] ), .A3(new_n6804_), .A4(new_n6975_), .ZN(new_n7194_));
  XOR2_X1    g07002(.A1(new_n7194_), .A2(new_n7193_), .Z(new_n7195_));
  NAND2_X1   g07003(.A1(new_n7195_), .A2(new_n3481_), .ZN(new_n7196_));
  AOI21_X1   g07004(.A1(new_n7192_), .A2(\asqrt[41] ), .B(new_n7196_), .ZN(new_n7197_));
  NOR2_X1    g07005(.A1(new_n7197_), .A2(new_n7191_), .ZN(new_n7198_));
  AOI22_X1   g07006(.A1(new_n7192_), .A2(\asqrt[41] ), .B1(new_n7190_), .B2(new_n7184_), .ZN(new_n7199_));
  NOR4_X1    g07007(.A1(new_n7110_), .A2(\asqrt[42] ), .A3(new_n6811_), .A4(new_n6816_), .ZN(new_n7200_));
  AOI21_X1   g07008(.A1(new_n7193_), .A2(new_n6973_), .B(new_n3481_), .ZN(new_n7201_));
  NOR2_X1    g07009(.A1(new_n7200_), .A2(new_n7201_), .ZN(new_n7202_));
  NAND2_X1   g07010(.A1(new_n7202_), .A2(new_n3208_), .ZN(new_n7203_));
  INV_X1     g07011(.I(new_n7203_), .ZN(new_n7204_));
  OAI21_X1   g07012(.A1(new_n7199_), .A2(new_n3481_), .B(new_n7204_), .ZN(new_n7205_));
  NAND2_X1   g07013(.A1(new_n7205_), .A2(new_n7198_), .ZN(new_n7206_));
  OAI22_X1   g07014(.A1(new_n7199_), .A2(new_n3481_), .B1(new_n7197_), .B2(new_n7191_), .ZN(new_n7207_));
  NAND2_X1   g07015(.A1(new_n6982_), .A2(\asqrt[43] ), .ZN(new_n7208_));
  NOR4_X1    g07016(.A1(new_n7110_), .A2(\asqrt[43] ), .A3(new_n6819_), .A4(new_n6982_), .ZN(new_n7209_));
  XOR2_X1    g07017(.A1(new_n7209_), .A2(new_n7208_), .Z(new_n7210_));
  NAND2_X1   g07018(.A1(new_n7210_), .A2(new_n2941_), .ZN(new_n7211_));
  AOI21_X1   g07019(.A1(new_n7207_), .A2(\asqrt[43] ), .B(new_n7211_), .ZN(new_n7212_));
  NOR2_X1    g07020(.A1(new_n7212_), .A2(new_n7206_), .ZN(new_n7213_));
  AOI22_X1   g07021(.A1(new_n7207_), .A2(\asqrt[43] ), .B1(new_n7205_), .B2(new_n7198_), .ZN(new_n7214_));
  NOR4_X1    g07022(.A1(new_n7110_), .A2(\asqrt[44] ), .A3(new_n6826_), .A4(new_n6831_), .ZN(new_n7215_));
  AOI21_X1   g07023(.A1(new_n7208_), .A2(new_n6981_), .B(new_n2941_), .ZN(new_n7216_));
  NOR2_X1    g07024(.A1(new_n7215_), .A2(new_n7216_), .ZN(new_n7217_));
  NAND2_X1   g07025(.A1(new_n7217_), .A2(new_n2728_), .ZN(new_n7218_));
  INV_X1     g07026(.I(new_n7218_), .ZN(new_n7219_));
  OAI21_X1   g07027(.A1(new_n7214_), .A2(new_n2941_), .B(new_n7219_), .ZN(new_n7220_));
  NAND2_X1   g07028(.A1(new_n7220_), .A2(new_n7213_), .ZN(new_n7221_));
  OAI22_X1   g07029(.A1(new_n7214_), .A2(new_n2941_), .B1(new_n7212_), .B2(new_n7206_), .ZN(new_n7222_));
  NAND2_X1   g07030(.A1(new_n6989_), .A2(\asqrt[45] ), .ZN(new_n7223_));
  NOR4_X1    g07031(.A1(new_n7110_), .A2(\asqrt[45] ), .A3(new_n6834_), .A4(new_n6989_), .ZN(new_n7224_));
  XOR2_X1    g07032(.A1(new_n7224_), .A2(new_n7223_), .Z(new_n7225_));
  NAND2_X1   g07033(.A1(new_n7225_), .A2(new_n2488_), .ZN(new_n7226_));
  AOI21_X1   g07034(.A1(new_n7222_), .A2(\asqrt[45] ), .B(new_n7226_), .ZN(new_n7227_));
  NOR2_X1    g07035(.A1(new_n7227_), .A2(new_n7221_), .ZN(new_n7228_));
  AOI22_X1   g07036(.A1(new_n7222_), .A2(\asqrt[45] ), .B1(new_n7220_), .B2(new_n7213_), .ZN(new_n7229_));
  NOR4_X1    g07037(.A1(new_n7110_), .A2(\asqrt[46] ), .A3(new_n6841_), .A4(new_n6846_), .ZN(new_n7230_));
  AOI21_X1   g07038(.A1(new_n7223_), .A2(new_n6988_), .B(new_n2488_), .ZN(new_n7231_));
  NOR2_X1    g07039(.A1(new_n7230_), .A2(new_n7231_), .ZN(new_n7232_));
  NAND2_X1   g07040(.A1(new_n7232_), .A2(new_n2253_), .ZN(new_n7233_));
  INV_X1     g07041(.I(new_n7233_), .ZN(new_n7234_));
  OAI21_X1   g07042(.A1(new_n7229_), .A2(new_n2488_), .B(new_n7234_), .ZN(new_n7235_));
  NAND2_X1   g07043(.A1(new_n7235_), .A2(new_n7228_), .ZN(new_n7236_));
  OAI22_X1   g07044(.A1(new_n7229_), .A2(new_n2488_), .B1(new_n7227_), .B2(new_n7221_), .ZN(new_n7237_));
  NAND2_X1   g07045(.A1(new_n6996_), .A2(\asqrt[47] ), .ZN(new_n7238_));
  NOR4_X1    g07046(.A1(new_n7110_), .A2(\asqrt[47] ), .A3(new_n6849_), .A4(new_n6996_), .ZN(new_n7239_));
  XOR2_X1    g07047(.A1(new_n7239_), .A2(new_n7238_), .Z(new_n7240_));
  NAND2_X1   g07048(.A1(new_n7240_), .A2(new_n2046_), .ZN(new_n7241_));
  AOI21_X1   g07049(.A1(new_n7237_), .A2(\asqrt[47] ), .B(new_n7241_), .ZN(new_n7242_));
  NOR2_X1    g07050(.A1(new_n7242_), .A2(new_n7236_), .ZN(new_n7243_));
  AOI22_X1   g07051(.A1(new_n7237_), .A2(\asqrt[47] ), .B1(new_n7235_), .B2(new_n7228_), .ZN(new_n7244_));
  NOR4_X1    g07052(.A1(new_n7110_), .A2(\asqrt[48] ), .A3(new_n6856_), .A4(new_n6861_), .ZN(new_n7245_));
  AOI21_X1   g07053(.A1(new_n7238_), .A2(new_n6995_), .B(new_n2046_), .ZN(new_n7246_));
  NOR2_X1    g07054(.A1(new_n7245_), .A2(new_n7246_), .ZN(new_n7247_));
  NAND2_X1   g07055(.A1(new_n7247_), .A2(new_n1854_), .ZN(new_n7248_));
  INV_X1     g07056(.I(new_n7248_), .ZN(new_n7249_));
  OAI21_X1   g07057(.A1(new_n7244_), .A2(new_n2046_), .B(new_n7249_), .ZN(new_n7250_));
  NAND2_X1   g07058(.A1(new_n7250_), .A2(new_n7243_), .ZN(new_n7251_));
  OAI22_X1   g07059(.A1(new_n7244_), .A2(new_n2046_), .B1(new_n7242_), .B2(new_n7236_), .ZN(new_n7252_));
  NAND2_X1   g07060(.A1(new_n7003_), .A2(\asqrt[49] ), .ZN(new_n7253_));
  NOR4_X1    g07061(.A1(new_n7110_), .A2(\asqrt[49] ), .A3(new_n6864_), .A4(new_n7003_), .ZN(new_n7254_));
  XOR2_X1    g07062(.A1(new_n7254_), .A2(new_n7253_), .Z(new_n7255_));
  NAND2_X1   g07063(.A1(new_n7255_), .A2(new_n1595_), .ZN(new_n7256_));
  AOI21_X1   g07064(.A1(new_n7252_), .A2(\asqrt[49] ), .B(new_n7256_), .ZN(new_n7257_));
  NOR2_X1    g07065(.A1(new_n7257_), .A2(new_n7251_), .ZN(new_n7258_));
  AOI22_X1   g07066(.A1(new_n7252_), .A2(\asqrt[49] ), .B1(new_n7250_), .B2(new_n7243_), .ZN(new_n7259_));
  NOR4_X1    g07067(.A1(new_n7110_), .A2(\asqrt[50] ), .A3(new_n6871_), .A4(new_n6876_), .ZN(new_n7260_));
  AOI21_X1   g07068(.A1(new_n7253_), .A2(new_n7002_), .B(new_n1595_), .ZN(new_n7261_));
  NOR2_X1    g07069(.A1(new_n7260_), .A2(new_n7261_), .ZN(new_n7262_));
  NAND2_X1   g07070(.A1(new_n7262_), .A2(new_n1436_), .ZN(new_n7263_));
  INV_X1     g07071(.I(new_n7263_), .ZN(new_n7264_));
  OAI21_X1   g07072(.A1(new_n7259_), .A2(new_n1595_), .B(new_n7264_), .ZN(new_n7265_));
  NAND2_X1   g07073(.A1(new_n7265_), .A2(new_n7258_), .ZN(new_n7266_));
  OAI22_X1   g07074(.A1(new_n7259_), .A2(new_n1595_), .B1(new_n7257_), .B2(new_n7251_), .ZN(new_n7267_));
  NAND2_X1   g07075(.A1(new_n7010_), .A2(\asqrt[51] ), .ZN(new_n7268_));
  NOR4_X1    g07076(.A1(new_n7110_), .A2(\asqrt[51] ), .A3(new_n6879_), .A4(new_n7010_), .ZN(new_n7269_));
  XOR2_X1    g07077(.A1(new_n7269_), .A2(new_n7268_), .Z(new_n7270_));
  NAND2_X1   g07078(.A1(new_n7270_), .A2(new_n1260_), .ZN(new_n7271_));
  AOI21_X1   g07079(.A1(new_n7267_), .A2(\asqrt[51] ), .B(new_n7271_), .ZN(new_n7272_));
  NOR2_X1    g07080(.A1(new_n7272_), .A2(new_n7266_), .ZN(new_n7273_));
  AOI22_X1   g07081(.A1(new_n7267_), .A2(\asqrt[51] ), .B1(new_n7265_), .B2(new_n7258_), .ZN(new_n7274_));
  NAND2_X1   g07082(.A1(new_n6891_), .A2(\asqrt[52] ), .ZN(new_n7275_));
  NOR4_X1    g07083(.A1(new_n7110_), .A2(\asqrt[52] ), .A3(new_n6886_), .A4(new_n6891_), .ZN(new_n7276_));
  XOR2_X1    g07084(.A1(new_n7276_), .A2(new_n7275_), .Z(new_n7277_));
  NAND2_X1   g07085(.A1(new_n7277_), .A2(new_n1096_), .ZN(new_n7278_));
  INV_X1     g07086(.I(new_n7278_), .ZN(new_n7279_));
  OAI21_X1   g07087(.A1(new_n7274_), .A2(new_n1260_), .B(new_n7279_), .ZN(new_n7280_));
  NAND2_X1   g07088(.A1(new_n7280_), .A2(new_n7273_), .ZN(new_n7281_));
  OAI22_X1   g07089(.A1(new_n7274_), .A2(new_n1260_), .B1(new_n7272_), .B2(new_n7266_), .ZN(new_n7282_));
  NOR4_X1    g07090(.A1(new_n7110_), .A2(\asqrt[53] ), .A3(new_n6894_), .A4(new_n7017_), .ZN(new_n7283_));
  XOR2_X1    g07091(.A1(new_n7283_), .A2(new_n7031_), .Z(new_n7284_));
  NAND2_X1   g07092(.A1(new_n7284_), .A2(new_n970_), .ZN(new_n7285_));
  AOI21_X1   g07093(.A1(new_n7282_), .A2(\asqrt[53] ), .B(new_n7285_), .ZN(new_n7286_));
  NOR2_X1    g07094(.A1(new_n7286_), .A2(new_n7281_), .ZN(new_n7287_));
  AOI22_X1   g07095(.A1(new_n7282_), .A2(\asqrt[53] ), .B1(new_n7280_), .B2(new_n7273_), .ZN(new_n7288_));
  NOR4_X1    g07096(.A1(new_n7110_), .A2(\asqrt[54] ), .A3(new_n6901_), .A4(new_n6906_), .ZN(new_n7289_));
  XOR2_X1    g07097(.A1(new_n7289_), .A2(new_n6944_), .Z(new_n7290_));
  NAND2_X1   g07098(.A1(new_n7290_), .A2(new_n825_), .ZN(new_n7291_));
  INV_X1     g07099(.I(new_n7291_), .ZN(new_n7292_));
  OAI21_X1   g07100(.A1(new_n7288_), .A2(new_n970_), .B(new_n7292_), .ZN(new_n7293_));
  NAND2_X1   g07101(.A1(new_n7293_), .A2(new_n7287_), .ZN(new_n7294_));
  OAI22_X1   g07102(.A1(new_n7288_), .A2(new_n970_), .B1(new_n7286_), .B2(new_n7281_), .ZN(new_n7295_));
  NOR4_X1    g07103(.A1(new_n7110_), .A2(\asqrt[55] ), .A3(new_n6908_), .A4(new_n7024_), .ZN(new_n7296_));
  XOR2_X1    g07104(.A1(new_n7296_), .A2(new_n7033_), .Z(new_n7297_));
  NAND2_X1   g07105(.A1(new_n7297_), .A2(new_n724_), .ZN(new_n7298_));
  AOI21_X1   g07106(.A1(new_n7295_), .A2(\asqrt[55] ), .B(new_n7298_), .ZN(new_n7299_));
  NOR2_X1    g07107(.A1(new_n7299_), .A2(new_n7294_), .ZN(new_n7300_));
  AOI22_X1   g07108(.A1(new_n7295_), .A2(\asqrt[55] ), .B1(new_n7293_), .B2(new_n7287_), .ZN(new_n7301_));
  NOR4_X1    g07109(.A1(new_n7110_), .A2(\asqrt[56] ), .A3(new_n6914_), .A4(new_n6919_), .ZN(new_n7302_));
  XOR2_X1    g07110(.A1(new_n7302_), .A2(new_n6946_), .Z(new_n7303_));
  NAND2_X1   g07111(.A1(new_n7303_), .A2(new_n587_), .ZN(new_n7304_));
  INV_X1     g07112(.I(new_n7304_), .ZN(new_n7305_));
  OAI21_X1   g07113(.A1(new_n7301_), .A2(new_n724_), .B(new_n7305_), .ZN(new_n7306_));
  NAND2_X1   g07114(.A1(new_n7306_), .A2(new_n7300_), .ZN(new_n7307_));
  OAI22_X1   g07115(.A1(new_n7301_), .A2(new_n724_), .B1(new_n7299_), .B2(new_n7294_), .ZN(new_n7308_));
  NOR4_X1    g07116(.A1(new_n7110_), .A2(\asqrt[57] ), .A3(new_n6921_), .A4(new_n7037_), .ZN(new_n7309_));
  XOR2_X1    g07117(.A1(new_n7309_), .A2(new_n7035_), .Z(new_n7310_));
  NAND2_X1   g07118(.A1(new_n7310_), .A2(new_n504_), .ZN(new_n7311_));
  AOI21_X1   g07119(.A1(new_n7308_), .A2(\asqrt[57] ), .B(new_n7311_), .ZN(new_n7312_));
  NOR2_X1    g07120(.A1(new_n7312_), .A2(new_n7307_), .ZN(new_n7313_));
  AOI22_X1   g07121(.A1(new_n7308_), .A2(\asqrt[57] ), .B1(new_n7306_), .B2(new_n7300_), .ZN(new_n7314_));
  NOR4_X1    g07122(.A1(new_n7110_), .A2(\asqrt[58] ), .A3(new_n6927_), .A4(new_n6932_), .ZN(new_n7315_));
  XOR2_X1    g07123(.A1(new_n7315_), .A2(new_n6948_), .Z(new_n7316_));
  NAND2_X1   g07124(.A1(new_n7316_), .A2(new_n376_), .ZN(new_n7317_));
  INV_X1     g07125(.I(new_n7317_), .ZN(new_n7318_));
  OAI21_X1   g07126(.A1(new_n7314_), .A2(new_n504_), .B(new_n7318_), .ZN(new_n7319_));
  NAND2_X1   g07127(.A1(new_n7319_), .A2(new_n7313_), .ZN(new_n7320_));
  OAI22_X1   g07128(.A1(new_n7314_), .A2(new_n504_), .B1(new_n7312_), .B2(new_n7307_), .ZN(new_n7321_));
  NOR4_X1    g07129(.A1(new_n7110_), .A2(\asqrt[59] ), .A3(new_n6934_), .A4(new_n7045_), .ZN(new_n7322_));
  XOR2_X1    g07130(.A1(new_n7322_), .A2(new_n7043_), .Z(new_n7323_));
  NAND2_X1   g07131(.A1(new_n7323_), .A2(new_n275_), .ZN(new_n7324_));
  AOI21_X1   g07132(.A1(new_n7321_), .A2(\asqrt[59] ), .B(new_n7324_), .ZN(new_n7325_));
  NOR2_X1    g07133(.A1(new_n7325_), .A2(new_n7320_), .ZN(new_n7326_));
  AOI22_X1   g07134(.A1(new_n7321_), .A2(\asqrt[59] ), .B1(new_n7319_), .B2(new_n7313_), .ZN(new_n7327_));
  OAI22_X1   g07135(.A1(new_n7327_), .A2(new_n275_), .B1(new_n7325_), .B2(new_n7320_), .ZN(new_n7328_));
  NOR4_X1    g07136(.A1(new_n7110_), .A2(\asqrt[60] ), .A3(new_n6940_), .A4(new_n7067_), .ZN(new_n7329_));
  XOR2_X1    g07137(.A1(new_n7329_), .A2(new_n6950_), .Z(new_n7330_));
  NAND2_X1   g07138(.A1(new_n7330_), .A2(new_n229_), .ZN(new_n7331_));
  INV_X1     g07139(.I(new_n7331_), .ZN(new_n7332_));
  OAI21_X1   g07140(.A1(new_n7327_), .A2(new_n275_), .B(new_n7332_), .ZN(new_n7333_));
  AOI22_X1   g07141(.A1(new_n7328_), .A2(\asqrt[61] ), .B1(new_n7333_), .B2(new_n7326_), .ZN(new_n7334_));
  NOR2_X1    g07142(.A1(new_n7334_), .A2(new_n196_), .ZN(new_n7335_));
  INV_X1     g07143(.I(new_n7087_), .ZN(new_n7336_));
  AOI21_X1   g07144(.A1(new_n7101_), .A2(new_n7336_), .B(new_n7089_), .ZN(new_n7337_));
  NOR3_X1    g07145(.A1(new_n7086_), .A2(new_n7081_), .A3(new_n7085_), .ZN(new_n7338_));
  NOR2_X1    g07146(.A1(new_n7338_), .A2(new_n7337_), .ZN(new_n7339_));
  NOR3_X1    g07147(.A1(new_n7124_), .A2(new_n6309_), .A3(\asqrt[31] ), .ZN(new_n7340_));
  AOI21_X1   g07148(.A1(new_n7118_), .A2(new_n6308_), .B(new_n7110_), .ZN(new_n7341_));
  NOR4_X1    g07149(.A1(new_n7341_), .A2(new_n7340_), .A3(\asqrt[33] ), .A4(new_n7108_), .ZN(new_n7342_));
  NOR2_X1    g07150(.A1(new_n7342_), .A2(new_n7339_), .ZN(new_n7343_));
  NOR3_X1    g07151(.A1(new_n7338_), .A2(new_n7337_), .A3(new_n7108_), .ZN(new_n7344_));
  NOR3_X1    g07152(.A1(new_n7110_), .A2(new_n6706_), .A3(new_n7134_), .ZN(new_n7345_));
  AOI21_X1   g07153(.A1(\asqrt[31] ), .A2(new_n7132_), .B(new_n6707_), .ZN(new_n7346_));
  NOR3_X1    g07154(.A1(new_n7346_), .A2(new_n7345_), .A3(\asqrt[34] ), .ZN(new_n7347_));
  OAI21_X1   g07155(.A1(new_n7344_), .A2(new_n6365_), .B(new_n7347_), .ZN(new_n7348_));
  NAND2_X1   g07156(.A1(new_n7343_), .A2(new_n7348_), .ZN(new_n7349_));
  OAI22_X1   g07157(.A1(new_n7342_), .A2(new_n7339_), .B1(new_n6365_), .B2(new_n7344_), .ZN(new_n7350_));
  INV_X1     g07158(.I(new_n7147_), .ZN(new_n7351_));
  AOI21_X1   g07159(.A1(new_n7350_), .A2(\asqrt[34] ), .B(new_n7351_), .ZN(new_n7352_));
  NOR2_X1    g07160(.A1(new_n7352_), .A2(new_n7349_), .ZN(new_n7353_));
  AOI22_X1   g07161(.A1(new_n7350_), .A2(\asqrt[34] ), .B1(new_n7343_), .B2(new_n7348_), .ZN(new_n7354_));
  INV_X1     g07162(.I(new_n7154_), .ZN(new_n7355_));
  OAI21_X1   g07163(.A1(new_n7354_), .A2(new_n5626_), .B(new_n7355_), .ZN(new_n7356_));
  NAND2_X1   g07164(.A1(new_n7356_), .A2(new_n7353_), .ZN(new_n7357_));
  OAI22_X1   g07165(.A1(new_n7354_), .A2(new_n5626_), .B1(new_n7352_), .B2(new_n7349_), .ZN(new_n7358_));
  AOI21_X1   g07166(.A1(new_n7358_), .A2(\asqrt[36] ), .B(new_n7161_), .ZN(new_n7359_));
  NOR2_X1    g07167(.A1(new_n7359_), .A2(new_n7357_), .ZN(new_n7360_));
  AOI22_X1   g07168(.A1(new_n7358_), .A2(\asqrt[36] ), .B1(new_n7356_), .B2(new_n7353_), .ZN(new_n7361_));
  INV_X1     g07169(.I(new_n7169_), .ZN(new_n7362_));
  OAI21_X1   g07170(.A1(new_n7361_), .A2(new_n4973_), .B(new_n7362_), .ZN(new_n7363_));
  NAND2_X1   g07171(.A1(new_n7363_), .A2(new_n7360_), .ZN(new_n7364_));
  OAI22_X1   g07172(.A1(new_n7361_), .A2(new_n4973_), .B1(new_n7359_), .B2(new_n7357_), .ZN(new_n7365_));
  AOI21_X1   g07173(.A1(new_n7365_), .A2(\asqrt[38] ), .B(new_n7175_), .ZN(new_n7366_));
  NOR2_X1    g07174(.A1(new_n7366_), .A2(new_n7364_), .ZN(new_n7367_));
  AOI22_X1   g07175(.A1(new_n7365_), .A2(\asqrt[38] ), .B1(new_n7363_), .B2(new_n7360_), .ZN(new_n7368_));
  INV_X1     g07176(.I(new_n7182_), .ZN(new_n7369_));
  OAI21_X1   g07177(.A1(new_n7368_), .A2(new_n4330_), .B(new_n7369_), .ZN(new_n7370_));
  NAND2_X1   g07178(.A1(new_n7370_), .A2(new_n7367_), .ZN(new_n7371_));
  OAI22_X1   g07179(.A1(new_n7368_), .A2(new_n4330_), .B1(new_n7366_), .B2(new_n7364_), .ZN(new_n7372_));
  AOI21_X1   g07180(.A1(new_n7372_), .A2(\asqrt[40] ), .B(new_n7188_), .ZN(new_n7373_));
  NOR2_X1    g07181(.A1(new_n7373_), .A2(new_n7371_), .ZN(new_n7374_));
  AOI22_X1   g07182(.A1(new_n7372_), .A2(\asqrt[40] ), .B1(new_n7370_), .B2(new_n7367_), .ZN(new_n7375_));
  INV_X1     g07183(.I(new_n7196_), .ZN(new_n7376_));
  OAI21_X1   g07184(.A1(new_n7375_), .A2(new_n3760_), .B(new_n7376_), .ZN(new_n7377_));
  NAND2_X1   g07185(.A1(new_n7377_), .A2(new_n7374_), .ZN(new_n7378_));
  OAI22_X1   g07186(.A1(new_n7375_), .A2(new_n3760_), .B1(new_n7373_), .B2(new_n7371_), .ZN(new_n7379_));
  AOI21_X1   g07187(.A1(new_n7379_), .A2(\asqrt[42] ), .B(new_n7203_), .ZN(new_n7380_));
  NOR2_X1    g07188(.A1(new_n7380_), .A2(new_n7378_), .ZN(new_n7381_));
  AOI22_X1   g07189(.A1(new_n7379_), .A2(\asqrt[42] ), .B1(new_n7377_), .B2(new_n7374_), .ZN(new_n7382_));
  INV_X1     g07190(.I(new_n7211_), .ZN(new_n7383_));
  OAI21_X1   g07191(.A1(new_n7382_), .A2(new_n3208_), .B(new_n7383_), .ZN(new_n7384_));
  NAND2_X1   g07192(.A1(new_n7384_), .A2(new_n7381_), .ZN(new_n7385_));
  OAI22_X1   g07193(.A1(new_n7382_), .A2(new_n3208_), .B1(new_n7380_), .B2(new_n7378_), .ZN(new_n7386_));
  AOI21_X1   g07194(.A1(new_n7386_), .A2(\asqrt[44] ), .B(new_n7218_), .ZN(new_n7387_));
  NOR2_X1    g07195(.A1(new_n7387_), .A2(new_n7385_), .ZN(new_n7388_));
  AOI22_X1   g07196(.A1(new_n7386_), .A2(\asqrt[44] ), .B1(new_n7384_), .B2(new_n7381_), .ZN(new_n7389_));
  INV_X1     g07197(.I(new_n7226_), .ZN(new_n7390_));
  OAI21_X1   g07198(.A1(new_n7389_), .A2(new_n2728_), .B(new_n7390_), .ZN(new_n7391_));
  NAND2_X1   g07199(.A1(new_n7391_), .A2(new_n7388_), .ZN(new_n7392_));
  OAI22_X1   g07200(.A1(new_n7389_), .A2(new_n2728_), .B1(new_n7387_), .B2(new_n7385_), .ZN(new_n7393_));
  AOI21_X1   g07201(.A1(new_n7393_), .A2(\asqrt[46] ), .B(new_n7233_), .ZN(new_n7394_));
  NOR2_X1    g07202(.A1(new_n7394_), .A2(new_n7392_), .ZN(new_n7395_));
  AOI22_X1   g07203(.A1(new_n7393_), .A2(\asqrt[46] ), .B1(new_n7391_), .B2(new_n7388_), .ZN(new_n7396_));
  INV_X1     g07204(.I(new_n7241_), .ZN(new_n7397_));
  OAI21_X1   g07205(.A1(new_n7396_), .A2(new_n2253_), .B(new_n7397_), .ZN(new_n7398_));
  NAND2_X1   g07206(.A1(new_n7398_), .A2(new_n7395_), .ZN(new_n7399_));
  OAI22_X1   g07207(.A1(new_n7396_), .A2(new_n2253_), .B1(new_n7394_), .B2(new_n7392_), .ZN(new_n7400_));
  AOI21_X1   g07208(.A1(new_n7400_), .A2(\asqrt[48] ), .B(new_n7248_), .ZN(new_n7401_));
  NOR2_X1    g07209(.A1(new_n7401_), .A2(new_n7399_), .ZN(new_n7402_));
  AOI22_X1   g07210(.A1(new_n7400_), .A2(\asqrt[48] ), .B1(new_n7398_), .B2(new_n7395_), .ZN(new_n7403_));
  INV_X1     g07211(.I(new_n7256_), .ZN(new_n7404_));
  OAI21_X1   g07212(.A1(new_n7403_), .A2(new_n1854_), .B(new_n7404_), .ZN(new_n7405_));
  NAND2_X1   g07213(.A1(new_n7405_), .A2(new_n7402_), .ZN(new_n7406_));
  OAI22_X1   g07214(.A1(new_n7403_), .A2(new_n1854_), .B1(new_n7401_), .B2(new_n7399_), .ZN(new_n7407_));
  AOI21_X1   g07215(.A1(new_n7407_), .A2(\asqrt[50] ), .B(new_n7263_), .ZN(new_n7408_));
  NOR2_X1    g07216(.A1(new_n7408_), .A2(new_n7406_), .ZN(new_n7409_));
  AOI22_X1   g07217(.A1(new_n7407_), .A2(\asqrt[50] ), .B1(new_n7405_), .B2(new_n7402_), .ZN(new_n7410_));
  INV_X1     g07218(.I(new_n7271_), .ZN(new_n7411_));
  OAI21_X1   g07219(.A1(new_n7410_), .A2(new_n1436_), .B(new_n7411_), .ZN(new_n7412_));
  NAND2_X1   g07220(.A1(new_n7412_), .A2(new_n7409_), .ZN(new_n7413_));
  OAI22_X1   g07221(.A1(new_n7410_), .A2(new_n1436_), .B1(new_n7408_), .B2(new_n7406_), .ZN(new_n7414_));
  AOI21_X1   g07222(.A1(new_n7414_), .A2(\asqrt[52] ), .B(new_n7278_), .ZN(new_n7415_));
  NOR2_X1    g07223(.A1(new_n7415_), .A2(new_n7413_), .ZN(new_n7416_));
  AOI22_X1   g07224(.A1(new_n7414_), .A2(\asqrt[52] ), .B1(new_n7412_), .B2(new_n7409_), .ZN(new_n7417_));
  INV_X1     g07225(.I(new_n7285_), .ZN(new_n7418_));
  OAI21_X1   g07226(.A1(new_n7417_), .A2(new_n1096_), .B(new_n7418_), .ZN(new_n7419_));
  NAND2_X1   g07227(.A1(new_n7419_), .A2(new_n7416_), .ZN(new_n7420_));
  OAI22_X1   g07228(.A1(new_n7417_), .A2(new_n1096_), .B1(new_n7415_), .B2(new_n7413_), .ZN(new_n7421_));
  AOI21_X1   g07229(.A1(new_n7421_), .A2(\asqrt[54] ), .B(new_n7291_), .ZN(new_n7422_));
  NOR2_X1    g07230(.A1(new_n7422_), .A2(new_n7420_), .ZN(new_n7423_));
  AOI22_X1   g07231(.A1(new_n7421_), .A2(\asqrt[54] ), .B1(new_n7419_), .B2(new_n7416_), .ZN(new_n7424_));
  INV_X1     g07232(.I(new_n7298_), .ZN(new_n7425_));
  OAI21_X1   g07233(.A1(new_n7424_), .A2(new_n825_), .B(new_n7425_), .ZN(new_n7426_));
  NAND2_X1   g07234(.A1(new_n7426_), .A2(new_n7423_), .ZN(new_n7427_));
  OAI22_X1   g07235(.A1(new_n7424_), .A2(new_n825_), .B1(new_n7422_), .B2(new_n7420_), .ZN(new_n7428_));
  AOI21_X1   g07236(.A1(new_n7428_), .A2(\asqrt[56] ), .B(new_n7304_), .ZN(new_n7429_));
  NOR2_X1    g07237(.A1(new_n7429_), .A2(new_n7427_), .ZN(new_n7430_));
  AOI22_X1   g07238(.A1(new_n7428_), .A2(\asqrt[56] ), .B1(new_n7426_), .B2(new_n7423_), .ZN(new_n7431_));
  INV_X1     g07239(.I(new_n7311_), .ZN(new_n7432_));
  OAI21_X1   g07240(.A1(new_n7431_), .A2(new_n587_), .B(new_n7432_), .ZN(new_n7433_));
  NAND2_X1   g07241(.A1(new_n7433_), .A2(new_n7430_), .ZN(new_n7434_));
  OAI22_X1   g07242(.A1(new_n7431_), .A2(new_n587_), .B1(new_n7429_), .B2(new_n7427_), .ZN(new_n7435_));
  AOI21_X1   g07243(.A1(new_n7435_), .A2(\asqrt[58] ), .B(new_n7317_), .ZN(new_n7436_));
  NOR2_X1    g07244(.A1(new_n7436_), .A2(new_n7434_), .ZN(new_n7437_));
  AOI22_X1   g07245(.A1(new_n7435_), .A2(\asqrt[58] ), .B1(new_n7433_), .B2(new_n7430_), .ZN(new_n7438_));
  INV_X1     g07246(.I(new_n7324_), .ZN(new_n7439_));
  OAI21_X1   g07247(.A1(new_n7438_), .A2(new_n376_), .B(new_n7439_), .ZN(new_n7440_));
  NAND2_X1   g07248(.A1(new_n7440_), .A2(new_n7437_), .ZN(new_n7441_));
  OAI22_X1   g07249(.A1(new_n7438_), .A2(new_n376_), .B1(new_n7436_), .B2(new_n7434_), .ZN(new_n7442_));
  AOI22_X1   g07250(.A1(new_n7442_), .A2(\asqrt[60] ), .B1(new_n7440_), .B2(new_n7437_), .ZN(new_n7443_));
  AOI21_X1   g07251(.A1(new_n7442_), .A2(\asqrt[60] ), .B(new_n7331_), .ZN(new_n7444_));
  OAI22_X1   g07252(.A1(new_n7443_), .A2(new_n229_), .B1(new_n7444_), .B2(new_n7441_), .ZN(new_n7445_));
  NOR2_X1    g07253(.A1(new_n7445_), .A2(\asqrt[62] ), .ZN(new_n7446_));
  NAND3_X1   g07254(.A1(new_n7104_), .A2(new_n6957_), .A3(new_n7073_), .ZN(new_n7447_));
  NOR2_X1    g07255(.A1(new_n7113_), .A2(new_n196_), .ZN(new_n7448_));
  INV_X1     g07256(.I(new_n7098_), .ZN(new_n7449_));
  NAND3_X1   g07257(.A1(\asqrt[31] ), .A2(new_n7448_), .A3(new_n7449_), .ZN(new_n7450_));
  OAI21_X1   g07258(.A1(new_n7070_), .A2(\asqrt[62] ), .B(new_n6959_), .ZN(new_n7451_));
  OAI21_X1   g07259(.A1(\asqrt[31] ), .A2(new_n7451_), .B(new_n7448_), .ZN(new_n7452_));
  NAND2_X1   g07260(.A1(new_n7452_), .A2(new_n7450_), .ZN(new_n7453_));
  INV_X1     g07261(.I(new_n7453_), .ZN(new_n7454_));
  NOR2_X1    g07262(.A1(new_n7078_), .A2(new_n196_), .ZN(new_n7455_));
  INV_X1     g07263(.I(new_n7455_), .ZN(new_n7456_));
  NAND2_X1   g07264(.A1(new_n7308_), .A2(\asqrt[57] ), .ZN(new_n7457_));
  AOI21_X1   g07265(.A1(new_n7457_), .A2(new_n7307_), .B(new_n504_), .ZN(new_n7458_));
  OAI21_X1   g07266(.A1(new_n7313_), .A2(new_n7458_), .B(\asqrt[59] ), .ZN(new_n7459_));
  AOI21_X1   g07267(.A1(new_n7320_), .A2(new_n7459_), .B(new_n275_), .ZN(new_n7460_));
  OAI21_X1   g07268(.A1(new_n7326_), .A2(new_n7460_), .B(\asqrt[61] ), .ZN(new_n7461_));
  NOR2_X1    g07269(.A1(new_n7079_), .A2(\asqrt[62] ), .ZN(new_n7462_));
  INV_X1     g07270(.I(new_n7462_), .ZN(new_n7463_));
  NAND3_X1   g07271(.A1(new_n7333_), .A2(new_n7326_), .A3(new_n7463_), .ZN(new_n7464_));
  OAI21_X1   g07272(.A1(new_n7464_), .A2(new_n7461_), .B(new_n7456_), .ZN(new_n7465_));
  NAND3_X1   g07273(.A1(new_n7110_), .A2(new_n7066_), .A3(new_n7114_), .ZN(new_n7466_));
  AOI21_X1   g07274(.A1(new_n7466_), .A2(new_n7057_), .B(\asqrt[63] ), .ZN(new_n7467_));
  INV_X1     g07275(.I(new_n7467_), .ZN(new_n7468_));
  OAI21_X1   g07276(.A1(new_n7465_), .A2(new_n7468_), .B(new_n7454_), .ZN(new_n7469_));
  NOR4_X1    g07277(.A1(new_n7445_), .A2(\asqrt[62] ), .A3(new_n7453_), .A4(new_n7078_), .ZN(new_n7470_));
  NAND2_X1   g07278(.A1(new_n7092_), .A2(new_n7066_), .ZN(new_n7471_));
  XOR2_X1    g07279(.A1(new_n7092_), .A2(\asqrt[63] ), .Z(new_n7472_));
  AOI21_X1   g07280(.A1(\asqrt[31] ), .A2(new_n7471_), .B(new_n7472_), .ZN(new_n7473_));
  NAND2_X1   g07281(.A1(new_n7470_), .A2(new_n7473_), .ZN(new_n7474_));
  NOR3_X1    g07282(.A1(new_n7474_), .A2(new_n7447_), .A3(new_n7469_), .ZN(\asqrt[30] ));
  NAND4_X1   g07283(.A1(\asqrt[30] ), .A2(new_n7079_), .A3(new_n7335_), .A4(new_n7446_), .ZN(new_n7476_));
  OAI21_X1   g07284(.A1(new_n7445_), .A2(\asqrt[62] ), .B(new_n7078_), .ZN(new_n7477_));
  OAI21_X1   g07285(.A1(\asqrt[30] ), .A2(new_n7477_), .B(new_n7335_), .ZN(new_n7478_));
  NAND2_X1   g07286(.A1(new_n7476_), .A2(new_n7478_), .ZN(new_n7479_));
  INV_X1     g07287(.I(new_n7479_), .ZN(new_n7480_));
  NAND2_X1   g07288(.A1(new_n7435_), .A2(\asqrt[58] ), .ZN(new_n7481_));
  AOI21_X1   g07289(.A1(new_n7481_), .A2(new_n7434_), .B(new_n376_), .ZN(new_n7482_));
  OAI21_X1   g07290(.A1(new_n7437_), .A2(new_n7482_), .B(\asqrt[60] ), .ZN(new_n7483_));
  AOI21_X1   g07291(.A1(new_n7441_), .A2(new_n7483_), .B(new_n229_), .ZN(new_n7484_));
  NOR3_X1    g07292(.A1(new_n7328_), .A2(\asqrt[61] ), .A3(new_n7330_), .ZN(new_n7485_));
  NAND2_X1   g07293(.A1(\asqrt[30] ), .A2(new_n7485_), .ZN(new_n7486_));
  XOR2_X1    g07294(.A1(new_n7486_), .A2(new_n7484_), .Z(new_n7487_));
  NOR2_X1    g07295(.A1(new_n7487_), .A2(new_n196_), .ZN(new_n7488_));
  INV_X1     g07296(.I(new_n7488_), .ZN(new_n7489_));
  INV_X1     g07297(.I(\a[60] ), .ZN(new_n7490_));
  NOR2_X1    g07298(.A1(\a[58] ), .A2(\a[59] ), .ZN(new_n7491_));
  INV_X1     g07299(.I(new_n7491_), .ZN(new_n7492_));
  NOR3_X1    g07300(.A1(new_n7116_), .A2(new_n7490_), .A3(new_n7492_), .ZN(new_n7493_));
  NAND2_X1   g07301(.A1(new_n7122_), .A2(new_n7493_), .ZN(new_n7494_));
  XOR2_X1    g07302(.A1(new_n7494_), .A2(\a[61] ), .Z(new_n7495_));
  INV_X1     g07303(.I(\a[61] ), .ZN(new_n7496_));
  NOR4_X1    g07304(.A1(new_n7474_), .A2(new_n7496_), .A3(new_n7447_), .A4(new_n7469_), .ZN(new_n7497_));
  NOR2_X1    g07305(.A1(new_n7496_), .A2(\a[60] ), .ZN(new_n7498_));
  OAI21_X1   g07306(.A1(new_n7497_), .A2(new_n7498_), .B(new_n7495_), .ZN(new_n7499_));
  INV_X1     g07307(.I(new_n7495_), .ZN(new_n7500_));
  INV_X1     g07308(.I(new_n7447_), .ZN(new_n7501_));
  NOR3_X1    g07309(.A1(new_n7444_), .A2(new_n7441_), .A3(new_n7462_), .ZN(new_n7502_));
  AOI21_X1   g07310(.A1(new_n7502_), .A2(new_n7484_), .B(new_n7455_), .ZN(new_n7503_));
  AOI21_X1   g07311(.A1(new_n7503_), .A2(new_n7467_), .B(new_n7453_), .ZN(new_n7504_));
  NAND4_X1   g07312(.A1(new_n7334_), .A2(new_n196_), .A3(new_n7454_), .A4(new_n7079_), .ZN(new_n7505_));
  INV_X1     g07313(.I(new_n7473_), .ZN(new_n7506_));
  NOR2_X1    g07314(.A1(new_n7505_), .A2(new_n7506_), .ZN(new_n7507_));
  NAND4_X1   g07315(.A1(new_n7507_), .A2(\a[61] ), .A3(new_n7504_), .A4(new_n7501_), .ZN(new_n7508_));
  NAND3_X1   g07316(.A1(new_n7508_), .A2(\a[60] ), .A3(new_n7500_), .ZN(new_n7509_));
  NAND2_X1   g07317(.A1(new_n7499_), .A2(new_n7509_), .ZN(new_n7510_));
  NOR2_X1    g07318(.A1(new_n7474_), .A2(new_n7469_), .ZN(new_n7511_));
  NOR4_X1    g07319(.A1(new_n7072_), .A2(new_n7066_), .A3(new_n7112_), .A4(new_n7073_), .ZN(new_n7512_));
  NAND2_X1   g07320(.A1(\asqrt[31] ), .A2(\a[60] ), .ZN(new_n7513_));
  XOR2_X1    g07321(.A1(new_n7513_), .A2(new_n7512_), .Z(new_n7514_));
  NOR2_X1    g07322(.A1(new_n7514_), .A2(new_n7492_), .ZN(new_n7515_));
  INV_X1     g07323(.I(new_n7515_), .ZN(new_n7516_));
  NAND3_X1   g07324(.A1(new_n7507_), .A2(new_n7501_), .A3(new_n7504_), .ZN(new_n7517_));
  NOR2_X1    g07325(.A1(new_n7501_), .A2(new_n7473_), .ZN(new_n7518_));
  INV_X1     g07326(.I(new_n7518_), .ZN(new_n7519_));
  NOR2_X1    g07327(.A1(new_n7519_), .A2(new_n7110_), .ZN(new_n7520_));
  NAND3_X1   g07328(.A1(new_n7469_), .A2(new_n7505_), .A3(new_n7520_), .ZN(new_n7521_));
  NAND2_X1   g07329(.A1(new_n7521_), .A2(new_n7081_), .ZN(new_n7522_));
  NAND3_X1   g07330(.A1(new_n7522_), .A2(new_n7082_), .A3(new_n7517_), .ZN(new_n7523_));
  INV_X1     g07331(.I(new_n7520_), .ZN(new_n7524_));
  NOR3_X1    g07332(.A1(new_n7504_), .A2(new_n7470_), .A3(new_n7524_), .ZN(new_n7525_));
  OAI21_X1   g07333(.A1(new_n7525_), .A2(\a[62] ), .B(new_n7082_), .ZN(new_n7526_));
  NAND2_X1   g07334(.A1(new_n7526_), .A2(\asqrt[30] ), .ZN(new_n7527_));
  NAND4_X1   g07335(.A1(new_n7527_), .A2(new_n6708_), .A3(new_n7523_), .A4(new_n7516_), .ZN(new_n7528_));
  NAND2_X1   g07336(.A1(new_n7528_), .A2(new_n7510_), .ZN(new_n7529_));
  NAND3_X1   g07337(.A1(new_n7499_), .A2(new_n7509_), .A3(new_n7516_), .ZN(new_n7530_));
  NAND2_X1   g07338(.A1(\asqrt[31] ), .A2(new_n7081_), .ZN(new_n7531_));
  AOI22_X1   g07339(.A1(new_n7531_), .A2(new_n7080_), .B1(new_n7081_), .B2(new_n7086_), .ZN(new_n7532_));
  OAI21_X1   g07340(.A1(new_n7110_), .A2(new_n7081_), .B(new_n7084_), .ZN(new_n7533_));
  NOR2_X1    g07341(.A1(new_n7532_), .A2(new_n7533_), .ZN(new_n7534_));
  NAND3_X1   g07342(.A1(\asqrt[30] ), .A2(new_n7109_), .A3(new_n7534_), .ZN(new_n7535_));
  INV_X1     g07343(.I(new_n7534_), .ZN(new_n7536_));
  OAI21_X1   g07344(.A1(new_n7517_), .A2(new_n7536_), .B(new_n7108_), .ZN(new_n7537_));
  NAND3_X1   g07345(.A1(new_n7535_), .A2(new_n7537_), .A3(new_n6365_), .ZN(new_n7538_));
  AOI21_X1   g07346(.A1(new_n7530_), .A2(\asqrt[32] ), .B(new_n7538_), .ZN(new_n7539_));
  NOR2_X1    g07347(.A1(new_n7529_), .A2(new_n7539_), .ZN(new_n7540_));
  NAND2_X1   g07348(.A1(new_n7530_), .A2(\asqrt[32] ), .ZN(new_n7541_));
  AOI21_X1   g07349(.A1(new_n7529_), .A2(new_n7541_), .B(new_n6365_), .ZN(new_n7542_));
  NOR2_X1    g07350(.A1(new_n7341_), .A2(new_n7340_), .ZN(new_n7543_));
  NOR4_X1    g07351(.A1(new_n7517_), .A2(\asqrt[33] ), .A3(new_n7543_), .A4(new_n7128_), .ZN(new_n7544_));
  AOI21_X1   g07352(.A1(new_n7339_), .A2(new_n7109_), .B(new_n6365_), .ZN(new_n7545_));
  NOR2_X1    g07353(.A1(new_n7544_), .A2(new_n7545_), .ZN(new_n7546_));
  NAND2_X1   g07354(.A1(new_n7546_), .A2(new_n5991_), .ZN(new_n7547_));
  OAI21_X1   g07355(.A1(new_n7542_), .A2(new_n7547_), .B(new_n7540_), .ZN(new_n7548_));
  AOI22_X1   g07356(.A1(new_n7528_), .A2(new_n7510_), .B1(\asqrt[32] ), .B2(new_n7530_), .ZN(new_n7549_));
  OAI22_X1   g07357(.A1(new_n7549_), .A2(new_n6365_), .B1(new_n7529_), .B2(new_n7539_), .ZN(new_n7550_));
  NOR2_X1    g07358(.A1(new_n7139_), .A2(new_n5991_), .ZN(new_n7551_));
  NAND2_X1   g07359(.A1(new_n7133_), .A2(new_n7135_), .ZN(new_n7552_));
  NAND4_X1   g07360(.A1(\asqrt[30] ), .A2(new_n5991_), .A3(new_n7552_), .A4(new_n7139_), .ZN(new_n7553_));
  XOR2_X1    g07361(.A1(new_n7553_), .A2(new_n7551_), .Z(new_n7554_));
  NAND2_X1   g07362(.A1(new_n7554_), .A2(new_n5626_), .ZN(new_n7555_));
  AOI21_X1   g07363(.A1(new_n7550_), .A2(\asqrt[34] ), .B(new_n7555_), .ZN(new_n7556_));
  OAI21_X1   g07364(.A1(new_n7542_), .A2(new_n7540_), .B(\asqrt[34] ), .ZN(new_n7557_));
  AOI21_X1   g07365(.A1(new_n7548_), .A2(new_n7557_), .B(new_n5626_), .ZN(new_n7558_));
  NAND2_X1   g07366(.A1(new_n7150_), .A2(\asqrt[35] ), .ZN(new_n7559_));
  NOR2_X1    g07367(.A1(new_n7145_), .A2(new_n7146_), .ZN(new_n7560_));
  NOR4_X1    g07368(.A1(new_n7517_), .A2(\asqrt[35] ), .A3(new_n7560_), .A4(new_n7150_), .ZN(new_n7561_));
  XOR2_X1    g07369(.A1(new_n7561_), .A2(new_n7559_), .Z(new_n7562_));
  NAND2_X1   g07370(.A1(new_n7562_), .A2(new_n5273_), .ZN(new_n7563_));
  NOR2_X1    g07371(.A1(new_n7558_), .A2(new_n7563_), .ZN(new_n7564_));
  NOR3_X1    g07372(.A1(new_n7564_), .A2(new_n7548_), .A3(new_n7556_), .ZN(new_n7565_));
  INV_X1     g07373(.I(new_n7555_), .ZN(new_n7566_));
  AOI21_X1   g07374(.A1(new_n7557_), .A2(new_n7566_), .B(new_n7548_), .ZN(new_n7567_));
  OAI21_X1   g07375(.A1(new_n7567_), .A2(new_n7558_), .B(\asqrt[36] ), .ZN(new_n7568_));
  NOR4_X1    g07376(.A1(new_n7517_), .A2(\asqrt[36] ), .A3(new_n7153_), .A4(new_n7358_), .ZN(new_n7569_));
  AOI21_X1   g07377(.A1(new_n7559_), .A2(new_n7149_), .B(new_n5273_), .ZN(new_n7570_));
  NOR2_X1    g07378(.A1(new_n7569_), .A2(new_n7570_), .ZN(new_n7571_));
  NAND2_X1   g07379(.A1(new_n7571_), .A2(new_n4973_), .ZN(new_n7572_));
  INV_X1     g07380(.I(new_n7572_), .ZN(new_n7573_));
  NAND2_X1   g07381(.A1(new_n7568_), .A2(new_n7573_), .ZN(new_n7574_));
  NAND2_X1   g07382(.A1(new_n7574_), .A2(new_n7565_), .ZN(new_n7575_));
  OAI21_X1   g07383(.A1(new_n7558_), .A2(new_n7563_), .B(new_n7567_), .ZN(new_n7576_));
  NAND2_X1   g07384(.A1(new_n7576_), .A2(new_n7568_), .ZN(new_n7577_));
  NAND2_X1   g07385(.A1(new_n7165_), .A2(\asqrt[37] ), .ZN(new_n7578_));
  NOR4_X1    g07386(.A1(new_n7517_), .A2(\asqrt[37] ), .A3(new_n7160_), .A4(new_n7165_), .ZN(new_n7579_));
  XOR2_X1    g07387(.A1(new_n7579_), .A2(new_n7578_), .Z(new_n7580_));
  NAND2_X1   g07388(.A1(new_n7580_), .A2(new_n4645_), .ZN(new_n7581_));
  AOI21_X1   g07389(.A1(new_n7577_), .A2(\asqrt[37] ), .B(new_n7581_), .ZN(new_n7582_));
  NOR2_X1    g07390(.A1(new_n7582_), .A2(new_n7575_), .ZN(new_n7583_));
  AOI21_X1   g07391(.A1(new_n7568_), .A2(new_n7573_), .B(new_n7576_), .ZN(new_n7584_));
  AOI21_X1   g07392(.A1(new_n7576_), .A2(new_n7568_), .B(new_n4973_), .ZN(new_n7585_));
  OAI21_X1   g07393(.A1(new_n7584_), .A2(new_n7585_), .B(\asqrt[38] ), .ZN(new_n7586_));
  NOR4_X1    g07394(.A1(new_n7517_), .A2(\asqrt[38] ), .A3(new_n7168_), .A4(new_n7365_), .ZN(new_n7587_));
  AOI21_X1   g07395(.A1(new_n7578_), .A2(new_n7164_), .B(new_n4645_), .ZN(new_n7588_));
  NOR2_X1    g07396(.A1(new_n7587_), .A2(new_n7588_), .ZN(new_n7589_));
  NAND2_X1   g07397(.A1(new_n7589_), .A2(new_n4330_), .ZN(new_n7590_));
  INV_X1     g07398(.I(new_n7590_), .ZN(new_n7591_));
  NAND2_X1   g07399(.A1(new_n7586_), .A2(new_n7591_), .ZN(new_n7592_));
  NAND2_X1   g07400(.A1(new_n7592_), .A2(new_n7583_), .ZN(new_n7593_));
  AOI22_X1   g07401(.A1(new_n7577_), .A2(\asqrt[37] ), .B1(new_n7574_), .B2(new_n7565_), .ZN(new_n7594_));
  OAI22_X1   g07402(.A1(new_n7594_), .A2(new_n4645_), .B1(new_n7582_), .B2(new_n7575_), .ZN(new_n7595_));
  NAND2_X1   g07403(.A1(new_n7179_), .A2(\asqrt[39] ), .ZN(new_n7596_));
  NOR4_X1    g07404(.A1(new_n7517_), .A2(\asqrt[39] ), .A3(new_n7174_), .A4(new_n7179_), .ZN(new_n7597_));
  XOR2_X1    g07405(.A1(new_n7597_), .A2(new_n7596_), .Z(new_n7598_));
  NAND2_X1   g07406(.A1(new_n7598_), .A2(new_n4018_), .ZN(new_n7599_));
  AOI21_X1   g07407(.A1(new_n7595_), .A2(\asqrt[39] ), .B(new_n7599_), .ZN(new_n7600_));
  NOR2_X1    g07408(.A1(new_n7600_), .A2(new_n7593_), .ZN(new_n7601_));
  AOI22_X1   g07409(.A1(new_n7595_), .A2(\asqrt[39] ), .B1(new_n7592_), .B2(new_n7583_), .ZN(new_n7602_));
  NOR4_X1    g07410(.A1(new_n7517_), .A2(\asqrt[40] ), .A3(new_n7181_), .A4(new_n7372_), .ZN(new_n7603_));
  AOI21_X1   g07411(.A1(new_n7596_), .A2(new_n7178_), .B(new_n4018_), .ZN(new_n7604_));
  NOR2_X1    g07412(.A1(new_n7603_), .A2(new_n7604_), .ZN(new_n7605_));
  NAND2_X1   g07413(.A1(new_n7605_), .A2(new_n3760_), .ZN(new_n7606_));
  INV_X1     g07414(.I(new_n7606_), .ZN(new_n7607_));
  OAI21_X1   g07415(.A1(new_n7602_), .A2(new_n4018_), .B(new_n7607_), .ZN(new_n7608_));
  NAND2_X1   g07416(.A1(new_n7608_), .A2(new_n7601_), .ZN(new_n7609_));
  OAI22_X1   g07417(.A1(new_n7602_), .A2(new_n4018_), .B1(new_n7600_), .B2(new_n7593_), .ZN(new_n7610_));
  NAND2_X1   g07418(.A1(new_n7192_), .A2(\asqrt[41] ), .ZN(new_n7611_));
  NOR4_X1    g07419(.A1(new_n7517_), .A2(\asqrt[41] ), .A3(new_n7187_), .A4(new_n7192_), .ZN(new_n7612_));
  XOR2_X1    g07420(.A1(new_n7612_), .A2(new_n7611_), .Z(new_n7613_));
  NAND2_X1   g07421(.A1(new_n7613_), .A2(new_n3481_), .ZN(new_n7614_));
  AOI21_X1   g07422(.A1(new_n7610_), .A2(\asqrt[41] ), .B(new_n7614_), .ZN(new_n7615_));
  NOR2_X1    g07423(.A1(new_n7615_), .A2(new_n7609_), .ZN(new_n7616_));
  AOI22_X1   g07424(.A1(new_n7610_), .A2(\asqrt[41] ), .B1(new_n7608_), .B2(new_n7601_), .ZN(new_n7617_));
  NAND2_X1   g07425(.A1(new_n7379_), .A2(\asqrt[42] ), .ZN(new_n7618_));
  NOR4_X1    g07426(.A1(new_n7517_), .A2(\asqrt[42] ), .A3(new_n7195_), .A4(new_n7379_), .ZN(new_n7619_));
  XOR2_X1    g07427(.A1(new_n7619_), .A2(new_n7618_), .Z(new_n7620_));
  NAND2_X1   g07428(.A1(new_n7620_), .A2(new_n3208_), .ZN(new_n7621_));
  INV_X1     g07429(.I(new_n7621_), .ZN(new_n7622_));
  OAI21_X1   g07430(.A1(new_n7617_), .A2(new_n3481_), .B(new_n7622_), .ZN(new_n7623_));
  NAND2_X1   g07431(.A1(new_n7623_), .A2(new_n7616_), .ZN(new_n7624_));
  OAI22_X1   g07432(.A1(new_n7617_), .A2(new_n3481_), .B1(new_n7615_), .B2(new_n7609_), .ZN(new_n7625_));
  NOR4_X1    g07433(.A1(new_n7517_), .A2(\asqrt[43] ), .A3(new_n7202_), .A4(new_n7207_), .ZN(new_n7626_));
  AOI21_X1   g07434(.A1(new_n7618_), .A2(new_n7378_), .B(new_n3208_), .ZN(new_n7627_));
  NOR2_X1    g07435(.A1(new_n7626_), .A2(new_n7627_), .ZN(new_n7628_));
  NAND2_X1   g07436(.A1(new_n7628_), .A2(new_n2941_), .ZN(new_n7629_));
  AOI21_X1   g07437(.A1(new_n7625_), .A2(\asqrt[43] ), .B(new_n7629_), .ZN(new_n7630_));
  NOR2_X1    g07438(.A1(new_n7630_), .A2(new_n7624_), .ZN(new_n7631_));
  AOI22_X1   g07439(.A1(new_n7625_), .A2(\asqrt[43] ), .B1(new_n7623_), .B2(new_n7616_), .ZN(new_n7632_));
  NAND2_X1   g07440(.A1(new_n7386_), .A2(\asqrt[44] ), .ZN(new_n7633_));
  NOR4_X1    g07441(.A1(new_n7517_), .A2(\asqrt[44] ), .A3(new_n7210_), .A4(new_n7386_), .ZN(new_n7634_));
  XOR2_X1    g07442(.A1(new_n7634_), .A2(new_n7633_), .Z(new_n7635_));
  NAND2_X1   g07443(.A1(new_n7635_), .A2(new_n2728_), .ZN(new_n7636_));
  INV_X1     g07444(.I(new_n7636_), .ZN(new_n7637_));
  OAI21_X1   g07445(.A1(new_n7632_), .A2(new_n2941_), .B(new_n7637_), .ZN(new_n7638_));
  NAND2_X1   g07446(.A1(new_n7638_), .A2(new_n7631_), .ZN(new_n7639_));
  OAI22_X1   g07447(.A1(new_n7632_), .A2(new_n2941_), .B1(new_n7630_), .B2(new_n7624_), .ZN(new_n7640_));
  NOR4_X1    g07448(.A1(new_n7517_), .A2(\asqrt[45] ), .A3(new_n7217_), .A4(new_n7222_), .ZN(new_n7641_));
  AOI21_X1   g07449(.A1(new_n7633_), .A2(new_n7385_), .B(new_n2728_), .ZN(new_n7642_));
  NOR2_X1    g07450(.A1(new_n7641_), .A2(new_n7642_), .ZN(new_n7643_));
  NAND2_X1   g07451(.A1(new_n7643_), .A2(new_n2488_), .ZN(new_n7644_));
  AOI21_X1   g07452(.A1(new_n7640_), .A2(\asqrt[45] ), .B(new_n7644_), .ZN(new_n7645_));
  NOR2_X1    g07453(.A1(new_n7645_), .A2(new_n7639_), .ZN(new_n7646_));
  AOI22_X1   g07454(.A1(new_n7640_), .A2(\asqrt[45] ), .B1(new_n7638_), .B2(new_n7631_), .ZN(new_n7647_));
  NAND2_X1   g07455(.A1(new_n7393_), .A2(\asqrt[46] ), .ZN(new_n7648_));
  NOR4_X1    g07456(.A1(new_n7517_), .A2(\asqrt[46] ), .A3(new_n7225_), .A4(new_n7393_), .ZN(new_n7649_));
  XOR2_X1    g07457(.A1(new_n7649_), .A2(new_n7648_), .Z(new_n7650_));
  NAND2_X1   g07458(.A1(new_n7650_), .A2(new_n2253_), .ZN(new_n7651_));
  INV_X1     g07459(.I(new_n7651_), .ZN(new_n7652_));
  OAI21_X1   g07460(.A1(new_n7647_), .A2(new_n2488_), .B(new_n7652_), .ZN(new_n7653_));
  NAND2_X1   g07461(.A1(new_n7653_), .A2(new_n7646_), .ZN(new_n7654_));
  OAI22_X1   g07462(.A1(new_n7647_), .A2(new_n2488_), .B1(new_n7645_), .B2(new_n7639_), .ZN(new_n7655_));
  NOR4_X1    g07463(.A1(new_n7517_), .A2(\asqrt[47] ), .A3(new_n7232_), .A4(new_n7237_), .ZN(new_n7656_));
  AOI21_X1   g07464(.A1(new_n7648_), .A2(new_n7392_), .B(new_n2253_), .ZN(new_n7657_));
  NOR2_X1    g07465(.A1(new_n7656_), .A2(new_n7657_), .ZN(new_n7658_));
  NAND2_X1   g07466(.A1(new_n7658_), .A2(new_n2046_), .ZN(new_n7659_));
  AOI21_X1   g07467(.A1(new_n7655_), .A2(\asqrt[47] ), .B(new_n7659_), .ZN(new_n7660_));
  NOR2_X1    g07468(.A1(new_n7660_), .A2(new_n7654_), .ZN(new_n7661_));
  AOI22_X1   g07469(.A1(new_n7655_), .A2(\asqrt[47] ), .B1(new_n7653_), .B2(new_n7646_), .ZN(new_n7662_));
  NAND2_X1   g07470(.A1(new_n7400_), .A2(\asqrt[48] ), .ZN(new_n7663_));
  NOR4_X1    g07471(.A1(new_n7517_), .A2(\asqrt[48] ), .A3(new_n7240_), .A4(new_n7400_), .ZN(new_n7664_));
  XOR2_X1    g07472(.A1(new_n7664_), .A2(new_n7663_), .Z(new_n7665_));
  NAND2_X1   g07473(.A1(new_n7665_), .A2(new_n1854_), .ZN(new_n7666_));
  INV_X1     g07474(.I(new_n7666_), .ZN(new_n7667_));
  OAI21_X1   g07475(.A1(new_n7662_), .A2(new_n2046_), .B(new_n7667_), .ZN(new_n7668_));
  NAND2_X1   g07476(.A1(new_n7668_), .A2(new_n7661_), .ZN(new_n7669_));
  OAI22_X1   g07477(.A1(new_n7662_), .A2(new_n2046_), .B1(new_n7660_), .B2(new_n7654_), .ZN(new_n7670_));
  NOR4_X1    g07478(.A1(new_n7517_), .A2(\asqrt[49] ), .A3(new_n7247_), .A4(new_n7252_), .ZN(new_n7671_));
  AOI21_X1   g07479(.A1(new_n7663_), .A2(new_n7399_), .B(new_n1854_), .ZN(new_n7672_));
  NOR2_X1    g07480(.A1(new_n7671_), .A2(new_n7672_), .ZN(new_n7673_));
  NAND2_X1   g07481(.A1(new_n7673_), .A2(new_n1595_), .ZN(new_n7674_));
  AOI21_X1   g07482(.A1(new_n7670_), .A2(\asqrt[49] ), .B(new_n7674_), .ZN(new_n7675_));
  NOR2_X1    g07483(.A1(new_n7675_), .A2(new_n7669_), .ZN(new_n7676_));
  AOI22_X1   g07484(.A1(new_n7670_), .A2(\asqrt[49] ), .B1(new_n7668_), .B2(new_n7661_), .ZN(new_n7677_));
  NAND2_X1   g07485(.A1(new_n7407_), .A2(\asqrt[50] ), .ZN(new_n7678_));
  NOR4_X1    g07486(.A1(new_n7517_), .A2(\asqrt[50] ), .A3(new_n7255_), .A4(new_n7407_), .ZN(new_n7679_));
  XOR2_X1    g07487(.A1(new_n7679_), .A2(new_n7678_), .Z(new_n7680_));
  NAND2_X1   g07488(.A1(new_n7680_), .A2(new_n1436_), .ZN(new_n7681_));
  INV_X1     g07489(.I(new_n7681_), .ZN(new_n7682_));
  OAI21_X1   g07490(.A1(new_n7677_), .A2(new_n1595_), .B(new_n7682_), .ZN(new_n7683_));
  NAND2_X1   g07491(.A1(new_n7683_), .A2(new_n7676_), .ZN(new_n7684_));
  OAI22_X1   g07492(.A1(new_n7677_), .A2(new_n1595_), .B1(new_n7675_), .B2(new_n7669_), .ZN(new_n7685_));
  NAND2_X1   g07493(.A1(new_n7267_), .A2(\asqrt[51] ), .ZN(new_n7686_));
  NOR4_X1    g07494(.A1(new_n7517_), .A2(\asqrt[51] ), .A3(new_n7262_), .A4(new_n7267_), .ZN(new_n7687_));
  XOR2_X1    g07495(.A1(new_n7687_), .A2(new_n7686_), .Z(new_n7688_));
  NAND2_X1   g07496(.A1(new_n7688_), .A2(new_n1260_), .ZN(new_n7689_));
  AOI21_X1   g07497(.A1(new_n7685_), .A2(\asqrt[51] ), .B(new_n7689_), .ZN(new_n7690_));
  NOR2_X1    g07498(.A1(new_n7690_), .A2(new_n7684_), .ZN(new_n7691_));
  AOI22_X1   g07499(.A1(new_n7685_), .A2(\asqrt[51] ), .B1(new_n7683_), .B2(new_n7676_), .ZN(new_n7692_));
  NOR4_X1    g07500(.A1(new_n7517_), .A2(\asqrt[52] ), .A3(new_n7270_), .A4(new_n7414_), .ZN(new_n7693_));
  AOI21_X1   g07501(.A1(new_n7686_), .A2(new_n7266_), .B(new_n1260_), .ZN(new_n7694_));
  NOR2_X1    g07502(.A1(new_n7693_), .A2(new_n7694_), .ZN(new_n7695_));
  NAND2_X1   g07503(.A1(new_n7695_), .A2(new_n1096_), .ZN(new_n7696_));
  INV_X1     g07504(.I(new_n7696_), .ZN(new_n7697_));
  OAI21_X1   g07505(.A1(new_n7692_), .A2(new_n1260_), .B(new_n7697_), .ZN(new_n7698_));
  NAND2_X1   g07506(.A1(new_n7698_), .A2(new_n7691_), .ZN(new_n7699_));
  OAI22_X1   g07507(.A1(new_n7692_), .A2(new_n1260_), .B1(new_n7690_), .B2(new_n7684_), .ZN(new_n7700_));
  NAND2_X1   g07508(.A1(new_n7282_), .A2(\asqrt[53] ), .ZN(new_n7701_));
  NOR4_X1    g07509(.A1(new_n7517_), .A2(\asqrt[53] ), .A3(new_n7277_), .A4(new_n7282_), .ZN(new_n7702_));
  XOR2_X1    g07510(.A1(new_n7702_), .A2(new_n7701_), .Z(new_n7703_));
  NAND2_X1   g07511(.A1(new_n7703_), .A2(new_n970_), .ZN(new_n7704_));
  AOI21_X1   g07512(.A1(new_n7700_), .A2(\asqrt[53] ), .B(new_n7704_), .ZN(new_n7705_));
  NOR2_X1    g07513(.A1(new_n7705_), .A2(new_n7699_), .ZN(new_n7706_));
  AOI22_X1   g07514(.A1(new_n7700_), .A2(\asqrt[53] ), .B1(new_n7698_), .B2(new_n7691_), .ZN(new_n7707_));
  NOR4_X1    g07515(.A1(new_n7517_), .A2(\asqrt[54] ), .A3(new_n7284_), .A4(new_n7421_), .ZN(new_n7708_));
  AOI21_X1   g07516(.A1(new_n7701_), .A2(new_n7281_), .B(new_n970_), .ZN(new_n7709_));
  NOR2_X1    g07517(.A1(new_n7708_), .A2(new_n7709_), .ZN(new_n7710_));
  NAND2_X1   g07518(.A1(new_n7710_), .A2(new_n825_), .ZN(new_n7711_));
  INV_X1     g07519(.I(new_n7711_), .ZN(new_n7712_));
  OAI21_X1   g07520(.A1(new_n7707_), .A2(new_n970_), .B(new_n7712_), .ZN(new_n7713_));
  NAND2_X1   g07521(.A1(new_n7713_), .A2(new_n7706_), .ZN(new_n7714_));
  OAI22_X1   g07522(.A1(new_n7707_), .A2(new_n970_), .B1(new_n7705_), .B2(new_n7699_), .ZN(new_n7715_));
  NAND2_X1   g07523(.A1(new_n7295_), .A2(\asqrt[55] ), .ZN(new_n7716_));
  NOR4_X1    g07524(.A1(new_n7517_), .A2(\asqrt[55] ), .A3(new_n7290_), .A4(new_n7295_), .ZN(new_n7717_));
  XOR2_X1    g07525(.A1(new_n7717_), .A2(new_n7716_), .Z(new_n7718_));
  NAND2_X1   g07526(.A1(new_n7718_), .A2(new_n724_), .ZN(new_n7719_));
  AOI21_X1   g07527(.A1(new_n7715_), .A2(\asqrt[55] ), .B(new_n7719_), .ZN(new_n7720_));
  NOR2_X1    g07528(.A1(new_n7720_), .A2(new_n7714_), .ZN(new_n7721_));
  AOI22_X1   g07529(.A1(new_n7715_), .A2(\asqrt[55] ), .B1(new_n7713_), .B2(new_n7706_), .ZN(new_n7722_));
  NAND2_X1   g07530(.A1(new_n7428_), .A2(\asqrt[56] ), .ZN(new_n7723_));
  NOR4_X1    g07531(.A1(new_n7517_), .A2(\asqrt[56] ), .A3(new_n7297_), .A4(new_n7428_), .ZN(new_n7724_));
  XOR2_X1    g07532(.A1(new_n7724_), .A2(new_n7723_), .Z(new_n7725_));
  NAND2_X1   g07533(.A1(new_n7725_), .A2(new_n587_), .ZN(new_n7726_));
  INV_X1     g07534(.I(new_n7726_), .ZN(new_n7727_));
  OAI21_X1   g07535(.A1(new_n7722_), .A2(new_n724_), .B(new_n7727_), .ZN(new_n7728_));
  NAND2_X1   g07536(.A1(new_n7728_), .A2(new_n7721_), .ZN(new_n7729_));
  NOR2_X1    g07537(.A1(new_n7722_), .A2(new_n724_), .ZN(new_n7730_));
  OAI21_X1   g07538(.A1(new_n7730_), .A2(new_n7721_), .B(\asqrt[57] ), .ZN(new_n7731_));
  NOR4_X1    g07539(.A1(new_n7517_), .A2(\asqrt[57] ), .A3(new_n7303_), .A4(new_n7308_), .ZN(new_n7732_));
  XOR2_X1    g07540(.A1(new_n7732_), .A2(new_n7457_), .Z(new_n7733_));
  NAND2_X1   g07541(.A1(new_n7733_), .A2(new_n504_), .ZN(new_n7734_));
  INV_X1     g07542(.I(new_n7734_), .ZN(new_n7735_));
  AOI21_X1   g07543(.A1(new_n7731_), .A2(new_n7735_), .B(new_n7729_), .ZN(new_n7736_));
  OAI22_X1   g07544(.A1(new_n7722_), .A2(new_n724_), .B1(new_n7720_), .B2(new_n7714_), .ZN(new_n7737_));
  AOI22_X1   g07545(.A1(new_n7737_), .A2(\asqrt[57] ), .B1(new_n7728_), .B2(new_n7721_), .ZN(new_n7738_));
  NOR4_X1    g07546(.A1(new_n7517_), .A2(\asqrt[58] ), .A3(new_n7310_), .A4(new_n7435_), .ZN(new_n7739_));
  XOR2_X1    g07547(.A1(new_n7739_), .A2(new_n7481_), .Z(new_n7740_));
  NAND2_X1   g07548(.A1(new_n7740_), .A2(new_n376_), .ZN(new_n7741_));
  INV_X1     g07549(.I(new_n7741_), .ZN(new_n7742_));
  OAI21_X1   g07550(.A1(new_n7738_), .A2(new_n504_), .B(new_n7742_), .ZN(new_n7743_));
  NAND2_X1   g07551(.A1(new_n7743_), .A2(new_n7736_), .ZN(new_n7744_));
  AOI21_X1   g07552(.A1(new_n7731_), .A2(new_n7729_), .B(new_n504_), .ZN(new_n7745_));
  OAI21_X1   g07553(.A1(new_n7736_), .A2(new_n7745_), .B(\asqrt[59] ), .ZN(new_n7746_));
  NOR4_X1    g07554(.A1(new_n7517_), .A2(\asqrt[59] ), .A3(new_n7316_), .A4(new_n7321_), .ZN(new_n7747_));
  XOR2_X1    g07555(.A1(new_n7747_), .A2(new_n7459_), .Z(new_n7748_));
  AND2_X2    g07556(.A1(new_n7748_), .A2(new_n275_), .Z(new_n7749_));
  AOI21_X1   g07557(.A1(new_n7746_), .A2(new_n7749_), .B(new_n7744_), .ZN(new_n7750_));
  INV_X1     g07558(.I(new_n7547_), .ZN(new_n7751_));
  OAI21_X1   g07559(.A1(new_n7549_), .A2(new_n6365_), .B(new_n7751_), .ZN(new_n7752_));
  AOI22_X1   g07560(.A1(new_n7550_), .A2(\asqrt[34] ), .B1(new_n7752_), .B2(new_n7540_), .ZN(new_n7753_));
  INV_X1     g07561(.I(new_n7563_), .ZN(new_n7754_));
  OAI21_X1   g07562(.A1(new_n7753_), .A2(new_n5626_), .B(new_n7754_), .ZN(new_n7755_));
  OAI22_X1   g07563(.A1(new_n7753_), .A2(new_n5626_), .B1(new_n7556_), .B2(new_n7548_), .ZN(new_n7756_));
  AOI22_X1   g07564(.A1(new_n7756_), .A2(\asqrt[36] ), .B1(new_n7755_), .B2(new_n7567_), .ZN(new_n7757_));
  INV_X1     g07565(.I(new_n7581_), .ZN(new_n7758_));
  OAI21_X1   g07566(.A1(new_n7757_), .A2(new_n4973_), .B(new_n7758_), .ZN(new_n7759_));
  NAND2_X1   g07567(.A1(new_n7759_), .A2(new_n7584_), .ZN(new_n7760_));
  AOI21_X1   g07568(.A1(new_n7756_), .A2(\asqrt[36] ), .B(new_n7572_), .ZN(new_n7761_));
  OAI22_X1   g07569(.A1(new_n7757_), .A2(new_n4973_), .B1(new_n7761_), .B2(new_n7576_), .ZN(new_n7762_));
  AOI21_X1   g07570(.A1(new_n7762_), .A2(\asqrt[38] ), .B(new_n7590_), .ZN(new_n7763_));
  NOR2_X1    g07571(.A1(new_n7763_), .A2(new_n7760_), .ZN(new_n7764_));
  AOI22_X1   g07572(.A1(new_n7762_), .A2(\asqrt[38] ), .B1(new_n7759_), .B2(new_n7584_), .ZN(new_n7765_));
  INV_X1     g07573(.I(new_n7599_), .ZN(new_n7766_));
  OAI21_X1   g07574(.A1(new_n7765_), .A2(new_n4330_), .B(new_n7766_), .ZN(new_n7767_));
  NAND2_X1   g07575(.A1(new_n7767_), .A2(new_n7764_), .ZN(new_n7768_));
  OAI22_X1   g07576(.A1(new_n7765_), .A2(new_n4330_), .B1(new_n7763_), .B2(new_n7760_), .ZN(new_n7769_));
  AOI21_X1   g07577(.A1(new_n7769_), .A2(\asqrt[40] ), .B(new_n7606_), .ZN(new_n7770_));
  NOR2_X1    g07578(.A1(new_n7770_), .A2(new_n7768_), .ZN(new_n7771_));
  AOI22_X1   g07579(.A1(new_n7769_), .A2(\asqrt[40] ), .B1(new_n7767_), .B2(new_n7764_), .ZN(new_n7772_));
  INV_X1     g07580(.I(new_n7614_), .ZN(new_n7773_));
  OAI21_X1   g07581(.A1(new_n7772_), .A2(new_n3760_), .B(new_n7773_), .ZN(new_n7774_));
  NAND2_X1   g07582(.A1(new_n7774_), .A2(new_n7771_), .ZN(new_n7775_));
  OAI22_X1   g07583(.A1(new_n7772_), .A2(new_n3760_), .B1(new_n7770_), .B2(new_n7768_), .ZN(new_n7776_));
  AOI21_X1   g07584(.A1(new_n7776_), .A2(\asqrt[42] ), .B(new_n7621_), .ZN(new_n7777_));
  NOR2_X1    g07585(.A1(new_n7777_), .A2(new_n7775_), .ZN(new_n7778_));
  AOI22_X1   g07586(.A1(new_n7776_), .A2(\asqrt[42] ), .B1(new_n7774_), .B2(new_n7771_), .ZN(new_n7779_));
  INV_X1     g07587(.I(new_n7629_), .ZN(new_n7780_));
  OAI21_X1   g07588(.A1(new_n7779_), .A2(new_n3208_), .B(new_n7780_), .ZN(new_n7781_));
  NAND2_X1   g07589(.A1(new_n7781_), .A2(new_n7778_), .ZN(new_n7782_));
  OAI22_X1   g07590(.A1(new_n7779_), .A2(new_n3208_), .B1(new_n7777_), .B2(new_n7775_), .ZN(new_n7783_));
  AOI21_X1   g07591(.A1(new_n7783_), .A2(\asqrt[44] ), .B(new_n7636_), .ZN(new_n7784_));
  NOR2_X1    g07592(.A1(new_n7784_), .A2(new_n7782_), .ZN(new_n7785_));
  AOI22_X1   g07593(.A1(new_n7783_), .A2(\asqrt[44] ), .B1(new_n7781_), .B2(new_n7778_), .ZN(new_n7786_));
  INV_X1     g07594(.I(new_n7644_), .ZN(new_n7787_));
  OAI21_X1   g07595(.A1(new_n7786_), .A2(new_n2728_), .B(new_n7787_), .ZN(new_n7788_));
  NAND2_X1   g07596(.A1(new_n7788_), .A2(new_n7785_), .ZN(new_n7789_));
  OAI22_X1   g07597(.A1(new_n7786_), .A2(new_n2728_), .B1(new_n7784_), .B2(new_n7782_), .ZN(new_n7790_));
  AOI21_X1   g07598(.A1(new_n7790_), .A2(\asqrt[46] ), .B(new_n7651_), .ZN(new_n7791_));
  NOR2_X1    g07599(.A1(new_n7791_), .A2(new_n7789_), .ZN(new_n7792_));
  AOI22_X1   g07600(.A1(new_n7790_), .A2(\asqrt[46] ), .B1(new_n7788_), .B2(new_n7785_), .ZN(new_n7793_));
  INV_X1     g07601(.I(new_n7659_), .ZN(new_n7794_));
  OAI21_X1   g07602(.A1(new_n7793_), .A2(new_n2253_), .B(new_n7794_), .ZN(new_n7795_));
  NAND2_X1   g07603(.A1(new_n7795_), .A2(new_n7792_), .ZN(new_n7796_));
  OAI22_X1   g07604(.A1(new_n7793_), .A2(new_n2253_), .B1(new_n7791_), .B2(new_n7789_), .ZN(new_n7797_));
  AOI21_X1   g07605(.A1(new_n7797_), .A2(\asqrt[48] ), .B(new_n7666_), .ZN(new_n7798_));
  NOR2_X1    g07606(.A1(new_n7798_), .A2(new_n7796_), .ZN(new_n7799_));
  AOI22_X1   g07607(.A1(new_n7797_), .A2(\asqrt[48] ), .B1(new_n7795_), .B2(new_n7792_), .ZN(new_n7800_));
  INV_X1     g07608(.I(new_n7674_), .ZN(new_n7801_));
  OAI21_X1   g07609(.A1(new_n7800_), .A2(new_n1854_), .B(new_n7801_), .ZN(new_n7802_));
  NAND2_X1   g07610(.A1(new_n7802_), .A2(new_n7799_), .ZN(new_n7803_));
  OAI22_X1   g07611(.A1(new_n7800_), .A2(new_n1854_), .B1(new_n7798_), .B2(new_n7796_), .ZN(new_n7804_));
  AOI21_X1   g07612(.A1(new_n7804_), .A2(\asqrt[50] ), .B(new_n7681_), .ZN(new_n7805_));
  NOR2_X1    g07613(.A1(new_n7805_), .A2(new_n7803_), .ZN(new_n7806_));
  AOI22_X1   g07614(.A1(new_n7804_), .A2(\asqrt[50] ), .B1(new_n7802_), .B2(new_n7799_), .ZN(new_n7807_));
  INV_X1     g07615(.I(new_n7689_), .ZN(new_n7808_));
  OAI21_X1   g07616(.A1(new_n7807_), .A2(new_n1436_), .B(new_n7808_), .ZN(new_n7809_));
  NAND2_X1   g07617(.A1(new_n7809_), .A2(new_n7806_), .ZN(new_n7810_));
  OAI22_X1   g07618(.A1(new_n7807_), .A2(new_n1436_), .B1(new_n7805_), .B2(new_n7803_), .ZN(new_n7811_));
  AOI21_X1   g07619(.A1(new_n7811_), .A2(\asqrt[52] ), .B(new_n7696_), .ZN(new_n7812_));
  NOR2_X1    g07620(.A1(new_n7812_), .A2(new_n7810_), .ZN(new_n7813_));
  AOI22_X1   g07621(.A1(new_n7811_), .A2(\asqrt[52] ), .B1(new_n7809_), .B2(new_n7806_), .ZN(new_n7814_));
  INV_X1     g07622(.I(new_n7704_), .ZN(new_n7815_));
  OAI21_X1   g07623(.A1(new_n7814_), .A2(new_n1096_), .B(new_n7815_), .ZN(new_n7816_));
  NAND2_X1   g07624(.A1(new_n7816_), .A2(new_n7813_), .ZN(new_n7817_));
  OAI22_X1   g07625(.A1(new_n7814_), .A2(new_n1096_), .B1(new_n7812_), .B2(new_n7810_), .ZN(new_n7818_));
  AOI21_X1   g07626(.A1(new_n7818_), .A2(\asqrt[54] ), .B(new_n7711_), .ZN(new_n7819_));
  NOR2_X1    g07627(.A1(new_n7819_), .A2(new_n7817_), .ZN(new_n7820_));
  AOI22_X1   g07628(.A1(new_n7818_), .A2(\asqrt[54] ), .B1(new_n7816_), .B2(new_n7813_), .ZN(new_n7821_));
  INV_X1     g07629(.I(new_n7719_), .ZN(new_n7822_));
  OAI21_X1   g07630(.A1(new_n7821_), .A2(new_n825_), .B(new_n7822_), .ZN(new_n7823_));
  NAND2_X1   g07631(.A1(new_n7823_), .A2(new_n7820_), .ZN(new_n7824_));
  OAI22_X1   g07632(.A1(new_n7821_), .A2(new_n825_), .B1(new_n7819_), .B2(new_n7817_), .ZN(new_n7825_));
  AOI21_X1   g07633(.A1(new_n7825_), .A2(\asqrt[56] ), .B(new_n7726_), .ZN(new_n7826_));
  NOR2_X1    g07634(.A1(new_n7826_), .A2(new_n7824_), .ZN(new_n7827_));
  AOI22_X1   g07635(.A1(new_n7825_), .A2(\asqrt[56] ), .B1(new_n7823_), .B2(new_n7820_), .ZN(new_n7828_));
  OAI21_X1   g07636(.A1(new_n7828_), .A2(new_n587_), .B(new_n7735_), .ZN(new_n7829_));
  NAND2_X1   g07637(.A1(new_n7829_), .A2(new_n7827_), .ZN(new_n7830_));
  NAND2_X1   g07638(.A1(new_n7818_), .A2(\asqrt[54] ), .ZN(new_n7831_));
  AOI21_X1   g07639(.A1(new_n7831_), .A2(new_n7817_), .B(new_n825_), .ZN(new_n7832_));
  OAI21_X1   g07640(.A1(new_n7820_), .A2(new_n7832_), .B(\asqrt[56] ), .ZN(new_n7833_));
  AOI21_X1   g07641(.A1(new_n7824_), .A2(new_n7833_), .B(new_n587_), .ZN(new_n7834_));
  OAI21_X1   g07642(.A1(new_n7827_), .A2(new_n7834_), .B(\asqrt[58] ), .ZN(new_n7835_));
  NAND2_X1   g07643(.A1(new_n7830_), .A2(new_n7835_), .ZN(new_n7836_));
  AOI22_X1   g07644(.A1(new_n7836_), .A2(\asqrt[59] ), .B1(new_n7743_), .B2(new_n7736_), .ZN(new_n7837_));
  NOR4_X1    g07645(.A1(new_n7517_), .A2(\asqrt[60] ), .A3(new_n7323_), .A4(new_n7442_), .ZN(new_n7838_));
  XOR2_X1    g07646(.A1(new_n7838_), .A2(new_n7483_), .Z(new_n7839_));
  NAND2_X1   g07647(.A1(new_n7839_), .A2(new_n229_), .ZN(new_n7840_));
  INV_X1     g07648(.I(new_n7840_), .ZN(new_n7841_));
  OAI21_X1   g07649(.A1(new_n7837_), .A2(new_n275_), .B(new_n7841_), .ZN(new_n7842_));
  OAI22_X1   g07650(.A1(new_n7828_), .A2(new_n587_), .B1(new_n7826_), .B2(new_n7824_), .ZN(new_n7843_));
  AOI21_X1   g07651(.A1(new_n7843_), .A2(\asqrt[58] ), .B(new_n7741_), .ZN(new_n7844_));
  NOR2_X1    g07652(.A1(new_n7844_), .A2(new_n7830_), .ZN(new_n7845_));
  AOI22_X1   g07653(.A1(new_n7843_), .A2(\asqrt[58] ), .B1(new_n7829_), .B2(new_n7827_), .ZN(new_n7846_));
  OAI21_X1   g07654(.A1(new_n7846_), .A2(new_n376_), .B(new_n7749_), .ZN(new_n7847_));
  NAND2_X1   g07655(.A1(new_n7847_), .A2(new_n7845_), .ZN(new_n7848_));
  AOI21_X1   g07656(.A1(new_n7830_), .A2(new_n7835_), .B(new_n376_), .ZN(new_n7849_));
  OAI21_X1   g07657(.A1(new_n7845_), .A2(new_n7849_), .B(\asqrt[60] ), .ZN(new_n7850_));
  AOI21_X1   g07658(.A1(new_n7848_), .A2(new_n7850_), .B(new_n229_), .ZN(new_n7851_));
  INV_X1     g07659(.I(new_n7487_), .ZN(new_n7852_));
  NOR2_X1    g07660(.A1(new_n7852_), .A2(\asqrt[62] ), .ZN(new_n7853_));
  INV_X1     g07661(.I(new_n7853_), .ZN(new_n7854_));
  NAND4_X1   g07662(.A1(new_n7851_), .A2(new_n7750_), .A3(new_n7842_), .A4(new_n7854_), .ZN(new_n7855_));
  NAND3_X1   g07663(.A1(new_n7517_), .A2(new_n7453_), .A3(new_n7505_), .ZN(new_n7856_));
  AOI21_X1   g07664(.A1(new_n7856_), .A2(new_n7465_), .B(\asqrt[63] ), .ZN(new_n7857_));
  NAND3_X1   g07665(.A1(new_n7855_), .A2(new_n7489_), .A3(new_n7857_), .ZN(new_n7858_));
  OAI22_X1   g07666(.A1(new_n7846_), .A2(new_n376_), .B1(new_n7844_), .B2(new_n7830_), .ZN(new_n7859_));
  AOI21_X1   g07667(.A1(new_n7859_), .A2(\asqrt[60] ), .B(new_n7840_), .ZN(new_n7860_));
  AOI22_X1   g07668(.A1(new_n7859_), .A2(\asqrt[60] ), .B1(new_n7847_), .B2(new_n7845_), .ZN(new_n7861_));
  OAI22_X1   g07669(.A1(new_n7861_), .A2(new_n229_), .B1(new_n7860_), .B2(new_n7848_), .ZN(new_n7862_));
  NOR4_X1    g07670(.A1(new_n7862_), .A2(\asqrt[62] ), .A3(new_n7479_), .A4(new_n7487_), .ZN(new_n7863_));
  AOI21_X1   g07671(.A1(new_n7480_), .A2(new_n7858_), .B(new_n7863_), .ZN(new_n7864_));
  INV_X1     g07672(.I(\a[56] ), .ZN(new_n7865_));
  OAI21_X1   g07673(.A1(new_n7454_), .A2(new_n7465_), .B(\asqrt[30] ), .ZN(new_n7866_));
  XOR2_X1    g07674(.A1(new_n7465_), .A2(\asqrt[63] ), .Z(new_n7867_));
  NAND2_X1   g07675(.A1(new_n7866_), .A2(new_n7867_), .ZN(new_n7868_));
  INV_X1     g07676(.I(new_n7868_), .ZN(new_n7869_));
  NAND3_X1   g07677(.A1(new_n7511_), .A2(new_n7447_), .A3(new_n7454_), .ZN(new_n7870_));
  INV_X1     g07678(.I(new_n7870_), .ZN(new_n7871_));
  NOR2_X1    g07679(.A1(new_n7869_), .A2(new_n7871_), .ZN(new_n7872_));
  NOR2_X1    g07680(.A1(\a[54] ), .A2(\a[55] ), .ZN(new_n7873_));
  INV_X1     g07681(.I(new_n7873_), .ZN(new_n7874_));
  NOR3_X1    g07682(.A1(new_n7872_), .A2(new_n7865_), .A3(new_n7874_), .ZN(new_n7875_));
  NAND2_X1   g07683(.A1(new_n7864_), .A2(new_n7875_), .ZN(new_n7876_));
  XOR2_X1    g07684(.A1(new_n7876_), .A2(\a[57] ), .Z(new_n7877_));
  INV_X1     g07685(.I(\a[57] ), .ZN(new_n7878_));
  NAND2_X1   g07686(.A1(new_n7842_), .A2(new_n7750_), .ZN(new_n7879_));
  NAND2_X1   g07687(.A1(new_n7851_), .A2(new_n7854_), .ZN(new_n7880_));
  OAI21_X1   g07688(.A1(new_n7880_), .A2(new_n7879_), .B(new_n7489_), .ZN(new_n7881_));
  INV_X1     g07689(.I(new_n7857_), .ZN(new_n7882_));
  OAI21_X1   g07690(.A1(new_n7881_), .A2(new_n7882_), .B(new_n7480_), .ZN(new_n7883_));
  NAND2_X1   g07691(.A1(new_n7863_), .A2(new_n7869_), .ZN(new_n7884_));
  NOR2_X1    g07692(.A1(new_n7884_), .A2(new_n7883_), .ZN(new_n7885_));
  NAND3_X1   g07693(.A1(new_n7885_), .A2(new_n7480_), .A3(new_n7870_), .ZN(new_n7886_));
  NAND2_X1   g07694(.A1(new_n7848_), .A2(new_n7850_), .ZN(new_n7887_));
  AOI22_X1   g07695(.A1(new_n7887_), .A2(\asqrt[61] ), .B1(new_n7842_), .B2(new_n7750_), .ZN(new_n7888_));
  NOR2_X1    g07696(.A1(new_n7888_), .A2(new_n196_), .ZN(new_n7889_));
  AOI21_X1   g07697(.A1(new_n7744_), .A2(new_n7746_), .B(new_n275_), .ZN(new_n7890_));
  OAI21_X1   g07698(.A1(new_n7750_), .A2(new_n7890_), .B(\asqrt[61] ), .ZN(new_n7891_));
  NAND4_X1   g07699(.A1(new_n7879_), .A2(new_n196_), .A3(new_n7891_), .A4(new_n7852_), .ZN(new_n7892_));
  INV_X1     g07700(.I(new_n7892_), .ZN(new_n7893_));
  NOR3_X1    g07701(.A1(new_n7884_), .A2(new_n7883_), .A3(new_n7870_), .ZN(\asqrt[29] ));
  NAND3_X1   g07702(.A1(\asqrt[29] ), .A2(new_n7889_), .A3(new_n7893_), .ZN(new_n7895_));
  OAI21_X1   g07703(.A1(new_n7862_), .A2(\asqrt[62] ), .B(new_n7487_), .ZN(new_n7896_));
  OAI21_X1   g07704(.A1(\asqrt[29] ), .A2(new_n7896_), .B(new_n7889_), .ZN(new_n7897_));
  NAND2_X1   g07705(.A1(new_n7897_), .A2(new_n7895_), .ZN(new_n7898_));
  INV_X1     g07706(.I(new_n7898_), .ZN(new_n7899_));
  NOR3_X1    g07707(.A1(new_n7887_), .A2(\asqrt[61] ), .A3(new_n7839_), .ZN(new_n7900_));
  NAND2_X1   g07708(.A1(\asqrt[29] ), .A2(new_n7900_), .ZN(new_n7901_));
  XOR2_X1    g07709(.A1(new_n7901_), .A2(new_n7851_), .Z(new_n7902_));
  NOR2_X1    g07710(.A1(new_n7902_), .A2(new_n196_), .ZN(new_n7903_));
  INV_X1     g07711(.I(new_n7903_), .ZN(new_n7904_));
  INV_X1     g07712(.I(\a[58] ), .ZN(new_n7905_));
  NOR2_X1    g07713(.A1(\a[56] ), .A2(\a[57] ), .ZN(new_n7906_));
  INV_X1     g07714(.I(new_n7906_), .ZN(new_n7907_));
  NOR2_X1    g07715(.A1(new_n7907_), .A2(new_n7905_), .ZN(new_n7908_));
  NAND4_X1   g07716(.A1(new_n7469_), .A2(new_n7505_), .A3(new_n7519_), .A4(new_n7908_), .ZN(new_n7909_));
  XOR2_X1    g07717(.A1(new_n7909_), .A2(\a[59] ), .Z(new_n7910_));
  INV_X1     g07718(.I(\a[59] ), .ZN(new_n7911_));
  NOR4_X1    g07719(.A1(new_n7884_), .A2(new_n7883_), .A3(new_n7911_), .A4(new_n7870_), .ZN(new_n7912_));
  NOR2_X1    g07720(.A1(new_n7910_), .A2(\a[58] ), .ZN(new_n7913_));
  OAI21_X1   g07721(.A1(new_n7912_), .A2(new_n7913_), .B(new_n7910_), .ZN(new_n7914_));
  INV_X1     g07722(.I(new_n7910_), .ZN(new_n7915_));
  NOR2_X1    g07723(.A1(new_n7860_), .A2(new_n7848_), .ZN(new_n7916_));
  NOR3_X1    g07724(.A1(new_n7861_), .A2(new_n229_), .A3(new_n7853_), .ZN(new_n7917_));
  AOI21_X1   g07725(.A1(new_n7917_), .A2(new_n7916_), .B(new_n7488_), .ZN(new_n7918_));
  AOI21_X1   g07726(.A1(new_n7918_), .A2(new_n7857_), .B(new_n7479_), .ZN(new_n7919_));
  AOI21_X1   g07727(.A1(new_n7862_), .A2(\asqrt[62] ), .B(new_n7480_), .ZN(new_n7920_));
  NOR3_X1    g07728(.A1(new_n7920_), .A2(new_n7892_), .A3(new_n7868_), .ZN(new_n7921_));
  NAND4_X1   g07729(.A1(new_n7921_), .A2(\a[59] ), .A3(new_n7919_), .A4(new_n7871_), .ZN(new_n7922_));
  NAND3_X1   g07730(.A1(new_n7922_), .A2(\a[58] ), .A3(new_n7915_), .ZN(new_n7923_));
  NAND2_X1   g07731(.A1(new_n7914_), .A2(new_n7923_), .ZN(new_n7924_));
  NAND2_X1   g07732(.A1(new_n7503_), .A2(new_n7467_), .ZN(new_n7925_));
  NAND4_X1   g07733(.A1(new_n7507_), .A2(new_n7501_), .A3(new_n7454_), .A4(new_n7925_), .ZN(new_n7926_));
  NOR2_X1    g07734(.A1(new_n7517_), .A2(new_n7905_), .ZN(new_n7927_));
  XOR2_X1    g07735(.A1(new_n7927_), .A2(new_n7926_), .Z(new_n7928_));
  NOR2_X1    g07736(.A1(new_n7928_), .A2(new_n7907_), .ZN(new_n7929_));
  INV_X1     g07737(.I(new_n7929_), .ZN(new_n7930_));
  NAND3_X1   g07738(.A1(new_n7921_), .A2(new_n7919_), .A3(new_n7871_), .ZN(new_n7931_));
  NOR4_X1    g07739(.A1(new_n7891_), .A2(new_n7848_), .A3(new_n7860_), .A4(new_n7853_), .ZN(new_n7932_));
  NOR3_X1    g07740(.A1(new_n7932_), .A2(new_n7488_), .A3(new_n7882_), .ZN(new_n7933_));
  NAND4_X1   g07741(.A1(new_n7888_), .A2(new_n196_), .A3(new_n7480_), .A4(new_n7852_), .ZN(new_n7934_));
  OAI21_X1   g07742(.A1(new_n7933_), .A2(new_n7479_), .B(new_n7934_), .ZN(new_n7935_));
  NAND2_X1   g07743(.A1(new_n7872_), .A2(\asqrt[30] ), .ZN(new_n7936_));
  OAI21_X1   g07744(.A1(new_n7935_), .A2(new_n7936_), .B(new_n7490_), .ZN(new_n7937_));
  NAND3_X1   g07745(.A1(new_n7937_), .A2(new_n7491_), .A3(new_n7931_), .ZN(new_n7938_));
  INV_X1     g07746(.I(new_n7936_), .ZN(new_n7939_));
  AOI21_X1   g07747(.A1(new_n7864_), .A2(new_n7939_), .B(\a[60] ), .ZN(new_n7940_));
  OAI21_X1   g07748(.A1(new_n7940_), .A2(new_n7492_), .B(\asqrt[29] ), .ZN(new_n7941_));
  NAND4_X1   g07749(.A1(new_n7938_), .A2(new_n7941_), .A3(new_n7110_), .A4(new_n7930_), .ZN(new_n7942_));
  NAND2_X1   g07750(.A1(new_n7942_), .A2(new_n7924_), .ZN(new_n7943_));
  NAND3_X1   g07751(.A1(new_n7914_), .A2(new_n7923_), .A3(new_n7930_), .ZN(new_n7944_));
  AOI21_X1   g07752(.A1(\asqrt[30] ), .A2(new_n7490_), .B(\a[61] ), .ZN(new_n7945_));
  NOR2_X1    g07753(.A1(new_n7508_), .A2(\a[60] ), .ZN(new_n7946_));
  AOI21_X1   g07754(.A1(\asqrt[30] ), .A2(\a[60] ), .B(new_n7494_), .ZN(new_n7947_));
  OAI21_X1   g07755(.A1(new_n7945_), .A2(new_n7946_), .B(new_n7947_), .ZN(new_n7948_));
  INV_X1     g07756(.I(new_n7948_), .ZN(new_n7949_));
  NAND3_X1   g07757(.A1(\asqrt[29] ), .A2(new_n7516_), .A3(new_n7949_), .ZN(new_n7950_));
  OAI21_X1   g07758(.A1(new_n7931_), .A2(new_n7948_), .B(new_n7515_), .ZN(new_n7951_));
  NAND3_X1   g07759(.A1(new_n7950_), .A2(new_n7951_), .A3(new_n6708_), .ZN(new_n7952_));
  AOI21_X1   g07760(.A1(new_n7944_), .A2(\asqrt[31] ), .B(new_n7952_), .ZN(new_n7953_));
  NOR2_X1    g07761(.A1(new_n7943_), .A2(new_n7953_), .ZN(new_n7954_));
  AOI22_X1   g07762(.A1(new_n7942_), .A2(new_n7924_), .B1(\asqrt[31] ), .B2(new_n7944_), .ZN(new_n7955_));
  INV_X1     g07763(.I(new_n7498_), .ZN(new_n7956_));
  AOI21_X1   g07764(.A1(new_n7508_), .A2(new_n7956_), .B(new_n7500_), .ZN(new_n7957_));
  INV_X1     g07765(.I(new_n7509_), .ZN(new_n7958_));
  NOR3_X1    g07766(.A1(new_n7958_), .A2(new_n7957_), .A3(new_n7515_), .ZN(new_n7959_));
  AOI21_X1   g07767(.A1(new_n7527_), .A2(new_n7523_), .B(\asqrt[32] ), .ZN(new_n7960_));
  AND4_X2    g07768(.A1(new_n7959_), .A2(\asqrt[29] ), .A3(new_n7541_), .A4(new_n7960_), .Z(new_n7961_));
  NOR2_X1    g07769(.A1(new_n7959_), .A2(new_n6708_), .ZN(new_n7962_));
  NOR3_X1    g07770(.A1(new_n7961_), .A2(\asqrt[33] ), .A3(new_n7962_), .ZN(new_n7963_));
  OAI21_X1   g07771(.A1(new_n7955_), .A2(new_n6708_), .B(new_n7963_), .ZN(new_n7964_));
  NAND2_X1   g07772(.A1(new_n7964_), .A2(new_n7954_), .ZN(new_n7965_));
  OAI22_X1   g07773(.A1(new_n7955_), .A2(new_n6708_), .B1(new_n7943_), .B2(new_n7953_), .ZN(new_n7966_));
  NAND2_X1   g07774(.A1(new_n7535_), .A2(new_n7537_), .ZN(new_n7967_));
  NAND4_X1   g07775(.A1(\asqrt[29] ), .A2(new_n6365_), .A3(new_n7967_), .A4(new_n7549_), .ZN(new_n7968_));
  XOR2_X1    g07776(.A1(new_n7968_), .A2(new_n7542_), .Z(new_n7969_));
  NAND2_X1   g07777(.A1(new_n7969_), .A2(new_n5991_), .ZN(new_n7970_));
  AOI21_X1   g07778(.A1(new_n7966_), .A2(\asqrt[33] ), .B(new_n7970_), .ZN(new_n7971_));
  NOR2_X1    g07779(.A1(new_n7971_), .A2(new_n7965_), .ZN(new_n7972_));
  AOI22_X1   g07780(.A1(new_n7966_), .A2(\asqrt[33] ), .B1(new_n7964_), .B2(new_n7954_), .ZN(new_n7973_));
  NOR4_X1    g07781(.A1(new_n7931_), .A2(\asqrt[34] ), .A3(new_n7546_), .A4(new_n7550_), .ZN(new_n7974_));
  XOR2_X1    g07782(.A1(new_n7974_), .A2(new_n7557_), .Z(new_n7975_));
  NAND2_X1   g07783(.A1(new_n7975_), .A2(new_n5626_), .ZN(new_n7976_));
  INV_X1     g07784(.I(new_n7976_), .ZN(new_n7977_));
  OAI21_X1   g07785(.A1(new_n7973_), .A2(new_n5991_), .B(new_n7977_), .ZN(new_n7978_));
  NAND2_X1   g07786(.A1(new_n7978_), .A2(new_n7972_), .ZN(new_n7979_));
  OAI22_X1   g07787(.A1(new_n7973_), .A2(new_n5991_), .B1(new_n7971_), .B2(new_n7965_), .ZN(new_n7980_));
  NOR2_X1    g07788(.A1(new_n7554_), .A2(\asqrt[35] ), .ZN(new_n7981_));
  NAND3_X1   g07789(.A1(\asqrt[29] ), .A2(new_n7753_), .A3(new_n7981_), .ZN(new_n7982_));
  XOR2_X1    g07790(.A1(new_n7982_), .A2(new_n7558_), .Z(new_n7983_));
  NAND2_X1   g07791(.A1(new_n7983_), .A2(new_n5273_), .ZN(new_n7984_));
  AOI21_X1   g07792(.A1(new_n7980_), .A2(\asqrt[35] ), .B(new_n7984_), .ZN(new_n7985_));
  NOR2_X1    g07793(.A1(new_n7985_), .A2(new_n7979_), .ZN(new_n7986_));
  AOI22_X1   g07794(.A1(new_n7980_), .A2(\asqrt[35] ), .B1(new_n7978_), .B2(new_n7972_), .ZN(new_n7987_));
  NOR4_X1    g07795(.A1(new_n7931_), .A2(\asqrt[36] ), .A3(new_n7562_), .A4(new_n7756_), .ZN(new_n7988_));
  XOR2_X1    g07796(.A1(new_n7988_), .A2(new_n7568_), .Z(new_n7989_));
  NAND2_X1   g07797(.A1(new_n7989_), .A2(new_n4973_), .ZN(new_n7990_));
  INV_X1     g07798(.I(new_n7990_), .ZN(new_n7991_));
  OAI21_X1   g07799(.A1(new_n7987_), .A2(new_n5273_), .B(new_n7991_), .ZN(new_n7992_));
  NAND2_X1   g07800(.A1(new_n7992_), .A2(new_n7986_), .ZN(new_n7993_));
  OAI22_X1   g07801(.A1(new_n7987_), .A2(new_n5273_), .B1(new_n7985_), .B2(new_n7979_), .ZN(new_n7994_));
  NOR4_X1    g07802(.A1(new_n7931_), .A2(\asqrt[37] ), .A3(new_n7571_), .A4(new_n7577_), .ZN(new_n7995_));
  XNOR2_X1   g07803(.A1(new_n7995_), .A2(new_n7585_), .ZN(new_n7996_));
  NAND2_X1   g07804(.A1(new_n7996_), .A2(new_n4645_), .ZN(new_n7997_));
  AOI21_X1   g07805(.A1(new_n7994_), .A2(\asqrt[37] ), .B(new_n7997_), .ZN(new_n7998_));
  NOR2_X1    g07806(.A1(new_n7998_), .A2(new_n7993_), .ZN(new_n7999_));
  AOI22_X1   g07807(.A1(new_n7994_), .A2(\asqrt[37] ), .B1(new_n7992_), .B2(new_n7986_), .ZN(new_n8000_));
  NOR4_X1    g07808(.A1(new_n7931_), .A2(\asqrt[38] ), .A3(new_n7580_), .A4(new_n7762_), .ZN(new_n8001_));
  XOR2_X1    g07809(.A1(new_n8001_), .A2(new_n7586_), .Z(new_n8002_));
  NAND2_X1   g07810(.A1(new_n8002_), .A2(new_n4330_), .ZN(new_n8003_));
  INV_X1     g07811(.I(new_n8003_), .ZN(new_n8004_));
  OAI21_X1   g07812(.A1(new_n8000_), .A2(new_n4645_), .B(new_n8004_), .ZN(new_n8005_));
  NAND2_X1   g07813(.A1(new_n8005_), .A2(new_n7999_), .ZN(new_n8006_));
  OAI22_X1   g07814(.A1(new_n8000_), .A2(new_n4645_), .B1(new_n7998_), .B2(new_n7993_), .ZN(new_n8007_));
  NAND2_X1   g07815(.A1(new_n7595_), .A2(\asqrt[39] ), .ZN(new_n8008_));
  NOR4_X1    g07816(.A1(new_n7931_), .A2(\asqrt[39] ), .A3(new_n7589_), .A4(new_n7595_), .ZN(new_n8009_));
  XOR2_X1    g07817(.A1(new_n8009_), .A2(new_n8008_), .Z(new_n8010_));
  NAND2_X1   g07818(.A1(new_n8010_), .A2(new_n4018_), .ZN(new_n8011_));
  AOI21_X1   g07819(.A1(new_n8007_), .A2(\asqrt[39] ), .B(new_n8011_), .ZN(new_n8012_));
  NOR2_X1    g07820(.A1(new_n8012_), .A2(new_n8006_), .ZN(new_n8013_));
  AOI22_X1   g07821(.A1(new_n8007_), .A2(\asqrt[39] ), .B1(new_n8005_), .B2(new_n7999_), .ZN(new_n8014_));
  NOR4_X1    g07822(.A1(new_n7931_), .A2(\asqrt[40] ), .A3(new_n7598_), .A4(new_n7769_), .ZN(new_n8015_));
  AOI21_X1   g07823(.A1(new_n8008_), .A2(new_n7593_), .B(new_n4018_), .ZN(new_n8016_));
  NOR2_X1    g07824(.A1(new_n8015_), .A2(new_n8016_), .ZN(new_n8017_));
  NAND2_X1   g07825(.A1(new_n8017_), .A2(new_n3760_), .ZN(new_n8018_));
  INV_X1     g07826(.I(new_n8018_), .ZN(new_n8019_));
  OAI21_X1   g07827(.A1(new_n8014_), .A2(new_n4018_), .B(new_n8019_), .ZN(new_n8020_));
  NAND2_X1   g07828(.A1(new_n8020_), .A2(new_n8013_), .ZN(new_n8021_));
  OAI22_X1   g07829(.A1(new_n8014_), .A2(new_n4018_), .B1(new_n8012_), .B2(new_n8006_), .ZN(new_n8022_));
  NAND2_X1   g07830(.A1(new_n7610_), .A2(\asqrt[41] ), .ZN(new_n8023_));
  NOR4_X1    g07831(.A1(new_n7931_), .A2(\asqrt[41] ), .A3(new_n7605_), .A4(new_n7610_), .ZN(new_n8024_));
  XOR2_X1    g07832(.A1(new_n8024_), .A2(new_n8023_), .Z(new_n8025_));
  NAND2_X1   g07833(.A1(new_n8025_), .A2(new_n3481_), .ZN(new_n8026_));
  AOI21_X1   g07834(.A1(new_n8022_), .A2(\asqrt[41] ), .B(new_n8026_), .ZN(new_n8027_));
  NOR2_X1    g07835(.A1(new_n8027_), .A2(new_n8021_), .ZN(new_n8028_));
  AOI22_X1   g07836(.A1(new_n8022_), .A2(\asqrt[41] ), .B1(new_n8020_), .B2(new_n8013_), .ZN(new_n8029_));
  NOR4_X1    g07837(.A1(new_n7931_), .A2(\asqrt[42] ), .A3(new_n7613_), .A4(new_n7776_), .ZN(new_n8030_));
  AOI21_X1   g07838(.A1(new_n8023_), .A2(new_n7609_), .B(new_n3481_), .ZN(new_n8031_));
  NOR2_X1    g07839(.A1(new_n8030_), .A2(new_n8031_), .ZN(new_n8032_));
  NAND2_X1   g07840(.A1(new_n8032_), .A2(new_n3208_), .ZN(new_n8033_));
  INV_X1     g07841(.I(new_n8033_), .ZN(new_n8034_));
  OAI21_X1   g07842(.A1(new_n8029_), .A2(new_n3481_), .B(new_n8034_), .ZN(new_n8035_));
  NAND2_X1   g07843(.A1(new_n8035_), .A2(new_n8028_), .ZN(new_n8036_));
  OAI22_X1   g07844(.A1(new_n8029_), .A2(new_n3481_), .B1(new_n8027_), .B2(new_n8021_), .ZN(new_n8037_));
  NAND2_X1   g07845(.A1(new_n7625_), .A2(\asqrt[43] ), .ZN(new_n8038_));
  NOR4_X1    g07846(.A1(new_n7931_), .A2(\asqrt[43] ), .A3(new_n7620_), .A4(new_n7625_), .ZN(new_n8039_));
  XOR2_X1    g07847(.A1(new_n8039_), .A2(new_n8038_), .Z(new_n8040_));
  NAND2_X1   g07848(.A1(new_n8040_), .A2(new_n2941_), .ZN(new_n8041_));
  AOI21_X1   g07849(.A1(new_n8037_), .A2(\asqrt[43] ), .B(new_n8041_), .ZN(new_n8042_));
  NOR2_X1    g07850(.A1(new_n8042_), .A2(new_n8036_), .ZN(new_n8043_));
  AOI22_X1   g07851(.A1(new_n8037_), .A2(\asqrt[43] ), .B1(new_n8035_), .B2(new_n8028_), .ZN(new_n8044_));
  NOR4_X1    g07852(.A1(new_n7931_), .A2(\asqrt[44] ), .A3(new_n7628_), .A4(new_n7783_), .ZN(new_n8045_));
  AOI21_X1   g07853(.A1(new_n8038_), .A2(new_n7624_), .B(new_n2941_), .ZN(new_n8046_));
  NOR2_X1    g07854(.A1(new_n8045_), .A2(new_n8046_), .ZN(new_n8047_));
  NAND2_X1   g07855(.A1(new_n8047_), .A2(new_n2728_), .ZN(new_n8048_));
  INV_X1     g07856(.I(new_n8048_), .ZN(new_n8049_));
  OAI21_X1   g07857(.A1(new_n8044_), .A2(new_n2941_), .B(new_n8049_), .ZN(new_n8050_));
  NAND2_X1   g07858(.A1(new_n8050_), .A2(new_n8043_), .ZN(new_n8051_));
  OAI22_X1   g07859(.A1(new_n8044_), .A2(new_n2941_), .B1(new_n8042_), .B2(new_n8036_), .ZN(new_n8052_));
  NAND2_X1   g07860(.A1(new_n7640_), .A2(\asqrt[45] ), .ZN(new_n8053_));
  NOR4_X1    g07861(.A1(new_n7931_), .A2(\asqrt[45] ), .A3(new_n7635_), .A4(new_n7640_), .ZN(new_n8054_));
  XOR2_X1    g07862(.A1(new_n8054_), .A2(new_n8053_), .Z(new_n8055_));
  NAND2_X1   g07863(.A1(new_n8055_), .A2(new_n2488_), .ZN(new_n8056_));
  AOI21_X1   g07864(.A1(new_n8052_), .A2(\asqrt[45] ), .B(new_n8056_), .ZN(new_n8057_));
  NOR2_X1    g07865(.A1(new_n8057_), .A2(new_n8051_), .ZN(new_n8058_));
  AOI22_X1   g07866(.A1(new_n8052_), .A2(\asqrt[45] ), .B1(new_n8050_), .B2(new_n8043_), .ZN(new_n8059_));
  NOR4_X1    g07867(.A1(new_n7931_), .A2(\asqrt[46] ), .A3(new_n7643_), .A4(new_n7790_), .ZN(new_n8060_));
  AOI21_X1   g07868(.A1(new_n8053_), .A2(new_n7639_), .B(new_n2488_), .ZN(new_n8061_));
  NOR2_X1    g07869(.A1(new_n8060_), .A2(new_n8061_), .ZN(new_n8062_));
  NAND2_X1   g07870(.A1(new_n8062_), .A2(new_n2253_), .ZN(new_n8063_));
  INV_X1     g07871(.I(new_n8063_), .ZN(new_n8064_));
  OAI21_X1   g07872(.A1(new_n8059_), .A2(new_n2488_), .B(new_n8064_), .ZN(new_n8065_));
  NAND2_X1   g07873(.A1(new_n8065_), .A2(new_n8058_), .ZN(new_n8066_));
  OAI22_X1   g07874(.A1(new_n8059_), .A2(new_n2488_), .B1(new_n8057_), .B2(new_n8051_), .ZN(new_n8067_));
  NAND2_X1   g07875(.A1(new_n7655_), .A2(\asqrt[47] ), .ZN(new_n8068_));
  NOR4_X1    g07876(.A1(new_n7931_), .A2(\asqrt[47] ), .A3(new_n7650_), .A4(new_n7655_), .ZN(new_n8069_));
  XOR2_X1    g07877(.A1(new_n8069_), .A2(new_n8068_), .Z(new_n8070_));
  NAND2_X1   g07878(.A1(new_n8070_), .A2(new_n2046_), .ZN(new_n8071_));
  AOI21_X1   g07879(.A1(new_n8067_), .A2(\asqrt[47] ), .B(new_n8071_), .ZN(new_n8072_));
  NOR2_X1    g07880(.A1(new_n8072_), .A2(new_n8066_), .ZN(new_n8073_));
  AOI22_X1   g07881(.A1(new_n8067_), .A2(\asqrt[47] ), .B1(new_n8065_), .B2(new_n8058_), .ZN(new_n8074_));
  NOR4_X1    g07882(.A1(new_n7931_), .A2(\asqrt[48] ), .A3(new_n7658_), .A4(new_n7797_), .ZN(new_n8075_));
  AOI21_X1   g07883(.A1(new_n8068_), .A2(new_n7654_), .B(new_n2046_), .ZN(new_n8076_));
  NOR2_X1    g07884(.A1(new_n8075_), .A2(new_n8076_), .ZN(new_n8077_));
  NAND2_X1   g07885(.A1(new_n8077_), .A2(new_n1854_), .ZN(new_n8078_));
  INV_X1     g07886(.I(new_n8078_), .ZN(new_n8079_));
  OAI21_X1   g07887(.A1(new_n8074_), .A2(new_n2046_), .B(new_n8079_), .ZN(new_n8080_));
  NAND2_X1   g07888(.A1(new_n8080_), .A2(new_n8073_), .ZN(new_n8081_));
  OAI22_X1   g07889(.A1(new_n8074_), .A2(new_n2046_), .B1(new_n8072_), .B2(new_n8066_), .ZN(new_n8082_));
  NAND2_X1   g07890(.A1(new_n7670_), .A2(\asqrt[49] ), .ZN(new_n8083_));
  NOR4_X1    g07891(.A1(new_n7931_), .A2(\asqrt[49] ), .A3(new_n7665_), .A4(new_n7670_), .ZN(new_n8084_));
  XOR2_X1    g07892(.A1(new_n8084_), .A2(new_n8083_), .Z(new_n8085_));
  NAND2_X1   g07893(.A1(new_n8085_), .A2(new_n1595_), .ZN(new_n8086_));
  AOI21_X1   g07894(.A1(new_n8082_), .A2(\asqrt[49] ), .B(new_n8086_), .ZN(new_n8087_));
  NOR2_X1    g07895(.A1(new_n8087_), .A2(new_n8081_), .ZN(new_n8088_));
  AOI22_X1   g07896(.A1(new_n8082_), .A2(\asqrt[49] ), .B1(new_n8080_), .B2(new_n8073_), .ZN(new_n8089_));
  NAND2_X1   g07897(.A1(new_n7804_), .A2(\asqrt[50] ), .ZN(new_n8090_));
  NOR4_X1    g07898(.A1(new_n7931_), .A2(\asqrt[50] ), .A3(new_n7673_), .A4(new_n7804_), .ZN(new_n8091_));
  XOR2_X1    g07899(.A1(new_n8091_), .A2(new_n8090_), .Z(new_n8092_));
  NAND2_X1   g07900(.A1(new_n8092_), .A2(new_n1436_), .ZN(new_n8093_));
  INV_X1     g07901(.I(new_n8093_), .ZN(new_n8094_));
  OAI21_X1   g07902(.A1(new_n8089_), .A2(new_n1595_), .B(new_n8094_), .ZN(new_n8095_));
  NAND2_X1   g07903(.A1(new_n8095_), .A2(new_n8088_), .ZN(new_n8096_));
  OAI22_X1   g07904(.A1(new_n8089_), .A2(new_n1595_), .B1(new_n8087_), .B2(new_n8081_), .ZN(new_n8097_));
  NOR4_X1    g07905(.A1(new_n7931_), .A2(\asqrt[51] ), .A3(new_n7680_), .A4(new_n7685_), .ZN(new_n8098_));
  AOI21_X1   g07906(.A1(new_n8090_), .A2(new_n7803_), .B(new_n1436_), .ZN(new_n8099_));
  NOR2_X1    g07907(.A1(new_n8098_), .A2(new_n8099_), .ZN(new_n8100_));
  NAND2_X1   g07908(.A1(new_n8100_), .A2(new_n1260_), .ZN(new_n8101_));
  AOI21_X1   g07909(.A1(new_n8097_), .A2(\asqrt[51] ), .B(new_n8101_), .ZN(new_n8102_));
  NOR2_X1    g07910(.A1(new_n8102_), .A2(new_n8096_), .ZN(new_n8103_));
  AOI22_X1   g07911(.A1(new_n8097_), .A2(\asqrt[51] ), .B1(new_n8095_), .B2(new_n8088_), .ZN(new_n8104_));
  NAND2_X1   g07912(.A1(new_n7811_), .A2(\asqrt[52] ), .ZN(new_n8105_));
  NOR4_X1    g07913(.A1(new_n7931_), .A2(\asqrt[52] ), .A3(new_n7688_), .A4(new_n7811_), .ZN(new_n8106_));
  XOR2_X1    g07914(.A1(new_n8106_), .A2(new_n8105_), .Z(new_n8107_));
  NAND2_X1   g07915(.A1(new_n8107_), .A2(new_n1096_), .ZN(new_n8108_));
  INV_X1     g07916(.I(new_n8108_), .ZN(new_n8109_));
  OAI21_X1   g07917(.A1(new_n8104_), .A2(new_n1260_), .B(new_n8109_), .ZN(new_n8110_));
  NAND2_X1   g07918(.A1(new_n8110_), .A2(new_n8103_), .ZN(new_n8111_));
  OAI22_X1   g07919(.A1(new_n8104_), .A2(new_n1260_), .B1(new_n8102_), .B2(new_n8096_), .ZN(new_n8112_));
  NOR2_X1    g07920(.A1(new_n7814_), .A2(new_n1096_), .ZN(new_n8113_));
  NOR4_X1    g07921(.A1(new_n7931_), .A2(\asqrt[53] ), .A3(new_n7695_), .A4(new_n7700_), .ZN(new_n8114_));
  XNOR2_X1   g07922(.A1(new_n8114_), .A2(new_n8113_), .ZN(new_n8115_));
  NAND2_X1   g07923(.A1(new_n8115_), .A2(new_n970_), .ZN(new_n8116_));
  AOI21_X1   g07924(.A1(new_n8112_), .A2(\asqrt[53] ), .B(new_n8116_), .ZN(new_n8117_));
  NOR2_X1    g07925(.A1(new_n8117_), .A2(new_n8111_), .ZN(new_n8118_));
  AOI22_X1   g07926(.A1(new_n8112_), .A2(\asqrt[53] ), .B1(new_n8110_), .B2(new_n8103_), .ZN(new_n8119_));
  NOR4_X1    g07927(.A1(new_n7931_), .A2(\asqrt[54] ), .A3(new_n7703_), .A4(new_n7818_), .ZN(new_n8120_));
  XOR2_X1    g07928(.A1(new_n8120_), .A2(new_n7831_), .Z(new_n8121_));
  NAND2_X1   g07929(.A1(new_n8121_), .A2(new_n825_), .ZN(new_n8122_));
  INV_X1     g07930(.I(new_n8122_), .ZN(new_n8123_));
  OAI21_X1   g07931(.A1(new_n8119_), .A2(new_n970_), .B(new_n8123_), .ZN(new_n8124_));
  NAND2_X1   g07932(.A1(new_n8124_), .A2(new_n8118_), .ZN(new_n8125_));
  OAI22_X1   g07933(.A1(new_n8119_), .A2(new_n970_), .B1(new_n8117_), .B2(new_n8111_), .ZN(new_n8126_));
  NOR4_X1    g07934(.A1(new_n7931_), .A2(\asqrt[55] ), .A3(new_n7710_), .A4(new_n7715_), .ZN(new_n8127_));
  XNOR2_X1   g07935(.A1(new_n8127_), .A2(new_n7832_), .ZN(new_n8128_));
  NAND2_X1   g07936(.A1(new_n8128_), .A2(new_n724_), .ZN(new_n8129_));
  AOI21_X1   g07937(.A1(new_n8126_), .A2(\asqrt[55] ), .B(new_n8129_), .ZN(new_n8130_));
  NOR2_X1    g07938(.A1(new_n8130_), .A2(new_n8125_), .ZN(new_n8131_));
  AOI22_X1   g07939(.A1(new_n8126_), .A2(\asqrt[55] ), .B1(new_n8124_), .B2(new_n8118_), .ZN(new_n8132_));
  NOR4_X1    g07940(.A1(new_n7931_), .A2(\asqrt[56] ), .A3(new_n7718_), .A4(new_n7825_), .ZN(new_n8133_));
  XOR2_X1    g07941(.A1(new_n8133_), .A2(new_n7833_), .Z(new_n8134_));
  NAND2_X1   g07942(.A1(new_n8134_), .A2(new_n587_), .ZN(new_n8135_));
  INV_X1     g07943(.I(new_n8135_), .ZN(new_n8136_));
  OAI21_X1   g07944(.A1(new_n8132_), .A2(new_n724_), .B(new_n8136_), .ZN(new_n8137_));
  NAND2_X1   g07945(.A1(new_n8137_), .A2(new_n8131_), .ZN(new_n8138_));
  OAI22_X1   g07946(.A1(new_n8132_), .A2(new_n724_), .B1(new_n8130_), .B2(new_n8125_), .ZN(new_n8139_));
  NOR4_X1    g07947(.A1(new_n7931_), .A2(\asqrt[57] ), .A3(new_n7725_), .A4(new_n7737_), .ZN(new_n8140_));
  XOR2_X1    g07948(.A1(new_n8140_), .A2(new_n7731_), .Z(new_n8141_));
  NAND2_X1   g07949(.A1(new_n8141_), .A2(new_n504_), .ZN(new_n8142_));
  AOI21_X1   g07950(.A1(new_n8139_), .A2(\asqrt[57] ), .B(new_n8142_), .ZN(new_n8143_));
  NOR2_X1    g07951(.A1(new_n8143_), .A2(new_n8138_), .ZN(new_n8144_));
  AOI22_X1   g07952(.A1(new_n8139_), .A2(\asqrt[57] ), .B1(new_n8137_), .B2(new_n8131_), .ZN(new_n8145_));
  NOR4_X1    g07953(.A1(new_n7931_), .A2(\asqrt[58] ), .A3(new_n7733_), .A4(new_n7843_), .ZN(new_n8146_));
  XOR2_X1    g07954(.A1(new_n8146_), .A2(new_n7835_), .Z(new_n8147_));
  NAND2_X1   g07955(.A1(new_n8147_), .A2(new_n376_), .ZN(new_n8148_));
  INV_X1     g07956(.I(new_n8148_), .ZN(new_n8149_));
  OAI21_X1   g07957(.A1(new_n8145_), .A2(new_n504_), .B(new_n8149_), .ZN(new_n8150_));
  NAND2_X1   g07958(.A1(new_n8150_), .A2(new_n8144_), .ZN(new_n8151_));
  OAI22_X1   g07959(.A1(new_n8145_), .A2(new_n504_), .B1(new_n8143_), .B2(new_n8138_), .ZN(new_n8152_));
  NOR4_X1    g07960(.A1(new_n7931_), .A2(\asqrt[59] ), .A3(new_n7740_), .A4(new_n7836_), .ZN(new_n8153_));
  XOR2_X1    g07961(.A1(new_n8153_), .A2(new_n7746_), .Z(new_n8154_));
  NAND2_X1   g07962(.A1(new_n8154_), .A2(new_n275_), .ZN(new_n8155_));
  AOI21_X1   g07963(.A1(new_n8152_), .A2(\asqrt[59] ), .B(new_n8155_), .ZN(new_n8156_));
  NOR2_X1    g07964(.A1(new_n8156_), .A2(new_n8151_), .ZN(new_n8157_));
  AOI22_X1   g07965(.A1(new_n8152_), .A2(\asqrt[59] ), .B1(new_n8150_), .B2(new_n8144_), .ZN(new_n8158_));
  NOR4_X1    g07966(.A1(new_n7931_), .A2(\asqrt[60] ), .A3(new_n7748_), .A4(new_n7859_), .ZN(new_n8159_));
  XOR2_X1    g07967(.A1(new_n8159_), .A2(new_n7850_), .Z(new_n8160_));
  NAND2_X1   g07968(.A1(new_n8160_), .A2(new_n229_), .ZN(new_n8161_));
  INV_X1     g07969(.I(new_n8161_), .ZN(new_n8162_));
  OAI21_X1   g07970(.A1(new_n8158_), .A2(new_n275_), .B(new_n8162_), .ZN(new_n8163_));
  NAND2_X1   g07971(.A1(new_n8163_), .A2(new_n8157_), .ZN(new_n8164_));
  OAI22_X1   g07972(.A1(new_n8158_), .A2(new_n275_), .B1(new_n8156_), .B2(new_n8151_), .ZN(new_n8165_));
  INV_X1     g07973(.I(new_n7902_), .ZN(new_n8166_));
  NOR2_X1    g07974(.A1(new_n8166_), .A2(\asqrt[62] ), .ZN(new_n8167_));
  INV_X1     g07975(.I(new_n8167_), .ZN(new_n8168_));
  NAND3_X1   g07976(.A1(new_n8165_), .A2(\asqrt[61] ), .A3(new_n8168_), .ZN(new_n8169_));
  OAI21_X1   g07977(.A1(new_n8169_), .A2(new_n8164_), .B(new_n7904_), .ZN(new_n8170_));
  NAND3_X1   g07978(.A1(new_n7931_), .A2(new_n7479_), .A3(new_n7934_), .ZN(new_n8171_));
  AOI21_X1   g07979(.A1(new_n8171_), .A2(new_n7881_), .B(\asqrt[63] ), .ZN(new_n8172_));
  INV_X1     g07980(.I(new_n8172_), .ZN(new_n8173_));
  OAI21_X1   g07981(.A1(new_n8170_), .A2(new_n8173_), .B(new_n7899_), .ZN(new_n8174_));
  INV_X1     g07982(.I(new_n7913_), .ZN(new_n8175_));
  AOI21_X1   g07983(.A1(new_n7922_), .A2(new_n8175_), .B(new_n7915_), .ZN(new_n8176_));
  NOR3_X1    g07984(.A1(new_n7912_), .A2(new_n7905_), .A3(new_n7910_), .ZN(new_n8177_));
  NOR2_X1    g07985(.A1(new_n8177_), .A2(new_n8176_), .ZN(new_n8178_));
  NOR3_X1    g07986(.A1(new_n7940_), .A2(new_n7492_), .A3(\asqrt[29] ), .ZN(new_n8179_));
  AOI21_X1   g07987(.A1(new_n7937_), .A2(new_n7491_), .B(new_n7931_), .ZN(new_n8180_));
  NOR4_X1    g07988(.A1(new_n8180_), .A2(new_n8179_), .A3(\asqrt[31] ), .A4(new_n7929_), .ZN(new_n8181_));
  NOR2_X1    g07989(.A1(new_n8181_), .A2(new_n8178_), .ZN(new_n8182_));
  NOR3_X1    g07990(.A1(new_n8177_), .A2(new_n8176_), .A3(new_n7929_), .ZN(new_n8183_));
  NOR3_X1    g07991(.A1(new_n7931_), .A2(new_n7515_), .A3(new_n7948_), .ZN(new_n8184_));
  AOI21_X1   g07992(.A1(\asqrt[29] ), .A2(new_n7949_), .B(new_n7516_), .ZN(new_n8185_));
  NOR3_X1    g07993(.A1(new_n8185_), .A2(new_n8184_), .A3(\asqrt[32] ), .ZN(new_n8186_));
  OAI21_X1   g07994(.A1(new_n8183_), .A2(new_n7110_), .B(new_n8186_), .ZN(new_n8187_));
  NAND2_X1   g07995(.A1(new_n8182_), .A2(new_n8187_), .ZN(new_n8188_));
  OAI22_X1   g07996(.A1(new_n8181_), .A2(new_n8178_), .B1(new_n7110_), .B2(new_n8183_), .ZN(new_n8189_));
  INV_X1     g07997(.I(new_n7963_), .ZN(new_n8190_));
  AOI21_X1   g07998(.A1(new_n8189_), .A2(\asqrt[32] ), .B(new_n8190_), .ZN(new_n8191_));
  NOR2_X1    g07999(.A1(new_n8191_), .A2(new_n8188_), .ZN(new_n8192_));
  AOI22_X1   g08000(.A1(new_n8189_), .A2(\asqrt[32] ), .B1(new_n8182_), .B2(new_n8187_), .ZN(new_n8193_));
  INV_X1     g08001(.I(new_n7970_), .ZN(new_n8194_));
  OAI21_X1   g08002(.A1(new_n8193_), .A2(new_n6365_), .B(new_n8194_), .ZN(new_n8195_));
  NAND2_X1   g08003(.A1(new_n8195_), .A2(new_n8192_), .ZN(new_n8196_));
  OAI22_X1   g08004(.A1(new_n8193_), .A2(new_n6365_), .B1(new_n8191_), .B2(new_n8188_), .ZN(new_n8197_));
  AOI21_X1   g08005(.A1(new_n8197_), .A2(\asqrt[34] ), .B(new_n7976_), .ZN(new_n8198_));
  NOR2_X1    g08006(.A1(new_n8198_), .A2(new_n8196_), .ZN(new_n8199_));
  AOI22_X1   g08007(.A1(new_n8197_), .A2(\asqrt[34] ), .B1(new_n8195_), .B2(new_n8192_), .ZN(new_n8200_));
  INV_X1     g08008(.I(new_n7984_), .ZN(new_n8201_));
  OAI21_X1   g08009(.A1(new_n8200_), .A2(new_n5626_), .B(new_n8201_), .ZN(new_n8202_));
  NAND2_X1   g08010(.A1(new_n8202_), .A2(new_n8199_), .ZN(new_n8203_));
  OAI22_X1   g08011(.A1(new_n8200_), .A2(new_n5626_), .B1(new_n8198_), .B2(new_n8196_), .ZN(new_n8204_));
  AOI21_X1   g08012(.A1(new_n8204_), .A2(\asqrt[36] ), .B(new_n7990_), .ZN(new_n8205_));
  NOR2_X1    g08013(.A1(new_n8205_), .A2(new_n8203_), .ZN(new_n8206_));
  AOI22_X1   g08014(.A1(new_n8204_), .A2(\asqrt[36] ), .B1(new_n8202_), .B2(new_n8199_), .ZN(new_n8207_));
  INV_X1     g08015(.I(new_n7997_), .ZN(new_n8208_));
  OAI21_X1   g08016(.A1(new_n8207_), .A2(new_n4973_), .B(new_n8208_), .ZN(new_n8209_));
  NAND2_X1   g08017(.A1(new_n8209_), .A2(new_n8206_), .ZN(new_n8210_));
  OAI22_X1   g08018(.A1(new_n8207_), .A2(new_n4973_), .B1(new_n8205_), .B2(new_n8203_), .ZN(new_n8211_));
  AOI21_X1   g08019(.A1(new_n8211_), .A2(\asqrt[38] ), .B(new_n8003_), .ZN(new_n8212_));
  NOR2_X1    g08020(.A1(new_n8212_), .A2(new_n8210_), .ZN(new_n8213_));
  AOI22_X1   g08021(.A1(new_n8211_), .A2(\asqrt[38] ), .B1(new_n8209_), .B2(new_n8206_), .ZN(new_n8214_));
  INV_X1     g08022(.I(new_n8011_), .ZN(new_n8215_));
  OAI21_X1   g08023(.A1(new_n8214_), .A2(new_n4330_), .B(new_n8215_), .ZN(new_n8216_));
  NAND2_X1   g08024(.A1(new_n8216_), .A2(new_n8213_), .ZN(new_n8217_));
  OAI22_X1   g08025(.A1(new_n8214_), .A2(new_n4330_), .B1(new_n8212_), .B2(new_n8210_), .ZN(new_n8218_));
  AOI21_X1   g08026(.A1(new_n8218_), .A2(\asqrt[40] ), .B(new_n8018_), .ZN(new_n8219_));
  NOR2_X1    g08027(.A1(new_n8219_), .A2(new_n8217_), .ZN(new_n8220_));
  AOI22_X1   g08028(.A1(new_n8218_), .A2(\asqrt[40] ), .B1(new_n8216_), .B2(new_n8213_), .ZN(new_n8221_));
  INV_X1     g08029(.I(new_n8026_), .ZN(new_n8222_));
  OAI21_X1   g08030(.A1(new_n8221_), .A2(new_n3760_), .B(new_n8222_), .ZN(new_n8223_));
  NAND2_X1   g08031(.A1(new_n8223_), .A2(new_n8220_), .ZN(new_n8224_));
  OAI22_X1   g08032(.A1(new_n8221_), .A2(new_n3760_), .B1(new_n8219_), .B2(new_n8217_), .ZN(new_n8225_));
  AOI21_X1   g08033(.A1(new_n8225_), .A2(\asqrt[42] ), .B(new_n8033_), .ZN(new_n8226_));
  NOR2_X1    g08034(.A1(new_n8226_), .A2(new_n8224_), .ZN(new_n8227_));
  AOI22_X1   g08035(.A1(new_n8225_), .A2(\asqrt[42] ), .B1(new_n8223_), .B2(new_n8220_), .ZN(new_n8228_));
  INV_X1     g08036(.I(new_n8041_), .ZN(new_n8229_));
  OAI21_X1   g08037(.A1(new_n8228_), .A2(new_n3208_), .B(new_n8229_), .ZN(new_n8230_));
  NAND2_X1   g08038(.A1(new_n8230_), .A2(new_n8227_), .ZN(new_n8231_));
  OAI22_X1   g08039(.A1(new_n8228_), .A2(new_n3208_), .B1(new_n8226_), .B2(new_n8224_), .ZN(new_n8232_));
  AOI21_X1   g08040(.A1(new_n8232_), .A2(\asqrt[44] ), .B(new_n8048_), .ZN(new_n8233_));
  NOR2_X1    g08041(.A1(new_n8233_), .A2(new_n8231_), .ZN(new_n8234_));
  AOI22_X1   g08042(.A1(new_n8232_), .A2(\asqrt[44] ), .B1(new_n8230_), .B2(new_n8227_), .ZN(new_n8235_));
  INV_X1     g08043(.I(new_n8056_), .ZN(new_n8236_));
  OAI21_X1   g08044(.A1(new_n8235_), .A2(new_n2728_), .B(new_n8236_), .ZN(new_n8237_));
  NAND2_X1   g08045(.A1(new_n8237_), .A2(new_n8234_), .ZN(new_n8238_));
  OAI22_X1   g08046(.A1(new_n8235_), .A2(new_n2728_), .B1(new_n8233_), .B2(new_n8231_), .ZN(new_n8239_));
  AOI21_X1   g08047(.A1(new_n8239_), .A2(\asqrt[46] ), .B(new_n8063_), .ZN(new_n8240_));
  NOR2_X1    g08048(.A1(new_n8240_), .A2(new_n8238_), .ZN(new_n8241_));
  AOI22_X1   g08049(.A1(new_n8239_), .A2(\asqrt[46] ), .B1(new_n8237_), .B2(new_n8234_), .ZN(new_n8242_));
  INV_X1     g08050(.I(new_n8071_), .ZN(new_n8243_));
  OAI21_X1   g08051(.A1(new_n8242_), .A2(new_n2253_), .B(new_n8243_), .ZN(new_n8244_));
  NAND2_X1   g08052(.A1(new_n8244_), .A2(new_n8241_), .ZN(new_n8245_));
  OAI22_X1   g08053(.A1(new_n8242_), .A2(new_n2253_), .B1(new_n8240_), .B2(new_n8238_), .ZN(new_n8246_));
  AOI21_X1   g08054(.A1(new_n8246_), .A2(\asqrt[48] ), .B(new_n8078_), .ZN(new_n8247_));
  NOR2_X1    g08055(.A1(new_n8247_), .A2(new_n8245_), .ZN(new_n8248_));
  AOI22_X1   g08056(.A1(new_n8246_), .A2(\asqrt[48] ), .B1(new_n8244_), .B2(new_n8241_), .ZN(new_n8249_));
  INV_X1     g08057(.I(new_n8086_), .ZN(new_n8250_));
  OAI21_X1   g08058(.A1(new_n8249_), .A2(new_n1854_), .B(new_n8250_), .ZN(new_n8251_));
  NAND2_X1   g08059(.A1(new_n8251_), .A2(new_n8248_), .ZN(new_n8252_));
  OAI22_X1   g08060(.A1(new_n8249_), .A2(new_n1854_), .B1(new_n8247_), .B2(new_n8245_), .ZN(new_n8253_));
  AOI21_X1   g08061(.A1(new_n8253_), .A2(\asqrt[50] ), .B(new_n8093_), .ZN(new_n8254_));
  NOR2_X1    g08062(.A1(new_n8254_), .A2(new_n8252_), .ZN(new_n8255_));
  AOI22_X1   g08063(.A1(new_n8253_), .A2(\asqrt[50] ), .B1(new_n8251_), .B2(new_n8248_), .ZN(new_n8256_));
  INV_X1     g08064(.I(new_n8101_), .ZN(new_n8257_));
  OAI21_X1   g08065(.A1(new_n8256_), .A2(new_n1436_), .B(new_n8257_), .ZN(new_n8258_));
  NAND2_X1   g08066(.A1(new_n8258_), .A2(new_n8255_), .ZN(new_n8259_));
  OAI22_X1   g08067(.A1(new_n8256_), .A2(new_n1436_), .B1(new_n8254_), .B2(new_n8252_), .ZN(new_n8260_));
  AOI21_X1   g08068(.A1(new_n8260_), .A2(\asqrt[52] ), .B(new_n8108_), .ZN(new_n8261_));
  NOR2_X1    g08069(.A1(new_n8261_), .A2(new_n8259_), .ZN(new_n8262_));
  AOI22_X1   g08070(.A1(new_n8260_), .A2(\asqrt[52] ), .B1(new_n8258_), .B2(new_n8255_), .ZN(new_n8263_));
  INV_X1     g08071(.I(new_n8116_), .ZN(new_n8264_));
  OAI21_X1   g08072(.A1(new_n8263_), .A2(new_n1096_), .B(new_n8264_), .ZN(new_n8265_));
  NAND2_X1   g08073(.A1(new_n8265_), .A2(new_n8262_), .ZN(new_n8266_));
  OAI22_X1   g08074(.A1(new_n8263_), .A2(new_n1096_), .B1(new_n8261_), .B2(new_n8259_), .ZN(new_n8267_));
  AOI21_X1   g08075(.A1(new_n8267_), .A2(\asqrt[54] ), .B(new_n8122_), .ZN(new_n8268_));
  NOR2_X1    g08076(.A1(new_n8268_), .A2(new_n8266_), .ZN(new_n8269_));
  AOI22_X1   g08077(.A1(new_n8267_), .A2(\asqrt[54] ), .B1(new_n8265_), .B2(new_n8262_), .ZN(new_n8270_));
  INV_X1     g08078(.I(new_n8129_), .ZN(new_n8271_));
  OAI21_X1   g08079(.A1(new_n8270_), .A2(new_n825_), .B(new_n8271_), .ZN(new_n8272_));
  NAND2_X1   g08080(.A1(new_n8272_), .A2(new_n8269_), .ZN(new_n8273_));
  OAI22_X1   g08081(.A1(new_n8270_), .A2(new_n825_), .B1(new_n8268_), .B2(new_n8266_), .ZN(new_n8274_));
  AOI21_X1   g08082(.A1(new_n8274_), .A2(\asqrt[56] ), .B(new_n8135_), .ZN(new_n8275_));
  NOR2_X1    g08083(.A1(new_n8275_), .A2(new_n8273_), .ZN(new_n8276_));
  AOI22_X1   g08084(.A1(new_n8274_), .A2(\asqrt[56] ), .B1(new_n8272_), .B2(new_n8269_), .ZN(new_n8277_));
  INV_X1     g08085(.I(new_n8142_), .ZN(new_n8278_));
  OAI21_X1   g08086(.A1(new_n8277_), .A2(new_n587_), .B(new_n8278_), .ZN(new_n8279_));
  NAND2_X1   g08087(.A1(new_n8279_), .A2(new_n8276_), .ZN(new_n8280_));
  OAI22_X1   g08088(.A1(new_n8277_), .A2(new_n587_), .B1(new_n8275_), .B2(new_n8273_), .ZN(new_n8281_));
  AOI21_X1   g08089(.A1(new_n8281_), .A2(\asqrt[58] ), .B(new_n8148_), .ZN(new_n8282_));
  NOR2_X1    g08090(.A1(new_n8282_), .A2(new_n8280_), .ZN(new_n8283_));
  AOI22_X1   g08091(.A1(new_n8281_), .A2(\asqrt[58] ), .B1(new_n8279_), .B2(new_n8276_), .ZN(new_n8284_));
  INV_X1     g08092(.I(new_n8155_), .ZN(new_n8285_));
  OAI21_X1   g08093(.A1(new_n8284_), .A2(new_n376_), .B(new_n8285_), .ZN(new_n8286_));
  NAND2_X1   g08094(.A1(new_n8286_), .A2(new_n8283_), .ZN(new_n8287_));
  OAI22_X1   g08095(.A1(new_n8284_), .A2(new_n376_), .B1(new_n8282_), .B2(new_n8280_), .ZN(new_n8288_));
  AOI21_X1   g08096(.A1(new_n8288_), .A2(\asqrt[60] ), .B(new_n8161_), .ZN(new_n8289_));
  AOI22_X1   g08097(.A1(new_n8288_), .A2(\asqrt[60] ), .B1(new_n8286_), .B2(new_n8283_), .ZN(new_n8290_));
  OAI22_X1   g08098(.A1(new_n8290_), .A2(new_n229_), .B1(new_n8289_), .B2(new_n8287_), .ZN(new_n8291_));
  NOR4_X1    g08099(.A1(new_n8291_), .A2(\asqrt[62] ), .A3(new_n7898_), .A4(new_n7902_), .ZN(new_n8292_));
  NAND2_X1   g08100(.A1(new_n7918_), .A2(new_n7479_), .ZN(new_n8293_));
  XOR2_X1    g08101(.A1(new_n7918_), .A2(\asqrt[63] ), .Z(new_n8294_));
  AOI21_X1   g08102(.A1(\asqrt[29] ), .A2(new_n8293_), .B(new_n8294_), .ZN(new_n8295_));
  NAND2_X1   g08103(.A1(new_n8292_), .A2(new_n8295_), .ZN(new_n8296_));
  NOR4_X1    g08104(.A1(new_n8296_), .A2(new_n7878_), .A3(new_n7886_), .A4(new_n8174_), .ZN(new_n8297_));
  NOR2_X1    g08105(.A1(new_n7878_), .A2(\a[56] ), .ZN(new_n8298_));
  OAI21_X1   g08106(.A1(new_n8297_), .A2(new_n8298_), .B(new_n7877_), .ZN(new_n8299_));
  INV_X1     g08107(.I(new_n7877_), .ZN(new_n8300_));
  INV_X1     g08108(.I(new_n7886_), .ZN(new_n8301_));
  NOR2_X1    g08109(.A1(new_n8289_), .A2(new_n8287_), .ZN(new_n8302_));
  NOR3_X1    g08110(.A1(new_n8290_), .A2(new_n229_), .A3(new_n8167_), .ZN(new_n8303_));
  AOI21_X1   g08111(.A1(new_n8303_), .A2(new_n8302_), .B(new_n7903_), .ZN(new_n8304_));
  AOI21_X1   g08112(.A1(new_n8304_), .A2(new_n8172_), .B(new_n7898_), .ZN(new_n8305_));
  AOI22_X1   g08113(.A1(new_n8165_), .A2(\asqrt[61] ), .B1(new_n8163_), .B2(new_n8157_), .ZN(new_n8306_));
  NAND4_X1   g08114(.A1(new_n8306_), .A2(new_n196_), .A3(new_n7899_), .A4(new_n8166_), .ZN(new_n8307_));
  INV_X1     g08115(.I(new_n8295_), .ZN(new_n8308_));
  NOR2_X1    g08116(.A1(new_n8307_), .A2(new_n8308_), .ZN(new_n8309_));
  NAND4_X1   g08117(.A1(new_n8309_), .A2(new_n8305_), .A3(\a[57] ), .A4(new_n8301_), .ZN(new_n8310_));
  NAND3_X1   g08118(.A1(new_n8310_), .A2(\a[56] ), .A3(new_n8300_), .ZN(new_n8311_));
  NAND2_X1   g08119(.A1(new_n8299_), .A2(new_n8311_), .ZN(new_n8312_));
  NOR2_X1    g08120(.A1(new_n8296_), .A2(new_n8174_), .ZN(new_n8313_));
  NOR4_X1    g08121(.A1(new_n7884_), .A2(new_n7479_), .A3(new_n7933_), .A4(new_n7870_), .ZN(new_n8314_));
  NAND2_X1   g08122(.A1(\asqrt[29] ), .A2(\a[56] ), .ZN(new_n8315_));
  XOR2_X1    g08123(.A1(new_n8315_), .A2(new_n8314_), .Z(new_n8316_));
  NOR2_X1    g08124(.A1(new_n8316_), .A2(new_n7874_), .ZN(new_n8317_));
  INV_X1     g08125(.I(new_n8317_), .ZN(new_n8318_));
  NAND3_X1   g08126(.A1(new_n8309_), .A2(new_n8305_), .A3(new_n8301_), .ZN(new_n8319_));
  NAND2_X1   g08127(.A1(new_n8126_), .A2(\asqrt[55] ), .ZN(new_n8320_));
  AOI21_X1   g08128(.A1(new_n8320_), .A2(new_n8125_), .B(new_n724_), .ZN(new_n8321_));
  OAI21_X1   g08129(.A1(new_n8131_), .A2(new_n8321_), .B(\asqrt[57] ), .ZN(new_n8322_));
  AOI21_X1   g08130(.A1(new_n8138_), .A2(new_n8322_), .B(new_n504_), .ZN(new_n8323_));
  OAI21_X1   g08131(.A1(new_n8144_), .A2(new_n8323_), .B(\asqrt[59] ), .ZN(new_n8324_));
  AOI21_X1   g08132(.A1(new_n8151_), .A2(new_n8324_), .B(new_n275_), .ZN(new_n8325_));
  OAI21_X1   g08133(.A1(new_n8157_), .A2(new_n8325_), .B(\asqrt[61] ), .ZN(new_n8326_));
  NOR3_X1    g08134(.A1(new_n8164_), .A2(new_n8326_), .A3(new_n8167_), .ZN(new_n8327_));
  NOR3_X1    g08135(.A1(new_n8327_), .A2(new_n7903_), .A3(new_n8173_), .ZN(new_n8328_));
  OAI21_X1   g08136(.A1(new_n8328_), .A2(new_n7898_), .B(new_n8307_), .ZN(new_n8329_));
  NOR2_X1    g08137(.A1(new_n8301_), .A2(new_n8295_), .ZN(new_n8330_));
  NAND2_X1   g08138(.A1(new_n8330_), .A2(\asqrt[29] ), .ZN(new_n8331_));
  OAI21_X1   g08139(.A1(new_n8329_), .A2(new_n8331_), .B(new_n7905_), .ZN(new_n8332_));
  NAND3_X1   g08140(.A1(new_n8332_), .A2(new_n7906_), .A3(new_n8319_), .ZN(new_n8333_));
  NOR3_X1    g08141(.A1(new_n8296_), .A2(new_n7886_), .A3(new_n8174_), .ZN(\asqrt[28] ));
  NAND2_X1   g08142(.A1(new_n8274_), .A2(\asqrt[56] ), .ZN(new_n8335_));
  AOI21_X1   g08143(.A1(new_n8335_), .A2(new_n8273_), .B(new_n587_), .ZN(new_n8336_));
  OAI21_X1   g08144(.A1(new_n8276_), .A2(new_n8336_), .B(\asqrt[58] ), .ZN(new_n8337_));
  AOI21_X1   g08145(.A1(new_n8280_), .A2(new_n8337_), .B(new_n376_), .ZN(new_n8338_));
  OAI21_X1   g08146(.A1(new_n8283_), .A2(new_n8338_), .B(\asqrt[60] ), .ZN(new_n8339_));
  AOI21_X1   g08147(.A1(new_n8287_), .A2(new_n8339_), .B(new_n229_), .ZN(new_n8340_));
  NAND4_X1   g08148(.A1(new_n8340_), .A2(new_n8157_), .A3(new_n8163_), .A4(new_n8168_), .ZN(new_n8341_));
  NAND3_X1   g08149(.A1(new_n8341_), .A2(new_n7904_), .A3(new_n8172_), .ZN(new_n8342_));
  AOI21_X1   g08150(.A1(new_n7899_), .A2(new_n8342_), .B(new_n8292_), .ZN(new_n8343_));
  INV_X1     g08151(.I(new_n8331_), .ZN(new_n8344_));
  AOI21_X1   g08152(.A1(new_n8343_), .A2(new_n8344_), .B(\a[58] ), .ZN(new_n8345_));
  OAI21_X1   g08153(.A1(new_n8345_), .A2(new_n7907_), .B(\asqrt[28] ), .ZN(new_n8346_));
  NAND4_X1   g08154(.A1(new_n8346_), .A2(new_n8333_), .A3(new_n7517_), .A4(new_n8318_), .ZN(new_n8347_));
  NAND2_X1   g08155(.A1(new_n8347_), .A2(new_n8312_), .ZN(new_n8348_));
  NAND3_X1   g08156(.A1(new_n8299_), .A2(new_n8311_), .A3(new_n8318_), .ZN(new_n8349_));
  AOI21_X1   g08157(.A1(\asqrt[29] ), .A2(new_n7905_), .B(\a[59] ), .ZN(new_n8350_));
  NOR2_X1    g08158(.A1(new_n7922_), .A2(\a[58] ), .ZN(new_n8351_));
  AOI21_X1   g08159(.A1(\asqrt[29] ), .A2(\a[58] ), .B(new_n7909_), .ZN(new_n8352_));
  OAI21_X1   g08160(.A1(new_n8351_), .A2(new_n8350_), .B(new_n8352_), .ZN(new_n8353_));
  INV_X1     g08161(.I(new_n8353_), .ZN(new_n8354_));
  NAND3_X1   g08162(.A1(\asqrt[28] ), .A2(new_n7930_), .A3(new_n8354_), .ZN(new_n8355_));
  OAI21_X1   g08163(.A1(new_n8319_), .A2(new_n8353_), .B(new_n7929_), .ZN(new_n8356_));
  NAND3_X1   g08164(.A1(new_n8355_), .A2(new_n8356_), .A3(new_n7110_), .ZN(new_n8357_));
  AOI21_X1   g08165(.A1(new_n8349_), .A2(\asqrt[30] ), .B(new_n8357_), .ZN(new_n8358_));
  NOR2_X1    g08166(.A1(new_n8348_), .A2(new_n8358_), .ZN(new_n8359_));
  NAND2_X1   g08167(.A1(new_n8349_), .A2(\asqrt[30] ), .ZN(new_n8360_));
  AOI21_X1   g08168(.A1(new_n8348_), .A2(new_n8360_), .B(new_n7110_), .ZN(new_n8361_));
  NAND2_X1   g08169(.A1(new_n7944_), .A2(\asqrt[31] ), .ZN(new_n8362_));
  NAND2_X1   g08170(.A1(new_n7938_), .A2(new_n7941_), .ZN(new_n8363_));
  NAND3_X1   g08171(.A1(new_n8363_), .A2(new_n8183_), .A3(new_n7110_), .ZN(new_n8364_));
  NOR2_X1    g08172(.A1(new_n8319_), .A2(new_n8364_), .ZN(new_n8365_));
  AND2_X2    g08173(.A1(new_n8365_), .A2(new_n8362_), .Z(new_n8366_));
  NOR2_X1    g08174(.A1(new_n8365_), .A2(new_n8362_), .ZN(new_n8367_));
  NOR3_X1    g08175(.A1(new_n8366_), .A2(\asqrt[32] ), .A3(new_n8367_), .ZN(new_n8368_));
  INV_X1     g08176(.I(new_n8368_), .ZN(new_n8369_));
  OAI21_X1   g08177(.A1(new_n8361_), .A2(new_n8369_), .B(new_n8359_), .ZN(new_n8370_));
  OAI21_X1   g08178(.A1(new_n8361_), .A2(new_n8359_), .B(\asqrt[32] ), .ZN(new_n8371_));
  NOR2_X1    g08179(.A1(new_n7955_), .A2(new_n6708_), .ZN(new_n8372_));
  NOR2_X1    g08180(.A1(new_n8185_), .A2(new_n8184_), .ZN(new_n8373_));
  NOR4_X1    g08181(.A1(new_n8319_), .A2(\asqrt[32] ), .A3(new_n8373_), .A4(new_n8189_), .ZN(new_n8374_));
  XNOR2_X1   g08182(.A1(new_n8374_), .A2(new_n8372_), .ZN(new_n8375_));
  NAND2_X1   g08183(.A1(new_n8375_), .A2(new_n6365_), .ZN(new_n8376_));
  INV_X1     g08184(.I(new_n8376_), .ZN(new_n8377_));
  AOI21_X1   g08185(.A1(new_n8371_), .A2(new_n8377_), .B(new_n8370_), .ZN(new_n8378_));
  AOI21_X1   g08186(.A1(new_n8370_), .A2(new_n8371_), .B(new_n6365_), .ZN(new_n8379_));
  NAND2_X1   g08187(.A1(new_n7966_), .A2(\asqrt[33] ), .ZN(new_n8380_));
  NOR2_X1    g08188(.A1(new_n7961_), .A2(new_n7962_), .ZN(new_n8381_));
  NOR4_X1    g08189(.A1(new_n8319_), .A2(\asqrt[33] ), .A3(new_n8381_), .A4(new_n7966_), .ZN(new_n8382_));
  XOR2_X1    g08190(.A1(new_n8382_), .A2(new_n8380_), .Z(new_n8383_));
  NAND2_X1   g08191(.A1(new_n8383_), .A2(new_n5991_), .ZN(new_n8384_));
  OAI21_X1   g08192(.A1(new_n8379_), .A2(new_n8384_), .B(new_n8378_), .ZN(new_n8385_));
  OAI21_X1   g08193(.A1(new_n8378_), .A2(new_n8379_), .B(\asqrt[34] ), .ZN(new_n8386_));
  NOR2_X1    g08194(.A1(new_n7973_), .A2(new_n5991_), .ZN(new_n8387_));
  NOR4_X1    g08195(.A1(new_n8319_), .A2(\asqrt[34] ), .A3(new_n7969_), .A4(new_n8197_), .ZN(new_n8388_));
  XNOR2_X1   g08196(.A1(new_n8388_), .A2(new_n8387_), .ZN(new_n8389_));
  NAND2_X1   g08197(.A1(new_n8389_), .A2(new_n5626_), .ZN(new_n8390_));
  INV_X1     g08198(.I(new_n8390_), .ZN(new_n8391_));
  AOI21_X1   g08199(.A1(new_n8386_), .A2(new_n8391_), .B(new_n8385_), .ZN(new_n8392_));
  AOI22_X1   g08200(.A1(new_n8347_), .A2(new_n8312_), .B1(\asqrt[30] ), .B2(new_n8349_), .ZN(new_n8393_));
  OAI21_X1   g08201(.A1(new_n8393_), .A2(new_n7110_), .B(new_n8368_), .ZN(new_n8394_));
  OAI22_X1   g08202(.A1(new_n8393_), .A2(new_n7110_), .B1(new_n8348_), .B2(new_n8358_), .ZN(new_n8395_));
  AOI22_X1   g08203(.A1(new_n8395_), .A2(\asqrt[32] ), .B1(new_n8394_), .B2(new_n8359_), .ZN(new_n8396_));
  INV_X1     g08204(.I(new_n8384_), .ZN(new_n8397_));
  OAI21_X1   g08205(.A1(new_n8396_), .A2(new_n6365_), .B(new_n8397_), .ZN(new_n8398_));
  AOI21_X1   g08206(.A1(new_n8395_), .A2(\asqrt[32] ), .B(new_n8376_), .ZN(new_n8399_));
  OAI22_X1   g08207(.A1(new_n8396_), .A2(new_n6365_), .B1(new_n8399_), .B2(new_n8370_), .ZN(new_n8400_));
  AOI22_X1   g08208(.A1(new_n8400_), .A2(\asqrt[34] ), .B1(new_n8398_), .B2(new_n8378_), .ZN(new_n8401_));
  NAND2_X1   g08209(.A1(new_n7980_), .A2(\asqrt[35] ), .ZN(new_n8402_));
  NOR4_X1    g08210(.A1(new_n8319_), .A2(\asqrt[35] ), .A3(new_n7975_), .A4(new_n7980_), .ZN(new_n8403_));
  XOR2_X1    g08211(.A1(new_n8403_), .A2(new_n8402_), .Z(new_n8404_));
  NAND2_X1   g08212(.A1(new_n8404_), .A2(new_n5273_), .ZN(new_n8405_));
  INV_X1     g08213(.I(new_n8405_), .ZN(new_n8406_));
  OAI21_X1   g08214(.A1(new_n8401_), .A2(new_n5626_), .B(new_n8406_), .ZN(new_n8407_));
  NAND2_X1   g08215(.A1(new_n8407_), .A2(new_n8392_), .ZN(new_n8408_));
  AOI21_X1   g08216(.A1(new_n8400_), .A2(\asqrt[34] ), .B(new_n8390_), .ZN(new_n8409_));
  OAI22_X1   g08217(.A1(new_n8401_), .A2(new_n5626_), .B1(new_n8409_), .B2(new_n8385_), .ZN(new_n8410_));
  NOR4_X1    g08218(.A1(new_n8319_), .A2(\asqrt[36] ), .A3(new_n7983_), .A4(new_n8204_), .ZN(new_n8411_));
  AOI21_X1   g08219(.A1(new_n8402_), .A2(new_n7979_), .B(new_n5273_), .ZN(new_n8412_));
  NOR2_X1    g08220(.A1(new_n8411_), .A2(new_n8412_), .ZN(new_n8413_));
  NAND2_X1   g08221(.A1(new_n8413_), .A2(new_n4973_), .ZN(new_n8414_));
  AOI21_X1   g08222(.A1(new_n8410_), .A2(\asqrt[36] ), .B(new_n8414_), .ZN(new_n8415_));
  NOR2_X1    g08223(.A1(new_n8415_), .A2(new_n8408_), .ZN(new_n8416_));
  AOI22_X1   g08224(.A1(new_n8410_), .A2(\asqrt[36] ), .B1(new_n8407_), .B2(new_n8392_), .ZN(new_n8417_));
  NAND2_X1   g08225(.A1(new_n7994_), .A2(\asqrt[37] ), .ZN(new_n8418_));
  NOR4_X1    g08226(.A1(new_n8319_), .A2(\asqrt[37] ), .A3(new_n7989_), .A4(new_n7994_), .ZN(new_n8419_));
  XOR2_X1    g08227(.A1(new_n8419_), .A2(new_n8418_), .Z(new_n8420_));
  NAND2_X1   g08228(.A1(new_n8420_), .A2(new_n4645_), .ZN(new_n8421_));
  INV_X1     g08229(.I(new_n8421_), .ZN(new_n8422_));
  OAI21_X1   g08230(.A1(new_n8417_), .A2(new_n4973_), .B(new_n8422_), .ZN(new_n8423_));
  NAND2_X1   g08231(.A1(new_n8423_), .A2(new_n8416_), .ZN(new_n8424_));
  OAI22_X1   g08232(.A1(new_n8417_), .A2(new_n4973_), .B1(new_n8415_), .B2(new_n8408_), .ZN(new_n8425_));
  NOR4_X1    g08233(.A1(new_n8319_), .A2(\asqrt[38] ), .A3(new_n7996_), .A4(new_n8211_), .ZN(new_n8426_));
  AOI21_X1   g08234(.A1(new_n8418_), .A2(new_n7993_), .B(new_n4645_), .ZN(new_n8427_));
  NOR2_X1    g08235(.A1(new_n8426_), .A2(new_n8427_), .ZN(new_n8428_));
  NAND2_X1   g08236(.A1(new_n8428_), .A2(new_n4330_), .ZN(new_n8429_));
  AOI21_X1   g08237(.A1(new_n8425_), .A2(\asqrt[38] ), .B(new_n8429_), .ZN(new_n8430_));
  NOR2_X1    g08238(.A1(new_n8430_), .A2(new_n8424_), .ZN(new_n8431_));
  AOI22_X1   g08239(.A1(new_n8425_), .A2(\asqrt[38] ), .B1(new_n8423_), .B2(new_n8416_), .ZN(new_n8432_));
  NAND2_X1   g08240(.A1(new_n8007_), .A2(\asqrt[39] ), .ZN(new_n8433_));
  NOR4_X1    g08241(.A1(new_n8319_), .A2(\asqrt[39] ), .A3(new_n8002_), .A4(new_n8007_), .ZN(new_n8434_));
  XOR2_X1    g08242(.A1(new_n8434_), .A2(new_n8433_), .Z(new_n8435_));
  NAND2_X1   g08243(.A1(new_n8435_), .A2(new_n4018_), .ZN(new_n8436_));
  INV_X1     g08244(.I(new_n8436_), .ZN(new_n8437_));
  OAI21_X1   g08245(.A1(new_n8432_), .A2(new_n4330_), .B(new_n8437_), .ZN(new_n8438_));
  NAND2_X1   g08246(.A1(new_n8438_), .A2(new_n8431_), .ZN(new_n8439_));
  OAI22_X1   g08247(.A1(new_n8432_), .A2(new_n4330_), .B1(new_n8430_), .B2(new_n8424_), .ZN(new_n8440_));
  NAND2_X1   g08248(.A1(new_n8218_), .A2(\asqrt[40] ), .ZN(new_n8441_));
  NOR4_X1    g08249(.A1(new_n8319_), .A2(\asqrt[40] ), .A3(new_n8010_), .A4(new_n8218_), .ZN(new_n8442_));
  XOR2_X1    g08250(.A1(new_n8442_), .A2(new_n8441_), .Z(new_n8443_));
  NAND2_X1   g08251(.A1(new_n8443_), .A2(new_n3760_), .ZN(new_n8444_));
  AOI21_X1   g08252(.A1(new_n8440_), .A2(\asqrt[40] ), .B(new_n8444_), .ZN(new_n8445_));
  NOR2_X1    g08253(.A1(new_n8445_), .A2(new_n8439_), .ZN(new_n8446_));
  AOI22_X1   g08254(.A1(new_n8440_), .A2(\asqrt[40] ), .B1(new_n8438_), .B2(new_n8431_), .ZN(new_n8447_));
  NOR4_X1    g08255(.A1(new_n8319_), .A2(\asqrt[41] ), .A3(new_n8017_), .A4(new_n8022_), .ZN(new_n8448_));
  AOI21_X1   g08256(.A1(new_n8441_), .A2(new_n8217_), .B(new_n3760_), .ZN(new_n8449_));
  NOR2_X1    g08257(.A1(new_n8448_), .A2(new_n8449_), .ZN(new_n8450_));
  NAND2_X1   g08258(.A1(new_n8450_), .A2(new_n3481_), .ZN(new_n8451_));
  INV_X1     g08259(.I(new_n8451_), .ZN(new_n8452_));
  OAI21_X1   g08260(.A1(new_n8447_), .A2(new_n3760_), .B(new_n8452_), .ZN(new_n8453_));
  NAND2_X1   g08261(.A1(new_n8453_), .A2(new_n8446_), .ZN(new_n8454_));
  OAI22_X1   g08262(.A1(new_n8447_), .A2(new_n3760_), .B1(new_n8445_), .B2(new_n8439_), .ZN(new_n8455_));
  NAND2_X1   g08263(.A1(new_n8225_), .A2(\asqrt[42] ), .ZN(new_n8456_));
  NOR4_X1    g08264(.A1(new_n8319_), .A2(\asqrt[42] ), .A3(new_n8025_), .A4(new_n8225_), .ZN(new_n8457_));
  XOR2_X1    g08265(.A1(new_n8457_), .A2(new_n8456_), .Z(new_n8458_));
  NAND2_X1   g08266(.A1(new_n8458_), .A2(new_n3208_), .ZN(new_n8459_));
  AOI21_X1   g08267(.A1(new_n8455_), .A2(\asqrt[42] ), .B(new_n8459_), .ZN(new_n8460_));
  NOR2_X1    g08268(.A1(new_n8460_), .A2(new_n8454_), .ZN(new_n8461_));
  AOI22_X1   g08269(.A1(new_n8455_), .A2(\asqrt[42] ), .B1(new_n8453_), .B2(new_n8446_), .ZN(new_n8462_));
  NOR4_X1    g08270(.A1(new_n8319_), .A2(\asqrt[43] ), .A3(new_n8032_), .A4(new_n8037_), .ZN(new_n8463_));
  AOI21_X1   g08271(.A1(new_n8456_), .A2(new_n8224_), .B(new_n3208_), .ZN(new_n8464_));
  NOR2_X1    g08272(.A1(new_n8463_), .A2(new_n8464_), .ZN(new_n8465_));
  NAND2_X1   g08273(.A1(new_n8465_), .A2(new_n2941_), .ZN(new_n8466_));
  INV_X1     g08274(.I(new_n8466_), .ZN(new_n8467_));
  OAI21_X1   g08275(.A1(new_n8462_), .A2(new_n3208_), .B(new_n8467_), .ZN(new_n8468_));
  NAND2_X1   g08276(.A1(new_n8468_), .A2(new_n8461_), .ZN(new_n8469_));
  OAI22_X1   g08277(.A1(new_n8462_), .A2(new_n3208_), .B1(new_n8460_), .B2(new_n8454_), .ZN(new_n8470_));
  NAND2_X1   g08278(.A1(new_n8232_), .A2(\asqrt[44] ), .ZN(new_n8471_));
  NOR4_X1    g08279(.A1(new_n8319_), .A2(\asqrt[44] ), .A3(new_n8040_), .A4(new_n8232_), .ZN(new_n8472_));
  XOR2_X1    g08280(.A1(new_n8472_), .A2(new_n8471_), .Z(new_n8473_));
  NAND2_X1   g08281(.A1(new_n8473_), .A2(new_n2728_), .ZN(new_n8474_));
  AOI21_X1   g08282(.A1(new_n8470_), .A2(\asqrt[44] ), .B(new_n8474_), .ZN(new_n8475_));
  NOR2_X1    g08283(.A1(new_n8475_), .A2(new_n8469_), .ZN(new_n8476_));
  AOI22_X1   g08284(.A1(new_n8470_), .A2(\asqrt[44] ), .B1(new_n8468_), .B2(new_n8461_), .ZN(new_n8477_));
  NOR4_X1    g08285(.A1(new_n8319_), .A2(\asqrt[45] ), .A3(new_n8047_), .A4(new_n8052_), .ZN(new_n8478_));
  AOI21_X1   g08286(.A1(new_n8471_), .A2(new_n8231_), .B(new_n2728_), .ZN(new_n8479_));
  NOR2_X1    g08287(.A1(new_n8478_), .A2(new_n8479_), .ZN(new_n8480_));
  NAND2_X1   g08288(.A1(new_n8480_), .A2(new_n2488_), .ZN(new_n8481_));
  INV_X1     g08289(.I(new_n8481_), .ZN(new_n8482_));
  OAI21_X1   g08290(.A1(new_n8477_), .A2(new_n2728_), .B(new_n8482_), .ZN(new_n8483_));
  NAND2_X1   g08291(.A1(new_n8483_), .A2(new_n8476_), .ZN(new_n8484_));
  OAI22_X1   g08292(.A1(new_n8477_), .A2(new_n2728_), .B1(new_n8475_), .B2(new_n8469_), .ZN(new_n8485_));
  NAND2_X1   g08293(.A1(new_n8239_), .A2(\asqrt[46] ), .ZN(new_n8486_));
  NOR4_X1    g08294(.A1(new_n8319_), .A2(\asqrt[46] ), .A3(new_n8055_), .A4(new_n8239_), .ZN(new_n8487_));
  XOR2_X1    g08295(.A1(new_n8487_), .A2(new_n8486_), .Z(new_n8488_));
  NAND2_X1   g08296(.A1(new_n8488_), .A2(new_n2253_), .ZN(new_n8489_));
  AOI21_X1   g08297(.A1(new_n8485_), .A2(\asqrt[46] ), .B(new_n8489_), .ZN(new_n8490_));
  NOR2_X1    g08298(.A1(new_n8490_), .A2(new_n8484_), .ZN(new_n8491_));
  AOI22_X1   g08299(.A1(new_n8485_), .A2(\asqrt[46] ), .B1(new_n8483_), .B2(new_n8476_), .ZN(new_n8492_));
  NOR4_X1    g08300(.A1(new_n8319_), .A2(\asqrt[47] ), .A3(new_n8062_), .A4(new_n8067_), .ZN(new_n8493_));
  AOI21_X1   g08301(.A1(new_n8486_), .A2(new_n8238_), .B(new_n2253_), .ZN(new_n8494_));
  NOR2_X1    g08302(.A1(new_n8493_), .A2(new_n8494_), .ZN(new_n8495_));
  NAND2_X1   g08303(.A1(new_n8495_), .A2(new_n2046_), .ZN(new_n8496_));
  INV_X1     g08304(.I(new_n8496_), .ZN(new_n8497_));
  OAI21_X1   g08305(.A1(new_n8492_), .A2(new_n2253_), .B(new_n8497_), .ZN(new_n8498_));
  NAND2_X1   g08306(.A1(new_n8498_), .A2(new_n8491_), .ZN(new_n8499_));
  OAI22_X1   g08307(.A1(new_n8492_), .A2(new_n2253_), .B1(new_n8490_), .B2(new_n8484_), .ZN(new_n8500_));
  NAND2_X1   g08308(.A1(new_n8246_), .A2(\asqrt[48] ), .ZN(new_n8501_));
  NOR4_X1    g08309(.A1(new_n8319_), .A2(\asqrt[48] ), .A3(new_n8070_), .A4(new_n8246_), .ZN(new_n8502_));
  XOR2_X1    g08310(.A1(new_n8502_), .A2(new_n8501_), .Z(new_n8503_));
  NAND2_X1   g08311(.A1(new_n8503_), .A2(new_n1854_), .ZN(new_n8504_));
  AOI21_X1   g08312(.A1(new_n8500_), .A2(\asqrt[48] ), .B(new_n8504_), .ZN(new_n8505_));
  NOR2_X1    g08313(.A1(new_n8505_), .A2(new_n8499_), .ZN(new_n8506_));
  AOI22_X1   g08314(.A1(new_n8500_), .A2(\asqrt[48] ), .B1(new_n8498_), .B2(new_n8491_), .ZN(new_n8507_));
  NAND2_X1   g08315(.A1(new_n8082_), .A2(\asqrt[49] ), .ZN(new_n8508_));
  NOR4_X1    g08316(.A1(new_n8319_), .A2(\asqrt[49] ), .A3(new_n8077_), .A4(new_n8082_), .ZN(new_n8509_));
  XOR2_X1    g08317(.A1(new_n8509_), .A2(new_n8508_), .Z(new_n8510_));
  NAND2_X1   g08318(.A1(new_n8510_), .A2(new_n1595_), .ZN(new_n8511_));
  INV_X1     g08319(.I(new_n8511_), .ZN(new_n8512_));
  OAI21_X1   g08320(.A1(new_n8507_), .A2(new_n1854_), .B(new_n8512_), .ZN(new_n8513_));
  NAND2_X1   g08321(.A1(new_n8513_), .A2(new_n8506_), .ZN(new_n8514_));
  OAI22_X1   g08322(.A1(new_n8507_), .A2(new_n1854_), .B1(new_n8505_), .B2(new_n8499_), .ZN(new_n8515_));
  NOR4_X1    g08323(.A1(new_n8319_), .A2(\asqrt[50] ), .A3(new_n8085_), .A4(new_n8253_), .ZN(new_n8516_));
  AOI21_X1   g08324(.A1(new_n8508_), .A2(new_n8081_), .B(new_n1595_), .ZN(new_n8517_));
  NOR2_X1    g08325(.A1(new_n8516_), .A2(new_n8517_), .ZN(new_n8518_));
  NAND2_X1   g08326(.A1(new_n8518_), .A2(new_n1436_), .ZN(new_n8519_));
  AOI21_X1   g08327(.A1(new_n8515_), .A2(\asqrt[50] ), .B(new_n8519_), .ZN(new_n8520_));
  NOR2_X1    g08328(.A1(new_n8520_), .A2(new_n8514_), .ZN(new_n8521_));
  AOI22_X1   g08329(.A1(new_n8515_), .A2(\asqrt[50] ), .B1(new_n8513_), .B2(new_n8506_), .ZN(new_n8522_));
  NAND2_X1   g08330(.A1(new_n8097_), .A2(\asqrt[51] ), .ZN(new_n8523_));
  NOR4_X1    g08331(.A1(new_n8319_), .A2(\asqrt[51] ), .A3(new_n8092_), .A4(new_n8097_), .ZN(new_n8524_));
  XOR2_X1    g08332(.A1(new_n8524_), .A2(new_n8523_), .Z(new_n8525_));
  NAND2_X1   g08333(.A1(new_n8525_), .A2(new_n1260_), .ZN(new_n8526_));
  INV_X1     g08334(.I(new_n8526_), .ZN(new_n8527_));
  OAI21_X1   g08335(.A1(new_n8522_), .A2(new_n1436_), .B(new_n8527_), .ZN(new_n8528_));
  NAND2_X1   g08336(.A1(new_n8528_), .A2(new_n8521_), .ZN(new_n8529_));
  OAI22_X1   g08337(.A1(new_n8522_), .A2(new_n1436_), .B1(new_n8520_), .B2(new_n8514_), .ZN(new_n8530_));
  NOR4_X1    g08338(.A1(new_n8319_), .A2(\asqrt[52] ), .A3(new_n8100_), .A4(new_n8260_), .ZN(new_n8531_));
  AOI21_X1   g08339(.A1(new_n8523_), .A2(new_n8096_), .B(new_n1260_), .ZN(new_n8532_));
  NOR2_X1    g08340(.A1(new_n8531_), .A2(new_n8532_), .ZN(new_n8533_));
  NAND2_X1   g08341(.A1(new_n8533_), .A2(new_n1096_), .ZN(new_n8534_));
  AOI21_X1   g08342(.A1(new_n8530_), .A2(\asqrt[52] ), .B(new_n8534_), .ZN(new_n8535_));
  NOR2_X1    g08343(.A1(new_n8535_), .A2(new_n8529_), .ZN(new_n8536_));
  AOI22_X1   g08344(.A1(new_n8530_), .A2(\asqrt[52] ), .B1(new_n8528_), .B2(new_n8521_), .ZN(new_n8537_));
  NAND2_X1   g08345(.A1(new_n8112_), .A2(\asqrt[53] ), .ZN(new_n8538_));
  NOR4_X1    g08346(.A1(new_n8319_), .A2(\asqrt[53] ), .A3(new_n8107_), .A4(new_n8112_), .ZN(new_n8539_));
  XOR2_X1    g08347(.A1(new_n8539_), .A2(new_n8538_), .Z(new_n8540_));
  NAND2_X1   g08348(.A1(new_n8540_), .A2(new_n970_), .ZN(new_n8541_));
  INV_X1     g08349(.I(new_n8541_), .ZN(new_n8542_));
  OAI21_X1   g08350(.A1(new_n8537_), .A2(new_n1096_), .B(new_n8542_), .ZN(new_n8543_));
  NAND2_X1   g08351(.A1(new_n8543_), .A2(new_n8536_), .ZN(new_n8544_));
  OAI22_X1   g08352(.A1(new_n8537_), .A2(new_n1096_), .B1(new_n8535_), .B2(new_n8529_), .ZN(new_n8545_));
  NOR2_X1    g08353(.A1(new_n8119_), .A2(new_n970_), .ZN(new_n8546_));
  NOR4_X1    g08354(.A1(new_n8319_), .A2(\asqrt[54] ), .A3(new_n8115_), .A4(new_n8267_), .ZN(new_n8547_));
  XNOR2_X1   g08355(.A1(new_n8547_), .A2(new_n8546_), .ZN(new_n8548_));
  NAND2_X1   g08356(.A1(new_n8548_), .A2(new_n825_), .ZN(new_n8549_));
  AOI21_X1   g08357(.A1(new_n8545_), .A2(\asqrt[54] ), .B(new_n8549_), .ZN(new_n8550_));
  NOR2_X1    g08358(.A1(new_n8550_), .A2(new_n8544_), .ZN(new_n8551_));
  AOI22_X1   g08359(.A1(new_n8545_), .A2(\asqrt[54] ), .B1(new_n8543_), .B2(new_n8536_), .ZN(new_n8552_));
  NOR4_X1    g08360(.A1(new_n8319_), .A2(\asqrt[55] ), .A3(new_n8121_), .A4(new_n8126_), .ZN(new_n8553_));
  XOR2_X1    g08361(.A1(new_n8553_), .A2(new_n8320_), .Z(new_n8554_));
  NAND2_X1   g08362(.A1(new_n8554_), .A2(new_n724_), .ZN(new_n8555_));
  INV_X1     g08363(.I(new_n8555_), .ZN(new_n8556_));
  OAI21_X1   g08364(.A1(new_n8552_), .A2(new_n825_), .B(new_n8556_), .ZN(new_n8557_));
  NAND2_X1   g08365(.A1(new_n8557_), .A2(new_n8551_), .ZN(new_n8558_));
  OAI22_X1   g08366(.A1(new_n8552_), .A2(new_n825_), .B1(new_n8550_), .B2(new_n8544_), .ZN(new_n8559_));
  NOR4_X1    g08367(.A1(new_n8319_), .A2(\asqrt[56] ), .A3(new_n8128_), .A4(new_n8274_), .ZN(new_n8560_));
  XOR2_X1    g08368(.A1(new_n8560_), .A2(new_n8335_), .Z(new_n8561_));
  NAND2_X1   g08369(.A1(new_n8561_), .A2(new_n587_), .ZN(new_n8562_));
  AOI21_X1   g08370(.A1(new_n8559_), .A2(\asqrt[56] ), .B(new_n8562_), .ZN(new_n8563_));
  NOR2_X1    g08371(.A1(new_n8563_), .A2(new_n8558_), .ZN(new_n8564_));
  AOI22_X1   g08372(.A1(new_n8559_), .A2(\asqrt[56] ), .B1(new_n8557_), .B2(new_n8551_), .ZN(new_n8565_));
  NOR4_X1    g08373(.A1(new_n8319_), .A2(\asqrt[57] ), .A3(new_n8134_), .A4(new_n8139_), .ZN(new_n8566_));
  XOR2_X1    g08374(.A1(new_n8566_), .A2(new_n8322_), .Z(new_n8567_));
  AND2_X2    g08375(.A1(new_n8567_), .A2(new_n504_), .Z(new_n8568_));
  OAI21_X1   g08376(.A1(new_n8565_), .A2(new_n587_), .B(new_n8568_), .ZN(new_n8569_));
  NAND2_X1   g08377(.A1(new_n8569_), .A2(new_n8564_), .ZN(new_n8570_));
  OAI22_X1   g08378(.A1(new_n8565_), .A2(new_n587_), .B1(new_n8563_), .B2(new_n8558_), .ZN(new_n8571_));
  NOR4_X1    g08379(.A1(new_n8319_), .A2(\asqrt[58] ), .A3(new_n8141_), .A4(new_n8281_), .ZN(new_n8572_));
  XOR2_X1    g08380(.A1(new_n8572_), .A2(new_n8337_), .Z(new_n8573_));
  NAND2_X1   g08381(.A1(new_n8573_), .A2(new_n376_), .ZN(new_n8574_));
  AOI21_X1   g08382(.A1(new_n8571_), .A2(\asqrt[58] ), .B(new_n8574_), .ZN(new_n8575_));
  NOR2_X1    g08383(.A1(new_n8575_), .A2(new_n8570_), .ZN(new_n8576_));
  AOI22_X1   g08384(.A1(new_n8571_), .A2(\asqrt[58] ), .B1(new_n8569_), .B2(new_n8564_), .ZN(new_n8577_));
  NOR4_X1    g08385(.A1(new_n8319_), .A2(\asqrt[59] ), .A3(new_n8147_), .A4(new_n8152_), .ZN(new_n8578_));
  XOR2_X1    g08386(.A1(new_n8578_), .A2(new_n8324_), .Z(new_n8579_));
  AND2_X2    g08387(.A1(new_n8579_), .A2(new_n275_), .Z(new_n8580_));
  OAI21_X1   g08388(.A1(new_n8577_), .A2(new_n376_), .B(new_n8580_), .ZN(new_n8581_));
  NAND2_X1   g08389(.A1(new_n8581_), .A2(new_n8576_), .ZN(new_n8582_));
  NAND2_X1   g08390(.A1(new_n8530_), .A2(\asqrt[52] ), .ZN(new_n8583_));
  AOI21_X1   g08391(.A1(new_n8583_), .A2(new_n8529_), .B(new_n1096_), .ZN(new_n8584_));
  OAI21_X1   g08392(.A1(new_n8536_), .A2(new_n8584_), .B(\asqrt[54] ), .ZN(new_n8585_));
  AOI21_X1   g08393(.A1(new_n8544_), .A2(new_n8585_), .B(new_n825_), .ZN(new_n8586_));
  OAI21_X1   g08394(.A1(new_n8551_), .A2(new_n8586_), .B(\asqrt[56] ), .ZN(new_n8587_));
  AOI21_X1   g08395(.A1(new_n8558_), .A2(new_n8587_), .B(new_n587_), .ZN(new_n8588_));
  OAI21_X1   g08396(.A1(new_n8564_), .A2(new_n8588_), .B(\asqrt[58] ), .ZN(new_n8589_));
  AOI21_X1   g08397(.A1(new_n8570_), .A2(new_n8589_), .B(new_n376_), .ZN(new_n8590_));
  OAI21_X1   g08398(.A1(new_n8576_), .A2(new_n8590_), .B(\asqrt[60] ), .ZN(new_n8591_));
  AOI21_X1   g08399(.A1(new_n8582_), .A2(new_n8591_), .B(new_n229_), .ZN(new_n8592_));
  NOR2_X1    g08400(.A1(new_n8306_), .A2(new_n196_), .ZN(new_n8593_));
  NOR2_X1    g08401(.A1(new_n8291_), .A2(\asqrt[62] ), .ZN(new_n8594_));
  NAND3_X1   g08402(.A1(new_n8594_), .A2(new_n8593_), .A3(new_n8166_), .ZN(new_n8595_));
  NOR2_X1    g08403(.A1(new_n8319_), .A2(new_n8595_), .ZN(new_n8596_));
  OR3_X2     g08404(.A1(\asqrt[28] ), .A2(new_n8166_), .A3(new_n8594_), .Z(new_n8597_));
  AOI21_X1   g08405(.A1(new_n8597_), .A2(new_n8593_), .B(new_n8596_), .ZN(new_n8598_));
  NOR4_X1    g08406(.A1(new_n8319_), .A2(\asqrt[61] ), .A3(new_n8160_), .A4(new_n8165_), .ZN(new_n8599_));
  XOR2_X1    g08407(.A1(new_n8599_), .A2(new_n8326_), .Z(new_n8600_));
  NOR2_X1    g08408(.A1(new_n8600_), .A2(new_n196_), .ZN(new_n8601_));
  INV_X1     g08409(.I(new_n8601_), .ZN(new_n8602_));
  NOR2_X1    g08410(.A1(new_n8379_), .A2(new_n8384_), .ZN(new_n8603_));
  NOR3_X1    g08411(.A1(new_n8603_), .A2(new_n8370_), .A3(new_n8399_), .ZN(new_n8604_));
  NAND2_X1   g08412(.A1(new_n8386_), .A2(new_n8391_), .ZN(new_n8605_));
  NAND2_X1   g08413(.A1(new_n8605_), .A2(new_n8604_), .ZN(new_n8606_));
  NAND2_X1   g08414(.A1(new_n8385_), .A2(new_n8386_), .ZN(new_n8607_));
  AOI21_X1   g08415(.A1(new_n8607_), .A2(\asqrt[35] ), .B(new_n8405_), .ZN(new_n8608_));
  NOR2_X1    g08416(.A1(new_n8608_), .A2(new_n8606_), .ZN(new_n8609_));
  AOI21_X1   g08417(.A1(new_n8385_), .A2(new_n8386_), .B(new_n5626_), .ZN(new_n8610_));
  OAI21_X1   g08418(.A1(new_n8392_), .A2(new_n8610_), .B(\asqrt[36] ), .ZN(new_n8611_));
  INV_X1     g08419(.I(new_n8414_), .ZN(new_n8612_));
  NAND2_X1   g08420(.A1(new_n8611_), .A2(new_n8612_), .ZN(new_n8613_));
  NAND2_X1   g08421(.A1(new_n8613_), .A2(new_n8609_), .ZN(new_n8614_));
  AOI22_X1   g08422(.A1(new_n8607_), .A2(\asqrt[35] ), .B1(new_n8605_), .B2(new_n8604_), .ZN(new_n8615_));
  OAI22_X1   g08423(.A1(new_n8615_), .A2(new_n5273_), .B1(new_n8608_), .B2(new_n8606_), .ZN(new_n8616_));
  AOI21_X1   g08424(.A1(new_n8616_), .A2(\asqrt[37] ), .B(new_n8421_), .ZN(new_n8617_));
  NOR2_X1    g08425(.A1(new_n8617_), .A2(new_n8614_), .ZN(new_n8618_));
  AOI22_X1   g08426(.A1(new_n8616_), .A2(\asqrt[37] ), .B1(new_n8613_), .B2(new_n8609_), .ZN(new_n8619_));
  INV_X1     g08427(.I(new_n8429_), .ZN(new_n8620_));
  OAI21_X1   g08428(.A1(new_n8619_), .A2(new_n4645_), .B(new_n8620_), .ZN(new_n8621_));
  NAND2_X1   g08429(.A1(new_n8621_), .A2(new_n8618_), .ZN(new_n8622_));
  OAI22_X1   g08430(.A1(new_n8619_), .A2(new_n4645_), .B1(new_n8617_), .B2(new_n8614_), .ZN(new_n8623_));
  AOI21_X1   g08431(.A1(new_n8623_), .A2(\asqrt[39] ), .B(new_n8436_), .ZN(new_n8624_));
  NOR2_X1    g08432(.A1(new_n8624_), .A2(new_n8622_), .ZN(new_n8625_));
  AOI22_X1   g08433(.A1(new_n8623_), .A2(\asqrt[39] ), .B1(new_n8621_), .B2(new_n8618_), .ZN(new_n8626_));
  INV_X1     g08434(.I(new_n8444_), .ZN(new_n8627_));
  OAI21_X1   g08435(.A1(new_n8626_), .A2(new_n4018_), .B(new_n8627_), .ZN(new_n8628_));
  NAND2_X1   g08436(.A1(new_n8628_), .A2(new_n8625_), .ZN(new_n8629_));
  OAI22_X1   g08437(.A1(new_n8626_), .A2(new_n4018_), .B1(new_n8624_), .B2(new_n8622_), .ZN(new_n8630_));
  AOI21_X1   g08438(.A1(new_n8630_), .A2(\asqrt[41] ), .B(new_n8451_), .ZN(new_n8631_));
  NOR2_X1    g08439(.A1(new_n8631_), .A2(new_n8629_), .ZN(new_n8632_));
  AOI22_X1   g08440(.A1(new_n8630_), .A2(\asqrt[41] ), .B1(new_n8628_), .B2(new_n8625_), .ZN(new_n8633_));
  INV_X1     g08441(.I(new_n8459_), .ZN(new_n8634_));
  OAI21_X1   g08442(.A1(new_n8633_), .A2(new_n3481_), .B(new_n8634_), .ZN(new_n8635_));
  NAND2_X1   g08443(.A1(new_n8635_), .A2(new_n8632_), .ZN(new_n8636_));
  OAI22_X1   g08444(.A1(new_n8633_), .A2(new_n3481_), .B1(new_n8631_), .B2(new_n8629_), .ZN(new_n8637_));
  AOI21_X1   g08445(.A1(new_n8637_), .A2(\asqrt[43] ), .B(new_n8466_), .ZN(new_n8638_));
  NOR2_X1    g08446(.A1(new_n8638_), .A2(new_n8636_), .ZN(new_n8639_));
  AOI22_X1   g08447(.A1(new_n8637_), .A2(\asqrt[43] ), .B1(new_n8635_), .B2(new_n8632_), .ZN(new_n8640_));
  INV_X1     g08448(.I(new_n8474_), .ZN(new_n8641_));
  OAI21_X1   g08449(.A1(new_n8640_), .A2(new_n2941_), .B(new_n8641_), .ZN(new_n8642_));
  NAND2_X1   g08450(.A1(new_n8642_), .A2(new_n8639_), .ZN(new_n8643_));
  OAI22_X1   g08451(.A1(new_n8640_), .A2(new_n2941_), .B1(new_n8638_), .B2(new_n8636_), .ZN(new_n8644_));
  AOI21_X1   g08452(.A1(new_n8644_), .A2(\asqrt[45] ), .B(new_n8481_), .ZN(new_n8645_));
  NOR2_X1    g08453(.A1(new_n8645_), .A2(new_n8643_), .ZN(new_n8646_));
  AOI22_X1   g08454(.A1(new_n8644_), .A2(\asqrt[45] ), .B1(new_n8642_), .B2(new_n8639_), .ZN(new_n8647_));
  INV_X1     g08455(.I(new_n8489_), .ZN(new_n8648_));
  OAI21_X1   g08456(.A1(new_n8647_), .A2(new_n2488_), .B(new_n8648_), .ZN(new_n8649_));
  NAND2_X1   g08457(.A1(new_n8649_), .A2(new_n8646_), .ZN(new_n8650_));
  OAI22_X1   g08458(.A1(new_n8647_), .A2(new_n2488_), .B1(new_n8645_), .B2(new_n8643_), .ZN(new_n8651_));
  AOI21_X1   g08459(.A1(new_n8651_), .A2(\asqrt[47] ), .B(new_n8496_), .ZN(new_n8652_));
  NOR2_X1    g08460(.A1(new_n8652_), .A2(new_n8650_), .ZN(new_n8653_));
  AOI22_X1   g08461(.A1(new_n8651_), .A2(\asqrt[47] ), .B1(new_n8649_), .B2(new_n8646_), .ZN(new_n8654_));
  INV_X1     g08462(.I(new_n8504_), .ZN(new_n8655_));
  OAI21_X1   g08463(.A1(new_n8654_), .A2(new_n2046_), .B(new_n8655_), .ZN(new_n8656_));
  NAND2_X1   g08464(.A1(new_n8656_), .A2(new_n8653_), .ZN(new_n8657_));
  OAI22_X1   g08465(.A1(new_n8654_), .A2(new_n2046_), .B1(new_n8652_), .B2(new_n8650_), .ZN(new_n8658_));
  AOI21_X1   g08466(.A1(new_n8658_), .A2(\asqrt[49] ), .B(new_n8511_), .ZN(new_n8659_));
  NOR2_X1    g08467(.A1(new_n8659_), .A2(new_n8657_), .ZN(new_n8660_));
  AOI22_X1   g08468(.A1(new_n8658_), .A2(\asqrt[49] ), .B1(new_n8656_), .B2(new_n8653_), .ZN(new_n8661_));
  INV_X1     g08469(.I(new_n8519_), .ZN(new_n8662_));
  OAI21_X1   g08470(.A1(new_n8661_), .A2(new_n1595_), .B(new_n8662_), .ZN(new_n8663_));
  NAND2_X1   g08471(.A1(new_n8663_), .A2(new_n8660_), .ZN(new_n8664_));
  OAI22_X1   g08472(.A1(new_n8661_), .A2(new_n1595_), .B1(new_n8659_), .B2(new_n8657_), .ZN(new_n8665_));
  AOI21_X1   g08473(.A1(new_n8665_), .A2(\asqrt[51] ), .B(new_n8526_), .ZN(new_n8666_));
  NOR2_X1    g08474(.A1(new_n8666_), .A2(new_n8664_), .ZN(new_n8667_));
  AOI22_X1   g08475(.A1(new_n8665_), .A2(\asqrt[51] ), .B1(new_n8663_), .B2(new_n8660_), .ZN(new_n8668_));
  INV_X1     g08476(.I(new_n8534_), .ZN(new_n8669_));
  OAI21_X1   g08477(.A1(new_n8668_), .A2(new_n1260_), .B(new_n8669_), .ZN(new_n8670_));
  NAND2_X1   g08478(.A1(new_n8670_), .A2(new_n8667_), .ZN(new_n8671_));
  OAI22_X1   g08479(.A1(new_n8668_), .A2(new_n1260_), .B1(new_n8666_), .B2(new_n8664_), .ZN(new_n8672_));
  AOI21_X1   g08480(.A1(new_n8672_), .A2(\asqrt[53] ), .B(new_n8541_), .ZN(new_n8673_));
  NOR2_X1    g08481(.A1(new_n8673_), .A2(new_n8671_), .ZN(new_n8674_));
  AOI22_X1   g08482(.A1(new_n8672_), .A2(\asqrt[53] ), .B1(new_n8670_), .B2(new_n8667_), .ZN(new_n8675_));
  INV_X1     g08483(.I(new_n8549_), .ZN(new_n8676_));
  OAI21_X1   g08484(.A1(new_n8675_), .A2(new_n970_), .B(new_n8676_), .ZN(new_n8677_));
  NAND2_X1   g08485(.A1(new_n8677_), .A2(new_n8674_), .ZN(new_n8678_));
  OAI22_X1   g08486(.A1(new_n8675_), .A2(new_n970_), .B1(new_n8673_), .B2(new_n8671_), .ZN(new_n8679_));
  AOI21_X1   g08487(.A1(new_n8679_), .A2(\asqrt[55] ), .B(new_n8555_), .ZN(new_n8680_));
  NOR2_X1    g08488(.A1(new_n8680_), .A2(new_n8678_), .ZN(new_n8681_));
  AOI22_X1   g08489(.A1(new_n8679_), .A2(\asqrt[55] ), .B1(new_n8677_), .B2(new_n8674_), .ZN(new_n8682_));
  INV_X1     g08490(.I(new_n8562_), .ZN(new_n8683_));
  OAI21_X1   g08491(.A1(new_n8682_), .A2(new_n724_), .B(new_n8683_), .ZN(new_n8684_));
  NAND2_X1   g08492(.A1(new_n8684_), .A2(new_n8681_), .ZN(new_n8685_));
  NAND2_X1   g08493(.A1(new_n8679_), .A2(\asqrt[55] ), .ZN(new_n8686_));
  AOI21_X1   g08494(.A1(new_n8686_), .A2(new_n8678_), .B(new_n724_), .ZN(new_n8687_));
  OAI21_X1   g08495(.A1(new_n8681_), .A2(new_n8687_), .B(\asqrt[57] ), .ZN(new_n8688_));
  AOI21_X1   g08496(.A1(new_n8688_), .A2(new_n8568_), .B(new_n8685_), .ZN(new_n8689_));
  OAI22_X1   g08497(.A1(new_n8682_), .A2(new_n724_), .B1(new_n8680_), .B2(new_n8678_), .ZN(new_n8690_));
  AOI22_X1   g08498(.A1(new_n8690_), .A2(\asqrt[57] ), .B1(new_n8684_), .B2(new_n8681_), .ZN(new_n8691_));
  INV_X1     g08499(.I(new_n8574_), .ZN(new_n8692_));
  OAI21_X1   g08500(.A1(new_n8691_), .A2(new_n504_), .B(new_n8692_), .ZN(new_n8693_));
  NAND2_X1   g08501(.A1(new_n8693_), .A2(new_n8689_), .ZN(new_n8694_));
  AOI21_X1   g08502(.A1(new_n8685_), .A2(new_n8688_), .B(new_n504_), .ZN(new_n8695_));
  OAI21_X1   g08503(.A1(new_n8689_), .A2(new_n8695_), .B(\asqrt[59] ), .ZN(new_n8696_));
  AOI21_X1   g08504(.A1(new_n8696_), .A2(new_n8580_), .B(new_n8694_), .ZN(new_n8697_));
  NAND2_X1   g08505(.A1(new_n8570_), .A2(new_n8589_), .ZN(new_n8698_));
  AOI22_X1   g08506(.A1(new_n8698_), .A2(\asqrt[59] ), .B1(new_n8693_), .B2(new_n8689_), .ZN(new_n8699_));
  NOR4_X1    g08507(.A1(new_n8319_), .A2(\asqrt[60] ), .A3(new_n8154_), .A4(new_n8288_), .ZN(new_n8700_));
  XOR2_X1    g08508(.A1(new_n8700_), .A2(new_n8339_), .Z(new_n8701_));
  NAND2_X1   g08509(.A1(new_n8701_), .A2(new_n229_), .ZN(new_n8702_));
  INV_X1     g08510(.I(new_n8702_), .ZN(new_n8703_));
  OAI21_X1   g08511(.A1(new_n8699_), .A2(new_n275_), .B(new_n8703_), .ZN(new_n8704_));
  NAND2_X1   g08512(.A1(new_n8704_), .A2(new_n8697_), .ZN(new_n8705_));
  INV_X1     g08513(.I(new_n8600_), .ZN(new_n8706_));
  NOR2_X1    g08514(.A1(new_n8706_), .A2(\asqrt[62] ), .ZN(new_n8707_));
  INV_X1     g08515(.I(new_n8707_), .ZN(new_n8708_));
  NAND2_X1   g08516(.A1(new_n8592_), .A2(new_n8708_), .ZN(new_n8709_));
  OAI21_X1   g08517(.A1(new_n8709_), .A2(new_n8705_), .B(new_n8602_), .ZN(new_n8710_));
  NOR3_X1    g08518(.A1(\asqrt[28] ), .A2(new_n7899_), .A3(new_n8292_), .ZN(new_n8711_));
  OAI21_X1   g08519(.A1(new_n8711_), .A2(new_n8304_), .B(new_n231_), .ZN(new_n8712_));
  OAI21_X1   g08520(.A1(new_n8710_), .A2(new_n8712_), .B(new_n8598_), .ZN(new_n8713_));
  OAI21_X1   g08521(.A1(new_n7899_), .A2(new_n8170_), .B(\asqrt[28] ), .ZN(new_n8714_));
  XOR2_X1    g08522(.A1(new_n8170_), .A2(\asqrt[63] ), .Z(new_n8715_));
  NAND2_X1   g08523(.A1(new_n8714_), .A2(new_n8715_), .ZN(new_n8716_));
  INV_X1     g08524(.I(new_n8716_), .ZN(new_n8717_));
  INV_X1     g08525(.I(new_n8598_), .ZN(new_n8718_));
  OAI22_X1   g08526(.A1(new_n8577_), .A2(new_n376_), .B1(new_n8575_), .B2(new_n8570_), .ZN(new_n8719_));
  AOI21_X1   g08527(.A1(new_n8719_), .A2(\asqrt[60] ), .B(new_n8702_), .ZN(new_n8720_));
  AOI22_X1   g08528(.A1(new_n8719_), .A2(\asqrt[60] ), .B1(new_n8581_), .B2(new_n8576_), .ZN(new_n8721_));
  OAI22_X1   g08529(.A1(new_n8721_), .A2(new_n229_), .B1(new_n8720_), .B2(new_n8582_), .ZN(new_n8722_));
  NOR4_X1    g08530(.A1(new_n8722_), .A2(\asqrt[62] ), .A3(new_n8718_), .A4(new_n8600_), .ZN(new_n8723_));
  NAND2_X1   g08531(.A1(new_n8723_), .A2(new_n8717_), .ZN(new_n8724_));
  NAND3_X1   g08532(.A1(new_n8313_), .A2(new_n7886_), .A3(new_n7899_), .ZN(new_n8725_));
  NOR3_X1    g08533(.A1(new_n8724_), .A2(new_n8713_), .A3(new_n8725_), .ZN(\asqrt[27] ));
  NAND2_X1   g08534(.A1(new_n8582_), .A2(new_n8591_), .ZN(new_n8727_));
  NOR3_X1    g08535(.A1(new_n8727_), .A2(\asqrt[61] ), .A3(new_n8701_), .ZN(new_n8728_));
  NAND2_X1   g08536(.A1(\asqrt[27] ), .A2(new_n8728_), .ZN(new_n8729_));
  XOR2_X1    g08537(.A1(new_n8729_), .A2(new_n8592_), .Z(new_n8730_));
  INV_X1     g08538(.I(new_n8730_), .ZN(new_n8731_));
  INV_X1     g08539(.I(\a[54] ), .ZN(new_n8732_));
  NOR2_X1    g08540(.A1(\a[52] ), .A2(\a[53] ), .ZN(new_n8733_));
  INV_X1     g08541(.I(new_n8733_), .ZN(new_n8734_));
  NOR3_X1    g08542(.A1(new_n8330_), .A2(new_n8732_), .A3(new_n8734_), .ZN(new_n8735_));
  NAND2_X1   g08543(.A1(new_n8343_), .A2(new_n8735_), .ZN(new_n8736_));
  XOR2_X1    g08544(.A1(new_n8736_), .A2(\a[55] ), .Z(new_n8737_));
  INV_X1     g08545(.I(\a[55] ), .ZN(new_n8738_));
  NOR4_X1    g08546(.A1(new_n8724_), .A2(new_n8713_), .A3(new_n8738_), .A4(new_n8725_), .ZN(new_n8739_));
  NOR2_X1    g08547(.A1(new_n8738_), .A2(\a[54] ), .ZN(new_n8740_));
  OAI21_X1   g08548(.A1(new_n8739_), .A2(new_n8740_), .B(new_n8737_), .ZN(new_n8741_));
  INV_X1     g08549(.I(new_n8737_), .ZN(new_n8742_));
  NOR2_X1    g08550(.A1(new_n8720_), .A2(new_n8582_), .ZN(new_n8743_));
  NOR3_X1    g08551(.A1(new_n8721_), .A2(new_n229_), .A3(new_n8707_), .ZN(new_n8744_));
  AOI21_X1   g08552(.A1(new_n8744_), .A2(new_n8743_), .B(new_n8601_), .ZN(new_n8745_));
  INV_X1     g08553(.I(new_n8712_), .ZN(new_n8746_));
  AOI21_X1   g08554(.A1(new_n8745_), .A2(new_n8746_), .B(new_n8718_), .ZN(new_n8747_));
  AOI21_X1   g08555(.A1(new_n8722_), .A2(\asqrt[62] ), .B(new_n8598_), .ZN(new_n8748_));
  AOI21_X1   g08556(.A1(new_n8694_), .A2(new_n8696_), .B(new_n275_), .ZN(new_n8749_));
  OAI21_X1   g08557(.A1(new_n8697_), .A2(new_n8749_), .B(\asqrt[61] ), .ZN(new_n8750_));
  NAND4_X1   g08558(.A1(new_n8705_), .A2(new_n196_), .A3(new_n8750_), .A4(new_n8706_), .ZN(new_n8751_));
  NOR3_X1    g08559(.A1(new_n8748_), .A2(new_n8716_), .A3(new_n8751_), .ZN(new_n8752_));
  INV_X1     g08560(.I(new_n8725_), .ZN(new_n8753_));
  NAND4_X1   g08561(.A1(new_n8752_), .A2(\a[55] ), .A3(new_n8747_), .A4(new_n8753_), .ZN(new_n8754_));
  NAND3_X1   g08562(.A1(new_n8754_), .A2(\a[54] ), .A3(new_n8742_), .ZN(new_n8755_));
  NAND2_X1   g08563(.A1(new_n8741_), .A2(new_n8755_), .ZN(new_n8756_));
  NOR2_X1    g08564(.A1(new_n8724_), .A2(new_n8713_), .ZN(new_n8757_));
  NAND4_X1   g08565(.A1(new_n8309_), .A2(new_n8301_), .A3(new_n7899_), .A4(new_n8342_), .ZN(new_n8758_));
  NOR2_X1    g08566(.A1(new_n8319_), .A2(new_n8732_), .ZN(new_n8759_));
  XOR2_X1    g08567(.A1(new_n8759_), .A2(new_n8758_), .Z(new_n8760_));
  NOR2_X1    g08568(.A1(new_n8760_), .A2(new_n8734_), .ZN(new_n8761_));
  INV_X1     g08569(.I(new_n8761_), .ZN(new_n8762_));
  NAND3_X1   g08570(.A1(new_n8752_), .A2(new_n8747_), .A3(new_n8753_), .ZN(new_n8763_));
  NOR4_X1    g08571(.A1(new_n8750_), .A2(new_n8582_), .A3(new_n8720_), .A4(new_n8707_), .ZN(new_n8764_));
  NOR3_X1    g08572(.A1(new_n8764_), .A2(new_n8601_), .A3(new_n8712_), .ZN(new_n8765_));
  AOI22_X1   g08573(.A1(new_n8727_), .A2(\asqrt[61] ), .B1(new_n8704_), .B2(new_n8697_), .ZN(new_n8766_));
  NAND4_X1   g08574(.A1(new_n8766_), .A2(new_n196_), .A3(new_n8598_), .A4(new_n8706_), .ZN(new_n8767_));
  OAI21_X1   g08575(.A1(new_n8765_), .A2(new_n8718_), .B(new_n8767_), .ZN(new_n8768_));
  NOR2_X1    g08576(.A1(new_n8717_), .A2(new_n8753_), .ZN(new_n8769_));
  NAND2_X1   g08577(.A1(new_n8769_), .A2(\asqrt[28] ), .ZN(new_n8770_));
  OAI21_X1   g08578(.A1(new_n8768_), .A2(new_n8770_), .B(new_n7865_), .ZN(new_n8771_));
  NAND3_X1   g08579(.A1(new_n8771_), .A2(new_n7873_), .A3(new_n8763_), .ZN(new_n8772_));
  NAND4_X1   g08580(.A1(new_n8592_), .A2(new_n8697_), .A3(new_n8704_), .A4(new_n8708_), .ZN(new_n8773_));
  NAND3_X1   g08581(.A1(new_n8773_), .A2(new_n8602_), .A3(new_n8746_), .ZN(new_n8774_));
  AOI21_X1   g08582(.A1(new_n8598_), .A2(new_n8774_), .B(new_n8723_), .ZN(new_n8775_));
  INV_X1     g08583(.I(new_n8770_), .ZN(new_n8776_));
  AOI21_X1   g08584(.A1(new_n8775_), .A2(new_n8776_), .B(\a[56] ), .ZN(new_n8777_));
  OAI21_X1   g08585(.A1(new_n8777_), .A2(new_n7874_), .B(\asqrt[27] ), .ZN(new_n8778_));
  NAND4_X1   g08586(.A1(new_n8772_), .A2(new_n8778_), .A3(new_n7931_), .A4(new_n8762_), .ZN(new_n8779_));
  NAND2_X1   g08587(.A1(new_n8779_), .A2(new_n8756_), .ZN(new_n8780_));
  NAND3_X1   g08588(.A1(new_n8741_), .A2(new_n8755_), .A3(new_n8762_), .ZN(new_n8781_));
  INV_X1     g08589(.I(new_n7876_), .ZN(new_n8782_));
  NOR2_X1    g08590(.A1(new_n8319_), .A2(\a[56] ), .ZN(new_n8783_));
  OAI22_X1   g08591(.A1(new_n8783_), .A2(\a[57] ), .B1(\a[56] ), .B2(new_n8310_), .ZN(new_n8784_));
  NAND2_X1   g08592(.A1(\asqrt[28] ), .A2(\a[56] ), .ZN(new_n8785_));
  AND3_X2    g08593(.A1(new_n8784_), .A2(new_n8782_), .A3(new_n8785_), .Z(new_n8786_));
  NAND3_X1   g08594(.A1(\asqrt[27] ), .A2(new_n8318_), .A3(new_n8786_), .ZN(new_n8787_));
  INV_X1     g08595(.I(new_n8786_), .ZN(new_n8788_));
  OAI21_X1   g08596(.A1(new_n8763_), .A2(new_n8788_), .B(new_n8317_), .ZN(new_n8789_));
  NAND3_X1   g08597(.A1(new_n8787_), .A2(new_n8789_), .A3(new_n7517_), .ZN(new_n8790_));
  AOI21_X1   g08598(.A1(new_n8781_), .A2(\asqrt[29] ), .B(new_n8790_), .ZN(new_n8791_));
  NOR2_X1    g08599(.A1(new_n8780_), .A2(new_n8791_), .ZN(new_n8792_));
  AOI22_X1   g08600(.A1(new_n8779_), .A2(new_n8756_), .B1(\asqrt[29] ), .B2(new_n8781_), .ZN(new_n8793_));
  INV_X1     g08601(.I(new_n8298_), .ZN(new_n8794_));
  AOI21_X1   g08602(.A1(new_n8310_), .A2(new_n8794_), .B(new_n8300_), .ZN(new_n8795_));
  INV_X1     g08603(.I(new_n8311_), .ZN(new_n8796_));
  NOR3_X1    g08604(.A1(new_n8796_), .A2(new_n8795_), .A3(new_n8317_), .ZN(new_n8797_));
  AOI21_X1   g08605(.A1(new_n8346_), .A2(new_n8333_), .B(\asqrt[30] ), .ZN(new_n8798_));
  AND4_X2    g08606(.A1(new_n8797_), .A2(\asqrt[27] ), .A3(new_n8360_), .A4(new_n8798_), .Z(new_n8799_));
  NOR2_X1    g08607(.A1(new_n8797_), .A2(new_n7517_), .ZN(new_n8800_));
  NOR3_X1    g08608(.A1(new_n8799_), .A2(\asqrt[31] ), .A3(new_n8800_), .ZN(new_n8801_));
  OAI21_X1   g08609(.A1(new_n8793_), .A2(new_n7517_), .B(new_n8801_), .ZN(new_n8802_));
  NAND2_X1   g08610(.A1(new_n8802_), .A2(new_n8792_), .ZN(new_n8803_));
  OAI22_X1   g08611(.A1(new_n8793_), .A2(new_n7517_), .B1(new_n8780_), .B2(new_n8791_), .ZN(new_n8804_));
  NAND2_X1   g08612(.A1(new_n8355_), .A2(new_n8356_), .ZN(new_n8805_));
  NAND4_X1   g08613(.A1(\asqrt[27] ), .A2(new_n7110_), .A3(new_n8805_), .A4(new_n8393_), .ZN(new_n8806_));
  XOR2_X1    g08614(.A1(new_n8806_), .A2(new_n8361_), .Z(new_n8807_));
  NAND2_X1   g08615(.A1(new_n8807_), .A2(new_n6708_), .ZN(new_n8808_));
  AOI21_X1   g08616(.A1(new_n8804_), .A2(\asqrt[31] ), .B(new_n8808_), .ZN(new_n8809_));
  NOR2_X1    g08617(.A1(new_n8809_), .A2(new_n8803_), .ZN(new_n8810_));
  AOI22_X1   g08618(.A1(new_n8804_), .A2(\asqrt[31] ), .B1(new_n8802_), .B2(new_n8792_), .ZN(new_n8811_));
  NOR2_X1    g08619(.A1(new_n8366_), .A2(new_n8367_), .ZN(new_n8812_));
  NOR4_X1    g08620(.A1(new_n8763_), .A2(\asqrt[32] ), .A3(new_n8812_), .A4(new_n8395_), .ZN(new_n8813_));
  XOR2_X1    g08621(.A1(new_n8813_), .A2(new_n8371_), .Z(new_n8814_));
  NAND2_X1   g08622(.A1(new_n8814_), .A2(new_n6365_), .ZN(new_n8815_));
  INV_X1     g08623(.I(new_n8815_), .ZN(new_n8816_));
  OAI21_X1   g08624(.A1(new_n8811_), .A2(new_n6708_), .B(new_n8816_), .ZN(new_n8817_));
  NAND2_X1   g08625(.A1(new_n8817_), .A2(new_n8810_), .ZN(new_n8818_));
  OAI22_X1   g08626(.A1(new_n8811_), .A2(new_n6708_), .B1(new_n8809_), .B2(new_n8803_), .ZN(new_n8819_));
  NOR2_X1    g08627(.A1(new_n8375_), .A2(\asqrt[33] ), .ZN(new_n8820_));
  NAND3_X1   g08628(.A1(\asqrt[27] ), .A2(new_n8396_), .A3(new_n8820_), .ZN(new_n8821_));
  XOR2_X1    g08629(.A1(new_n8821_), .A2(new_n8379_), .Z(new_n8822_));
  NAND2_X1   g08630(.A1(new_n8822_), .A2(new_n5991_), .ZN(new_n8823_));
  AOI21_X1   g08631(.A1(new_n8819_), .A2(\asqrt[33] ), .B(new_n8823_), .ZN(new_n8824_));
  NOR2_X1    g08632(.A1(new_n8824_), .A2(new_n8818_), .ZN(new_n8825_));
  AOI22_X1   g08633(.A1(new_n8819_), .A2(\asqrt[33] ), .B1(new_n8817_), .B2(new_n8810_), .ZN(new_n8826_));
  NOR4_X1    g08634(.A1(new_n8763_), .A2(\asqrt[34] ), .A3(new_n8383_), .A4(new_n8400_), .ZN(new_n8827_));
  XOR2_X1    g08635(.A1(new_n8827_), .A2(new_n8386_), .Z(new_n8828_));
  NAND2_X1   g08636(.A1(new_n8828_), .A2(new_n5626_), .ZN(new_n8829_));
  INV_X1     g08637(.I(new_n8829_), .ZN(new_n8830_));
  OAI21_X1   g08638(.A1(new_n8826_), .A2(new_n5991_), .B(new_n8830_), .ZN(new_n8831_));
  NAND2_X1   g08639(.A1(new_n8831_), .A2(new_n8825_), .ZN(new_n8832_));
  OAI22_X1   g08640(.A1(new_n8826_), .A2(new_n5991_), .B1(new_n8824_), .B2(new_n8818_), .ZN(new_n8833_));
  NOR4_X1    g08641(.A1(new_n8763_), .A2(\asqrt[35] ), .A3(new_n8389_), .A4(new_n8607_), .ZN(new_n8834_));
  XNOR2_X1   g08642(.A1(new_n8834_), .A2(new_n8610_), .ZN(new_n8835_));
  NAND2_X1   g08643(.A1(new_n8835_), .A2(new_n5273_), .ZN(new_n8836_));
  AOI21_X1   g08644(.A1(new_n8833_), .A2(\asqrt[35] ), .B(new_n8836_), .ZN(new_n8837_));
  NOR2_X1    g08645(.A1(new_n8837_), .A2(new_n8832_), .ZN(new_n8838_));
  AOI22_X1   g08646(.A1(new_n8833_), .A2(\asqrt[35] ), .B1(new_n8831_), .B2(new_n8825_), .ZN(new_n8839_));
  NOR4_X1    g08647(.A1(new_n8763_), .A2(\asqrt[36] ), .A3(new_n8404_), .A4(new_n8410_), .ZN(new_n8840_));
  XOR2_X1    g08648(.A1(new_n8840_), .A2(new_n8611_), .Z(new_n8841_));
  NAND2_X1   g08649(.A1(new_n8841_), .A2(new_n4973_), .ZN(new_n8842_));
  INV_X1     g08650(.I(new_n8842_), .ZN(new_n8843_));
  OAI21_X1   g08651(.A1(new_n8839_), .A2(new_n5273_), .B(new_n8843_), .ZN(new_n8844_));
  NAND2_X1   g08652(.A1(new_n8844_), .A2(new_n8838_), .ZN(new_n8845_));
  OAI22_X1   g08653(.A1(new_n8839_), .A2(new_n5273_), .B1(new_n8837_), .B2(new_n8832_), .ZN(new_n8846_));
  NAND2_X1   g08654(.A1(new_n8616_), .A2(\asqrt[37] ), .ZN(new_n8847_));
  NOR4_X1    g08655(.A1(new_n8763_), .A2(\asqrt[37] ), .A3(new_n8413_), .A4(new_n8616_), .ZN(new_n8848_));
  XOR2_X1    g08656(.A1(new_n8848_), .A2(new_n8847_), .Z(new_n8849_));
  NAND2_X1   g08657(.A1(new_n8849_), .A2(new_n4645_), .ZN(new_n8850_));
  AOI21_X1   g08658(.A1(new_n8846_), .A2(\asqrt[37] ), .B(new_n8850_), .ZN(new_n8851_));
  NOR2_X1    g08659(.A1(new_n8851_), .A2(new_n8845_), .ZN(new_n8852_));
  AOI22_X1   g08660(.A1(new_n8846_), .A2(\asqrt[37] ), .B1(new_n8844_), .B2(new_n8838_), .ZN(new_n8853_));
  NOR4_X1    g08661(.A1(new_n8763_), .A2(\asqrt[38] ), .A3(new_n8420_), .A4(new_n8425_), .ZN(new_n8854_));
  AOI21_X1   g08662(.A1(new_n8847_), .A2(new_n8614_), .B(new_n4645_), .ZN(new_n8855_));
  NOR2_X1    g08663(.A1(new_n8854_), .A2(new_n8855_), .ZN(new_n8856_));
  NAND2_X1   g08664(.A1(new_n8856_), .A2(new_n4330_), .ZN(new_n8857_));
  INV_X1     g08665(.I(new_n8857_), .ZN(new_n8858_));
  OAI21_X1   g08666(.A1(new_n8853_), .A2(new_n4645_), .B(new_n8858_), .ZN(new_n8859_));
  NAND2_X1   g08667(.A1(new_n8859_), .A2(new_n8852_), .ZN(new_n8860_));
  OAI22_X1   g08668(.A1(new_n8853_), .A2(new_n4645_), .B1(new_n8851_), .B2(new_n8845_), .ZN(new_n8861_));
  NAND2_X1   g08669(.A1(new_n8623_), .A2(\asqrt[39] ), .ZN(new_n8862_));
  NOR4_X1    g08670(.A1(new_n8763_), .A2(\asqrt[39] ), .A3(new_n8428_), .A4(new_n8623_), .ZN(new_n8863_));
  XOR2_X1    g08671(.A1(new_n8863_), .A2(new_n8862_), .Z(new_n8864_));
  NAND2_X1   g08672(.A1(new_n8864_), .A2(new_n4018_), .ZN(new_n8865_));
  AOI21_X1   g08673(.A1(new_n8861_), .A2(\asqrt[39] ), .B(new_n8865_), .ZN(new_n8866_));
  NOR2_X1    g08674(.A1(new_n8866_), .A2(new_n8860_), .ZN(new_n8867_));
  AOI22_X1   g08675(.A1(new_n8861_), .A2(\asqrt[39] ), .B1(new_n8859_), .B2(new_n8852_), .ZN(new_n8868_));
  NOR4_X1    g08676(.A1(new_n8763_), .A2(\asqrt[40] ), .A3(new_n8435_), .A4(new_n8440_), .ZN(new_n8869_));
  AOI21_X1   g08677(.A1(new_n8862_), .A2(new_n8622_), .B(new_n4018_), .ZN(new_n8870_));
  NOR2_X1    g08678(.A1(new_n8869_), .A2(new_n8870_), .ZN(new_n8871_));
  NAND2_X1   g08679(.A1(new_n8871_), .A2(new_n3760_), .ZN(new_n8872_));
  INV_X1     g08680(.I(new_n8872_), .ZN(new_n8873_));
  OAI21_X1   g08681(.A1(new_n8868_), .A2(new_n4018_), .B(new_n8873_), .ZN(new_n8874_));
  NAND2_X1   g08682(.A1(new_n8874_), .A2(new_n8867_), .ZN(new_n8875_));
  OAI22_X1   g08683(.A1(new_n8868_), .A2(new_n4018_), .B1(new_n8866_), .B2(new_n8860_), .ZN(new_n8876_));
  NAND2_X1   g08684(.A1(new_n8630_), .A2(\asqrt[41] ), .ZN(new_n8877_));
  NOR4_X1    g08685(.A1(new_n8763_), .A2(\asqrt[41] ), .A3(new_n8443_), .A4(new_n8630_), .ZN(new_n8878_));
  XOR2_X1    g08686(.A1(new_n8878_), .A2(new_n8877_), .Z(new_n8879_));
  NAND2_X1   g08687(.A1(new_n8879_), .A2(new_n3481_), .ZN(new_n8880_));
  AOI21_X1   g08688(.A1(new_n8876_), .A2(\asqrt[41] ), .B(new_n8880_), .ZN(new_n8881_));
  NOR2_X1    g08689(.A1(new_n8881_), .A2(new_n8875_), .ZN(new_n8882_));
  AOI22_X1   g08690(.A1(new_n8876_), .A2(\asqrt[41] ), .B1(new_n8874_), .B2(new_n8867_), .ZN(new_n8883_));
  NOR4_X1    g08691(.A1(new_n8763_), .A2(\asqrt[42] ), .A3(new_n8450_), .A4(new_n8455_), .ZN(new_n8884_));
  AOI21_X1   g08692(.A1(new_n8877_), .A2(new_n8629_), .B(new_n3481_), .ZN(new_n8885_));
  NOR2_X1    g08693(.A1(new_n8884_), .A2(new_n8885_), .ZN(new_n8886_));
  NAND2_X1   g08694(.A1(new_n8886_), .A2(new_n3208_), .ZN(new_n8887_));
  INV_X1     g08695(.I(new_n8887_), .ZN(new_n8888_));
  OAI21_X1   g08696(.A1(new_n8883_), .A2(new_n3481_), .B(new_n8888_), .ZN(new_n8889_));
  NAND2_X1   g08697(.A1(new_n8889_), .A2(new_n8882_), .ZN(new_n8890_));
  OAI22_X1   g08698(.A1(new_n8883_), .A2(new_n3481_), .B1(new_n8881_), .B2(new_n8875_), .ZN(new_n8891_));
  NAND2_X1   g08699(.A1(new_n8637_), .A2(\asqrt[43] ), .ZN(new_n8892_));
  NOR4_X1    g08700(.A1(new_n8763_), .A2(\asqrt[43] ), .A3(new_n8458_), .A4(new_n8637_), .ZN(new_n8893_));
  XOR2_X1    g08701(.A1(new_n8893_), .A2(new_n8892_), .Z(new_n8894_));
  NAND2_X1   g08702(.A1(new_n8894_), .A2(new_n2941_), .ZN(new_n8895_));
  AOI21_X1   g08703(.A1(new_n8891_), .A2(\asqrt[43] ), .B(new_n8895_), .ZN(new_n8896_));
  NOR2_X1    g08704(.A1(new_n8896_), .A2(new_n8890_), .ZN(new_n8897_));
  AOI22_X1   g08705(.A1(new_n8891_), .A2(\asqrt[43] ), .B1(new_n8889_), .B2(new_n8882_), .ZN(new_n8898_));
  NOR4_X1    g08706(.A1(new_n8763_), .A2(\asqrt[44] ), .A3(new_n8465_), .A4(new_n8470_), .ZN(new_n8899_));
  AOI21_X1   g08707(.A1(new_n8892_), .A2(new_n8636_), .B(new_n2941_), .ZN(new_n8900_));
  NOR2_X1    g08708(.A1(new_n8899_), .A2(new_n8900_), .ZN(new_n8901_));
  NAND2_X1   g08709(.A1(new_n8901_), .A2(new_n2728_), .ZN(new_n8902_));
  INV_X1     g08710(.I(new_n8902_), .ZN(new_n8903_));
  OAI21_X1   g08711(.A1(new_n8898_), .A2(new_n2941_), .B(new_n8903_), .ZN(new_n8904_));
  NAND2_X1   g08712(.A1(new_n8904_), .A2(new_n8897_), .ZN(new_n8905_));
  OAI22_X1   g08713(.A1(new_n8898_), .A2(new_n2941_), .B1(new_n8896_), .B2(new_n8890_), .ZN(new_n8906_));
  NAND2_X1   g08714(.A1(new_n8644_), .A2(\asqrt[45] ), .ZN(new_n8907_));
  NOR4_X1    g08715(.A1(new_n8763_), .A2(\asqrt[45] ), .A3(new_n8473_), .A4(new_n8644_), .ZN(new_n8908_));
  XOR2_X1    g08716(.A1(new_n8908_), .A2(new_n8907_), .Z(new_n8909_));
  NAND2_X1   g08717(.A1(new_n8909_), .A2(new_n2488_), .ZN(new_n8910_));
  AOI21_X1   g08718(.A1(new_n8906_), .A2(\asqrt[45] ), .B(new_n8910_), .ZN(new_n8911_));
  NOR2_X1    g08719(.A1(new_n8911_), .A2(new_n8905_), .ZN(new_n8912_));
  AOI22_X1   g08720(.A1(new_n8906_), .A2(\asqrt[45] ), .B1(new_n8904_), .B2(new_n8897_), .ZN(new_n8913_));
  NOR4_X1    g08721(.A1(new_n8763_), .A2(\asqrt[46] ), .A3(new_n8480_), .A4(new_n8485_), .ZN(new_n8914_));
  AOI21_X1   g08722(.A1(new_n8907_), .A2(new_n8643_), .B(new_n2488_), .ZN(new_n8915_));
  NOR2_X1    g08723(.A1(new_n8914_), .A2(new_n8915_), .ZN(new_n8916_));
  NAND2_X1   g08724(.A1(new_n8916_), .A2(new_n2253_), .ZN(new_n8917_));
  INV_X1     g08725(.I(new_n8917_), .ZN(new_n8918_));
  OAI21_X1   g08726(.A1(new_n8913_), .A2(new_n2488_), .B(new_n8918_), .ZN(new_n8919_));
  NAND2_X1   g08727(.A1(new_n8919_), .A2(new_n8912_), .ZN(new_n8920_));
  OAI22_X1   g08728(.A1(new_n8913_), .A2(new_n2488_), .B1(new_n8911_), .B2(new_n8905_), .ZN(new_n8921_));
  NAND2_X1   g08729(.A1(new_n8651_), .A2(\asqrt[47] ), .ZN(new_n8922_));
  NOR4_X1    g08730(.A1(new_n8763_), .A2(\asqrt[47] ), .A3(new_n8488_), .A4(new_n8651_), .ZN(new_n8923_));
  XOR2_X1    g08731(.A1(new_n8923_), .A2(new_n8922_), .Z(new_n8924_));
  NAND2_X1   g08732(.A1(new_n8924_), .A2(new_n2046_), .ZN(new_n8925_));
  AOI21_X1   g08733(.A1(new_n8921_), .A2(\asqrt[47] ), .B(new_n8925_), .ZN(new_n8926_));
  NOR2_X1    g08734(.A1(new_n8926_), .A2(new_n8920_), .ZN(new_n8927_));
  AOI22_X1   g08735(.A1(new_n8921_), .A2(\asqrt[47] ), .B1(new_n8919_), .B2(new_n8912_), .ZN(new_n8928_));
  NAND2_X1   g08736(.A1(new_n8500_), .A2(\asqrt[48] ), .ZN(new_n8929_));
  NOR4_X1    g08737(.A1(new_n8763_), .A2(\asqrt[48] ), .A3(new_n8495_), .A4(new_n8500_), .ZN(new_n8930_));
  XOR2_X1    g08738(.A1(new_n8930_), .A2(new_n8929_), .Z(new_n8931_));
  NAND2_X1   g08739(.A1(new_n8931_), .A2(new_n1854_), .ZN(new_n8932_));
  INV_X1     g08740(.I(new_n8932_), .ZN(new_n8933_));
  OAI21_X1   g08741(.A1(new_n8928_), .A2(new_n2046_), .B(new_n8933_), .ZN(new_n8934_));
  NAND2_X1   g08742(.A1(new_n8934_), .A2(new_n8927_), .ZN(new_n8935_));
  OAI22_X1   g08743(.A1(new_n8928_), .A2(new_n2046_), .B1(new_n8926_), .B2(new_n8920_), .ZN(new_n8936_));
  NOR4_X1    g08744(.A1(new_n8763_), .A2(\asqrt[49] ), .A3(new_n8503_), .A4(new_n8658_), .ZN(new_n8937_));
  AOI21_X1   g08745(.A1(new_n8929_), .A2(new_n8499_), .B(new_n1854_), .ZN(new_n8938_));
  NOR2_X1    g08746(.A1(new_n8937_), .A2(new_n8938_), .ZN(new_n8939_));
  NAND2_X1   g08747(.A1(new_n8939_), .A2(new_n1595_), .ZN(new_n8940_));
  AOI21_X1   g08748(.A1(new_n8936_), .A2(\asqrt[49] ), .B(new_n8940_), .ZN(new_n8941_));
  NOR2_X1    g08749(.A1(new_n8941_), .A2(new_n8935_), .ZN(new_n8942_));
  AOI22_X1   g08750(.A1(new_n8936_), .A2(\asqrt[49] ), .B1(new_n8934_), .B2(new_n8927_), .ZN(new_n8943_));
  NAND2_X1   g08751(.A1(new_n8515_), .A2(\asqrt[50] ), .ZN(new_n8944_));
  NOR4_X1    g08752(.A1(new_n8763_), .A2(\asqrt[50] ), .A3(new_n8510_), .A4(new_n8515_), .ZN(new_n8945_));
  XOR2_X1    g08753(.A1(new_n8945_), .A2(new_n8944_), .Z(new_n8946_));
  NAND2_X1   g08754(.A1(new_n8946_), .A2(new_n1436_), .ZN(new_n8947_));
  INV_X1     g08755(.I(new_n8947_), .ZN(new_n8948_));
  OAI21_X1   g08756(.A1(new_n8943_), .A2(new_n1595_), .B(new_n8948_), .ZN(new_n8949_));
  NAND2_X1   g08757(.A1(new_n8949_), .A2(new_n8942_), .ZN(new_n8950_));
  OAI22_X1   g08758(.A1(new_n8943_), .A2(new_n1595_), .B1(new_n8941_), .B2(new_n8935_), .ZN(new_n8951_));
  NOR4_X1    g08759(.A1(new_n8763_), .A2(\asqrt[51] ), .A3(new_n8518_), .A4(new_n8665_), .ZN(new_n8952_));
  AOI21_X1   g08760(.A1(new_n8944_), .A2(new_n8514_), .B(new_n1436_), .ZN(new_n8953_));
  NOR2_X1    g08761(.A1(new_n8952_), .A2(new_n8953_), .ZN(new_n8954_));
  NAND2_X1   g08762(.A1(new_n8954_), .A2(new_n1260_), .ZN(new_n8955_));
  AOI21_X1   g08763(.A1(new_n8951_), .A2(\asqrt[51] ), .B(new_n8955_), .ZN(new_n8956_));
  NOR2_X1    g08764(.A1(new_n8956_), .A2(new_n8950_), .ZN(new_n8957_));
  AOI22_X1   g08765(.A1(new_n8951_), .A2(\asqrt[51] ), .B1(new_n8949_), .B2(new_n8942_), .ZN(new_n8958_));
  NOR4_X1    g08766(.A1(new_n8763_), .A2(\asqrt[52] ), .A3(new_n8525_), .A4(new_n8530_), .ZN(new_n8959_));
  XOR2_X1    g08767(.A1(new_n8959_), .A2(new_n8583_), .Z(new_n8960_));
  NAND2_X1   g08768(.A1(new_n8960_), .A2(new_n1096_), .ZN(new_n8961_));
  INV_X1     g08769(.I(new_n8961_), .ZN(new_n8962_));
  OAI21_X1   g08770(.A1(new_n8958_), .A2(new_n1260_), .B(new_n8962_), .ZN(new_n8963_));
  NAND2_X1   g08771(.A1(new_n8963_), .A2(new_n8957_), .ZN(new_n8964_));
  OAI22_X1   g08772(.A1(new_n8958_), .A2(new_n1260_), .B1(new_n8956_), .B2(new_n8950_), .ZN(new_n8965_));
  NOR4_X1    g08773(.A1(new_n8763_), .A2(\asqrt[53] ), .A3(new_n8533_), .A4(new_n8672_), .ZN(new_n8966_));
  XNOR2_X1   g08774(.A1(new_n8966_), .A2(new_n8584_), .ZN(new_n8967_));
  NAND2_X1   g08775(.A1(new_n8967_), .A2(new_n970_), .ZN(new_n8968_));
  AOI21_X1   g08776(.A1(new_n8965_), .A2(\asqrt[53] ), .B(new_n8968_), .ZN(new_n8969_));
  NOR2_X1    g08777(.A1(new_n8969_), .A2(new_n8964_), .ZN(new_n8970_));
  AOI22_X1   g08778(.A1(new_n8965_), .A2(\asqrt[53] ), .B1(new_n8963_), .B2(new_n8957_), .ZN(new_n8971_));
  NOR4_X1    g08779(.A1(new_n8763_), .A2(\asqrt[54] ), .A3(new_n8540_), .A4(new_n8545_), .ZN(new_n8972_));
  XOR2_X1    g08780(.A1(new_n8972_), .A2(new_n8585_), .Z(new_n8973_));
  NAND2_X1   g08781(.A1(new_n8973_), .A2(new_n825_), .ZN(new_n8974_));
  INV_X1     g08782(.I(new_n8974_), .ZN(new_n8975_));
  OAI21_X1   g08783(.A1(new_n8971_), .A2(new_n970_), .B(new_n8975_), .ZN(new_n8976_));
  NAND2_X1   g08784(.A1(new_n8976_), .A2(new_n8970_), .ZN(new_n8977_));
  OAI22_X1   g08785(.A1(new_n8971_), .A2(new_n970_), .B1(new_n8969_), .B2(new_n8964_), .ZN(new_n8978_));
  NOR4_X1    g08786(.A1(new_n8763_), .A2(\asqrt[55] ), .A3(new_n8548_), .A4(new_n8679_), .ZN(new_n8979_));
  XOR2_X1    g08787(.A1(new_n8979_), .A2(new_n8686_), .Z(new_n8980_));
  NAND2_X1   g08788(.A1(new_n8980_), .A2(new_n724_), .ZN(new_n8981_));
  AOI21_X1   g08789(.A1(new_n8978_), .A2(\asqrt[55] ), .B(new_n8981_), .ZN(new_n8982_));
  NOR2_X1    g08790(.A1(new_n8982_), .A2(new_n8977_), .ZN(new_n8983_));
  AOI22_X1   g08791(.A1(new_n8978_), .A2(\asqrt[55] ), .B1(new_n8976_), .B2(new_n8970_), .ZN(new_n8984_));
  NOR4_X1    g08792(.A1(new_n8763_), .A2(\asqrt[56] ), .A3(new_n8554_), .A4(new_n8559_), .ZN(new_n8985_));
  XOR2_X1    g08793(.A1(new_n8985_), .A2(new_n8587_), .Z(new_n8986_));
  NAND2_X1   g08794(.A1(new_n8986_), .A2(new_n587_), .ZN(new_n8987_));
  INV_X1     g08795(.I(new_n8987_), .ZN(new_n8988_));
  OAI21_X1   g08796(.A1(new_n8984_), .A2(new_n724_), .B(new_n8988_), .ZN(new_n8989_));
  NAND2_X1   g08797(.A1(new_n8989_), .A2(new_n8983_), .ZN(new_n8990_));
  OAI22_X1   g08798(.A1(new_n8984_), .A2(new_n724_), .B1(new_n8982_), .B2(new_n8977_), .ZN(new_n8991_));
  NOR4_X1    g08799(.A1(new_n8763_), .A2(\asqrt[57] ), .A3(new_n8561_), .A4(new_n8690_), .ZN(new_n8992_));
  XOR2_X1    g08800(.A1(new_n8992_), .A2(new_n8688_), .Z(new_n8993_));
  NAND2_X1   g08801(.A1(new_n8993_), .A2(new_n504_), .ZN(new_n8994_));
  AOI21_X1   g08802(.A1(new_n8991_), .A2(\asqrt[57] ), .B(new_n8994_), .ZN(new_n8995_));
  NOR2_X1    g08803(.A1(new_n8995_), .A2(new_n8990_), .ZN(new_n8996_));
  AOI22_X1   g08804(.A1(new_n8991_), .A2(\asqrt[57] ), .B1(new_n8989_), .B2(new_n8983_), .ZN(new_n8997_));
  NOR4_X1    g08805(.A1(new_n8763_), .A2(\asqrt[58] ), .A3(new_n8567_), .A4(new_n8571_), .ZN(new_n8998_));
  XOR2_X1    g08806(.A1(new_n8998_), .A2(new_n8589_), .Z(new_n8999_));
  NAND2_X1   g08807(.A1(new_n8999_), .A2(new_n376_), .ZN(new_n9000_));
  INV_X1     g08808(.I(new_n9000_), .ZN(new_n9001_));
  OAI21_X1   g08809(.A1(new_n8997_), .A2(new_n504_), .B(new_n9001_), .ZN(new_n9002_));
  NAND2_X1   g08810(.A1(new_n9002_), .A2(new_n8996_), .ZN(new_n9003_));
  OAI22_X1   g08811(.A1(new_n8997_), .A2(new_n504_), .B1(new_n8995_), .B2(new_n8990_), .ZN(new_n9004_));
  NOR4_X1    g08812(.A1(new_n8763_), .A2(\asqrt[59] ), .A3(new_n8573_), .A4(new_n8698_), .ZN(new_n9005_));
  XOR2_X1    g08813(.A1(new_n9005_), .A2(new_n8696_), .Z(new_n9006_));
  NAND2_X1   g08814(.A1(new_n9006_), .A2(new_n275_), .ZN(new_n9007_));
  AOI21_X1   g08815(.A1(new_n9004_), .A2(\asqrt[59] ), .B(new_n9007_), .ZN(new_n9008_));
  NOR2_X1    g08816(.A1(new_n9008_), .A2(new_n9003_), .ZN(new_n9009_));
  AOI22_X1   g08817(.A1(new_n9004_), .A2(\asqrt[59] ), .B1(new_n9002_), .B2(new_n8996_), .ZN(new_n9010_));
  OAI22_X1   g08818(.A1(new_n9010_), .A2(new_n275_), .B1(new_n9008_), .B2(new_n9003_), .ZN(new_n9011_));
  NOR4_X1    g08819(.A1(new_n8763_), .A2(\asqrt[60] ), .A3(new_n8579_), .A4(new_n8719_), .ZN(new_n9012_));
  XOR2_X1    g08820(.A1(new_n9012_), .A2(new_n8591_), .Z(new_n9013_));
  NAND2_X1   g08821(.A1(new_n9013_), .A2(new_n229_), .ZN(new_n9014_));
  INV_X1     g08822(.I(new_n9014_), .ZN(new_n9015_));
  OAI21_X1   g08823(.A1(new_n9010_), .A2(new_n275_), .B(new_n9015_), .ZN(new_n9016_));
  AOI22_X1   g08824(.A1(new_n9011_), .A2(\asqrt[61] ), .B1(new_n9016_), .B2(new_n9009_), .ZN(new_n9017_));
  NOR2_X1    g08825(.A1(new_n9017_), .A2(new_n196_), .ZN(new_n9018_));
  INV_X1     g08826(.I(new_n8740_), .ZN(new_n9019_));
  AOI21_X1   g08827(.A1(new_n8754_), .A2(new_n9019_), .B(new_n8742_), .ZN(new_n9020_));
  NOR3_X1    g08828(.A1(new_n8739_), .A2(new_n8732_), .A3(new_n8737_), .ZN(new_n9021_));
  NOR2_X1    g08829(.A1(new_n9021_), .A2(new_n9020_), .ZN(new_n9022_));
  NOR3_X1    g08830(.A1(new_n8777_), .A2(new_n7874_), .A3(\asqrt[27] ), .ZN(new_n9023_));
  AOI21_X1   g08831(.A1(new_n8771_), .A2(new_n7873_), .B(new_n8763_), .ZN(new_n9024_));
  NOR4_X1    g08832(.A1(new_n9024_), .A2(new_n9023_), .A3(\asqrt[29] ), .A4(new_n8761_), .ZN(new_n9025_));
  NOR2_X1    g08833(.A1(new_n9025_), .A2(new_n9022_), .ZN(new_n9026_));
  NOR3_X1    g08834(.A1(new_n9021_), .A2(new_n9020_), .A3(new_n8761_), .ZN(new_n9027_));
  NOR3_X1    g08835(.A1(new_n8763_), .A2(new_n8317_), .A3(new_n8788_), .ZN(new_n9028_));
  AOI21_X1   g08836(.A1(\asqrt[27] ), .A2(new_n8786_), .B(new_n8318_), .ZN(new_n9029_));
  NOR3_X1    g08837(.A1(new_n9029_), .A2(new_n9028_), .A3(\asqrt[30] ), .ZN(new_n9030_));
  OAI21_X1   g08838(.A1(new_n9027_), .A2(new_n7931_), .B(new_n9030_), .ZN(new_n9031_));
  NAND2_X1   g08839(.A1(new_n9026_), .A2(new_n9031_), .ZN(new_n9032_));
  OAI22_X1   g08840(.A1(new_n9025_), .A2(new_n9022_), .B1(new_n7931_), .B2(new_n9027_), .ZN(new_n9033_));
  INV_X1     g08841(.I(new_n8801_), .ZN(new_n9034_));
  AOI21_X1   g08842(.A1(new_n9033_), .A2(\asqrt[30] ), .B(new_n9034_), .ZN(new_n9035_));
  NOR2_X1    g08843(.A1(new_n9035_), .A2(new_n9032_), .ZN(new_n9036_));
  AOI22_X1   g08844(.A1(new_n9033_), .A2(\asqrt[30] ), .B1(new_n9026_), .B2(new_n9031_), .ZN(new_n9037_));
  INV_X1     g08845(.I(new_n8808_), .ZN(new_n9038_));
  OAI21_X1   g08846(.A1(new_n9037_), .A2(new_n7110_), .B(new_n9038_), .ZN(new_n9039_));
  NAND2_X1   g08847(.A1(new_n9039_), .A2(new_n9036_), .ZN(new_n9040_));
  OAI22_X1   g08848(.A1(new_n9037_), .A2(new_n7110_), .B1(new_n9035_), .B2(new_n9032_), .ZN(new_n9041_));
  AOI21_X1   g08849(.A1(new_n9041_), .A2(\asqrt[32] ), .B(new_n8815_), .ZN(new_n9042_));
  NOR2_X1    g08850(.A1(new_n9042_), .A2(new_n9040_), .ZN(new_n9043_));
  AOI22_X1   g08851(.A1(new_n9041_), .A2(\asqrt[32] ), .B1(new_n9039_), .B2(new_n9036_), .ZN(new_n9044_));
  INV_X1     g08852(.I(new_n8823_), .ZN(new_n9045_));
  OAI21_X1   g08853(.A1(new_n9044_), .A2(new_n6365_), .B(new_n9045_), .ZN(new_n9046_));
  NAND2_X1   g08854(.A1(new_n9046_), .A2(new_n9043_), .ZN(new_n9047_));
  OAI22_X1   g08855(.A1(new_n9044_), .A2(new_n6365_), .B1(new_n9042_), .B2(new_n9040_), .ZN(new_n9048_));
  AOI21_X1   g08856(.A1(new_n9048_), .A2(\asqrt[34] ), .B(new_n8829_), .ZN(new_n9049_));
  NOR2_X1    g08857(.A1(new_n9049_), .A2(new_n9047_), .ZN(new_n9050_));
  AOI22_X1   g08858(.A1(new_n9048_), .A2(\asqrt[34] ), .B1(new_n9046_), .B2(new_n9043_), .ZN(new_n9051_));
  INV_X1     g08859(.I(new_n8836_), .ZN(new_n9052_));
  OAI21_X1   g08860(.A1(new_n9051_), .A2(new_n5626_), .B(new_n9052_), .ZN(new_n9053_));
  NAND2_X1   g08861(.A1(new_n9053_), .A2(new_n9050_), .ZN(new_n9054_));
  OAI22_X1   g08862(.A1(new_n9051_), .A2(new_n5626_), .B1(new_n9049_), .B2(new_n9047_), .ZN(new_n9055_));
  AOI21_X1   g08863(.A1(new_n9055_), .A2(\asqrt[36] ), .B(new_n8842_), .ZN(new_n9056_));
  NOR2_X1    g08864(.A1(new_n9056_), .A2(new_n9054_), .ZN(new_n9057_));
  AOI22_X1   g08865(.A1(new_n9055_), .A2(\asqrt[36] ), .B1(new_n9053_), .B2(new_n9050_), .ZN(new_n9058_));
  INV_X1     g08866(.I(new_n8850_), .ZN(new_n9059_));
  OAI21_X1   g08867(.A1(new_n9058_), .A2(new_n4973_), .B(new_n9059_), .ZN(new_n9060_));
  NAND2_X1   g08868(.A1(new_n9060_), .A2(new_n9057_), .ZN(new_n9061_));
  OAI22_X1   g08869(.A1(new_n9058_), .A2(new_n4973_), .B1(new_n9056_), .B2(new_n9054_), .ZN(new_n9062_));
  AOI21_X1   g08870(.A1(new_n9062_), .A2(\asqrt[38] ), .B(new_n8857_), .ZN(new_n9063_));
  NOR2_X1    g08871(.A1(new_n9063_), .A2(new_n9061_), .ZN(new_n9064_));
  AOI22_X1   g08872(.A1(new_n9062_), .A2(\asqrt[38] ), .B1(new_n9060_), .B2(new_n9057_), .ZN(new_n9065_));
  INV_X1     g08873(.I(new_n8865_), .ZN(new_n9066_));
  OAI21_X1   g08874(.A1(new_n9065_), .A2(new_n4330_), .B(new_n9066_), .ZN(new_n9067_));
  NAND2_X1   g08875(.A1(new_n9067_), .A2(new_n9064_), .ZN(new_n9068_));
  OAI22_X1   g08876(.A1(new_n9065_), .A2(new_n4330_), .B1(new_n9063_), .B2(new_n9061_), .ZN(new_n9069_));
  AOI21_X1   g08877(.A1(new_n9069_), .A2(\asqrt[40] ), .B(new_n8872_), .ZN(new_n9070_));
  NOR2_X1    g08878(.A1(new_n9070_), .A2(new_n9068_), .ZN(new_n9071_));
  AOI22_X1   g08879(.A1(new_n9069_), .A2(\asqrt[40] ), .B1(new_n9067_), .B2(new_n9064_), .ZN(new_n9072_));
  INV_X1     g08880(.I(new_n8880_), .ZN(new_n9073_));
  OAI21_X1   g08881(.A1(new_n9072_), .A2(new_n3760_), .B(new_n9073_), .ZN(new_n9074_));
  NAND2_X1   g08882(.A1(new_n9074_), .A2(new_n9071_), .ZN(new_n9075_));
  OAI22_X1   g08883(.A1(new_n9072_), .A2(new_n3760_), .B1(new_n9070_), .B2(new_n9068_), .ZN(new_n9076_));
  AOI21_X1   g08884(.A1(new_n9076_), .A2(\asqrt[42] ), .B(new_n8887_), .ZN(new_n9077_));
  NOR2_X1    g08885(.A1(new_n9077_), .A2(new_n9075_), .ZN(new_n9078_));
  AOI22_X1   g08886(.A1(new_n9076_), .A2(\asqrt[42] ), .B1(new_n9074_), .B2(new_n9071_), .ZN(new_n9079_));
  INV_X1     g08887(.I(new_n8895_), .ZN(new_n9080_));
  OAI21_X1   g08888(.A1(new_n9079_), .A2(new_n3208_), .B(new_n9080_), .ZN(new_n9081_));
  NAND2_X1   g08889(.A1(new_n9081_), .A2(new_n9078_), .ZN(new_n9082_));
  OAI22_X1   g08890(.A1(new_n9079_), .A2(new_n3208_), .B1(new_n9077_), .B2(new_n9075_), .ZN(new_n9083_));
  AOI21_X1   g08891(.A1(new_n9083_), .A2(\asqrt[44] ), .B(new_n8902_), .ZN(new_n9084_));
  NOR2_X1    g08892(.A1(new_n9084_), .A2(new_n9082_), .ZN(new_n9085_));
  AOI22_X1   g08893(.A1(new_n9083_), .A2(\asqrt[44] ), .B1(new_n9081_), .B2(new_n9078_), .ZN(new_n9086_));
  INV_X1     g08894(.I(new_n8910_), .ZN(new_n9087_));
  OAI21_X1   g08895(.A1(new_n9086_), .A2(new_n2728_), .B(new_n9087_), .ZN(new_n9088_));
  NAND2_X1   g08896(.A1(new_n9088_), .A2(new_n9085_), .ZN(new_n9089_));
  OAI22_X1   g08897(.A1(new_n9086_), .A2(new_n2728_), .B1(new_n9084_), .B2(new_n9082_), .ZN(new_n9090_));
  AOI21_X1   g08898(.A1(new_n9090_), .A2(\asqrt[46] ), .B(new_n8917_), .ZN(new_n9091_));
  NOR2_X1    g08899(.A1(new_n9091_), .A2(new_n9089_), .ZN(new_n9092_));
  AOI22_X1   g08900(.A1(new_n9090_), .A2(\asqrt[46] ), .B1(new_n9088_), .B2(new_n9085_), .ZN(new_n9093_));
  INV_X1     g08901(.I(new_n8925_), .ZN(new_n9094_));
  OAI21_X1   g08902(.A1(new_n9093_), .A2(new_n2253_), .B(new_n9094_), .ZN(new_n9095_));
  NAND2_X1   g08903(.A1(new_n9095_), .A2(new_n9092_), .ZN(new_n9096_));
  OAI22_X1   g08904(.A1(new_n9093_), .A2(new_n2253_), .B1(new_n9091_), .B2(new_n9089_), .ZN(new_n9097_));
  AOI21_X1   g08905(.A1(new_n9097_), .A2(\asqrt[48] ), .B(new_n8932_), .ZN(new_n9098_));
  NOR2_X1    g08906(.A1(new_n9098_), .A2(new_n9096_), .ZN(new_n9099_));
  AOI22_X1   g08907(.A1(new_n9097_), .A2(\asqrt[48] ), .B1(new_n9095_), .B2(new_n9092_), .ZN(new_n9100_));
  INV_X1     g08908(.I(new_n8940_), .ZN(new_n9101_));
  OAI21_X1   g08909(.A1(new_n9100_), .A2(new_n1854_), .B(new_n9101_), .ZN(new_n9102_));
  NAND2_X1   g08910(.A1(new_n9102_), .A2(new_n9099_), .ZN(new_n9103_));
  OAI22_X1   g08911(.A1(new_n9100_), .A2(new_n1854_), .B1(new_n9098_), .B2(new_n9096_), .ZN(new_n9104_));
  AOI21_X1   g08912(.A1(new_n9104_), .A2(\asqrt[50] ), .B(new_n8947_), .ZN(new_n9105_));
  NOR2_X1    g08913(.A1(new_n9105_), .A2(new_n9103_), .ZN(new_n9106_));
  AOI22_X1   g08914(.A1(new_n9104_), .A2(\asqrt[50] ), .B1(new_n9102_), .B2(new_n9099_), .ZN(new_n9107_));
  INV_X1     g08915(.I(new_n8955_), .ZN(new_n9108_));
  OAI21_X1   g08916(.A1(new_n9107_), .A2(new_n1436_), .B(new_n9108_), .ZN(new_n9109_));
  NAND2_X1   g08917(.A1(new_n9109_), .A2(new_n9106_), .ZN(new_n9110_));
  OAI22_X1   g08918(.A1(new_n9107_), .A2(new_n1436_), .B1(new_n9105_), .B2(new_n9103_), .ZN(new_n9111_));
  AOI21_X1   g08919(.A1(new_n9111_), .A2(\asqrt[52] ), .B(new_n8961_), .ZN(new_n9112_));
  NOR2_X1    g08920(.A1(new_n9112_), .A2(new_n9110_), .ZN(new_n9113_));
  AOI22_X1   g08921(.A1(new_n9111_), .A2(\asqrt[52] ), .B1(new_n9109_), .B2(new_n9106_), .ZN(new_n9114_));
  INV_X1     g08922(.I(new_n8968_), .ZN(new_n9115_));
  OAI21_X1   g08923(.A1(new_n9114_), .A2(new_n1096_), .B(new_n9115_), .ZN(new_n9116_));
  NAND2_X1   g08924(.A1(new_n9116_), .A2(new_n9113_), .ZN(new_n9117_));
  OAI22_X1   g08925(.A1(new_n9114_), .A2(new_n1096_), .B1(new_n9112_), .B2(new_n9110_), .ZN(new_n9118_));
  AOI21_X1   g08926(.A1(new_n9118_), .A2(\asqrt[54] ), .B(new_n8974_), .ZN(new_n9119_));
  NOR2_X1    g08927(.A1(new_n9119_), .A2(new_n9117_), .ZN(new_n9120_));
  AOI22_X1   g08928(.A1(new_n9118_), .A2(\asqrt[54] ), .B1(new_n9116_), .B2(new_n9113_), .ZN(new_n9121_));
  INV_X1     g08929(.I(new_n8981_), .ZN(new_n9122_));
  OAI21_X1   g08930(.A1(new_n9121_), .A2(new_n825_), .B(new_n9122_), .ZN(new_n9123_));
  NAND2_X1   g08931(.A1(new_n9123_), .A2(new_n9120_), .ZN(new_n9124_));
  OAI22_X1   g08932(.A1(new_n9121_), .A2(new_n825_), .B1(new_n9119_), .B2(new_n9117_), .ZN(new_n9125_));
  AOI21_X1   g08933(.A1(new_n9125_), .A2(\asqrt[56] ), .B(new_n8987_), .ZN(new_n9126_));
  NOR2_X1    g08934(.A1(new_n9126_), .A2(new_n9124_), .ZN(new_n9127_));
  AOI22_X1   g08935(.A1(new_n9125_), .A2(\asqrt[56] ), .B1(new_n9123_), .B2(new_n9120_), .ZN(new_n9128_));
  INV_X1     g08936(.I(new_n8994_), .ZN(new_n9129_));
  OAI21_X1   g08937(.A1(new_n9128_), .A2(new_n587_), .B(new_n9129_), .ZN(new_n9130_));
  NAND2_X1   g08938(.A1(new_n9130_), .A2(new_n9127_), .ZN(new_n9131_));
  OAI22_X1   g08939(.A1(new_n9128_), .A2(new_n587_), .B1(new_n9126_), .B2(new_n9124_), .ZN(new_n9132_));
  AOI21_X1   g08940(.A1(new_n9132_), .A2(\asqrt[58] ), .B(new_n9000_), .ZN(new_n9133_));
  NOR2_X1    g08941(.A1(new_n9133_), .A2(new_n9131_), .ZN(new_n9134_));
  AOI22_X1   g08942(.A1(new_n9132_), .A2(\asqrt[58] ), .B1(new_n9130_), .B2(new_n9127_), .ZN(new_n9135_));
  INV_X1     g08943(.I(new_n9007_), .ZN(new_n9136_));
  OAI21_X1   g08944(.A1(new_n9135_), .A2(new_n376_), .B(new_n9136_), .ZN(new_n9137_));
  NAND2_X1   g08945(.A1(new_n9137_), .A2(new_n9134_), .ZN(new_n9138_));
  OAI22_X1   g08946(.A1(new_n9135_), .A2(new_n376_), .B1(new_n9133_), .B2(new_n9131_), .ZN(new_n9139_));
  AOI22_X1   g08947(.A1(new_n9139_), .A2(\asqrt[60] ), .B1(new_n9137_), .B2(new_n9134_), .ZN(new_n9140_));
  AOI21_X1   g08948(.A1(new_n9139_), .A2(\asqrt[60] ), .B(new_n9014_), .ZN(new_n9141_));
  OAI22_X1   g08949(.A1(new_n9140_), .A2(new_n229_), .B1(new_n9141_), .B2(new_n9138_), .ZN(new_n9142_));
  NOR2_X1    g08950(.A1(new_n9142_), .A2(\asqrt[62] ), .ZN(new_n9143_));
  NAND3_X1   g08951(.A1(new_n8757_), .A2(new_n8598_), .A3(new_n8725_), .ZN(new_n9144_));
  NOR2_X1    g08952(.A1(new_n8766_), .A2(new_n196_), .ZN(new_n9145_));
  INV_X1     g08953(.I(new_n8751_), .ZN(new_n9146_));
  NAND3_X1   g08954(.A1(\asqrt[27] ), .A2(new_n9145_), .A3(new_n9146_), .ZN(new_n9147_));
  OAI21_X1   g08955(.A1(new_n8722_), .A2(\asqrt[62] ), .B(new_n8600_), .ZN(new_n9148_));
  OAI21_X1   g08956(.A1(\asqrt[27] ), .A2(new_n9148_), .B(new_n9145_), .ZN(new_n9149_));
  NAND2_X1   g08957(.A1(new_n9149_), .A2(new_n9147_), .ZN(new_n9150_));
  INV_X1     g08958(.I(new_n9150_), .ZN(new_n9151_));
  NOR2_X1    g08959(.A1(new_n8730_), .A2(new_n196_), .ZN(new_n9152_));
  INV_X1     g08960(.I(new_n9152_), .ZN(new_n9153_));
  NAND2_X1   g08961(.A1(new_n9004_), .A2(\asqrt[59] ), .ZN(new_n9154_));
  AOI21_X1   g08962(.A1(new_n9154_), .A2(new_n9003_), .B(new_n275_), .ZN(new_n9155_));
  OAI21_X1   g08963(.A1(new_n9009_), .A2(new_n9155_), .B(\asqrt[61] ), .ZN(new_n9156_));
  NOR2_X1    g08964(.A1(new_n8731_), .A2(\asqrt[62] ), .ZN(new_n9157_));
  INV_X1     g08965(.I(new_n9157_), .ZN(new_n9158_));
  NAND3_X1   g08966(.A1(new_n9016_), .A2(new_n9009_), .A3(new_n9158_), .ZN(new_n9159_));
  OAI21_X1   g08967(.A1(new_n9159_), .A2(new_n9156_), .B(new_n9153_), .ZN(new_n9160_));
  NAND3_X1   g08968(.A1(new_n8763_), .A2(new_n8718_), .A3(new_n8767_), .ZN(new_n9161_));
  AOI21_X1   g08969(.A1(new_n9161_), .A2(new_n8710_), .B(\asqrt[63] ), .ZN(new_n9162_));
  INV_X1     g08970(.I(new_n9162_), .ZN(new_n9163_));
  OAI21_X1   g08971(.A1(new_n9160_), .A2(new_n9163_), .B(new_n9151_), .ZN(new_n9164_));
  NOR4_X1    g08972(.A1(new_n9142_), .A2(\asqrt[62] ), .A3(new_n9150_), .A4(new_n8730_), .ZN(new_n9165_));
  NAND2_X1   g08973(.A1(new_n8745_), .A2(new_n8718_), .ZN(new_n9166_));
  XOR2_X1    g08974(.A1(new_n8745_), .A2(\asqrt[63] ), .Z(new_n9167_));
  AOI21_X1   g08975(.A1(\asqrt[27] ), .A2(new_n9166_), .B(new_n9167_), .ZN(new_n9168_));
  NAND2_X1   g08976(.A1(new_n9165_), .A2(new_n9168_), .ZN(new_n9169_));
  NOR3_X1    g08977(.A1(new_n9169_), .A2(new_n9144_), .A3(new_n9164_), .ZN(\asqrt[26] ));
  NAND4_X1   g08978(.A1(\asqrt[26] ), .A2(new_n8731_), .A3(new_n9018_), .A4(new_n9143_), .ZN(new_n9171_));
  OAI21_X1   g08979(.A1(new_n9142_), .A2(\asqrt[62] ), .B(new_n8730_), .ZN(new_n9172_));
  OAI21_X1   g08980(.A1(\asqrt[26] ), .A2(new_n9172_), .B(new_n9018_), .ZN(new_n9173_));
  NAND2_X1   g08981(.A1(new_n9171_), .A2(new_n9173_), .ZN(new_n9174_));
  INV_X1     g08982(.I(new_n9174_), .ZN(new_n9175_));
  NAND2_X1   g08983(.A1(new_n9132_), .A2(\asqrt[58] ), .ZN(new_n9176_));
  AOI21_X1   g08984(.A1(new_n9176_), .A2(new_n9131_), .B(new_n376_), .ZN(new_n9177_));
  OAI21_X1   g08985(.A1(new_n9134_), .A2(new_n9177_), .B(\asqrt[60] ), .ZN(new_n9178_));
  AOI21_X1   g08986(.A1(new_n9138_), .A2(new_n9178_), .B(new_n229_), .ZN(new_n9179_));
  NOR3_X1    g08987(.A1(new_n9011_), .A2(\asqrt[61] ), .A3(new_n9013_), .ZN(new_n9180_));
  NAND2_X1   g08988(.A1(\asqrt[26] ), .A2(new_n9180_), .ZN(new_n9181_));
  XOR2_X1    g08989(.A1(new_n9181_), .A2(new_n9179_), .Z(new_n9182_));
  NOR2_X1    g08990(.A1(new_n9182_), .A2(new_n196_), .ZN(new_n9183_));
  INV_X1     g08991(.I(new_n9183_), .ZN(new_n9184_));
  INV_X1     g08992(.I(\a[52] ), .ZN(new_n9185_));
  NOR2_X1    g08993(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n9186_));
  INV_X1     g08994(.I(new_n9186_), .ZN(new_n9187_));
  NOR3_X1    g08995(.A1(new_n8769_), .A2(new_n9185_), .A3(new_n9187_), .ZN(new_n9188_));
  NAND2_X1   g08996(.A1(new_n8775_), .A2(new_n9188_), .ZN(new_n9189_));
  XOR2_X1    g08997(.A1(new_n9189_), .A2(\a[53] ), .Z(new_n9190_));
  INV_X1     g08998(.I(\a[53] ), .ZN(new_n9191_));
  NOR4_X1    g08999(.A1(new_n9169_), .A2(new_n9191_), .A3(new_n9144_), .A4(new_n9164_), .ZN(new_n9192_));
  NOR2_X1    g09000(.A1(new_n9191_), .A2(\a[52] ), .ZN(new_n9193_));
  OAI21_X1   g09001(.A1(new_n9192_), .A2(new_n9193_), .B(new_n9190_), .ZN(new_n9194_));
  INV_X1     g09002(.I(new_n9190_), .ZN(new_n9195_));
  INV_X1     g09003(.I(new_n9144_), .ZN(new_n9196_));
  NOR3_X1    g09004(.A1(new_n9141_), .A2(new_n9138_), .A3(new_n9157_), .ZN(new_n9197_));
  AOI21_X1   g09005(.A1(new_n9197_), .A2(new_n9179_), .B(new_n9152_), .ZN(new_n9198_));
  AOI21_X1   g09006(.A1(new_n9198_), .A2(new_n9162_), .B(new_n9150_), .ZN(new_n9199_));
  NAND4_X1   g09007(.A1(new_n9017_), .A2(new_n196_), .A3(new_n9151_), .A4(new_n8731_), .ZN(new_n9200_));
  INV_X1     g09008(.I(new_n9168_), .ZN(new_n9201_));
  NOR2_X1    g09009(.A1(new_n9200_), .A2(new_n9201_), .ZN(new_n9202_));
  NAND4_X1   g09010(.A1(new_n9202_), .A2(\a[53] ), .A3(new_n9199_), .A4(new_n9196_), .ZN(new_n9203_));
  NAND3_X1   g09011(.A1(new_n9203_), .A2(\a[52] ), .A3(new_n9195_), .ZN(new_n9204_));
  NAND2_X1   g09012(.A1(new_n9194_), .A2(new_n9204_), .ZN(new_n9205_));
  NOR2_X1    g09013(.A1(new_n9169_), .A2(new_n9164_), .ZN(new_n9206_));
  NOR4_X1    g09014(.A1(new_n8724_), .A2(new_n8718_), .A3(new_n8765_), .A4(new_n8725_), .ZN(new_n9207_));
  NAND2_X1   g09015(.A1(\asqrt[27] ), .A2(\a[52] ), .ZN(new_n9208_));
  XOR2_X1    g09016(.A1(new_n9208_), .A2(new_n9207_), .Z(new_n9209_));
  NOR2_X1    g09017(.A1(new_n9209_), .A2(new_n9187_), .ZN(new_n9210_));
  INV_X1     g09018(.I(new_n9210_), .ZN(new_n9211_));
  NAND3_X1   g09019(.A1(new_n9202_), .A2(new_n9196_), .A3(new_n9199_), .ZN(new_n9212_));
  NOR2_X1    g09020(.A1(new_n9196_), .A2(new_n9168_), .ZN(new_n9213_));
  NAND2_X1   g09021(.A1(new_n9213_), .A2(\asqrt[27] ), .ZN(new_n9214_));
  INV_X1     g09022(.I(new_n9214_), .ZN(new_n9215_));
  NAND3_X1   g09023(.A1(new_n9164_), .A2(new_n9200_), .A3(new_n9215_), .ZN(new_n9216_));
  NAND2_X1   g09024(.A1(new_n9216_), .A2(new_n8732_), .ZN(new_n9217_));
  NAND3_X1   g09025(.A1(new_n9217_), .A2(new_n8733_), .A3(new_n9212_), .ZN(new_n9218_));
  NOR3_X1    g09026(.A1(new_n9199_), .A2(new_n9165_), .A3(new_n9214_), .ZN(new_n9219_));
  OAI21_X1   g09027(.A1(new_n9219_), .A2(\a[54] ), .B(new_n8733_), .ZN(new_n9220_));
  NAND2_X1   g09028(.A1(new_n9220_), .A2(\asqrt[26] ), .ZN(new_n9221_));
  NAND4_X1   g09029(.A1(new_n9221_), .A2(new_n8319_), .A3(new_n9218_), .A4(new_n9211_), .ZN(new_n9222_));
  NAND2_X1   g09030(.A1(new_n9222_), .A2(new_n9205_), .ZN(new_n9223_));
  NAND3_X1   g09031(.A1(new_n9194_), .A2(new_n9204_), .A3(new_n9211_), .ZN(new_n9224_));
  AOI21_X1   g09032(.A1(\asqrt[27] ), .A2(new_n8732_), .B(\a[55] ), .ZN(new_n9225_));
  NOR2_X1    g09033(.A1(new_n8754_), .A2(\a[54] ), .ZN(new_n9226_));
  AOI21_X1   g09034(.A1(\asqrt[27] ), .A2(\a[54] ), .B(new_n8736_), .ZN(new_n9227_));
  OAI21_X1   g09035(.A1(new_n9226_), .A2(new_n9225_), .B(new_n9227_), .ZN(new_n9228_));
  INV_X1     g09036(.I(new_n9228_), .ZN(new_n9229_));
  NAND3_X1   g09037(.A1(\asqrt[26] ), .A2(new_n8762_), .A3(new_n9229_), .ZN(new_n9230_));
  OAI21_X1   g09038(.A1(new_n9212_), .A2(new_n9228_), .B(new_n8761_), .ZN(new_n9231_));
  NAND3_X1   g09039(.A1(new_n9230_), .A2(new_n9231_), .A3(new_n7931_), .ZN(new_n9232_));
  AOI21_X1   g09040(.A1(new_n9224_), .A2(\asqrt[28] ), .B(new_n9232_), .ZN(new_n9233_));
  NOR2_X1    g09041(.A1(new_n9223_), .A2(new_n9233_), .ZN(new_n9234_));
  NAND2_X1   g09042(.A1(new_n9224_), .A2(\asqrt[28] ), .ZN(new_n9235_));
  AOI21_X1   g09043(.A1(new_n9223_), .A2(new_n9235_), .B(new_n7931_), .ZN(new_n9236_));
  NOR2_X1    g09044(.A1(new_n9024_), .A2(new_n9023_), .ZN(new_n9237_));
  NOR4_X1    g09045(.A1(new_n9212_), .A2(\asqrt[29] ), .A3(new_n9237_), .A4(new_n8781_), .ZN(new_n9238_));
  AOI21_X1   g09046(.A1(new_n9022_), .A2(new_n8762_), .B(new_n7931_), .ZN(new_n9239_));
  NOR2_X1    g09047(.A1(new_n9238_), .A2(new_n9239_), .ZN(new_n9240_));
  NAND2_X1   g09048(.A1(new_n9240_), .A2(new_n7517_), .ZN(new_n9241_));
  OAI21_X1   g09049(.A1(new_n9236_), .A2(new_n9241_), .B(new_n9234_), .ZN(new_n9242_));
  AOI22_X1   g09050(.A1(new_n9222_), .A2(new_n9205_), .B1(\asqrt[28] ), .B2(new_n9224_), .ZN(new_n9243_));
  OAI22_X1   g09051(.A1(new_n9243_), .A2(new_n7931_), .B1(new_n9223_), .B2(new_n9233_), .ZN(new_n9244_));
  NOR2_X1    g09052(.A1(new_n8793_), .A2(new_n7517_), .ZN(new_n9245_));
  NAND2_X1   g09053(.A1(new_n8787_), .A2(new_n8789_), .ZN(new_n9246_));
  NAND4_X1   g09054(.A1(\asqrt[26] ), .A2(new_n7517_), .A3(new_n9246_), .A4(new_n8793_), .ZN(new_n9247_));
  XOR2_X1    g09055(.A1(new_n9247_), .A2(new_n9245_), .Z(new_n9248_));
  NAND2_X1   g09056(.A1(new_n9248_), .A2(new_n7110_), .ZN(new_n9249_));
  AOI21_X1   g09057(.A1(new_n9244_), .A2(\asqrt[30] ), .B(new_n9249_), .ZN(new_n9250_));
  OAI21_X1   g09058(.A1(new_n9236_), .A2(new_n9234_), .B(\asqrt[30] ), .ZN(new_n9251_));
  AOI21_X1   g09059(.A1(new_n9242_), .A2(new_n9251_), .B(new_n7110_), .ZN(new_n9252_));
  NAND2_X1   g09060(.A1(new_n8804_), .A2(\asqrt[31] ), .ZN(new_n9253_));
  NOR2_X1    g09061(.A1(new_n8799_), .A2(new_n8800_), .ZN(new_n9254_));
  NOR4_X1    g09062(.A1(new_n9212_), .A2(\asqrt[31] ), .A3(new_n9254_), .A4(new_n8804_), .ZN(new_n9255_));
  XOR2_X1    g09063(.A1(new_n9255_), .A2(new_n9253_), .Z(new_n9256_));
  NAND2_X1   g09064(.A1(new_n9256_), .A2(new_n6708_), .ZN(new_n9257_));
  NOR2_X1    g09065(.A1(new_n9252_), .A2(new_n9257_), .ZN(new_n9258_));
  NOR3_X1    g09066(.A1(new_n9258_), .A2(new_n9242_), .A3(new_n9250_), .ZN(new_n9259_));
  INV_X1     g09067(.I(new_n9249_), .ZN(new_n9260_));
  AOI21_X1   g09068(.A1(new_n9251_), .A2(new_n9260_), .B(new_n9242_), .ZN(new_n9261_));
  OAI21_X1   g09069(.A1(new_n9261_), .A2(new_n9252_), .B(\asqrt[32] ), .ZN(new_n9262_));
  NOR4_X1    g09070(.A1(new_n9212_), .A2(\asqrt[32] ), .A3(new_n8807_), .A4(new_n9041_), .ZN(new_n9263_));
  AOI21_X1   g09071(.A1(new_n9253_), .A2(new_n8803_), .B(new_n6708_), .ZN(new_n9264_));
  NOR2_X1    g09072(.A1(new_n9263_), .A2(new_n9264_), .ZN(new_n9265_));
  NAND2_X1   g09073(.A1(new_n9265_), .A2(new_n6365_), .ZN(new_n9266_));
  INV_X1     g09074(.I(new_n9266_), .ZN(new_n9267_));
  NAND2_X1   g09075(.A1(new_n9262_), .A2(new_n9267_), .ZN(new_n9268_));
  NAND2_X1   g09076(.A1(new_n9268_), .A2(new_n9259_), .ZN(new_n9269_));
  OAI21_X1   g09077(.A1(new_n9252_), .A2(new_n9257_), .B(new_n9261_), .ZN(new_n9270_));
  NAND2_X1   g09078(.A1(new_n9270_), .A2(new_n9262_), .ZN(new_n9271_));
  NAND2_X1   g09079(.A1(new_n8819_), .A2(\asqrt[33] ), .ZN(new_n9272_));
  NOR4_X1    g09080(.A1(new_n9212_), .A2(\asqrt[33] ), .A3(new_n8814_), .A4(new_n8819_), .ZN(new_n9273_));
  XOR2_X1    g09081(.A1(new_n9273_), .A2(new_n9272_), .Z(new_n9274_));
  NAND2_X1   g09082(.A1(new_n9274_), .A2(new_n5991_), .ZN(new_n9275_));
  AOI21_X1   g09083(.A1(new_n9271_), .A2(\asqrt[33] ), .B(new_n9275_), .ZN(new_n9276_));
  NOR2_X1    g09084(.A1(new_n9276_), .A2(new_n9269_), .ZN(new_n9277_));
  AOI21_X1   g09085(.A1(new_n9262_), .A2(new_n9267_), .B(new_n9270_), .ZN(new_n9278_));
  AOI21_X1   g09086(.A1(new_n9270_), .A2(new_n9262_), .B(new_n6365_), .ZN(new_n9279_));
  OAI21_X1   g09087(.A1(new_n9278_), .A2(new_n9279_), .B(\asqrt[34] ), .ZN(new_n9280_));
  NOR4_X1    g09088(.A1(new_n9212_), .A2(\asqrt[34] ), .A3(new_n8822_), .A4(new_n9048_), .ZN(new_n9281_));
  AOI21_X1   g09089(.A1(new_n9272_), .A2(new_n8818_), .B(new_n5991_), .ZN(new_n9282_));
  NOR2_X1    g09090(.A1(new_n9281_), .A2(new_n9282_), .ZN(new_n9283_));
  NAND2_X1   g09091(.A1(new_n9283_), .A2(new_n5626_), .ZN(new_n9284_));
  INV_X1     g09092(.I(new_n9284_), .ZN(new_n9285_));
  NAND2_X1   g09093(.A1(new_n9280_), .A2(new_n9285_), .ZN(new_n9286_));
  NAND2_X1   g09094(.A1(new_n9286_), .A2(new_n9277_), .ZN(new_n9287_));
  AOI22_X1   g09095(.A1(new_n9271_), .A2(\asqrt[33] ), .B1(new_n9268_), .B2(new_n9259_), .ZN(new_n9288_));
  OAI22_X1   g09096(.A1(new_n9288_), .A2(new_n5991_), .B1(new_n9276_), .B2(new_n9269_), .ZN(new_n9289_));
  NAND2_X1   g09097(.A1(new_n8833_), .A2(\asqrt[35] ), .ZN(new_n9290_));
  NOR4_X1    g09098(.A1(new_n9212_), .A2(\asqrt[35] ), .A3(new_n8828_), .A4(new_n8833_), .ZN(new_n9291_));
  XOR2_X1    g09099(.A1(new_n9291_), .A2(new_n9290_), .Z(new_n9292_));
  NAND2_X1   g09100(.A1(new_n9292_), .A2(new_n5273_), .ZN(new_n9293_));
  AOI21_X1   g09101(.A1(new_n9289_), .A2(\asqrt[35] ), .B(new_n9293_), .ZN(new_n9294_));
  NOR2_X1    g09102(.A1(new_n9294_), .A2(new_n9287_), .ZN(new_n9295_));
  AOI22_X1   g09103(.A1(new_n9289_), .A2(\asqrt[35] ), .B1(new_n9286_), .B2(new_n9277_), .ZN(new_n9296_));
  NOR4_X1    g09104(.A1(new_n9212_), .A2(\asqrt[36] ), .A3(new_n8835_), .A4(new_n9055_), .ZN(new_n9297_));
  AOI21_X1   g09105(.A1(new_n9290_), .A2(new_n8832_), .B(new_n5273_), .ZN(new_n9298_));
  NOR2_X1    g09106(.A1(new_n9297_), .A2(new_n9298_), .ZN(new_n9299_));
  NAND2_X1   g09107(.A1(new_n9299_), .A2(new_n4973_), .ZN(new_n9300_));
  INV_X1     g09108(.I(new_n9300_), .ZN(new_n9301_));
  OAI21_X1   g09109(.A1(new_n9296_), .A2(new_n5273_), .B(new_n9301_), .ZN(new_n9302_));
  NAND2_X1   g09110(.A1(new_n9302_), .A2(new_n9295_), .ZN(new_n9303_));
  OAI22_X1   g09111(.A1(new_n9296_), .A2(new_n5273_), .B1(new_n9294_), .B2(new_n9287_), .ZN(new_n9304_));
  NAND2_X1   g09112(.A1(new_n8846_), .A2(\asqrt[37] ), .ZN(new_n9305_));
  NOR4_X1    g09113(.A1(new_n9212_), .A2(\asqrt[37] ), .A3(new_n8841_), .A4(new_n8846_), .ZN(new_n9306_));
  XOR2_X1    g09114(.A1(new_n9306_), .A2(new_n9305_), .Z(new_n9307_));
  NAND2_X1   g09115(.A1(new_n9307_), .A2(new_n4645_), .ZN(new_n9308_));
  AOI21_X1   g09116(.A1(new_n9304_), .A2(\asqrt[37] ), .B(new_n9308_), .ZN(new_n9309_));
  NOR2_X1    g09117(.A1(new_n9309_), .A2(new_n9303_), .ZN(new_n9310_));
  AOI22_X1   g09118(.A1(new_n9304_), .A2(\asqrt[37] ), .B1(new_n9302_), .B2(new_n9295_), .ZN(new_n9311_));
  NAND2_X1   g09119(.A1(new_n9062_), .A2(\asqrt[38] ), .ZN(new_n9312_));
  NOR4_X1    g09120(.A1(new_n9212_), .A2(\asqrt[38] ), .A3(new_n8849_), .A4(new_n9062_), .ZN(new_n9313_));
  XOR2_X1    g09121(.A1(new_n9313_), .A2(new_n9312_), .Z(new_n9314_));
  NAND2_X1   g09122(.A1(new_n9314_), .A2(new_n4330_), .ZN(new_n9315_));
  INV_X1     g09123(.I(new_n9315_), .ZN(new_n9316_));
  OAI21_X1   g09124(.A1(new_n9311_), .A2(new_n4645_), .B(new_n9316_), .ZN(new_n9317_));
  NAND2_X1   g09125(.A1(new_n9317_), .A2(new_n9310_), .ZN(new_n9318_));
  OAI22_X1   g09126(.A1(new_n9311_), .A2(new_n4645_), .B1(new_n9309_), .B2(new_n9303_), .ZN(new_n9319_));
  NOR4_X1    g09127(.A1(new_n9212_), .A2(\asqrt[39] ), .A3(new_n8856_), .A4(new_n8861_), .ZN(new_n9320_));
  AOI21_X1   g09128(.A1(new_n9312_), .A2(new_n9061_), .B(new_n4330_), .ZN(new_n9321_));
  NOR2_X1    g09129(.A1(new_n9320_), .A2(new_n9321_), .ZN(new_n9322_));
  NAND2_X1   g09130(.A1(new_n9322_), .A2(new_n4018_), .ZN(new_n9323_));
  AOI21_X1   g09131(.A1(new_n9319_), .A2(\asqrt[39] ), .B(new_n9323_), .ZN(new_n9324_));
  NOR2_X1    g09132(.A1(new_n9324_), .A2(new_n9318_), .ZN(new_n9325_));
  AOI22_X1   g09133(.A1(new_n9319_), .A2(\asqrt[39] ), .B1(new_n9317_), .B2(new_n9310_), .ZN(new_n9326_));
  NAND2_X1   g09134(.A1(new_n9069_), .A2(\asqrt[40] ), .ZN(new_n9327_));
  NOR4_X1    g09135(.A1(new_n9212_), .A2(\asqrt[40] ), .A3(new_n8864_), .A4(new_n9069_), .ZN(new_n9328_));
  XOR2_X1    g09136(.A1(new_n9328_), .A2(new_n9327_), .Z(new_n9329_));
  NAND2_X1   g09137(.A1(new_n9329_), .A2(new_n3760_), .ZN(new_n9330_));
  INV_X1     g09138(.I(new_n9330_), .ZN(new_n9331_));
  OAI21_X1   g09139(.A1(new_n9326_), .A2(new_n4018_), .B(new_n9331_), .ZN(new_n9332_));
  NAND2_X1   g09140(.A1(new_n9332_), .A2(new_n9325_), .ZN(new_n9333_));
  OAI22_X1   g09141(.A1(new_n9326_), .A2(new_n4018_), .B1(new_n9324_), .B2(new_n9318_), .ZN(new_n9334_));
  NOR4_X1    g09142(.A1(new_n9212_), .A2(\asqrt[41] ), .A3(new_n8871_), .A4(new_n8876_), .ZN(new_n9335_));
  AOI21_X1   g09143(.A1(new_n9327_), .A2(new_n9068_), .B(new_n3760_), .ZN(new_n9336_));
  NOR2_X1    g09144(.A1(new_n9335_), .A2(new_n9336_), .ZN(new_n9337_));
  NAND2_X1   g09145(.A1(new_n9337_), .A2(new_n3481_), .ZN(new_n9338_));
  AOI21_X1   g09146(.A1(new_n9334_), .A2(\asqrt[41] ), .B(new_n9338_), .ZN(new_n9339_));
  NOR2_X1    g09147(.A1(new_n9339_), .A2(new_n9333_), .ZN(new_n9340_));
  AOI22_X1   g09148(.A1(new_n9334_), .A2(\asqrt[41] ), .B1(new_n9332_), .B2(new_n9325_), .ZN(new_n9341_));
  NAND2_X1   g09149(.A1(new_n9076_), .A2(\asqrt[42] ), .ZN(new_n9342_));
  NOR4_X1    g09150(.A1(new_n9212_), .A2(\asqrt[42] ), .A3(new_n8879_), .A4(new_n9076_), .ZN(new_n9343_));
  XOR2_X1    g09151(.A1(new_n9343_), .A2(new_n9342_), .Z(new_n9344_));
  NAND2_X1   g09152(.A1(new_n9344_), .A2(new_n3208_), .ZN(new_n9345_));
  INV_X1     g09153(.I(new_n9345_), .ZN(new_n9346_));
  OAI21_X1   g09154(.A1(new_n9341_), .A2(new_n3481_), .B(new_n9346_), .ZN(new_n9347_));
  NAND2_X1   g09155(.A1(new_n9347_), .A2(new_n9340_), .ZN(new_n9348_));
  OAI22_X1   g09156(.A1(new_n9341_), .A2(new_n3481_), .B1(new_n9339_), .B2(new_n9333_), .ZN(new_n9349_));
  NOR4_X1    g09157(.A1(new_n9212_), .A2(\asqrt[43] ), .A3(new_n8886_), .A4(new_n8891_), .ZN(new_n9350_));
  AOI21_X1   g09158(.A1(new_n9342_), .A2(new_n9075_), .B(new_n3208_), .ZN(new_n9351_));
  NOR2_X1    g09159(.A1(new_n9350_), .A2(new_n9351_), .ZN(new_n9352_));
  NAND2_X1   g09160(.A1(new_n9352_), .A2(new_n2941_), .ZN(new_n9353_));
  AOI21_X1   g09161(.A1(new_n9349_), .A2(\asqrt[43] ), .B(new_n9353_), .ZN(new_n9354_));
  NOR2_X1    g09162(.A1(new_n9354_), .A2(new_n9348_), .ZN(new_n9355_));
  AOI22_X1   g09163(.A1(new_n9349_), .A2(\asqrt[43] ), .B1(new_n9347_), .B2(new_n9340_), .ZN(new_n9356_));
  NAND2_X1   g09164(.A1(new_n9083_), .A2(\asqrt[44] ), .ZN(new_n9357_));
  NOR4_X1    g09165(.A1(new_n9212_), .A2(\asqrt[44] ), .A3(new_n8894_), .A4(new_n9083_), .ZN(new_n9358_));
  XOR2_X1    g09166(.A1(new_n9358_), .A2(new_n9357_), .Z(new_n9359_));
  NAND2_X1   g09167(.A1(new_n9359_), .A2(new_n2728_), .ZN(new_n9360_));
  INV_X1     g09168(.I(new_n9360_), .ZN(new_n9361_));
  OAI21_X1   g09169(.A1(new_n9356_), .A2(new_n2941_), .B(new_n9361_), .ZN(new_n9362_));
  NAND2_X1   g09170(.A1(new_n9362_), .A2(new_n9355_), .ZN(new_n9363_));
  OAI22_X1   g09171(.A1(new_n9356_), .A2(new_n2941_), .B1(new_n9354_), .B2(new_n9348_), .ZN(new_n9364_));
  NOR4_X1    g09172(.A1(new_n9212_), .A2(\asqrt[45] ), .A3(new_n8901_), .A4(new_n8906_), .ZN(new_n9365_));
  AOI21_X1   g09173(.A1(new_n9357_), .A2(new_n9082_), .B(new_n2728_), .ZN(new_n9366_));
  NOR2_X1    g09174(.A1(new_n9365_), .A2(new_n9366_), .ZN(new_n9367_));
  NAND2_X1   g09175(.A1(new_n9367_), .A2(new_n2488_), .ZN(new_n9368_));
  AOI21_X1   g09176(.A1(new_n9364_), .A2(\asqrt[45] ), .B(new_n9368_), .ZN(new_n9369_));
  NOR2_X1    g09177(.A1(new_n9369_), .A2(new_n9363_), .ZN(new_n9370_));
  AOI22_X1   g09178(.A1(new_n9364_), .A2(\asqrt[45] ), .B1(new_n9362_), .B2(new_n9355_), .ZN(new_n9371_));
  NAND2_X1   g09179(.A1(new_n9090_), .A2(\asqrt[46] ), .ZN(new_n9372_));
  NOR4_X1    g09180(.A1(new_n9212_), .A2(\asqrt[46] ), .A3(new_n8909_), .A4(new_n9090_), .ZN(new_n9373_));
  XOR2_X1    g09181(.A1(new_n9373_), .A2(new_n9372_), .Z(new_n9374_));
  NAND2_X1   g09182(.A1(new_n9374_), .A2(new_n2253_), .ZN(new_n9375_));
  INV_X1     g09183(.I(new_n9375_), .ZN(new_n9376_));
  OAI21_X1   g09184(.A1(new_n9371_), .A2(new_n2488_), .B(new_n9376_), .ZN(new_n9377_));
  NAND2_X1   g09185(.A1(new_n9377_), .A2(new_n9370_), .ZN(new_n9378_));
  OAI22_X1   g09186(.A1(new_n9371_), .A2(new_n2488_), .B1(new_n9369_), .B2(new_n9363_), .ZN(new_n9379_));
  NAND2_X1   g09187(.A1(new_n8921_), .A2(\asqrt[47] ), .ZN(new_n9380_));
  NOR4_X1    g09188(.A1(new_n9212_), .A2(\asqrt[47] ), .A3(new_n8916_), .A4(new_n8921_), .ZN(new_n9381_));
  XOR2_X1    g09189(.A1(new_n9381_), .A2(new_n9380_), .Z(new_n9382_));
  NAND2_X1   g09190(.A1(new_n9382_), .A2(new_n2046_), .ZN(new_n9383_));
  AOI21_X1   g09191(.A1(new_n9379_), .A2(\asqrt[47] ), .B(new_n9383_), .ZN(new_n9384_));
  NOR2_X1    g09192(.A1(new_n9384_), .A2(new_n9378_), .ZN(new_n9385_));
  AOI22_X1   g09193(.A1(new_n9379_), .A2(\asqrt[47] ), .B1(new_n9377_), .B2(new_n9370_), .ZN(new_n9386_));
  NOR4_X1    g09194(.A1(new_n9212_), .A2(\asqrt[48] ), .A3(new_n8924_), .A4(new_n9097_), .ZN(new_n9387_));
  AOI21_X1   g09195(.A1(new_n9380_), .A2(new_n8920_), .B(new_n2046_), .ZN(new_n9388_));
  NOR2_X1    g09196(.A1(new_n9387_), .A2(new_n9388_), .ZN(new_n9389_));
  NAND2_X1   g09197(.A1(new_n9389_), .A2(new_n1854_), .ZN(new_n9390_));
  INV_X1     g09198(.I(new_n9390_), .ZN(new_n9391_));
  OAI21_X1   g09199(.A1(new_n9386_), .A2(new_n2046_), .B(new_n9391_), .ZN(new_n9392_));
  NAND2_X1   g09200(.A1(new_n9392_), .A2(new_n9385_), .ZN(new_n9393_));
  OAI22_X1   g09201(.A1(new_n9386_), .A2(new_n2046_), .B1(new_n9384_), .B2(new_n9378_), .ZN(new_n9394_));
  NAND2_X1   g09202(.A1(new_n8936_), .A2(\asqrt[49] ), .ZN(new_n9395_));
  NOR4_X1    g09203(.A1(new_n9212_), .A2(\asqrt[49] ), .A3(new_n8931_), .A4(new_n8936_), .ZN(new_n9396_));
  XOR2_X1    g09204(.A1(new_n9396_), .A2(new_n9395_), .Z(new_n9397_));
  NAND2_X1   g09205(.A1(new_n9397_), .A2(new_n1595_), .ZN(new_n9398_));
  AOI21_X1   g09206(.A1(new_n9394_), .A2(\asqrt[49] ), .B(new_n9398_), .ZN(new_n9399_));
  NOR2_X1    g09207(.A1(new_n9399_), .A2(new_n9393_), .ZN(new_n9400_));
  AOI22_X1   g09208(.A1(new_n9394_), .A2(\asqrt[49] ), .B1(new_n9392_), .B2(new_n9385_), .ZN(new_n9401_));
  NOR4_X1    g09209(.A1(new_n9212_), .A2(\asqrt[50] ), .A3(new_n8939_), .A4(new_n9104_), .ZN(new_n9402_));
  AOI21_X1   g09210(.A1(new_n9395_), .A2(new_n8935_), .B(new_n1595_), .ZN(new_n9403_));
  NOR2_X1    g09211(.A1(new_n9402_), .A2(new_n9403_), .ZN(new_n9404_));
  NAND2_X1   g09212(.A1(new_n9404_), .A2(new_n1436_), .ZN(new_n9405_));
  INV_X1     g09213(.I(new_n9405_), .ZN(new_n9406_));
  OAI21_X1   g09214(.A1(new_n9401_), .A2(new_n1595_), .B(new_n9406_), .ZN(new_n9407_));
  NAND2_X1   g09215(.A1(new_n9407_), .A2(new_n9400_), .ZN(new_n9408_));
  OAI22_X1   g09216(.A1(new_n9401_), .A2(new_n1595_), .B1(new_n9399_), .B2(new_n9393_), .ZN(new_n9409_));
  NAND2_X1   g09217(.A1(new_n8951_), .A2(\asqrt[51] ), .ZN(new_n9410_));
  NOR4_X1    g09218(.A1(new_n9212_), .A2(\asqrt[51] ), .A3(new_n8946_), .A4(new_n8951_), .ZN(new_n9411_));
  XOR2_X1    g09219(.A1(new_n9411_), .A2(new_n9410_), .Z(new_n9412_));
  NAND2_X1   g09220(.A1(new_n9412_), .A2(new_n1260_), .ZN(new_n9413_));
  AOI21_X1   g09221(.A1(new_n9409_), .A2(\asqrt[51] ), .B(new_n9413_), .ZN(new_n9414_));
  NOR2_X1    g09222(.A1(new_n9414_), .A2(new_n9408_), .ZN(new_n9415_));
  AOI22_X1   g09223(.A1(new_n9409_), .A2(\asqrt[51] ), .B1(new_n9407_), .B2(new_n9400_), .ZN(new_n9416_));
  NAND2_X1   g09224(.A1(new_n9111_), .A2(\asqrt[52] ), .ZN(new_n9417_));
  NOR4_X1    g09225(.A1(new_n9212_), .A2(\asqrt[52] ), .A3(new_n8954_), .A4(new_n9111_), .ZN(new_n9418_));
  XOR2_X1    g09226(.A1(new_n9418_), .A2(new_n9417_), .Z(new_n9419_));
  NAND2_X1   g09227(.A1(new_n9419_), .A2(new_n1096_), .ZN(new_n9420_));
  INV_X1     g09228(.I(new_n9420_), .ZN(new_n9421_));
  OAI21_X1   g09229(.A1(new_n9416_), .A2(new_n1260_), .B(new_n9421_), .ZN(new_n9422_));
  NAND2_X1   g09230(.A1(new_n9422_), .A2(new_n9415_), .ZN(new_n9423_));
  OAI22_X1   g09231(.A1(new_n9416_), .A2(new_n1260_), .B1(new_n9414_), .B2(new_n9408_), .ZN(new_n9424_));
  NOR4_X1    g09232(.A1(new_n9212_), .A2(\asqrt[53] ), .A3(new_n8960_), .A4(new_n8965_), .ZN(new_n9425_));
  AOI21_X1   g09233(.A1(new_n9417_), .A2(new_n9110_), .B(new_n1096_), .ZN(new_n9426_));
  NOR2_X1    g09234(.A1(new_n9425_), .A2(new_n9426_), .ZN(new_n9427_));
  NAND2_X1   g09235(.A1(new_n9427_), .A2(new_n970_), .ZN(new_n9428_));
  AOI21_X1   g09236(.A1(new_n9424_), .A2(\asqrt[53] ), .B(new_n9428_), .ZN(new_n9429_));
  NOR2_X1    g09237(.A1(new_n9429_), .A2(new_n9423_), .ZN(new_n9430_));
  AOI22_X1   g09238(.A1(new_n9424_), .A2(\asqrt[53] ), .B1(new_n9422_), .B2(new_n9415_), .ZN(new_n9431_));
  NAND2_X1   g09239(.A1(new_n9118_), .A2(\asqrt[54] ), .ZN(new_n9432_));
  NOR4_X1    g09240(.A1(new_n9212_), .A2(\asqrt[54] ), .A3(new_n8967_), .A4(new_n9118_), .ZN(new_n9433_));
  XOR2_X1    g09241(.A1(new_n9433_), .A2(new_n9432_), .Z(new_n9434_));
  NAND2_X1   g09242(.A1(new_n9434_), .A2(new_n825_), .ZN(new_n9435_));
  INV_X1     g09243(.I(new_n9435_), .ZN(new_n9436_));
  OAI21_X1   g09244(.A1(new_n9431_), .A2(new_n970_), .B(new_n9436_), .ZN(new_n9437_));
  NAND2_X1   g09245(.A1(new_n9437_), .A2(new_n9430_), .ZN(new_n9438_));
  OAI22_X1   g09246(.A1(new_n9431_), .A2(new_n970_), .B1(new_n9429_), .B2(new_n9423_), .ZN(new_n9439_));
  NOR4_X1    g09247(.A1(new_n9212_), .A2(\asqrt[55] ), .A3(new_n8973_), .A4(new_n8978_), .ZN(new_n9440_));
  AOI21_X1   g09248(.A1(new_n9432_), .A2(new_n9117_), .B(new_n825_), .ZN(new_n9441_));
  NOR2_X1    g09249(.A1(new_n9440_), .A2(new_n9441_), .ZN(new_n9442_));
  NAND2_X1   g09250(.A1(new_n9442_), .A2(new_n724_), .ZN(new_n9443_));
  AOI21_X1   g09251(.A1(new_n9439_), .A2(\asqrt[55] ), .B(new_n9443_), .ZN(new_n9444_));
  NOR2_X1    g09252(.A1(new_n9444_), .A2(new_n9438_), .ZN(new_n9445_));
  AOI22_X1   g09253(.A1(new_n9439_), .A2(\asqrt[55] ), .B1(new_n9437_), .B2(new_n9430_), .ZN(new_n9446_));
  NAND2_X1   g09254(.A1(new_n9125_), .A2(\asqrt[56] ), .ZN(new_n9447_));
  NOR4_X1    g09255(.A1(new_n9212_), .A2(\asqrt[56] ), .A3(new_n8980_), .A4(new_n9125_), .ZN(new_n9448_));
  XOR2_X1    g09256(.A1(new_n9448_), .A2(new_n9447_), .Z(new_n9449_));
  NAND2_X1   g09257(.A1(new_n9449_), .A2(new_n587_), .ZN(new_n9450_));
  INV_X1     g09258(.I(new_n9450_), .ZN(new_n9451_));
  OAI21_X1   g09259(.A1(new_n9446_), .A2(new_n724_), .B(new_n9451_), .ZN(new_n9452_));
  NAND2_X1   g09260(.A1(new_n9452_), .A2(new_n9445_), .ZN(new_n9453_));
  NAND2_X1   g09261(.A1(new_n9439_), .A2(\asqrt[55] ), .ZN(new_n9454_));
  AOI21_X1   g09262(.A1(new_n9454_), .A2(new_n9438_), .B(new_n724_), .ZN(new_n9455_));
  OAI21_X1   g09263(.A1(new_n9445_), .A2(new_n9455_), .B(\asqrt[57] ), .ZN(new_n9456_));
  NOR2_X1    g09264(.A1(new_n9128_), .A2(new_n587_), .ZN(new_n9457_));
  NOR4_X1    g09265(.A1(new_n9212_), .A2(\asqrt[57] ), .A3(new_n8986_), .A4(new_n8991_), .ZN(new_n9458_));
  XNOR2_X1   g09266(.A1(new_n9458_), .A2(new_n9457_), .ZN(new_n9459_));
  NAND2_X1   g09267(.A1(new_n9459_), .A2(new_n504_), .ZN(new_n9460_));
  INV_X1     g09268(.I(new_n9460_), .ZN(new_n9461_));
  AOI21_X1   g09269(.A1(new_n9456_), .A2(new_n9461_), .B(new_n9453_), .ZN(new_n9462_));
  OAI22_X1   g09270(.A1(new_n9446_), .A2(new_n724_), .B1(new_n9444_), .B2(new_n9438_), .ZN(new_n9463_));
  AOI22_X1   g09271(.A1(new_n9463_), .A2(\asqrt[57] ), .B1(new_n9452_), .B2(new_n9445_), .ZN(new_n9464_));
  NOR4_X1    g09272(.A1(new_n9212_), .A2(\asqrt[58] ), .A3(new_n8993_), .A4(new_n9132_), .ZN(new_n9465_));
  XOR2_X1    g09273(.A1(new_n9465_), .A2(new_n9176_), .Z(new_n9466_));
  NAND2_X1   g09274(.A1(new_n9466_), .A2(new_n376_), .ZN(new_n9467_));
  INV_X1     g09275(.I(new_n9467_), .ZN(new_n9468_));
  OAI21_X1   g09276(.A1(new_n9464_), .A2(new_n504_), .B(new_n9468_), .ZN(new_n9469_));
  NAND2_X1   g09277(.A1(new_n9469_), .A2(new_n9462_), .ZN(new_n9470_));
  AOI21_X1   g09278(.A1(new_n9453_), .A2(new_n9456_), .B(new_n504_), .ZN(new_n9471_));
  OAI21_X1   g09279(.A1(new_n9462_), .A2(new_n9471_), .B(\asqrt[59] ), .ZN(new_n9472_));
  NOR4_X1    g09280(.A1(new_n9212_), .A2(\asqrt[59] ), .A3(new_n8999_), .A4(new_n9004_), .ZN(new_n9473_));
  XOR2_X1    g09281(.A1(new_n9473_), .A2(new_n9154_), .Z(new_n9474_));
  AND2_X2    g09282(.A1(new_n9474_), .A2(new_n275_), .Z(new_n9475_));
  AOI21_X1   g09283(.A1(new_n9472_), .A2(new_n9475_), .B(new_n9470_), .ZN(new_n9476_));
  INV_X1     g09284(.I(new_n9241_), .ZN(new_n9477_));
  OAI21_X1   g09285(.A1(new_n9243_), .A2(new_n7931_), .B(new_n9477_), .ZN(new_n9478_));
  AOI22_X1   g09286(.A1(new_n9244_), .A2(\asqrt[30] ), .B1(new_n9478_), .B2(new_n9234_), .ZN(new_n9479_));
  INV_X1     g09287(.I(new_n9257_), .ZN(new_n9480_));
  OAI21_X1   g09288(.A1(new_n9479_), .A2(new_n7110_), .B(new_n9480_), .ZN(new_n9481_));
  OAI22_X1   g09289(.A1(new_n9479_), .A2(new_n7110_), .B1(new_n9250_), .B2(new_n9242_), .ZN(new_n9482_));
  AOI22_X1   g09290(.A1(new_n9482_), .A2(\asqrt[32] ), .B1(new_n9481_), .B2(new_n9261_), .ZN(new_n9483_));
  INV_X1     g09291(.I(new_n9275_), .ZN(new_n9484_));
  OAI21_X1   g09292(.A1(new_n9483_), .A2(new_n6365_), .B(new_n9484_), .ZN(new_n9485_));
  NAND2_X1   g09293(.A1(new_n9485_), .A2(new_n9278_), .ZN(new_n9486_));
  AOI21_X1   g09294(.A1(new_n9482_), .A2(\asqrt[32] ), .B(new_n9266_), .ZN(new_n9487_));
  OAI22_X1   g09295(.A1(new_n9483_), .A2(new_n6365_), .B1(new_n9487_), .B2(new_n9270_), .ZN(new_n9488_));
  AOI21_X1   g09296(.A1(new_n9488_), .A2(\asqrt[34] ), .B(new_n9284_), .ZN(new_n9489_));
  NOR2_X1    g09297(.A1(new_n9489_), .A2(new_n9486_), .ZN(new_n9490_));
  AOI22_X1   g09298(.A1(new_n9488_), .A2(\asqrt[34] ), .B1(new_n9485_), .B2(new_n9278_), .ZN(new_n9491_));
  INV_X1     g09299(.I(new_n9293_), .ZN(new_n9492_));
  OAI21_X1   g09300(.A1(new_n9491_), .A2(new_n5626_), .B(new_n9492_), .ZN(new_n9493_));
  NAND2_X1   g09301(.A1(new_n9493_), .A2(new_n9490_), .ZN(new_n9494_));
  OAI22_X1   g09302(.A1(new_n9491_), .A2(new_n5626_), .B1(new_n9489_), .B2(new_n9486_), .ZN(new_n9495_));
  AOI21_X1   g09303(.A1(new_n9495_), .A2(\asqrt[36] ), .B(new_n9300_), .ZN(new_n9496_));
  NOR2_X1    g09304(.A1(new_n9496_), .A2(new_n9494_), .ZN(new_n9497_));
  AOI22_X1   g09305(.A1(new_n9495_), .A2(\asqrt[36] ), .B1(new_n9493_), .B2(new_n9490_), .ZN(new_n9498_));
  INV_X1     g09306(.I(new_n9308_), .ZN(new_n9499_));
  OAI21_X1   g09307(.A1(new_n9498_), .A2(new_n4973_), .B(new_n9499_), .ZN(new_n9500_));
  NAND2_X1   g09308(.A1(new_n9500_), .A2(new_n9497_), .ZN(new_n9501_));
  OAI22_X1   g09309(.A1(new_n9498_), .A2(new_n4973_), .B1(new_n9496_), .B2(new_n9494_), .ZN(new_n9502_));
  AOI21_X1   g09310(.A1(new_n9502_), .A2(\asqrt[38] ), .B(new_n9315_), .ZN(new_n9503_));
  NOR2_X1    g09311(.A1(new_n9503_), .A2(new_n9501_), .ZN(new_n9504_));
  AOI22_X1   g09312(.A1(new_n9502_), .A2(\asqrt[38] ), .B1(new_n9500_), .B2(new_n9497_), .ZN(new_n9505_));
  INV_X1     g09313(.I(new_n9323_), .ZN(new_n9506_));
  OAI21_X1   g09314(.A1(new_n9505_), .A2(new_n4330_), .B(new_n9506_), .ZN(new_n9507_));
  NAND2_X1   g09315(.A1(new_n9507_), .A2(new_n9504_), .ZN(new_n9508_));
  OAI22_X1   g09316(.A1(new_n9505_), .A2(new_n4330_), .B1(new_n9503_), .B2(new_n9501_), .ZN(new_n9509_));
  AOI21_X1   g09317(.A1(new_n9509_), .A2(\asqrt[40] ), .B(new_n9330_), .ZN(new_n9510_));
  NOR2_X1    g09318(.A1(new_n9510_), .A2(new_n9508_), .ZN(new_n9511_));
  AOI22_X1   g09319(.A1(new_n9509_), .A2(\asqrt[40] ), .B1(new_n9507_), .B2(new_n9504_), .ZN(new_n9512_));
  INV_X1     g09320(.I(new_n9338_), .ZN(new_n9513_));
  OAI21_X1   g09321(.A1(new_n9512_), .A2(new_n3760_), .B(new_n9513_), .ZN(new_n9514_));
  NAND2_X1   g09322(.A1(new_n9514_), .A2(new_n9511_), .ZN(new_n9515_));
  OAI22_X1   g09323(.A1(new_n9512_), .A2(new_n3760_), .B1(new_n9510_), .B2(new_n9508_), .ZN(new_n9516_));
  AOI21_X1   g09324(.A1(new_n9516_), .A2(\asqrt[42] ), .B(new_n9345_), .ZN(new_n9517_));
  NOR2_X1    g09325(.A1(new_n9517_), .A2(new_n9515_), .ZN(new_n9518_));
  AOI22_X1   g09326(.A1(new_n9516_), .A2(\asqrt[42] ), .B1(new_n9514_), .B2(new_n9511_), .ZN(new_n9519_));
  INV_X1     g09327(.I(new_n9353_), .ZN(new_n9520_));
  OAI21_X1   g09328(.A1(new_n9519_), .A2(new_n3208_), .B(new_n9520_), .ZN(new_n9521_));
  NAND2_X1   g09329(.A1(new_n9521_), .A2(new_n9518_), .ZN(new_n9522_));
  OAI22_X1   g09330(.A1(new_n9519_), .A2(new_n3208_), .B1(new_n9517_), .B2(new_n9515_), .ZN(new_n9523_));
  AOI21_X1   g09331(.A1(new_n9523_), .A2(\asqrt[44] ), .B(new_n9360_), .ZN(new_n9524_));
  NOR2_X1    g09332(.A1(new_n9524_), .A2(new_n9522_), .ZN(new_n9525_));
  AOI22_X1   g09333(.A1(new_n9523_), .A2(\asqrt[44] ), .B1(new_n9521_), .B2(new_n9518_), .ZN(new_n9526_));
  INV_X1     g09334(.I(new_n9368_), .ZN(new_n9527_));
  OAI21_X1   g09335(.A1(new_n9526_), .A2(new_n2728_), .B(new_n9527_), .ZN(new_n9528_));
  NAND2_X1   g09336(.A1(new_n9528_), .A2(new_n9525_), .ZN(new_n9529_));
  OAI22_X1   g09337(.A1(new_n9526_), .A2(new_n2728_), .B1(new_n9524_), .B2(new_n9522_), .ZN(new_n9530_));
  AOI21_X1   g09338(.A1(new_n9530_), .A2(\asqrt[46] ), .B(new_n9375_), .ZN(new_n9531_));
  NOR2_X1    g09339(.A1(new_n9531_), .A2(new_n9529_), .ZN(new_n9532_));
  AOI22_X1   g09340(.A1(new_n9530_), .A2(\asqrt[46] ), .B1(new_n9528_), .B2(new_n9525_), .ZN(new_n9533_));
  INV_X1     g09341(.I(new_n9383_), .ZN(new_n9534_));
  OAI21_X1   g09342(.A1(new_n9533_), .A2(new_n2253_), .B(new_n9534_), .ZN(new_n9535_));
  NAND2_X1   g09343(.A1(new_n9535_), .A2(new_n9532_), .ZN(new_n9536_));
  OAI22_X1   g09344(.A1(new_n9533_), .A2(new_n2253_), .B1(new_n9531_), .B2(new_n9529_), .ZN(new_n9537_));
  AOI21_X1   g09345(.A1(new_n9537_), .A2(\asqrt[48] ), .B(new_n9390_), .ZN(new_n9538_));
  NOR2_X1    g09346(.A1(new_n9538_), .A2(new_n9536_), .ZN(new_n9539_));
  AOI22_X1   g09347(.A1(new_n9537_), .A2(\asqrt[48] ), .B1(new_n9535_), .B2(new_n9532_), .ZN(new_n9540_));
  INV_X1     g09348(.I(new_n9398_), .ZN(new_n9541_));
  OAI21_X1   g09349(.A1(new_n9540_), .A2(new_n1854_), .B(new_n9541_), .ZN(new_n9542_));
  NAND2_X1   g09350(.A1(new_n9542_), .A2(new_n9539_), .ZN(new_n9543_));
  OAI22_X1   g09351(.A1(new_n9540_), .A2(new_n1854_), .B1(new_n9538_), .B2(new_n9536_), .ZN(new_n9544_));
  AOI21_X1   g09352(.A1(new_n9544_), .A2(\asqrt[50] ), .B(new_n9405_), .ZN(new_n9545_));
  NOR2_X1    g09353(.A1(new_n9545_), .A2(new_n9543_), .ZN(new_n9546_));
  AOI22_X1   g09354(.A1(new_n9544_), .A2(\asqrt[50] ), .B1(new_n9542_), .B2(new_n9539_), .ZN(new_n9547_));
  INV_X1     g09355(.I(new_n9413_), .ZN(new_n9548_));
  OAI21_X1   g09356(.A1(new_n9547_), .A2(new_n1436_), .B(new_n9548_), .ZN(new_n9549_));
  NAND2_X1   g09357(.A1(new_n9549_), .A2(new_n9546_), .ZN(new_n9550_));
  OAI22_X1   g09358(.A1(new_n9547_), .A2(new_n1436_), .B1(new_n9545_), .B2(new_n9543_), .ZN(new_n9551_));
  AOI21_X1   g09359(.A1(new_n9551_), .A2(\asqrt[52] ), .B(new_n9420_), .ZN(new_n9552_));
  NOR2_X1    g09360(.A1(new_n9552_), .A2(new_n9550_), .ZN(new_n9553_));
  AOI22_X1   g09361(.A1(new_n9551_), .A2(\asqrt[52] ), .B1(new_n9549_), .B2(new_n9546_), .ZN(new_n9554_));
  INV_X1     g09362(.I(new_n9428_), .ZN(new_n9555_));
  OAI21_X1   g09363(.A1(new_n9554_), .A2(new_n1096_), .B(new_n9555_), .ZN(new_n9556_));
  NAND2_X1   g09364(.A1(new_n9556_), .A2(new_n9553_), .ZN(new_n9557_));
  OAI22_X1   g09365(.A1(new_n9554_), .A2(new_n1096_), .B1(new_n9552_), .B2(new_n9550_), .ZN(new_n9558_));
  AOI21_X1   g09366(.A1(new_n9558_), .A2(\asqrt[54] ), .B(new_n9435_), .ZN(new_n9559_));
  NOR2_X1    g09367(.A1(new_n9559_), .A2(new_n9557_), .ZN(new_n9560_));
  AOI22_X1   g09368(.A1(new_n9558_), .A2(\asqrt[54] ), .B1(new_n9556_), .B2(new_n9553_), .ZN(new_n9561_));
  INV_X1     g09369(.I(new_n9443_), .ZN(new_n9562_));
  OAI21_X1   g09370(.A1(new_n9561_), .A2(new_n825_), .B(new_n9562_), .ZN(new_n9563_));
  NAND2_X1   g09371(.A1(new_n9563_), .A2(new_n9560_), .ZN(new_n9564_));
  OAI22_X1   g09372(.A1(new_n9561_), .A2(new_n825_), .B1(new_n9559_), .B2(new_n9557_), .ZN(new_n9565_));
  AOI21_X1   g09373(.A1(new_n9565_), .A2(\asqrt[56] ), .B(new_n9450_), .ZN(new_n9566_));
  NOR2_X1    g09374(.A1(new_n9566_), .A2(new_n9564_), .ZN(new_n9567_));
  AOI22_X1   g09375(.A1(new_n9565_), .A2(\asqrt[56] ), .B1(new_n9563_), .B2(new_n9560_), .ZN(new_n9568_));
  OAI21_X1   g09376(.A1(new_n9568_), .A2(new_n587_), .B(new_n9461_), .ZN(new_n9569_));
  NAND2_X1   g09377(.A1(new_n9569_), .A2(new_n9567_), .ZN(new_n9570_));
  NAND2_X1   g09378(.A1(new_n9558_), .A2(\asqrt[54] ), .ZN(new_n9571_));
  AOI21_X1   g09379(.A1(new_n9571_), .A2(new_n9557_), .B(new_n825_), .ZN(new_n9572_));
  OAI21_X1   g09380(.A1(new_n9560_), .A2(new_n9572_), .B(\asqrt[56] ), .ZN(new_n9573_));
  AOI21_X1   g09381(.A1(new_n9564_), .A2(new_n9573_), .B(new_n587_), .ZN(new_n9574_));
  OAI21_X1   g09382(.A1(new_n9567_), .A2(new_n9574_), .B(\asqrt[58] ), .ZN(new_n9575_));
  NAND2_X1   g09383(.A1(new_n9570_), .A2(new_n9575_), .ZN(new_n9576_));
  AOI22_X1   g09384(.A1(new_n9576_), .A2(\asqrt[59] ), .B1(new_n9469_), .B2(new_n9462_), .ZN(new_n9577_));
  NOR4_X1    g09385(.A1(new_n9212_), .A2(\asqrt[60] ), .A3(new_n9006_), .A4(new_n9139_), .ZN(new_n9578_));
  XOR2_X1    g09386(.A1(new_n9578_), .A2(new_n9178_), .Z(new_n9579_));
  NAND2_X1   g09387(.A1(new_n9579_), .A2(new_n229_), .ZN(new_n9580_));
  INV_X1     g09388(.I(new_n9580_), .ZN(new_n9581_));
  OAI21_X1   g09389(.A1(new_n9577_), .A2(new_n275_), .B(new_n9581_), .ZN(new_n9582_));
  OAI22_X1   g09390(.A1(new_n9568_), .A2(new_n587_), .B1(new_n9566_), .B2(new_n9564_), .ZN(new_n9583_));
  AOI21_X1   g09391(.A1(new_n9583_), .A2(\asqrt[58] ), .B(new_n9467_), .ZN(new_n9584_));
  NOR2_X1    g09392(.A1(new_n9584_), .A2(new_n9570_), .ZN(new_n9585_));
  AOI22_X1   g09393(.A1(new_n9583_), .A2(\asqrt[58] ), .B1(new_n9569_), .B2(new_n9567_), .ZN(new_n9586_));
  OAI21_X1   g09394(.A1(new_n9586_), .A2(new_n376_), .B(new_n9475_), .ZN(new_n9587_));
  NAND2_X1   g09395(.A1(new_n9587_), .A2(new_n9585_), .ZN(new_n9588_));
  AOI21_X1   g09396(.A1(new_n9570_), .A2(new_n9575_), .B(new_n376_), .ZN(new_n9589_));
  OAI21_X1   g09397(.A1(new_n9585_), .A2(new_n9589_), .B(\asqrt[60] ), .ZN(new_n9590_));
  AOI21_X1   g09398(.A1(new_n9588_), .A2(new_n9590_), .B(new_n229_), .ZN(new_n9591_));
  INV_X1     g09399(.I(new_n9182_), .ZN(new_n9592_));
  NOR2_X1    g09400(.A1(new_n9592_), .A2(\asqrt[62] ), .ZN(new_n9593_));
  INV_X1     g09401(.I(new_n9593_), .ZN(new_n9594_));
  NAND4_X1   g09402(.A1(new_n9591_), .A2(new_n9476_), .A3(new_n9582_), .A4(new_n9594_), .ZN(new_n9595_));
  NAND2_X1   g09403(.A1(new_n9200_), .A2(new_n9150_), .ZN(new_n9596_));
  OAI21_X1   g09404(.A1(\asqrt[26] ), .A2(new_n9596_), .B(new_n9160_), .ZN(new_n9597_));
  NAND2_X1   g09405(.A1(new_n9597_), .A2(new_n231_), .ZN(new_n9598_));
  INV_X1     g09406(.I(new_n9598_), .ZN(new_n9599_));
  NAND3_X1   g09407(.A1(new_n9595_), .A2(new_n9184_), .A3(new_n9599_), .ZN(new_n9600_));
  OAI22_X1   g09408(.A1(new_n9586_), .A2(new_n376_), .B1(new_n9584_), .B2(new_n9570_), .ZN(new_n9601_));
  AOI21_X1   g09409(.A1(new_n9601_), .A2(\asqrt[60] ), .B(new_n9580_), .ZN(new_n9602_));
  AOI22_X1   g09410(.A1(new_n9601_), .A2(\asqrt[60] ), .B1(new_n9587_), .B2(new_n9585_), .ZN(new_n9603_));
  OAI22_X1   g09411(.A1(new_n9603_), .A2(new_n229_), .B1(new_n9602_), .B2(new_n9588_), .ZN(new_n9604_));
  NOR4_X1    g09412(.A1(new_n9604_), .A2(\asqrt[62] ), .A3(new_n9174_), .A4(new_n9182_), .ZN(new_n9605_));
  AOI21_X1   g09413(.A1(new_n9175_), .A2(new_n9600_), .B(new_n9605_), .ZN(new_n9606_));
  INV_X1     g09414(.I(\a[48] ), .ZN(new_n9607_));
  OAI21_X1   g09415(.A1(new_n9151_), .A2(new_n9160_), .B(\asqrt[26] ), .ZN(new_n9608_));
  XOR2_X1    g09416(.A1(new_n9160_), .A2(\asqrt[63] ), .Z(new_n9609_));
  NAND2_X1   g09417(.A1(new_n9608_), .A2(new_n9609_), .ZN(new_n9610_));
  INV_X1     g09418(.I(new_n9610_), .ZN(new_n9611_));
  NAND3_X1   g09419(.A1(new_n9206_), .A2(new_n9144_), .A3(new_n9151_), .ZN(new_n9612_));
  INV_X1     g09420(.I(new_n9612_), .ZN(new_n9613_));
  NOR2_X1    g09421(.A1(new_n9611_), .A2(new_n9613_), .ZN(new_n9614_));
  NOR2_X1    g09422(.A1(\a[46] ), .A2(\a[47] ), .ZN(new_n9615_));
  INV_X1     g09423(.I(new_n9615_), .ZN(new_n9616_));
  NOR3_X1    g09424(.A1(new_n9614_), .A2(new_n9607_), .A3(new_n9616_), .ZN(new_n9617_));
  NAND2_X1   g09425(.A1(new_n9606_), .A2(new_n9617_), .ZN(new_n9618_));
  XOR2_X1    g09426(.A1(new_n9618_), .A2(\a[49] ), .Z(new_n9619_));
  INV_X1     g09427(.I(\a[49] ), .ZN(new_n9620_));
  NAND2_X1   g09428(.A1(new_n9582_), .A2(new_n9476_), .ZN(new_n9621_));
  NAND2_X1   g09429(.A1(new_n9591_), .A2(new_n9594_), .ZN(new_n9622_));
  OAI21_X1   g09430(.A1(new_n9622_), .A2(new_n9621_), .B(new_n9184_), .ZN(new_n9623_));
  OAI21_X1   g09431(.A1(new_n9623_), .A2(new_n9598_), .B(new_n9175_), .ZN(new_n9624_));
  NAND2_X1   g09432(.A1(new_n9605_), .A2(new_n9611_), .ZN(new_n9625_));
  NOR2_X1    g09433(.A1(new_n9625_), .A2(new_n9624_), .ZN(new_n9626_));
  NAND3_X1   g09434(.A1(new_n9626_), .A2(new_n9175_), .A3(new_n9612_), .ZN(new_n9627_));
  NAND2_X1   g09435(.A1(new_n9588_), .A2(new_n9590_), .ZN(new_n9628_));
  AOI22_X1   g09436(.A1(new_n9628_), .A2(\asqrt[61] ), .B1(new_n9582_), .B2(new_n9476_), .ZN(new_n9629_));
  NOR2_X1    g09437(.A1(new_n9629_), .A2(new_n196_), .ZN(new_n9630_));
  AOI21_X1   g09438(.A1(new_n9470_), .A2(new_n9472_), .B(new_n275_), .ZN(new_n9631_));
  OAI21_X1   g09439(.A1(new_n9476_), .A2(new_n9631_), .B(\asqrt[61] ), .ZN(new_n9632_));
  NAND4_X1   g09440(.A1(new_n9621_), .A2(new_n196_), .A3(new_n9632_), .A4(new_n9592_), .ZN(new_n9633_));
  INV_X1     g09441(.I(new_n9633_), .ZN(new_n9634_));
  NOR3_X1    g09442(.A1(new_n9625_), .A2(new_n9624_), .A3(new_n9612_), .ZN(\asqrt[25] ));
  NAND3_X1   g09443(.A1(\asqrt[25] ), .A2(new_n9630_), .A3(new_n9634_), .ZN(new_n9636_));
  OAI21_X1   g09444(.A1(new_n9604_), .A2(\asqrt[62] ), .B(new_n9182_), .ZN(new_n9637_));
  OAI21_X1   g09445(.A1(\asqrt[25] ), .A2(new_n9637_), .B(new_n9630_), .ZN(new_n9638_));
  NAND2_X1   g09446(.A1(new_n9638_), .A2(new_n9636_), .ZN(new_n9639_));
  INV_X1     g09447(.I(new_n9639_), .ZN(new_n9640_));
  NOR3_X1    g09448(.A1(new_n9628_), .A2(\asqrt[61] ), .A3(new_n9579_), .ZN(new_n9641_));
  NAND2_X1   g09449(.A1(\asqrt[25] ), .A2(new_n9641_), .ZN(new_n9642_));
  XOR2_X1    g09450(.A1(new_n9642_), .A2(new_n9591_), .Z(new_n9643_));
  NOR2_X1    g09451(.A1(new_n9643_), .A2(new_n196_), .ZN(new_n9644_));
  INV_X1     g09452(.I(new_n9644_), .ZN(new_n9645_));
  INV_X1     g09453(.I(\a[50] ), .ZN(new_n9646_));
  NOR2_X1    g09454(.A1(\a[48] ), .A2(\a[49] ), .ZN(new_n9647_));
  INV_X1     g09455(.I(new_n9647_), .ZN(new_n9648_));
  NOR3_X1    g09456(.A1(new_n9213_), .A2(new_n9646_), .A3(new_n9648_), .ZN(new_n9649_));
  NAND3_X1   g09457(.A1(new_n9164_), .A2(new_n9200_), .A3(new_n9649_), .ZN(new_n9650_));
  XOR2_X1    g09458(.A1(new_n9650_), .A2(\a[51] ), .Z(new_n9651_));
  INV_X1     g09459(.I(\a[51] ), .ZN(new_n9652_));
  NOR4_X1    g09460(.A1(new_n9625_), .A2(new_n9624_), .A3(new_n9652_), .A4(new_n9612_), .ZN(new_n9653_));
  NOR2_X1    g09461(.A1(new_n9651_), .A2(\a[50] ), .ZN(new_n9654_));
  OAI21_X1   g09462(.A1(new_n9653_), .A2(new_n9654_), .B(new_n9651_), .ZN(new_n9655_));
  INV_X1     g09463(.I(new_n9651_), .ZN(new_n9656_));
  NOR2_X1    g09464(.A1(new_n9602_), .A2(new_n9588_), .ZN(new_n9657_));
  NOR3_X1    g09465(.A1(new_n9603_), .A2(new_n229_), .A3(new_n9593_), .ZN(new_n9658_));
  AOI21_X1   g09466(.A1(new_n9658_), .A2(new_n9657_), .B(new_n9183_), .ZN(new_n9659_));
  AOI21_X1   g09467(.A1(new_n9659_), .A2(new_n9599_), .B(new_n9174_), .ZN(new_n9660_));
  AOI21_X1   g09468(.A1(new_n9604_), .A2(\asqrt[62] ), .B(new_n9175_), .ZN(new_n9661_));
  NOR3_X1    g09469(.A1(new_n9661_), .A2(new_n9633_), .A3(new_n9610_), .ZN(new_n9662_));
  NAND4_X1   g09470(.A1(new_n9662_), .A2(\a[51] ), .A3(new_n9660_), .A4(new_n9613_), .ZN(new_n9663_));
  NAND3_X1   g09471(.A1(new_n9663_), .A2(\a[50] ), .A3(new_n9656_), .ZN(new_n9664_));
  NAND2_X1   g09472(.A1(new_n9655_), .A2(new_n9664_), .ZN(new_n9665_));
  NAND2_X1   g09473(.A1(new_n9198_), .A2(new_n9162_), .ZN(new_n9666_));
  NAND4_X1   g09474(.A1(new_n9202_), .A2(new_n9196_), .A3(new_n9151_), .A4(new_n9666_), .ZN(new_n9667_));
  NOR2_X1    g09475(.A1(new_n9212_), .A2(new_n9646_), .ZN(new_n9668_));
  XOR2_X1    g09476(.A1(new_n9668_), .A2(new_n9667_), .Z(new_n9669_));
  NOR2_X1    g09477(.A1(new_n9669_), .A2(new_n9648_), .ZN(new_n9670_));
  INV_X1     g09478(.I(new_n9670_), .ZN(new_n9671_));
  NAND3_X1   g09479(.A1(new_n9662_), .A2(new_n9660_), .A3(new_n9613_), .ZN(new_n9672_));
  NOR4_X1    g09480(.A1(new_n9632_), .A2(new_n9588_), .A3(new_n9602_), .A4(new_n9593_), .ZN(new_n9673_));
  NOR3_X1    g09481(.A1(new_n9673_), .A2(new_n9183_), .A3(new_n9598_), .ZN(new_n9674_));
  NAND4_X1   g09482(.A1(new_n9629_), .A2(new_n196_), .A3(new_n9175_), .A4(new_n9592_), .ZN(new_n9675_));
  OAI21_X1   g09483(.A1(new_n9674_), .A2(new_n9174_), .B(new_n9675_), .ZN(new_n9676_));
  NAND2_X1   g09484(.A1(new_n9614_), .A2(\asqrt[26] ), .ZN(new_n9677_));
  OAI21_X1   g09485(.A1(new_n9676_), .A2(new_n9677_), .B(new_n9185_), .ZN(new_n9678_));
  NAND3_X1   g09486(.A1(new_n9678_), .A2(new_n9186_), .A3(new_n9672_), .ZN(new_n9679_));
  INV_X1     g09487(.I(new_n9677_), .ZN(new_n9680_));
  AOI21_X1   g09488(.A1(new_n9606_), .A2(new_n9680_), .B(\a[52] ), .ZN(new_n9681_));
  OAI21_X1   g09489(.A1(new_n9681_), .A2(new_n9187_), .B(\asqrt[25] ), .ZN(new_n9682_));
  NAND4_X1   g09490(.A1(new_n9679_), .A2(new_n9682_), .A3(new_n8763_), .A4(new_n9671_), .ZN(new_n9683_));
  NAND2_X1   g09491(.A1(new_n9683_), .A2(new_n9665_), .ZN(new_n9684_));
  NAND3_X1   g09492(.A1(new_n9655_), .A2(new_n9664_), .A3(new_n9671_), .ZN(new_n9685_));
  AOI21_X1   g09493(.A1(\asqrt[26] ), .A2(new_n9185_), .B(\a[53] ), .ZN(new_n9686_));
  NOR2_X1    g09494(.A1(new_n9203_), .A2(\a[52] ), .ZN(new_n9687_));
  AOI21_X1   g09495(.A1(\asqrt[26] ), .A2(\a[52] ), .B(new_n9189_), .ZN(new_n9688_));
  OAI21_X1   g09496(.A1(new_n9686_), .A2(new_n9687_), .B(new_n9688_), .ZN(new_n9689_));
  INV_X1     g09497(.I(new_n9689_), .ZN(new_n9690_));
  NAND3_X1   g09498(.A1(\asqrt[25] ), .A2(new_n9211_), .A3(new_n9690_), .ZN(new_n9691_));
  OAI21_X1   g09499(.A1(new_n9672_), .A2(new_n9689_), .B(new_n9210_), .ZN(new_n9692_));
  NAND3_X1   g09500(.A1(new_n9691_), .A2(new_n9692_), .A3(new_n8319_), .ZN(new_n9693_));
  AOI21_X1   g09501(.A1(new_n9685_), .A2(\asqrt[27] ), .B(new_n9693_), .ZN(new_n9694_));
  NOR2_X1    g09502(.A1(new_n9684_), .A2(new_n9694_), .ZN(new_n9695_));
  AOI22_X1   g09503(.A1(new_n9683_), .A2(new_n9665_), .B1(\asqrt[27] ), .B2(new_n9685_), .ZN(new_n9696_));
  INV_X1     g09504(.I(new_n9193_), .ZN(new_n9697_));
  AOI21_X1   g09505(.A1(new_n9203_), .A2(new_n9697_), .B(new_n9195_), .ZN(new_n9698_));
  INV_X1     g09506(.I(new_n9204_), .ZN(new_n9699_));
  NOR3_X1    g09507(.A1(new_n9699_), .A2(new_n9698_), .A3(new_n9210_), .ZN(new_n9700_));
  AOI21_X1   g09508(.A1(new_n9221_), .A2(new_n9218_), .B(\asqrt[28] ), .ZN(new_n9701_));
  AND4_X2    g09509(.A1(new_n9700_), .A2(\asqrt[25] ), .A3(new_n9235_), .A4(new_n9701_), .Z(new_n9702_));
  NOR2_X1    g09510(.A1(new_n9700_), .A2(new_n8319_), .ZN(new_n9703_));
  NOR3_X1    g09511(.A1(new_n9702_), .A2(\asqrt[29] ), .A3(new_n9703_), .ZN(new_n9704_));
  OAI21_X1   g09512(.A1(new_n9696_), .A2(new_n8319_), .B(new_n9704_), .ZN(new_n9705_));
  NAND2_X1   g09513(.A1(new_n9705_), .A2(new_n9695_), .ZN(new_n9706_));
  OAI22_X1   g09514(.A1(new_n9696_), .A2(new_n8319_), .B1(new_n9684_), .B2(new_n9694_), .ZN(new_n9707_));
  NAND2_X1   g09515(.A1(new_n9230_), .A2(new_n9231_), .ZN(new_n9708_));
  NAND4_X1   g09516(.A1(\asqrt[25] ), .A2(new_n7931_), .A3(new_n9708_), .A4(new_n9243_), .ZN(new_n9709_));
  XOR2_X1    g09517(.A1(new_n9709_), .A2(new_n9236_), .Z(new_n9710_));
  NAND2_X1   g09518(.A1(new_n9710_), .A2(new_n7517_), .ZN(new_n9711_));
  AOI21_X1   g09519(.A1(new_n9707_), .A2(\asqrt[29] ), .B(new_n9711_), .ZN(new_n9712_));
  NOR2_X1    g09520(.A1(new_n9712_), .A2(new_n9706_), .ZN(new_n9713_));
  AOI22_X1   g09521(.A1(new_n9707_), .A2(\asqrt[29] ), .B1(new_n9705_), .B2(new_n9695_), .ZN(new_n9714_));
  NOR4_X1    g09522(.A1(new_n9672_), .A2(\asqrt[30] ), .A3(new_n9240_), .A4(new_n9244_), .ZN(new_n9715_));
  XOR2_X1    g09523(.A1(new_n9715_), .A2(new_n9251_), .Z(new_n9716_));
  NAND2_X1   g09524(.A1(new_n9716_), .A2(new_n7110_), .ZN(new_n9717_));
  INV_X1     g09525(.I(new_n9717_), .ZN(new_n9718_));
  OAI21_X1   g09526(.A1(new_n9714_), .A2(new_n7517_), .B(new_n9718_), .ZN(new_n9719_));
  NAND2_X1   g09527(.A1(new_n9719_), .A2(new_n9713_), .ZN(new_n9720_));
  OAI22_X1   g09528(.A1(new_n9714_), .A2(new_n7517_), .B1(new_n9712_), .B2(new_n9706_), .ZN(new_n9721_));
  NAND2_X1   g09529(.A1(new_n9242_), .A2(new_n9251_), .ZN(new_n9722_));
  NOR4_X1    g09530(.A1(new_n9672_), .A2(\asqrt[31] ), .A3(new_n9248_), .A4(new_n9722_), .ZN(new_n9723_));
  XNOR2_X1   g09531(.A1(new_n9723_), .A2(new_n9252_), .ZN(new_n9724_));
  NAND2_X1   g09532(.A1(new_n9724_), .A2(new_n6708_), .ZN(new_n9725_));
  AOI21_X1   g09533(.A1(new_n9721_), .A2(\asqrt[31] ), .B(new_n9725_), .ZN(new_n9726_));
  NOR2_X1    g09534(.A1(new_n9726_), .A2(new_n9720_), .ZN(new_n9727_));
  AOI22_X1   g09535(.A1(new_n9721_), .A2(\asqrt[31] ), .B1(new_n9719_), .B2(new_n9713_), .ZN(new_n9728_));
  NOR4_X1    g09536(.A1(new_n9672_), .A2(\asqrt[32] ), .A3(new_n9256_), .A4(new_n9482_), .ZN(new_n9729_));
  XOR2_X1    g09537(.A1(new_n9729_), .A2(new_n9262_), .Z(new_n9730_));
  NAND2_X1   g09538(.A1(new_n9730_), .A2(new_n6365_), .ZN(new_n9731_));
  INV_X1     g09539(.I(new_n9731_), .ZN(new_n9732_));
  OAI21_X1   g09540(.A1(new_n9728_), .A2(new_n6708_), .B(new_n9732_), .ZN(new_n9733_));
  NAND2_X1   g09541(.A1(new_n9733_), .A2(new_n9727_), .ZN(new_n9734_));
  OAI22_X1   g09542(.A1(new_n9728_), .A2(new_n6708_), .B1(new_n9726_), .B2(new_n9720_), .ZN(new_n9735_));
  NOR4_X1    g09543(.A1(new_n9672_), .A2(\asqrt[33] ), .A3(new_n9265_), .A4(new_n9271_), .ZN(new_n9736_));
  XNOR2_X1   g09544(.A1(new_n9736_), .A2(new_n9279_), .ZN(new_n9737_));
  NAND2_X1   g09545(.A1(new_n9737_), .A2(new_n5991_), .ZN(new_n9738_));
  AOI21_X1   g09546(.A1(new_n9735_), .A2(\asqrt[33] ), .B(new_n9738_), .ZN(new_n9739_));
  NOR2_X1    g09547(.A1(new_n9739_), .A2(new_n9734_), .ZN(new_n9740_));
  AOI22_X1   g09548(.A1(new_n9735_), .A2(\asqrt[33] ), .B1(new_n9733_), .B2(new_n9727_), .ZN(new_n9741_));
  NOR4_X1    g09549(.A1(new_n9672_), .A2(\asqrt[34] ), .A3(new_n9274_), .A4(new_n9488_), .ZN(new_n9742_));
  XOR2_X1    g09550(.A1(new_n9742_), .A2(new_n9280_), .Z(new_n9743_));
  NAND2_X1   g09551(.A1(new_n9743_), .A2(new_n5626_), .ZN(new_n9744_));
  INV_X1     g09552(.I(new_n9744_), .ZN(new_n9745_));
  OAI21_X1   g09553(.A1(new_n9741_), .A2(new_n5991_), .B(new_n9745_), .ZN(new_n9746_));
  NAND2_X1   g09554(.A1(new_n9746_), .A2(new_n9740_), .ZN(new_n9747_));
  OAI22_X1   g09555(.A1(new_n9741_), .A2(new_n5991_), .B1(new_n9739_), .B2(new_n9734_), .ZN(new_n9748_));
  NAND2_X1   g09556(.A1(new_n9289_), .A2(\asqrt[35] ), .ZN(new_n9749_));
  NOR4_X1    g09557(.A1(new_n9672_), .A2(\asqrt[35] ), .A3(new_n9283_), .A4(new_n9289_), .ZN(new_n9750_));
  XOR2_X1    g09558(.A1(new_n9750_), .A2(new_n9749_), .Z(new_n9751_));
  NAND2_X1   g09559(.A1(new_n9751_), .A2(new_n5273_), .ZN(new_n9752_));
  AOI21_X1   g09560(.A1(new_n9748_), .A2(\asqrt[35] ), .B(new_n9752_), .ZN(new_n9753_));
  NOR2_X1    g09561(.A1(new_n9753_), .A2(new_n9747_), .ZN(new_n9754_));
  AOI22_X1   g09562(.A1(new_n9748_), .A2(\asqrt[35] ), .B1(new_n9746_), .B2(new_n9740_), .ZN(new_n9755_));
  NOR4_X1    g09563(.A1(new_n9672_), .A2(\asqrt[36] ), .A3(new_n9292_), .A4(new_n9495_), .ZN(new_n9756_));
  AOI21_X1   g09564(.A1(new_n9749_), .A2(new_n9287_), .B(new_n5273_), .ZN(new_n9757_));
  NOR2_X1    g09565(.A1(new_n9756_), .A2(new_n9757_), .ZN(new_n9758_));
  NAND2_X1   g09566(.A1(new_n9758_), .A2(new_n4973_), .ZN(new_n9759_));
  INV_X1     g09567(.I(new_n9759_), .ZN(new_n9760_));
  OAI21_X1   g09568(.A1(new_n9755_), .A2(new_n5273_), .B(new_n9760_), .ZN(new_n9761_));
  NAND2_X1   g09569(.A1(new_n9761_), .A2(new_n9754_), .ZN(new_n9762_));
  OAI22_X1   g09570(.A1(new_n9755_), .A2(new_n5273_), .B1(new_n9753_), .B2(new_n9747_), .ZN(new_n9763_));
  NAND2_X1   g09571(.A1(new_n9304_), .A2(\asqrt[37] ), .ZN(new_n9764_));
  NOR4_X1    g09572(.A1(new_n9672_), .A2(\asqrt[37] ), .A3(new_n9299_), .A4(new_n9304_), .ZN(new_n9765_));
  XOR2_X1    g09573(.A1(new_n9765_), .A2(new_n9764_), .Z(new_n9766_));
  NAND2_X1   g09574(.A1(new_n9766_), .A2(new_n4645_), .ZN(new_n9767_));
  AOI21_X1   g09575(.A1(new_n9763_), .A2(\asqrt[37] ), .B(new_n9767_), .ZN(new_n9768_));
  NOR2_X1    g09576(.A1(new_n9768_), .A2(new_n9762_), .ZN(new_n9769_));
  AOI22_X1   g09577(.A1(new_n9763_), .A2(\asqrt[37] ), .B1(new_n9761_), .B2(new_n9754_), .ZN(new_n9770_));
  NOR4_X1    g09578(.A1(new_n9672_), .A2(\asqrt[38] ), .A3(new_n9307_), .A4(new_n9502_), .ZN(new_n9771_));
  AOI21_X1   g09579(.A1(new_n9764_), .A2(new_n9303_), .B(new_n4645_), .ZN(new_n9772_));
  NOR2_X1    g09580(.A1(new_n9771_), .A2(new_n9772_), .ZN(new_n9773_));
  NAND2_X1   g09581(.A1(new_n9773_), .A2(new_n4330_), .ZN(new_n9774_));
  INV_X1     g09582(.I(new_n9774_), .ZN(new_n9775_));
  OAI21_X1   g09583(.A1(new_n9770_), .A2(new_n4645_), .B(new_n9775_), .ZN(new_n9776_));
  NAND2_X1   g09584(.A1(new_n9776_), .A2(new_n9769_), .ZN(new_n9777_));
  OAI22_X1   g09585(.A1(new_n9770_), .A2(new_n4645_), .B1(new_n9768_), .B2(new_n9762_), .ZN(new_n9778_));
  NAND2_X1   g09586(.A1(new_n9319_), .A2(\asqrt[39] ), .ZN(new_n9779_));
  NOR4_X1    g09587(.A1(new_n9672_), .A2(\asqrt[39] ), .A3(new_n9314_), .A4(new_n9319_), .ZN(new_n9780_));
  XOR2_X1    g09588(.A1(new_n9780_), .A2(new_n9779_), .Z(new_n9781_));
  NAND2_X1   g09589(.A1(new_n9781_), .A2(new_n4018_), .ZN(new_n9782_));
  AOI21_X1   g09590(.A1(new_n9778_), .A2(\asqrt[39] ), .B(new_n9782_), .ZN(new_n9783_));
  NOR2_X1    g09591(.A1(new_n9783_), .A2(new_n9777_), .ZN(new_n9784_));
  AOI22_X1   g09592(.A1(new_n9778_), .A2(\asqrt[39] ), .B1(new_n9776_), .B2(new_n9769_), .ZN(new_n9785_));
  NOR4_X1    g09593(.A1(new_n9672_), .A2(\asqrt[40] ), .A3(new_n9322_), .A4(new_n9509_), .ZN(new_n9786_));
  AOI21_X1   g09594(.A1(new_n9779_), .A2(new_n9318_), .B(new_n4018_), .ZN(new_n9787_));
  NOR2_X1    g09595(.A1(new_n9786_), .A2(new_n9787_), .ZN(new_n9788_));
  NAND2_X1   g09596(.A1(new_n9788_), .A2(new_n3760_), .ZN(new_n9789_));
  INV_X1     g09597(.I(new_n9789_), .ZN(new_n9790_));
  OAI21_X1   g09598(.A1(new_n9785_), .A2(new_n4018_), .B(new_n9790_), .ZN(new_n9791_));
  NAND2_X1   g09599(.A1(new_n9791_), .A2(new_n9784_), .ZN(new_n9792_));
  OAI22_X1   g09600(.A1(new_n9785_), .A2(new_n4018_), .B1(new_n9783_), .B2(new_n9777_), .ZN(new_n9793_));
  NAND2_X1   g09601(.A1(new_n9334_), .A2(\asqrt[41] ), .ZN(new_n9794_));
  NOR4_X1    g09602(.A1(new_n9672_), .A2(\asqrt[41] ), .A3(new_n9329_), .A4(new_n9334_), .ZN(new_n9795_));
  XOR2_X1    g09603(.A1(new_n9795_), .A2(new_n9794_), .Z(new_n9796_));
  NAND2_X1   g09604(.A1(new_n9796_), .A2(new_n3481_), .ZN(new_n9797_));
  AOI21_X1   g09605(.A1(new_n9793_), .A2(\asqrt[41] ), .B(new_n9797_), .ZN(new_n9798_));
  NOR2_X1    g09606(.A1(new_n9798_), .A2(new_n9792_), .ZN(new_n9799_));
  AOI22_X1   g09607(.A1(new_n9793_), .A2(\asqrt[41] ), .B1(new_n9791_), .B2(new_n9784_), .ZN(new_n9800_));
  NOR4_X1    g09608(.A1(new_n9672_), .A2(\asqrt[42] ), .A3(new_n9337_), .A4(new_n9516_), .ZN(new_n9801_));
  AOI21_X1   g09609(.A1(new_n9794_), .A2(new_n9333_), .B(new_n3481_), .ZN(new_n9802_));
  NOR2_X1    g09610(.A1(new_n9801_), .A2(new_n9802_), .ZN(new_n9803_));
  NAND2_X1   g09611(.A1(new_n9803_), .A2(new_n3208_), .ZN(new_n9804_));
  INV_X1     g09612(.I(new_n9804_), .ZN(new_n9805_));
  OAI21_X1   g09613(.A1(new_n9800_), .A2(new_n3481_), .B(new_n9805_), .ZN(new_n9806_));
  NAND2_X1   g09614(.A1(new_n9806_), .A2(new_n9799_), .ZN(new_n9807_));
  OAI22_X1   g09615(.A1(new_n9800_), .A2(new_n3481_), .B1(new_n9798_), .B2(new_n9792_), .ZN(new_n9808_));
  NAND2_X1   g09616(.A1(new_n9349_), .A2(\asqrt[43] ), .ZN(new_n9809_));
  NOR4_X1    g09617(.A1(new_n9672_), .A2(\asqrt[43] ), .A3(new_n9344_), .A4(new_n9349_), .ZN(new_n9810_));
  XOR2_X1    g09618(.A1(new_n9810_), .A2(new_n9809_), .Z(new_n9811_));
  NAND2_X1   g09619(.A1(new_n9811_), .A2(new_n2941_), .ZN(new_n9812_));
  AOI21_X1   g09620(.A1(new_n9808_), .A2(\asqrt[43] ), .B(new_n9812_), .ZN(new_n9813_));
  NOR2_X1    g09621(.A1(new_n9813_), .A2(new_n9807_), .ZN(new_n9814_));
  AOI22_X1   g09622(.A1(new_n9808_), .A2(\asqrt[43] ), .B1(new_n9806_), .B2(new_n9799_), .ZN(new_n9815_));
  NOR4_X1    g09623(.A1(new_n9672_), .A2(\asqrt[44] ), .A3(new_n9352_), .A4(new_n9523_), .ZN(new_n9816_));
  AOI21_X1   g09624(.A1(new_n9809_), .A2(new_n9348_), .B(new_n2941_), .ZN(new_n9817_));
  NOR2_X1    g09625(.A1(new_n9816_), .A2(new_n9817_), .ZN(new_n9818_));
  NAND2_X1   g09626(.A1(new_n9818_), .A2(new_n2728_), .ZN(new_n9819_));
  INV_X1     g09627(.I(new_n9819_), .ZN(new_n9820_));
  OAI21_X1   g09628(.A1(new_n9815_), .A2(new_n2941_), .B(new_n9820_), .ZN(new_n9821_));
  NAND2_X1   g09629(.A1(new_n9821_), .A2(new_n9814_), .ZN(new_n9822_));
  OAI22_X1   g09630(.A1(new_n9815_), .A2(new_n2941_), .B1(new_n9813_), .B2(new_n9807_), .ZN(new_n9823_));
  NAND2_X1   g09631(.A1(new_n9364_), .A2(\asqrt[45] ), .ZN(new_n9824_));
  NOR4_X1    g09632(.A1(new_n9672_), .A2(\asqrt[45] ), .A3(new_n9359_), .A4(new_n9364_), .ZN(new_n9825_));
  XOR2_X1    g09633(.A1(new_n9825_), .A2(new_n9824_), .Z(new_n9826_));
  NAND2_X1   g09634(.A1(new_n9826_), .A2(new_n2488_), .ZN(new_n9827_));
  AOI21_X1   g09635(.A1(new_n9823_), .A2(\asqrt[45] ), .B(new_n9827_), .ZN(new_n9828_));
  NOR2_X1    g09636(.A1(new_n9828_), .A2(new_n9822_), .ZN(new_n9829_));
  AOI22_X1   g09637(.A1(new_n9823_), .A2(\asqrt[45] ), .B1(new_n9821_), .B2(new_n9814_), .ZN(new_n9830_));
  NAND2_X1   g09638(.A1(new_n9530_), .A2(\asqrt[46] ), .ZN(new_n9831_));
  NOR4_X1    g09639(.A1(new_n9672_), .A2(\asqrt[46] ), .A3(new_n9367_), .A4(new_n9530_), .ZN(new_n9832_));
  XOR2_X1    g09640(.A1(new_n9832_), .A2(new_n9831_), .Z(new_n9833_));
  NAND2_X1   g09641(.A1(new_n9833_), .A2(new_n2253_), .ZN(new_n9834_));
  INV_X1     g09642(.I(new_n9834_), .ZN(new_n9835_));
  OAI21_X1   g09643(.A1(new_n9830_), .A2(new_n2488_), .B(new_n9835_), .ZN(new_n9836_));
  NAND2_X1   g09644(.A1(new_n9836_), .A2(new_n9829_), .ZN(new_n9837_));
  OAI22_X1   g09645(.A1(new_n9830_), .A2(new_n2488_), .B1(new_n9828_), .B2(new_n9822_), .ZN(new_n9838_));
  NOR4_X1    g09646(.A1(new_n9672_), .A2(\asqrt[47] ), .A3(new_n9374_), .A4(new_n9379_), .ZN(new_n9839_));
  AOI21_X1   g09647(.A1(new_n9831_), .A2(new_n9529_), .B(new_n2253_), .ZN(new_n9840_));
  NOR2_X1    g09648(.A1(new_n9839_), .A2(new_n9840_), .ZN(new_n9841_));
  NAND2_X1   g09649(.A1(new_n9841_), .A2(new_n2046_), .ZN(new_n9842_));
  AOI21_X1   g09650(.A1(new_n9838_), .A2(\asqrt[47] ), .B(new_n9842_), .ZN(new_n9843_));
  NOR2_X1    g09651(.A1(new_n9843_), .A2(new_n9837_), .ZN(new_n9844_));
  AOI22_X1   g09652(.A1(new_n9838_), .A2(\asqrt[47] ), .B1(new_n9836_), .B2(new_n9829_), .ZN(new_n9845_));
  NAND2_X1   g09653(.A1(new_n9537_), .A2(\asqrt[48] ), .ZN(new_n9846_));
  NOR4_X1    g09654(.A1(new_n9672_), .A2(\asqrt[48] ), .A3(new_n9382_), .A4(new_n9537_), .ZN(new_n9847_));
  XOR2_X1    g09655(.A1(new_n9847_), .A2(new_n9846_), .Z(new_n9848_));
  NAND2_X1   g09656(.A1(new_n9848_), .A2(new_n1854_), .ZN(new_n9849_));
  INV_X1     g09657(.I(new_n9849_), .ZN(new_n9850_));
  OAI21_X1   g09658(.A1(new_n9845_), .A2(new_n2046_), .B(new_n9850_), .ZN(new_n9851_));
  NAND2_X1   g09659(.A1(new_n9851_), .A2(new_n9844_), .ZN(new_n9852_));
  OAI22_X1   g09660(.A1(new_n9845_), .A2(new_n2046_), .B1(new_n9843_), .B2(new_n9837_), .ZN(new_n9853_));
  NOR4_X1    g09661(.A1(new_n9672_), .A2(\asqrt[49] ), .A3(new_n9389_), .A4(new_n9394_), .ZN(new_n9854_));
  AOI21_X1   g09662(.A1(new_n9846_), .A2(new_n9536_), .B(new_n1854_), .ZN(new_n9855_));
  NOR2_X1    g09663(.A1(new_n9854_), .A2(new_n9855_), .ZN(new_n9856_));
  NAND2_X1   g09664(.A1(new_n9856_), .A2(new_n1595_), .ZN(new_n9857_));
  AOI21_X1   g09665(.A1(new_n9853_), .A2(\asqrt[49] ), .B(new_n9857_), .ZN(new_n9858_));
  NOR2_X1    g09666(.A1(new_n9858_), .A2(new_n9852_), .ZN(new_n9859_));
  AOI22_X1   g09667(.A1(new_n9853_), .A2(\asqrt[49] ), .B1(new_n9851_), .B2(new_n9844_), .ZN(new_n9860_));
  NAND2_X1   g09668(.A1(new_n9544_), .A2(\asqrt[50] ), .ZN(new_n9861_));
  NOR4_X1    g09669(.A1(new_n9672_), .A2(\asqrt[50] ), .A3(new_n9397_), .A4(new_n9544_), .ZN(new_n9862_));
  XOR2_X1    g09670(.A1(new_n9862_), .A2(new_n9861_), .Z(new_n9863_));
  NAND2_X1   g09671(.A1(new_n9863_), .A2(new_n1436_), .ZN(new_n9864_));
  INV_X1     g09672(.I(new_n9864_), .ZN(new_n9865_));
  OAI21_X1   g09673(.A1(new_n9860_), .A2(new_n1595_), .B(new_n9865_), .ZN(new_n9866_));
  NAND2_X1   g09674(.A1(new_n9866_), .A2(new_n9859_), .ZN(new_n9867_));
  OAI22_X1   g09675(.A1(new_n9860_), .A2(new_n1595_), .B1(new_n9858_), .B2(new_n9852_), .ZN(new_n9868_));
  NAND2_X1   g09676(.A1(new_n9409_), .A2(\asqrt[51] ), .ZN(new_n9869_));
  NOR4_X1    g09677(.A1(new_n9672_), .A2(\asqrt[51] ), .A3(new_n9404_), .A4(new_n9409_), .ZN(new_n9870_));
  XOR2_X1    g09678(.A1(new_n9870_), .A2(new_n9869_), .Z(new_n9871_));
  NAND2_X1   g09679(.A1(new_n9871_), .A2(new_n1260_), .ZN(new_n9872_));
  AOI21_X1   g09680(.A1(new_n9868_), .A2(\asqrt[51] ), .B(new_n9872_), .ZN(new_n9873_));
  NOR2_X1    g09681(.A1(new_n9873_), .A2(new_n9867_), .ZN(new_n9874_));
  AOI22_X1   g09682(.A1(new_n9868_), .A2(\asqrt[51] ), .B1(new_n9866_), .B2(new_n9859_), .ZN(new_n9875_));
  NOR4_X1    g09683(.A1(new_n9672_), .A2(\asqrt[52] ), .A3(new_n9412_), .A4(new_n9551_), .ZN(new_n9876_));
  AOI21_X1   g09684(.A1(new_n9869_), .A2(new_n9408_), .B(new_n1260_), .ZN(new_n9877_));
  NOR2_X1    g09685(.A1(new_n9876_), .A2(new_n9877_), .ZN(new_n9878_));
  NAND2_X1   g09686(.A1(new_n9878_), .A2(new_n1096_), .ZN(new_n9879_));
  INV_X1     g09687(.I(new_n9879_), .ZN(new_n9880_));
  OAI21_X1   g09688(.A1(new_n9875_), .A2(new_n1260_), .B(new_n9880_), .ZN(new_n9881_));
  NAND2_X1   g09689(.A1(new_n9881_), .A2(new_n9874_), .ZN(new_n9882_));
  OAI22_X1   g09690(.A1(new_n9875_), .A2(new_n1260_), .B1(new_n9873_), .B2(new_n9867_), .ZN(new_n9883_));
  NOR2_X1    g09691(.A1(new_n9554_), .A2(new_n1096_), .ZN(new_n9884_));
  NOR4_X1    g09692(.A1(new_n9672_), .A2(\asqrt[53] ), .A3(new_n9419_), .A4(new_n9424_), .ZN(new_n9885_));
  XNOR2_X1   g09693(.A1(new_n9885_), .A2(new_n9884_), .ZN(new_n9886_));
  NAND2_X1   g09694(.A1(new_n9886_), .A2(new_n970_), .ZN(new_n9887_));
  AOI21_X1   g09695(.A1(new_n9883_), .A2(\asqrt[53] ), .B(new_n9887_), .ZN(new_n9888_));
  NOR2_X1    g09696(.A1(new_n9888_), .A2(new_n9882_), .ZN(new_n9889_));
  AOI22_X1   g09697(.A1(new_n9883_), .A2(\asqrt[53] ), .B1(new_n9881_), .B2(new_n9874_), .ZN(new_n9890_));
  NOR4_X1    g09698(.A1(new_n9672_), .A2(\asqrt[54] ), .A3(new_n9427_), .A4(new_n9558_), .ZN(new_n9891_));
  XOR2_X1    g09699(.A1(new_n9891_), .A2(new_n9571_), .Z(new_n9892_));
  NAND2_X1   g09700(.A1(new_n9892_), .A2(new_n825_), .ZN(new_n9893_));
  INV_X1     g09701(.I(new_n9893_), .ZN(new_n9894_));
  OAI21_X1   g09702(.A1(new_n9890_), .A2(new_n970_), .B(new_n9894_), .ZN(new_n9895_));
  NAND2_X1   g09703(.A1(new_n9895_), .A2(new_n9889_), .ZN(new_n9896_));
  OAI22_X1   g09704(.A1(new_n9890_), .A2(new_n970_), .B1(new_n9888_), .B2(new_n9882_), .ZN(new_n9897_));
  NOR4_X1    g09705(.A1(new_n9672_), .A2(\asqrt[55] ), .A3(new_n9434_), .A4(new_n9439_), .ZN(new_n9898_));
  XOR2_X1    g09706(.A1(new_n9898_), .A2(new_n9454_), .Z(new_n9899_));
  NAND2_X1   g09707(.A1(new_n9899_), .A2(new_n724_), .ZN(new_n9900_));
  AOI21_X1   g09708(.A1(new_n9897_), .A2(\asqrt[55] ), .B(new_n9900_), .ZN(new_n9901_));
  NOR2_X1    g09709(.A1(new_n9901_), .A2(new_n9896_), .ZN(new_n9902_));
  AOI22_X1   g09710(.A1(new_n9897_), .A2(\asqrt[55] ), .B1(new_n9895_), .B2(new_n9889_), .ZN(new_n9903_));
  NOR4_X1    g09711(.A1(new_n9672_), .A2(\asqrt[56] ), .A3(new_n9442_), .A4(new_n9565_), .ZN(new_n9904_));
  XOR2_X1    g09712(.A1(new_n9904_), .A2(new_n9573_), .Z(new_n9905_));
  NAND2_X1   g09713(.A1(new_n9905_), .A2(new_n587_), .ZN(new_n9906_));
  INV_X1     g09714(.I(new_n9906_), .ZN(new_n9907_));
  OAI21_X1   g09715(.A1(new_n9903_), .A2(new_n724_), .B(new_n9907_), .ZN(new_n9908_));
  NAND2_X1   g09716(.A1(new_n9908_), .A2(new_n9902_), .ZN(new_n9909_));
  OAI22_X1   g09717(.A1(new_n9903_), .A2(new_n724_), .B1(new_n9901_), .B2(new_n9896_), .ZN(new_n9910_));
  NOR4_X1    g09718(.A1(new_n9672_), .A2(\asqrt[57] ), .A3(new_n9449_), .A4(new_n9463_), .ZN(new_n9911_));
  XOR2_X1    g09719(.A1(new_n9911_), .A2(new_n9456_), .Z(new_n9912_));
  NAND2_X1   g09720(.A1(new_n9912_), .A2(new_n504_), .ZN(new_n9913_));
  AOI21_X1   g09721(.A1(new_n9910_), .A2(\asqrt[57] ), .B(new_n9913_), .ZN(new_n9914_));
  NOR2_X1    g09722(.A1(new_n9914_), .A2(new_n9909_), .ZN(new_n9915_));
  AOI22_X1   g09723(.A1(new_n9910_), .A2(\asqrt[57] ), .B1(new_n9908_), .B2(new_n9902_), .ZN(new_n9916_));
  NOR4_X1    g09724(.A1(new_n9672_), .A2(\asqrt[58] ), .A3(new_n9459_), .A4(new_n9583_), .ZN(new_n9917_));
  XOR2_X1    g09725(.A1(new_n9917_), .A2(new_n9575_), .Z(new_n9918_));
  NAND2_X1   g09726(.A1(new_n9918_), .A2(new_n376_), .ZN(new_n9919_));
  INV_X1     g09727(.I(new_n9919_), .ZN(new_n9920_));
  OAI21_X1   g09728(.A1(new_n9916_), .A2(new_n504_), .B(new_n9920_), .ZN(new_n9921_));
  NAND2_X1   g09729(.A1(new_n9921_), .A2(new_n9915_), .ZN(new_n9922_));
  OAI22_X1   g09730(.A1(new_n9916_), .A2(new_n504_), .B1(new_n9914_), .B2(new_n9909_), .ZN(new_n9923_));
  NOR4_X1    g09731(.A1(new_n9672_), .A2(\asqrt[59] ), .A3(new_n9466_), .A4(new_n9576_), .ZN(new_n9924_));
  XOR2_X1    g09732(.A1(new_n9924_), .A2(new_n9472_), .Z(new_n9925_));
  NAND2_X1   g09733(.A1(new_n9925_), .A2(new_n275_), .ZN(new_n9926_));
  AOI21_X1   g09734(.A1(new_n9923_), .A2(\asqrt[59] ), .B(new_n9926_), .ZN(new_n9927_));
  NOR2_X1    g09735(.A1(new_n9927_), .A2(new_n9922_), .ZN(new_n9928_));
  AOI22_X1   g09736(.A1(new_n9923_), .A2(\asqrt[59] ), .B1(new_n9921_), .B2(new_n9915_), .ZN(new_n9929_));
  NOR4_X1    g09737(.A1(new_n9672_), .A2(\asqrt[60] ), .A3(new_n9474_), .A4(new_n9601_), .ZN(new_n9930_));
  XOR2_X1    g09738(.A1(new_n9930_), .A2(new_n9590_), .Z(new_n9931_));
  NAND2_X1   g09739(.A1(new_n9931_), .A2(new_n229_), .ZN(new_n9932_));
  INV_X1     g09740(.I(new_n9932_), .ZN(new_n9933_));
  OAI21_X1   g09741(.A1(new_n9929_), .A2(new_n275_), .B(new_n9933_), .ZN(new_n9934_));
  NAND2_X1   g09742(.A1(new_n9934_), .A2(new_n9928_), .ZN(new_n9935_));
  OAI22_X1   g09743(.A1(new_n9929_), .A2(new_n275_), .B1(new_n9927_), .B2(new_n9922_), .ZN(new_n9936_));
  INV_X1     g09744(.I(new_n9643_), .ZN(new_n9937_));
  NOR2_X1    g09745(.A1(new_n9937_), .A2(\asqrt[62] ), .ZN(new_n9938_));
  INV_X1     g09746(.I(new_n9938_), .ZN(new_n9939_));
  NAND3_X1   g09747(.A1(new_n9936_), .A2(\asqrt[61] ), .A3(new_n9939_), .ZN(new_n9940_));
  OAI21_X1   g09748(.A1(new_n9940_), .A2(new_n9935_), .B(new_n9645_), .ZN(new_n9941_));
  NAND3_X1   g09749(.A1(new_n9672_), .A2(new_n9174_), .A3(new_n9675_), .ZN(new_n9942_));
  AOI21_X1   g09750(.A1(new_n9942_), .A2(new_n9623_), .B(\asqrt[63] ), .ZN(new_n9943_));
  INV_X1     g09751(.I(new_n9943_), .ZN(new_n9944_));
  OAI21_X1   g09752(.A1(new_n9941_), .A2(new_n9944_), .B(new_n9640_), .ZN(new_n9945_));
  INV_X1     g09753(.I(new_n9654_), .ZN(new_n9946_));
  AOI21_X1   g09754(.A1(new_n9663_), .A2(new_n9946_), .B(new_n9656_), .ZN(new_n9947_));
  NOR3_X1    g09755(.A1(new_n9653_), .A2(new_n9646_), .A3(new_n9651_), .ZN(new_n9948_));
  NOR2_X1    g09756(.A1(new_n9948_), .A2(new_n9947_), .ZN(new_n9949_));
  NOR3_X1    g09757(.A1(new_n9681_), .A2(new_n9187_), .A3(\asqrt[25] ), .ZN(new_n9950_));
  AOI21_X1   g09758(.A1(new_n9678_), .A2(new_n9186_), .B(new_n9672_), .ZN(new_n9951_));
  NOR4_X1    g09759(.A1(new_n9951_), .A2(new_n9950_), .A3(\asqrt[27] ), .A4(new_n9670_), .ZN(new_n9952_));
  NOR2_X1    g09760(.A1(new_n9952_), .A2(new_n9949_), .ZN(new_n9953_));
  NOR3_X1    g09761(.A1(new_n9948_), .A2(new_n9947_), .A3(new_n9670_), .ZN(new_n9954_));
  NOR3_X1    g09762(.A1(new_n9672_), .A2(new_n9210_), .A3(new_n9689_), .ZN(new_n9955_));
  AOI21_X1   g09763(.A1(\asqrt[25] ), .A2(new_n9690_), .B(new_n9211_), .ZN(new_n9956_));
  NOR3_X1    g09764(.A1(new_n9956_), .A2(new_n9955_), .A3(\asqrt[28] ), .ZN(new_n9957_));
  OAI21_X1   g09765(.A1(new_n9954_), .A2(new_n8763_), .B(new_n9957_), .ZN(new_n9958_));
  NAND2_X1   g09766(.A1(new_n9953_), .A2(new_n9958_), .ZN(new_n9959_));
  OAI22_X1   g09767(.A1(new_n9952_), .A2(new_n9949_), .B1(new_n8763_), .B2(new_n9954_), .ZN(new_n9960_));
  INV_X1     g09768(.I(new_n9704_), .ZN(new_n9961_));
  AOI21_X1   g09769(.A1(new_n9960_), .A2(\asqrt[28] ), .B(new_n9961_), .ZN(new_n9962_));
  NOR2_X1    g09770(.A1(new_n9962_), .A2(new_n9959_), .ZN(new_n9963_));
  AOI22_X1   g09771(.A1(new_n9960_), .A2(\asqrt[28] ), .B1(new_n9953_), .B2(new_n9958_), .ZN(new_n9964_));
  INV_X1     g09772(.I(new_n9711_), .ZN(new_n9965_));
  OAI21_X1   g09773(.A1(new_n9964_), .A2(new_n7931_), .B(new_n9965_), .ZN(new_n9966_));
  NAND2_X1   g09774(.A1(new_n9966_), .A2(new_n9963_), .ZN(new_n9967_));
  OAI22_X1   g09775(.A1(new_n9964_), .A2(new_n7931_), .B1(new_n9962_), .B2(new_n9959_), .ZN(new_n9968_));
  AOI21_X1   g09776(.A1(new_n9968_), .A2(\asqrt[30] ), .B(new_n9717_), .ZN(new_n9969_));
  NOR2_X1    g09777(.A1(new_n9969_), .A2(new_n9967_), .ZN(new_n9970_));
  AOI22_X1   g09778(.A1(new_n9968_), .A2(\asqrt[30] ), .B1(new_n9966_), .B2(new_n9963_), .ZN(new_n9971_));
  INV_X1     g09779(.I(new_n9725_), .ZN(new_n9972_));
  OAI21_X1   g09780(.A1(new_n9971_), .A2(new_n7110_), .B(new_n9972_), .ZN(new_n9973_));
  NAND2_X1   g09781(.A1(new_n9973_), .A2(new_n9970_), .ZN(new_n9974_));
  OAI22_X1   g09782(.A1(new_n9971_), .A2(new_n7110_), .B1(new_n9969_), .B2(new_n9967_), .ZN(new_n9975_));
  AOI21_X1   g09783(.A1(new_n9975_), .A2(\asqrt[32] ), .B(new_n9731_), .ZN(new_n9976_));
  NOR2_X1    g09784(.A1(new_n9976_), .A2(new_n9974_), .ZN(new_n9977_));
  AOI22_X1   g09785(.A1(new_n9975_), .A2(\asqrt[32] ), .B1(new_n9973_), .B2(new_n9970_), .ZN(new_n9978_));
  INV_X1     g09786(.I(new_n9738_), .ZN(new_n9979_));
  OAI21_X1   g09787(.A1(new_n9978_), .A2(new_n6365_), .B(new_n9979_), .ZN(new_n9980_));
  NAND2_X1   g09788(.A1(new_n9980_), .A2(new_n9977_), .ZN(new_n9981_));
  OAI22_X1   g09789(.A1(new_n9978_), .A2(new_n6365_), .B1(new_n9976_), .B2(new_n9974_), .ZN(new_n9982_));
  AOI21_X1   g09790(.A1(new_n9982_), .A2(\asqrt[34] ), .B(new_n9744_), .ZN(new_n9983_));
  NOR2_X1    g09791(.A1(new_n9983_), .A2(new_n9981_), .ZN(new_n9984_));
  AOI22_X1   g09792(.A1(new_n9982_), .A2(\asqrt[34] ), .B1(new_n9980_), .B2(new_n9977_), .ZN(new_n9985_));
  INV_X1     g09793(.I(new_n9752_), .ZN(new_n9986_));
  OAI21_X1   g09794(.A1(new_n9985_), .A2(new_n5626_), .B(new_n9986_), .ZN(new_n9987_));
  NAND2_X1   g09795(.A1(new_n9987_), .A2(new_n9984_), .ZN(new_n9988_));
  OAI22_X1   g09796(.A1(new_n9985_), .A2(new_n5626_), .B1(new_n9983_), .B2(new_n9981_), .ZN(new_n9989_));
  AOI21_X1   g09797(.A1(new_n9989_), .A2(\asqrt[36] ), .B(new_n9759_), .ZN(new_n9990_));
  NOR2_X1    g09798(.A1(new_n9990_), .A2(new_n9988_), .ZN(new_n9991_));
  AOI22_X1   g09799(.A1(new_n9989_), .A2(\asqrt[36] ), .B1(new_n9987_), .B2(new_n9984_), .ZN(new_n9992_));
  INV_X1     g09800(.I(new_n9767_), .ZN(new_n9993_));
  OAI21_X1   g09801(.A1(new_n9992_), .A2(new_n4973_), .B(new_n9993_), .ZN(new_n9994_));
  NAND2_X1   g09802(.A1(new_n9994_), .A2(new_n9991_), .ZN(new_n9995_));
  OAI22_X1   g09803(.A1(new_n9992_), .A2(new_n4973_), .B1(new_n9990_), .B2(new_n9988_), .ZN(new_n9996_));
  AOI21_X1   g09804(.A1(new_n9996_), .A2(\asqrt[38] ), .B(new_n9774_), .ZN(new_n9997_));
  NOR2_X1    g09805(.A1(new_n9997_), .A2(new_n9995_), .ZN(new_n9998_));
  AOI22_X1   g09806(.A1(new_n9996_), .A2(\asqrt[38] ), .B1(new_n9994_), .B2(new_n9991_), .ZN(new_n9999_));
  INV_X1     g09807(.I(new_n9782_), .ZN(new_n10000_));
  OAI21_X1   g09808(.A1(new_n9999_), .A2(new_n4330_), .B(new_n10000_), .ZN(new_n10001_));
  NAND2_X1   g09809(.A1(new_n10001_), .A2(new_n9998_), .ZN(new_n10002_));
  OAI22_X1   g09810(.A1(new_n9999_), .A2(new_n4330_), .B1(new_n9997_), .B2(new_n9995_), .ZN(new_n10003_));
  AOI21_X1   g09811(.A1(new_n10003_), .A2(\asqrt[40] ), .B(new_n9789_), .ZN(new_n10004_));
  NOR2_X1    g09812(.A1(new_n10004_), .A2(new_n10002_), .ZN(new_n10005_));
  AOI22_X1   g09813(.A1(new_n10003_), .A2(\asqrt[40] ), .B1(new_n10001_), .B2(new_n9998_), .ZN(new_n10006_));
  INV_X1     g09814(.I(new_n9797_), .ZN(new_n10007_));
  OAI21_X1   g09815(.A1(new_n10006_), .A2(new_n3760_), .B(new_n10007_), .ZN(new_n10008_));
  NAND2_X1   g09816(.A1(new_n10008_), .A2(new_n10005_), .ZN(new_n10009_));
  OAI22_X1   g09817(.A1(new_n10006_), .A2(new_n3760_), .B1(new_n10004_), .B2(new_n10002_), .ZN(new_n10010_));
  AOI21_X1   g09818(.A1(new_n10010_), .A2(\asqrt[42] ), .B(new_n9804_), .ZN(new_n10011_));
  NOR2_X1    g09819(.A1(new_n10011_), .A2(new_n10009_), .ZN(new_n10012_));
  AOI22_X1   g09820(.A1(new_n10010_), .A2(\asqrt[42] ), .B1(new_n10008_), .B2(new_n10005_), .ZN(new_n10013_));
  INV_X1     g09821(.I(new_n9812_), .ZN(new_n10014_));
  OAI21_X1   g09822(.A1(new_n10013_), .A2(new_n3208_), .B(new_n10014_), .ZN(new_n10015_));
  NAND2_X1   g09823(.A1(new_n10015_), .A2(new_n10012_), .ZN(new_n10016_));
  OAI22_X1   g09824(.A1(new_n10013_), .A2(new_n3208_), .B1(new_n10011_), .B2(new_n10009_), .ZN(new_n10017_));
  AOI21_X1   g09825(.A1(new_n10017_), .A2(\asqrt[44] ), .B(new_n9819_), .ZN(new_n10018_));
  NOR2_X1    g09826(.A1(new_n10018_), .A2(new_n10016_), .ZN(new_n10019_));
  AOI22_X1   g09827(.A1(new_n10017_), .A2(\asqrt[44] ), .B1(new_n10015_), .B2(new_n10012_), .ZN(new_n10020_));
  INV_X1     g09828(.I(new_n9827_), .ZN(new_n10021_));
  OAI21_X1   g09829(.A1(new_n10020_), .A2(new_n2728_), .B(new_n10021_), .ZN(new_n10022_));
  NAND2_X1   g09830(.A1(new_n10022_), .A2(new_n10019_), .ZN(new_n10023_));
  OAI22_X1   g09831(.A1(new_n10020_), .A2(new_n2728_), .B1(new_n10018_), .B2(new_n10016_), .ZN(new_n10024_));
  AOI21_X1   g09832(.A1(new_n10024_), .A2(\asqrt[46] ), .B(new_n9834_), .ZN(new_n10025_));
  NOR2_X1    g09833(.A1(new_n10025_), .A2(new_n10023_), .ZN(new_n10026_));
  AOI22_X1   g09834(.A1(new_n10024_), .A2(\asqrt[46] ), .B1(new_n10022_), .B2(new_n10019_), .ZN(new_n10027_));
  INV_X1     g09835(.I(new_n9842_), .ZN(new_n10028_));
  OAI21_X1   g09836(.A1(new_n10027_), .A2(new_n2253_), .B(new_n10028_), .ZN(new_n10029_));
  NAND2_X1   g09837(.A1(new_n10029_), .A2(new_n10026_), .ZN(new_n10030_));
  OAI22_X1   g09838(.A1(new_n10027_), .A2(new_n2253_), .B1(new_n10025_), .B2(new_n10023_), .ZN(new_n10031_));
  AOI21_X1   g09839(.A1(new_n10031_), .A2(\asqrt[48] ), .B(new_n9849_), .ZN(new_n10032_));
  NOR2_X1    g09840(.A1(new_n10032_), .A2(new_n10030_), .ZN(new_n10033_));
  AOI22_X1   g09841(.A1(new_n10031_), .A2(\asqrt[48] ), .B1(new_n10029_), .B2(new_n10026_), .ZN(new_n10034_));
  INV_X1     g09842(.I(new_n9857_), .ZN(new_n10035_));
  OAI21_X1   g09843(.A1(new_n10034_), .A2(new_n1854_), .B(new_n10035_), .ZN(new_n10036_));
  NAND2_X1   g09844(.A1(new_n10036_), .A2(new_n10033_), .ZN(new_n10037_));
  OAI22_X1   g09845(.A1(new_n10034_), .A2(new_n1854_), .B1(new_n10032_), .B2(new_n10030_), .ZN(new_n10038_));
  AOI21_X1   g09846(.A1(new_n10038_), .A2(\asqrt[50] ), .B(new_n9864_), .ZN(new_n10039_));
  NOR2_X1    g09847(.A1(new_n10039_), .A2(new_n10037_), .ZN(new_n10040_));
  AOI22_X1   g09848(.A1(new_n10038_), .A2(\asqrt[50] ), .B1(new_n10036_), .B2(new_n10033_), .ZN(new_n10041_));
  INV_X1     g09849(.I(new_n9872_), .ZN(new_n10042_));
  OAI21_X1   g09850(.A1(new_n10041_), .A2(new_n1436_), .B(new_n10042_), .ZN(new_n10043_));
  NAND2_X1   g09851(.A1(new_n10043_), .A2(new_n10040_), .ZN(new_n10044_));
  OAI22_X1   g09852(.A1(new_n10041_), .A2(new_n1436_), .B1(new_n10039_), .B2(new_n10037_), .ZN(new_n10045_));
  AOI21_X1   g09853(.A1(new_n10045_), .A2(\asqrt[52] ), .B(new_n9879_), .ZN(new_n10046_));
  NOR2_X1    g09854(.A1(new_n10046_), .A2(new_n10044_), .ZN(new_n10047_));
  AOI22_X1   g09855(.A1(new_n10045_), .A2(\asqrt[52] ), .B1(new_n10043_), .B2(new_n10040_), .ZN(new_n10048_));
  INV_X1     g09856(.I(new_n9887_), .ZN(new_n10049_));
  OAI21_X1   g09857(.A1(new_n10048_), .A2(new_n1096_), .B(new_n10049_), .ZN(new_n10050_));
  NAND2_X1   g09858(.A1(new_n10050_), .A2(new_n10047_), .ZN(new_n10051_));
  OAI22_X1   g09859(.A1(new_n10048_), .A2(new_n1096_), .B1(new_n10046_), .B2(new_n10044_), .ZN(new_n10052_));
  AOI21_X1   g09860(.A1(new_n10052_), .A2(\asqrt[54] ), .B(new_n9893_), .ZN(new_n10053_));
  NOR2_X1    g09861(.A1(new_n10053_), .A2(new_n10051_), .ZN(new_n10054_));
  AOI22_X1   g09862(.A1(new_n10052_), .A2(\asqrt[54] ), .B1(new_n10050_), .B2(new_n10047_), .ZN(new_n10055_));
  INV_X1     g09863(.I(new_n9900_), .ZN(new_n10056_));
  OAI21_X1   g09864(.A1(new_n10055_), .A2(new_n825_), .B(new_n10056_), .ZN(new_n10057_));
  NAND2_X1   g09865(.A1(new_n10057_), .A2(new_n10054_), .ZN(new_n10058_));
  OAI22_X1   g09866(.A1(new_n10055_), .A2(new_n825_), .B1(new_n10053_), .B2(new_n10051_), .ZN(new_n10059_));
  AOI21_X1   g09867(.A1(new_n10059_), .A2(\asqrt[56] ), .B(new_n9906_), .ZN(new_n10060_));
  NOR2_X1    g09868(.A1(new_n10060_), .A2(new_n10058_), .ZN(new_n10061_));
  AOI22_X1   g09869(.A1(new_n10059_), .A2(\asqrt[56] ), .B1(new_n10057_), .B2(new_n10054_), .ZN(new_n10062_));
  INV_X1     g09870(.I(new_n9913_), .ZN(new_n10063_));
  OAI21_X1   g09871(.A1(new_n10062_), .A2(new_n587_), .B(new_n10063_), .ZN(new_n10064_));
  NAND2_X1   g09872(.A1(new_n10064_), .A2(new_n10061_), .ZN(new_n10065_));
  OAI22_X1   g09873(.A1(new_n10062_), .A2(new_n587_), .B1(new_n10060_), .B2(new_n10058_), .ZN(new_n10066_));
  AOI21_X1   g09874(.A1(new_n10066_), .A2(\asqrt[58] ), .B(new_n9919_), .ZN(new_n10067_));
  NOR2_X1    g09875(.A1(new_n10067_), .A2(new_n10065_), .ZN(new_n10068_));
  AOI22_X1   g09876(.A1(new_n10066_), .A2(\asqrt[58] ), .B1(new_n10064_), .B2(new_n10061_), .ZN(new_n10069_));
  INV_X1     g09877(.I(new_n9926_), .ZN(new_n10070_));
  OAI21_X1   g09878(.A1(new_n10069_), .A2(new_n376_), .B(new_n10070_), .ZN(new_n10071_));
  NAND2_X1   g09879(.A1(new_n10071_), .A2(new_n10068_), .ZN(new_n10072_));
  OAI22_X1   g09880(.A1(new_n10069_), .A2(new_n376_), .B1(new_n10067_), .B2(new_n10065_), .ZN(new_n10073_));
  AOI21_X1   g09881(.A1(new_n10073_), .A2(\asqrt[60] ), .B(new_n9932_), .ZN(new_n10074_));
  AOI22_X1   g09882(.A1(new_n10073_), .A2(\asqrt[60] ), .B1(new_n10071_), .B2(new_n10068_), .ZN(new_n10075_));
  OAI22_X1   g09883(.A1(new_n10075_), .A2(new_n229_), .B1(new_n10074_), .B2(new_n10072_), .ZN(new_n10076_));
  NOR4_X1    g09884(.A1(new_n10076_), .A2(\asqrt[62] ), .A3(new_n9639_), .A4(new_n9643_), .ZN(new_n10077_));
  NAND2_X1   g09885(.A1(new_n9659_), .A2(new_n9174_), .ZN(new_n10078_));
  XOR2_X1    g09886(.A1(new_n9659_), .A2(\asqrt[63] ), .Z(new_n10079_));
  AOI21_X1   g09887(.A1(\asqrt[25] ), .A2(new_n10078_), .B(new_n10079_), .ZN(new_n10080_));
  NAND2_X1   g09888(.A1(new_n10077_), .A2(new_n10080_), .ZN(new_n10081_));
  NOR4_X1    g09889(.A1(new_n10081_), .A2(new_n9620_), .A3(new_n9945_), .A4(new_n9627_), .ZN(new_n10082_));
  NOR2_X1    g09890(.A1(new_n9620_), .A2(\a[48] ), .ZN(new_n10083_));
  OAI21_X1   g09891(.A1(new_n10082_), .A2(new_n10083_), .B(new_n9619_), .ZN(new_n10084_));
  INV_X1     g09892(.I(new_n9619_), .ZN(new_n10085_));
  INV_X1     g09893(.I(new_n9627_), .ZN(new_n10086_));
  NOR2_X1    g09894(.A1(new_n10074_), .A2(new_n10072_), .ZN(new_n10087_));
  NOR3_X1    g09895(.A1(new_n10075_), .A2(new_n229_), .A3(new_n9938_), .ZN(new_n10088_));
  AOI21_X1   g09896(.A1(new_n10088_), .A2(new_n10087_), .B(new_n9644_), .ZN(new_n10089_));
  AOI21_X1   g09897(.A1(new_n10089_), .A2(new_n9943_), .B(new_n9639_), .ZN(new_n10090_));
  AOI22_X1   g09898(.A1(new_n9936_), .A2(\asqrt[61] ), .B1(new_n9934_), .B2(new_n9928_), .ZN(new_n10091_));
  NAND4_X1   g09899(.A1(new_n10091_), .A2(new_n196_), .A3(new_n9640_), .A4(new_n9937_), .ZN(new_n10092_));
  INV_X1     g09900(.I(new_n10080_), .ZN(new_n10093_));
  NOR2_X1    g09901(.A1(new_n10092_), .A2(new_n10093_), .ZN(new_n10094_));
  NAND4_X1   g09902(.A1(new_n10094_), .A2(new_n10090_), .A3(\a[49] ), .A4(new_n10086_), .ZN(new_n10095_));
  NAND3_X1   g09903(.A1(new_n10095_), .A2(\a[48] ), .A3(new_n10085_), .ZN(new_n10096_));
  NAND2_X1   g09904(.A1(new_n10084_), .A2(new_n10096_), .ZN(new_n10097_));
  NOR2_X1    g09905(.A1(new_n10081_), .A2(new_n9945_), .ZN(new_n10098_));
  NOR4_X1    g09906(.A1(new_n9625_), .A2(new_n9174_), .A3(new_n9674_), .A4(new_n9612_), .ZN(new_n10099_));
  NAND2_X1   g09907(.A1(\asqrt[25] ), .A2(\a[48] ), .ZN(new_n10100_));
  XOR2_X1    g09908(.A1(new_n10100_), .A2(new_n10099_), .Z(new_n10101_));
  NOR2_X1    g09909(.A1(new_n10101_), .A2(new_n9616_), .ZN(new_n10102_));
  INV_X1     g09910(.I(new_n10102_), .ZN(new_n10103_));
  NAND3_X1   g09911(.A1(new_n10094_), .A2(new_n10090_), .A3(new_n10086_), .ZN(new_n10104_));
  NAND2_X1   g09912(.A1(new_n9897_), .A2(\asqrt[55] ), .ZN(new_n10105_));
  AOI21_X1   g09913(.A1(new_n10105_), .A2(new_n9896_), .B(new_n724_), .ZN(new_n10106_));
  OAI21_X1   g09914(.A1(new_n9902_), .A2(new_n10106_), .B(\asqrt[57] ), .ZN(new_n10107_));
  AOI21_X1   g09915(.A1(new_n9909_), .A2(new_n10107_), .B(new_n504_), .ZN(new_n10108_));
  OAI21_X1   g09916(.A1(new_n9915_), .A2(new_n10108_), .B(\asqrt[59] ), .ZN(new_n10109_));
  AOI21_X1   g09917(.A1(new_n9922_), .A2(new_n10109_), .B(new_n275_), .ZN(new_n10110_));
  OAI21_X1   g09918(.A1(new_n9928_), .A2(new_n10110_), .B(\asqrt[61] ), .ZN(new_n10111_));
  NOR3_X1    g09919(.A1(new_n9935_), .A2(new_n10111_), .A3(new_n9938_), .ZN(new_n10112_));
  NOR3_X1    g09920(.A1(new_n10112_), .A2(new_n9644_), .A3(new_n9944_), .ZN(new_n10113_));
  OAI21_X1   g09921(.A1(new_n10113_), .A2(new_n9639_), .B(new_n10092_), .ZN(new_n10114_));
  NOR2_X1    g09922(.A1(new_n10086_), .A2(new_n10080_), .ZN(new_n10115_));
  NAND2_X1   g09923(.A1(new_n10115_), .A2(\asqrt[25] ), .ZN(new_n10116_));
  OAI21_X1   g09924(.A1(new_n10114_), .A2(new_n10116_), .B(new_n9646_), .ZN(new_n10117_));
  NAND3_X1   g09925(.A1(new_n10117_), .A2(new_n9647_), .A3(new_n10104_), .ZN(new_n10118_));
  NOR3_X1    g09926(.A1(new_n10081_), .A2(new_n9627_), .A3(new_n9945_), .ZN(\asqrt[24] ));
  NAND2_X1   g09927(.A1(new_n10052_), .A2(\asqrt[54] ), .ZN(new_n10120_));
  AOI21_X1   g09928(.A1(new_n10120_), .A2(new_n10051_), .B(new_n825_), .ZN(new_n10121_));
  OAI21_X1   g09929(.A1(new_n10054_), .A2(new_n10121_), .B(\asqrt[56] ), .ZN(new_n10122_));
  AOI21_X1   g09930(.A1(new_n10058_), .A2(new_n10122_), .B(new_n587_), .ZN(new_n10123_));
  OAI21_X1   g09931(.A1(new_n10061_), .A2(new_n10123_), .B(\asqrt[58] ), .ZN(new_n10124_));
  AOI21_X1   g09932(.A1(new_n10065_), .A2(new_n10124_), .B(new_n376_), .ZN(new_n10125_));
  OAI21_X1   g09933(.A1(new_n10068_), .A2(new_n10125_), .B(\asqrt[60] ), .ZN(new_n10126_));
  AOI21_X1   g09934(.A1(new_n10072_), .A2(new_n10126_), .B(new_n229_), .ZN(new_n10127_));
  NAND4_X1   g09935(.A1(new_n10127_), .A2(new_n9928_), .A3(new_n9934_), .A4(new_n9939_), .ZN(new_n10128_));
  NAND3_X1   g09936(.A1(new_n10128_), .A2(new_n9645_), .A3(new_n9943_), .ZN(new_n10129_));
  AOI21_X1   g09937(.A1(new_n9640_), .A2(new_n10129_), .B(new_n10077_), .ZN(new_n10130_));
  INV_X1     g09938(.I(new_n10116_), .ZN(new_n10131_));
  AOI21_X1   g09939(.A1(new_n10130_), .A2(new_n10131_), .B(\a[50] ), .ZN(new_n10132_));
  OAI21_X1   g09940(.A1(new_n10132_), .A2(new_n9648_), .B(\asqrt[24] ), .ZN(new_n10133_));
  NAND4_X1   g09941(.A1(new_n10133_), .A2(new_n10118_), .A3(new_n9212_), .A4(new_n10103_), .ZN(new_n10134_));
  NAND2_X1   g09942(.A1(new_n10134_), .A2(new_n10097_), .ZN(new_n10135_));
  NAND3_X1   g09943(.A1(new_n10084_), .A2(new_n10096_), .A3(new_n10103_), .ZN(new_n10136_));
  AOI21_X1   g09944(.A1(\asqrt[25] ), .A2(new_n9646_), .B(\a[51] ), .ZN(new_n10137_));
  NOR2_X1    g09945(.A1(new_n9663_), .A2(\a[50] ), .ZN(new_n10138_));
  AOI21_X1   g09946(.A1(\asqrt[25] ), .A2(\a[50] ), .B(new_n9650_), .ZN(new_n10139_));
  OAI21_X1   g09947(.A1(new_n10138_), .A2(new_n10137_), .B(new_n10139_), .ZN(new_n10140_));
  INV_X1     g09948(.I(new_n10140_), .ZN(new_n10141_));
  NAND3_X1   g09949(.A1(\asqrt[24] ), .A2(new_n9671_), .A3(new_n10141_), .ZN(new_n10142_));
  OAI21_X1   g09950(.A1(new_n10104_), .A2(new_n10140_), .B(new_n9670_), .ZN(new_n10143_));
  NAND3_X1   g09951(.A1(new_n10142_), .A2(new_n10143_), .A3(new_n8763_), .ZN(new_n10144_));
  AOI21_X1   g09952(.A1(new_n10136_), .A2(\asqrt[26] ), .B(new_n10144_), .ZN(new_n10145_));
  NOR2_X1    g09953(.A1(new_n10135_), .A2(new_n10145_), .ZN(new_n10146_));
  NAND2_X1   g09954(.A1(new_n10136_), .A2(\asqrt[26] ), .ZN(new_n10147_));
  AOI21_X1   g09955(.A1(new_n10135_), .A2(new_n10147_), .B(new_n8763_), .ZN(new_n10148_));
  NAND2_X1   g09956(.A1(new_n9685_), .A2(\asqrt[27] ), .ZN(new_n10149_));
  INV_X1     g09957(.I(new_n10149_), .ZN(new_n10150_));
  NAND2_X1   g09958(.A1(new_n9679_), .A2(new_n9682_), .ZN(new_n10151_));
  NAND3_X1   g09959(.A1(new_n10151_), .A2(new_n9954_), .A3(new_n8763_), .ZN(new_n10152_));
  NOR3_X1    g09960(.A1(new_n10104_), .A2(new_n10150_), .A3(new_n10152_), .ZN(new_n10153_));
  NOR2_X1    g09961(.A1(new_n10104_), .A2(new_n10152_), .ZN(new_n10154_));
  NOR2_X1    g09962(.A1(new_n10154_), .A2(new_n10149_), .ZN(new_n10155_));
  NOR3_X1    g09963(.A1(new_n10155_), .A2(\asqrt[28] ), .A3(new_n10153_), .ZN(new_n10156_));
  INV_X1     g09964(.I(new_n10156_), .ZN(new_n10157_));
  OAI21_X1   g09965(.A1(new_n10148_), .A2(new_n10157_), .B(new_n10146_), .ZN(new_n10158_));
  OAI21_X1   g09966(.A1(new_n10148_), .A2(new_n10146_), .B(\asqrt[28] ), .ZN(new_n10159_));
  NOR2_X1    g09967(.A1(new_n9956_), .A2(new_n9955_), .ZN(new_n10160_));
  NOR4_X1    g09968(.A1(new_n10104_), .A2(\asqrt[28] ), .A3(new_n10160_), .A4(new_n9960_), .ZN(new_n10161_));
  AOI21_X1   g09969(.A1(new_n9684_), .A2(new_n10149_), .B(new_n8319_), .ZN(new_n10162_));
  NOR2_X1    g09970(.A1(new_n10161_), .A2(new_n10162_), .ZN(new_n10163_));
  NAND2_X1   g09971(.A1(new_n10163_), .A2(new_n7931_), .ZN(new_n10164_));
  INV_X1     g09972(.I(new_n10164_), .ZN(new_n10165_));
  AOI21_X1   g09973(.A1(new_n10159_), .A2(new_n10165_), .B(new_n10158_), .ZN(new_n10166_));
  AOI21_X1   g09974(.A1(new_n10158_), .A2(new_n10159_), .B(new_n7931_), .ZN(new_n10167_));
  NAND2_X1   g09975(.A1(new_n9707_), .A2(\asqrt[29] ), .ZN(new_n10168_));
  NOR2_X1    g09976(.A1(new_n9702_), .A2(new_n9703_), .ZN(new_n10169_));
  NOR4_X1    g09977(.A1(new_n10104_), .A2(\asqrt[29] ), .A3(new_n10169_), .A4(new_n9707_), .ZN(new_n10170_));
  XOR2_X1    g09978(.A1(new_n10170_), .A2(new_n10168_), .Z(new_n10171_));
  NAND2_X1   g09979(.A1(new_n10171_), .A2(new_n7517_), .ZN(new_n10172_));
  OAI21_X1   g09980(.A1(new_n10167_), .A2(new_n10172_), .B(new_n10166_), .ZN(new_n10173_));
  OAI21_X1   g09981(.A1(new_n10166_), .A2(new_n10167_), .B(\asqrt[30] ), .ZN(new_n10174_));
  NOR4_X1    g09982(.A1(new_n10104_), .A2(\asqrt[30] ), .A3(new_n9710_), .A4(new_n9968_), .ZN(new_n10175_));
  AOI21_X1   g09983(.A1(new_n10168_), .A2(new_n9706_), .B(new_n7517_), .ZN(new_n10176_));
  NOR2_X1    g09984(.A1(new_n10175_), .A2(new_n10176_), .ZN(new_n10177_));
  NAND2_X1   g09985(.A1(new_n10177_), .A2(new_n7110_), .ZN(new_n10178_));
  INV_X1     g09986(.I(new_n10178_), .ZN(new_n10179_));
  AOI21_X1   g09987(.A1(new_n10174_), .A2(new_n10179_), .B(new_n10173_), .ZN(new_n10180_));
  AOI22_X1   g09988(.A1(new_n10134_), .A2(new_n10097_), .B1(\asqrt[26] ), .B2(new_n10136_), .ZN(new_n10181_));
  OAI21_X1   g09989(.A1(new_n10181_), .A2(new_n8763_), .B(new_n10156_), .ZN(new_n10182_));
  OAI22_X1   g09990(.A1(new_n10181_), .A2(new_n8763_), .B1(new_n10135_), .B2(new_n10145_), .ZN(new_n10183_));
  AOI22_X1   g09991(.A1(new_n10183_), .A2(\asqrt[28] ), .B1(new_n10182_), .B2(new_n10146_), .ZN(new_n10184_));
  INV_X1     g09992(.I(new_n10172_), .ZN(new_n10185_));
  OAI21_X1   g09993(.A1(new_n10184_), .A2(new_n7931_), .B(new_n10185_), .ZN(new_n10186_));
  AOI21_X1   g09994(.A1(new_n10183_), .A2(\asqrt[28] ), .B(new_n10164_), .ZN(new_n10187_));
  OAI22_X1   g09995(.A1(new_n10184_), .A2(new_n7931_), .B1(new_n10187_), .B2(new_n10158_), .ZN(new_n10188_));
  AOI22_X1   g09996(.A1(new_n10188_), .A2(\asqrt[30] ), .B1(new_n10186_), .B2(new_n10166_), .ZN(new_n10189_));
  NAND2_X1   g09997(.A1(new_n9721_), .A2(\asqrt[31] ), .ZN(new_n10190_));
  NOR4_X1    g09998(.A1(new_n10104_), .A2(\asqrt[31] ), .A3(new_n9716_), .A4(new_n9721_), .ZN(new_n10191_));
  XOR2_X1    g09999(.A1(new_n10191_), .A2(new_n10190_), .Z(new_n10192_));
  NAND2_X1   g10000(.A1(new_n10192_), .A2(new_n6708_), .ZN(new_n10193_));
  INV_X1     g10001(.I(new_n10193_), .ZN(new_n10194_));
  OAI21_X1   g10002(.A1(new_n10189_), .A2(new_n7110_), .B(new_n10194_), .ZN(new_n10195_));
  NAND2_X1   g10003(.A1(new_n10195_), .A2(new_n10180_), .ZN(new_n10196_));
  AOI21_X1   g10004(.A1(new_n10188_), .A2(\asqrt[30] ), .B(new_n10178_), .ZN(new_n10197_));
  OAI22_X1   g10005(.A1(new_n10189_), .A2(new_n7110_), .B1(new_n10197_), .B2(new_n10173_), .ZN(new_n10198_));
  NOR4_X1    g10006(.A1(new_n10104_), .A2(\asqrt[32] ), .A3(new_n9724_), .A4(new_n9975_), .ZN(new_n10199_));
  AOI21_X1   g10007(.A1(new_n10190_), .A2(new_n9720_), .B(new_n6708_), .ZN(new_n10200_));
  NOR2_X1    g10008(.A1(new_n10199_), .A2(new_n10200_), .ZN(new_n10201_));
  NAND2_X1   g10009(.A1(new_n10201_), .A2(new_n6365_), .ZN(new_n10202_));
  AOI21_X1   g10010(.A1(new_n10198_), .A2(\asqrt[32] ), .B(new_n10202_), .ZN(new_n10203_));
  NOR2_X1    g10011(.A1(new_n10203_), .A2(new_n10196_), .ZN(new_n10204_));
  AOI22_X1   g10012(.A1(new_n10198_), .A2(\asqrt[32] ), .B1(new_n10195_), .B2(new_n10180_), .ZN(new_n10205_));
  NAND2_X1   g10013(.A1(new_n9735_), .A2(\asqrt[33] ), .ZN(new_n10206_));
  NOR4_X1    g10014(.A1(new_n10104_), .A2(\asqrt[33] ), .A3(new_n9730_), .A4(new_n9735_), .ZN(new_n10207_));
  XOR2_X1    g10015(.A1(new_n10207_), .A2(new_n10206_), .Z(new_n10208_));
  NAND2_X1   g10016(.A1(new_n10208_), .A2(new_n5991_), .ZN(new_n10209_));
  INV_X1     g10017(.I(new_n10209_), .ZN(new_n10210_));
  OAI21_X1   g10018(.A1(new_n10205_), .A2(new_n6365_), .B(new_n10210_), .ZN(new_n10211_));
  NAND2_X1   g10019(.A1(new_n10211_), .A2(new_n10204_), .ZN(new_n10212_));
  OAI22_X1   g10020(.A1(new_n10205_), .A2(new_n6365_), .B1(new_n10203_), .B2(new_n10196_), .ZN(new_n10213_));
  NOR4_X1    g10021(.A1(new_n10104_), .A2(\asqrt[34] ), .A3(new_n9737_), .A4(new_n9982_), .ZN(new_n10214_));
  AOI21_X1   g10022(.A1(new_n10206_), .A2(new_n9734_), .B(new_n5991_), .ZN(new_n10215_));
  NOR2_X1    g10023(.A1(new_n10214_), .A2(new_n10215_), .ZN(new_n10216_));
  NAND2_X1   g10024(.A1(new_n10216_), .A2(new_n5626_), .ZN(new_n10217_));
  AOI21_X1   g10025(.A1(new_n10213_), .A2(\asqrt[34] ), .B(new_n10217_), .ZN(new_n10218_));
  NOR2_X1    g10026(.A1(new_n10218_), .A2(new_n10212_), .ZN(new_n10219_));
  AOI22_X1   g10027(.A1(new_n10213_), .A2(\asqrt[34] ), .B1(new_n10211_), .B2(new_n10204_), .ZN(new_n10220_));
  NAND2_X1   g10028(.A1(new_n9748_), .A2(\asqrt[35] ), .ZN(new_n10221_));
  NOR4_X1    g10029(.A1(new_n10104_), .A2(\asqrt[35] ), .A3(new_n9743_), .A4(new_n9748_), .ZN(new_n10222_));
  XOR2_X1    g10030(.A1(new_n10222_), .A2(new_n10221_), .Z(new_n10223_));
  NAND2_X1   g10031(.A1(new_n10223_), .A2(new_n5273_), .ZN(new_n10224_));
  INV_X1     g10032(.I(new_n10224_), .ZN(new_n10225_));
  OAI21_X1   g10033(.A1(new_n10220_), .A2(new_n5626_), .B(new_n10225_), .ZN(new_n10226_));
  NAND2_X1   g10034(.A1(new_n10226_), .A2(new_n10219_), .ZN(new_n10227_));
  OAI22_X1   g10035(.A1(new_n10220_), .A2(new_n5626_), .B1(new_n10218_), .B2(new_n10212_), .ZN(new_n10228_));
  NAND2_X1   g10036(.A1(new_n9989_), .A2(\asqrt[36] ), .ZN(new_n10229_));
  NOR4_X1    g10037(.A1(new_n10104_), .A2(\asqrt[36] ), .A3(new_n9751_), .A4(new_n9989_), .ZN(new_n10230_));
  XOR2_X1    g10038(.A1(new_n10230_), .A2(new_n10229_), .Z(new_n10231_));
  NAND2_X1   g10039(.A1(new_n10231_), .A2(new_n4973_), .ZN(new_n10232_));
  AOI21_X1   g10040(.A1(new_n10228_), .A2(\asqrt[36] ), .B(new_n10232_), .ZN(new_n10233_));
  NOR2_X1    g10041(.A1(new_n10233_), .A2(new_n10227_), .ZN(new_n10234_));
  AOI22_X1   g10042(.A1(new_n10228_), .A2(\asqrt[36] ), .B1(new_n10226_), .B2(new_n10219_), .ZN(new_n10235_));
  NOR4_X1    g10043(.A1(new_n10104_), .A2(\asqrt[37] ), .A3(new_n9758_), .A4(new_n9763_), .ZN(new_n10236_));
  AOI21_X1   g10044(.A1(new_n10229_), .A2(new_n9988_), .B(new_n4973_), .ZN(new_n10237_));
  NOR2_X1    g10045(.A1(new_n10236_), .A2(new_n10237_), .ZN(new_n10238_));
  NAND2_X1   g10046(.A1(new_n10238_), .A2(new_n4645_), .ZN(new_n10239_));
  INV_X1     g10047(.I(new_n10239_), .ZN(new_n10240_));
  OAI21_X1   g10048(.A1(new_n10235_), .A2(new_n4973_), .B(new_n10240_), .ZN(new_n10241_));
  NAND2_X1   g10049(.A1(new_n10241_), .A2(new_n10234_), .ZN(new_n10242_));
  OAI22_X1   g10050(.A1(new_n10235_), .A2(new_n4973_), .B1(new_n10233_), .B2(new_n10227_), .ZN(new_n10243_));
  NAND2_X1   g10051(.A1(new_n9996_), .A2(\asqrt[38] ), .ZN(new_n10244_));
  NOR4_X1    g10052(.A1(new_n10104_), .A2(\asqrt[38] ), .A3(new_n9766_), .A4(new_n9996_), .ZN(new_n10245_));
  XOR2_X1    g10053(.A1(new_n10245_), .A2(new_n10244_), .Z(new_n10246_));
  NAND2_X1   g10054(.A1(new_n10246_), .A2(new_n4330_), .ZN(new_n10247_));
  AOI21_X1   g10055(.A1(new_n10243_), .A2(\asqrt[38] ), .B(new_n10247_), .ZN(new_n10248_));
  NOR2_X1    g10056(.A1(new_n10248_), .A2(new_n10242_), .ZN(new_n10249_));
  AOI22_X1   g10057(.A1(new_n10243_), .A2(\asqrt[38] ), .B1(new_n10241_), .B2(new_n10234_), .ZN(new_n10250_));
  NOR4_X1    g10058(.A1(new_n10104_), .A2(\asqrt[39] ), .A3(new_n9773_), .A4(new_n9778_), .ZN(new_n10251_));
  AOI21_X1   g10059(.A1(new_n10244_), .A2(new_n9995_), .B(new_n4330_), .ZN(new_n10252_));
  NOR2_X1    g10060(.A1(new_n10251_), .A2(new_n10252_), .ZN(new_n10253_));
  NAND2_X1   g10061(.A1(new_n10253_), .A2(new_n4018_), .ZN(new_n10254_));
  INV_X1     g10062(.I(new_n10254_), .ZN(new_n10255_));
  OAI21_X1   g10063(.A1(new_n10250_), .A2(new_n4330_), .B(new_n10255_), .ZN(new_n10256_));
  NAND2_X1   g10064(.A1(new_n10256_), .A2(new_n10249_), .ZN(new_n10257_));
  OAI22_X1   g10065(.A1(new_n10250_), .A2(new_n4330_), .B1(new_n10248_), .B2(new_n10242_), .ZN(new_n10258_));
  NAND2_X1   g10066(.A1(new_n10003_), .A2(\asqrt[40] ), .ZN(new_n10259_));
  NOR4_X1    g10067(.A1(new_n10104_), .A2(\asqrt[40] ), .A3(new_n9781_), .A4(new_n10003_), .ZN(new_n10260_));
  XOR2_X1    g10068(.A1(new_n10260_), .A2(new_n10259_), .Z(new_n10261_));
  NAND2_X1   g10069(.A1(new_n10261_), .A2(new_n3760_), .ZN(new_n10262_));
  AOI21_X1   g10070(.A1(new_n10258_), .A2(\asqrt[40] ), .B(new_n10262_), .ZN(new_n10263_));
  NOR2_X1    g10071(.A1(new_n10263_), .A2(new_n10257_), .ZN(new_n10264_));
  AOI22_X1   g10072(.A1(new_n10258_), .A2(\asqrt[40] ), .B1(new_n10256_), .B2(new_n10249_), .ZN(new_n10265_));
  NOR4_X1    g10073(.A1(new_n10104_), .A2(\asqrt[41] ), .A3(new_n9788_), .A4(new_n9793_), .ZN(new_n10266_));
  AOI21_X1   g10074(.A1(new_n10259_), .A2(new_n10002_), .B(new_n3760_), .ZN(new_n10267_));
  NOR2_X1    g10075(.A1(new_n10266_), .A2(new_n10267_), .ZN(new_n10268_));
  NAND2_X1   g10076(.A1(new_n10268_), .A2(new_n3481_), .ZN(new_n10269_));
  INV_X1     g10077(.I(new_n10269_), .ZN(new_n10270_));
  OAI21_X1   g10078(.A1(new_n10265_), .A2(new_n3760_), .B(new_n10270_), .ZN(new_n10271_));
  NAND2_X1   g10079(.A1(new_n10271_), .A2(new_n10264_), .ZN(new_n10272_));
  OAI22_X1   g10080(.A1(new_n10265_), .A2(new_n3760_), .B1(new_n10263_), .B2(new_n10257_), .ZN(new_n10273_));
  NAND2_X1   g10081(.A1(new_n10010_), .A2(\asqrt[42] ), .ZN(new_n10274_));
  NOR4_X1    g10082(.A1(new_n10104_), .A2(\asqrt[42] ), .A3(new_n9796_), .A4(new_n10010_), .ZN(new_n10275_));
  XOR2_X1    g10083(.A1(new_n10275_), .A2(new_n10274_), .Z(new_n10276_));
  NAND2_X1   g10084(.A1(new_n10276_), .A2(new_n3208_), .ZN(new_n10277_));
  AOI21_X1   g10085(.A1(new_n10273_), .A2(\asqrt[42] ), .B(new_n10277_), .ZN(new_n10278_));
  NOR2_X1    g10086(.A1(new_n10278_), .A2(new_n10272_), .ZN(new_n10279_));
  AOI22_X1   g10087(.A1(new_n10273_), .A2(\asqrt[42] ), .B1(new_n10271_), .B2(new_n10264_), .ZN(new_n10280_));
  NOR4_X1    g10088(.A1(new_n10104_), .A2(\asqrt[43] ), .A3(new_n9803_), .A4(new_n9808_), .ZN(new_n10281_));
  AOI21_X1   g10089(.A1(new_n10274_), .A2(new_n10009_), .B(new_n3208_), .ZN(new_n10282_));
  NOR2_X1    g10090(.A1(new_n10281_), .A2(new_n10282_), .ZN(new_n10283_));
  NAND2_X1   g10091(.A1(new_n10283_), .A2(new_n2941_), .ZN(new_n10284_));
  INV_X1     g10092(.I(new_n10284_), .ZN(new_n10285_));
  OAI21_X1   g10093(.A1(new_n10280_), .A2(new_n3208_), .B(new_n10285_), .ZN(new_n10286_));
  NAND2_X1   g10094(.A1(new_n10286_), .A2(new_n10279_), .ZN(new_n10287_));
  OAI22_X1   g10095(.A1(new_n10280_), .A2(new_n3208_), .B1(new_n10278_), .B2(new_n10272_), .ZN(new_n10288_));
  NAND2_X1   g10096(.A1(new_n10017_), .A2(\asqrt[44] ), .ZN(new_n10289_));
  NOR4_X1    g10097(.A1(new_n10104_), .A2(\asqrt[44] ), .A3(new_n9811_), .A4(new_n10017_), .ZN(new_n10290_));
  XOR2_X1    g10098(.A1(new_n10290_), .A2(new_n10289_), .Z(new_n10291_));
  NAND2_X1   g10099(.A1(new_n10291_), .A2(new_n2728_), .ZN(new_n10292_));
  AOI21_X1   g10100(.A1(new_n10288_), .A2(\asqrt[44] ), .B(new_n10292_), .ZN(new_n10293_));
  NOR2_X1    g10101(.A1(new_n10293_), .A2(new_n10287_), .ZN(new_n10294_));
  AOI22_X1   g10102(.A1(new_n10288_), .A2(\asqrt[44] ), .B1(new_n10286_), .B2(new_n10279_), .ZN(new_n10295_));
  NAND2_X1   g10103(.A1(new_n9823_), .A2(\asqrt[45] ), .ZN(new_n10296_));
  NOR4_X1    g10104(.A1(new_n10104_), .A2(\asqrt[45] ), .A3(new_n9818_), .A4(new_n9823_), .ZN(new_n10297_));
  XOR2_X1    g10105(.A1(new_n10297_), .A2(new_n10296_), .Z(new_n10298_));
  NAND2_X1   g10106(.A1(new_n10298_), .A2(new_n2488_), .ZN(new_n10299_));
  INV_X1     g10107(.I(new_n10299_), .ZN(new_n10300_));
  OAI21_X1   g10108(.A1(new_n10295_), .A2(new_n2728_), .B(new_n10300_), .ZN(new_n10301_));
  NAND2_X1   g10109(.A1(new_n10301_), .A2(new_n10294_), .ZN(new_n10302_));
  OAI22_X1   g10110(.A1(new_n10295_), .A2(new_n2728_), .B1(new_n10293_), .B2(new_n10287_), .ZN(new_n10303_));
  NOR4_X1    g10111(.A1(new_n10104_), .A2(\asqrt[46] ), .A3(new_n9826_), .A4(new_n10024_), .ZN(new_n10304_));
  AOI21_X1   g10112(.A1(new_n10296_), .A2(new_n9822_), .B(new_n2488_), .ZN(new_n10305_));
  NOR2_X1    g10113(.A1(new_n10304_), .A2(new_n10305_), .ZN(new_n10306_));
  NAND2_X1   g10114(.A1(new_n10306_), .A2(new_n2253_), .ZN(new_n10307_));
  AOI21_X1   g10115(.A1(new_n10303_), .A2(\asqrt[46] ), .B(new_n10307_), .ZN(new_n10308_));
  NOR2_X1    g10116(.A1(new_n10308_), .A2(new_n10302_), .ZN(new_n10309_));
  AOI22_X1   g10117(.A1(new_n10303_), .A2(\asqrt[46] ), .B1(new_n10301_), .B2(new_n10294_), .ZN(new_n10310_));
  NAND2_X1   g10118(.A1(new_n9838_), .A2(\asqrt[47] ), .ZN(new_n10311_));
  NOR4_X1    g10119(.A1(new_n10104_), .A2(\asqrt[47] ), .A3(new_n9833_), .A4(new_n9838_), .ZN(new_n10312_));
  XOR2_X1    g10120(.A1(new_n10312_), .A2(new_n10311_), .Z(new_n10313_));
  NAND2_X1   g10121(.A1(new_n10313_), .A2(new_n2046_), .ZN(new_n10314_));
  INV_X1     g10122(.I(new_n10314_), .ZN(new_n10315_));
  OAI21_X1   g10123(.A1(new_n10310_), .A2(new_n2253_), .B(new_n10315_), .ZN(new_n10316_));
  NAND2_X1   g10124(.A1(new_n10316_), .A2(new_n10309_), .ZN(new_n10317_));
  OAI22_X1   g10125(.A1(new_n10310_), .A2(new_n2253_), .B1(new_n10308_), .B2(new_n10302_), .ZN(new_n10318_));
  NOR4_X1    g10126(.A1(new_n10104_), .A2(\asqrt[48] ), .A3(new_n9841_), .A4(new_n10031_), .ZN(new_n10319_));
  AOI21_X1   g10127(.A1(new_n10311_), .A2(new_n9837_), .B(new_n2046_), .ZN(new_n10320_));
  NOR2_X1    g10128(.A1(new_n10319_), .A2(new_n10320_), .ZN(new_n10321_));
  NAND2_X1   g10129(.A1(new_n10321_), .A2(new_n1854_), .ZN(new_n10322_));
  AOI21_X1   g10130(.A1(new_n10318_), .A2(\asqrt[48] ), .B(new_n10322_), .ZN(new_n10323_));
  NOR2_X1    g10131(.A1(new_n10323_), .A2(new_n10317_), .ZN(new_n10324_));
  AOI22_X1   g10132(.A1(new_n10318_), .A2(\asqrt[48] ), .B1(new_n10316_), .B2(new_n10309_), .ZN(new_n10325_));
  NAND2_X1   g10133(.A1(new_n9853_), .A2(\asqrt[49] ), .ZN(new_n10326_));
  NOR4_X1    g10134(.A1(new_n10104_), .A2(\asqrt[49] ), .A3(new_n9848_), .A4(new_n9853_), .ZN(new_n10327_));
  XOR2_X1    g10135(.A1(new_n10327_), .A2(new_n10326_), .Z(new_n10328_));
  NAND2_X1   g10136(.A1(new_n10328_), .A2(new_n1595_), .ZN(new_n10329_));
  INV_X1     g10137(.I(new_n10329_), .ZN(new_n10330_));
  OAI21_X1   g10138(.A1(new_n10325_), .A2(new_n1854_), .B(new_n10330_), .ZN(new_n10331_));
  NAND2_X1   g10139(.A1(new_n10331_), .A2(new_n10324_), .ZN(new_n10332_));
  OAI22_X1   g10140(.A1(new_n10325_), .A2(new_n1854_), .B1(new_n10323_), .B2(new_n10317_), .ZN(new_n10333_));
  NOR4_X1    g10141(.A1(new_n10104_), .A2(\asqrt[50] ), .A3(new_n9856_), .A4(new_n10038_), .ZN(new_n10334_));
  AOI21_X1   g10142(.A1(new_n10326_), .A2(new_n9852_), .B(new_n1595_), .ZN(new_n10335_));
  NOR2_X1    g10143(.A1(new_n10334_), .A2(new_n10335_), .ZN(new_n10336_));
  NAND2_X1   g10144(.A1(new_n10336_), .A2(new_n1436_), .ZN(new_n10337_));
  AOI21_X1   g10145(.A1(new_n10333_), .A2(\asqrt[50] ), .B(new_n10337_), .ZN(new_n10338_));
  NOR2_X1    g10146(.A1(new_n10338_), .A2(new_n10332_), .ZN(new_n10339_));
  AOI22_X1   g10147(.A1(new_n10333_), .A2(\asqrt[50] ), .B1(new_n10331_), .B2(new_n10324_), .ZN(new_n10340_));
  NAND2_X1   g10148(.A1(new_n9868_), .A2(\asqrt[51] ), .ZN(new_n10341_));
  NOR4_X1    g10149(.A1(new_n10104_), .A2(\asqrt[51] ), .A3(new_n9863_), .A4(new_n9868_), .ZN(new_n10342_));
  XOR2_X1    g10150(.A1(new_n10342_), .A2(new_n10341_), .Z(new_n10343_));
  NAND2_X1   g10151(.A1(new_n10343_), .A2(new_n1260_), .ZN(new_n10344_));
  INV_X1     g10152(.I(new_n10344_), .ZN(new_n10345_));
  OAI21_X1   g10153(.A1(new_n10340_), .A2(new_n1436_), .B(new_n10345_), .ZN(new_n10346_));
  NAND2_X1   g10154(.A1(new_n10346_), .A2(new_n10339_), .ZN(new_n10347_));
  OAI22_X1   g10155(.A1(new_n10340_), .A2(new_n1436_), .B1(new_n10338_), .B2(new_n10332_), .ZN(new_n10348_));
  NAND2_X1   g10156(.A1(new_n10045_), .A2(\asqrt[52] ), .ZN(new_n10349_));
  NOR4_X1    g10157(.A1(new_n10104_), .A2(\asqrt[52] ), .A3(new_n9871_), .A4(new_n10045_), .ZN(new_n10350_));
  XOR2_X1    g10158(.A1(new_n10350_), .A2(new_n10349_), .Z(new_n10351_));
  NAND2_X1   g10159(.A1(new_n10351_), .A2(new_n1096_), .ZN(new_n10352_));
  AOI21_X1   g10160(.A1(new_n10348_), .A2(\asqrt[52] ), .B(new_n10352_), .ZN(new_n10353_));
  NOR2_X1    g10161(.A1(new_n10353_), .A2(new_n10347_), .ZN(new_n10354_));
  AOI22_X1   g10162(.A1(new_n10348_), .A2(\asqrt[52] ), .B1(new_n10346_), .B2(new_n10339_), .ZN(new_n10355_));
  NOR4_X1    g10163(.A1(new_n10104_), .A2(\asqrt[53] ), .A3(new_n9878_), .A4(new_n9883_), .ZN(new_n10356_));
  AOI21_X1   g10164(.A1(new_n10349_), .A2(new_n10044_), .B(new_n1096_), .ZN(new_n10357_));
  NOR2_X1    g10165(.A1(new_n10356_), .A2(new_n10357_), .ZN(new_n10358_));
  NAND2_X1   g10166(.A1(new_n10358_), .A2(new_n970_), .ZN(new_n10359_));
  INV_X1     g10167(.I(new_n10359_), .ZN(new_n10360_));
  OAI21_X1   g10168(.A1(new_n10355_), .A2(new_n1096_), .B(new_n10360_), .ZN(new_n10361_));
  NAND2_X1   g10169(.A1(new_n10361_), .A2(new_n10354_), .ZN(new_n10362_));
  OAI22_X1   g10170(.A1(new_n10355_), .A2(new_n1096_), .B1(new_n10353_), .B2(new_n10347_), .ZN(new_n10363_));
  NOR4_X1    g10171(.A1(new_n10104_), .A2(\asqrt[54] ), .A3(new_n9886_), .A4(new_n10052_), .ZN(new_n10364_));
  XOR2_X1    g10172(.A1(new_n10364_), .A2(new_n10120_), .Z(new_n10365_));
  NAND2_X1   g10173(.A1(new_n10365_), .A2(new_n825_), .ZN(new_n10366_));
  AOI21_X1   g10174(.A1(new_n10363_), .A2(\asqrt[54] ), .B(new_n10366_), .ZN(new_n10367_));
  NOR2_X1    g10175(.A1(new_n10367_), .A2(new_n10362_), .ZN(new_n10368_));
  AOI22_X1   g10176(.A1(new_n10363_), .A2(\asqrt[54] ), .B1(new_n10361_), .B2(new_n10354_), .ZN(new_n10369_));
  NOR4_X1    g10177(.A1(new_n10104_), .A2(\asqrt[55] ), .A3(new_n9892_), .A4(new_n9897_), .ZN(new_n10370_));
  XOR2_X1    g10178(.A1(new_n10370_), .A2(new_n10105_), .Z(new_n10371_));
  NAND2_X1   g10179(.A1(new_n10371_), .A2(new_n724_), .ZN(new_n10372_));
  INV_X1     g10180(.I(new_n10372_), .ZN(new_n10373_));
  OAI21_X1   g10181(.A1(new_n10369_), .A2(new_n825_), .B(new_n10373_), .ZN(new_n10374_));
  NAND2_X1   g10182(.A1(new_n10374_), .A2(new_n10368_), .ZN(new_n10375_));
  OAI22_X1   g10183(.A1(new_n10369_), .A2(new_n825_), .B1(new_n10367_), .B2(new_n10362_), .ZN(new_n10376_));
  NOR4_X1    g10184(.A1(new_n10104_), .A2(\asqrt[56] ), .A3(new_n9899_), .A4(new_n10059_), .ZN(new_n10377_));
  XOR2_X1    g10185(.A1(new_n10377_), .A2(new_n10122_), .Z(new_n10378_));
  NAND2_X1   g10186(.A1(new_n10378_), .A2(new_n587_), .ZN(new_n10379_));
  AOI21_X1   g10187(.A1(new_n10376_), .A2(\asqrt[56] ), .B(new_n10379_), .ZN(new_n10380_));
  NOR2_X1    g10188(.A1(new_n10380_), .A2(new_n10375_), .ZN(new_n10381_));
  AOI22_X1   g10189(.A1(new_n10376_), .A2(\asqrt[56] ), .B1(new_n10374_), .B2(new_n10368_), .ZN(new_n10382_));
  NOR4_X1    g10190(.A1(new_n10104_), .A2(\asqrt[57] ), .A3(new_n9905_), .A4(new_n9910_), .ZN(new_n10383_));
  XOR2_X1    g10191(.A1(new_n10383_), .A2(new_n10107_), .Z(new_n10384_));
  NAND2_X1   g10192(.A1(new_n10384_), .A2(new_n504_), .ZN(new_n10385_));
  INV_X1     g10193(.I(new_n10385_), .ZN(new_n10386_));
  OAI21_X1   g10194(.A1(new_n10382_), .A2(new_n587_), .B(new_n10386_), .ZN(new_n10387_));
  NAND2_X1   g10195(.A1(new_n10387_), .A2(new_n10381_), .ZN(new_n10388_));
  OAI22_X1   g10196(.A1(new_n10382_), .A2(new_n587_), .B1(new_n10380_), .B2(new_n10375_), .ZN(new_n10389_));
  NOR4_X1    g10197(.A1(new_n10104_), .A2(\asqrt[58] ), .A3(new_n9912_), .A4(new_n10066_), .ZN(new_n10390_));
  XOR2_X1    g10198(.A1(new_n10390_), .A2(new_n10124_), .Z(new_n10391_));
  NAND2_X1   g10199(.A1(new_n10391_), .A2(new_n376_), .ZN(new_n10392_));
  AOI21_X1   g10200(.A1(new_n10389_), .A2(\asqrt[58] ), .B(new_n10392_), .ZN(new_n10393_));
  NOR2_X1    g10201(.A1(new_n10393_), .A2(new_n10388_), .ZN(new_n10394_));
  AOI22_X1   g10202(.A1(new_n10389_), .A2(\asqrt[58] ), .B1(new_n10387_), .B2(new_n10381_), .ZN(new_n10395_));
  NOR4_X1    g10203(.A1(new_n10104_), .A2(\asqrt[59] ), .A3(new_n9918_), .A4(new_n9923_), .ZN(new_n10396_));
  XOR2_X1    g10204(.A1(new_n10396_), .A2(new_n10109_), .Z(new_n10397_));
  AND2_X2    g10205(.A1(new_n10397_), .A2(new_n275_), .Z(new_n10398_));
  OAI21_X1   g10206(.A1(new_n10395_), .A2(new_n376_), .B(new_n10398_), .ZN(new_n10399_));
  NAND2_X1   g10207(.A1(new_n10399_), .A2(new_n10394_), .ZN(new_n10400_));
  NAND2_X1   g10208(.A1(new_n10376_), .A2(\asqrt[56] ), .ZN(new_n10401_));
  AOI21_X1   g10209(.A1(new_n10401_), .A2(new_n10375_), .B(new_n587_), .ZN(new_n10402_));
  OAI21_X1   g10210(.A1(new_n10381_), .A2(new_n10402_), .B(\asqrt[58] ), .ZN(new_n10403_));
  AOI21_X1   g10211(.A1(new_n10388_), .A2(new_n10403_), .B(new_n376_), .ZN(new_n10404_));
  OAI21_X1   g10212(.A1(new_n10394_), .A2(new_n10404_), .B(\asqrt[60] ), .ZN(new_n10405_));
  AOI21_X1   g10213(.A1(new_n10400_), .A2(new_n10405_), .B(new_n229_), .ZN(new_n10406_));
  NOR2_X1    g10214(.A1(new_n10091_), .A2(new_n196_), .ZN(new_n10407_));
  NOR2_X1    g10215(.A1(new_n10076_), .A2(\asqrt[62] ), .ZN(new_n10408_));
  NAND3_X1   g10216(.A1(new_n10408_), .A2(new_n10407_), .A3(new_n9937_), .ZN(new_n10409_));
  NOR2_X1    g10217(.A1(new_n10104_), .A2(new_n10409_), .ZN(new_n10410_));
  OR3_X2     g10218(.A1(\asqrt[24] ), .A2(new_n9937_), .A3(new_n10408_), .Z(new_n10411_));
  AOI21_X1   g10219(.A1(new_n10411_), .A2(new_n10407_), .B(new_n10410_), .ZN(new_n10412_));
  NOR4_X1    g10220(.A1(new_n10104_), .A2(\asqrt[61] ), .A3(new_n9931_), .A4(new_n9936_), .ZN(new_n10413_));
  XOR2_X1    g10221(.A1(new_n10413_), .A2(new_n10111_), .Z(new_n10414_));
  NOR2_X1    g10222(.A1(new_n10414_), .A2(new_n196_), .ZN(new_n10415_));
  INV_X1     g10223(.I(new_n10415_), .ZN(new_n10416_));
  NAND2_X1   g10224(.A1(new_n10159_), .A2(new_n10165_), .ZN(new_n10417_));
  NAND3_X1   g10225(.A1(new_n10417_), .A2(new_n10146_), .A3(new_n10182_), .ZN(new_n10418_));
  INV_X1     g10226(.I(new_n10083_), .ZN(new_n10419_));
  AOI21_X1   g10227(.A1(new_n10095_), .A2(new_n10419_), .B(new_n10085_), .ZN(new_n10420_));
  NOR3_X1    g10228(.A1(new_n10082_), .A2(new_n9607_), .A3(new_n9619_), .ZN(new_n10421_));
  NOR2_X1    g10229(.A1(new_n10421_), .A2(new_n10420_), .ZN(new_n10422_));
  NOR3_X1    g10230(.A1(new_n10132_), .A2(new_n9648_), .A3(\asqrt[24] ), .ZN(new_n10423_));
  AOI21_X1   g10231(.A1(new_n10117_), .A2(new_n9647_), .B(new_n10104_), .ZN(new_n10424_));
  NOR4_X1    g10232(.A1(new_n10423_), .A2(new_n10424_), .A3(\asqrt[26] ), .A4(new_n10102_), .ZN(new_n10425_));
  NOR2_X1    g10233(.A1(new_n10425_), .A2(new_n10422_), .ZN(new_n10426_));
  NOR3_X1    g10234(.A1(new_n10421_), .A2(new_n10420_), .A3(new_n10102_), .ZN(new_n10427_));
  NOR3_X1    g10235(.A1(new_n10104_), .A2(new_n9670_), .A3(new_n10140_), .ZN(new_n10428_));
  AOI21_X1   g10236(.A1(\asqrt[24] ), .A2(new_n10141_), .B(new_n9671_), .ZN(new_n10429_));
  NOR3_X1    g10237(.A1(new_n10429_), .A2(new_n10428_), .A3(\asqrt[27] ), .ZN(new_n10430_));
  OAI21_X1   g10238(.A1(new_n10427_), .A2(new_n9212_), .B(new_n10430_), .ZN(new_n10431_));
  NAND2_X1   g10239(.A1(new_n10426_), .A2(new_n10431_), .ZN(new_n10432_));
  OAI22_X1   g10240(.A1(new_n10425_), .A2(new_n10422_), .B1(new_n9212_), .B2(new_n10427_), .ZN(new_n10433_));
  AOI21_X1   g10241(.A1(new_n10433_), .A2(\asqrt[27] ), .B(new_n10157_), .ZN(new_n10434_));
  AOI22_X1   g10242(.A1(new_n10433_), .A2(\asqrt[27] ), .B1(new_n10426_), .B2(new_n10431_), .ZN(new_n10435_));
  OAI22_X1   g10243(.A1(new_n10435_), .A2(new_n8319_), .B1(new_n10434_), .B2(new_n10432_), .ZN(new_n10436_));
  AOI21_X1   g10244(.A1(new_n10436_), .A2(\asqrt[29] ), .B(new_n10172_), .ZN(new_n10437_));
  NOR2_X1    g10245(.A1(new_n10437_), .A2(new_n10418_), .ZN(new_n10438_));
  NAND2_X1   g10246(.A1(new_n10174_), .A2(new_n10179_), .ZN(new_n10439_));
  NAND2_X1   g10247(.A1(new_n10439_), .A2(new_n10438_), .ZN(new_n10440_));
  NAND2_X1   g10248(.A1(new_n10173_), .A2(new_n10174_), .ZN(new_n10441_));
  AOI21_X1   g10249(.A1(new_n10441_), .A2(\asqrt[31] ), .B(new_n10193_), .ZN(new_n10442_));
  NOR2_X1    g10250(.A1(new_n10442_), .A2(new_n10440_), .ZN(new_n10443_));
  AOI21_X1   g10251(.A1(new_n10173_), .A2(new_n10174_), .B(new_n7110_), .ZN(new_n10444_));
  OAI21_X1   g10252(.A1(new_n10180_), .A2(new_n10444_), .B(\asqrt[32] ), .ZN(new_n10445_));
  INV_X1     g10253(.I(new_n10202_), .ZN(new_n10446_));
  NAND2_X1   g10254(.A1(new_n10445_), .A2(new_n10446_), .ZN(new_n10447_));
  NAND2_X1   g10255(.A1(new_n10447_), .A2(new_n10443_), .ZN(new_n10448_));
  AOI22_X1   g10256(.A1(new_n10441_), .A2(\asqrt[31] ), .B1(new_n10439_), .B2(new_n10438_), .ZN(new_n10449_));
  OAI22_X1   g10257(.A1(new_n10449_), .A2(new_n6708_), .B1(new_n10442_), .B2(new_n10440_), .ZN(new_n10450_));
  AOI21_X1   g10258(.A1(new_n10450_), .A2(\asqrt[33] ), .B(new_n10209_), .ZN(new_n10451_));
  NOR2_X1    g10259(.A1(new_n10451_), .A2(new_n10448_), .ZN(new_n10452_));
  AOI22_X1   g10260(.A1(new_n10450_), .A2(\asqrt[33] ), .B1(new_n10447_), .B2(new_n10443_), .ZN(new_n10453_));
  INV_X1     g10261(.I(new_n10217_), .ZN(new_n10454_));
  OAI21_X1   g10262(.A1(new_n10453_), .A2(new_n5991_), .B(new_n10454_), .ZN(new_n10455_));
  NAND2_X1   g10263(.A1(new_n10455_), .A2(new_n10452_), .ZN(new_n10456_));
  OAI22_X1   g10264(.A1(new_n10453_), .A2(new_n5991_), .B1(new_n10451_), .B2(new_n10448_), .ZN(new_n10457_));
  AOI21_X1   g10265(.A1(new_n10457_), .A2(\asqrt[35] ), .B(new_n10224_), .ZN(new_n10458_));
  NOR2_X1    g10266(.A1(new_n10458_), .A2(new_n10456_), .ZN(new_n10459_));
  AOI22_X1   g10267(.A1(new_n10457_), .A2(\asqrt[35] ), .B1(new_n10455_), .B2(new_n10452_), .ZN(new_n10460_));
  INV_X1     g10268(.I(new_n10232_), .ZN(new_n10461_));
  OAI21_X1   g10269(.A1(new_n10460_), .A2(new_n5273_), .B(new_n10461_), .ZN(new_n10462_));
  NAND2_X1   g10270(.A1(new_n10462_), .A2(new_n10459_), .ZN(new_n10463_));
  OAI22_X1   g10271(.A1(new_n10460_), .A2(new_n5273_), .B1(new_n10458_), .B2(new_n10456_), .ZN(new_n10464_));
  AOI21_X1   g10272(.A1(new_n10464_), .A2(\asqrt[37] ), .B(new_n10239_), .ZN(new_n10465_));
  NOR2_X1    g10273(.A1(new_n10465_), .A2(new_n10463_), .ZN(new_n10466_));
  AOI22_X1   g10274(.A1(new_n10464_), .A2(\asqrt[37] ), .B1(new_n10462_), .B2(new_n10459_), .ZN(new_n10467_));
  INV_X1     g10275(.I(new_n10247_), .ZN(new_n10468_));
  OAI21_X1   g10276(.A1(new_n10467_), .A2(new_n4645_), .B(new_n10468_), .ZN(new_n10469_));
  NAND2_X1   g10277(.A1(new_n10469_), .A2(new_n10466_), .ZN(new_n10470_));
  OAI22_X1   g10278(.A1(new_n10467_), .A2(new_n4645_), .B1(new_n10465_), .B2(new_n10463_), .ZN(new_n10471_));
  AOI21_X1   g10279(.A1(new_n10471_), .A2(\asqrt[39] ), .B(new_n10254_), .ZN(new_n10472_));
  NOR2_X1    g10280(.A1(new_n10472_), .A2(new_n10470_), .ZN(new_n10473_));
  AOI22_X1   g10281(.A1(new_n10471_), .A2(\asqrt[39] ), .B1(new_n10469_), .B2(new_n10466_), .ZN(new_n10474_));
  INV_X1     g10282(.I(new_n10262_), .ZN(new_n10475_));
  OAI21_X1   g10283(.A1(new_n10474_), .A2(new_n4018_), .B(new_n10475_), .ZN(new_n10476_));
  NAND2_X1   g10284(.A1(new_n10476_), .A2(new_n10473_), .ZN(new_n10477_));
  OAI22_X1   g10285(.A1(new_n10474_), .A2(new_n4018_), .B1(new_n10472_), .B2(new_n10470_), .ZN(new_n10478_));
  AOI21_X1   g10286(.A1(new_n10478_), .A2(\asqrt[41] ), .B(new_n10269_), .ZN(new_n10479_));
  NOR2_X1    g10287(.A1(new_n10479_), .A2(new_n10477_), .ZN(new_n10480_));
  AOI22_X1   g10288(.A1(new_n10478_), .A2(\asqrt[41] ), .B1(new_n10476_), .B2(new_n10473_), .ZN(new_n10481_));
  INV_X1     g10289(.I(new_n10277_), .ZN(new_n10482_));
  OAI21_X1   g10290(.A1(new_n10481_), .A2(new_n3481_), .B(new_n10482_), .ZN(new_n10483_));
  NAND2_X1   g10291(.A1(new_n10483_), .A2(new_n10480_), .ZN(new_n10484_));
  OAI22_X1   g10292(.A1(new_n10481_), .A2(new_n3481_), .B1(new_n10479_), .B2(new_n10477_), .ZN(new_n10485_));
  AOI21_X1   g10293(.A1(new_n10485_), .A2(\asqrt[43] ), .B(new_n10284_), .ZN(new_n10486_));
  NOR2_X1    g10294(.A1(new_n10486_), .A2(new_n10484_), .ZN(new_n10487_));
  AOI22_X1   g10295(.A1(new_n10485_), .A2(\asqrt[43] ), .B1(new_n10483_), .B2(new_n10480_), .ZN(new_n10488_));
  INV_X1     g10296(.I(new_n10292_), .ZN(new_n10489_));
  OAI21_X1   g10297(.A1(new_n10488_), .A2(new_n2941_), .B(new_n10489_), .ZN(new_n10490_));
  NAND2_X1   g10298(.A1(new_n10490_), .A2(new_n10487_), .ZN(new_n10491_));
  OAI22_X1   g10299(.A1(new_n10488_), .A2(new_n2941_), .B1(new_n10486_), .B2(new_n10484_), .ZN(new_n10492_));
  AOI21_X1   g10300(.A1(new_n10492_), .A2(\asqrt[45] ), .B(new_n10299_), .ZN(new_n10493_));
  NOR2_X1    g10301(.A1(new_n10493_), .A2(new_n10491_), .ZN(new_n10494_));
  AOI22_X1   g10302(.A1(new_n10492_), .A2(\asqrt[45] ), .B1(new_n10490_), .B2(new_n10487_), .ZN(new_n10495_));
  INV_X1     g10303(.I(new_n10307_), .ZN(new_n10496_));
  OAI21_X1   g10304(.A1(new_n10495_), .A2(new_n2488_), .B(new_n10496_), .ZN(new_n10497_));
  NAND2_X1   g10305(.A1(new_n10497_), .A2(new_n10494_), .ZN(new_n10498_));
  OAI22_X1   g10306(.A1(new_n10495_), .A2(new_n2488_), .B1(new_n10493_), .B2(new_n10491_), .ZN(new_n10499_));
  AOI21_X1   g10307(.A1(new_n10499_), .A2(\asqrt[47] ), .B(new_n10314_), .ZN(new_n10500_));
  NOR2_X1    g10308(.A1(new_n10500_), .A2(new_n10498_), .ZN(new_n10501_));
  AOI22_X1   g10309(.A1(new_n10499_), .A2(\asqrt[47] ), .B1(new_n10497_), .B2(new_n10494_), .ZN(new_n10502_));
  INV_X1     g10310(.I(new_n10322_), .ZN(new_n10503_));
  OAI21_X1   g10311(.A1(new_n10502_), .A2(new_n2046_), .B(new_n10503_), .ZN(new_n10504_));
  NAND2_X1   g10312(.A1(new_n10504_), .A2(new_n10501_), .ZN(new_n10505_));
  OAI22_X1   g10313(.A1(new_n10502_), .A2(new_n2046_), .B1(new_n10500_), .B2(new_n10498_), .ZN(new_n10506_));
  AOI21_X1   g10314(.A1(new_n10506_), .A2(\asqrt[49] ), .B(new_n10329_), .ZN(new_n10507_));
  NOR2_X1    g10315(.A1(new_n10507_), .A2(new_n10505_), .ZN(new_n10508_));
  AOI22_X1   g10316(.A1(new_n10506_), .A2(\asqrt[49] ), .B1(new_n10504_), .B2(new_n10501_), .ZN(new_n10509_));
  INV_X1     g10317(.I(new_n10337_), .ZN(new_n10510_));
  OAI21_X1   g10318(.A1(new_n10509_), .A2(new_n1595_), .B(new_n10510_), .ZN(new_n10511_));
  NAND2_X1   g10319(.A1(new_n10511_), .A2(new_n10508_), .ZN(new_n10512_));
  OAI22_X1   g10320(.A1(new_n10509_), .A2(new_n1595_), .B1(new_n10507_), .B2(new_n10505_), .ZN(new_n10513_));
  AOI21_X1   g10321(.A1(new_n10513_), .A2(\asqrt[51] ), .B(new_n10344_), .ZN(new_n10514_));
  NOR2_X1    g10322(.A1(new_n10514_), .A2(new_n10512_), .ZN(new_n10515_));
  AOI22_X1   g10323(.A1(new_n10513_), .A2(\asqrt[51] ), .B1(new_n10511_), .B2(new_n10508_), .ZN(new_n10516_));
  INV_X1     g10324(.I(new_n10352_), .ZN(new_n10517_));
  OAI21_X1   g10325(.A1(new_n10516_), .A2(new_n1260_), .B(new_n10517_), .ZN(new_n10518_));
  NAND2_X1   g10326(.A1(new_n10518_), .A2(new_n10515_), .ZN(new_n10519_));
  OAI22_X1   g10327(.A1(new_n10516_), .A2(new_n1260_), .B1(new_n10514_), .B2(new_n10512_), .ZN(new_n10520_));
  AOI21_X1   g10328(.A1(new_n10520_), .A2(\asqrt[53] ), .B(new_n10359_), .ZN(new_n10521_));
  NOR2_X1    g10329(.A1(new_n10521_), .A2(new_n10519_), .ZN(new_n10522_));
  AOI22_X1   g10330(.A1(new_n10520_), .A2(\asqrt[53] ), .B1(new_n10518_), .B2(new_n10515_), .ZN(new_n10523_));
  INV_X1     g10331(.I(new_n10366_), .ZN(new_n10524_));
  OAI21_X1   g10332(.A1(new_n10523_), .A2(new_n970_), .B(new_n10524_), .ZN(new_n10525_));
  NAND2_X1   g10333(.A1(new_n10525_), .A2(new_n10522_), .ZN(new_n10526_));
  OAI22_X1   g10334(.A1(new_n10523_), .A2(new_n970_), .B1(new_n10521_), .B2(new_n10519_), .ZN(new_n10527_));
  AOI21_X1   g10335(.A1(new_n10527_), .A2(\asqrt[55] ), .B(new_n10372_), .ZN(new_n10528_));
  NOR2_X1    g10336(.A1(new_n10528_), .A2(new_n10526_), .ZN(new_n10529_));
  AOI22_X1   g10337(.A1(new_n10527_), .A2(\asqrt[55] ), .B1(new_n10525_), .B2(new_n10522_), .ZN(new_n10530_));
  INV_X1     g10338(.I(new_n10379_), .ZN(new_n10531_));
  OAI21_X1   g10339(.A1(new_n10530_), .A2(new_n724_), .B(new_n10531_), .ZN(new_n10532_));
  NAND2_X1   g10340(.A1(new_n10532_), .A2(new_n10529_), .ZN(new_n10533_));
  OAI22_X1   g10341(.A1(new_n10530_), .A2(new_n724_), .B1(new_n10528_), .B2(new_n10526_), .ZN(new_n10534_));
  AOI21_X1   g10342(.A1(new_n10534_), .A2(\asqrt[57] ), .B(new_n10385_), .ZN(new_n10535_));
  NOR2_X1    g10343(.A1(new_n10535_), .A2(new_n10533_), .ZN(new_n10536_));
  AOI22_X1   g10344(.A1(new_n10534_), .A2(\asqrt[57] ), .B1(new_n10532_), .B2(new_n10529_), .ZN(new_n10537_));
  INV_X1     g10345(.I(new_n10392_), .ZN(new_n10538_));
  OAI21_X1   g10346(.A1(new_n10537_), .A2(new_n504_), .B(new_n10538_), .ZN(new_n10539_));
  NAND2_X1   g10347(.A1(new_n10539_), .A2(new_n10536_), .ZN(new_n10540_));
  NAND2_X1   g10348(.A1(new_n10520_), .A2(\asqrt[53] ), .ZN(new_n10541_));
  AOI21_X1   g10349(.A1(new_n10541_), .A2(new_n10519_), .B(new_n970_), .ZN(new_n10542_));
  OAI21_X1   g10350(.A1(new_n10522_), .A2(new_n10542_), .B(\asqrt[55] ), .ZN(new_n10543_));
  AOI21_X1   g10351(.A1(new_n10526_), .A2(new_n10543_), .B(new_n724_), .ZN(new_n10544_));
  OAI21_X1   g10352(.A1(new_n10529_), .A2(new_n10544_), .B(\asqrt[57] ), .ZN(new_n10545_));
  AOI21_X1   g10353(.A1(new_n10533_), .A2(new_n10545_), .B(new_n504_), .ZN(new_n10546_));
  OAI21_X1   g10354(.A1(new_n10536_), .A2(new_n10546_), .B(\asqrt[59] ), .ZN(new_n10547_));
  AOI21_X1   g10355(.A1(new_n10547_), .A2(new_n10398_), .B(new_n10540_), .ZN(new_n10548_));
  OAI22_X1   g10356(.A1(new_n10537_), .A2(new_n504_), .B1(new_n10535_), .B2(new_n10533_), .ZN(new_n10549_));
  AOI22_X1   g10357(.A1(new_n10549_), .A2(\asqrt[59] ), .B1(new_n10539_), .B2(new_n10536_), .ZN(new_n10550_));
  NOR4_X1    g10358(.A1(new_n10104_), .A2(\asqrt[60] ), .A3(new_n9925_), .A4(new_n10073_), .ZN(new_n10551_));
  XOR2_X1    g10359(.A1(new_n10551_), .A2(new_n10126_), .Z(new_n10552_));
  NAND2_X1   g10360(.A1(new_n10552_), .A2(new_n229_), .ZN(new_n10553_));
  INV_X1     g10361(.I(new_n10553_), .ZN(new_n10554_));
  OAI21_X1   g10362(.A1(new_n10550_), .A2(new_n275_), .B(new_n10554_), .ZN(new_n10555_));
  NAND2_X1   g10363(.A1(new_n10555_), .A2(new_n10548_), .ZN(new_n10556_));
  INV_X1     g10364(.I(new_n10414_), .ZN(new_n10557_));
  NOR2_X1    g10365(.A1(new_n10557_), .A2(\asqrt[62] ), .ZN(new_n10558_));
  INV_X1     g10366(.I(new_n10558_), .ZN(new_n10559_));
  NAND2_X1   g10367(.A1(new_n10406_), .A2(new_n10559_), .ZN(new_n10560_));
  OAI21_X1   g10368(.A1(new_n10560_), .A2(new_n10556_), .B(new_n10416_), .ZN(new_n10561_));
  NOR3_X1    g10369(.A1(\asqrt[24] ), .A2(new_n9640_), .A3(new_n10077_), .ZN(new_n10562_));
  OAI21_X1   g10370(.A1(new_n10562_), .A2(new_n10089_), .B(new_n231_), .ZN(new_n10563_));
  OAI21_X1   g10371(.A1(new_n10561_), .A2(new_n10563_), .B(new_n10412_), .ZN(new_n10564_));
  OAI21_X1   g10372(.A1(new_n9640_), .A2(new_n9941_), .B(\asqrt[24] ), .ZN(new_n10565_));
  XOR2_X1    g10373(.A1(new_n9941_), .A2(\asqrt[63] ), .Z(new_n10566_));
  NAND2_X1   g10374(.A1(new_n10565_), .A2(new_n10566_), .ZN(new_n10567_));
  INV_X1     g10375(.I(new_n10567_), .ZN(new_n10568_));
  INV_X1     g10376(.I(new_n10412_), .ZN(new_n10569_));
  OAI22_X1   g10377(.A1(new_n10395_), .A2(new_n376_), .B1(new_n10393_), .B2(new_n10388_), .ZN(new_n10570_));
  AOI21_X1   g10378(.A1(new_n10570_), .A2(\asqrt[60] ), .B(new_n10553_), .ZN(new_n10571_));
  AOI22_X1   g10379(.A1(new_n10570_), .A2(\asqrt[60] ), .B1(new_n10399_), .B2(new_n10394_), .ZN(new_n10572_));
  OAI22_X1   g10380(.A1(new_n10572_), .A2(new_n229_), .B1(new_n10571_), .B2(new_n10400_), .ZN(new_n10573_));
  NOR4_X1    g10381(.A1(new_n10573_), .A2(\asqrt[62] ), .A3(new_n10569_), .A4(new_n10414_), .ZN(new_n10574_));
  NAND2_X1   g10382(.A1(new_n10574_), .A2(new_n10568_), .ZN(new_n10575_));
  NAND3_X1   g10383(.A1(new_n10098_), .A2(new_n9627_), .A3(new_n9640_), .ZN(new_n10576_));
  NOR3_X1    g10384(.A1(new_n10575_), .A2(new_n10564_), .A3(new_n10576_), .ZN(\asqrt[23] ));
  NAND2_X1   g10385(.A1(new_n10400_), .A2(new_n10405_), .ZN(new_n10578_));
  NOR3_X1    g10386(.A1(new_n10578_), .A2(\asqrt[61] ), .A3(new_n10552_), .ZN(new_n10579_));
  NAND2_X1   g10387(.A1(\asqrt[23] ), .A2(new_n10579_), .ZN(new_n10580_));
  XOR2_X1    g10388(.A1(new_n10580_), .A2(new_n10406_), .Z(new_n10581_));
  INV_X1     g10389(.I(new_n10581_), .ZN(new_n10582_));
  INV_X1     g10390(.I(\a[46] ), .ZN(new_n10583_));
  NOR2_X1    g10391(.A1(\a[44] ), .A2(\a[45] ), .ZN(new_n10584_));
  INV_X1     g10392(.I(new_n10584_), .ZN(new_n10585_));
  NOR3_X1    g10393(.A1(new_n10115_), .A2(new_n10583_), .A3(new_n10585_), .ZN(new_n10586_));
  NAND2_X1   g10394(.A1(new_n10130_), .A2(new_n10586_), .ZN(new_n10587_));
  XOR2_X1    g10395(.A1(new_n10587_), .A2(\a[47] ), .Z(new_n10588_));
  INV_X1     g10396(.I(\a[47] ), .ZN(new_n10589_));
  NOR4_X1    g10397(.A1(new_n10575_), .A2(new_n10564_), .A3(new_n10589_), .A4(new_n10576_), .ZN(new_n10590_));
  NOR2_X1    g10398(.A1(new_n10589_), .A2(\a[46] ), .ZN(new_n10591_));
  OAI21_X1   g10399(.A1(new_n10590_), .A2(new_n10591_), .B(new_n10588_), .ZN(new_n10592_));
  INV_X1     g10400(.I(new_n10588_), .ZN(new_n10593_));
  NOR2_X1    g10401(.A1(new_n10571_), .A2(new_n10400_), .ZN(new_n10594_));
  NOR3_X1    g10402(.A1(new_n10572_), .A2(new_n229_), .A3(new_n10558_), .ZN(new_n10595_));
  AOI21_X1   g10403(.A1(new_n10595_), .A2(new_n10594_), .B(new_n10415_), .ZN(new_n10596_));
  INV_X1     g10404(.I(new_n10563_), .ZN(new_n10597_));
  AOI21_X1   g10405(.A1(new_n10596_), .A2(new_n10597_), .B(new_n10569_), .ZN(new_n10598_));
  AOI21_X1   g10406(.A1(new_n10573_), .A2(\asqrt[62] ), .B(new_n10412_), .ZN(new_n10599_));
  AOI21_X1   g10407(.A1(new_n10540_), .A2(new_n10547_), .B(new_n275_), .ZN(new_n10600_));
  OAI21_X1   g10408(.A1(new_n10548_), .A2(new_n10600_), .B(\asqrt[61] ), .ZN(new_n10601_));
  NAND4_X1   g10409(.A1(new_n10556_), .A2(new_n10601_), .A3(new_n196_), .A4(new_n10557_), .ZN(new_n10602_));
  NOR3_X1    g10410(.A1(new_n10599_), .A2(new_n10567_), .A3(new_n10602_), .ZN(new_n10603_));
  INV_X1     g10411(.I(new_n10576_), .ZN(new_n10604_));
  NAND4_X1   g10412(.A1(new_n10603_), .A2(\a[47] ), .A3(new_n10598_), .A4(new_n10604_), .ZN(new_n10605_));
  NAND3_X1   g10413(.A1(new_n10605_), .A2(\a[46] ), .A3(new_n10593_), .ZN(new_n10606_));
  NAND2_X1   g10414(.A1(new_n10592_), .A2(new_n10606_), .ZN(new_n10607_));
  NOR2_X1    g10415(.A1(new_n10575_), .A2(new_n10564_), .ZN(new_n10608_));
  NAND4_X1   g10416(.A1(new_n10094_), .A2(new_n10086_), .A3(new_n9640_), .A4(new_n10129_), .ZN(new_n10609_));
  NOR2_X1    g10417(.A1(new_n10104_), .A2(new_n10583_), .ZN(new_n10610_));
  XOR2_X1    g10418(.A1(new_n10610_), .A2(new_n10609_), .Z(new_n10611_));
  NOR2_X1    g10419(.A1(new_n10611_), .A2(new_n10585_), .ZN(new_n10612_));
  INV_X1     g10420(.I(new_n10612_), .ZN(new_n10613_));
  NAND3_X1   g10421(.A1(new_n10603_), .A2(new_n10598_), .A3(new_n10604_), .ZN(new_n10614_));
  NOR4_X1    g10422(.A1(new_n10601_), .A2(new_n10400_), .A3(new_n10571_), .A4(new_n10558_), .ZN(new_n10615_));
  NOR3_X1    g10423(.A1(new_n10615_), .A2(new_n10415_), .A3(new_n10563_), .ZN(new_n10616_));
  AOI22_X1   g10424(.A1(new_n10578_), .A2(\asqrt[61] ), .B1(new_n10555_), .B2(new_n10548_), .ZN(new_n10617_));
  NAND4_X1   g10425(.A1(new_n10617_), .A2(new_n196_), .A3(new_n10412_), .A4(new_n10557_), .ZN(new_n10618_));
  OAI21_X1   g10426(.A1(new_n10616_), .A2(new_n10569_), .B(new_n10618_), .ZN(new_n10619_));
  NOR2_X1    g10427(.A1(new_n10568_), .A2(new_n10604_), .ZN(new_n10620_));
  NAND2_X1   g10428(.A1(new_n10620_), .A2(\asqrt[24] ), .ZN(new_n10621_));
  OAI21_X1   g10429(.A1(new_n10619_), .A2(new_n10621_), .B(new_n9607_), .ZN(new_n10622_));
  NAND3_X1   g10430(.A1(new_n10622_), .A2(new_n9615_), .A3(new_n10614_), .ZN(new_n10623_));
  NAND4_X1   g10431(.A1(new_n10406_), .A2(new_n10548_), .A3(new_n10555_), .A4(new_n10559_), .ZN(new_n10624_));
  NAND3_X1   g10432(.A1(new_n10624_), .A2(new_n10416_), .A3(new_n10597_), .ZN(new_n10625_));
  AOI21_X1   g10433(.A1(new_n10412_), .A2(new_n10625_), .B(new_n10574_), .ZN(new_n10626_));
  INV_X1     g10434(.I(new_n10621_), .ZN(new_n10627_));
  AOI21_X1   g10435(.A1(new_n10626_), .A2(new_n10627_), .B(\a[48] ), .ZN(new_n10628_));
  OAI21_X1   g10436(.A1(new_n10628_), .A2(new_n9616_), .B(\asqrt[23] ), .ZN(new_n10629_));
  NAND4_X1   g10437(.A1(new_n10623_), .A2(new_n10629_), .A3(new_n9672_), .A4(new_n10613_), .ZN(new_n10630_));
  NAND2_X1   g10438(.A1(new_n10630_), .A2(new_n10607_), .ZN(new_n10631_));
  NAND3_X1   g10439(.A1(new_n10592_), .A2(new_n10606_), .A3(new_n10613_), .ZN(new_n10632_));
  INV_X1     g10440(.I(new_n9618_), .ZN(new_n10633_));
  NOR2_X1    g10441(.A1(new_n10104_), .A2(\a[48] ), .ZN(new_n10634_));
  OAI22_X1   g10442(.A1(new_n10634_), .A2(\a[49] ), .B1(\a[48] ), .B2(new_n10095_), .ZN(new_n10635_));
  NAND2_X1   g10443(.A1(\asqrt[24] ), .A2(\a[48] ), .ZN(new_n10636_));
  AND3_X2    g10444(.A1(new_n10635_), .A2(new_n10633_), .A3(new_n10636_), .Z(new_n10637_));
  NAND3_X1   g10445(.A1(\asqrt[23] ), .A2(new_n10103_), .A3(new_n10637_), .ZN(new_n10638_));
  INV_X1     g10446(.I(new_n10637_), .ZN(new_n10639_));
  OAI21_X1   g10447(.A1(new_n10614_), .A2(new_n10639_), .B(new_n10102_), .ZN(new_n10640_));
  NAND3_X1   g10448(.A1(new_n10638_), .A2(new_n10640_), .A3(new_n9212_), .ZN(new_n10641_));
  AOI21_X1   g10449(.A1(new_n10632_), .A2(\asqrt[25] ), .B(new_n10641_), .ZN(new_n10642_));
  NOR2_X1    g10450(.A1(new_n10631_), .A2(new_n10642_), .ZN(new_n10643_));
  AOI22_X1   g10451(.A1(new_n10630_), .A2(new_n10607_), .B1(\asqrt[25] ), .B2(new_n10632_), .ZN(new_n10644_));
  AOI21_X1   g10452(.A1(new_n10133_), .A2(new_n10118_), .B(\asqrt[26] ), .ZN(new_n10645_));
  AND4_X2    g10453(.A1(new_n10427_), .A2(\asqrt[23] ), .A3(new_n10147_), .A4(new_n10645_), .Z(new_n10646_));
  NOR2_X1    g10454(.A1(new_n10427_), .A2(new_n9212_), .ZN(new_n10647_));
  NOR3_X1    g10455(.A1(new_n10646_), .A2(\asqrt[27] ), .A3(new_n10647_), .ZN(new_n10648_));
  OAI21_X1   g10456(.A1(new_n10644_), .A2(new_n9212_), .B(new_n10648_), .ZN(new_n10649_));
  NAND2_X1   g10457(.A1(new_n10649_), .A2(new_n10643_), .ZN(new_n10650_));
  OAI22_X1   g10458(.A1(new_n10644_), .A2(new_n9212_), .B1(new_n10631_), .B2(new_n10642_), .ZN(new_n10651_));
  NAND2_X1   g10459(.A1(new_n10142_), .A2(new_n10143_), .ZN(new_n10652_));
  NAND4_X1   g10460(.A1(\asqrt[23] ), .A2(new_n8763_), .A3(new_n10652_), .A4(new_n10181_), .ZN(new_n10653_));
  XOR2_X1    g10461(.A1(new_n10653_), .A2(new_n10148_), .Z(new_n10654_));
  NAND2_X1   g10462(.A1(new_n10654_), .A2(new_n8319_), .ZN(new_n10655_));
  AOI21_X1   g10463(.A1(new_n10651_), .A2(\asqrt[27] ), .B(new_n10655_), .ZN(new_n10656_));
  NOR2_X1    g10464(.A1(new_n10656_), .A2(new_n10650_), .ZN(new_n10657_));
  AOI22_X1   g10465(.A1(new_n10651_), .A2(\asqrt[27] ), .B1(new_n10649_), .B2(new_n10643_), .ZN(new_n10658_));
  NOR2_X1    g10466(.A1(new_n10155_), .A2(new_n10153_), .ZN(new_n10659_));
  NOR4_X1    g10467(.A1(new_n10614_), .A2(\asqrt[28] ), .A3(new_n10659_), .A4(new_n10183_), .ZN(new_n10660_));
  XOR2_X1    g10468(.A1(new_n10660_), .A2(new_n10159_), .Z(new_n10661_));
  NAND2_X1   g10469(.A1(new_n10661_), .A2(new_n7931_), .ZN(new_n10662_));
  INV_X1     g10470(.I(new_n10662_), .ZN(new_n10663_));
  OAI21_X1   g10471(.A1(new_n10658_), .A2(new_n8319_), .B(new_n10663_), .ZN(new_n10664_));
  NAND2_X1   g10472(.A1(new_n10664_), .A2(new_n10657_), .ZN(new_n10665_));
  OAI22_X1   g10473(.A1(new_n10658_), .A2(new_n8319_), .B1(new_n10656_), .B2(new_n10650_), .ZN(new_n10666_));
  NOR4_X1    g10474(.A1(new_n10614_), .A2(\asqrt[29] ), .A3(new_n10163_), .A4(new_n10436_), .ZN(new_n10667_));
  XNOR2_X1   g10475(.A1(new_n10667_), .A2(new_n10167_), .ZN(new_n10668_));
  NAND2_X1   g10476(.A1(new_n10668_), .A2(new_n7517_), .ZN(new_n10669_));
  AOI21_X1   g10477(.A1(new_n10666_), .A2(\asqrt[29] ), .B(new_n10669_), .ZN(new_n10670_));
  NOR2_X1    g10478(.A1(new_n10670_), .A2(new_n10665_), .ZN(new_n10671_));
  AOI22_X1   g10479(.A1(new_n10666_), .A2(\asqrt[29] ), .B1(new_n10664_), .B2(new_n10657_), .ZN(new_n10672_));
  NOR4_X1    g10480(.A1(new_n10614_), .A2(\asqrt[30] ), .A3(new_n10171_), .A4(new_n10188_), .ZN(new_n10673_));
  XOR2_X1    g10481(.A1(new_n10673_), .A2(new_n10174_), .Z(new_n10674_));
  NAND2_X1   g10482(.A1(new_n10674_), .A2(new_n7110_), .ZN(new_n10675_));
  INV_X1     g10483(.I(new_n10675_), .ZN(new_n10676_));
  OAI21_X1   g10484(.A1(new_n10672_), .A2(new_n7517_), .B(new_n10676_), .ZN(new_n10677_));
  NAND2_X1   g10485(.A1(new_n10677_), .A2(new_n10671_), .ZN(new_n10678_));
  OAI22_X1   g10486(.A1(new_n10672_), .A2(new_n7517_), .B1(new_n10670_), .B2(new_n10665_), .ZN(new_n10679_));
  NOR4_X1    g10487(.A1(new_n10614_), .A2(\asqrt[31] ), .A3(new_n10177_), .A4(new_n10441_), .ZN(new_n10680_));
  XNOR2_X1   g10488(.A1(new_n10680_), .A2(new_n10444_), .ZN(new_n10681_));
  NAND2_X1   g10489(.A1(new_n10681_), .A2(new_n6708_), .ZN(new_n10682_));
  AOI21_X1   g10490(.A1(new_n10679_), .A2(\asqrt[31] ), .B(new_n10682_), .ZN(new_n10683_));
  NOR2_X1    g10491(.A1(new_n10683_), .A2(new_n10678_), .ZN(new_n10684_));
  AOI22_X1   g10492(.A1(new_n10679_), .A2(\asqrt[31] ), .B1(new_n10677_), .B2(new_n10671_), .ZN(new_n10685_));
  NOR4_X1    g10493(.A1(new_n10614_), .A2(\asqrt[32] ), .A3(new_n10192_), .A4(new_n10198_), .ZN(new_n10686_));
  XOR2_X1    g10494(.A1(new_n10686_), .A2(new_n10445_), .Z(new_n10687_));
  NAND2_X1   g10495(.A1(new_n10687_), .A2(new_n6365_), .ZN(new_n10688_));
  INV_X1     g10496(.I(new_n10688_), .ZN(new_n10689_));
  OAI21_X1   g10497(.A1(new_n10685_), .A2(new_n6708_), .B(new_n10689_), .ZN(new_n10690_));
  NAND2_X1   g10498(.A1(new_n10690_), .A2(new_n10684_), .ZN(new_n10691_));
  OAI22_X1   g10499(.A1(new_n10685_), .A2(new_n6708_), .B1(new_n10683_), .B2(new_n10678_), .ZN(new_n10692_));
  NAND2_X1   g10500(.A1(new_n10450_), .A2(\asqrt[33] ), .ZN(new_n10693_));
  NOR4_X1    g10501(.A1(new_n10614_), .A2(\asqrt[33] ), .A3(new_n10201_), .A4(new_n10450_), .ZN(new_n10694_));
  XOR2_X1    g10502(.A1(new_n10694_), .A2(new_n10693_), .Z(new_n10695_));
  NAND2_X1   g10503(.A1(new_n10695_), .A2(new_n5991_), .ZN(new_n10696_));
  AOI21_X1   g10504(.A1(new_n10692_), .A2(\asqrt[33] ), .B(new_n10696_), .ZN(new_n10697_));
  NOR2_X1    g10505(.A1(new_n10697_), .A2(new_n10691_), .ZN(new_n10698_));
  AOI22_X1   g10506(.A1(new_n10692_), .A2(\asqrt[33] ), .B1(new_n10690_), .B2(new_n10684_), .ZN(new_n10699_));
  NOR4_X1    g10507(.A1(new_n10614_), .A2(\asqrt[34] ), .A3(new_n10208_), .A4(new_n10213_), .ZN(new_n10700_));
  AOI21_X1   g10508(.A1(new_n10693_), .A2(new_n10448_), .B(new_n5991_), .ZN(new_n10701_));
  NOR2_X1    g10509(.A1(new_n10700_), .A2(new_n10701_), .ZN(new_n10702_));
  NAND2_X1   g10510(.A1(new_n10702_), .A2(new_n5626_), .ZN(new_n10703_));
  INV_X1     g10511(.I(new_n10703_), .ZN(new_n10704_));
  OAI21_X1   g10512(.A1(new_n10699_), .A2(new_n5991_), .B(new_n10704_), .ZN(new_n10705_));
  NAND2_X1   g10513(.A1(new_n10705_), .A2(new_n10698_), .ZN(new_n10706_));
  OAI22_X1   g10514(.A1(new_n10699_), .A2(new_n5991_), .B1(new_n10697_), .B2(new_n10691_), .ZN(new_n10707_));
  NAND2_X1   g10515(.A1(new_n10457_), .A2(\asqrt[35] ), .ZN(new_n10708_));
  NOR4_X1    g10516(.A1(new_n10614_), .A2(\asqrt[35] ), .A3(new_n10216_), .A4(new_n10457_), .ZN(new_n10709_));
  XOR2_X1    g10517(.A1(new_n10709_), .A2(new_n10708_), .Z(new_n10710_));
  NAND2_X1   g10518(.A1(new_n10710_), .A2(new_n5273_), .ZN(new_n10711_));
  AOI21_X1   g10519(.A1(new_n10707_), .A2(\asqrt[35] ), .B(new_n10711_), .ZN(new_n10712_));
  NOR2_X1    g10520(.A1(new_n10712_), .A2(new_n10706_), .ZN(new_n10713_));
  AOI22_X1   g10521(.A1(new_n10707_), .A2(\asqrt[35] ), .B1(new_n10705_), .B2(new_n10698_), .ZN(new_n10714_));
  NOR4_X1    g10522(.A1(new_n10614_), .A2(\asqrt[36] ), .A3(new_n10223_), .A4(new_n10228_), .ZN(new_n10715_));
  AOI21_X1   g10523(.A1(new_n10708_), .A2(new_n10456_), .B(new_n5273_), .ZN(new_n10716_));
  NOR2_X1    g10524(.A1(new_n10715_), .A2(new_n10716_), .ZN(new_n10717_));
  NAND2_X1   g10525(.A1(new_n10717_), .A2(new_n4973_), .ZN(new_n10718_));
  INV_X1     g10526(.I(new_n10718_), .ZN(new_n10719_));
  OAI21_X1   g10527(.A1(new_n10714_), .A2(new_n5273_), .B(new_n10719_), .ZN(new_n10720_));
  NAND2_X1   g10528(.A1(new_n10720_), .A2(new_n10713_), .ZN(new_n10721_));
  OAI22_X1   g10529(.A1(new_n10714_), .A2(new_n5273_), .B1(new_n10712_), .B2(new_n10706_), .ZN(new_n10722_));
  NAND2_X1   g10530(.A1(new_n10464_), .A2(\asqrt[37] ), .ZN(new_n10723_));
  NOR4_X1    g10531(.A1(new_n10614_), .A2(\asqrt[37] ), .A3(new_n10231_), .A4(new_n10464_), .ZN(new_n10724_));
  XOR2_X1    g10532(.A1(new_n10724_), .A2(new_n10723_), .Z(new_n10725_));
  NAND2_X1   g10533(.A1(new_n10725_), .A2(new_n4645_), .ZN(new_n10726_));
  AOI21_X1   g10534(.A1(new_n10722_), .A2(\asqrt[37] ), .B(new_n10726_), .ZN(new_n10727_));
  NOR2_X1    g10535(.A1(new_n10727_), .A2(new_n10721_), .ZN(new_n10728_));
  AOI22_X1   g10536(.A1(new_n10722_), .A2(\asqrt[37] ), .B1(new_n10720_), .B2(new_n10713_), .ZN(new_n10729_));
  NOR4_X1    g10537(.A1(new_n10614_), .A2(\asqrt[38] ), .A3(new_n10238_), .A4(new_n10243_), .ZN(new_n10730_));
  AOI21_X1   g10538(.A1(new_n10723_), .A2(new_n10463_), .B(new_n4645_), .ZN(new_n10731_));
  NOR2_X1    g10539(.A1(new_n10730_), .A2(new_n10731_), .ZN(new_n10732_));
  NAND2_X1   g10540(.A1(new_n10732_), .A2(new_n4330_), .ZN(new_n10733_));
  INV_X1     g10541(.I(new_n10733_), .ZN(new_n10734_));
  OAI21_X1   g10542(.A1(new_n10729_), .A2(new_n4645_), .B(new_n10734_), .ZN(new_n10735_));
  NAND2_X1   g10543(.A1(new_n10735_), .A2(new_n10728_), .ZN(new_n10736_));
  OAI22_X1   g10544(.A1(new_n10729_), .A2(new_n4645_), .B1(new_n10727_), .B2(new_n10721_), .ZN(new_n10737_));
  NAND2_X1   g10545(.A1(new_n10471_), .A2(\asqrt[39] ), .ZN(new_n10738_));
  NOR4_X1    g10546(.A1(new_n10614_), .A2(\asqrt[39] ), .A3(new_n10246_), .A4(new_n10471_), .ZN(new_n10739_));
  XOR2_X1    g10547(.A1(new_n10739_), .A2(new_n10738_), .Z(new_n10740_));
  NAND2_X1   g10548(.A1(new_n10740_), .A2(new_n4018_), .ZN(new_n10741_));
  AOI21_X1   g10549(.A1(new_n10737_), .A2(\asqrt[39] ), .B(new_n10741_), .ZN(new_n10742_));
  NOR2_X1    g10550(.A1(new_n10742_), .A2(new_n10736_), .ZN(new_n10743_));
  AOI22_X1   g10551(.A1(new_n10737_), .A2(\asqrt[39] ), .B1(new_n10735_), .B2(new_n10728_), .ZN(new_n10744_));
  NOR4_X1    g10552(.A1(new_n10614_), .A2(\asqrt[40] ), .A3(new_n10253_), .A4(new_n10258_), .ZN(new_n10745_));
  AOI21_X1   g10553(.A1(new_n10738_), .A2(new_n10470_), .B(new_n4018_), .ZN(new_n10746_));
  NOR2_X1    g10554(.A1(new_n10745_), .A2(new_n10746_), .ZN(new_n10747_));
  NAND2_X1   g10555(.A1(new_n10747_), .A2(new_n3760_), .ZN(new_n10748_));
  INV_X1     g10556(.I(new_n10748_), .ZN(new_n10749_));
  OAI21_X1   g10557(.A1(new_n10744_), .A2(new_n4018_), .B(new_n10749_), .ZN(new_n10750_));
  NAND2_X1   g10558(.A1(new_n10750_), .A2(new_n10743_), .ZN(new_n10751_));
  OAI22_X1   g10559(.A1(new_n10744_), .A2(new_n4018_), .B1(new_n10742_), .B2(new_n10736_), .ZN(new_n10752_));
  NAND2_X1   g10560(.A1(new_n10478_), .A2(\asqrt[41] ), .ZN(new_n10753_));
  NOR4_X1    g10561(.A1(new_n10614_), .A2(\asqrt[41] ), .A3(new_n10261_), .A4(new_n10478_), .ZN(new_n10754_));
  XOR2_X1    g10562(.A1(new_n10754_), .A2(new_n10753_), .Z(new_n10755_));
  NAND2_X1   g10563(.A1(new_n10755_), .A2(new_n3481_), .ZN(new_n10756_));
  AOI21_X1   g10564(.A1(new_n10752_), .A2(\asqrt[41] ), .B(new_n10756_), .ZN(new_n10757_));
  NOR2_X1    g10565(.A1(new_n10757_), .A2(new_n10751_), .ZN(new_n10758_));
  AOI22_X1   g10566(.A1(new_n10752_), .A2(\asqrt[41] ), .B1(new_n10750_), .B2(new_n10743_), .ZN(new_n10759_));
  NOR4_X1    g10567(.A1(new_n10614_), .A2(\asqrt[42] ), .A3(new_n10268_), .A4(new_n10273_), .ZN(new_n10760_));
  AOI21_X1   g10568(.A1(new_n10753_), .A2(new_n10477_), .B(new_n3481_), .ZN(new_n10761_));
  NOR2_X1    g10569(.A1(new_n10760_), .A2(new_n10761_), .ZN(new_n10762_));
  NAND2_X1   g10570(.A1(new_n10762_), .A2(new_n3208_), .ZN(new_n10763_));
  INV_X1     g10571(.I(new_n10763_), .ZN(new_n10764_));
  OAI21_X1   g10572(.A1(new_n10759_), .A2(new_n3481_), .B(new_n10764_), .ZN(new_n10765_));
  NAND2_X1   g10573(.A1(new_n10765_), .A2(new_n10758_), .ZN(new_n10766_));
  OAI22_X1   g10574(.A1(new_n10759_), .A2(new_n3481_), .B1(new_n10757_), .B2(new_n10751_), .ZN(new_n10767_));
  NAND2_X1   g10575(.A1(new_n10485_), .A2(\asqrt[43] ), .ZN(new_n10768_));
  NOR4_X1    g10576(.A1(new_n10614_), .A2(\asqrt[43] ), .A3(new_n10276_), .A4(new_n10485_), .ZN(new_n10769_));
  XOR2_X1    g10577(.A1(new_n10769_), .A2(new_n10768_), .Z(new_n10770_));
  NAND2_X1   g10578(.A1(new_n10770_), .A2(new_n2941_), .ZN(new_n10771_));
  AOI21_X1   g10579(.A1(new_n10767_), .A2(\asqrt[43] ), .B(new_n10771_), .ZN(new_n10772_));
  NOR2_X1    g10580(.A1(new_n10772_), .A2(new_n10766_), .ZN(new_n10773_));
  AOI22_X1   g10581(.A1(new_n10767_), .A2(\asqrt[43] ), .B1(new_n10765_), .B2(new_n10758_), .ZN(new_n10774_));
  NAND2_X1   g10582(.A1(new_n10288_), .A2(\asqrt[44] ), .ZN(new_n10775_));
  NOR4_X1    g10583(.A1(new_n10614_), .A2(\asqrt[44] ), .A3(new_n10283_), .A4(new_n10288_), .ZN(new_n10776_));
  XOR2_X1    g10584(.A1(new_n10776_), .A2(new_n10775_), .Z(new_n10777_));
  NAND2_X1   g10585(.A1(new_n10777_), .A2(new_n2728_), .ZN(new_n10778_));
  INV_X1     g10586(.I(new_n10778_), .ZN(new_n10779_));
  OAI21_X1   g10587(.A1(new_n10774_), .A2(new_n2941_), .B(new_n10779_), .ZN(new_n10780_));
  NAND2_X1   g10588(.A1(new_n10780_), .A2(new_n10773_), .ZN(new_n10781_));
  OAI22_X1   g10589(.A1(new_n10774_), .A2(new_n2941_), .B1(new_n10772_), .B2(new_n10766_), .ZN(new_n10782_));
  NOR4_X1    g10590(.A1(new_n10614_), .A2(\asqrt[45] ), .A3(new_n10291_), .A4(new_n10492_), .ZN(new_n10783_));
  AOI21_X1   g10591(.A1(new_n10775_), .A2(new_n10287_), .B(new_n2728_), .ZN(new_n10784_));
  NOR2_X1    g10592(.A1(new_n10783_), .A2(new_n10784_), .ZN(new_n10785_));
  NAND2_X1   g10593(.A1(new_n10785_), .A2(new_n2488_), .ZN(new_n10786_));
  AOI21_X1   g10594(.A1(new_n10782_), .A2(\asqrt[45] ), .B(new_n10786_), .ZN(new_n10787_));
  NOR2_X1    g10595(.A1(new_n10787_), .A2(new_n10781_), .ZN(new_n10788_));
  AOI22_X1   g10596(.A1(new_n10782_), .A2(\asqrt[45] ), .B1(new_n10780_), .B2(new_n10773_), .ZN(new_n10789_));
  NAND2_X1   g10597(.A1(new_n10303_), .A2(\asqrt[46] ), .ZN(new_n10790_));
  NOR4_X1    g10598(.A1(new_n10614_), .A2(\asqrt[46] ), .A3(new_n10298_), .A4(new_n10303_), .ZN(new_n10791_));
  XOR2_X1    g10599(.A1(new_n10791_), .A2(new_n10790_), .Z(new_n10792_));
  NAND2_X1   g10600(.A1(new_n10792_), .A2(new_n2253_), .ZN(new_n10793_));
  INV_X1     g10601(.I(new_n10793_), .ZN(new_n10794_));
  OAI21_X1   g10602(.A1(new_n10789_), .A2(new_n2488_), .B(new_n10794_), .ZN(new_n10795_));
  NAND2_X1   g10603(.A1(new_n10795_), .A2(new_n10788_), .ZN(new_n10796_));
  OAI22_X1   g10604(.A1(new_n10789_), .A2(new_n2488_), .B1(new_n10787_), .B2(new_n10781_), .ZN(new_n10797_));
  NOR4_X1    g10605(.A1(new_n10614_), .A2(\asqrt[47] ), .A3(new_n10306_), .A4(new_n10499_), .ZN(new_n10798_));
  AOI21_X1   g10606(.A1(new_n10790_), .A2(new_n10302_), .B(new_n2253_), .ZN(new_n10799_));
  NOR2_X1    g10607(.A1(new_n10798_), .A2(new_n10799_), .ZN(new_n10800_));
  NAND2_X1   g10608(.A1(new_n10800_), .A2(new_n2046_), .ZN(new_n10801_));
  AOI21_X1   g10609(.A1(new_n10797_), .A2(\asqrt[47] ), .B(new_n10801_), .ZN(new_n10802_));
  NOR2_X1    g10610(.A1(new_n10802_), .A2(new_n10796_), .ZN(new_n10803_));
  AOI22_X1   g10611(.A1(new_n10797_), .A2(\asqrt[47] ), .B1(new_n10795_), .B2(new_n10788_), .ZN(new_n10804_));
  NAND2_X1   g10612(.A1(new_n10318_), .A2(\asqrt[48] ), .ZN(new_n10805_));
  NOR4_X1    g10613(.A1(new_n10614_), .A2(\asqrt[48] ), .A3(new_n10313_), .A4(new_n10318_), .ZN(new_n10806_));
  XOR2_X1    g10614(.A1(new_n10806_), .A2(new_n10805_), .Z(new_n10807_));
  NAND2_X1   g10615(.A1(new_n10807_), .A2(new_n1854_), .ZN(new_n10808_));
  INV_X1     g10616(.I(new_n10808_), .ZN(new_n10809_));
  OAI21_X1   g10617(.A1(new_n10804_), .A2(new_n2046_), .B(new_n10809_), .ZN(new_n10810_));
  NAND2_X1   g10618(.A1(new_n10810_), .A2(new_n10803_), .ZN(new_n10811_));
  OAI22_X1   g10619(.A1(new_n10804_), .A2(new_n2046_), .B1(new_n10802_), .B2(new_n10796_), .ZN(new_n10812_));
  NAND2_X1   g10620(.A1(new_n10506_), .A2(\asqrt[49] ), .ZN(new_n10813_));
  NOR4_X1    g10621(.A1(new_n10614_), .A2(\asqrt[49] ), .A3(new_n10321_), .A4(new_n10506_), .ZN(new_n10814_));
  XOR2_X1    g10622(.A1(new_n10814_), .A2(new_n10813_), .Z(new_n10815_));
  NAND2_X1   g10623(.A1(new_n10815_), .A2(new_n1595_), .ZN(new_n10816_));
  AOI21_X1   g10624(.A1(new_n10812_), .A2(\asqrt[49] ), .B(new_n10816_), .ZN(new_n10817_));
  NOR2_X1    g10625(.A1(new_n10817_), .A2(new_n10811_), .ZN(new_n10818_));
  AOI22_X1   g10626(.A1(new_n10812_), .A2(\asqrt[49] ), .B1(new_n10810_), .B2(new_n10803_), .ZN(new_n10819_));
  NOR4_X1    g10627(.A1(new_n10614_), .A2(\asqrt[50] ), .A3(new_n10328_), .A4(new_n10333_), .ZN(new_n10820_));
  AOI21_X1   g10628(.A1(new_n10813_), .A2(new_n10505_), .B(new_n1595_), .ZN(new_n10821_));
  NOR2_X1    g10629(.A1(new_n10820_), .A2(new_n10821_), .ZN(new_n10822_));
  NAND2_X1   g10630(.A1(new_n10822_), .A2(new_n1436_), .ZN(new_n10823_));
  INV_X1     g10631(.I(new_n10823_), .ZN(new_n10824_));
  OAI21_X1   g10632(.A1(new_n10819_), .A2(new_n1595_), .B(new_n10824_), .ZN(new_n10825_));
  NAND2_X1   g10633(.A1(new_n10825_), .A2(new_n10818_), .ZN(new_n10826_));
  OAI22_X1   g10634(.A1(new_n10819_), .A2(new_n1595_), .B1(new_n10817_), .B2(new_n10811_), .ZN(new_n10827_));
  NAND2_X1   g10635(.A1(new_n10513_), .A2(\asqrt[51] ), .ZN(new_n10828_));
  NOR4_X1    g10636(.A1(new_n10614_), .A2(\asqrt[51] ), .A3(new_n10336_), .A4(new_n10513_), .ZN(new_n10829_));
  XOR2_X1    g10637(.A1(new_n10829_), .A2(new_n10828_), .Z(new_n10830_));
  NAND2_X1   g10638(.A1(new_n10830_), .A2(new_n1260_), .ZN(new_n10831_));
  AOI21_X1   g10639(.A1(new_n10827_), .A2(\asqrt[51] ), .B(new_n10831_), .ZN(new_n10832_));
  NOR2_X1    g10640(.A1(new_n10832_), .A2(new_n10826_), .ZN(new_n10833_));
  AOI22_X1   g10641(.A1(new_n10827_), .A2(\asqrt[51] ), .B1(new_n10825_), .B2(new_n10818_), .ZN(new_n10834_));
  NOR4_X1    g10642(.A1(new_n10614_), .A2(\asqrt[52] ), .A3(new_n10343_), .A4(new_n10348_), .ZN(new_n10835_));
  AOI21_X1   g10643(.A1(new_n10828_), .A2(new_n10512_), .B(new_n1260_), .ZN(new_n10836_));
  NOR2_X1    g10644(.A1(new_n10835_), .A2(new_n10836_), .ZN(new_n10837_));
  NAND2_X1   g10645(.A1(new_n10837_), .A2(new_n1096_), .ZN(new_n10838_));
  INV_X1     g10646(.I(new_n10838_), .ZN(new_n10839_));
  OAI21_X1   g10647(.A1(new_n10834_), .A2(new_n1260_), .B(new_n10839_), .ZN(new_n10840_));
  NAND2_X1   g10648(.A1(new_n10840_), .A2(new_n10833_), .ZN(new_n10841_));
  OAI22_X1   g10649(.A1(new_n10834_), .A2(new_n1260_), .B1(new_n10832_), .B2(new_n10826_), .ZN(new_n10842_));
  NOR4_X1    g10650(.A1(new_n10614_), .A2(\asqrt[53] ), .A3(new_n10351_), .A4(new_n10520_), .ZN(new_n10843_));
  XOR2_X1    g10651(.A1(new_n10843_), .A2(new_n10541_), .Z(new_n10844_));
  NAND2_X1   g10652(.A1(new_n10844_), .A2(new_n970_), .ZN(new_n10845_));
  AOI21_X1   g10653(.A1(new_n10842_), .A2(\asqrt[53] ), .B(new_n10845_), .ZN(new_n10846_));
  NOR2_X1    g10654(.A1(new_n10846_), .A2(new_n10841_), .ZN(new_n10847_));
  AOI22_X1   g10655(.A1(new_n10842_), .A2(\asqrt[53] ), .B1(new_n10840_), .B2(new_n10833_), .ZN(new_n10848_));
  NOR4_X1    g10656(.A1(new_n10614_), .A2(\asqrt[54] ), .A3(new_n10358_), .A4(new_n10363_), .ZN(new_n10849_));
  XNOR2_X1   g10657(.A1(new_n10849_), .A2(new_n10542_), .ZN(new_n10850_));
  NAND2_X1   g10658(.A1(new_n10850_), .A2(new_n825_), .ZN(new_n10851_));
  INV_X1     g10659(.I(new_n10851_), .ZN(new_n10852_));
  OAI21_X1   g10660(.A1(new_n10848_), .A2(new_n970_), .B(new_n10852_), .ZN(new_n10853_));
  NAND2_X1   g10661(.A1(new_n10853_), .A2(new_n10847_), .ZN(new_n10854_));
  OAI22_X1   g10662(.A1(new_n10848_), .A2(new_n970_), .B1(new_n10846_), .B2(new_n10841_), .ZN(new_n10855_));
  NOR4_X1    g10663(.A1(new_n10614_), .A2(\asqrt[55] ), .A3(new_n10365_), .A4(new_n10527_), .ZN(new_n10856_));
  XOR2_X1    g10664(.A1(new_n10856_), .A2(new_n10543_), .Z(new_n10857_));
  NAND2_X1   g10665(.A1(new_n10857_), .A2(new_n724_), .ZN(new_n10858_));
  AOI21_X1   g10666(.A1(new_n10855_), .A2(\asqrt[55] ), .B(new_n10858_), .ZN(new_n10859_));
  NOR2_X1    g10667(.A1(new_n10859_), .A2(new_n10854_), .ZN(new_n10860_));
  AOI22_X1   g10668(.A1(new_n10855_), .A2(\asqrt[55] ), .B1(new_n10853_), .B2(new_n10847_), .ZN(new_n10861_));
  NOR4_X1    g10669(.A1(new_n10614_), .A2(\asqrt[56] ), .A3(new_n10371_), .A4(new_n10376_), .ZN(new_n10862_));
  XOR2_X1    g10670(.A1(new_n10862_), .A2(new_n10401_), .Z(new_n10863_));
  NAND2_X1   g10671(.A1(new_n10863_), .A2(new_n587_), .ZN(new_n10864_));
  INV_X1     g10672(.I(new_n10864_), .ZN(new_n10865_));
  OAI21_X1   g10673(.A1(new_n10861_), .A2(new_n724_), .B(new_n10865_), .ZN(new_n10866_));
  NAND2_X1   g10674(.A1(new_n10866_), .A2(new_n10860_), .ZN(new_n10867_));
  OAI22_X1   g10675(.A1(new_n10861_), .A2(new_n724_), .B1(new_n10859_), .B2(new_n10854_), .ZN(new_n10868_));
  NOR4_X1    g10676(.A1(new_n10614_), .A2(\asqrt[57] ), .A3(new_n10378_), .A4(new_n10534_), .ZN(new_n10869_));
  XOR2_X1    g10677(.A1(new_n10869_), .A2(new_n10545_), .Z(new_n10870_));
  NAND2_X1   g10678(.A1(new_n10870_), .A2(new_n504_), .ZN(new_n10871_));
  AOI21_X1   g10679(.A1(new_n10868_), .A2(\asqrt[57] ), .B(new_n10871_), .ZN(new_n10872_));
  NOR2_X1    g10680(.A1(new_n10872_), .A2(new_n10867_), .ZN(new_n10873_));
  AOI22_X1   g10681(.A1(new_n10868_), .A2(\asqrt[57] ), .B1(new_n10866_), .B2(new_n10860_), .ZN(new_n10874_));
  NOR4_X1    g10682(.A1(new_n10614_), .A2(\asqrt[58] ), .A3(new_n10384_), .A4(new_n10389_), .ZN(new_n10875_));
  XOR2_X1    g10683(.A1(new_n10875_), .A2(new_n10403_), .Z(new_n10876_));
  NAND2_X1   g10684(.A1(new_n10876_), .A2(new_n376_), .ZN(new_n10877_));
  INV_X1     g10685(.I(new_n10877_), .ZN(new_n10878_));
  OAI21_X1   g10686(.A1(new_n10874_), .A2(new_n504_), .B(new_n10878_), .ZN(new_n10879_));
  NAND2_X1   g10687(.A1(new_n10879_), .A2(new_n10873_), .ZN(new_n10880_));
  OAI22_X1   g10688(.A1(new_n10874_), .A2(new_n504_), .B1(new_n10872_), .B2(new_n10867_), .ZN(new_n10881_));
  NOR4_X1    g10689(.A1(new_n10614_), .A2(\asqrt[59] ), .A3(new_n10391_), .A4(new_n10549_), .ZN(new_n10882_));
  XOR2_X1    g10690(.A1(new_n10882_), .A2(new_n10547_), .Z(new_n10883_));
  NAND2_X1   g10691(.A1(new_n10883_), .A2(new_n275_), .ZN(new_n10884_));
  AOI21_X1   g10692(.A1(new_n10881_), .A2(\asqrt[59] ), .B(new_n10884_), .ZN(new_n10885_));
  NOR2_X1    g10693(.A1(new_n10885_), .A2(new_n10880_), .ZN(new_n10886_));
  AOI22_X1   g10694(.A1(new_n10881_), .A2(\asqrt[59] ), .B1(new_n10879_), .B2(new_n10873_), .ZN(new_n10887_));
  OAI22_X1   g10695(.A1(new_n10887_), .A2(new_n275_), .B1(new_n10885_), .B2(new_n10880_), .ZN(new_n10888_));
  NOR4_X1    g10696(.A1(new_n10614_), .A2(\asqrt[60] ), .A3(new_n10397_), .A4(new_n10570_), .ZN(new_n10889_));
  XOR2_X1    g10697(.A1(new_n10889_), .A2(new_n10405_), .Z(new_n10890_));
  NAND2_X1   g10698(.A1(new_n10890_), .A2(new_n229_), .ZN(new_n10891_));
  INV_X1     g10699(.I(new_n10891_), .ZN(new_n10892_));
  OAI21_X1   g10700(.A1(new_n10887_), .A2(new_n275_), .B(new_n10892_), .ZN(new_n10893_));
  AOI22_X1   g10701(.A1(new_n10888_), .A2(\asqrt[61] ), .B1(new_n10893_), .B2(new_n10886_), .ZN(new_n10894_));
  NOR2_X1    g10702(.A1(new_n10894_), .A2(new_n196_), .ZN(new_n10895_));
  INV_X1     g10703(.I(new_n10591_), .ZN(new_n10896_));
  AOI21_X1   g10704(.A1(new_n10605_), .A2(new_n10896_), .B(new_n10593_), .ZN(new_n10897_));
  NOR3_X1    g10705(.A1(new_n10590_), .A2(new_n10583_), .A3(new_n10588_), .ZN(new_n10898_));
  NOR2_X1    g10706(.A1(new_n10898_), .A2(new_n10897_), .ZN(new_n10899_));
  NOR3_X1    g10707(.A1(new_n10628_), .A2(new_n9616_), .A3(\asqrt[23] ), .ZN(new_n10900_));
  AOI21_X1   g10708(.A1(new_n10622_), .A2(new_n9615_), .B(new_n10614_), .ZN(new_n10901_));
  NOR4_X1    g10709(.A1(new_n10901_), .A2(new_n10900_), .A3(\asqrt[25] ), .A4(new_n10612_), .ZN(new_n10902_));
  NOR2_X1    g10710(.A1(new_n10902_), .A2(new_n10899_), .ZN(new_n10903_));
  NOR3_X1    g10711(.A1(new_n10898_), .A2(new_n10897_), .A3(new_n10612_), .ZN(new_n10904_));
  NOR3_X1    g10712(.A1(new_n10614_), .A2(new_n10102_), .A3(new_n10639_), .ZN(new_n10905_));
  AOI21_X1   g10713(.A1(\asqrt[23] ), .A2(new_n10637_), .B(new_n10103_), .ZN(new_n10906_));
  NOR3_X1    g10714(.A1(new_n10906_), .A2(new_n10905_), .A3(\asqrt[26] ), .ZN(new_n10907_));
  OAI21_X1   g10715(.A1(new_n10904_), .A2(new_n9672_), .B(new_n10907_), .ZN(new_n10908_));
  NAND2_X1   g10716(.A1(new_n10903_), .A2(new_n10908_), .ZN(new_n10909_));
  OAI22_X1   g10717(.A1(new_n10902_), .A2(new_n10899_), .B1(new_n9672_), .B2(new_n10904_), .ZN(new_n10910_));
  INV_X1     g10718(.I(new_n10648_), .ZN(new_n10911_));
  AOI21_X1   g10719(.A1(new_n10910_), .A2(\asqrt[26] ), .B(new_n10911_), .ZN(new_n10912_));
  NOR2_X1    g10720(.A1(new_n10912_), .A2(new_n10909_), .ZN(new_n10913_));
  AOI22_X1   g10721(.A1(new_n10910_), .A2(\asqrt[26] ), .B1(new_n10903_), .B2(new_n10908_), .ZN(new_n10914_));
  INV_X1     g10722(.I(new_n10655_), .ZN(new_n10915_));
  OAI21_X1   g10723(.A1(new_n10914_), .A2(new_n8763_), .B(new_n10915_), .ZN(new_n10916_));
  NAND2_X1   g10724(.A1(new_n10916_), .A2(new_n10913_), .ZN(new_n10917_));
  OAI22_X1   g10725(.A1(new_n10914_), .A2(new_n8763_), .B1(new_n10912_), .B2(new_n10909_), .ZN(new_n10918_));
  AOI21_X1   g10726(.A1(new_n10918_), .A2(\asqrt[28] ), .B(new_n10662_), .ZN(new_n10919_));
  NOR2_X1    g10727(.A1(new_n10919_), .A2(new_n10917_), .ZN(new_n10920_));
  AOI22_X1   g10728(.A1(new_n10918_), .A2(\asqrt[28] ), .B1(new_n10916_), .B2(new_n10913_), .ZN(new_n10921_));
  INV_X1     g10729(.I(new_n10669_), .ZN(new_n10922_));
  OAI21_X1   g10730(.A1(new_n10921_), .A2(new_n7931_), .B(new_n10922_), .ZN(new_n10923_));
  NAND2_X1   g10731(.A1(new_n10923_), .A2(new_n10920_), .ZN(new_n10924_));
  OAI22_X1   g10732(.A1(new_n10921_), .A2(new_n7931_), .B1(new_n10919_), .B2(new_n10917_), .ZN(new_n10925_));
  AOI21_X1   g10733(.A1(new_n10925_), .A2(\asqrt[30] ), .B(new_n10675_), .ZN(new_n10926_));
  NOR2_X1    g10734(.A1(new_n10926_), .A2(new_n10924_), .ZN(new_n10927_));
  AOI22_X1   g10735(.A1(new_n10925_), .A2(\asqrt[30] ), .B1(new_n10923_), .B2(new_n10920_), .ZN(new_n10928_));
  INV_X1     g10736(.I(new_n10682_), .ZN(new_n10929_));
  OAI21_X1   g10737(.A1(new_n10928_), .A2(new_n7110_), .B(new_n10929_), .ZN(new_n10930_));
  NAND2_X1   g10738(.A1(new_n10930_), .A2(new_n10927_), .ZN(new_n10931_));
  OAI22_X1   g10739(.A1(new_n10928_), .A2(new_n7110_), .B1(new_n10926_), .B2(new_n10924_), .ZN(new_n10932_));
  AOI21_X1   g10740(.A1(new_n10932_), .A2(\asqrt[32] ), .B(new_n10688_), .ZN(new_n10933_));
  NOR2_X1    g10741(.A1(new_n10933_), .A2(new_n10931_), .ZN(new_n10934_));
  AOI22_X1   g10742(.A1(new_n10932_), .A2(\asqrt[32] ), .B1(new_n10930_), .B2(new_n10927_), .ZN(new_n10935_));
  INV_X1     g10743(.I(new_n10696_), .ZN(new_n10936_));
  OAI21_X1   g10744(.A1(new_n10935_), .A2(new_n6365_), .B(new_n10936_), .ZN(new_n10937_));
  NAND2_X1   g10745(.A1(new_n10937_), .A2(new_n10934_), .ZN(new_n10938_));
  OAI22_X1   g10746(.A1(new_n10935_), .A2(new_n6365_), .B1(new_n10933_), .B2(new_n10931_), .ZN(new_n10939_));
  AOI21_X1   g10747(.A1(new_n10939_), .A2(\asqrt[34] ), .B(new_n10703_), .ZN(new_n10940_));
  NOR2_X1    g10748(.A1(new_n10940_), .A2(new_n10938_), .ZN(new_n10941_));
  AOI22_X1   g10749(.A1(new_n10939_), .A2(\asqrt[34] ), .B1(new_n10937_), .B2(new_n10934_), .ZN(new_n10942_));
  INV_X1     g10750(.I(new_n10711_), .ZN(new_n10943_));
  OAI21_X1   g10751(.A1(new_n10942_), .A2(new_n5626_), .B(new_n10943_), .ZN(new_n10944_));
  NAND2_X1   g10752(.A1(new_n10944_), .A2(new_n10941_), .ZN(new_n10945_));
  OAI22_X1   g10753(.A1(new_n10942_), .A2(new_n5626_), .B1(new_n10940_), .B2(new_n10938_), .ZN(new_n10946_));
  AOI21_X1   g10754(.A1(new_n10946_), .A2(\asqrt[36] ), .B(new_n10718_), .ZN(new_n10947_));
  NOR2_X1    g10755(.A1(new_n10947_), .A2(new_n10945_), .ZN(new_n10948_));
  AOI22_X1   g10756(.A1(new_n10946_), .A2(\asqrt[36] ), .B1(new_n10944_), .B2(new_n10941_), .ZN(new_n10949_));
  INV_X1     g10757(.I(new_n10726_), .ZN(new_n10950_));
  OAI21_X1   g10758(.A1(new_n10949_), .A2(new_n4973_), .B(new_n10950_), .ZN(new_n10951_));
  NAND2_X1   g10759(.A1(new_n10951_), .A2(new_n10948_), .ZN(new_n10952_));
  OAI22_X1   g10760(.A1(new_n10949_), .A2(new_n4973_), .B1(new_n10947_), .B2(new_n10945_), .ZN(new_n10953_));
  AOI21_X1   g10761(.A1(new_n10953_), .A2(\asqrt[38] ), .B(new_n10733_), .ZN(new_n10954_));
  NOR2_X1    g10762(.A1(new_n10954_), .A2(new_n10952_), .ZN(new_n10955_));
  AOI22_X1   g10763(.A1(new_n10953_), .A2(\asqrt[38] ), .B1(new_n10951_), .B2(new_n10948_), .ZN(new_n10956_));
  INV_X1     g10764(.I(new_n10741_), .ZN(new_n10957_));
  OAI21_X1   g10765(.A1(new_n10956_), .A2(new_n4330_), .B(new_n10957_), .ZN(new_n10958_));
  NAND2_X1   g10766(.A1(new_n10958_), .A2(new_n10955_), .ZN(new_n10959_));
  OAI22_X1   g10767(.A1(new_n10956_), .A2(new_n4330_), .B1(new_n10954_), .B2(new_n10952_), .ZN(new_n10960_));
  AOI21_X1   g10768(.A1(new_n10960_), .A2(\asqrt[40] ), .B(new_n10748_), .ZN(new_n10961_));
  NOR2_X1    g10769(.A1(new_n10961_), .A2(new_n10959_), .ZN(new_n10962_));
  AOI22_X1   g10770(.A1(new_n10960_), .A2(\asqrt[40] ), .B1(new_n10958_), .B2(new_n10955_), .ZN(new_n10963_));
  INV_X1     g10771(.I(new_n10756_), .ZN(new_n10964_));
  OAI21_X1   g10772(.A1(new_n10963_), .A2(new_n3760_), .B(new_n10964_), .ZN(new_n10965_));
  NAND2_X1   g10773(.A1(new_n10965_), .A2(new_n10962_), .ZN(new_n10966_));
  OAI22_X1   g10774(.A1(new_n10963_), .A2(new_n3760_), .B1(new_n10961_), .B2(new_n10959_), .ZN(new_n10967_));
  AOI21_X1   g10775(.A1(new_n10967_), .A2(\asqrt[42] ), .B(new_n10763_), .ZN(new_n10968_));
  NOR2_X1    g10776(.A1(new_n10968_), .A2(new_n10966_), .ZN(new_n10969_));
  AOI22_X1   g10777(.A1(new_n10967_), .A2(\asqrt[42] ), .B1(new_n10965_), .B2(new_n10962_), .ZN(new_n10970_));
  INV_X1     g10778(.I(new_n10771_), .ZN(new_n10971_));
  OAI21_X1   g10779(.A1(new_n10970_), .A2(new_n3208_), .B(new_n10971_), .ZN(new_n10972_));
  NAND2_X1   g10780(.A1(new_n10972_), .A2(new_n10969_), .ZN(new_n10973_));
  OAI22_X1   g10781(.A1(new_n10970_), .A2(new_n3208_), .B1(new_n10968_), .B2(new_n10966_), .ZN(new_n10974_));
  AOI21_X1   g10782(.A1(new_n10974_), .A2(\asqrt[44] ), .B(new_n10778_), .ZN(new_n10975_));
  NOR2_X1    g10783(.A1(new_n10975_), .A2(new_n10973_), .ZN(new_n10976_));
  AOI22_X1   g10784(.A1(new_n10974_), .A2(\asqrt[44] ), .B1(new_n10972_), .B2(new_n10969_), .ZN(new_n10977_));
  INV_X1     g10785(.I(new_n10786_), .ZN(new_n10978_));
  OAI21_X1   g10786(.A1(new_n10977_), .A2(new_n2728_), .B(new_n10978_), .ZN(new_n10979_));
  NAND2_X1   g10787(.A1(new_n10979_), .A2(new_n10976_), .ZN(new_n10980_));
  OAI22_X1   g10788(.A1(new_n10977_), .A2(new_n2728_), .B1(new_n10975_), .B2(new_n10973_), .ZN(new_n10981_));
  AOI21_X1   g10789(.A1(new_n10981_), .A2(\asqrt[46] ), .B(new_n10793_), .ZN(new_n10982_));
  NOR2_X1    g10790(.A1(new_n10982_), .A2(new_n10980_), .ZN(new_n10983_));
  AOI22_X1   g10791(.A1(new_n10981_), .A2(\asqrt[46] ), .B1(new_n10979_), .B2(new_n10976_), .ZN(new_n10984_));
  INV_X1     g10792(.I(new_n10801_), .ZN(new_n10985_));
  OAI21_X1   g10793(.A1(new_n10984_), .A2(new_n2253_), .B(new_n10985_), .ZN(new_n10986_));
  NAND2_X1   g10794(.A1(new_n10986_), .A2(new_n10983_), .ZN(new_n10987_));
  OAI22_X1   g10795(.A1(new_n10984_), .A2(new_n2253_), .B1(new_n10982_), .B2(new_n10980_), .ZN(new_n10988_));
  AOI21_X1   g10796(.A1(new_n10988_), .A2(\asqrt[48] ), .B(new_n10808_), .ZN(new_n10989_));
  NOR2_X1    g10797(.A1(new_n10989_), .A2(new_n10987_), .ZN(new_n10990_));
  AOI22_X1   g10798(.A1(new_n10988_), .A2(\asqrt[48] ), .B1(new_n10986_), .B2(new_n10983_), .ZN(new_n10991_));
  INV_X1     g10799(.I(new_n10816_), .ZN(new_n10992_));
  OAI21_X1   g10800(.A1(new_n10991_), .A2(new_n1854_), .B(new_n10992_), .ZN(new_n10993_));
  NAND2_X1   g10801(.A1(new_n10993_), .A2(new_n10990_), .ZN(new_n10994_));
  OAI22_X1   g10802(.A1(new_n10991_), .A2(new_n1854_), .B1(new_n10989_), .B2(new_n10987_), .ZN(new_n10995_));
  AOI21_X1   g10803(.A1(new_n10995_), .A2(\asqrt[50] ), .B(new_n10823_), .ZN(new_n10996_));
  NOR2_X1    g10804(.A1(new_n10996_), .A2(new_n10994_), .ZN(new_n10997_));
  AOI22_X1   g10805(.A1(new_n10995_), .A2(\asqrt[50] ), .B1(new_n10993_), .B2(new_n10990_), .ZN(new_n10998_));
  INV_X1     g10806(.I(new_n10831_), .ZN(new_n10999_));
  OAI21_X1   g10807(.A1(new_n10998_), .A2(new_n1436_), .B(new_n10999_), .ZN(new_n11000_));
  NAND2_X1   g10808(.A1(new_n11000_), .A2(new_n10997_), .ZN(new_n11001_));
  OAI22_X1   g10809(.A1(new_n10998_), .A2(new_n1436_), .B1(new_n10996_), .B2(new_n10994_), .ZN(new_n11002_));
  AOI21_X1   g10810(.A1(new_n11002_), .A2(\asqrt[52] ), .B(new_n10838_), .ZN(new_n11003_));
  NOR2_X1    g10811(.A1(new_n11003_), .A2(new_n11001_), .ZN(new_n11004_));
  AOI22_X1   g10812(.A1(new_n11002_), .A2(\asqrt[52] ), .B1(new_n11000_), .B2(new_n10997_), .ZN(new_n11005_));
  INV_X1     g10813(.I(new_n10845_), .ZN(new_n11006_));
  OAI21_X1   g10814(.A1(new_n11005_), .A2(new_n1096_), .B(new_n11006_), .ZN(new_n11007_));
  NAND2_X1   g10815(.A1(new_n11007_), .A2(new_n11004_), .ZN(new_n11008_));
  OAI22_X1   g10816(.A1(new_n11005_), .A2(new_n1096_), .B1(new_n11003_), .B2(new_n11001_), .ZN(new_n11009_));
  AOI21_X1   g10817(.A1(new_n11009_), .A2(\asqrt[54] ), .B(new_n10851_), .ZN(new_n11010_));
  NOR2_X1    g10818(.A1(new_n11010_), .A2(new_n11008_), .ZN(new_n11011_));
  AOI22_X1   g10819(.A1(new_n11009_), .A2(\asqrt[54] ), .B1(new_n11007_), .B2(new_n11004_), .ZN(new_n11012_));
  INV_X1     g10820(.I(new_n10858_), .ZN(new_n11013_));
  OAI21_X1   g10821(.A1(new_n11012_), .A2(new_n825_), .B(new_n11013_), .ZN(new_n11014_));
  NAND2_X1   g10822(.A1(new_n11014_), .A2(new_n11011_), .ZN(new_n11015_));
  OAI22_X1   g10823(.A1(new_n11012_), .A2(new_n825_), .B1(new_n11010_), .B2(new_n11008_), .ZN(new_n11016_));
  AOI21_X1   g10824(.A1(new_n11016_), .A2(\asqrt[56] ), .B(new_n10864_), .ZN(new_n11017_));
  NOR2_X1    g10825(.A1(new_n11017_), .A2(new_n11015_), .ZN(new_n11018_));
  AOI22_X1   g10826(.A1(new_n11016_), .A2(\asqrt[56] ), .B1(new_n11014_), .B2(new_n11011_), .ZN(new_n11019_));
  INV_X1     g10827(.I(new_n10871_), .ZN(new_n11020_));
  OAI21_X1   g10828(.A1(new_n11019_), .A2(new_n587_), .B(new_n11020_), .ZN(new_n11021_));
  NAND2_X1   g10829(.A1(new_n11021_), .A2(new_n11018_), .ZN(new_n11022_));
  OAI22_X1   g10830(.A1(new_n11019_), .A2(new_n587_), .B1(new_n11017_), .B2(new_n11015_), .ZN(new_n11023_));
  AOI21_X1   g10831(.A1(new_n11023_), .A2(\asqrt[58] ), .B(new_n10877_), .ZN(new_n11024_));
  NOR2_X1    g10832(.A1(new_n11024_), .A2(new_n11022_), .ZN(new_n11025_));
  AOI22_X1   g10833(.A1(new_n11023_), .A2(\asqrt[58] ), .B1(new_n11021_), .B2(new_n11018_), .ZN(new_n11026_));
  INV_X1     g10834(.I(new_n10884_), .ZN(new_n11027_));
  OAI21_X1   g10835(.A1(new_n11026_), .A2(new_n376_), .B(new_n11027_), .ZN(new_n11028_));
  NAND2_X1   g10836(.A1(new_n11028_), .A2(new_n11025_), .ZN(new_n11029_));
  OAI22_X1   g10837(.A1(new_n11026_), .A2(new_n376_), .B1(new_n11024_), .B2(new_n11022_), .ZN(new_n11030_));
  AOI22_X1   g10838(.A1(new_n11030_), .A2(\asqrt[60] ), .B1(new_n11028_), .B2(new_n11025_), .ZN(new_n11031_));
  AOI21_X1   g10839(.A1(new_n11030_), .A2(\asqrt[60] ), .B(new_n10891_), .ZN(new_n11032_));
  OAI22_X1   g10840(.A1(new_n11031_), .A2(new_n229_), .B1(new_n11032_), .B2(new_n11029_), .ZN(new_n11033_));
  NOR2_X1    g10841(.A1(new_n11033_), .A2(\asqrt[62] ), .ZN(new_n11034_));
  NAND3_X1   g10842(.A1(new_n10608_), .A2(new_n10412_), .A3(new_n10576_), .ZN(new_n11035_));
  NOR2_X1    g10843(.A1(new_n10617_), .A2(new_n196_), .ZN(new_n11036_));
  INV_X1     g10844(.I(new_n10602_), .ZN(new_n11037_));
  NAND3_X1   g10845(.A1(\asqrt[23] ), .A2(new_n11036_), .A3(new_n11037_), .ZN(new_n11038_));
  OAI21_X1   g10846(.A1(new_n10573_), .A2(\asqrt[62] ), .B(new_n10414_), .ZN(new_n11039_));
  OAI21_X1   g10847(.A1(\asqrt[23] ), .A2(new_n11039_), .B(new_n11036_), .ZN(new_n11040_));
  NAND2_X1   g10848(.A1(new_n11040_), .A2(new_n11038_), .ZN(new_n11041_));
  INV_X1     g10849(.I(new_n11041_), .ZN(new_n11042_));
  NOR2_X1    g10850(.A1(new_n10581_), .A2(new_n196_), .ZN(new_n11043_));
  INV_X1     g10851(.I(new_n11043_), .ZN(new_n11044_));
  NAND2_X1   g10852(.A1(new_n10868_), .A2(\asqrt[57] ), .ZN(new_n11045_));
  AOI21_X1   g10853(.A1(new_n11045_), .A2(new_n10867_), .B(new_n504_), .ZN(new_n11046_));
  OAI21_X1   g10854(.A1(new_n10873_), .A2(new_n11046_), .B(\asqrt[59] ), .ZN(new_n11047_));
  AOI21_X1   g10855(.A1(new_n10880_), .A2(new_n11047_), .B(new_n275_), .ZN(new_n11048_));
  OAI21_X1   g10856(.A1(new_n10886_), .A2(new_n11048_), .B(\asqrt[61] ), .ZN(new_n11049_));
  NOR2_X1    g10857(.A1(new_n10582_), .A2(\asqrt[62] ), .ZN(new_n11050_));
  INV_X1     g10858(.I(new_n11050_), .ZN(new_n11051_));
  NAND3_X1   g10859(.A1(new_n10893_), .A2(new_n10886_), .A3(new_n11051_), .ZN(new_n11052_));
  OAI21_X1   g10860(.A1(new_n11052_), .A2(new_n11049_), .B(new_n11044_), .ZN(new_n11053_));
  NAND3_X1   g10861(.A1(new_n10614_), .A2(new_n10569_), .A3(new_n10618_), .ZN(new_n11054_));
  AOI21_X1   g10862(.A1(new_n11054_), .A2(new_n10561_), .B(\asqrt[63] ), .ZN(new_n11055_));
  INV_X1     g10863(.I(new_n11055_), .ZN(new_n11056_));
  OAI21_X1   g10864(.A1(new_n11053_), .A2(new_n11056_), .B(new_n11042_), .ZN(new_n11057_));
  NOR4_X1    g10865(.A1(new_n11033_), .A2(\asqrt[62] ), .A3(new_n11041_), .A4(new_n10581_), .ZN(new_n11058_));
  NAND2_X1   g10866(.A1(new_n10596_), .A2(new_n10569_), .ZN(new_n11059_));
  XOR2_X1    g10867(.A1(new_n10596_), .A2(\asqrt[63] ), .Z(new_n11060_));
  AOI21_X1   g10868(.A1(\asqrt[23] ), .A2(new_n11059_), .B(new_n11060_), .ZN(new_n11061_));
  NAND2_X1   g10869(.A1(new_n11058_), .A2(new_n11061_), .ZN(new_n11062_));
  NOR3_X1    g10870(.A1(new_n11062_), .A2(new_n11035_), .A3(new_n11057_), .ZN(\asqrt[22] ));
  NAND4_X1   g10871(.A1(\asqrt[22] ), .A2(new_n10582_), .A3(new_n10895_), .A4(new_n11034_), .ZN(new_n11064_));
  OAI21_X1   g10872(.A1(new_n11033_), .A2(\asqrt[62] ), .B(new_n10581_), .ZN(new_n11065_));
  OAI21_X1   g10873(.A1(\asqrt[22] ), .A2(new_n11065_), .B(new_n10895_), .ZN(new_n11066_));
  NAND2_X1   g10874(.A1(new_n11064_), .A2(new_n11066_), .ZN(new_n11067_));
  INV_X1     g10875(.I(new_n11067_), .ZN(new_n11068_));
  NAND2_X1   g10876(.A1(new_n11023_), .A2(\asqrt[58] ), .ZN(new_n11069_));
  AOI21_X1   g10877(.A1(new_n11069_), .A2(new_n11022_), .B(new_n376_), .ZN(new_n11070_));
  OAI21_X1   g10878(.A1(new_n11025_), .A2(new_n11070_), .B(\asqrt[60] ), .ZN(new_n11071_));
  AOI21_X1   g10879(.A1(new_n11029_), .A2(new_n11071_), .B(new_n229_), .ZN(new_n11072_));
  NOR3_X1    g10880(.A1(new_n10888_), .A2(\asqrt[61] ), .A3(new_n10890_), .ZN(new_n11073_));
  NAND2_X1   g10881(.A1(\asqrt[22] ), .A2(new_n11073_), .ZN(new_n11074_));
  XOR2_X1    g10882(.A1(new_n11074_), .A2(new_n11072_), .Z(new_n11075_));
  NOR2_X1    g10883(.A1(new_n11075_), .A2(new_n196_), .ZN(new_n11076_));
  INV_X1     g10884(.I(new_n11076_), .ZN(new_n11077_));
  INV_X1     g10885(.I(\a[44] ), .ZN(new_n11078_));
  NOR2_X1    g10886(.A1(\a[42] ), .A2(\a[43] ), .ZN(new_n11079_));
  INV_X1     g10887(.I(new_n11079_), .ZN(new_n11080_));
  NOR3_X1    g10888(.A1(new_n10620_), .A2(new_n11078_), .A3(new_n11080_), .ZN(new_n11081_));
  NAND2_X1   g10889(.A1(new_n10626_), .A2(new_n11081_), .ZN(new_n11082_));
  XOR2_X1    g10890(.A1(new_n11082_), .A2(\a[45] ), .Z(new_n11083_));
  INV_X1     g10891(.I(\a[45] ), .ZN(new_n11084_));
  NOR4_X1    g10892(.A1(new_n11062_), .A2(new_n11084_), .A3(new_n11035_), .A4(new_n11057_), .ZN(new_n11085_));
  NOR2_X1    g10893(.A1(new_n11084_), .A2(\a[44] ), .ZN(new_n11086_));
  OAI21_X1   g10894(.A1(new_n11085_), .A2(new_n11086_), .B(new_n11083_), .ZN(new_n11087_));
  INV_X1     g10895(.I(new_n11083_), .ZN(new_n11088_));
  INV_X1     g10896(.I(new_n11035_), .ZN(new_n11089_));
  NOR3_X1    g10897(.A1(new_n11032_), .A2(new_n11029_), .A3(new_n11050_), .ZN(new_n11090_));
  AOI21_X1   g10898(.A1(new_n11090_), .A2(new_n11072_), .B(new_n11043_), .ZN(new_n11091_));
  AOI21_X1   g10899(.A1(new_n11091_), .A2(new_n11055_), .B(new_n11041_), .ZN(new_n11092_));
  NAND4_X1   g10900(.A1(new_n10894_), .A2(new_n196_), .A3(new_n11042_), .A4(new_n10582_), .ZN(new_n11093_));
  INV_X1     g10901(.I(new_n11061_), .ZN(new_n11094_));
  NOR2_X1    g10902(.A1(new_n11093_), .A2(new_n11094_), .ZN(new_n11095_));
  NAND4_X1   g10903(.A1(new_n11095_), .A2(\a[45] ), .A3(new_n11092_), .A4(new_n11089_), .ZN(new_n11096_));
  NAND3_X1   g10904(.A1(new_n11096_), .A2(\a[44] ), .A3(new_n11088_), .ZN(new_n11097_));
  NAND2_X1   g10905(.A1(new_n11087_), .A2(new_n11097_), .ZN(new_n11098_));
  NOR2_X1    g10906(.A1(new_n11062_), .A2(new_n11057_), .ZN(new_n11099_));
  NOR4_X1    g10907(.A1(new_n10575_), .A2(new_n10569_), .A3(new_n10616_), .A4(new_n10576_), .ZN(new_n11100_));
  NAND2_X1   g10908(.A1(\asqrt[23] ), .A2(\a[44] ), .ZN(new_n11101_));
  XOR2_X1    g10909(.A1(new_n11101_), .A2(new_n11100_), .Z(new_n11102_));
  NOR2_X1    g10910(.A1(new_n11102_), .A2(new_n11080_), .ZN(new_n11103_));
  INV_X1     g10911(.I(new_n11103_), .ZN(new_n11104_));
  NAND3_X1   g10912(.A1(new_n11095_), .A2(new_n11092_), .A3(new_n11089_), .ZN(new_n11105_));
  NOR2_X1    g10913(.A1(new_n11089_), .A2(new_n11061_), .ZN(new_n11106_));
  NAND2_X1   g10914(.A1(new_n11106_), .A2(\asqrt[23] ), .ZN(new_n11107_));
  INV_X1     g10915(.I(new_n11107_), .ZN(new_n11108_));
  NAND3_X1   g10916(.A1(new_n11057_), .A2(new_n11093_), .A3(new_n11108_), .ZN(new_n11109_));
  NAND2_X1   g10917(.A1(new_n11109_), .A2(new_n10583_), .ZN(new_n11110_));
  NAND3_X1   g10918(.A1(new_n11110_), .A2(new_n10584_), .A3(new_n11105_), .ZN(new_n11111_));
  NOR3_X1    g10919(.A1(new_n11092_), .A2(new_n11058_), .A3(new_n11107_), .ZN(new_n11112_));
  OAI21_X1   g10920(.A1(new_n11112_), .A2(\a[46] ), .B(new_n10584_), .ZN(new_n11113_));
  NAND2_X1   g10921(.A1(new_n11113_), .A2(\asqrt[22] ), .ZN(new_n11114_));
  NAND4_X1   g10922(.A1(new_n11114_), .A2(new_n10104_), .A3(new_n11111_), .A4(new_n11104_), .ZN(new_n11115_));
  NAND2_X1   g10923(.A1(new_n11115_), .A2(new_n11098_), .ZN(new_n11116_));
  NAND3_X1   g10924(.A1(new_n11087_), .A2(new_n11097_), .A3(new_n11104_), .ZN(new_n11117_));
  AOI21_X1   g10925(.A1(\asqrt[23] ), .A2(new_n10583_), .B(\a[47] ), .ZN(new_n11118_));
  NOR2_X1    g10926(.A1(new_n10605_), .A2(\a[46] ), .ZN(new_n11119_));
  AOI21_X1   g10927(.A1(\asqrt[23] ), .A2(\a[46] ), .B(new_n10587_), .ZN(new_n11120_));
  OAI21_X1   g10928(.A1(new_n11119_), .A2(new_n11118_), .B(new_n11120_), .ZN(new_n11121_));
  INV_X1     g10929(.I(new_n11121_), .ZN(new_n11122_));
  NAND3_X1   g10930(.A1(\asqrt[22] ), .A2(new_n10613_), .A3(new_n11122_), .ZN(new_n11123_));
  OAI21_X1   g10931(.A1(new_n11105_), .A2(new_n11121_), .B(new_n10612_), .ZN(new_n11124_));
  NAND3_X1   g10932(.A1(new_n11123_), .A2(new_n11124_), .A3(new_n9672_), .ZN(new_n11125_));
  AOI21_X1   g10933(.A1(new_n11117_), .A2(\asqrt[24] ), .B(new_n11125_), .ZN(new_n11126_));
  NOR2_X1    g10934(.A1(new_n11116_), .A2(new_n11126_), .ZN(new_n11127_));
  AOI22_X1   g10935(.A1(new_n11115_), .A2(new_n11098_), .B1(\asqrt[24] ), .B2(new_n11117_), .ZN(new_n11128_));
  NOR2_X1    g10936(.A1(new_n10901_), .A2(new_n10900_), .ZN(new_n11129_));
  NOR4_X1    g10937(.A1(new_n11105_), .A2(\asqrt[25] ), .A3(new_n11129_), .A4(new_n10632_), .ZN(new_n11130_));
  AOI21_X1   g10938(.A1(new_n10899_), .A2(new_n10613_), .B(new_n9672_), .ZN(new_n11131_));
  NOR2_X1    g10939(.A1(new_n11130_), .A2(new_n11131_), .ZN(new_n11132_));
  NAND2_X1   g10940(.A1(new_n11132_), .A2(new_n9212_), .ZN(new_n11133_));
  INV_X1     g10941(.I(new_n11133_), .ZN(new_n11134_));
  OAI21_X1   g10942(.A1(new_n11128_), .A2(new_n9672_), .B(new_n11134_), .ZN(new_n11135_));
  NAND2_X1   g10943(.A1(new_n11117_), .A2(\asqrt[24] ), .ZN(new_n11136_));
  AOI21_X1   g10944(.A1(new_n11116_), .A2(new_n11136_), .B(new_n9672_), .ZN(new_n11137_));
  OAI21_X1   g10945(.A1(new_n11137_), .A2(new_n11127_), .B(\asqrt[26] ), .ZN(new_n11138_));
  NOR2_X1    g10946(.A1(new_n10644_), .A2(new_n9212_), .ZN(new_n11139_));
  NAND2_X1   g10947(.A1(new_n10638_), .A2(new_n10640_), .ZN(new_n11140_));
  NAND4_X1   g10948(.A1(\asqrt[22] ), .A2(new_n9212_), .A3(new_n11140_), .A4(new_n10644_), .ZN(new_n11141_));
  XOR2_X1    g10949(.A1(new_n11141_), .A2(new_n11139_), .Z(new_n11142_));
  NAND2_X1   g10950(.A1(new_n11142_), .A2(new_n8763_), .ZN(new_n11143_));
  INV_X1     g10951(.I(new_n11143_), .ZN(new_n11144_));
  NAND2_X1   g10952(.A1(new_n11138_), .A2(new_n11144_), .ZN(new_n11145_));
  NAND3_X1   g10953(.A1(new_n11145_), .A2(new_n11127_), .A3(new_n11135_), .ZN(new_n11146_));
  INV_X1     g10954(.I(new_n11086_), .ZN(new_n11147_));
  AOI21_X1   g10955(.A1(new_n11096_), .A2(new_n11147_), .B(new_n11088_), .ZN(new_n11148_));
  NOR3_X1    g10956(.A1(new_n11085_), .A2(new_n11078_), .A3(new_n11083_), .ZN(new_n11149_));
  NOR2_X1    g10957(.A1(new_n11149_), .A2(new_n11148_), .ZN(new_n11150_));
  NOR2_X1    g10958(.A1(new_n11113_), .A2(\asqrt[22] ), .ZN(new_n11151_));
  AOI21_X1   g10959(.A1(new_n11110_), .A2(new_n10584_), .B(new_n11105_), .ZN(new_n11152_));
  NOR4_X1    g10960(.A1(new_n11151_), .A2(\asqrt[24] ), .A3(new_n11152_), .A4(new_n11103_), .ZN(new_n11153_));
  NOR2_X1    g10961(.A1(new_n11153_), .A2(new_n11150_), .ZN(new_n11154_));
  NOR3_X1    g10962(.A1(new_n11149_), .A2(new_n11148_), .A3(new_n11103_), .ZN(new_n11155_));
  NOR3_X1    g10963(.A1(new_n11105_), .A2(new_n10612_), .A3(new_n11121_), .ZN(new_n11156_));
  AOI21_X1   g10964(.A1(\asqrt[22] ), .A2(new_n11122_), .B(new_n10613_), .ZN(new_n11157_));
  NOR3_X1    g10965(.A1(new_n11157_), .A2(new_n11156_), .A3(\asqrt[25] ), .ZN(new_n11158_));
  OAI21_X1   g10966(.A1(new_n11155_), .A2(new_n10104_), .B(new_n11158_), .ZN(new_n11159_));
  NAND2_X1   g10967(.A1(new_n11154_), .A2(new_n11159_), .ZN(new_n11160_));
  OAI22_X1   g10968(.A1(new_n11153_), .A2(new_n11150_), .B1(new_n10104_), .B2(new_n11155_), .ZN(new_n11161_));
  AOI21_X1   g10969(.A1(new_n11161_), .A2(\asqrt[25] ), .B(new_n11133_), .ZN(new_n11162_));
  AOI22_X1   g10970(.A1(new_n11161_), .A2(\asqrt[25] ), .B1(new_n11154_), .B2(new_n11159_), .ZN(new_n11163_));
  OAI22_X1   g10971(.A1(new_n11163_), .A2(new_n9212_), .B1(new_n11162_), .B2(new_n11160_), .ZN(new_n11164_));
  NAND2_X1   g10972(.A1(new_n10651_), .A2(\asqrt[27] ), .ZN(new_n11165_));
  NOR2_X1    g10973(.A1(new_n10646_), .A2(new_n10647_), .ZN(new_n11166_));
  NOR4_X1    g10974(.A1(new_n11105_), .A2(\asqrt[27] ), .A3(new_n11166_), .A4(new_n10651_), .ZN(new_n11167_));
  XOR2_X1    g10975(.A1(new_n11167_), .A2(new_n11165_), .Z(new_n11168_));
  NAND2_X1   g10976(.A1(new_n11168_), .A2(new_n8319_), .ZN(new_n11169_));
  AOI21_X1   g10977(.A1(new_n11164_), .A2(\asqrt[27] ), .B(new_n11169_), .ZN(new_n11170_));
  NOR2_X1    g10978(.A1(new_n11170_), .A2(new_n11146_), .ZN(new_n11171_));
  OAI21_X1   g10979(.A1(new_n11137_), .A2(new_n11133_), .B(new_n11127_), .ZN(new_n11172_));
  AOI21_X1   g10980(.A1(new_n11138_), .A2(new_n11144_), .B(new_n11172_), .ZN(new_n11173_));
  AOI21_X1   g10981(.A1(new_n11172_), .A2(new_n11138_), .B(new_n8763_), .ZN(new_n11174_));
  OAI21_X1   g10982(.A1(new_n11173_), .A2(new_n11174_), .B(\asqrt[28] ), .ZN(new_n11175_));
  NOR4_X1    g10983(.A1(new_n11105_), .A2(\asqrt[28] ), .A3(new_n10654_), .A4(new_n10918_), .ZN(new_n11176_));
  AOI21_X1   g10984(.A1(new_n11165_), .A2(new_n10650_), .B(new_n8319_), .ZN(new_n11177_));
  NOR2_X1    g10985(.A1(new_n11176_), .A2(new_n11177_), .ZN(new_n11178_));
  NAND2_X1   g10986(.A1(new_n11178_), .A2(new_n7931_), .ZN(new_n11179_));
  INV_X1     g10987(.I(new_n11179_), .ZN(new_n11180_));
  NAND2_X1   g10988(.A1(new_n11175_), .A2(new_n11180_), .ZN(new_n11181_));
  NAND2_X1   g10989(.A1(new_n11181_), .A2(new_n11171_), .ZN(new_n11182_));
  NOR2_X1    g10990(.A1(new_n11173_), .A2(new_n11174_), .ZN(new_n11183_));
  OAI22_X1   g10991(.A1(new_n11183_), .A2(new_n8319_), .B1(new_n11170_), .B2(new_n11146_), .ZN(new_n11184_));
  NAND2_X1   g10992(.A1(new_n10666_), .A2(\asqrt[29] ), .ZN(new_n11185_));
  NOR4_X1    g10993(.A1(new_n11105_), .A2(\asqrt[29] ), .A3(new_n10661_), .A4(new_n10666_), .ZN(new_n11186_));
  XOR2_X1    g10994(.A1(new_n11186_), .A2(new_n11185_), .Z(new_n11187_));
  NAND2_X1   g10995(.A1(new_n11187_), .A2(new_n7517_), .ZN(new_n11188_));
  AOI21_X1   g10996(.A1(new_n11184_), .A2(\asqrt[29] ), .B(new_n11188_), .ZN(new_n11189_));
  NOR2_X1    g10997(.A1(new_n11189_), .A2(new_n11182_), .ZN(new_n11190_));
  OAI21_X1   g10998(.A1(new_n11174_), .A2(new_n11169_), .B(new_n11173_), .ZN(new_n11191_));
  AOI21_X1   g10999(.A1(new_n11175_), .A2(new_n11180_), .B(new_n11191_), .ZN(new_n11192_));
  AOI21_X1   g11000(.A1(new_n11191_), .A2(new_n11175_), .B(new_n7931_), .ZN(new_n11193_));
  OAI21_X1   g11001(.A1(new_n11192_), .A2(new_n11193_), .B(\asqrt[30] ), .ZN(new_n11194_));
  NOR4_X1    g11002(.A1(new_n11105_), .A2(\asqrt[30] ), .A3(new_n10668_), .A4(new_n10925_), .ZN(new_n11195_));
  AOI21_X1   g11003(.A1(new_n11185_), .A2(new_n10665_), .B(new_n7517_), .ZN(new_n11196_));
  NOR2_X1    g11004(.A1(new_n11195_), .A2(new_n11196_), .ZN(new_n11197_));
  NAND2_X1   g11005(.A1(new_n11197_), .A2(new_n7110_), .ZN(new_n11198_));
  INV_X1     g11006(.I(new_n11198_), .ZN(new_n11199_));
  NAND2_X1   g11007(.A1(new_n11194_), .A2(new_n11199_), .ZN(new_n11200_));
  NAND2_X1   g11008(.A1(new_n11200_), .A2(new_n11190_), .ZN(new_n11201_));
  AOI22_X1   g11009(.A1(new_n11184_), .A2(\asqrt[29] ), .B1(new_n11181_), .B2(new_n11171_), .ZN(new_n11202_));
  OAI22_X1   g11010(.A1(new_n11202_), .A2(new_n7517_), .B1(new_n11189_), .B2(new_n11182_), .ZN(new_n11203_));
  NAND2_X1   g11011(.A1(new_n10679_), .A2(\asqrt[31] ), .ZN(new_n11204_));
  NOR4_X1    g11012(.A1(new_n11105_), .A2(\asqrt[31] ), .A3(new_n10674_), .A4(new_n10679_), .ZN(new_n11205_));
  XOR2_X1    g11013(.A1(new_n11205_), .A2(new_n11204_), .Z(new_n11206_));
  NAND2_X1   g11014(.A1(new_n11206_), .A2(new_n6708_), .ZN(new_n11207_));
  AOI21_X1   g11015(.A1(new_n11203_), .A2(\asqrt[31] ), .B(new_n11207_), .ZN(new_n11208_));
  NOR2_X1    g11016(.A1(new_n11208_), .A2(new_n11201_), .ZN(new_n11209_));
  AOI22_X1   g11017(.A1(new_n11203_), .A2(\asqrt[31] ), .B1(new_n11200_), .B2(new_n11190_), .ZN(new_n11210_));
  NOR4_X1    g11018(.A1(new_n11105_), .A2(\asqrt[32] ), .A3(new_n10681_), .A4(new_n10932_), .ZN(new_n11211_));
  AOI21_X1   g11019(.A1(new_n11204_), .A2(new_n10678_), .B(new_n6708_), .ZN(new_n11212_));
  NOR2_X1    g11020(.A1(new_n11211_), .A2(new_n11212_), .ZN(new_n11213_));
  NAND2_X1   g11021(.A1(new_n11213_), .A2(new_n6365_), .ZN(new_n11214_));
  INV_X1     g11022(.I(new_n11214_), .ZN(new_n11215_));
  OAI21_X1   g11023(.A1(new_n11210_), .A2(new_n6708_), .B(new_n11215_), .ZN(new_n11216_));
  NAND2_X1   g11024(.A1(new_n11216_), .A2(new_n11209_), .ZN(new_n11217_));
  OAI22_X1   g11025(.A1(new_n11210_), .A2(new_n6708_), .B1(new_n11208_), .B2(new_n11201_), .ZN(new_n11218_));
  NAND2_X1   g11026(.A1(new_n10692_), .A2(\asqrt[33] ), .ZN(new_n11219_));
  NOR4_X1    g11027(.A1(new_n11105_), .A2(\asqrt[33] ), .A3(new_n10687_), .A4(new_n10692_), .ZN(new_n11220_));
  XOR2_X1    g11028(.A1(new_n11220_), .A2(new_n11219_), .Z(new_n11221_));
  NAND2_X1   g11029(.A1(new_n11221_), .A2(new_n5991_), .ZN(new_n11222_));
  AOI21_X1   g11030(.A1(new_n11218_), .A2(\asqrt[33] ), .B(new_n11222_), .ZN(new_n11223_));
  NOR2_X1    g11031(.A1(new_n11223_), .A2(new_n11217_), .ZN(new_n11224_));
  AOI22_X1   g11032(.A1(new_n11218_), .A2(\asqrt[33] ), .B1(new_n11216_), .B2(new_n11209_), .ZN(new_n11225_));
  NAND2_X1   g11033(.A1(new_n10939_), .A2(\asqrt[34] ), .ZN(new_n11226_));
  NOR4_X1    g11034(.A1(new_n11105_), .A2(\asqrt[34] ), .A3(new_n10695_), .A4(new_n10939_), .ZN(new_n11227_));
  XOR2_X1    g11035(.A1(new_n11227_), .A2(new_n11226_), .Z(new_n11228_));
  NAND2_X1   g11036(.A1(new_n11228_), .A2(new_n5626_), .ZN(new_n11229_));
  INV_X1     g11037(.I(new_n11229_), .ZN(new_n11230_));
  OAI21_X1   g11038(.A1(new_n11225_), .A2(new_n5991_), .B(new_n11230_), .ZN(new_n11231_));
  NAND2_X1   g11039(.A1(new_n11231_), .A2(new_n11224_), .ZN(new_n11232_));
  OAI22_X1   g11040(.A1(new_n11225_), .A2(new_n5991_), .B1(new_n11223_), .B2(new_n11217_), .ZN(new_n11233_));
  NOR4_X1    g11041(.A1(new_n11105_), .A2(\asqrt[35] ), .A3(new_n10702_), .A4(new_n10707_), .ZN(new_n11234_));
  AOI21_X1   g11042(.A1(new_n11226_), .A2(new_n10938_), .B(new_n5626_), .ZN(new_n11235_));
  NOR2_X1    g11043(.A1(new_n11234_), .A2(new_n11235_), .ZN(new_n11236_));
  NAND2_X1   g11044(.A1(new_n11236_), .A2(new_n5273_), .ZN(new_n11237_));
  AOI21_X1   g11045(.A1(new_n11233_), .A2(\asqrt[35] ), .B(new_n11237_), .ZN(new_n11238_));
  NOR2_X1    g11046(.A1(new_n11238_), .A2(new_n11232_), .ZN(new_n11239_));
  AOI22_X1   g11047(.A1(new_n11233_), .A2(\asqrt[35] ), .B1(new_n11231_), .B2(new_n11224_), .ZN(new_n11240_));
  NAND2_X1   g11048(.A1(new_n10946_), .A2(\asqrt[36] ), .ZN(new_n11241_));
  NOR4_X1    g11049(.A1(new_n11105_), .A2(\asqrt[36] ), .A3(new_n10710_), .A4(new_n10946_), .ZN(new_n11242_));
  XOR2_X1    g11050(.A1(new_n11242_), .A2(new_n11241_), .Z(new_n11243_));
  NAND2_X1   g11051(.A1(new_n11243_), .A2(new_n4973_), .ZN(new_n11244_));
  INV_X1     g11052(.I(new_n11244_), .ZN(new_n11245_));
  OAI21_X1   g11053(.A1(new_n11240_), .A2(new_n5273_), .B(new_n11245_), .ZN(new_n11246_));
  NAND2_X1   g11054(.A1(new_n11246_), .A2(new_n11239_), .ZN(new_n11247_));
  OAI22_X1   g11055(.A1(new_n11240_), .A2(new_n5273_), .B1(new_n11238_), .B2(new_n11232_), .ZN(new_n11248_));
  NOR4_X1    g11056(.A1(new_n11105_), .A2(\asqrt[37] ), .A3(new_n10717_), .A4(new_n10722_), .ZN(new_n11249_));
  AOI21_X1   g11057(.A1(new_n11241_), .A2(new_n10945_), .B(new_n4973_), .ZN(new_n11250_));
  NOR2_X1    g11058(.A1(new_n11249_), .A2(new_n11250_), .ZN(new_n11251_));
  NAND2_X1   g11059(.A1(new_n11251_), .A2(new_n4645_), .ZN(new_n11252_));
  AOI21_X1   g11060(.A1(new_n11248_), .A2(\asqrt[37] ), .B(new_n11252_), .ZN(new_n11253_));
  NOR2_X1    g11061(.A1(new_n11253_), .A2(new_n11247_), .ZN(new_n11254_));
  AOI22_X1   g11062(.A1(new_n11248_), .A2(\asqrt[37] ), .B1(new_n11246_), .B2(new_n11239_), .ZN(new_n11255_));
  NAND2_X1   g11063(.A1(new_n10953_), .A2(\asqrt[38] ), .ZN(new_n11256_));
  NOR4_X1    g11064(.A1(new_n11105_), .A2(\asqrt[38] ), .A3(new_n10725_), .A4(new_n10953_), .ZN(new_n11257_));
  XOR2_X1    g11065(.A1(new_n11257_), .A2(new_n11256_), .Z(new_n11258_));
  NAND2_X1   g11066(.A1(new_n11258_), .A2(new_n4330_), .ZN(new_n11259_));
  INV_X1     g11067(.I(new_n11259_), .ZN(new_n11260_));
  OAI21_X1   g11068(.A1(new_n11255_), .A2(new_n4645_), .B(new_n11260_), .ZN(new_n11261_));
  NAND2_X1   g11069(.A1(new_n11261_), .A2(new_n11254_), .ZN(new_n11262_));
  OAI22_X1   g11070(.A1(new_n11255_), .A2(new_n4645_), .B1(new_n11253_), .B2(new_n11247_), .ZN(new_n11263_));
  NOR4_X1    g11071(.A1(new_n11105_), .A2(\asqrt[39] ), .A3(new_n10732_), .A4(new_n10737_), .ZN(new_n11264_));
  AOI21_X1   g11072(.A1(new_n11256_), .A2(new_n10952_), .B(new_n4330_), .ZN(new_n11265_));
  NOR2_X1    g11073(.A1(new_n11264_), .A2(new_n11265_), .ZN(new_n11266_));
  NAND2_X1   g11074(.A1(new_n11266_), .A2(new_n4018_), .ZN(new_n11267_));
  AOI21_X1   g11075(.A1(new_n11263_), .A2(\asqrt[39] ), .B(new_n11267_), .ZN(new_n11268_));
  NOR2_X1    g11076(.A1(new_n11268_), .A2(new_n11262_), .ZN(new_n11269_));
  AOI22_X1   g11077(.A1(new_n11263_), .A2(\asqrt[39] ), .B1(new_n11261_), .B2(new_n11254_), .ZN(new_n11270_));
  NAND2_X1   g11078(.A1(new_n10960_), .A2(\asqrt[40] ), .ZN(new_n11271_));
  NOR4_X1    g11079(.A1(new_n11105_), .A2(\asqrt[40] ), .A3(new_n10740_), .A4(new_n10960_), .ZN(new_n11272_));
  XOR2_X1    g11080(.A1(new_n11272_), .A2(new_n11271_), .Z(new_n11273_));
  NAND2_X1   g11081(.A1(new_n11273_), .A2(new_n3760_), .ZN(new_n11274_));
  INV_X1     g11082(.I(new_n11274_), .ZN(new_n11275_));
  OAI21_X1   g11083(.A1(new_n11270_), .A2(new_n4018_), .B(new_n11275_), .ZN(new_n11276_));
  NAND2_X1   g11084(.A1(new_n11276_), .A2(new_n11269_), .ZN(new_n11277_));
  OAI22_X1   g11085(.A1(new_n11270_), .A2(new_n4018_), .B1(new_n11268_), .B2(new_n11262_), .ZN(new_n11278_));
  NOR4_X1    g11086(.A1(new_n11105_), .A2(\asqrt[41] ), .A3(new_n10747_), .A4(new_n10752_), .ZN(new_n11279_));
  AOI21_X1   g11087(.A1(new_n11271_), .A2(new_n10959_), .B(new_n3760_), .ZN(new_n11280_));
  NOR2_X1    g11088(.A1(new_n11279_), .A2(new_n11280_), .ZN(new_n11281_));
  NAND2_X1   g11089(.A1(new_n11281_), .A2(new_n3481_), .ZN(new_n11282_));
  AOI21_X1   g11090(.A1(new_n11278_), .A2(\asqrt[41] ), .B(new_n11282_), .ZN(new_n11283_));
  NOR2_X1    g11091(.A1(new_n11283_), .A2(new_n11277_), .ZN(new_n11284_));
  AOI22_X1   g11092(.A1(new_n11278_), .A2(\asqrt[41] ), .B1(new_n11276_), .B2(new_n11269_), .ZN(new_n11285_));
  NAND2_X1   g11093(.A1(new_n10967_), .A2(\asqrt[42] ), .ZN(new_n11286_));
  NOR4_X1    g11094(.A1(new_n11105_), .A2(\asqrt[42] ), .A3(new_n10755_), .A4(new_n10967_), .ZN(new_n11287_));
  XOR2_X1    g11095(.A1(new_n11287_), .A2(new_n11286_), .Z(new_n11288_));
  NAND2_X1   g11096(.A1(new_n11288_), .A2(new_n3208_), .ZN(new_n11289_));
  INV_X1     g11097(.I(new_n11289_), .ZN(new_n11290_));
  OAI21_X1   g11098(.A1(new_n11285_), .A2(new_n3481_), .B(new_n11290_), .ZN(new_n11291_));
  NAND2_X1   g11099(.A1(new_n11291_), .A2(new_n11284_), .ZN(new_n11292_));
  OAI22_X1   g11100(.A1(new_n11285_), .A2(new_n3481_), .B1(new_n11283_), .B2(new_n11277_), .ZN(new_n11293_));
  NAND2_X1   g11101(.A1(new_n10767_), .A2(\asqrt[43] ), .ZN(new_n11294_));
  NOR4_X1    g11102(.A1(new_n11105_), .A2(\asqrt[43] ), .A3(new_n10762_), .A4(new_n10767_), .ZN(new_n11295_));
  XOR2_X1    g11103(.A1(new_n11295_), .A2(new_n11294_), .Z(new_n11296_));
  NAND2_X1   g11104(.A1(new_n11296_), .A2(new_n2941_), .ZN(new_n11297_));
  AOI21_X1   g11105(.A1(new_n11293_), .A2(\asqrt[43] ), .B(new_n11297_), .ZN(new_n11298_));
  NOR2_X1    g11106(.A1(new_n11298_), .A2(new_n11292_), .ZN(new_n11299_));
  AOI22_X1   g11107(.A1(new_n11293_), .A2(\asqrt[43] ), .B1(new_n11291_), .B2(new_n11284_), .ZN(new_n11300_));
  NOR4_X1    g11108(.A1(new_n11105_), .A2(\asqrt[44] ), .A3(new_n10770_), .A4(new_n10974_), .ZN(new_n11301_));
  AOI21_X1   g11109(.A1(new_n11294_), .A2(new_n10766_), .B(new_n2941_), .ZN(new_n11302_));
  NOR2_X1    g11110(.A1(new_n11301_), .A2(new_n11302_), .ZN(new_n11303_));
  NAND2_X1   g11111(.A1(new_n11303_), .A2(new_n2728_), .ZN(new_n11304_));
  INV_X1     g11112(.I(new_n11304_), .ZN(new_n11305_));
  OAI21_X1   g11113(.A1(new_n11300_), .A2(new_n2941_), .B(new_n11305_), .ZN(new_n11306_));
  NAND2_X1   g11114(.A1(new_n11306_), .A2(new_n11299_), .ZN(new_n11307_));
  OAI22_X1   g11115(.A1(new_n11300_), .A2(new_n2941_), .B1(new_n11298_), .B2(new_n11292_), .ZN(new_n11308_));
  NAND2_X1   g11116(.A1(new_n10782_), .A2(\asqrt[45] ), .ZN(new_n11309_));
  NOR4_X1    g11117(.A1(new_n11105_), .A2(\asqrt[45] ), .A3(new_n10777_), .A4(new_n10782_), .ZN(new_n11310_));
  XOR2_X1    g11118(.A1(new_n11310_), .A2(new_n11309_), .Z(new_n11311_));
  NAND2_X1   g11119(.A1(new_n11311_), .A2(new_n2488_), .ZN(new_n11312_));
  AOI21_X1   g11120(.A1(new_n11308_), .A2(\asqrt[45] ), .B(new_n11312_), .ZN(new_n11313_));
  NOR2_X1    g11121(.A1(new_n11313_), .A2(new_n11307_), .ZN(new_n11314_));
  AOI22_X1   g11122(.A1(new_n11308_), .A2(\asqrt[45] ), .B1(new_n11306_), .B2(new_n11299_), .ZN(new_n11315_));
  NOR4_X1    g11123(.A1(new_n11105_), .A2(\asqrt[46] ), .A3(new_n10785_), .A4(new_n10981_), .ZN(new_n11316_));
  AOI21_X1   g11124(.A1(new_n11309_), .A2(new_n10781_), .B(new_n2488_), .ZN(new_n11317_));
  NOR2_X1    g11125(.A1(new_n11316_), .A2(new_n11317_), .ZN(new_n11318_));
  NAND2_X1   g11126(.A1(new_n11318_), .A2(new_n2253_), .ZN(new_n11319_));
  INV_X1     g11127(.I(new_n11319_), .ZN(new_n11320_));
  OAI21_X1   g11128(.A1(new_n11315_), .A2(new_n2488_), .B(new_n11320_), .ZN(new_n11321_));
  NAND2_X1   g11129(.A1(new_n11321_), .A2(new_n11314_), .ZN(new_n11322_));
  OAI22_X1   g11130(.A1(new_n11315_), .A2(new_n2488_), .B1(new_n11313_), .B2(new_n11307_), .ZN(new_n11323_));
  NAND2_X1   g11131(.A1(new_n10797_), .A2(\asqrt[47] ), .ZN(new_n11324_));
  NOR4_X1    g11132(.A1(new_n11105_), .A2(\asqrt[47] ), .A3(new_n10792_), .A4(new_n10797_), .ZN(new_n11325_));
  XOR2_X1    g11133(.A1(new_n11325_), .A2(new_n11324_), .Z(new_n11326_));
  NAND2_X1   g11134(.A1(new_n11326_), .A2(new_n2046_), .ZN(new_n11327_));
  AOI21_X1   g11135(.A1(new_n11323_), .A2(\asqrt[47] ), .B(new_n11327_), .ZN(new_n11328_));
  NOR2_X1    g11136(.A1(new_n11328_), .A2(new_n11322_), .ZN(new_n11329_));
  AOI22_X1   g11137(.A1(new_n11323_), .A2(\asqrt[47] ), .B1(new_n11321_), .B2(new_n11314_), .ZN(new_n11330_));
  NAND2_X1   g11138(.A1(new_n10988_), .A2(\asqrt[48] ), .ZN(new_n11331_));
  NOR4_X1    g11139(.A1(new_n11105_), .A2(\asqrt[48] ), .A3(new_n10800_), .A4(new_n10988_), .ZN(new_n11332_));
  XOR2_X1    g11140(.A1(new_n11332_), .A2(new_n11331_), .Z(new_n11333_));
  NAND2_X1   g11141(.A1(new_n11333_), .A2(new_n1854_), .ZN(new_n11334_));
  INV_X1     g11142(.I(new_n11334_), .ZN(new_n11335_));
  OAI21_X1   g11143(.A1(new_n11330_), .A2(new_n2046_), .B(new_n11335_), .ZN(new_n11336_));
  NAND2_X1   g11144(.A1(new_n11336_), .A2(new_n11329_), .ZN(new_n11337_));
  OAI22_X1   g11145(.A1(new_n11330_), .A2(new_n2046_), .B1(new_n11328_), .B2(new_n11322_), .ZN(new_n11338_));
  NOR4_X1    g11146(.A1(new_n11105_), .A2(\asqrt[49] ), .A3(new_n10807_), .A4(new_n10812_), .ZN(new_n11339_));
  AOI21_X1   g11147(.A1(new_n11331_), .A2(new_n10987_), .B(new_n1854_), .ZN(new_n11340_));
  NOR2_X1    g11148(.A1(new_n11339_), .A2(new_n11340_), .ZN(new_n11341_));
  NAND2_X1   g11149(.A1(new_n11341_), .A2(new_n1595_), .ZN(new_n11342_));
  AOI21_X1   g11150(.A1(new_n11338_), .A2(\asqrt[49] ), .B(new_n11342_), .ZN(new_n11343_));
  NOR2_X1    g11151(.A1(new_n11343_), .A2(new_n11337_), .ZN(new_n11344_));
  AOI22_X1   g11152(.A1(new_n11338_), .A2(\asqrt[49] ), .B1(new_n11336_), .B2(new_n11329_), .ZN(new_n11345_));
  NAND2_X1   g11153(.A1(new_n10995_), .A2(\asqrt[50] ), .ZN(new_n11346_));
  NOR4_X1    g11154(.A1(new_n11105_), .A2(\asqrt[50] ), .A3(new_n10815_), .A4(new_n10995_), .ZN(new_n11347_));
  XOR2_X1    g11155(.A1(new_n11347_), .A2(new_n11346_), .Z(new_n11348_));
  NAND2_X1   g11156(.A1(new_n11348_), .A2(new_n1436_), .ZN(new_n11349_));
  INV_X1     g11157(.I(new_n11349_), .ZN(new_n11350_));
  OAI21_X1   g11158(.A1(new_n11345_), .A2(new_n1595_), .B(new_n11350_), .ZN(new_n11351_));
  NAND2_X1   g11159(.A1(new_n11351_), .A2(new_n11344_), .ZN(new_n11352_));
  OAI22_X1   g11160(.A1(new_n11345_), .A2(new_n1595_), .B1(new_n11343_), .B2(new_n11337_), .ZN(new_n11353_));
  NOR4_X1    g11161(.A1(new_n11105_), .A2(\asqrt[51] ), .A3(new_n10822_), .A4(new_n10827_), .ZN(new_n11354_));
  AOI21_X1   g11162(.A1(new_n11346_), .A2(new_n10994_), .B(new_n1436_), .ZN(new_n11355_));
  NOR2_X1    g11163(.A1(new_n11354_), .A2(new_n11355_), .ZN(new_n11356_));
  NAND2_X1   g11164(.A1(new_n11356_), .A2(new_n1260_), .ZN(new_n11357_));
  AOI21_X1   g11165(.A1(new_n11353_), .A2(\asqrt[51] ), .B(new_n11357_), .ZN(new_n11358_));
  NOR2_X1    g11166(.A1(new_n11358_), .A2(new_n11352_), .ZN(new_n11359_));
  AOI22_X1   g11167(.A1(new_n11353_), .A2(\asqrt[51] ), .B1(new_n11351_), .B2(new_n11344_), .ZN(new_n11360_));
  NAND2_X1   g11168(.A1(new_n11002_), .A2(\asqrt[52] ), .ZN(new_n11361_));
  NOR4_X1    g11169(.A1(new_n11105_), .A2(\asqrt[52] ), .A3(new_n10830_), .A4(new_n11002_), .ZN(new_n11362_));
  XOR2_X1    g11170(.A1(new_n11362_), .A2(new_n11361_), .Z(new_n11363_));
  NAND2_X1   g11171(.A1(new_n11363_), .A2(new_n1096_), .ZN(new_n11364_));
  INV_X1     g11172(.I(new_n11364_), .ZN(new_n11365_));
  OAI21_X1   g11173(.A1(new_n11360_), .A2(new_n1260_), .B(new_n11365_), .ZN(new_n11366_));
  NAND2_X1   g11174(.A1(new_n11366_), .A2(new_n11359_), .ZN(new_n11367_));
  OAI22_X1   g11175(.A1(new_n11360_), .A2(new_n1260_), .B1(new_n11358_), .B2(new_n11352_), .ZN(new_n11368_));
  NOR4_X1    g11176(.A1(new_n11105_), .A2(\asqrt[53] ), .A3(new_n10837_), .A4(new_n10842_), .ZN(new_n11369_));
  AOI21_X1   g11177(.A1(new_n11361_), .A2(new_n11001_), .B(new_n1096_), .ZN(new_n11370_));
  NOR2_X1    g11178(.A1(new_n11369_), .A2(new_n11370_), .ZN(new_n11371_));
  NAND2_X1   g11179(.A1(new_n11371_), .A2(new_n970_), .ZN(new_n11372_));
  AOI21_X1   g11180(.A1(new_n11368_), .A2(\asqrt[53] ), .B(new_n11372_), .ZN(new_n11373_));
  NOR2_X1    g11181(.A1(new_n11373_), .A2(new_n11367_), .ZN(new_n11374_));
  AOI22_X1   g11182(.A1(new_n11368_), .A2(\asqrt[53] ), .B1(new_n11366_), .B2(new_n11359_), .ZN(new_n11375_));
  NAND2_X1   g11183(.A1(new_n11009_), .A2(\asqrt[54] ), .ZN(new_n11376_));
  NOR4_X1    g11184(.A1(new_n11105_), .A2(\asqrt[54] ), .A3(new_n10844_), .A4(new_n11009_), .ZN(new_n11377_));
  XOR2_X1    g11185(.A1(new_n11377_), .A2(new_n11376_), .Z(new_n11378_));
  NAND2_X1   g11186(.A1(new_n11378_), .A2(new_n825_), .ZN(new_n11379_));
  INV_X1     g11187(.I(new_n11379_), .ZN(new_n11380_));
  OAI21_X1   g11188(.A1(new_n11375_), .A2(new_n970_), .B(new_n11380_), .ZN(new_n11381_));
  NAND2_X1   g11189(.A1(new_n11381_), .A2(new_n11374_), .ZN(new_n11382_));
  OAI22_X1   g11190(.A1(new_n11375_), .A2(new_n970_), .B1(new_n11373_), .B2(new_n11367_), .ZN(new_n11383_));
  NAND2_X1   g11191(.A1(new_n10855_), .A2(\asqrt[55] ), .ZN(new_n11384_));
  NOR4_X1    g11192(.A1(new_n11105_), .A2(\asqrt[55] ), .A3(new_n10850_), .A4(new_n10855_), .ZN(new_n11385_));
  XOR2_X1    g11193(.A1(new_n11385_), .A2(new_n11384_), .Z(new_n11386_));
  NAND2_X1   g11194(.A1(new_n11386_), .A2(new_n724_), .ZN(new_n11387_));
  AOI21_X1   g11195(.A1(new_n11383_), .A2(\asqrt[55] ), .B(new_n11387_), .ZN(new_n11388_));
  NOR2_X1    g11196(.A1(new_n11388_), .A2(new_n11382_), .ZN(new_n11389_));
  AOI22_X1   g11197(.A1(new_n11383_), .A2(\asqrt[55] ), .B1(new_n11381_), .B2(new_n11374_), .ZN(new_n11390_));
  NOR4_X1    g11198(.A1(new_n11105_), .A2(\asqrt[56] ), .A3(new_n10857_), .A4(new_n11016_), .ZN(new_n11391_));
  AOI21_X1   g11199(.A1(new_n11384_), .A2(new_n10854_), .B(new_n724_), .ZN(new_n11392_));
  NOR2_X1    g11200(.A1(new_n11391_), .A2(new_n11392_), .ZN(new_n11393_));
  NAND2_X1   g11201(.A1(new_n11393_), .A2(new_n587_), .ZN(new_n11394_));
  INV_X1     g11202(.I(new_n11394_), .ZN(new_n11395_));
  OAI21_X1   g11203(.A1(new_n11390_), .A2(new_n724_), .B(new_n11395_), .ZN(new_n11396_));
  NAND2_X1   g11204(.A1(new_n11396_), .A2(new_n11389_), .ZN(new_n11397_));
  NAND2_X1   g11205(.A1(new_n11368_), .A2(\asqrt[53] ), .ZN(new_n11398_));
  AOI21_X1   g11206(.A1(new_n11398_), .A2(new_n11367_), .B(new_n970_), .ZN(new_n11399_));
  OAI21_X1   g11207(.A1(new_n11374_), .A2(new_n11399_), .B(\asqrt[55] ), .ZN(new_n11400_));
  AOI21_X1   g11208(.A1(new_n11382_), .A2(new_n11400_), .B(new_n724_), .ZN(new_n11401_));
  OAI21_X1   g11209(.A1(new_n11389_), .A2(new_n11401_), .B(\asqrt[57] ), .ZN(new_n11402_));
  NOR4_X1    g11210(.A1(new_n11105_), .A2(\asqrt[57] ), .A3(new_n10863_), .A4(new_n10868_), .ZN(new_n11403_));
  XOR2_X1    g11211(.A1(new_n11403_), .A2(new_n11045_), .Z(new_n11404_));
  NAND2_X1   g11212(.A1(new_n11404_), .A2(new_n504_), .ZN(new_n11405_));
  INV_X1     g11213(.I(new_n11405_), .ZN(new_n11406_));
  AOI21_X1   g11214(.A1(new_n11402_), .A2(new_n11406_), .B(new_n11397_), .ZN(new_n11407_));
  OAI22_X1   g11215(.A1(new_n11390_), .A2(new_n724_), .B1(new_n11388_), .B2(new_n11382_), .ZN(new_n11408_));
  AOI22_X1   g11216(.A1(new_n11408_), .A2(\asqrt[57] ), .B1(new_n11396_), .B2(new_n11389_), .ZN(new_n11409_));
  NOR4_X1    g11217(.A1(new_n11105_), .A2(\asqrt[58] ), .A3(new_n10870_), .A4(new_n11023_), .ZN(new_n11410_));
  XOR2_X1    g11218(.A1(new_n11410_), .A2(new_n11069_), .Z(new_n11411_));
  NAND2_X1   g11219(.A1(new_n11411_), .A2(new_n376_), .ZN(new_n11412_));
  INV_X1     g11220(.I(new_n11412_), .ZN(new_n11413_));
  OAI21_X1   g11221(.A1(new_n11409_), .A2(new_n504_), .B(new_n11413_), .ZN(new_n11414_));
  NAND2_X1   g11222(.A1(new_n11414_), .A2(new_n11407_), .ZN(new_n11415_));
  AOI21_X1   g11223(.A1(new_n11397_), .A2(new_n11402_), .B(new_n504_), .ZN(new_n11416_));
  OAI21_X1   g11224(.A1(new_n11407_), .A2(new_n11416_), .B(\asqrt[59] ), .ZN(new_n11417_));
  NOR4_X1    g11225(.A1(new_n11105_), .A2(\asqrt[59] ), .A3(new_n10876_), .A4(new_n10881_), .ZN(new_n11418_));
  XOR2_X1    g11226(.A1(new_n11418_), .A2(new_n11047_), .Z(new_n11419_));
  AND2_X2    g11227(.A1(new_n11419_), .A2(new_n275_), .Z(new_n11420_));
  AOI21_X1   g11228(.A1(new_n11417_), .A2(new_n11420_), .B(new_n11415_), .ZN(new_n11421_));
  OAI22_X1   g11229(.A1(new_n11128_), .A2(new_n9672_), .B1(new_n11116_), .B2(new_n11126_), .ZN(new_n11422_));
  AOI22_X1   g11230(.A1(new_n11422_), .A2(\asqrt[26] ), .B1(new_n11135_), .B2(new_n11127_), .ZN(new_n11423_));
  INV_X1     g11231(.I(new_n11169_), .ZN(new_n11424_));
  OAI21_X1   g11232(.A1(new_n11423_), .A2(new_n8763_), .B(new_n11424_), .ZN(new_n11425_));
  AOI21_X1   g11233(.A1(new_n11422_), .A2(\asqrt[26] ), .B(new_n11143_), .ZN(new_n11426_));
  OAI22_X1   g11234(.A1(new_n11423_), .A2(new_n8763_), .B1(new_n11426_), .B2(new_n11172_), .ZN(new_n11427_));
  AOI22_X1   g11235(.A1(new_n11427_), .A2(\asqrt[28] ), .B1(new_n11425_), .B2(new_n11173_), .ZN(new_n11428_));
  INV_X1     g11236(.I(new_n11188_), .ZN(new_n11429_));
  OAI21_X1   g11237(.A1(new_n11428_), .A2(new_n7931_), .B(new_n11429_), .ZN(new_n11430_));
  NAND2_X1   g11238(.A1(new_n11430_), .A2(new_n11192_), .ZN(new_n11431_));
  AOI21_X1   g11239(.A1(new_n11427_), .A2(\asqrt[28] ), .B(new_n11179_), .ZN(new_n11432_));
  OAI22_X1   g11240(.A1(new_n11428_), .A2(new_n7931_), .B1(new_n11432_), .B2(new_n11191_), .ZN(new_n11433_));
  AOI21_X1   g11241(.A1(new_n11433_), .A2(\asqrt[30] ), .B(new_n11198_), .ZN(new_n11434_));
  NOR2_X1    g11242(.A1(new_n11434_), .A2(new_n11431_), .ZN(new_n11435_));
  AOI22_X1   g11243(.A1(new_n11433_), .A2(\asqrt[30] ), .B1(new_n11430_), .B2(new_n11192_), .ZN(new_n11436_));
  INV_X1     g11244(.I(new_n11207_), .ZN(new_n11437_));
  OAI21_X1   g11245(.A1(new_n11436_), .A2(new_n7110_), .B(new_n11437_), .ZN(new_n11438_));
  NAND2_X1   g11246(.A1(new_n11438_), .A2(new_n11435_), .ZN(new_n11439_));
  OAI22_X1   g11247(.A1(new_n11436_), .A2(new_n7110_), .B1(new_n11434_), .B2(new_n11431_), .ZN(new_n11440_));
  AOI21_X1   g11248(.A1(new_n11440_), .A2(\asqrt[32] ), .B(new_n11214_), .ZN(new_n11441_));
  NOR2_X1    g11249(.A1(new_n11441_), .A2(new_n11439_), .ZN(new_n11442_));
  AOI22_X1   g11250(.A1(new_n11440_), .A2(\asqrt[32] ), .B1(new_n11438_), .B2(new_n11435_), .ZN(new_n11443_));
  INV_X1     g11251(.I(new_n11222_), .ZN(new_n11444_));
  OAI21_X1   g11252(.A1(new_n11443_), .A2(new_n6365_), .B(new_n11444_), .ZN(new_n11445_));
  NAND2_X1   g11253(.A1(new_n11445_), .A2(new_n11442_), .ZN(new_n11446_));
  OAI22_X1   g11254(.A1(new_n11443_), .A2(new_n6365_), .B1(new_n11441_), .B2(new_n11439_), .ZN(new_n11447_));
  AOI21_X1   g11255(.A1(new_n11447_), .A2(\asqrt[34] ), .B(new_n11229_), .ZN(new_n11448_));
  NOR2_X1    g11256(.A1(new_n11448_), .A2(new_n11446_), .ZN(new_n11449_));
  AOI22_X1   g11257(.A1(new_n11447_), .A2(\asqrt[34] ), .B1(new_n11445_), .B2(new_n11442_), .ZN(new_n11450_));
  INV_X1     g11258(.I(new_n11237_), .ZN(new_n11451_));
  OAI21_X1   g11259(.A1(new_n11450_), .A2(new_n5626_), .B(new_n11451_), .ZN(new_n11452_));
  NAND2_X1   g11260(.A1(new_n11452_), .A2(new_n11449_), .ZN(new_n11453_));
  OAI22_X1   g11261(.A1(new_n11450_), .A2(new_n5626_), .B1(new_n11448_), .B2(new_n11446_), .ZN(new_n11454_));
  AOI21_X1   g11262(.A1(new_n11454_), .A2(\asqrt[36] ), .B(new_n11244_), .ZN(new_n11455_));
  NOR2_X1    g11263(.A1(new_n11455_), .A2(new_n11453_), .ZN(new_n11456_));
  AOI22_X1   g11264(.A1(new_n11454_), .A2(\asqrt[36] ), .B1(new_n11452_), .B2(new_n11449_), .ZN(new_n11457_));
  INV_X1     g11265(.I(new_n11252_), .ZN(new_n11458_));
  OAI21_X1   g11266(.A1(new_n11457_), .A2(new_n4973_), .B(new_n11458_), .ZN(new_n11459_));
  NAND2_X1   g11267(.A1(new_n11459_), .A2(new_n11456_), .ZN(new_n11460_));
  OAI22_X1   g11268(.A1(new_n11457_), .A2(new_n4973_), .B1(new_n11455_), .B2(new_n11453_), .ZN(new_n11461_));
  AOI21_X1   g11269(.A1(new_n11461_), .A2(\asqrt[38] ), .B(new_n11259_), .ZN(new_n11462_));
  NOR2_X1    g11270(.A1(new_n11462_), .A2(new_n11460_), .ZN(new_n11463_));
  AOI22_X1   g11271(.A1(new_n11461_), .A2(\asqrt[38] ), .B1(new_n11459_), .B2(new_n11456_), .ZN(new_n11464_));
  INV_X1     g11272(.I(new_n11267_), .ZN(new_n11465_));
  OAI21_X1   g11273(.A1(new_n11464_), .A2(new_n4330_), .B(new_n11465_), .ZN(new_n11466_));
  NAND2_X1   g11274(.A1(new_n11466_), .A2(new_n11463_), .ZN(new_n11467_));
  OAI22_X1   g11275(.A1(new_n11464_), .A2(new_n4330_), .B1(new_n11462_), .B2(new_n11460_), .ZN(new_n11468_));
  AOI21_X1   g11276(.A1(new_n11468_), .A2(\asqrt[40] ), .B(new_n11274_), .ZN(new_n11469_));
  NOR2_X1    g11277(.A1(new_n11469_), .A2(new_n11467_), .ZN(new_n11470_));
  AOI22_X1   g11278(.A1(new_n11468_), .A2(\asqrt[40] ), .B1(new_n11466_), .B2(new_n11463_), .ZN(new_n11471_));
  INV_X1     g11279(.I(new_n11282_), .ZN(new_n11472_));
  OAI21_X1   g11280(.A1(new_n11471_), .A2(new_n3760_), .B(new_n11472_), .ZN(new_n11473_));
  NAND2_X1   g11281(.A1(new_n11473_), .A2(new_n11470_), .ZN(new_n11474_));
  OAI22_X1   g11282(.A1(new_n11471_), .A2(new_n3760_), .B1(new_n11469_), .B2(new_n11467_), .ZN(new_n11475_));
  AOI21_X1   g11283(.A1(new_n11475_), .A2(\asqrt[42] ), .B(new_n11289_), .ZN(new_n11476_));
  NOR2_X1    g11284(.A1(new_n11476_), .A2(new_n11474_), .ZN(new_n11477_));
  AOI22_X1   g11285(.A1(new_n11475_), .A2(\asqrt[42] ), .B1(new_n11473_), .B2(new_n11470_), .ZN(new_n11478_));
  INV_X1     g11286(.I(new_n11297_), .ZN(new_n11479_));
  OAI21_X1   g11287(.A1(new_n11478_), .A2(new_n3208_), .B(new_n11479_), .ZN(new_n11480_));
  NAND2_X1   g11288(.A1(new_n11480_), .A2(new_n11477_), .ZN(new_n11481_));
  OAI22_X1   g11289(.A1(new_n11478_), .A2(new_n3208_), .B1(new_n11476_), .B2(new_n11474_), .ZN(new_n11482_));
  AOI21_X1   g11290(.A1(new_n11482_), .A2(\asqrt[44] ), .B(new_n11304_), .ZN(new_n11483_));
  NOR2_X1    g11291(.A1(new_n11483_), .A2(new_n11481_), .ZN(new_n11484_));
  AOI22_X1   g11292(.A1(new_n11482_), .A2(\asqrt[44] ), .B1(new_n11480_), .B2(new_n11477_), .ZN(new_n11485_));
  INV_X1     g11293(.I(new_n11312_), .ZN(new_n11486_));
  OAI21_X1   g11294(.A1(new_n11485_), .A2(new_n2728_), .B(new_n11486_), .ZN(new_n11487_));
  NAND2_X1   g11295(.A1(new_n11487_), .A2(new_n11484_), .ZN(new_n11488_));
  OAI22_X1   g11296(.A1(new_n11485_), .A2(new_n2728_), .B1(new_n11483_), .B2(new_n11481_), .ZN(new_n11489_));
  AOI21_X1   g11297(.A1(new_n11489_), .A2(\asqrt[46] ), .B(new_n11319_), .ZN(new_n11490_));
  NOR2_X1    g11298(.A1(new_n11490_), .A2(new_n11488_), .ZN(new_n11491_));
  AOI22_X1   g11299(.A1(new_n11489_), .A2(\asqrt[46] ), .B1(new_n11487_), .B2(new_n11484_), .ZN(new_n11492_));
  INV_X1     g11300(.I(new_n11327_), .ZN(new_n11493_));
  OAI21_X1   g11301(.A1(new_n11492_), .A2(new_n2253_), .B(new_n11493_), .ZN(new_n11494_));
  NAND2_X1   g11302(.A1(new_n11494_), .A2(new_n11491_), .ZN(new_n11495_));
  OAI22_X1   g11303(.A1(new_n11492_), .A2(new_n2253_), .B1(new_n11490_), .B2(new_n11488_), .ZN(new_n11496_));
  AOI21_X1   g11304(.A1(new_n11496_), .A2(\asqrt[48] ), .B(new_n11334_), .ZN(new_n11497_));
  NOR2_X1    g11305(.A1(new_n11497_), .A2(new_n11495_), .ZN(new_n11498_));
  AOI22_X1   g11306(.A1(new_n11496_), .A2(\asqrt[48] ), .B1(new_n11494_), .B2(new_n11491_), .ZN(new_n11499_));
  INV_X1     g11307(.I(new_n11342_), .ZN(new_n11500_));
  OAI21_X1   g11308(.A1(new_n11499_), .A2(new_n1854_), .B(new_n11500_), .ZN(new_n11501_));
  NAND2_X1   g11309(.A1(new_n11501_), .A2(new_n11498_), .ZN(new_n11502_));
  OAI22_X1   g11310(.A1(new_n11499_), .A2(new_n1854_), .B1(new_n11497_), .B2(new_n11495_), .ZN(new_n11503_));
  AOI21_X1   g11311(.A1(new_n11503_), .A2(\asqrt[50] ), .B(new_n11349_), .ZN(new_n11504_));
  NOR2_X1    g11312(.A1(new_n11504_), .A2(new_n11502_), .ZN(new_n11505_));
  AOI22_X1   g11313(.A1(new_n11503_), .A2(\asqrt[50] ), .B1(new_n11501_), .B2(new_n11498_), .ZN(new_n11506_));
  INV_X1     g11314(.I(new_n11357_), .ZN(new_n11507_));
  OAI21_X1   g11315(.A1(new_n11506_), .A2(new_n1436_), .B(new_n11507_), .ZN(new_n11508_));
  NAND2_X1   g11316(.A1(new_n11508_), .A2(new_n11505_), .ZN(new_n11509_));
  OAI22_X1   g11317(.A1(new_n11506_), .A2(new_n1436_), .B1(new_n11504_), .B2(new_n11502_), .ZN(new_n11510_));
  AOI21_X1   g11318(.A1(new_n11510_), .A2(\asqrt[52] ), .B(new_n11364_), .ZN(new_n11511_));
  NOR2_X1    g11319(.A1(new_n11511_), .A2(new_n11509_), .ZN(new_n11512_));
  AOI22_X1   g11320(.A1(new_n11510_), .A2(\asqrt[52] ), .B1(new_n11508_), .B2(new_n11505_), .ZN(new_n11513_));
  INV_X1     g11321(.I(new_n11372_), .ZN(new_n11514_));
  OAI21_X1   g11322(.A1(new_n11513_), .A2(new_n1096_), .B(new_n11514_), .ZN(new_n11515_));
  NAND2_X1   g11323(.A1(new_n11515_), .A2(new_n11512_), .ZN(new_n11516_));
  OAI22_X1   g11324(.A1(new_n11513_), .A2(new_n1096_), .B1(new_n11511_), .B2(new_n11509_), .ZN(new_n11517_));
  AOI21_X1   g11325(.A1(new_n11517_), .A2(\asqrt[54] ), .B(new_n11379_), .ZN(new_n11518_));
  NOR2_X1    g11326(.A1(new_n11518_), .A2(new_n11516_), .ZN(new_n11519_));
  AOI22_X1   g11327(.A1(new_n11517_), .A2(\asqrt[54] ), .B1(new_n11515_), .B2(new_n11512_), .ZN(new_n11520_));
  INV_X1     g11328(.I(new_n11387_), .ZN(new_n11521_));
  OAI21_X1   g11329(.A1(new_n11520_), .A2(new_n825_), .B(new_n11521_), .ZN(new_n11522_));
  NAND2_X1   g11330(.A1(new_n11522_), .A2(new_n11519_), .ZN(new_n11523_));
  OAI22_X1   g11331(.A1(new_n11520_), .A2(new_n825_), .B1(new_n11518_), .B2(new_n11516_), .ZN(new_n11524_));
  AOI21_X1   g11332(.A1(new_n11524_), .A2(\asqrt[56] ), .B(new_n11394_), .ZN(new_n11525_));
  NOR2_X1    g11333(.A1(new_n11525_), .A2(new_n11523_), .ZN(new_n11526_));
  AOI22_X1   g11334(.A1(new_n11524_), .A2(\asqrt[56] ), .B1(new_n11522_), .B2(new_n11519_), .ZN(new_n11527_));
  OAI21_X1   g11335(.A1(new_n11527_), .A2(new_n587_), .B(new_n11406_), .ZN(new_n11528_));
  NAND2_X1   g11336(.A1(new_n11528_), .A2(new_n11526_), .ZN(new_n11529_));
  NAND2_X1   g11337(.A1(new_n11517_), .A2(\asqrt[54] ), .ZN(new_n11530_));
  AOI21_X1   g11338(.A1(new_n11530_), .A2(new_n11516_), .B(new_n825_), .ZN(new_n11531_));
  OAI21_X1   g11339(.A1(new_n11519_), .A2(new_n11531_), .B(\asqrt[56] ), .ZN(new_n11532_));
  AOI21_X1   g11340(.A1(new_n11523_), .A2(new_n11532_), .B(new_n587_), .ZN(new_n11533_));
  OAI21_X1   g11341(.A1(new_n11526_), .A2(new_n11533_), .B(\asqrt[58] ), .ZN(new_n11534_));
  NAND2_X1   g11342(.A1(new_n11529_), .A2(new_n11534_), .ZN(new_n11535_));
  AOI22_X1   g11343(.A1(new_n11535_), .A2(\asqrt[59] ), .B1(new_n11414_), .B2(new_n11407_), .ZN(new_n11536_));
  NOR4_X1    g11344(.A1(new_n11105_), .A2(\asqrt[60] ), .A3(new_n10883_), .A4(new_n11030_), .ZN(new_n11537_));
  XOR2_X1    g11345(.A1(new_n11537_), .A2(new_n11071_), .Z(new_n11538_));
  NAND2_X1   g11346(.A1(new_n11538_), .A2(new_n229_), .ZN(new_n11539_));
  INV_X1     g11347(.I(new_n11539_), .ZN(new_n11540_));
  OAI21_X1   g11348(.A1(new_n11536_), .A2(new_n275_), .B(new_n11540_), .ZN(new_n11541_));
  OAI22_X1   g11349(.A1(new_n11527_), .A2(new_n587_), .B1(new_n11525_), .B2(new_n11523_), .ZN(new_n11542_));
  AOI21_X1   g11350(.A1(new_n11542_), .A2(\asqrt[58] ), .B(new_n11412_), .ZN(new_n11543_));
  NOR2_X1    g11351(.A1(new_n11543_), .A2(new_n11529_), .ZN(new_n11544_));
  AOI22_X1   g11352(.A1(new_n11542_), .A2(\asqrt[58] ), .B1(new_n11528_), .B2(new_n11526_), .ZN(new_n11545_));
  OAI21_X1   g11353(.A1(new_n11545_), .A2(new_n376_), .B(new_n11420_), .ZN(new_n11546_));
  NAND2_X1   g11354(.A1(new_n11546_), .A2(new_n11544_), .ZN(new_n11547_));
  AOI21_X1   g11355(.A1(new_n11529_), .A2(new_n11534_), .B(new_n376_), .ZN(new_n11548_));
  OAI21_X1   g11356(.A1(new_n11544_), .A2(new_n11548_), .B(\asqrt[60] ), .ZN(new_n11549_));
  AOI21_X1   g11357(.A1(new_n11547_), .A2(new_n11549_), .B(new_n229_), .ZN(new_n11550_));
  INV_X1     g11358(.I(new_n11075_), .ZN(new_n11551_));
  NOR2_X1    g11359(.A1(new_n11551_), .A2(\asqrt[62] ), .ZN(new_n11552_));
  INV_X1     g11360(.I(new_n11552_), .ZN(new_n11553_));
  NAND4_X1   g11361(.A1(new_n11550_), .A2(new_n11421_), .A3(new_n11541_), .A4(new_n11553_), .ZN(new_n11554_));
  NAND2_X1   g11362(.A1(new_n11093_), .A2(new_n11041_), .ZN(new_n11555_));
  OAI21_X1   g11363(.A1(\asqrt[22] ), .A2(new_n11555_), .B(new_n11053_), .ZN(new_n11556_));
  NAND2_X1   g11364(.A1(new_n11556_), .A2(new_n231_), .ZN(new_n11557_));
  INV_X1     g11365(.I(new_n11557_), .ZN(new_n11558_));
  NAND3_X1   g11366(.A1(new_n11554_), .A2(new_n11077_), .A3(new_n11558_), .ZN(new_n11559_));
  OAI22_X1   g11367(.A1(new_n11545_), .A2(new_n376_), .B1(new_n11543_), .B2(new_n11529_), .ZN(new_n11560_));
  AOI21_X1   g11368(.A1(new_n11560_), .A2(\asqrt[60] ), .B(new_n11539_), .ZN(new_n11561_));
  AOI22_X1   g11369(.A1(new_n11560_), .A2(\asqrt[60] ), .B1(new_n11546_), .B2(new_n11544_), .ZN(new_n11562_));
  OAI22_X1   g11370(.A1(new_n11562_), .A2(new_n229_), .B1(new_n11561_), .B2(new_n11547_), .ZN(new_n11563_));
  NOR4_X1    g11371(.A1(new_n11563_), .A2(\asqrt[62] ), .A3(new_n11067_), .A4(new_n11075_), .ZN(new_n11564_));
  AOI21_X1   g11372(.A1(new_n11068_), .A2(new_n11559_), .B(new_n11564_), .ZN(new_n11565_));
  INV_X1     g11373(.I(\a[40] ), .ZN(new_n11566_));
  OAI21_X1   g11374(.A1(new_n11042_), .A2(new_n11053_), .B(\asqrt[22] ), .ZN(new_n11567_));
  XOR2_X1    g11375(.A1(new_n11053_), .A2(\asqrt[63] ), .Z(new_n11568_));
  NAND2_X1   g11376(.A1(new_n11567_), .A2(new_n11568_), .ZN(new_n11569_));
  INV_X1     g11377(.I(new_n11569_), .ZN(new_n11570_));
  NAND3_X1   g11378(.A1(new_n11099_), .A2(new_n11035_), .A3(new_n11042_), .ZN(new_n11571_));
  INV_X1     g11379(.I(new_n11571_), .ZN(new_n11572_));
  NOR2_X1    g11380(.A1(new_n11570_), .A2(new_n11572_), .ZN(new_n11573_));
  NOR2_X1    g11381(.A1(\a[38] ), .A2(\a[39] ), .ZN(new_n11574_));
  INV_X1     g11382(.I(new_n11574_), .ZN(new_n11575_));
  NOR3_X1    g11383(.A1(new_n11573_), .A2(new_n11566_), .A3(new_n11575_), .ZN(new_n11576_));
  NAND2_X1   g11384(.A1(new_n11565_), .A2(new_n11576_), .ZN(new_n11577_));
  XOR2_X1    g11385(.A1(new_n11577_), .A2(\a[41] ), .Z(new_n11578_));
  INV_X1     g11386(.I(\a[41] ), .ZN(new_n11579_));
  NAND2_X1   g11387(.A1(new_n11541_), .A2(new_n11421_), .ZN(new_n11580_));
  NAND2_X1   g11388(.A1(new_n11550_), .A2(new_n11553_), .ZN(new_n11581_));
  OAI21_X1   g11389(.A1(new_n11581_), .A2(new_n11580_), .B(new_n11077_), .ZN(new_n11582_));
  OAI21_X1   g11390(.A1(new_n11582_), .A2(new_n11557_), .B(new_n11068_), .ZN(new_n11583_));
  NAND2_X1   g11391(.A1(new_n11564_), .A2(new_n11570_), .ZN(new_n11584_));
  NOR2_X1    g11392(.A1(new_n11584_), .A2(new_n11583_), .ZN(new_n11585_));
  NAND3_X1   g11393(.A1(new_n11585_), .A2(new_n11068_), .A3(new_n11571_), .ZN(new_n11586_));
  NAND2_X1   g11394(.A1(new_n11547_), .A2(new_n11549_), .ZN(new_n11587_));
  AOI22_X1   g11395(.A1(new_n11587_), .A2(\asqrt[61] ), .B1(new_n11541_), .B2(new_n11421_), .ZN(new_n11588_));
  NOR2_X1    g11396(.A1(new_n11588_), .A2(new_n196_), .ZN(new_n11589_));
  AOI21_X1   g11397(.A1(new_n11415_), .A2(new_n11417_), .B(new_n275_), .ZN(new_n11590_));
  OAI21_X1   g11398(.A1(new_n11421_), .A2(new_n11590_), .B(\asqrt[61] ), .ZN(new_n11591_));
  NAND4_X1   g11399(.A1(new_n11580_), .A2(new_n196_), .A3(new_n11591_), .A4(new_n11551_), .ZN(new_n11592_));
  INV_X1     g11400(.I(new_n11592_), .ZN(new_n11593_));
  NOR3_X1    g11401(.A1(new_n11584_), .A2(new_n11583_), .A3(new_n11571_), .ZN(\asqrt[21] ));
  NAND3_X1   g11402(.A1(\asqrt[21] ), .A2(new_n11589_), .A3(new_n11593_), .ZN(new_n11595_));
  OAI21_X1   g11403(.A1(new_n11563_), .A2(\asqrt[62] ), .B(new_n11075_), .ZN(new_n11596_));
  OAI21_X1   g11404(.A1(\asqrt[21] ), .A2(new_n11596_), .B(new_n11589_), .ZN(new_n11597_));
  NAND2_X1   g11405(.A1(new_n11597_), .A2(new_n11595_), .ZN(new_n11598_));
  INV_X1     g11406(.I(new_n11598_), .ZN(new_n11599_));
  NOR3_X1    g11407(.A1(new_n11587_), .A2(\asqrt[61] ), .A3(new_n11538_), .ZN(new_n11600_));
  NAND2_X1   g11408(.A1(\asqrt[21] ), .A2(new_n11600_), .ZN(new_n11601_));
  XOR2_X1    g11409(.A1(new_n11601_), .A2(new_n11550_), .Z(new_n11602_));
  NOR2_X1    g11410(.A1(new_n11602_), .A2(new_n196_), .ZN(new_n11603_));
  INV_X1     g11411(.I(new_n11603_), .ZN(new_n11604_));
  INV_X1     g11412(.I(\a[42] ), .ZN(new_n11605_));
  NOR2_X1    g11413(.A1(\a[40] ), .A2(\a[41] ), .ZN(new_n11606_));
  INV_X1     g11414(.I(new_n11606_), .ZN(new_n11607_));
  NOR3_X1    g11415(.A1(new_n11106_), .A2(new_n11605_), .A3(new_n11607_), .ZN(new_n11608_));
  NAND3_X1   g11416(.A1(new_n11057_), .A2(new_n11093_), .A3(new_n11608_), .ZN(new_n11609_));
  XOR2_X1    g11417(.A1(new_n11609_), .A2(\a[43] ), .Z(new_n11610_));
  INV_X1     g11418(.I(\a[43] ), .ZN(new_n11611_));
  NOR4_X1    g11419(.A1(new_n11584_), .A2(new_n11583_), .A3(new_n11611_), .A4(new_n11571_), .ZN(new_n11612_));
  NOR2_X1    g11420(.A1(new_n11610_), .A2(\a[42] ), .ZN(new_n11613_));
  OAI21_X1   g11421(.A1(new_n11612_), .A2(new_n11613_), .B(new_n11610_), .ZN(new_n11614_));
  INV_X1     g11422(.I(new_n11610_), .ZN(new_n11615_));
  NOR2_X1    g11423(.A1(new_n11561_), .A2(new_n11547_), .ZN(new_n11616_));
  NOR3_X1    g11424(.A1(new_n11562_), .A2(new_n229_), .A3(new_n11552_), .ZN(new_n11617_));
  AOI21_X1   g11425(.A1(new_n11617_), .A2(new_n11616_), .B(new_n11076_), .ZN(new_n11618_));
  AOI21_X1   g11426(.A1(new_n11618_), .A2(new_n11558_), .B(new_n11067_), .ZN(new_n11619_));
  AOI21_X1   g11427(.A1(new_n11563_), .A2(\asqrt[62] ), .B(new_n11068_), .ZN(new_n11620_));
  NOR3_X1    g11428(.A1(new_n11620_), .A2(new_n11592_), .A3(new_n11569_), .ZN(new_n11621_));
  NAND4_X1   g11429(.A1(new_n11621_), .A2(\a[43] ), .A3(new_n11619_), .A4(new_n11572_), .ZN(new_n11622_));
  NAND3_X1   g11430(.A1(new_n11622_), .A2(\a[42] ), .A3(new_n11615_), .ZN(new_n11623_));
  NAND2_X1   g11431(.A1(new_n11614_), .A2(new_n11623_), .ZN(new_n11624_));
  NAND2_X1   g11432(.A1(new_n11091_), .A2(new_n11055_), .ZN(new_n11625_));
  NAND4_X1   g11433(.A1(new_n11095_), .A2(new_n11089_), .A3(new_n11042_), .A4(new_n11625_), .ZN(new_n11626_));
  NOR2_X1    g11434(.A1(new_n11105_), .A2(new_n11605_), .ZN(new_n11627_));
  XOR2_X1    g11435(.A1(new_n11627_), .A2(new_n11626_), .Z(new_n11628_));
  NOR2_X1    g11436(.A1(new_n11628_), .A2(new_n11607_), .ZN(new_n11629_));
  INV_X1     g11437(.I(new_n11629_), .ZN(new_n11630_));
  NAND3_X1   g11438(.A1(new_n11621_), .A2(new_n11619_), .A3(new_n11572_), .ZN(new_n11631_));
  NOR4_X1    g11439(.A1(new_n11591_), .A2(new_n11547_), .A3(new_n11561_), .A4(new_n11552_), .ZN(new_n11632_));
  NOR3_X1    g11440(.A1(new_n11632_), .A2(new_n11076_), .A3(new_n11557_), .ZN(new_n11633_));
  NAND4_X1   g11441(.A1(new_n11588_), .A2(new_n196_), .A3(new_n11068_), .A4(new_n11551_), .ZN(new_n11634_));
  OAI21_X1   g11442(.A1(new_n11633_), .A2(new_n11067_), .B(new_n11634_), .ZN(new_n11635_));
  NAND2_X1   g11443(.A1(new_n11573_), .A2(\asqrt[22] ), .ZN(new_n11636_));
  OAI21_X1   g11444(.A1(new_n11635_), .A2(new_n11636_), .B(new_n11078_), .ZN(new_n11637_));
  NAND3_X1   g11445(.A1(new_n11637_), .A2(new_n11079_), .A3(new_n11631_), .ZN(new_n11638_));
  INV_X1     g11446(.I(new_n11636_), .ZN(new_n11639_));
  AOI21_X1   g11447(.A1(new_n11565_), .A2(new_n11639_), .B(\a[44] ), .ZN(new_n11640_));
  OAI21_X1   g11448(.A1(new_n11640_), .A2(new_n11080_), .B(\asqrt[21] ), .ZN(new_n11641_));
  NAND4_X1   g11449(.A1(new_n11638_), .A2(new_n11641_), .A3(new_n10614_), .A4(new_n11630_), .ZN(new_n11642_));
  NAND2_X1   g11450(.A1(new_n11642_), .A2(new_n11624_), .ZN(new_n11643_));
  NAND3_X1   g11451(.A1(new_n11614_), .A2(new_n11623_), .A3(new_n11630_), .ZN(new_n11644_));
  AOI21_X1   g11452(.A1(\asqrt[22] ), .A2(new_n11078_), .B(\a[45] ), .ZN(new_n11645_));
  NOR2_X1    g11453(.A1(new_n11096_), .A2(\a[44] ), .ZN(new_n11646_));
  AOI21_X1   g11454(.A1(\asqrt[22] ), .A2(\a[44] ), .B(new_n11082_), .ZN(new_n11647_));
  OAI21_X1   g11455(.A1(new_n11645_), .A2(new_n11646_), .B(new_n11647_), .ZN(new_n11648_));
  INV_X1     g11456(.I(new_n11648_), .ZN(new_n11649_));
  NAND3_X1   g11457(.A1(\asqrt[21] ), .A2(new_n11104_), .A3(new_n11649_), .ZN(new_n11650_));
  OAI21_X1   g11458(.A1(new_n11631_), .A2(new_n11648_), .B(new_n11103_), .ZN(new_n11651_));
  NAND3_X1   g11459(.A1(new_n11650_), .A2(new_n11651_), .A3(new_n10104_), .ZN(new_n11652_));
  AOI21_X1   g11460(.A1(new_n11644_), .A2(\asqrt[23] ), .B(new_n11652_), .ZN(new_n11653_));
  NOR2_X1    g11461(.A1(new_n11643_), .A2(new_n11653_), .ZN(new_n11654_));
  AOI22_X1   g11462(.A1(new_n11642_), .A2(new_n11624_), .B1(\asqrt[23] ), .B2(new_n11644_), .ZN(new_n11655_));
  AOI21_X1   g11463(.A1(new_n11114_), .A2(new_n11111_), .B(\asqrt[24] ), .ZN(new_n11656_));
  AND4_X2    g11464(.A1(new_n11155_), .A2(\asqrt[21] ), .A3(new_n11136_), .A4(new_n11656_), .Z(new_n11657_));
  NOR2_X1    g11465(.A1(new_n11155_), .A2(new_n10104_), .ZN(new_n11658_));
  NOR3_X1    g11466(.A1(new_n11657_), .A2(\asqrt[25] ), .A3(new_n11658_), .ZN(new_n11659_));
  OAI21_X1   g11467(.A1(new_n11655_), .A2(new_n10104_), .B(new_n11659_), .ZN(new_n11660_));
  NAND2_X1   g11468(.A1(new_n11660_), .A2(new_n11654_), .ZN(new_n11661_));
  OAI22_X1   g11469(.A1(new_n11655_), .A2(new_n10104_), .B1(new_n11643_), .B2(new_n11653_), .ZN(new_n11662_));
  NAND2_X1   g11470(.A1(new_n11123_), .A2(new_n11124_), .ZN(new_n11663_));
  NAND4_X1   g11471(.A1(\asqrt[21] ), .A2(new_n9672_), .A3(new_n11663_), .A4(new_n11128_), .ZN(new_n11664_));
  XOR2_X1    g11472(.A1(new_n11664_), .A2(new_n11137_), .Z(new_n11665_));
  NAND2_X1   g11473(.A1(new_n11665_), .A2(new_n9212_), .ZN(new_n11666_));
  AOI21_X1   g11474(.A1(new_n11662_), .A2(\asqrt[25] ), .B(new_n11666_), .ZN(new_n11667_));
  NOR2_X1    g11475(.A1(new_n11667_), .A2(new_n11661_), .ZN(new_n11668_));
  AOI22_X1   g11476(.A1(new_n11662_), .A2(\asqrt[25] ), .B1(new_n11660_), .B2(new_n11654_), .ZN(new_n11669_));
  NOR4_X1    g11477(.A1(new_n11631_), .A2(\asqrt[26] ), .A3(new_n11132_), .A4(new_n11422_), .ZN(new_n11670_));
  XOR2_X1    g11478(.A1(new_n11670_), .A2(new_n11138_), .Z(new_n11671_));
  NAND2_X1   g11479(.A1(new_n11671_), .A2(new_n8763_), .ZN(new_n11672_));
  INV_X1     g11480(.I(new_n11672_), .ZN(new_n11673_));
  OAI21_X1   g11481(.A1(new_n11669_), .A2(new_n9212_), .B(new_n11673_), .ZN(new_n11674_));
  NAND2_X1   g11482(.A1(new_n11674_), .A2(new_n11668_), .ZN(new_n11675_));
  OAI22_X1   g11483(.A1(new_n11669_), .A2(new_n9212_), .B1(new_n11667_), .B2(new_n11661_), .ZN(new_n11676_));
  NOR4_X1    g11484(.A1(new_n11631_), .A2(\asqrt[27] ), .A3(new_n11142_), .A4(new_n11164_), .ZN(new_n11677_));
  XNOR2_X1   g11485(.A1(new_n11677_), .A2(new_n11174_), .ZN(new_n11678_));
  NAND2_X1   g11486(.A1(new_n11678_), .A2(new_n8319_), .ZN(new_n11679_));
  AOI21_X1   g11487(.A1(new_n11676_), .A2(\asqrt[27] ), .B(new_n11679_), .ZN(new_n11680_));
  NOR2_X1    g11488(.A1(new_n11680_), .A2(new_n11675_), .ZN(new_n11681_));
  AOI22_X1   g11489(.A1(new_n11676_), .A2(\asqrt[27] ), .B1(new_n11674_), .B2(new_n11668_), .ZN(new_n11682_));
  NOR4_X1    g11490(.A1(new_n11631_), .A2(\asqrt[28] ), .A3(new_n11168_), .A4(new_n11427_), .ZN(new_n11683_));
  XOR2_X1    g11491(.A1(new_n11683_), .A2(new_n11175_), .Z(new_n11684_));
  NAND2_X1   g11492(.A1(new_n11684_), .A2(new_n7931_), .ZN(new_n11685_));
  INV_X1     g11493(.I(new_n11685_), .ZN(new_n11686_));
  OAI21_X1   g11494(.A1(new_n11682_), .A2(new_n8319_), .B(new_n11686_), .ZN(new_n11687_));
  NAND2_X1   g11495(.A1(new_n11687_), .A2(new_n11681_), .ZN(new_n11688_));
  OAI22_X1   g11496(.A1(new_n11682_), .A2(new_n8319_), .B1(new_n11680_), .B2(new_n11675_), .ZN(new_n11689_));
  NOR4_X1    g11497(.A1(new_n11631_), .A2(\asqrt[29] ), .A3(new_n11178_), .A4(new_n11184_), .ZN(new_n11690_));
  XNOR2_X1   g11498(.A1(new_n11690_), .A2(new_n11193_), .ZN(new_n11691_));
  NAND2_X1   g11499(.A1(new_n11691_), .A2(new_n7517_), .ZN(new_n11692_));
  AOI21_X1   g11500(.A1(new_n11689_), .A2(\asqrt[29] ), .B(new_n11692_), .ZN(new_n11693_));
  NOR2_X1    g11501(.A1(new_n11693_), .A2(new_n11688_), .ZN(new_n11694_));
  AOI22_X1   g11502(.A1(new_n11689_), .A2(\asqrt[29] ), .B1(new_n11687_), .B2(new_n11681_), .ZN(new_n11695_));
  NOR4_X1    g11503(.A1(new_n11631_), .A2(\asqrt[30] ), .A3(new_n11187_), .A4(new_n11433_), .ZN(new_n11696_));
  XOR2_X1    g11504(.A1(new_n11696_), .A2(new_n11194_), .Z(new_n11697_));
  NAND2_X1   g11505(.A1(new_n11697_), .A2(new_n7110_), .ZN(new_n11698_));
  INV_X1     g11506(.I(new_n11698_), .ZN(new_n11699_));
  OAI21_X1   g11507(.A1(new_n11695_), .A2(new_n7517_), .B(new_n11699_), .ZN(new_n11700_));
  NAND2_X1   g11508(.A1(new_n11700_), .A2(new_n11694_), .ZN(new_n11701_));
  OAI22_X1   g11509(.A1(new_n11695_), .A2(new_n7517_), .B1(new_n11693_), .B2(new_n11688_), .ZN(new_n11702_));
  NAND2_X1   g11510(.A1(new_n11203_), .A2(\asqrt[31] ), .ZN(new_n11703_));
  NOR4_X1    g11511(.A1(new_n11631_), .A2(\asqrt[31] ), .A3(new_n11197_), .A4(new_n11203_), .ZN(new_n11704_));
  XOR2_X1    g11512(.A1(new_n11704_), .A2(new_n11703_), .Z(new_n11705_));
  NAND2_X1   g11513(.A1(new_n11705_), .A2(new_n6708_), .ZN(new_n11706_));
  AOI21_X1   g11514(.A1(new_n11702_), .A2(\asqrt[31] ), .B(new_n11706_), .ZN(new_n11707_));
  NOR2_X1    g11515(.A1(new_n11707_), .A2(new_n11701_), .ZN(new_n11708_));
  AOI22_X1   g11516(.A1(new_n11702_), .A2(\asqrt[31] ), .B1(new_n11700_), .B2(new_n11694_), .ZN(new_n11709_));
  NOR4_X1    g11517(.A1(new_n11631_), .A2(\asqrt[32] ), .A3(new_n11206_), .A4(new_n11440_), .ZN(new_n11710_));
  AOI21_X1   g11518(.A1(new_n11703_), .A2(new_n11201_), .B(new_n6708_), .ZN(new_n11711_));
  NOR2_X1    g11519(.A1(new_n11710_), .A2(new_n11711_), .ZN(new_n11712_));
  NAND2_X1   g11520(.A1(new_n11712_), .A2(new_n6365_), .ZN(new_n11713_));
  INV_X1     g11521(.I(new_n11713_), .ZN(new_n11714_));
  OAI21_X1   g11522(.A1(new_n11709_), .A2(new_n6708_), .B(new_n11714_), .ZN(new_n11715_));
  NAND2_X1   g11523(.A1(new_n11715_), .A2(new_n11708_), .ZN(new_n11716_));
  OAI22_X1   g11524(.A1(new_n11709_), .A2(new_n6708_), .B1(new_n11707_), .B2(new_n11701_), .ZN(new_n11717_));
  NAND2_X1   g11525(.A1(new_n11218_), .A2(\asqrt[33] ), .ZN(new_n11718_));
  NOR4_X1    g11526(.A1(new_n11631_), .A2(\asqrt[33] ), .A3(new_n11213_), .A4(new_n11218_), .ZN(new_n11719_));
  XOR2_X1    g11527(.A1(new_n11719_), .A2(new_n11718_), .Z(new_n11720_));
  NAND2_X1   g11528(.A1(new_n11720_), .A2(new_n5991_), .ZN(new_n11721_));
  AOI21_X1   g11529(.A1(new_n11717_), .A2(\asqrt[33] ), .B(new_n11721_), .ZN(new_n11722_));
  NOR2_X1    g11530(.A1(new_n11722_), .A2(new_n11716_), .ZN(new_n11723_));
  AOI22_X1   g11531(.A1(new_n11717_), .A2(\asqrt[33] ), .B1(new_n11715_), .B2(new_n11708_), .ZN(new_n11724_));
  NOR4_X1    g11532(.A1(new_n11631_), .A2(\asqrt[34] ), .A3(new_n11221_), .A4(new_n11447_), .ZN(new_n11725_));
  AOI21_X1   g11533(.A1(new_n11718_), .A2(new_n11217_), .B(new_n5991_), .ZN(new_n11726_));
  NOR2_X1    g11534(.A1(new_n11725_), .A2(new_n11726_), .ZN(new_n11727_));
  NAND2_X1   g11535(.A1(new_n11727_), .A2(new_n5626_), .ZN(new_n11728_));
  INV_X1     g11536(.I(new_n11728_), .ZN(new_n11729_));
  OAI21_X1   g11537(.A1(new_n11724_), .A2(new_n5991_), .B(new_n11729_), .ZN(new_n11730_));
  NAND2_X1   g11538(.A1(new_n11730_), .A2(new_n11723_), .ZN(new_n11731_));
  OAI22_X1   g11539(.A1(new_n11724_), .A2(new_n5991_), .B1(new_n11722_), .B2(new_n11716_), .ZN(new_n11732_));
  NAND2_X1   g11540(.A1(new_n11233_), .A2(\asqrt[35] ), .ZN(new_n11733_));
  NOR4_X1    g11541(.A1(new_n11631_), .A2(\asqrt[35] ), .A3(new_n11228_), .A4(new_n11233_), .ZN(new_n11734_));
  XOR2_X1    g11542(.A1(new_n11734_), .A2(new_n11733_), .Z(new_n11735_));
  NAND2_X1   g11543(.A1(new_n11735_), .A2(new_n5273_), .ZN(new_n11736_));
  AOI21_X1   g11544(.A1(new_n11732_), .A2(\asqrt[35] ), .B(new_n11736_), .ZN(new_n11737_));
  NOR2_X1    g11545(.A1(new_n11737_), .A2(new_n11731_), .ZN(new_n11738_));
  AOI22_X1   g11546(.A1(new_n11732_), .A2(\asqrt[35] ), .B1(new_n11730_), .B2(new_n11723_), .ZN(new_n11739_));
  NOR4_X1    g11547(.A1(new_n11631_), .A2(\asqrt[36] ), .A3(new_n11236_), .A4(new_n11454_), .ZN(new_n11740_));
  AOI21_X1   g11548(.A1(new_n11733_), .A2(new_n11232_), .B(new_n5273_), .ZN(new_n11741_));
  NOR2_X1    g11549(.A1(new_n11740_), .A2(new_n11741_), .ZN(new_n11742_));
  NAND2_X1   g11550(.A1(new_n11742_), .A2(new_n4973_), .ZN(new_n11743_));
  INV_X1     g11551(.I(new_n11743_), .ZN(new_n11744_));
  OAI21_X1   g11552(.A1(new_n11739_), .A2(new_n5273_), .B(new_n11744_), .ZN(new_n11745_));
  NAND2_X1   g11553(.A1(new_n11745_), .A2(new_n11738_), .ZN(new_n11746_));
  OAI22_X1   g11554(.A1(new_n11739_), .A2(new_n5273_), .B1(new_n11737_), .B2(new_n11731_), .ZN(new_n11747_));
  NAND2_X1   g11555(.A1(new_n11248_), .A2(\asqrt[37] ), .ZN(new_n11748_));
  NOR4_X1    g11556(.A1(new_n11631_), .A2(\asqrt[37] ), .A3(new_n11243_), .A4(new_n11248_), .ZN(new_n11749_));
  XOR2_X1    g11557(.A1(new_n11749_), .A2(new_n11748_), .Z(new_n11750_));
  NAND2_X1   g11558(.A1(new_n11750_), .A2(new_n4645_), .ZN(new_n11751_));
  AOI21_X1   g11559(.A1(new_n11747_), .A2(\asqrt[37] ), .B(new_n11751_), .ZN(new_n11752_));
  NOR2_X1    g11560(.A1(new_n11752_), .A2(new_n11746_), .ZN(new_n11753_));
  AOI22_X1   g11561(.A1(new_n11747_), .A2(\asqrt[37] ), .B1(new_n11745_), .B2(new_n11738_), .ZN(new_n11754_));
  NOR4_X1    g11562(.A1(new_n11631_), .A2(\asqrt[38] ), .A3(new_n11251_), .A4(new_n11461_), .ZN(new_n11755_));
  AOI21_X1   g11563(.A1(new_n11748_), .A2(new_n11247_), .B(new_n4645_), .ZN(new_n11756_));
  NOR2_X1    g11564(.A1(new_n11755_), .A2(new_n11756_), .ZN(new_n11757_));
  NAND2_X1   g11565(.A1(new_n11757_), .A2(new_n4330_), .ZN(new_n11758_));
  INV_X1     g11566(.I(new_n11758_), .ZN(new_n11759_));
  OAI21_X1   g11567(.A1(new_n11754_), .A2(new_n4645_), .B(new_n11759_), .ZN(new_n11760_));
  NAND2_X1   g11568(.A1(new_n11760_), .A2(new_n11753_), .ZN(new_n11761_));
  OAI22_X1   g11569(.A1(new_n11754_), .A2(new_n4645_), .B1(new_n11752_), .B2(new_n11746_), .ZN(new_n11762_));
  NAND2_X1   g11570(.A1(new_n11263_), .A2(\asqrt[39] ), .ZN(new_n11763_));
  NOR4_X1    g11571(.A1(new_n11631_), .A2(\asqrt[39] ), .A3(new_n11258_), .A4(new_n11263_), .ZN(new_n11764_));
  XOR2_X1    g11572(.A1(new_n11764_), .A2(new_n11763_), .Z(new_n11765_));
  NAND2_X1   g11573(.A1(new_n11765_), .A2(new_n4018_), .ZN(new_n11766_));
  AOI21_X1   g11574(.A1(new_n11762_), .A2(\asqrt[39] ), .B(new_n11766_), .ZN(new_n11767_));
  NOR2_X1    g11575(.A1(new_n11767_), .A2(new_n11761_), .ZN(new_n11768_));
  AOI22_X1   g11576(.A1(new_n11762_), .A2(\asqrt[39] ), .B1(new_n11760_), .B2(new_n11753_), .ZN(new_n11769_));
  NOR4_X1    g11577(.A1(new_n11631_), .A2(\asqrt[40] ), .A3(new_n11266_), .A4(new_n11468_), .ZN(new_n11770_));
  AOI21_X1   g11578(.A1(new_n11763_), .A2(new_n11262_), .B(new_n4018_), .ZN(new_n11771_));
  NOR2_X1    g11579(.A1(new_n11770_), .A2(new_n11771_), .ZN(new_n11772_));
  NAND2_X1   g11580(.A1(new_n11772_), .A2(new_n3760_), .ZN(new_n11773_));
  INV_X1     g11581(.I(new_n11773_), .ZN(new_n11774_));
  OAI21_X1   g11582(.A1(new_n11769_), .A2(new_n4018_), .B(new_n11774_), .ZN(new_n11775_));
  NAND2_X1   g11583(.A1(new_n11775_), .A2(new_n11768_), .ZN(new_n11776_));
  OAI22_X1   g11584(.A1(new_n11769_), .A2(new_n4018_), .B1(new_n11767_), .B2(new_n11761_), .ZN(new_n11777_));
  NAND2_X1   g11585(.A1(new_n11278_), .A2(\asqrt[41] ), .ZN(new_n11778_));
  NOR4_X1    g11586(.A1(new_n11631_), .A2(\asqrt[41] ), .A3(new_n11273_), .A4(new_n11278_), .ZN(new_n11779_));
  XOR2_X1    g11587(.A1(new_n11779_), .A2(new_n11778_), .Z(new_n11780_));
  NAND2_X1   g11588(.A1(new_n11780_), .A2(new_n3481_), .ZN(new_n11781_));
  AOI21_X1   g11589(.A1(new_n11777_), .A2(\asqrt[41] ), .B(new_n11781_), .ZN(new_n11782_));
  NOR2_X1    g11590(.A1(new_n11782_), .A2(new_n11776_), .ZN(new_n11783_));
  AOI22_X1   g11591(.A1(new_n11777_), .A2(\asqrt[41] ), .B1(new_n11775_), .B2(new_n11768_), .ZN(new_n11784_));
  NAND2_X1   g11592(.A1(new_n11475_), .A2(\asqrt[42] ), .ZN(new_n11785_));
  NOR4_X1    g11593(.A1(new_n11631_), .A2(\asqrt[42] ), .A3(new_n11281_), .A4(new_n11475_), .ZN(new_n11786_));
  XOR2_X1    g11594(.A1(new_n11786_), .A2(new_n11785_), .Z(new_n11787_));
  NAND2_X1   g11595(.A1(new_n11787_), .A2(new_n3208_), .ZN(new_n11788_));
  INV_X1     g11596(.I(new_n11788_), .ZN(new_n11789_));
  OAI21_X1   g11597(.A1(new_n11784_), .A2(new_n3481_), .B(new_n11789_), .ZN(new_n11790_));
  NAND2_X1   g11598(.A1(new_n11790_), .A2(new_n11783_), .ZN(new_n11791_));
  OAI22_X1   g11599(.A1(new_n11784_), .A2(new_n3481_), .B1(new_n11782_), .B2(new_n11776_), .ZN(new_n11792_));
  NOR4_X1    g11600(.A1(new_n11631_), .A2(\asqrt[43] ), .A3(new_n11288_), .A4(new_n11293_), .ZN(new_n11793_));
  AOI21_X1   g11601(.A1(new_n11785_), .A2(new_n11474_), .B(new_n3208_), .ZN(new_n11794_));
  NOR2_X1    g11602(.A1(new_n11793_), .A2(new_n11794_), .ZN(new_n11795_));
  NAND2_X1   g11603(.A1(new_n11795_), .A2(new_n2941_), .ZN(new_n11796_));
  AOI21_X1   g11604(.A1(new_n11792_), .A2(\asqrt[43] ), .B(new_n11796_), .ZN(new_n11797_));
  NOR2_X1    g11605(.A1(new_n11797_), .A2(new_n11791_), .ZN(new_n11798_));
  AOI22_X1   g11606(.A1(new_n11792_), .A2(\asqrt[43] ), .B1(new_n11790_), .B2(new_n11783_), .ZN(new_n11799_));
  NAND2_X1   g11607(.A1(new_n11482_), .A2(\asqrt[44] ), .ZN(new_n11800_));
  NOR4_X1    g11608(.A1(new_n11631_), .A2(\asqrt[44] ), .A3(new_n11296_), .A4(new_n11482_), .ZN(new_n11801_));
  XOR2_X1    g11609(.A1(new_n11801_), .A2(new_n11800_), .Z(new_n11802_));
  NAND2_X1   g11610(.A1(new_n11802_), .A2(new_n2728_), .ZN(new_n11803_));
  INV_X1     g11611(.I(new_n11803_), .ZN(new_n11804_));
  OAI21_X1   g11612(.A1(new_n11799_), .A2(new_n2941_), .B(new_n11804_), .ZN(new_n11805_));
  NAND2_X1   g11613(.A1(new_n11805_), .A2(new_n11798_), .ZN(new_n11806_));
  OAI22_X1   g11614(.A1(new_n11799_), .A2(new_n2941_), .B1(new_n11797_), .B2(new_n11791_), .ZN(new_n11807_));
  NOR4_X1    g11615(.A1(new_n11631_), .A2(\asqrt[45] ), .A3(new_n11303_), .A4(new_n11308_), .ZN(new_n11808_));
  AOI21_X1   g11616(.A1(new_n11800_), .A2(new_n11481_), .B(new_n2728_), .ZN(new_n11809_));
  NOR2_X1    g11617(.A1(new_n11808_), .A2(new_n11809_), .ZN(new_n11810_));
  NAND2_X1   g11618(.A1(new_n11810_), .A2(new_n2488_), .ZN(new_n11811_));
  AOI21_X1   g11619(.A1(new_n11807_), .A2(\asqrt[45] ), .B(new_n11811_), .ZN(new_n11812_));
  NOR2_X1    g11620(.A1(new_n11812_), .A2(new_n11806_), .ZN(new_n11813_));
  AOI22_X1   g11621(.A1(new_n11807_), .A2(\asqrt[45] ), .B1(new_n11805_), .B2(new_n11798_), .ZN(new_n11814_));
  NAND2_X1   g11622(.A1(new_n11489_), .A2(\asqrt[46] ), .ZN(new_n11815_));
  NOR4_X1    g11623(.A1(new_n11631_), .A2(\asqrt[46] ), .A3(new_n11311_), .A4(new_n11489_), .ZN(new_n11816_));
  XOR2_X1    g11624(.A1(new_n11816_), .A2(new_n11815_), .Z(new_n11817_));
  NAND2_X1   g11625(.A1(new_n11817_), .A2(new_n2253_), .ZN(new_n11818_));
  INV_X1     g11626(.I(new_n11818_), .ZN(new_n11819_));
  OAI21_X1   g11627(.A1(new_n11814_), .A2(new_n2488_), .B(new_n11819_), .ZN(new_n11820_));
  NAND2_X1   g11628(.A1(new_n11820_), .A2(new_n11813_), .ZN(new_n11821_));
  OAI22_X1   g11629(.A1(new_n11814_), .A2(new_n2488_), .B1(new_n11812_), .B2(new_n11806_), .ZN(new_n11822_));
  NAND2_X1   g11630(.A1(new_n11323_), .A2(\asqrt[47] ), .ZN(new_n11823_));
  NOR4_X1    g11631(.A1(new_n11631_), .A2(\asqrt[47] ), .A3(new_n11318_), .A4(new_n11323_), .ZN(new_n11824_));
  XOR2_X1    g11632(.A1(new_n11824_), .A2(new_n11823_), .Z(new_n11825_));
  NAND2_X1   g11633(.A1(new_n11825_), .A2(new_n2046_), .ZN(new_n11826_));
  AOI21_X1   g11634(.A1(new_n11822_), .A2(\asqrt[47] ), .B(new_n11826_), .ZN(new_n11827_));
  NOR2_X1    g11635(.A1(new_n11827_), .A2(new_n11821_), .ZN(new_n11828_));
  AOI22_X1   g11636(.A1(new_n11822_), .A2(\asqrt[47] ), .B1(new_n11820_), .B2(new_n11813_), .ZN(new_n11829_));
  NOR4_X1    g11637(.A1(new_n11631_), .A2(\asqrt[48] ), .A3(new_n11326_), .A4(new_n11496_), .ZN(new_n11830_));
  AOI21_X1   g11638(.A1(new_n11823_), .A2(new_n11322_), .B(new_n2046_), .ZN(new_n11831_));
  NOR2_X1    g11639(.A1(new_n11830_), .A2(new_n11831_), .ZN(new_n11832_));
  NAND2_X1   g11640(.A1(new_n11832_), .A2(new_n1854_), .ZN(new_n11833_));
  INV_X1     g11641(.I(new_n11833_), .ZN(new_n11834_));
  OAI21_X1   g11642(.A1(new_n11829_), .A2(new_n2046_), .B(new_n11834_), .ZN(new_n11835_));
  NAND2_X1   g11643(.A1(new_n11835_), .A2(new_n11828_), .ZN(new_n11836_));
  OAI22_X1   g11644(.A1(new_n11829_), .A2(new_n2046_), .B1(new_n11827_), .B2(new_n11821_), .ZN(new_n11837_));
  NAND2_X1   g11645(.A1(new_n11338_), .A2(\asqrt[49] ), .ZN(new_n11838_));
  NOR4_X1    g11646(.A1(new_n11631_), .A2(\asqrt[49] ), .A3(new_n11333_), .A4(new_n11338_), .ZN(new_n11839_));
  XOR2_X1    g11647(.A1(new_n11839_), .A2(new_n11838_), .Z(new_n11840_));
  NAND2_X1   g11648(.A1(new_n11840_), .A2(new_n1595_), .ZN(new_n11841_));
  AOI21_X1   g11649(.A1(new_n11837_), .A2(\asqrt[49] ), .B(new_n11841_), .ZN(new_n11842_));
  NOR2_X1    g11650(.A1(new_n11842_), .A2(new_n11836_), .ZN(new_n11843_));
  AOI22_X1   g11651(.A1(new_n11837_), .A2(\asqrt[49] ), .B1(new_n11835_), .B2(new_n11828_), .ZN(new_n11844_));
  NOR4_X1    g11652(.A1(new_n11631_), .A2(\asqrt[50] ), .A3(new_n11341_), .A4(new_n11503_), .ZN(new_n11845_));
  AOI21_X1   g11653(.A1(new_n11838_), .A2(new_n11337_), .B(new_n1595_), .ZN(new_n11846_));
  NOR2_X1    g11654(.A1(new_n11845_), .A2(new_n11846_), .ZN(new_n11847_));
  NAND2_X1   g11655(.A1(new_n11847_), .A2(new_n1436_), .ZN(new_n11848_));
  INV_X1     g11656(.I(new_n11848_), .ZN(new_n11849_));
  OAI21_X1   g11657(.A1(new_n11844_), .A2(new_n1595_), .B(new_n11849_), .ZN(new_n11850_));
  NAND2_X1   g11658(.A1(new_n11850_), .A2(new_n11843_), .ZN(new_n11851_));
  OAI22_X1   g11659(.A1(new_n11844_), .A2(new_n1595_), .B1(new_n11842_), .B2(new_n11836_), .ZN(new_n11852_));
  NAND2_X1   g11660(.A1(new_n11353_), .A2(\asqrt[51] ), .ZN(new_n11853_));
  NOR4_X1    g11661(.A1(new_n11631_), .A2(\asqrt[51] ), .A3(new_n11348_), .A4(new_n11353_), .ZN(new_n11854_));
  XOR2_X1    g11662(.A1(new_n11854_), .A2(new_n11853_), .Z(new_n11855_));
  NAND2_X1   g11663(.A1(new_n11855_), .A2(new_n1260_), .ZN(new_n11856_));
  AOI21_X1   g11664(.A1(new_n11852_), .A2(\asqrt[51] ), .B(new_n11856_), .ZN(new_n11857_));
  NOR2_X1    g11665(.A1(new_n11857_), .A2(new_n11851_), .ZN(new_n11858_));
  AOI22_X1   g11666(.A1(new_n11852_), .A2(\asqrt[51] ), .B1(new_n11850_), .B2(new_n11843_), .ZN(new_n11859_));
  NOR4_X1    g11667(.A1(new_n11631_), .A2(\asqrt[52] ), .A3(new_n11356_), .A4(new_n11510_), .ZN(new_n11860_));
  AOI21_X1   g11668(.A1(new_n11853_), .A2(new_n11352_), .B(new_n1260_), .ZN(new_n11861_));
  NOR2_X1    g11669(.A1(new_n11860_), .A2(new_n11861_), .ZN(new_n11862_));
  NAND2_X1   g11670(.A1(new_n11862_), .A2(new_n1096_), .ZN(new_n11863_));
  INV_X1     g11671(.I(new_n11863_), .ZN(new_n11864_));
  OAI21_X1   g11672(.A1(new_n11859_), .A2(new_n1260_), .B(new_n11864_), .ZN(new_n11865_));
  NAND2_X1   g11673(.A1(new_n11865_), .A2(new_n11858_), .ZN(new_n11866_));
  OAI22_X1   g11674(.A1(new_n11859_), .A2(new_n1260_), .B1(new_n11857_), .B2(new_n11851_), .ZN(new_n11867_));
  NOR4_X1    g11675(.A1(new_n11631_), .A2(\asqrt[53] ), .A3(new_n11363_), .A4(new_n11368_), .ZN(new_n11868_));
  XOR2_X1    g11676(.A1(new_n11868_), .A2(new_n11398_), .Z(new_n11869_));
  NAND2_X1   g11677(.A1(new_n11869_), .A2(new_n970_), .ZN(new_n11870_));
  AOI21_X1   g11678(.A1(new_n11867_), .A2(\asqrt[53] ), .B(new_n11870_), .ZN(new_n11871_));
  NOR2_X1    g11679(.A1(new_n11871_), .A2(new_n11866_), .ZN(new_n11872_));
  AOI22_X1   g11680(.A1(new_n11867_), .A2(\asqrt[53] ), .B1(new_n11865_), .B2(new_n11858_), .ZN(new_n11873_));
  NOR4_X1    g11681(.A1(new_n11631_), .A2(\asqrt[54] ), .A3(new_n11371_), .A4(new_n11517_), .ZN(new_n11874_));
  XOR2_X1    g11682(.A1(new_n11874_), .A2(new_n11530_), .Z(new_n11875_));
  NAND2_X1   g11683(.A1(new_n11875_), .A2(new_n825_), .ZN(new_n11876_));
  INV_X1     g11684(.I(new_n11876_), .ZN(new_n11877_));
  OAI21_X1   g11685(.A1(new_n11873_), .A2(new_n970_), .B(new_n11877_), .ZN(new_n11878_));
  NAND2_X1   g11686(.A1(new_n11878_), .A2(new_n11872_), .ZN(new_n11879_));
  OAI22_X1   g11687(.A1(new_n11873_), .A2(new_n970_), .B1(new_n11871_), .B2(new_n11866_), .ZN(new_n11880_));
  NOR4_X1    g11688(.A1(new_n11631_), .A2(\asqrt[55] ), .A3(new_n11378_), .A4(new_n11383_), .ZN(new_n11881_));
  XOR2_X1    g11689(.A1(new_n11881_), .A2(new_n11400_), .Z(new_n11882_));
  NAND2_X1   g11690(.A1(new_n11882_), .A2(new_n724_), .ZN(new_n11883_));
  AOI21_X1   g11691(.A1(new_n11880_), .A2(\asqrt[55] ), .B(new_n11883_), .ZN(new_n11884_));
  NOR2_X1    g11692(.A1(new_n11884_), .A2(new_n11879_), .ZN(new_n11885_));
  AOI22_X1   g11693(.A1(new_n11880_), .A2(\asqrt[55] ), .B1(new_n11878_), .B2(new_n11872_), .ZN(new_n11886_));
  NOR4_X1    g11694(.A1(new_n11631_), .A2(\asqrt[56] ), .A3(new_n11386_), .A4(new_n11524_), .ZN(new_n11887_));
  XOR2_X1    g11695(.A1(new_n11887_), .A2(new_n11532_), .Z(new_n11888_));
  NAND2_X1   g11696(.A1(new_n11888_), .A2(new_n587_), .ZN(new_n11889_));
  INV_X1     g11697(.I(new_n11889_), .ZN(new_n11890_));
  OAI21_X1   g11698(.A1(new_n11886_), .A2(new_n724_), .B(new_n11890_), .ZN(new_n11891_));
  NAND2_X1   g11699(.A1(new_n11891_), .A2(new_n11885_), .ZN(new_n11892_));
  OAI22_X1   g11700(.A1(new_n11886_), .A2(new_n724_), .B1(new_n11884_), .B2(new_n11879_), .ZN(new_n11893_));
  NOR4_X1    g11701(.A1(new_n11631_), .A2(\asqrt[57] ), .A3(new_n11393_), .A4(new_n11408_), .ZN(new_n11894_));
  XOR2_X1    g11702(.A1(new_n11894_), .A2(new_n11402_), .Z(new_n11895_));
  NAND2_X1   g11703(.A1(new_n11895_), .A2(new_n504_), .ZN(new_n11896_));
  AOI21_X1   g11704(.A1(new_n11893_), .A2(\asqrt[57] ), .B(new_n11896_), .ZN(new_n11897_));
  NOR2_X1    g11705(.A1(new_n11897_), .A2(new_n11892_), .ZN(new_n11898_));
  AOI22_X1   g11706(.A1(new_n11893_), .A2(\asqrt[57] ), .B1(new_n11891_), .B2(new_n11885_), .ZN(new_n11899_));
  NOR4_X1    g11707(.A1(new_n11631_), .A2(\asqrt[58] ), .A3(new_n11404_), .A4(new_n11542_), .ZN(new_n11900_));
  XOR2_X1    g11708(.A1(new_n11900_), .A2(new_n11534_), .Z(new_n11901_));
  NAND2_X1   g11709(.A1(new_n11901_), .A2(new_n376_), .ZN(new_n11902_));
  INV_X1     g11710(.I(new_n11902_), .ZN(new_n11903_));
  OAI21_X1   g11711(.A1(new_n11899_), .A2(new_n504_), .B(new_n11903_), .ZN(new_n11904_));
  NAND2_X1   g11712(.A1(new_n11904_), .A2(new_n11898_), .ZN(new_n11905_));
  OAI22_X1   g11713(.A1(new_n11899_), .A2(new_n504_), .B1(new_n11897_), .B2(new_n11892_), .ZN(new_n11906_));
  NOR4_X1    g11714(.A1(new_n11631_), .A2(\asqrt[59] ), .A3(new_n11411_), .A4(new_n11535_), .ZN(new_n11907_));
  XOR2_X1    g11715(.A1(new_n11907_), .A2(new_n11417_), .Z(new_n11908_));
  NAND2_X1   g11716(.A1(new_n11908_), .A2(new_n275_), .ZN(new_n11909_));
  AOI21_X1   g11717(.A1(new_n11906_), .A2(\asqrt[59] ), .B(new_n11909_), .ZN(new_n11910_));
  NOR2_X1    g11718(.A1(new_n11910_), .A2(new_n11905_), .ZN(new_n11911_));
  AOI22_X1   g11719(.A1(new_n11906_), .A2(\asqrt[59] ), .B1(new_n11904_), .B2(new_n11898_), .ZN(new_n11912_));
  NOR4_X1    g11720(.A1(new_n11631_), .A2(\asqrt[60] ), .A3(new_n11419_), .A4(new_n11560_), .ZN(new_n11913_));
  XOR2_X1    g11721(.A1(new_n11913_), .A2(new_n11549_), .Z(new_n11914_));
  NAND2_X1   g11722(.A1(new_n11914_), .A2(new_n229_), .ZN(new_n11915_));
  INV_X1     g11723(.I(new_n11915_), .ZN(new_n11916_));
  OAI21_X1   g11724(.A1(new_n11912_), .A2(new_n275_), .B(new_n11916_), .ZN(new_n11917_));
  NAND2_X1   g11725(.A1(new_n11917_), .A2(new_n11911_), .ZN(new_n11918_));
  OAI22_X1   g11726(.A1(new_n11912_), .A2(new_n275_), .B1(new_n11910_), .B2(new_n11905_), .ZN(new_n11919_));
  INV_X1     g11727(.I(new_n11602_), .ZN(new_n11920_));
  NOR2_X1    g11728(.A1(new_n11920_), .A2(\asqrt[62] ), .ZN(new_n11921_));
  INV_X1     g11729(.I(new_n11921_), .ZN(new_n11922_));
  NAND3_X1   g11730(.A1(new_n11919_), .A2(\asqrt[61] ), .A3(new_n11922_), .ZN(new_n11923_));
  OAI21_X1   g11731(.A1(new_n11923_), .A2(new_n11918_), .B(new_n11604_), .ZN(new_n11924_));
  NAND3_X1   g11732(.A1(new_n11631_), .A2(new_n11067_), .A3(new_n11634_), .ZN(new_n11925_));
  AOI21_X1   g11733(.A1(new_n11925_), .A2(new_n11582_), .B(\asqrt[63] ), .ZN(new_n11926_));
  INV_X1     g11734(.I(new_n11926_), .ZN(new_n11927_));
  OAI21_X1   g11735(.A1(new_n11924_), .A2(new_n11927_), .B(new_n11599_), .ZN(new_n11928_));
  INV_X1     g11736(.I(new_n11613_), .ZN(new_n11929_));
  AOI21_X1   g11737(.A1(new_n11622_), .A2(new_n11929_), .B(new_n11615_), .ZN(new_n11930_));
  NOR3_X1    g11738(.A1(new_n11612_), .A2(new_n11605_), .A3(new_n11610_), .ZN(new_n11931_));
  NOR2_X1    g11739(.A1(new_n11931_), .A2(new_n11930_), .ZN(new_n11932_));
  NOR3_X1    g11740(.A1(new_n11640_), .A2(new_n11080_), .A3(\asqrt[21] ), .ZN(new_n11933_));
  AOI21_X1   g11741(.A1(new_n11637_), .A2(new_n11079_), .B(new_n11631_), .ZN(new_n11934_));
  NOR4_X1    g11742(.A1(new_n11934_), .A2(new_n11933_), .A3(\asqrt[23] ), .A4(new_n11629_), .ZN(new_n11935_));
  NOR2_X1    g11743(.A1(new_n11935_), .A2(new_n11932_), .ZN(new_n11936_));
  NOR3_X1    g11744(.A1(new_n11931_), .A2(new_n11930_), .A3(new_n11629_), .ZN(new_n11937_));
  NOR3_X1    g11745(.A1(new_n11631_), .A2(new_n11103_), .A3(new_n11648_), .ZN(new_n11938_));
  AOI21_X1   g11746(.A1(\asqrt[21] ), .A2(new_n11649_), .B(new_n11104_), .ZN(new_n11939_));
  NOR3_X1    g11747(.A1(new_n11939_), .A2(new_n11938_), .A3(\asqrt[24] ), .ZN(new_n11940_));
  OAI21_X1   g11748(.A1(new_n11937_), .A2(new_n10614_), .B(new_n11940_), .ZN(new_n11941_));
  NAND2_X1   g11749(.A1(new_n11936_), .A2(new_n11941_), .ZN(new_n11942_));
  OAI22_X1   g11750(.A1(new_n11935_), .A2(new_n11932_), .B1(new_n10614_), .B2(new_n11937_), .ZN(new_n11943_));
  INV_X1     g11751(.I(new_n11659_), .ZN(new_n11944_));
  AOI21_X1   g11752(.A1(new_n11943_), .A2(\asqrt[24] ), .B(new_n11944_), .ZN(new_n11945_));
  NOR2_X1    g11753(.A1(new_n11945_), .A2(new_n11942_), .ZN(new_n11946_));
  AOI22_X1   g11754(.A1(new_n11943_), .A2(\asqrt[24] ), .B1(new_n11936_), .B2(new_n11941_), .ZN(new_n11947_));
  INV_X1     g11755(.I(new_n11666_), .ZN(new_n11948_));
  OAI21_X1   g11756(.A1(new_n11947_), .A2(new_n9672_), .B(new_n11948_), .ZN(new_n11949_));
  NAND2_X1   g11757(.A1(new_n11949_), .A2(new_n11946_), .ZN(new_n11950_));
  OAI22_X1   g11758(.A1(new_n11947_), .A2(new_n9672_), .B1(new_n11945_), .B2(new_n11942_), .ZN(new_n11951_));
  AOI21_X1   g11759(.A1(new_n11951_), .A2(\asqrt[26] ), .B(new_n11672_), .ZN(new_n11952_));
  NOR2_X1    g11760(.A1(new_n11952_), .A2(new_n11950_), .ZN(new_n11953_));
  AOI22_X1   g11761(.A1(new_n11951_), .A2(\asqrt[26] ), .B1(new_n11949_), .B2(new_n11946_), .ZN(new_n11954_));
  INV_X1     g11762(.I(new_n11679_), .ZN(new_n11955_));
  OAI21_X1   g11763(.A1(new_n11954_), .A2(new_n8763_), .B(new_n11955_), .ZN(new_n11956_));
  NAND2_X1   g11764(.A1(new_n11956_), .A2(new_n11953_), .ZN(new_n11957_));
  OAI22_X1   g11765(.A1(new_n11954_), .A2(new_n8763_), .B1(new_n11952_), .B2(new_n11950_), .ZN(new_n11958_));
  AOI21_X1   g11766(.A1(new_n11958_), .A2(\asqrt[28] ), .B(new_n11685_), .ZN(new_n11959_));
  NOR2_X1    g11767(.A1(new_n11959_), .A2(new_n11957_), .ZN(new_n11960_));
  AOI22_X1   g11768(.A1(new_n11958_), .A2(\asqrt[28] ), .B1(new_n11956_), .B2(new_n11953_), .ZN(new_n11961_));
  INV_X1     g11769(.I(new_n11692_), .ZN(new_n11962_));
  OAI21_X1   g11770(.A1(new_n11961_), .A2(new_n7931_), .B(new_n11962_), .ZN(new_n11963_));
  NAND2_X1   g11771(.A1(new_n11963_), .A2(new_n11960_), .ZN(new_n11964_));
  OAI22_X1   g11772(.A1(new_n11961_), .A2(new_n7931_), .B1(new_n11959_), .B2(new_n11957_), .ZN(new_n11965_));
  AOI21_X1   g11773(.A1(new_n11965_), .A2(\asqrt[30] ), .B(new_n11698_), .ZN(new_n11966_));
  NOR2_X1    g11774(.A1(new_n11966_), .A2(new_n11964_), .ZN(new_n11967_));
  AOI22_X1   g11775(.A1(new_n11965_), .A2(\asqrt[30] ), .B1(new_n11963_), .B2(new_n11960_), .ZN(new_n11968_));
  INV_X1     g11776(.I(new_n11706_), .ZN(new_n11969_));
  OAI21_X1   g11777(.A1(new_n11968_), .A2(new_n7110_), .B(new_n11969_), .ZN(new_n11970_));
  NAND2_X1   g11778(.A1(new_n11970_), .A2(new_n11967_), .ZN(new_n11971_));
  OAI22_X1   g11779(.A1(new_n11968_), .A2(new_n7110_), .B1(new_n11966_), .B2(new_n11964_), .ZN(new_n11972_));
  AOI21_X1   g11780(.A1(new_n11972_), .A2(\asqrt[32] ), .B(new_n11713_), .ZN(new_n11973_));
  NOR2_X1    g11781(.A1(new_n11973_), .A2(new_n11971_), .ZN(new_n11974_));
  AOI22_X1   g11782(.A1(new_n11972_), .A2(\asqrt[32] ), .B1(new_n11970_), .B2(new_n11967_), .ZN(new_n11975_));
  INV_X1     g11783(.I(new_n11721_), .ZN(new_n11976_));
  OAI21_X1   g11784(.A1(new_n11975_), .A2(new_n6365_), .B(new_n11976_), .ZN(new_n11977_));
  NAND2_X1   g11785(.A1(new_n11977_), .A2(new_n11974_), .ZN(new_n11978_));
  OAI22_X1   g11786(.A1(new_n11975_), .A2(new_n6365_), .B1(new_n11973_), .B2(new_n11971_), .ZN(new_n11979_));
  AOI21_X1   g11787(.A1(new_n11979_), .A2(\asqrt[34] ), .B(new_n11728_), .ZN(new_n11980_));
  NOR2_X1    g11788(.A1(new_n11980_), .A2(new_n11978_), .ZN(new_n11981_));
  AOI22_X1   g11789(.A1(new_n11979_), .A2(\asqrt[34] ), .B1(new_n11977_), .B2(new_n11974_), .ZN(new_n11982_));
  INV_X1     g11790(.I(new_n11736_), .ZN(new_n11983_));
  OAI21_X1   g11791(.A1(new_n11982_), .A2(new_n5626_), .B(new_n11983_), .ZN(new_n11984_));
  NAND2_X1   g11792(.A1(new_n11984_), .A2(new_n11981_), .ZN(new_n11985_));
  OAI22_X1   g11793(.A1(new_n11982_), .A2(new_n5626_), .B1(new_n11980_), .B2(new_n11978_), .ZN(new_n11986_));
  AOI21_X1   g11794(.A1(new_n11986_), .A2(\asqrt[36] ), .B(new_n11743_), .ZN(new_n11987_));
  NOR2_X1    g11795(.A1(new_n11987_), .A2(new_n11985_), .ZN(new_n11988_));
  AOI22_X1   g11796(.A1(new_n11986_), .A2(\asqrt[36] ), .B1(new_n11984_), .B2(new_n11981_), .ZN(new_n11989_));
  INV_X1     g11797(.I(new_n11751_), .ZN(new_n11990_));
  OAI21_X1   g11798(.A1(new_n11989_), .A2(new_n4973_), .B(new_n11990_), .ZN(new_n11991_));
  NAND2_X1   g11799(.A1(new_n11991_), .A2(new_n11988_), .ZN(new_n11992_));
  OAI22_X1   g11800(.A1(new_n11989_), .A2(new_n4973_), .B1(new_n11987_), .B2(new_n11985_), .ZN(new_n11993_));
  AOI21_X1   g11801(.A1(new_n11993_), .A2(\asqrt[38] ), .B(new_n11758_), .ZN(new_n11994_));
  NOR2_X1    g11802(.A1(new_n11994_), .A2(new_n11992_), .ZN(new_n11995_));
  AOI22_X1   g11803(.A1(new_n11993_), .A2(\asqrt[38] ), .B1(new_n11991_), .B2(new_n11988_), .ZN(new_n11996_));
  INV_X1     g11804(.I(new_n11766_), .ZN(new_n11997_));
  OAI21_X1   g11805(.A1(new_n11996_), .A2(new_n4330_), .B(new_n11997_), .ZN(new_n11998_));
  NAND2_X1   g11806(.A1(new_n11998_), .A2(new_n11995_), .ZN(new_n11999_));
  OAI22_X1   g11807(.A1(new_n11996_), .A2(new_n4330_), .B1(new_n11994_), .B2(new_n11992_), .ZN(new_n12000_));
  AOI21_X1   g11808(.A1(new_n12000_), .A2(\asqrt[40] ), .B(new_n11773_), .ZN(new_n12001_));
  NOR2_X1    g11809(.A1(new_n12001_), .A2(new_n11999_), .ZN(new_n12002_));
  AOI22_X1   g11810(.A1(new_n12000_), .A2(\asqrt[40] ), .B1(new_n11998_), .B2(new_n11995_), .ZN(new_n12003_));
  INV_X1     g11811(.I(new_n11781_), .ZN(new_n12004_));
  OAI21_X1   g11812(.A1(new_n12003_), .A2(new_n3760_), .B(new_n12004_), .ZN(new_n12005_));
  NAND2_X1   g11813(.A1(new_n12005_), .A2(new_n12002_), .ZN(new_n12006_));
  OAI22_X1   g11814(.A1(new_n12003_), .A2(new_n3760_), .B1(new_n12001_), .B2(new_n11999_), .ZN(new_n12007_));
  AOI21_X1   g11815(.A1(new_n12007_), .A2(\asqrt[42] ), .B(new_n11788_), .ZN(new_n12008_));
  NOR2_X1    g11816(.A1(new_n12008_), .A2(new_n12006_), .ZN(new_n12009_));
  AOI22_X1   g11817(.A1(new_n12007_), .A2(\asqrt[42] ), .B1(new_n12005_), .B2(new_n12002_), .ZN(new_n12010_));
  INV_X1     g11818(.I(new_n11796_), .ZN(new_n12011_));
  OAI21_X1   g11819(.A1(new_n12010_), .A2(new_n3208_), .B(new_n12011_), .ZN(new_n12012_));
  NAND2_X1   g11820(.A1(new_n12012_), .A2(new_n12009_), .ZN(new_n12013_));
  OAI22_X1   g11821(.A1(new_n12010_), .A2(new_n3208_), .B1(new_n12008_), .B2(new_n12006_), .ZN(new_n12014_));
  AOI21_X1   g11822(.A1(new_n12014_), .A2(\asqrt[44] ), .B(new_n11803_), .ZN(new_n12015_));
  NOR2_X1    g11823(.A1(new_n12015_), .A2(new_n12013_), .ZN(new_n12016_));
  AOI22_X1   g11824(.A1(new_n12014_), .A2(\asqrt[44] ), .B1(new_n12012_), .B2(new_n12009_), .ZN(new_n12017_));
  INV_X1     g11825(.I(new_n11811_), .ZN(new_n12018_));
  OAI21_X1   g11826(.A1(new_n12017_), .A2(new_n2728_), .B(new_n12018_), .ZN(new_n12019_));
  NAND2_X1   g11827(.A1(new_n12019_), .A2(new_n12016_), .ZN(new_n12020_));
  OAI22_X1   g11828(.A1(new_n12017_), .A2(new_n2728_), .B1(new_n12015_), .B2(new_n12013_), .ZN(new_n12021_));
  AOI21_X1   g11829(.A1(new_n12021_), .A2(\asqrt[46] ), .B(new_n11818_), .ZN(new_n12022_));
  NOR2_X1    g11830(.A1(new_n12022_), .A2(new_n12020_), .ZN(new_n12023_));
  AOI22_X1   g11831(.A1(new_n12021_), .A2(\asqrt[46] ), .B1(new_n12019_), .B2(new_n12016_), .ZN(new_n12024_));
  INV_X1     g11832(.I(new_n11826_), .ZN(new_n12025_));
  OAI21_X1   g11833(.A1(new_n12024_), .A2(new_n2253_), .B(new_n12025_), .ZN(new_n12026_));
  NAND2_X1   g11834(.A1(new_n12026_), .A2(new_n12023_), .ZN(new_n12027_));
  OAI22_X1   g11835(.A1(new_n12024_), .A2(new_n2253_), .B1(new_n12022_), .B2(new_n12020_), .ZN(new_n12028_));
  AOI21_X1   g11836(.A1(new_n12028_), .A2(\asqrt[48] ), .B(new_n11833_), .ZN(new_n12029_));
  NOR2_X1    g11837(.A1(new_n12029_), .A2(new_n12027_), .ZN(new_n12030_));
  AOI22_X1   g11838(.A1(new_n12028_), .A2(\asqrt[48] ), .B1(new_n12026_), .B2(new_n12023_), .ZN(new_n12031_));
  INV_X1     g11839(.I(new_n11841_), .ZN(new_n12032_));
  OAI21_X1   g11840(.A1(new_n12031_), .A2(new_n1854_), .B(new_n12032_), .ZN(new_n12033_));
  NAND2_X1   g11841(.A1(new_n12033_), .A2(new_n12030_), .ZN(new_n12034_));
  OAI22_X1   g11842(.A1(new_n12031_), .A2(new_n1854_), .B1(new_n12029_), .B2(new_n12027_), .ZN(new_n12035_));
  AOI21_X1   g11843(.A1(new_n12035_), .A2(\asqrt[50] ), .B(new_n11848_), .ZN(new_n12036_));
  NOR2_X1    g11844(.A1(new_n12036_), .A2(new_n12034_), .ZN(new_n12037_));
  AOI22_X1   g11845(.A1(new_n12035_), .A2(\asqrt[50] ), .B1(new_n12033_), .B2(new_n12030_), .ZN(new_n12038_));
  INV_X1     g11846(.I(new_n11856_), .ZN(new_n12039_));
  OAI21_X1   g11847(.A1(new_n12038_), .A2(new_n1436_), .B(new_n12039_), .ZN(new_n12040_));
  NAND2_X1   g11848(.A1(new_n12040_), .A2(new_n12037_), .ZN(new_n12041_));
  OAI22_X1   g11849(.A1(new_n12038_), .A2(new_n1436_), .B1(new_n12036_), .B2(new_n12034_), .ZN(new_n12042_));
  AOI21_X1   g11850(.A1(new_n12042_), .A2(\asqrt[52] ), .B(new_n11863_), .ZN(new_n12043_));
  NOR2_X1    g11851(.A1(new_n12043_), .A2(new_n12041_), .ZN(new_n12044_));
  AOI22_X1   g11852(.A1(new_n12042_), .A2(\asqrt[52] ), .B1(new_n12040_), .B2(new_n12037_), .ZN(new_n12045_));
  INV_X1     g11853(.I(new_n11870_), .ZN(new_n12046_));
  OAI21_X1   g11854(.A1(new_n12045_), .A2(new_n1096_), .B(new_n12046_), .ZN(new_n12047_));
  NAND2_X1   g11855(.A1(new_n12047_), .A2(new_n12044_), .ZN(new_n12048_));
  OAI22_X1   g11856(.A1(new_n12045_), .A2(new_n1096_), .B1(new_n12043_), .B2(new_n12041_), .ZN(new_n12049_));
  AOI21_X1   g11857(.A1(new_n12049_), .A2(\asqrt[54] ), .B(new_n11876_), .ZN(new_n12050_));
  NOR2_X1    g11858(.A1(new_n12050_), .A2(new_n12048_), .ZN(new_n12051_));
  AOI22_X1   g11859(.A1(new_n12049_), .A2(\asqrt[54] ), .B1(new_n12047_), .B2(new_n12044_), .ZN(new_n12052_));
  INV_X1     g11860(.I(new_n11883_), .ZN(new_n12053_));
  OAI21_X1   g11861(.A1(new_n12052_), .A2(new_n825_), .B(new_n12053_), .ZN(new_n12054_));
  NAND2_X1   g11862(.A1(new_n12054_), .A2(new_n12051_), .ZN(new_n12055_));
  OAI22_X1   g11863(.A1(new_n12052_), .A2(new_n825_), .B1(new_n12050_), .B2(new_n12048_), .ZN(new_n12056_));
  AOI21_X1   g11864(.A1(new_n12056_), .A2(\asqrt[56] ), .B(new_n11889_), .ZN(new_n12057_));
  NOR2_X1    g11865(.A1(new_n12057_), .A2(new_n12055_), .ZN(new_n12058_));
  AOI22_X1   g11866(.A1(new_n12056_), .A2(\asqrt[56] ), .B1(new_n12054_), .B2(new_n12051_), .ZN(new_n12059_));
  INV_X1     g11867(.I(new_n11896_), .ZN(new_n12060_));
  OAI21_X1   g11868(.A1(new_n12059_), .A2(new_n587_), .B(new_n12060_), .ZN(new_n12061_));
  NAND2_X1   g11869(.A1(new_n12061_), .A2(new_n12058_), .ZN(new_n12062_));
  OAI22_X1   g11870(.A1(new_n12059_), .A2(new_n587_), .B1(new_n12057_), .B2(new_n12055_), .ZN(new_n12063_));
  AOI21_X1   g11871(.A1(new_n12063_), .A2(\asqrt[58] ), .B(new_n11902_), .ZN(new_n12064_));
  NOR2_X1    g11872(.A1(new_n12064_), .A2(new_n12062_), .ZN(new_n12065_));
  AOI22_X1   g11873(.A1(new_n12063_), .A2(\asqrt[58] ), .B1(new_n12061_), .B2(new_n12058_), .ZN(new_n12066_));
  INV_X1     g11874(.I(new_n11909_), .ZN(new_n12067_));
  OAI21_X1   g11875(.A1(new_n12066_), .A2(new_n376_), .B(new_n12067_), .ZN(new_n12068_));
  NAND2_X1   g11876(.A1(new_n12068_), .A2(new_n12065_), .ZN(new_n12069_));
  OAI22_X1   g11877(.A1(new_n12066_), .A2(new_n376_), .B1(new_n12064_), .B2(new_n12062_), .ZN(new_n12070_));
  AOI21_X1   g11878(.A1(new_n12070_), .A2(\asqrt[60] ), .B(new_n11915_), .ZN(new_n12071_));
  AOI22_X1   g11879(.A1(new_n12070_), .A2(\asqrt[60] ), .B1(new_n12068_), .B2(new_n12065_), .ZN(new_n12072_));
  OAI22_X1   g11880(.A1(new_n12072_), .A2(new_n229_), .B1(new_n12071_), .B2(new_n12069_), .ZN(new_n12073_));
  NOR4_X1    g11881(.A1(new_n12073_), .A2(\asqrt[62] ), .A3(new_n11598_), .A4(new_n11602_), .ZN(new_n12074_));
  NAND2_X1   g11882(.A1(new_n11618_), .A2(new_n11067_), .ZN(new_n12075_));
  XOR2_X1    g11883(.A1(new_n11618_), .A2(\asqrt[63] ), .Z(new_n12076_));
  AOI21_X1   g11884(.A1(\asqrt[21] ), .A2(new_n12075_), .B(new_n12076_), .ZN(new_n12077_));
  NAND2_X1   g11885(.A1(new_n12074_), .A2(new_n12077_), .ZN(new_n12078_));
  NOR4_X1    g11886(.A1(new_n12078_), .A2(new_n11579_), .A3(new_n11928_), .A4(new_n11586_), .ZN(new_n12079_));
  NOR2_X1    g11887(.A1(new_n11579_), .A2(\a[40] ), .ZN(new_n12080_));
  OAI21_X1   g11888(.A1(new_n12079_), .A2(new_n12080_), .B(new_n11578_), .ZN(new_n12081_));
  INV_X1     g11889(.I(new_n11578_), .ZN(new_n12082_));
  INV_X1     g11890(.I(new_n11586_), .ZN(new_n12083_));
  NOR2_X1    g11891(.A1(new_n12071_), .A2(new_n12069_), .ZN(new_n12084_));
  NOR3_X1    g11892(.A1(new_n12072_), .A2(new_n229_), .A3(new_n11921_), .ZN(new_n12085_));
  AOI21_X1   g11893(.A1(new_n12085_), .A2(new_n12084_), .B(new_n11603_), .ZN(new_n12086_));
  AOI21_X1   g11894(.A1(new_n12086_), .A2(new_n11926_), .B(new_n11598_), .ZN(new_n12087_));
  AOI22_X1   g11895(.A1(new_n11919_), .A2(\asqrt[61] ), .B1(new_n11917_), .B2(new_n11911_), .ZN(new_n12088_));
  NAND4_X1   g11896(.A1(new_n12088_), .A2(new_n196_), .A3(new_n11599_), .A4(new_n11920_), .ZN(new_n12089_));
  INV_X1     g11897(.I(new_n12077_), .ZN(new_n12090_));
  NOR2_X1    g11898(.A1(new_n12089_), .A2(new_n12090_), .ZN(new_n12091_));
  NAND4_X1   g11899(.A1(new_n12091_), .A2(new_n12087_), .A3(\a[41] ), .A4(new_n12083_), .ZN(new_n12092_));
  NAND3_X1   g11900(.A1(new_n12092_), .A2(\a[40] ), .A3(new_n12082_), .ZN(new_n12093_));
  NAND2_X1   g11901(.A1(new_n12081_), .A2(new_n12093_), .ZN(new_n12094_));
  NOR2_X1    g11902(.A1(new_n12078_), .A2(new_n11928_), .ZN(new_n12095_));
  NOR4_X1    g11903(.A1(new_n11584_), .A2(new_n11067_), .A3(new_n11633_), .A4(new_n11571_), .ZN(new_n12096_));
  NAND2_X1   g11904(.A1(\asqrt[21] ), .A2(\a[40] ), .ZN(new_n12097_));
  XOR2_X1    g11905(.A1(new_n12097_), .A2(new_n12096_), .Z(new_n12098_));
  NOR2_X1    g11906(.A1(new_n12098_), .A2(new_n11575_), .ZN(new_n12099_));
  INV_X1     g11907(.I(new_n12099_), .ZN(new_n12100_));
  NAND3_X1   g11908(.A1(new_n12091_), .A2(new_n12087_), .A3(new_n12083_), .ZN(new_n12101_));
  NAND2_X1   g11909(.A1(new_n11880_), .A2(\asqrt[55] ), .ZN(new_n12102_));
  AOI21_X1   g11910(.A1(new_n12102_), .A2(new_n11879_), .B(new_n724_), .ZN(new_n12103_));
  OAI21_X1   g11911(.A1(new_n11885_), .A2(new_n12103_), .B(\asqrt[57] ), .ZN(new_n12104_));
  AOI21_X1   g11912(.A1(new_n11892_), .A2(new_n12104_), .B(new_n504_), .ZN(new_n12105_));
  OAI21_X1   g11913(.A1(new_n11898_), .A2(new_n12105_), .B(\asqrt[59] ), .ZN(new_n12106_));
  AOI21_X1   g11914(.A1(new_n11905_), .A2(new_n12106_), .B(new_n275_), .ZN(new_n12107_));
  OAI21_X1   g11915(.A1(new_n11911_), .A2(new_n12107_), .B(\asqrt[61] ), .ZN(new_n12108_));
  NOR3_X1    g11916(.A1(new_n11918_), .A2(new_n12108_), .A3(new_n11921_), .ZN(new_n12109_));
  NOR3_X1    g11917(.A1(new_n12109_), .A2(new_n11603_), .A3(new_n11927_), .ZN(new_n12110_));
  OAI21_X1   g11918(.A1(new_n12110_), .A2(new_n11598_), .B(new_n12089_), .ZN(new_n12111_));
  NOR2_X1    g11919(.A1(new_n12083_), .A2(new_n12077_), .ZN(new_n12112_));
  NAND2_X1   g11920(.A1(new_n12112_), .A2(\asqrt[21] ), .ZN(new_n12113_));
  OAI21_X1   g11921(.A1(new_n12111_), .A2(new_n12113_), .B(new_n11605_), .ZN(new_n12114_));
  NAND3_X1   g11922(.A1(new_n12114_), .A2(new_n11606_), .A3(new_n12101_), .ZN(new_n12115_));
  NOR4_X1    g11923(.A1(new_n11928_), .A2(new_n11586_), .A3(new_n12089_), .A4(new_n12090_), .ZN(\asqrt[20] ));
  NAND2_X1   g11924(.A1(new_n12049_), .A2(\asqrt[54] ), .ZN(new_n12117_));
  AOI21_X1   g11925(.A1(new_n12117_), .A2(new_n12048_), .B(new_n825_), .ZN(new_n12118_));
  OAI21_X1   g11926(.A1(new_n12051_), .A2(new_n12118_), .B(\asqrt[56] ), .ZN(new_n12119_));
  AOI21_X1   g11927(.A1(new_n12055_), .A2(new_n12119_), .B(new_n587_), .ZN(new_n12120_));
  OAI21_X1   g11928(.A1(new_n12058_), .A2(new_n12120_), .B(\asqrt[58] ), .ZN(new_n12121_));
  AOI21_X1   g11929(.A1(new_n12062_), .A2(new_n12121_), .B(new_n376_), .ZN(new_n12122_));
  OAI21_X1   g11930(.A1(new_n12065_), .A2(new_n12122_), .B(\asqrt[60] ), .ZN(new_n12123_));
  AOI21_X1   g11931(.A1(new_n12069_), .A2(new_n12123_), .B(new_n229_), .ZN(new_n12124_));
  NAND4_X1   g11932(.A1(new_n12124_), .A2(new_n11911_), .A3(new_n11917_), .A4(new_n11922_), .ZN(new_n12125_));
  NAND3_X1   g11933(.A1(new_n12125_), .A2(new_n11604_), .A3(new_n11926_), .ZN(new_n12126_));
  AOI21_X1   g11934(.A1(new_n11599_), .A2(new_n12126_), .B(new_n12074_), .ZN(new_n12127_));
  INV_X1     g11935(.I(new_n12113_), .ZN(new_n12128_));
  AOI21_X1   g11936(.A1(new_n12127_), .A2(new_n12128_), .B(\a[42] ), .ZN(new_n12129_));
  OAI21_X1   g11937(.A1(new_n12129_), .A2(new_n11607_), .B(\asqrt[20] ), .ZN(new_n12130_));
  NAND4_X1   g11938(.A1(new_n12130_), .A2(new_n12115_), .A3(new_n11105_), .A4(new_n12100_), .ZN(new_n12131_));
  NAND2_X1   g11939(.A1(new_n12131_), .A2(new_n12094_), .ZN(new_n12132_));
  NAND3_X1   g11940(.A1(new_n12081_), .A2(new_n12093_), .A3(new_n12100_), .ZN(new_n12133_));
  AOI21_X1   g11941(.A1(\asqrt[21] ), .A2(new_n11605_), .B(\a[43] ), .ZN(new_n12134_));
  NOR2_X1    g11942(.A1(new_n11622_), .A2(\a[42] ), .ZN(new_n12135_));
  AOI21_X1   g11943(.A1(\asqrt[21] ), .A2(\a[42] ), .B(new_n11609_), .ZN(new_n12136_));
  OAI21_X1   g11944(.A1(new_n12135_), .A2(new_n12134_), .B(new_n12136_), .ZN(new_n12137_));
  INV_X1     g11945(.I(new_n12137_), .ZN(new_n12138_));
  NAND3_X1   g11946(.A1(\asqrt[20] ), .A2(new_n11630_), .A3(new_n12138_), .ZN(new_n12139_));
  OAI21_X1   g11947(.A1(new_n12101_), .A2(new_n12137_), .B(new_n11629_), .ZN(new_n12140_));
  NAND3_X1   g11948(.A1(new_n12140_), .A2(new_n12139_), .A3(new_n10614_), .ZN(new_n12141_));
  AOI21_X1   g11949(.A1(new_n12133_), .A2(\asqrt[22] ), .B(new_n12141_), .ZN(new_n12142_));
  NOR2_X1    g11950(.A1(new_n12132_), .A2(new_n12142_), .ZN(new_n12143_));
  NAND2_X1   g11951(.A1(new_n12133_), .A2(\asqrt[22] ), .ZN(new_n12144_));
  AOI21_X1   g11952(.A1(new_n12132_), .A2(new_n12144_), .B(new_n10614_), .ZN(new_n12145_));
  NAND2_X1   g11953(.A1(new_n11644_), .A2(\asqrt[23] ), .ZN(new_n12146_));
  INV_X1     g11954(.I(new_n12146_), .ZN(new_n12147_));
  NAND2_X1   g11955(.A1(new_n11638_), .A2(new_n11641_), .ZN(new_n12148_));
  NAND3_X1   g11956(.A1(new_n12148_), .A2(new_n11937_), .A3(new_n10614_), .ZN(new_n12149_));
  NOR3_X1    g11957(.A1(new_n12101_), .A2(new_n12147_), .A3(new_n12149_), .ZN(new_n12150_));
  NOR2_X1    g11958(.A1(new_n12101_), .A2(new_n12149_), .ZN(new_n12151_));
  NOR2_X1    g11959(.A1(new_n12151_), .A2(new_n12146_), .ZN(new_n12152_));
  NOR3_X1    g11960(.A1(new_n12152_), .A2(\asqrt[24] ), .A3(new_n12150_), .ZN(new_n12153_));
  INV_X1     g11961(.I(new_n12153_), .ZN(new_n12154_));
  OAI21_X1   g11962(.A1(new_n12145_), .A2(new_n12154_), .B(new_n12143_), .ZN(new_n12155_));
  OAI21_X1   g11963(.A1(new_n12145_), .A2(new_n12143_), .B(\asqrt[24] ), .ZN(new_n12156_));
  NAND2_X1   g11964(.A1(new_n11943_), .A2(\asqrt[24] ), .ZN(new_n12157_));
  NOR2_X1    g11965(.A1(new_n11939_), .A2(new_n11938_), .ZN(new_n12158_));
  NOR4_X1    g11966(.A1(new_n12101_), .A2(\asqrt[24] ), .A3(new_n12158_), .A4(new_n11943_), .ZN(new_n12159_));
  XOR2_X1    g11967(.A1(new_n12159_), .A2(new_n12157_), .Z(new_n12160_));
  NAND2_X1   g11968(.A1(new_n12160_), .A2(new_n9672_), .ZN(new_n12161_));
  INV_X1     g11969(.I(new_n12161_), .ZN(new_n12162_));
  AOI21_X1   g11970(.A1(new_n12156_), .A2(new_n12162_), .B(new_n12155_), .ZN(new_n12163_));
  AOI21_X1   g11971(.A1(new_n12155_), .A2(new_n12156_), .B(new_n9672_), .ZN(new_n12164_));
  NAND2_X1   g11972(.A1(new_n11662_), .A2(\asqrt[25] ), .ZN(new_n12165_));
  NOR2_X1    g11973(.A1(new_n11657_), .A2(new_n11658_), .ZN(new_n12166_));
  NOR4_X1    g11974(.A1(new_n12101_), .A2(\asqrt[25] ), .A3(new_n12166_), .A4(new_n11662_), .ZN(new_n12167_));
  XOR2_X1    g11975(.A1(new_n12167_), .A2(new_n12165_), .Z(new_n12168_));
  NAND2_X1   g11976(.A1(new_n12168_), .A2(new_n9212_), .ZN(new_n12169_));
  OAI21_X1   g11977(.A1(new_n12164_), .A2(new_n12169_), .B(new_n12163_), .ZN(new_n12170_));
  OAI21_X1   g11978(.A1(new_n12163_), .A2(new_n12164_), .B(\asqrt[26] ), .ZN(new_n12171_));
  NOR4_X1    g11979(.A1(new_n12101_), .A2(\asqrt[26] ), .A3(new_n11665_), .A4(new_n11951_), .ZN(new_n12172_));
  AOI21_X1   g11980(.A1(new_n12165_), .A2(new_n11661_), .B(new_n9212_), .ZN(new_n12173_));
  NOR2_X1    g11981(.A1(new_n12172_), .A2(new_n12173_), .ZN(new_n12174_));
  NAND2_X1   g11982(.A1(new_n12174_), .A2(new_n8763_), .ZN(new_n12175_));
  INV_X1     g11983(.I(new_n12175_), .ZN(new_n12176_));
  AOI21_X1   g11984(.A1(new_n12171_), .A2(new_n12176_), .B(new_n12170_), .ZN(new_n12177_));
  AOI22_X1   g11985(.A1(new_n12131_), .A2(new_n12094_), .B1(\asqrt[22] ), .B2(new_n12133_), .ZN(new_n12178_));
  OAI21_X1   g11986(.A1(new_n12178_), .A2(new_n10614_), .B(new_n12153_), .ZN(new_n12179_));
  OAI22_X1   g11987(.A1(new_n12178_), .A2(new_n10614_), .B1(new_n12132_), .B2(new_n12142_), .ZN(new_n12180_));
  AOI22_X1   g11988(.A1(new_n12180_), .A2(\asqrt[24] ), .B1(new_n12179_), .B2(new_n12143_), .ZN(new_n12181_));
  INV_X1     g11989(.I(new_n12169_), .ZN(new_n12182_));
  OAI21_X1   g11990(.A1(new_n12181_), .A2(new_n9672_), .B(new_n12182_), .ZN(new_n12183_));
  AOI21_X1   g11991(.A1(new_n12180_), .A2(\asqrt[24] ), .B(new_n12161_), .ZN(new_n12184_));
  OAI22_X1   g11992(.A1(new_n12181_), .A2(new_n9672_), .B1(new_n12184_), .B2(new_n12155_), .ZN(new_n12185_));
  AOI22_X1   g11993(.A1(new_n12185_), .A2(\asqrt[26] ), .B1(new_n12183_), .B2(new_n12163_), .ZN(new_n12186_));
  NAND2_X1   g11994(.A1(new_n11676_), .A2(\asqrt[27] ), .ZN(new_n12187_));
  NOR4_X1    g11995(.A1(new_n12101_), .A2(\asqrt[27] ), .A3(new_n11671_), .A4(new_n11676_), .ZN(new_n12188_));
  XOR2_X1    g11996(.A1(new_n12188_), .A2(new_n12187_), .Z(new_n12189_));
  NAND2_X1   g11997(.A1(new_n12189_), .A2(new_n8319_), .ZN(new_n12190_));
  INV_X1     g11998(.I(new_n12190_), .ZN(new_n12191_));
  OAI21_X1   g11999(.A1(new_n12186_), .A2(new_n8763_), .B(new_n12191_), .ZN(new_n12192_));
  NAND2_X1   g12000(.A1(new_n12192_), .A2(new_n12177_), .ZN(new_n12193_));
  AOI21_X1   g12001(.A1(new_n12185_), .A2(\asqrt[26] ), .B(new_n12175_), .ZN(new_n12194_));
  OAI22_X1   g12002(.A1(new_n12186_), .A2(new_n8763_), .B1(new_n12194_), .B2(new_n12170_), .ZN(new_n12195_));
  NOR4_X1    g12003(.A1(new_n12101_), .A2(\asqrt[28] ), .A3(new_n11678_), .A4(new_n11958_), .ZN(new_n12196_));
  AOI21_X1   g12004(.A1(new_n12187_), .A2(new_n11675_), .B(new_n8319_), .ZN(new_n12197_));
  NOR2_X1    g12005(.A1(new_n12196_), .A2(new_n12197_), .ZN(new_n12198_));
  NAND2_X1   g12006(.A1(new_n12198_), .A2(new_n7931_), .ZN(new_n12199_));
  AOI21_X1   g12007(.A1(new_n12195_), .A2(\asqrt[28] ), .B(new_n12199_), .ZN(new_n12200_));
  NOR2_X1    g12008(.A1(new_n12200_), .A2(new_n12193_), .ZN(new_n12201_));
  AOI22_X1   g12009(.A1(new_n12195_), .A2(\asqrt[28] ), .B1(new_n12192_), .B2(new_n12177_), .ZN(new_n12202_));
  NAND2_X1   g12010(.A1(new_n11689_), .A2(\asqrt[29] ), .ZN(new_n12203_));
  NOR4_X1    g12011(.A1(new_n12101_), .A2(\asqrt[29] ), .A3(new_n11684_), .A4(new_n11689_), .ZN(new_n12204_));
  XOR2_X1    g12012(.A1(new_n12204_), .A2(new_n12203_), .Z(new_n12205_));
  NAND2_X1   g12013(.A1(new_n12205_), .A2(new_n7517_), .ZN(new_n12206_));
  INV_X1     g12014(.I(new_n12206_), .ZN(new_n12207_));
  OAI21_X1   g12015(.A1(new_n12202_), .A2(new_n7931_), .B(new_n12207_), .ZN(new_n12208_));
  NAND2_X1   g12016(.A1(new_n12208_), .A2(new_n12201_), .ZN(new_n12209_));
  OAI22_X1   g12017(.A1(new_n12202_), .A2(new_n7931_), .B1(new_n12200_), .B2(new_n12193_), .ZN(new_n12210_));
  NOR4_X1    g12018(.A1(new_n12101_), .A2(\asqrt[30] ), .A3(new_n11691_), .A4(new_n11965_), .ZN(new_n12211_));
  AOI21_X1   g12019(.A1(new_n12203_), .A2(new_n11688_), .B(new_n7517_), .ZN(new_n12212_));
  NOR2_X1    g12020(.A1(new_n12211_), .A2(new_n12212_), .ZN(new_n12213_));
  NAND2_X1   g12021(.A1(new_n12213_), .A2(new_n7110_), .ZN(new_n12214_));
  AOI21_X1   g12022(.A1(new_n12210_), .A2(\asqrt[30] ), .B(new_n12214_), .ZN(new_n12215_));
  NOR2_X1    g12023(.A1(new_n12215_), .A2(new_n12209_), .ZN(new_n12216_));
  AOI22_X1   g12024(.A1(new_n12210_), .A2(\asqrt[30] ), .B1(new_n12208_), .B2(new_n12201_), .ZN(new_n12217_));
  NAND2_X1   g12025(.A1(new_n11702_), .A2(\asqrt[31] ), .ZN(new_n12218_));
  NOR4_X1    g12026(.A1(new_n12101_), .A2(\asqrt[31] ), .A3(new_n11697_), .A4(new_n11702_), .ZN(new_n12219_));
  XOR2_X1    g12027(.A1(new_n12219_), .A2(new_n12218_), .Z(new_n12220_));
  NAND2_X1   g12028(.A1(new_n12220_), .A2(new_n6708_), .ZN(new_n12221_));
  INV_X1     g12029(.I(new_n12221_), .ZN(new_n12222_));
  OAI21_X1   g12030(.A1(new_n12217_), .A2(new_n7110_), .B(new_n12222_), .ZN(new_n12223_));
  NAND2_X1   g12031(.A1(new_n12223_), .A2(new_n12216_), .ZN(new_n12224_));
  OAI22_X1   g12032(.A1(new_n12217_), .A2(new_n7110_), .B1(new_n12215_), .B2(new_n12209_), .ZN(new_n12225_));
  NAND2_X1   g12033(.A1(new_n11972_), .A2(\asqrt[32] ), .ZN(new_n12226_));
  NOR4_X1    g12034(.A1(new_n12101_), .A2(\asqrt[32] ), .A3(new_n11705_), .A4(new_n11972_), .ZN(new_n12227_));
  XOR2_X1    g12035(.A1(new_n12227_), .A2(new_n12226_), .Z(new_n12228_));
  NAND2_X1   g12036(.A1(new_n12228_), .A2(new_n6365_), .ZN(new_n12229_));
  AOI21_X1   g12037(.A1(new_n12225_), .A2(\asqrt[32] ), .B(new_n12229_), .ZN(new_n12230_));
  NOR2_X1    g12038(.A1(new_n12230_), .A2(new_n12224_), .ZN(new_n12231_));
  AOI22_X1   g12039(.A1(new_n12225_), .A2(\asqrt[32] ), .B1(new_n12223_), .B2(new_n12216_), .ZN(new_n12232_));
  NOR4_X1    g12040(.A1(new_n12101_), .A2(\asqrt[33] ), .A3(new_n11712_), .A4(new_n11717_), .ZN(new_n12233_));
  AOI21_X1   g12041(.A1(new_n12226_), .A2(new_n11971_), .B(new_n6365_), .ZN(new_n12234_));
  NOR2_X1    g12042(.A1(new_n12233_), .A2(new_n12234_), .ZN(new_n12235_));
  NAND2_X1   g12043(.A1(new_n12235_), .A2(new_n5991_), .ZN(new_n12236_));
  INV_X1     g12044(.I(new_n12236_), .ZN(new_n12237_));
  OAI21_X1   g12045(.A1(new_n12232_), .A2(new_n6365_), .B(new_n12237_), .ZN(new_n12238_));
  NAND2_X1   g12046(.A1(new_n12238_), .A2(new_n12231_), .ZN(new_n12239_));
  OAI22_X1   g12047(.A1(new_n12232_), .A2(new_n6365_), .B1(new_n12230_), .B2(new_n12224_), .ZN(new_n12240_));
  NAND2_X1   g12048(.A1(new_n11979_), .A2(\asqrt[34] ), .ZN(new_n12241_));
  NOR4_X1    g12049(.A1(new_n12101_), .A2(\asqrt[34] ), .A3(new_n11720_), .A4(new_n11979_), .ZN(new_n12242_));
  XOR2_X1    g12050(.A1(new_n12242_), .A2(new_n12241_), .Z(new_n12243_));
  NAND2_X1   g12051(.A1(new_n12243_), .A2(new_n5626_), .ZN(new_n12244_));
  AOI21_X1   g12052(.A1(new_n12240_), .A2(\asqrt[34] ), .B(new_n12244_), .ZN(new_n12245_));
  NOR2_X1    g12053(.A1(new_n12245_), .A2(new_n12239_), .ZN(new_n12246_));
  AOI22_X1   g12054(.A1(new_n12240_), .A2(\asqrt[34] ), .B1(new_n12238_), .B2(new_n12231_), .ZN(new_n12247_));
  NOR4_X1    g12055(.A1(new_n12101_), .A2(\asqrt[35] ), .A3(new_n11727_), .A4(new_n11732_), .ZN(new_n12248_));
  AOI21_X1   g12056(.A1(new_n12241_), .A2(new_n11978_), .B(new_n5626_), .ZN(new_n12249_));
  NOR2_X1    g12057(.A1(new_n12248_), .A2(new_n12249_), .ZN(new_n12250_));
  NAND2_X1   g12058(.A1(new_n12250_), .A2(new_n5273_), .ZN(new_n12251_));
  INV_X1     g12059(.I(new_n12251_), .ZN(new_n12252_));
  OAI21_X1   g12060(.A1(new_n12247_), .A2(new_n5626_), .B(new_n12252_), .ZN(new_n12253_));
  NAND2_X1   g12061(.A1(new_n12253_), .A2(new_n12246_), .ZN(new_n12254_));
  OAI22_X1   g12062(.A1(new_n12247_), .A2(new_n5626_), .B1(new_n12245_), .B2(new_n12239_), .ZN(new_n12255_));
  NAND2_X1   g12063(.A1(new_n11986_), .A2(\asqrt[36] ), .ZN(new_n12256_));
  NOR4_X1    g12064(.A1(new_n12101_), .A2(\asqrt[36] ), .A3(new_n11735_), .A4(new_n11986_), .ZN(new_n12257_));
  XOR2_X1    g12065(.A1(new_n12257_), .A2(new_n12256_), .Z(new_n12258_));
  NAND2_X1   g12066(.A1(new_n12258_), .A2(new_n4973_), .ZN(new_n12259_));
  AOI21_X1   g12067(.A1(new_n12255_), .A2(\asqrt[36] ), .B(new_n12259_), .ZN(new_n12260_));
  NOR2_X1    g12068(.A1(new_n12260_), .A2(new_n12254_), .ZN(new_n12261_));
  AOI22_X1   g12069(.A1(new_n12255_), .A2(\asqrt[36] ), .B1(new_n12253_), .B2(new_n12246_), .ZN(new_n12262_));
  NOR4_X1    g12070(.A1(new_n12101_), .A2(\asqrt[37] ), .A3(new_n11742_), .A4(new_n11747_), .ZN(new_n12263_));
  AOI21_X1   g12071(.A1(new_n12256_), .A2(new_n11985_), .B(new_n4973_), .ZN(new_n12264_));
  NOR2_X1    g12072(.A1(new_n12263_), .A2(new_n12264_), .ZN(new_n12265_));
  NAND2_X1   g12073(.A1(new_n12265_), .A2(new_n4645_), .ZN(new_n12266_));
  INV_X1     g12074(.I(new_n12266_), .ZN(new_n12267_));
  OAI21_X1   g12075(.A1(new_n12262_), .A2(new_n4973_), .B(new_n12267_), .ZN(new_n12268_));
  NAND2_X1   g12076(.A1(new_n12268_), .A2(new_n12261_), .ZN(new_n12269_));
  OAI22_X1   g12077(.A1(new_n12262_), .A2(new_n4973_), .B1(new_n12260_), .B2(new_n12254_), .ZN(new_n12270_));
  NAND2_X1   g12078(.A1(new_n11993_), .A2(\asqrt[38] ), .ZN(new_n12271_));
  NOR4_X1    g12079(.A1(new_n12101_), .A2(\asqrt[38] ), .A3(new_n11750_), .A4(new_n11993_), .ZN(new_n12272_));
  XOR2_X1    g12080(.A1(new_n12272_), .A2(new_n12271_), .Z(new_n12273_));
  NAND2_X1   g12081(.A1(new_n12273_), .A2(new_n4330_), .ZN(new_n12274_));
  AOI21_X1   g12082(.A1(new_n12270_), .A2(\asqrt[38] ), .B(new_n12274_), .ZN(new_n12275_));
  NOR2_X1    g12083(.A1(new_n12275_), .A2(new_n12269_), .ZN(new_n12276_));
  AOI22_X1   g12084(.A1(new_n12270_), .A2(\asqrt[38] ), .B1(new_n12268_), .B2(new_n12261_), .ZN(new_n12277_));
  NOR4_X1    g12085(.A1(new_n12101_), .A2(\asqrt[39] ), .A3(new_n11757_), .A4(new_n11762_), .ZN(new_n12278_));
  AOI21_X1   g12086(.A1(new_n12271_), .A2(new_n11992_), .B(new_n4330_), .ZN(new_n12279_));
  NOR2_X1    g12087(.A1(new_n12278_), .A2(new_n12279_), .ZN(new_n12280_));
  NAND2_X1   g12088(.A1(new_n12280_), .A2(new_n4018_), .ZN(new_n12281_));
  INV_X1     g12089(.I(new_n12281_), .ZN(new_n12282_));
  OAI21_X1   g12090(.A1(new_n12277_), .A2(new_n4330_), .B(new_n12282_), .ZN(new_n12283_));
  NAND2_X1   g12091(.A1(new_n12283_), .A2(new_n12276_), .ZN(new_n12284_));
  OAI22_X1   g12092(.A1(new_n12277_), .A2(new_n4330_), .B1(new_n12275_), .B2(new_n12269_), .ZN(new_n12285_));
  NAND2_X1   g12093(.A1(new_n12000_), .A2(\asqrt[40] ), .ZN(new_n12286_));
  NOR4_X1    g12094(.A1(new_n12101_), .A2(\asqrt[40] ), .A3(new_n11765_), .A4(new_n12000_), .ZN(new_n12287_));
  XOR2_X1    g12095(.A1(new_n12287_), .A2(new_n12286_), .Z(new_n12288_));
  NAND2_X1   g12096(.A1(new_n12288_), .A2(new_n3760_), .ZN(new_n12289_));
  AOI21_X1   g12097(.A1(new_n12285_), .A2(\asqrt[40] ), .B(new_n12289_), .ZN(new_n12290_));
  NOR2_X1    g12098(.A1(new_n12290_), .A2(new_n12284_), .ZN(new_n12291_));
  AOI22_X1   g12099(.A1(new_n12285_), .A2(\asqrt[40] ), .B1(new_n12283_), .B2(new_n12276_), .ZN(new_n12292_));
  NAND2_X1   g12100(.A1(new_n11777_), .A2(\asqrt[41] ), .ZN(new_n12293_));
  NOR4_X1    g12101(.A1(new_n12101_), .A2(\asqrt[41] ), .A3(new_n11772_), .A4(new_n11777_), .ZN(new_n12294_));
  XOR2_X1    g12102(.A1(new_n12294_), .A2(new_n12293_), .Z(new_n12295_));
  NAND2_X1   g12103(.A1(new_n12295_), .A2(new_n3481_), .ZN(new_n12296_));
  INV_X1     g12104(.I(new_n12296_), .ZN(new_n12297_));
  OAI21_X1   g12105(.A1(new_n12292_), .A2(new_n3760_), .B(new_n12297_), .ZN(new_n12298_));
  NAND2_X1   g12106(.A1(new_n12298_), .A2(new_n12291_), .ZN(new_n12299_));
  OAI22_X1   g12107(.A1(new_n12292_), .A2(new_n3760_), .B1(new_n12290_), .B2(new_n12284_), .ZN(new_n12300_));
  NOR4_X1    g12108(.A1(new_n12101_), .A2(\asqrt[42] ), .A3(new_n11780_), .A4(new_n12007_), .ZN(new_n12301_));
  AOI21_X1   g12109(.A1(new_n12293_), .A2(new_n11776_), .B(new_n3481_), .ZN(new_n12302_));
  NOR2_X1    g12110(.A1(new_n12301_), .A2(new_n12302_), .ZN(new_n12303_));
  NAND2_X1   g12111(.A1(new_n12303_), .A2(new_n3208_), .ZN(new_n12304_));
  AOI21_X1   g12112(.A1(new_n12300_), .A2(\asqrt[42] ), .B(new_n12304_), .ZN(new_n12305_));
  NOR2_X1    g12113(.A1(new_n12305_), .A2(new_n12299_), .ZN(new_n12306_));
  AOI22_X1   g12114(.A1(new_n12300_), .A2(\asqrt[42] ), .B1(new_n12298_), .B2(new_n12291_), .ZN(new_n12307_));
  NAND2_X1   g12115(.A1(new_n11792_), .A2(\asqrt[43] ), .ZN(new_n12308_));
  NOR4_X1    g12116(.A1(new_n12101_), .A2(\asqrt[43] ), .A3(new_n11787_), .A4(new_n11792_), .ZN(new_n12309_));
  XOR2_X1    g12117(.A1(new_n12309_), .A2(new_n12308_), .Z(new_n12310_));
  NAND2_X1   g12118(.A1(new_n12310_), .A2(new_n2941_), .ZN(new_n12311_));
  INV_X1     g12119(.I(new_n12311_), .ZN(new_n12312_));
  OAI21_X1   g12120(.A1(new_n12307_), .A2(new_n3208_), .B(new_n12312_), .ZN(new_n12313_));
  NAND2_X1   g12121(.A1(new_n12313_), .A2(new_n12306_), .ZN(new_n12314_));
  OAI22_X1   g12122(.A1(new_n12307_), .A2(new_n3208_), .B1(new_n12305_), .B2(new_n12299_), .ZN(new_n12315_));
  NOR4_X1    g12123(.A1(new_n12101_), .A2(\asqrt[44] ), .A3(new_n11795_), .A4(new_n12014_), .ZN(new_n12316_));
  AOI21_X1   g12124(.A1(new_n12308_), .A2(new_n11791_), .B(new_n2941_), .ZN(new_n12317_));
  NOR2_X1    g12125(.A1(new_n12316_), .A2(new_n12317_), .ZN(new_n12318_));
  NAND2_X1   g12126(.A1(new_n12318_), .A2(new_n2728_), .ZN(new_n12319_));
  AOI21_X1   g12127(.A1(new_n12315_), .A2(\asqrt[44] ), .B(new_n12319_), .ZN(new_n12320_));
  NOR2_X1    g12128(.A1(new_n12320_), .A2(new_n12314_), .ZN(new_n12321_));
  AOI22_X1   g12129(.A1(new_n12315_), .A2(\asqrt[44] ), .B1(new_n12313_), .B2(new_n12306_), .ZN(new_n12322_));
  NAND2_X1   g12130(.A1(new_n11807_), .A2(\asqrt[45] ), .ZN(new_n12323_));
  NOR4_X1    g12131(.A1(new_n12101_), .A2(\asqrt[45] ), .A3(new_n11802_), .A4(new_n11807_), .ZN(new_n12324_));
  XOR2_X1    g12132(.A1(new_n12324_), .A2(new_n12323_), .Z(new_n12325_));
  NAND2_X1   g12133(.A1(new_n12325_), .A2(new_n2488_), .ZN(new_n12326_));
  INV_X1     g12134(.I(new_n12326_), .ZN(new_n12327_));
  OAI21_X1   g12135(.A1(new_n12322_), .A2(new_n2728_), .B(new_n12327_), .ZN(new_n12328_));
  NAND2_X1   g12136(.A1(new_n12328_), .A2(new_n12321_), .ZN(new_n12329_));
  OAI22_X1   g12137(.A1(new_n12322_), .A2(new_n2728_), .B1(new_n12320_), .B2(new_n12314_), .ZN(new_n12330_));
  NOR4_X1    g12138(.A1(new_n12101_), .A2(\asqrt[46] ), .A3(new_n11810_), .A4(new_n12021_), .ZN(new_n12331_));
  AOI21_X1   g12139(.A1(new_n12323_), .A2(new_n11806_), .B(new_n2488_), .ZN(new_n12332_));
  NOR2_X1    g12140(.A1(new_n12331_), .A2(new_n12332_), .ZN(new_n12333_));
  NAND2_X1   g12141(.A1(new_n12333_), .A2(new_n2253_), .ZN(new_n12334_));
  AOI21_X1   g12142(.A1(new_n12330_), .A2(\asqrt[46] ), .B(new_n12334_), .ZN(new_n12335_));
  NOR2_X1    g12143(.A1(new_n12335_), .A2(new_n12329_), .ZN(new_n12336_));
  AOI22_X1   g12144(.A1(new_n12330_), .A2(\asqrt[46] ), .B1(new_n12328_), .B2(new_n12321_), .ZN(new_n12337_));
  NAND2_X1   g12145(.A1(new_n11822_), .A2(\asqrt[47] ), .ZN(new_n12338_));
  NOR4_X1    g12146(.A1(new_n12101_), .A2(\asqrt[47] ), .A3(new_n11817_), .A4(new_n11822_), .ZN(new_n12339_));
  XOR2_X1    g12147(.A1(new_n12339_), .A2(new_n12338_), .Z(new_n12340_));
  NAND2_X1   g12148(.A1(new_n12340_), .A2(new_n2046_), .ZN(new_n12341_));
  INV_X1     g12149(.I(new_n12341_), .ZN(new_n12342_));
  OAI21_X1   g12150(.A1(new_n12337_), .A2(new_n2253_), .B(new_n12342_), .ZN(new_n12343_));
  NAND2_X1   g12151(.A1(new_n12343_), .A2(new_n12336_), .ZN(new_n12344_));
  OAI22_X1   g12152(.A1(new_n12337_), .A2(new_n2253_), .B1(new_n12335_), .B2(new_n12329_), .ZN(new_n12345_));
  NAND2_X1   g12153(.A1(new_n12028_), .A2(\asqrt[48] ), .ZN(new_n12346_));
  NOR4_X1    g12154(.A1(new_n12101_), .A2(\asqrt[48] ), .A3(new_n11825_), .A4(new_n12028_), .ZN(new_n12347_));
  XOR2_X1    g12155(.A1(new_n12347_), .A2(new_n12346_), .Z(new_n12348_));
  NAND2_X1   g12156(.A1(new_n12348_), .A2(new_n1854_), .ZN(new_n12349_));
  AOI21_X1   g12157(.A1(new_n12345_), .A2(\asqrt[48] ), .B(new_n12349_), .ZN(new_n12350_));
  NOR2_X1    g12158(.A1(new_n12350_), .A2(new_n12344_), .ZN(new_n12351_));
  AOI22_X1   g12159(.A1(new_n12345_), .A2(\asqrt[48] ), .B1(new_n12343_), .B2(new_n12336_), .ZN(new_n12352_));
  NOR4_X1    g12160(.A1(new_n12101_), .A2(\asqrt[49] ), .A3(new_n11832_), .A4(new_n11837_), .ZN(new_n12353_));
  AOI21_X1   g12161(.A1(new_n12346_), .A2(new_n12027_), .B(new_n1854_), .ZN(new_n12354_));
  NOR2_X1    g12162(.A1(new_n12353_), .A2(new_n12354_), .ZN(new_n12355_));
  NAND2_X1   g12163(.A1(new_n12355_), .A2(new_n1595_), .ZN(new_n12356_));
  INV_X1     g12164(.I(new_n12356_), .ZN(new_n12357_));
  OAI21_X1   g12165(.A1(new_n12352_), .A2(new_n1854_), .B(new_n12357_), .ZN(new_n12358_));
  NAND2_X1   g12166(.A1(new_n12358_), .A2(new_n12351_), .ZN(new_n12359_));
  OAI22_X1   g12167(.A1(new_n12352_), .A2(new_n1854_), .B1(new_n12350_), .B2(new_n12344_), .ZN(new_n12360_));
  NAND2_X1   g12168(.A1(new_n12035_), .A2(\asqrt[50] ), .ZN(new_n12361_));
  NOR4_X1    g12169(.A1(new_n12101_), .A2(\asqrt[50] ), .A3(new_n11840_), .A4(new_n12035_), .ZN(new_n12362_));
  XOR2_X1    g12170(.A1(new_n12362_), .A2(new_n12361_), .Z(new_n12363_));
  NAND2_X1   g12171(.A1(new_n12363_), .A2(new_n1436_), .ZN(new_n12364_));
  AOI21_X1   g12172(.A1(new_n12360_), .A2(\asqrt[50] ), .B(new_n12364_), .ZN(new_n12365_));
  NOR2_X1    g12173(.A1(new_n12365_), .A2(new_n12359_), .ZN(new_n12366_));
  AOI22_X1   g12174(.A1(new_n12360_), .A2(\asqrt[50] ), .B1(new_n12358_), .B2(new_n12351_), .ZN(new_n12367_));
  NOR4_X1    g12175(.A1(new_n12101_), .A2(\asqrt[51] ), .A3(new_n11847_), .A4(new_n11852_), .ZN(new_n12368_));
  AOI21_X1   g12176(.A1(new_n12361_), .A2(new_n12034_), .B(new_n1436_), .ZN(new_n12369_));
  NOR2_X1    g12177(.A1(new_n12368_), .A2(new_n12369_), .ZN(new_n12370_));
  NAND2_X1   g12178(.A1(new_n12370_), .A2(new_n1260_), .ZN(new_n12371_));
  INV_X1     g12179(.I(new_n12371_), .ZN(new_n12372_));
  OAI21_X1   g12180(.A1(new_n12367_), .A2(new_n1436_), .B(new_n12372_), .ZN(new_n12373_));
  NAND2_X1   g12181(.A1(new_n12373_), .A2(new_n12366_), .ZN(new_n12374_));
  OAI22_X1   g12182(.A1(new_n12367_), .A2(new_n1436_), .B1(new_n12365_), .B2(new_n12359_), .ZN(new_n12375_));
  NAND2_X1   g12183(.A1(new_n12042_), .A2(\asqrt[52] ), .ZN(new_n12376_));
  NOR4_X1    g12184(.A1(new_n12101_), .A2(\asqrt[52] ), .A3(new_n11855_), .A4(new_n12042_), .ZN(new_n12377_));
  XOR2_X1    g12185(.A1(new_n12377_), .A2(new_n12376_), .Z(new_n12378_));
  NAND2_X1   g12186(.A1(new_n12378_), .A2(new_n1096_), .ZN(new_n12379_));
  AOI21_X1   g12187(.A1(new_n12375_), .A2(\asqrt[52] ), .B(new_n12379_), .ZN(new_n12380_));
  NOR2_X1    g12188(.A1(new_n12380_), .A2(new_n12374_), .ZN(new_n12381_));
  AOI22_X1   g12189(.A1(new_n12375_), .A2(\asqrt[52] ), .B1(new_n12373_), .B2(new_n12366_), .ZN(new_n12382_));
  NOR2_X1    g12190(.A1(new_n12045_), .A2(new_n1096_), .ZN(new_n12383_));
  NOR4_X1    g12191(.A1(new_n12101_), .A2(\asqrt[53] ), .A3(new_n11862_), .A4(new_n11867_), .ZN(new_n12384_));
  XNOR2_X1   g12192(.A1(new_n12384_), .A2(new_n12383_), .ZN(new_n12385_));
  NAND2_X1   g12193(.A1(new_n12385_), .A2(new_n970_), .ZN(new_n12386_));
  INV_X1     g12194(.I(new_n12386_), .ZN(new_n12387_));
  OAI21_X1   g12195(.A1(new_n12382_), .A2(new_n1096_), .B(new_n12387_), .ZN(new_n12388_));
  NAND2_X1   g12196(.A1(new_n12388_), .A2(new_n12381_), .ZN(new_n12389_));
  OAI22_X1   g12197(.A1(new_n12382_), .A2(new_n1096_), .B1(new_n12380_), .B2(new_n12374_), .ZN(new_n12390_));
  NOR4_X1    g12198(.A1(new_n12101_), .A2(\asqrt[54] ), .A3(new_n11869_), .A4(new_n12049_), .ZN(new_n12391_));
  XOR2_X1    g12199(.A1(new_n12391_), .A2(new_n12117_), .Z(new_n12392_));
  NAND2_X1   g12200(.A1(new_n12392_), .A2(new_n825_), .ZN(new_n12393_));
  AOI21_X1   g12201(.A1(new_n12390_), .A2(\asqrt[54] ), .B(new_n12393_), .ZN(new_n12394_));
  NOR2_X1    g12202(.A1(new_n12394_), .A2(new_n12389_), .ZN(new_n12395_));
  AOI22_X1   g12203(.A1(new_n12390_), .A2(\asqrt[54] ), .B1(new_n12388_), .B2(new_n12381_), .ZN(new_n12396_));
  NOR4_X1    g12204(.A1(new_n12101_), .A2(\asqrt[55] ), .A3(new_n11875_), .A4(new_n11880_), .ZN(new_n12397_));
  XOR2_X1    g12205(.A1(new_n12397_), .A2(new_n12102_), .Z(new_n12398_));
  NAND2_X1   g12206(.A1(new_n12398_), .A2(new_n724_), .ZN(new_n12399_));
  INV_X1     g12207(.I(new_n12399_), .ZN(new_n12400_));
  OAI21_X1   g12208(.A1(new_n12396_), .A2(new_n825_), .B(new_n12400_), .ZN(new_n12401_));
  NAND2_X1   g12209(.A1(new_n12401_), .A2(new_n12395_), .ZN(new_n12402_));
  OAI22_X1   g12210(.A1(new_n12396_), .A2(new_n825_), .B1(new_n12394_), .B2(new_n12389_), .ZN(new_n12403_));
  NOR4_X1    g12211(.A1(new_n12101_), .A2(\asqrt[56] ), .A3(new_n11882_), .A4(new_n12056_), .ZN(new_n12404_));
  XOR2_X1    g12212(.A1(new_n12404_), .A2(new_n12119_), .Z(new_n12405_));
  NAND2_X1   g12213(.A1(new_n12405_), .A2(new_n587_), .ZN(new_n12406_));
  AOI21_X1   g12214(.A1(new_n12403_), .A2(\asqrt[56] ), .B(new_n12406_), .ZN(new_n12407_));
  NOR2_X1    g12215(.A1(new_n12407_), .A2(new_n12402_), .ZN(new_n12408_));
  AOI22_X1   g12216(.A1(new_n12403_), .A2(\asqrt[56] ), .B1(new_n12401_), .B2(new_n12395_), .ZN(new_n12409_));
  NOR4_X1    g12217(.A1(new_n12101_), .A2(\asqrt[57] ), .A3(new_n11888_), .A4(new_n11893_), .ZN(new_n12410_));
  XOR2_X1    g12218(.A1(new_n12410_), .A2(new_n12104_), .Z(new_n12411_));
  NAND2_X1   g12219(.A1(new_n12411_), .A2(new_n504_), .ZN(new_n12412_));
  INV_X1     g12220(.I(new_n12412_), .ZN(new_n12413_));
  OAI21_X1   g12221(.A1(new_n12409_), .A2(new_n587_), .B(new_n12413_), .ZN(new_n12414_));
  NAND2_X1   g12222(.A1(new_n12414_), .A2(new_n12408_), .ZN(new_n12415_));
  OAI22_X1   g12223(.A1(new_n12409_), .A2(new_n587_), .B1(new_n12407_), .B2(new_n12402_), .ZN(new_n12416_));
  NOR4_X1    g12224(.A1(new_n12101_), .A2(\asqrt[58] ), .A3(new_n11895_), .A4(new_n12063_), .ZN(new_n12417_));
  XOR2_X1    g12225(.A1(new_n12417_), .A2(new_n12121_), .Z(new_n12418_));
  NAND2_X1   g12226(.A1(new_n12418_), .A2(new_n376_), .ZN(new_n12419_));
  AOI21_X1   g12227(.A1(new_n12416_), .A2(\asqrt[58] ), .B(new_n12419_), .ZN(new_n12420_));
  NOR2_X1    g12228(.A1(new_n12420_), .A2(new_n12415_), .ZN(new_n12421_));
  AOI22_X1   g12229(.A1(new_n12416_), .A2(\asqrt[58] ), .B1(new_n12414_), .B2(new_n12408_), .ZN(new_n12422_));
  NOR4_X1    g12230(.A1(new_n12101_), .A2(\asqrt[59] ), .A3(new_n11901_), .A4(new_n11906_), .ZN(new_n12423_));
  XOR2_X1    g12231(.A1(new_n12423_), .A2(new_n12106_), .Z(new_n12424_));
  AND2_X2    g12232(.A1(new_n12424_), .A2(new_n275_), .Z(new_n12425_));
  OAI21_X1   g12233(.A1(new_n12422_), .A2(new_n376_), .B(new_n12425_), .ZN(new_n12426_));
  NAND2_X1   g12234(.A1(new_n12426_), .A2(new_n12421_), .ZN(new_n12427_));
  NAND2_X1   g12235(.A1(new_n12390_), .A2(\asqrt[54] ), .ZN(new_n12428_));
  AOI21_X1   g12236(.A1(new_n12428_), .A2(new_n12389_), .B(new_n825_), .ZN(new_n12429_));
  OAI21_X1   g12237(.A1(new_n12395_), .A2(new_n12429_), .B(\asqrt[56] ), .ZN(new_n12430_));
  AOI21_X1   g12238(.A1(new_n12402_), .A2(new_n12430_), .B(new_n587_), .ZN(new_n12431_));
  OAI21_X1   g12239(.A1(new_n12408_), .A2(new_n12431_), .B(\asqrt[58] ), .ZN(new_n12432_));
  AOI21_X1   g12240(.A1(new_n12415_), .A2(new_n12432_), .B(new_n376_), .ZN(new_n12433_));
  OAI21_X1   g12241(.A1(new_n12421_), .A2(new_n12433_), .B(\asqrt[60] ), .ZN(new_n12434_));
  AOI21_X1   g12242(.A1(new_n12427_), .A2(new_n12434_), .B(new_n229_), .ZN(new_n12435_));
  NOR2_X1    g12243(.A1(new_n12088_), .A2(new_n196_), .ZN(new_n12436_));
  NOR2_X1    g12244(.A1(new_n12073_), .A2(\asqrt[62] ), .ZN(new_n12437_));
  NAND3_X1   g12245(.A1(new_n12437_), .A2(new_n12436_), .A3(new_n11920_), .ZN(new_n12438_));
  NOR2_X1    g12246(.A1(new_n12101_), .A2(new_n12438_), .ZN(new_n12439_));
  OR3_X2     g12247(.A1(\asqrt[20] ), .A2(new_n11920_), .A3(new_n12437_), .Z(new_n12440_));
  AOI21_X1   g12248(.A1(new_n12440_), .A2(new_n12436_), .B(new_n12439_), .ZN(new_n12441_));
  NOR4_X1    g12249(.A1(new_n12101_), .A2(\asqrt[61] ), .A3(new_n11914_), .A4(new_n11919_), .ZN(new_n12442_));
  XOR2_X1    g12250(.A1(new_n12442_), .A2(new_n12108_), .Z(new_n12443_));
  NOR2_X1    g12251(.A1(new_n12443_), .A2(new_n196_), .ZN(new_n12444_));
  INV_X1     g12252(.I(new_n12444_), .ZN(new_n12445_));
  NAND2_X1   g12253(.A1(new_n12156_), .A2(new_n12162_), .ZN(new_n12446_));
  NAND3_X1   g12254(.A1(new_n12446_), .A2(new_n12143_), .A3(new_n12179_), .ZN(new_n12447_));
  INV_X1     g12255(.I(new_n12080_), .ZN(new_n12448_));
  AOI21_X1   g12256(.A1(new_n12092_), .A2(new_n12448_), .B(new_n12082_), .ZN(new_n12449_));
  NOR3_X1    g12257(.A1(new_n12079_), .A2(new_n11566_), .A3(new_n11578_), .ZN(new_n12450_));
  NOR2_X1    g12258(.A1(new_n12450_), .A2(new_n12449_), .ZN(new_n12451_));
  NOR3_X1    g12259(.A1(new_n12129_), .A2(new_n11607_), .A3(\asqrt[20] ), .ZN(new_n12452_));
  AOI21_X1   g12260(.A1(new_n12114_), .A2(new_n11606_), .B(new_n12101_), .ZN(new_n12453_));
  NOR4_X1    g12261(.A1(new_n12452_), .A2(new_n12453_), .A3(\asqrt[22] ), .A4(new_n12099_), .ZN(new_n12454_));
  NOR2_X1    g12262(.A1(new_n12454_), .A2(new_n12451_), .ZN(new_n12455_));
  NOR3_X1    g12263(.A1(new_n12450_), .A2(new_n12449_), .A3(new_n12099_), .ZN(new_n12456_));
  NOR3_X1    g12264(.A1(new_n12101_), .A2(new_n11629_), .A3(new_n12137_), .ZN(new_n12457_));
  AOI21_X1   g12265(.A1(\asqrt[20] ), .A2(new_n12138_), .B(new_n11630_), .ZN(new_n12458_));
  NOR3_X1    g12266(.A1(new_n12457_), .A2(new_n12458_), .A3(\asqrt[23] ), .ZN(new_n12459_));
  OAI21_X1   g12267(.A1(new_n12456_), .A2(new_n11105_), .B(new_n12459_), .ZN(new_n12460_));
  NAND2_X1   g12268(.A1(new_n12455_), .A2(new_n12460_), .ZN(new_n12461_));
  OAI22_X1   g12269(.A1(new_n12454_), .A2(new_n12451_), .B1(new_n11105_), .B2(new_n12456_), .ZN(new_n12462_));
  AOI21_X1   g12270(.A1(new_n12462_), .A2(\asqrt[23] ), .B(new_n12154_), .ZN(new_n12463_));
  AOI22_X1   g12271(.A1(new_n12462_), .A2(\asqrt[23] ), .B1(new_n12455_), .B2(new_n12460_), .ZN(new_n12464_));
  OAI22_X1   g12272(.A1(new_n12464_), .A2(new_n10104_), .B1(new_n12463_), .B2(new_n12461_), .ZN(new_n12465_));
  AOI21_X1   g12273(.A1(new_n12465_), .A2(\asqrt[25] ), .B(new_n12169_), .ZN(new_n12466_));
  NOR2_X1    g12274(.A1(new_n12466_), .A2(new_n12447_), .ZN(new_n12467_));
  NAND2_X1   g12275(.A1(new_n12171_), .A2(new_n12176_), .ZN(new_n12468_));
  NAND2_X1   g12276(.A1(new_n12468_), .A2(new_n12467_), .ZN(new_n12469_));
  NOR2_X1    g12277(.A1(new_n12163_), .A2(new_n12164_), .ZN(new_n12470_));
  OAI22_X1   g12278(.A1(new_n12470_), .A2(new_n9212_), .B1(new_n12466_), .B2(new_n12447_), .ZN(new_n12471_));
  AOI21_X1   g12279(.A1(new_n12471_), .A2(\asqrt[27] ), .B(new_n12190_), .ZN(new_n12472_));
  NOR2_X1    g12280(.A1(new_n12472_), .A2(new_n12469_), .ZN(new_n12473_));
  AOI21_X1   g12281(.A1(new_n12170_), .A2(new_n12171_), .B(new_n8763_), .ZN(new_n12474_));
  OAI21_X1   g12282(.A1(new_n12177_), .A2(new_n12474_), .B(\asqrt[28] ), .ZN(new_n12475_));
  INV_X1     g12283(.I(new_n12199_), .ZN(new_n12476_));
  NAND2_X1   g12284(.A1(new_n12475_), .A2(new_n12476_), .ZN(new_n12477_));
  NAND2_X1   g12285(.A1(new_n12477_), .A2(new_n12473_), .ZN(new_n12478_));
  AOI22_X1   g12286(.A1(new_n12471_), .A2(\asqrt[27] ), .B1(new_n12468_), .B2(new_n12467_), .ZN(new_n12479_));
  OAI22_X1   g12287(.A1(new_n12479_), .A2(new_n8319_), .B1(new_n12472_), .B2(new_n12469_), .ZN(new_n12480_));
  AOI21_X1   g12288(.A1(new_n12480_), .A2(\asqrt[29] ), .B(new_n12206_), .ZN(new_n12481_));
  NOR2_X1    g12289(.A1(new_n12481_), .A2(new_n12478_), .ZN(new_n12482_));
  AOI22_X1   g12290(.A1(new_n12480_), .A2(\asqrt[29] ), .B1(new_n12477_), .B2(new_n12473_), .ZN(new_n12483_));
  INV_X1     g12291(.I(new_n12214_), .ZN(new_n12484_));
  OAI21_X1   g12292(.A1(new_n12483_), .A2(new_n7517_), .B(new_n12484_), .ZN(new_n12485_));
  NAND2_X1   g12293(.A1(new_n12485_), .A2(new_n12482_), .ZN(new_n12486_));
  OAI22_X1   g12294(.A1(new_n12483_), .A2(new_n7517_), .B1(new_n12481_), .B2(new_n12478_), .ZN(new_n12487_));
  AOI21_X1   g12295(.A1(new_n12487_), .A2(\asqrt[31] ), .B(new_n12221_), .ZN(new_n12488_));
  NOR2_X1    g12296(.A1(new_n12488_), .A2(new_n12486_), .ZN(new_n12489_));
  AOI22_X1   g12297(.A1(new_n12487_), .A2(\asqrt[31] ), .B1(new_n12485_), .B2(new_n12482_), .ZN(new_n12490_));
  INV_X1     g12298(.I(new_n12229_), .ZN(new_n12491_));
  OAI21_X1   g12299(.A1(new_n12490_), .A2(new_n6708_), .B(new_n12491_), .ZN(new_n12492_));
  NAND2_X1   g12300(.A1(new_n12492_), .A2(new_n12489_), .ZN(new_n12493_));
  OAI22_X1   g12301(.A1(new_n12490_), .A2(new_n6708_), .B1(new_n12488_), .B2(new_n12486_), .ZN(new_n12494_));
  AOI21_X1   g12302(.A1(new_n12494_), .A2(\asqrt[33] ), .B(new_n12236_), .ZN(new_n12495_));
  NOR2_X1    g12303(.A1(new_n12495_), .A2(new_n12493_), .ZN(new_n12496_));
  AOI22_X1   g12304(.A1(new_n12494_), .A2(\asqrt[33] ), .B1(new_n12492_), .B2(new_n12489_), .ZN(new_n12497_));
  INV_X1     g12305(.I(new_n12244_), .ZN(new_n12498_));
  OAI21_X1   g12306(.A1(new_n12497_), .A2(new_n5991_), .B(new_n12498_), .ZN(new_n12499_));
  NAND2_X1   g12307(.A1(new_n12499_), .A2(new_n12496_), .ZN(new_n12500_));
  OAI22_X1   g12308(.A1(new_n12497_), .A2(new_n5991_), .B1(new_n12495_), .B2(new_n12493_), .ZN(new_n12501_));
  AOI21_X1   g12309(.A1(new_n12501_), .A2(\asqrt[35] ), .B(new_n12251_), .ZN(new_n12502_));
  NOR2_X1    g12310(.A1(new_n12502_), .A2(new_n12500_), .ZN(new_n12503_));
  AOI22_X1   g12311(.A1(new_n12501_), .A2(\asqrt[35] ), .B1(new_n12499_), .B2(new_n12496_), .ZN(new_n12504_));
  INV_X1     g12312(.I(new_n12259_), .ZN(new_n12505_));
  OAI21_X1   g12313(.A1(new_n12504_), .A2(new_n5273_), .B(new_n12505_), .ZN(new_n12506_));
  NAND2_X1   g12314(.A1(new_n12506_), .A2(new_n12503_), .ZN(new_n12507_));
  OAI22_X1   g12315(.A1(new_n12504_), .A2(new_n5273_), .B1(new_n12502_), .B2(new_n12500_), .ZN(new_n12508_));
  AOI21_X1   g12316(.A1(new_n12508_), .A2(\asqrt[37] ), .B(new_n12266_), .ZN(new_n12509_));
  NOR2_X1    g12317(.A1(new_n12509_), .A2(new_n12507_), .ZN(new_n12510_));
  AOI22_X1   g12318(.A1(new_n12508_), .A2(\asqrt[37] ), .B1(new_n12506_), .B2(new_n12503_), .ZN(new_n12511_));
  INV_X1     g12319(.I(new_n12274_), .ZN(new_n12512_));
  OAI21_X1   g12320(.A1(new_n12511_), .A2(new_n4645_), .B(new_n12512_), .ZN(new_n12513_));
  NAND2_X1   g12321(.A1(new_n12513_), .A2(new_n12510_), .ZN(new_n12514_));
  OAI22_X1   g12322(.A1(new_n12511_), .A2(new_n4645_), .B1(new_n12509_), .B2(new_n12507_), .ZN(new_n12515_));
  AOI21_X1   g12323(.A1(new_n12515_), .A2(\asqrt[39] ), .B(new_n12281_), .ZN(new_n12516_));
  NOR2_X1    g12324(.A1(new_n12516_), .A2(new_n12514_), .ZN(new_n12517_));
  AOI22_X1   g12325(.A1(new_n12515_), .A2(\asqrt[39] ), .B1(new_n12513_), .B2(new_n12510_), .ZN(new_n12518_));
  INV_X1     g12326(.I(new_n12289_), .ZN(new_n12519_));
  OAI21_X1   g12327(.A1(new_n12518_), .A2(new_n4018_), .B(new_n12519_), .ZN(new_n12520_));
  NAND2_X1   g12328(.A1(new_n12520_), .A2(new_n12517_), .ZN(new_n12521_));
  OAI22_X1   g12329(.A1(new_n12518_), .A2(new_n4018_), .B1(new_n12516_), .B2(new_n12514_), .ZN(new_n12522_));
  AOI21_X1   g12330(.A1(new_n12522_), .A2(\asqrt[41] ), .B(new_n12296_), .ZN(new_n12523_));
  NOR2_X1    g12331(.A1(new_n12523_), .A2(new_n12521_), .ZN(new_n12524_));
  AOI22_X1   g12332(.A1(new_n12522_), .A2(\asqrt[41] ), .B1(new_n12520_), .B2(new_n12517_), .ZN(new_n12525_));
  INV_X1     g12333(.I(new_n12304_), .ZN(new_n12526_));
  OAI21_X1   g12334(.A1(new_n12525_), .A2(new_n3481_), .B(new_n12526_), .ZN(new_n12527_));
  NAND2_X1   g12335(.A1(new_n12527_), .A2(new_n12524_), .ZN(new_n12528_));
  OAI22_X1   g12336(.A1(new_n12525_), .A2(new_n3481_), .B1(new_n12523_), .B2(new_n12521_), .ZN(new_n12529_));
  AOI21_X1   g12337(.A1(new_n12529_), .A2(\asqrt[43] ), .B(new_n12311_), .ZN(new_n12530_));
  NOR2_X1    g12338(.A1(new_n12530_), .A2(new_n12528_), .ZN(new_n12531_));
  AOI22_X1   g12339(.A1(new_n12529_), .A2(\asqrt[43] ), .B1(new_n12527_), .B2(new_n12524_), .ZN(new_n12532_));
  INV_X1     g12340(.I(new_n12319_), .ZN(new_n12533_));
  OAI21_X1   g12341(.A1(new_n12532_), .A2(new_n2941_), .B(new_n12533_), .ZN(new_n12534_));
  NAND2_X1   g12342(.A1(new_n12534_), .A2(new_n12531_), .ZN(new_n12535_));
  OAI22_X1   g12343(.A1(new_n12532_), .A2(new_n2941_), .B1(new_n12530_), .B2(new_n12528_), .ZN(new_n12536_));
  AOI21_X1   g12344(.A1(new_n12536_), .A2(\asqrt[45] ), .B(new_n12326_), .ZN(new_n12537_));
  NOR2_X1    g12345(.A1(new_n12537_), .A2(new_n12535_), .ZN(new_n12538_));
  AOI22_X1   g12346(.A1(new_n12536_), .A2(\asqrt[45] ), .B1(new_n12534_), .B2(new_n12531_), .ZN(new_n12539_));
  INV_X1     g12347(.I(new_n12334_), .ZN(new_n12540_));
  OAI21_X1   g12348(.A1(new_n12539_), .A2(new_n2488_), .B(new_n12540_), .ZN(new_n12541_));
  NAND2_X1   g12349(.A1(new_n12541_), .A2(new_n12538_), .ZN(new_n12542_));
  OAI22_X1   g12350(.A1(new_n12539_), .A2(new_n2488_), .B1(new_n12537_), .B2(new_n12535_), .ZN(new_n12543_));
  AOI21_X1   g12351(.A1(new_n12543_), .A2(\asqrt[47] ), .B(new_n12341_), .ZN(new_n12544_));
  NOR2_X1    g12352(.A1(new_n12544_), .A2(new_n12542_), .ZN(new_n12545_));
  AOI22_X1   g12353(.A1(new_n12543_), .A2(\asqrt[47] ), .B1(new_n12541_), .B2(new_n12538_), .ZN(new_n12546_));
  INV_X1     g12354(.I(new_n12349_), .ZN(new_n12547_));
  OAI21_X1   g12355(.A1(new_n12546_), .A2(new_n2046_), .B(new_n12547_), .ZN(new_n12548_));
  NAND2_X1   g12356(.A1(new_n12548_), .A2(new_n12545_), .ZN(new_n12549_));
  OAI22_X1   g12357(.A1(new_n12546_), .A2(new_n2046_), .B1(new_n12544_), .B2(new_n12542_), .ZN(new_n12550_));
  AOI21_X1   g12358(.A1(new_n12550_), .A2(\asqrt[49] ), .B(new_n12356_), .ZN(new_n12551_));
  NOR2_X1    g12359(.A1(new_n12551_), .A2(new_n12549_), .ZN(new_n12552_));
  AOI22_X1   g12360(.A1(new_n12550_), .A2(\asqrt[49] ), .B1(new_n12548_), .B2(new_n12545_), .ZN(new_n12553_));
  INV_X1     g12361(.I(new_n12364_), .ZN(new_n12554_));
  OAI21_X1   g12362(.A1(new_n12553_), .A2(new_n1595_), .B(new_n12554_), .ZN(new_n12555_));
  NAND2_X1   g12363(.A1(new_n12555_), .A2(new_n12552_), .ZN(new_n12556_));
  OAI22_X1   g12364(.A1(new_n12553_), .A2(new_n1595_), .B1(new_n12551_), .B2(new_n12549_), .ZN(new_n12557_));
  AOI21_X1   g12365(.A1(new_n12557_), .A2(\asqrt[51] ), .B(new_n12371_), .ZN(new_n12558_));
  NOR2_X1    g12366(.A1(new_n12558_), .A2(new_n12556_), .ZN(new_n12559_));
  AOI22_X1   g12367(.A1(new_n12557_), .A2(\asqrt[51] ), .B1(new_n12555_), .B2(new_n12552_), .ZN(new_n12560_));
  INV_X1     g12368(.I(new_n12379_), .ZN(new_n12561_));
  OAI21_X1   g12369(.A1(new_n12560_), .A2(new_n1260_), .B(new_n12561_), .ZN(new_n12562_));
  NAND2_X1   g12370(.A1(new_n12562_), .A2(new_n12559_), .ZN(new_n12563_));
  OAI22_X1   g12371(.A1(new_n12560_), .A2(new_n1260_), .B1(new_n12558_), .B2(new_n12556_), .ZN(new_n12564_));
  AOI21_X1   g12372(.A1(new_n12564_), .A2(\asqrt[53] ), .B(new_n12386_), .ZN(new_n12565_));
  NOR2_X1    g12373(.A1(new_n12565_), .A2(new_n12563_), .ZN(new_n12566_));
  AOI22_X1   g12374(.A1(new_n12564_), .A2(\asqrt[53] ), .B1(new_n12562_), .B2(new_n12559_), .ZN(new_n12567_));
  INV_X1     g12375(.I(new_n12393_), .ZN(new_n12568_));
  OAI21_X1   g12376(.A1(new_n12567_), .A2(new_n970_), .B(new_n12568_), .ZN(new_n12569_));
  NAND2_X1   g12377(.A1(new_n12569_), .A2(new_n12566_), .ZN(new_n12570_));
  OAI22_X1   g12378(.A1(new_n12567_), .A2(new_n970_), .B1(new_n12565_), .B2(new_n12563_), .ZN(new_n12571_));
  AOI21_X1   g12379(.A1(new_n12571_), .A2(\asqrt[55] ), .B(new_n12399_), .ZN(new_n12572_));
  NOR2_X1    g12380(.A1(new_n12572_), .A2(new_n12570_), .ZN(new_n12573_));
  AOI22_X1   g12381(.A1(new_n12571_), .A2(\asqrt[55] ), .B1(new_n12569_), .B2(new_n12566_), .ZN(new_n12574_));
  INV_X1     g12382(.I(new_n12406_), .ZN(new_n12575_));
  OAI21_X1   g12383(.A1(new_n12574_), .A2(new_n724_), .B(new_n12575_), .ZN(new_n12576_));
  NAND2_X1   g12384(.A1(new_n12576_), .A2(new_n12573_), .ZN(new_n12577_));
  NAND2_X1   g12385(.A1(new_n12564_), .A2(\asqrt[53] ), .ZN(new_n12578_));
  AOI21_X1   g12386(.A1(new_n12578_), .A2(new_n12563_), .B(new_n970_), .ZN(new_n12579_));
  OAI21_X1   g12387(.A1(new_n12566_), .A2(new_n12579_), .B(\asqrt[55] ), .ZN(new_n12580_));
  AOI21_X1   g12388(.A1(new_n12570_), .A2(new_n12580_), .B(new_n724_), .ZN(new_n12581_));
  OAI21_X1   g12389(.A1(new_n12573_), .A2(new_n12581_), .B(\asqrt[57] ), .ZN(new_n12582_));
  AOI21_X1   g12390(.A1(new_n12582_), .A2(new_n12413_), .B(new_n12577_), .ZN(new_n12583_));
  OAI22_X1   g12391(.A1(new_n12574_), .A2(new_n724_), .B1(new_n12572_), .B2(new_n12570_), .ZN(new_n12584_));
  AOI22_X1   g12392(.A1(new_n12584_), .A2(\asqrt[57] ), .B1(new_n12576_), .B2(new_n12573_), .ZN(new_n12585_));
  INV_X1     g12393(.I(new_n12419_), .ZN(new_n12586_));
  OAI21_X1   g12394(.A1(new_n12585_), .A2(new_n504_), .B(new_n12586_), .ZN(new_n12587_));
  NAND2_X1   g12395(.A1(new_n12587_), .A2(new_n12583_), .ZN(new_n12588_));
  AOI21_X1   g12396(.A1(new_n12577_), .A2(new_n12582_), .B(new_n504_), .ZN(new_n12589_));
  OAI21_X1   g12397(.A1(new_n12583_), .A2(new_n12589_), .B(\asqrt[59] ), .ZN(new_n12590_));
  AOI21_X1   g12398(.A1(new_n12590_), .A2(new_n12425_), .B(new_n12588_), .ZN(new_n12591_));
  NAND2_X1   g12399(.A1(new_n12415_), .A2(new_n12432_), .ZN(new_n12592_));
  AOI22_X1   g12400(.A1(new_n12592_), .A2(\asqrt[59] ), .B1(new_n12587_), .B2(new_n12583_), .ZN(new_n12593_));
  NOR4_X1    g12401(.A1(new_n12101_), .A2(\asqrt[60] ), .A3(new_n11908_), .A4(new_n12070_), .ZN(new_n12594_));
  XOR2_X1    g12402(.A1(new_n12594_), .A2(new_n12123_), .Z(new_n12595_));
  NAND2_X1   g12403(.A1(new_n12595_), .A2(new_n229_), .ZN(new_n12596_));
  INV_X1     g12404(.I(new_n12596_), .ZN(new_n12597_));
  OAI21_X1   g12405(.A1(new_n12593_), .A2(new_n275_), .B(new_n12597_), .ZN(new_n12598_));
  NAND2_X1   g12406(.A1(new_n12598_), .A2(new_n12591_), .ZN(new_n12599_));
  INV_X1     g12407(.I(new_n12443_), .ZN(new_n12600_));
  NOR2_X1    g12408(.A1(new_n12600_), .A2(\asqrt[62] ), .ZN(new_n12601_));
  INV_X1     g12409(.I(new_n12601_), .ZN(new_n12602_));
  NAND2_X1   g12410(.A1(new_n12435_), .A2(new_n12602_), .ZN(new_n12603_));
  OAI21_X1   g12411(.A1(new_n12603_), .A2(new_n12599_), .B(new_n12445_), .ZN(new_n12604_));
  NOR3_X1    g12412(.A1(\asqrt[20] ), .A2(new_n11599_), .A3(new_n12074_), .ZN(new_n12605_));
  OAI21_X1   g12413(.A1(new_n12605_), .A2(new_n12086_), .B(new_n231_), .ZN(new_n12606_));
  OAI21_X1   g12414(.A1(new_n12604_), .A2(new_n12606_), .B(new_n12441_), .ZN(new_n12607_));
  OAI21_X1   g12415(.A1(new_n11599_), .A2(new_n11924_), .B(\asqrt[20] ), .ZN(new_n12608_));
  XOR2_X1    g12416(.A1(new_n11924_), .A2(\asqrt[63] ), .Z(new_n12609_));
  NAND2_X1   g12417(.A1(new_n12608_), .A2(new_n12609_), .ZN(new_n12610_));
  INV_X1     g12418(.I(new_n12610_), .ZN(new_n12611_));
  INV_X1     g12419(.I(new_n12441_), .ZN(new_n12612_));
  OAI22_X1   g12420(.A1(new_n12422_), .A2(new_n376_), .B1(new_n12420_), .B2(new_n12415_), .ZN(new_n12613_));
  AOI21_X1   g12421(.A1(new_n12613_), .A2(\asqrt[60] ), .B(new_n12596_), .ZN(new_n12614_));
  AOI22_X1   g12422(.A1(new_n12613_), .A2(\asqrt[60] ), .B1(new_n12426_), .B2(new_n12421_), .ZN(new_n12615_));
  OAI22_X1   g12423(.A1(new_n12615_), .A2(new_n229_), .B1(new_n12614_), .B2(new_n12427_), .ZN(new_n12616_));
  NOR4_X1    g12424(.A1(new_n12616_), .A2(\asqrt[62] ), .A3(new_n12612_), .A4(new_n12443_), .ZN(new_n12617_));
  NAND2_X1   g12425(.A1(new_n12617_), .A2(new_n12611_), .ZN(new_n12618_));
  NAND3_X1   g12426(.A1(new_n12095_), .A2(new_n11586_), .A3(new_n11599_), .ZN(new_n12619_));
  NOR3_X1    g12427(.A1(new_n12618_), .A2(new_n12607_), .A3(new_n12619_), .ZN(\asqrt[19] ));
  NAND2_X1   g12428(.A1(new_n12427_), .A2(new_n12434_), .ZN(new_n12621_));
  NOR3_X1    g12429(.A1(new_n12621_), .A2(\asqrt[61] ), .A3(new_n12595_), .ZN(new_n12622_));
  NAND2_X1   g12430(.A1(\asqrt[19] ), .A2(new_n12622_), .ZN(new_n12623_));
  XOR2_X1    g12431(.A1(new_n12623_), .A2(new_n12435_), .Z(new_n12624_));
  INV_X1     g12432(.I(new_n12624_), .ZN(new_n12625_));
  INV_X1     g12433(.I(\a[38] ), .ZN(new_n12626_));
  NOR2_X1    g12434(.A1(\a[36] ), .A2(\a[37] ), .ZN(new_n12627_));
  INV_X1     g12435(.I(new_n12627_), .ZN(new_n12628_));
  NOR3_X1    g12436(.A1(new_n12112_), .A2(new_n12626_), .A3(new_n12628_), .ZN(new_n12629_));
  NAND2_X1   g12437(.A1(new_n12127_), .A2(new_n12629_), .ZN(new_n12630_));
  XOR2_X1    g12438(.A1(new_n12630_), .A2(\a[39] ), .Z(new_n12631_));
  INV_X1     g12439(.I(\a[39] ), .ZN(new_n12632_));
  NOR4_X1    g12440(.A1(new_n12618_), .A2(new_n12607_), .A3(new_n12632_), .A4(new_n12619_), .ZN(new_n12633_));
  NOR2_X1    g12441(.A1(new_n12632_), .A2(\a[38] ), .ZN(new_n12634_));
  OAI21_X1   g12442(.A1(new_n12633_), .A2(new_n12634_), .B(new_n12631_), .ZN(new_n12635_));
  INV_X1     g12443(.I(new_n12631_), .ZN(new_n12636_));
  NOR2_X1    g12444(.A1(new_n12614_), .A2(new_n12427_), .ZN(new_n12637_));
  NOR3_X1    g12445(.A1(new_n12615_), .A2(new_n229_), .A3(new_n12601_), .ZN(new_n12638_));
  AOI21_X1   g12446(.A1(new_n12638_), .A2(new_n12637_), .B(new_n12444_), .ZN(new_n12639_));
  INV_X1     g12447(.I(new_n12606_), .ZN(new_n12640_));
  AOI21_X1   g12448(.A1(new_n12639_), .A2(new_n12640_), .B(new_n12612_), .ZN(new_n12641_));
  AOI21_X1   g12449(.A1(new_n12616_), .A2(\asqrt[62] ), .B(new_n12441_), .ZN(new_n12642_));
  AOI21_X1   g12450(.A1(new_n12588_), .A2(new_n12590_), .B(new_n275_), .ZN(new_n12643_));
  OAI21_X1   g12451(.A1(new_n12591_), .A2(new_n12643_), .B(\asqrt[61] ), .ZN(new_n12644_));
  NAND4_X1   g12452(.A1(new_n12599_), .A2(new_n196_), .A3(new_n12644_), .A4(new_n12600_), .ZN(new_n12645_));
  NOR3_X1    g12453(.A1(new_n12642_), .A2(new_n12610_), .A3(new_n12645_), .ZN(new_n12646_));
  INV_X1     g12454(.I(new_n12619_), .ZN(new_n12647_));
  NAND4_X1   g12455(.A1(new_n12646_), .A2(\a[39] ), .A3(new_n12641_), .A4(new_n12647_), .ZN(new_n12648_));
  NAND3_X1   g12456(.A1(new_n12648_), .A2(\a[38] ), .A3(new_n12636_), .ZN(new_n12649_));
  NAND2_X1   g12457(.A1(new_n12635_), .A2(new_n12649_), .ZN(new_n12650_));
  NOR2_X1    g12458(.A1(new_n12618_), .A2(new_n12607_), .ZN(new_n12651_));
  NAND4_X1   g12459(.A1(new_n12091_), .A2(new_n12083_), .A3(new_n11599_), .A4(new_n12126_), .ZN(new_n12652_));
  NOR2_X1    g12460(.A1(new_n12101_), .A2(new_n12626_), .ZN(new_n12653_));
  XOR2_X1    g12461(.A1(new_n12653_), .A2(new_n12652_), .Z(new_n12654_));
  NOR2_X1    g12462(.A1(new_n12654_), .A2(new_n12628_), .ZN(new_n12655_));
  INV_X1     g12463(.I(new_n12655_), .ZN(new_n12656_));
  NAND3_X1   g12464(.A1(new_n12646_), .A2(new_n12641_), .A3(new_n12647_), .ZN(new_n12657_));
  NOR4_X1    g12465(.A1(new_n12644_), .A2(new_n12427_), .A3(new_n12614_), .A4(new_n12601_), .ZN(new_n12658_));
  NOR3_X1    g12466(.A1(new_n12658_), .A2(new_n12444_), .A3(new_n12606_), .ZN(new_n12659_));
  AOI22_X1   g12467(.A1(new_n12621_), .A2(\asqrt[61] ), .B1(new_n12598_), .B2(new_n12591_), .ZN(new_n12660_));
  NAND4_X1   g12468(.A1(new_n12660_), .A2(new_n196_), .A3(new_n12441_), .A4(new_n12600_), .ZN(new_n12661_));
  OAI21_X1   g12469(.A1(new_n12659_), .A2(new_n12612_), .B(new_n12661_), .ZN(new_n12662_));
  NOR2_X1    g12470(.A1(new_n12611_), .A2(new_n12647_), .ZN(new_n12663_));
  NAND2_X1   g12471(.A1(new_n12663_), .A2(\asqrt[20] ), .ZN(new_n12664_));
  OAI21_X1   g12472(.A1(new_n12662_), .A2(new_n12664_), .B(new_n11566_), .ZN(new_n12665_));
  NAND3_X1   g12473(.A1(new_n12665_), .A2(new_n11574_), .A3(new_n12657_), .ZN(new_n12666_));
  NAND4_X1   g12474(.A1(new_n12435_), .A2(new_n12591_), .A3(new_n12598_), .A4(new_n12602_), .ZN(new_n12667_));
  NAND3_X1   g12475(.A1(new_n12667_), .A2(new_n12445_), .A3(new_n12640_), .ZN(new_n12668_));
  AOI21_X1   g12476(.A1(new_n12441_), .A2(new_n12668_), .B(new_n12617_), .ZN(new_n12669_));
  INV_X1     g12477(.I(new_n12664_), .ZN(new_n12670_));
  AOI21_X1   g12478(.A1(new_n12669_), .A2(new_n12670_), .B(\a[40] ), .ZN(new_n12671_));
  OAI21_X1   g12479(.A1(new_n12671_), .A2(new_n11575_), .B(\asqrt[19] ), .ZN(new_n12672_));
  NAND4_X1   g12480(.A1(new_n12666_), .A2(new_n12672_), .A3(new_n11631_), .A4(new_n12656_), .ZN(new_n12673_));
  NAND2_X1   g12481(.A1(new_n12673_), .A2(new_n12650_), .ZN(new_n12674_));
  NAND3_X1   g12482(.A1(new_n12635_), .A2(new_n12649_), .A3(new_n12656_), .ZN(new_n12675_));
  INV_X1     g12483(.I(new_n11577_), .ZN(new_n12676_));
  NOR2_X1    g12484(.A1(new_n12101_), .A2(\a[40] ), .ZN(new_n12677_));
  OAI22_X1   g12485(.A1(new_n12677_), .A2(\a[41] ), .B1(\a[40] ), .B2(new_n12092_), .ZN(new_n12678_));
  NAND2_X1   g12486(.A1(\asqrt[20] ), .A2(\a[40] ), .ZN(new_n12679_));
  AND3_X2    g12487(.A1(new_n12678_), .A2(new_n12676_), .A3(new_n12679_), .Z(new_n12680_));
  NAND3_X1   g12488(.A1(\asqrt[19] ), .A2(new_n12100_), .A3(new_n12680_), .ZN(new_n12681_));
  INV_X1     g12489(.I(new_n12680_), .ZN(new_n12682_));
  OAI21_X1   g12490(.A1(new_n12657_), .A2(new_n12682_), .B(new_n12099_), .ZN(new_n12683_));
  NAND3_X1   g12491(.A1(new_n12681_), .A2(new_n12683_), .A3(new_n11105_), .ZN(new_n12684_));
  AOI21_X1   g12492(.A1(new_n12675_), .A2(\asqrt[21] ), .B(new_n12684_), .ZN(new_n12685_));
  NOR2_X1    g12493(.A1(new_n12674_), .A2(new_n12685_), .ZN(new_n12686_));
  AOI22_X1   g12494(.A1(new_n12673_), .A2(new_n12650_), .B1(\asqrt[21] ), .B2(new_n12675_), .ZN(new_n12687_));
  AOI21_X1   g12495(.A1(new_n12130_), .A2(new_n12115_), .B(\asqrt[22] ), .ZN(new_n12688_));
  AND4_X2    g12496(.A1(new_n12456_), .A2(\asqrt[19] ), .A3(new_n12144_), .A4(new_n12688_), .Z(new_n12689_));
  NOR2_X1    g12497(.A1(new_n12456_), .A2(new_n11105_), .ZN(new_n12690_));
  NOR3_X1    g12498(.A1(new_n12689_), .A2(\asqrt[23] ), .A3(new_n12690_), .ZN(new_n12691_));
  OAI21_X1   g12499(.A1(new_n12687_), .A2(new_n11105_), .B(new_n12691_), .ZN(new_n12692_));
  NAND2_X1   g12500(.A1(new_n12692_), .A2(new_n12686_), .ZN(new_n12693_));
  OAI22_X1   g12501(.A1(new_n12687_), .A2(new_n11105_), .B1(new_n12674_), .B2(new_n12685_), .ZN(new_n12694_));
  NAND2_X1   g12502(.A1(new_n12140_), .A2(new_n12139_), .ZN(new_n12695_));
  NAND4_X1   g12503(.A1(\asqrt[19] ), .A2(new_n10614_), .A3(new_n12695_), .A4(new_n12178_), .ZN(new_n12696_));
  XOR2_X1    g12504(.A1(new_n12696_), .A2(new_n12145_), .Z(new_n12697_));
  NAND2_X1   g12505(.A1(new_n12697_), .A2(new_n10104_), .ZN(new_n12698_));
  AOI21_X1   g12506(.A1(new_n12694_), .A2(\asqrt[23] ), .B(new_n12698_), .ZN(new_n12699_));
  NOR2_X1    g12507(.A1(new_n12699_), .A2(new_n12693_), .ZN(new_n12700_));
  AOI22_X1   g12508(.A1(new_n12694_), .A2(\asqrt[23] ), .B1(new_n12692_), .B2(new_n12686_), .ZN(new_n12701_));
  NOR2_X1    g12509(.A1(new_n12152_), .A2(new_n12150_), .ZN(new_n12702_));
  NOR4_X1    g12510(.A1(new_n12657_), .A2(\asqrt[24] ), .A3(new_n12702_), .A4(new_n12180_), .ZN(new_n12703_));
  XOR2_X1    g12511(.A1(new_n12703_), .A2(new_n12156_), .Z(new_n12704_));
  NAND2_X1   g12512(.A1(new_n12704_), .A2(new_n9672_), .ZN(new_n12705_));
  INV_X1     g12513(.I(new_n12705_), .ZN(new_n12706_));
  OAI21_X1   g12514(.A1(new_n12701_), .A2(new_n10104_), .B(new_n12706_), .ZN(new_n12707_));
  NAND2_X1   g12515(.A1(new_n12707_), .A2(new_n12700_), .ZN(new_n12708_));
  OAI22_X1   g12516(.A1(new_n12701_), .A2(new_n10104_), .B1(new_n12699_), .B2(new_n12693_), .ZN(new_n12709_));
  NOR4_X1    g12517(.A1(new_n12657_), .A2(\asqrt[25] ), .A3(new_n12160_), .A4(new_n12465_), .ZN(new_n12710_));
  XNOR2_X1   g12518(.A1(new_n12710_), .A2(new_n12164_), .ZN(new_n12711_));
  NAND2_X1   g12519(.A1(new_n12711_), .A2(new_n9212_), .ZN(new_n12712_));
  AOI21_X1   g12520(.A1(new_n12709_), .A2(\asqrt[25] ), .B(new_n12712_), .ZN(new_n12713_));
  NOR2_X1    g12521(.A1(new_n12713_), .A2(new_n12708_), .ZN(new_n12714_));
  AOI22_X1   g12522(.A1(new_n12709_), .A2(\asqrt[25] ), .B1(new_n12707_), .B2(new_n12700_), .ZN(new_n12715_));
  NOR4_X1    g12523(.A1(new_n12657_), .A2(\asqrt[26] ), .A3(new_n12168_), .A4(new_n12185_), .ZN(new_n12716_));
  XOR2_X1    g12524(.A1(new_n12716_), .A2(new_n12171_), .Z(new_n12717_));
  NAND2_X1   g12525(.A1(new_n12717_), .A2(new_n8763_), .ZN(new_n12718_));
  INV_X1     g12526(.I(new_n12718_), .ZN(new_n12719_));
  OAI21_X1   g12527(.A1(new_n12715_), .A2(new_n9212_), .B(new_n12719_), .ZN(new_n12720_));
  NAND2_X1   g12528(.A1(new_n12720_), .A2(new_n12714_), .ZN(new_n12721_));
  OAI22_X1   g12529(.A1(new_n12715_), .A2(new_n9212_), .B1(new_n12713_), .B2(new_n12708_), .ZN(new_n12722_));
  NOR4_X1    g12530(.A1(new_n12657_), .A2(\asqrt[27] ), .A3(new_n12174_), .A4(new_n12471_), .ZN(new_n12723_));
  XNOR2_X1   g12531(.A1(new_n12723_), .A2(new_n12474_), .ZN(new_n12724_));
  NAND2_X1   g12532(.A1(new_n12724_), .A2(new_n8319_), .ZN(new_n12725_));
  AOI21_X1   g12533(.A1(new_n12722_), .A2(\asqrt[27] ), .B(new_n12725_), .ZN(new_n12726_));
  NOR2_X1    g12534(.A1(new_n12726_), .A2(new_n12721_), .ZN(new_n12727_));
  AOI22_X1   g12535(.A1(new_n12722_), .A2(\asqrt[27] ), .B1(new_n12720_), .B2(new_n12714_), .ZN(new_n12728_));
  NOR4_X1    g12536(.A1(new_n12657_), .A2(\asqrt[28] ), .A3(new_n12189_), .A4(new_n12195_), .ZN(new_n12729_));
  XOR2_X1    g12537(.A1(new_n12729_), .A2(new_n12475_), .Z(new_n12730_));
  NAND2_X1   g12538(.A1(new_n12730_), .A2(new_n7931_), .ZN(new_n12731_));
  INV_X1     g12539(.I(new_n12731_), .ZN(new_n12732_));
  OAI21_X1   g12540(.A1(new_n12728_), .A2(new_n8319_), .B(new_n12732_), .ZN(new_n12733_));
  NAND2_X1   g12541(.A1(new_n12733_), .A2(new_n12727_), .ZN(new_n12734_));
  OAI22_X1   g12542(.A1(new_n12728_), .A2(new_n8319_), .B1(new_n12726_), .B2(new_n12721_), .ZN(new_n12735_));
  NAND2_X1   g12543(.A1(new_n12480_), .A2(\asqrt[29] ), .ZN(new_n12736_));
  NOR4_X1    g12544(.A1(new_n12657_), .A2(\asqrt[29] ), .A3(new_n12198_), .A4(new_n12480_), .ZN(new_n12737_));
  XOR2_X1    g12545(.A1(new_n12737_), .A2(new_n12736_), .Z(new_n12738_));
  NAND2_X1   g12546(.A1(new_n12738_), .A2(new_n7517_), .ZN(new_n12739_));
  AOI21_X1   g12547(.A1(new_n12735_), .A2(\asqrt[29] ), .B(new_n12739_), .ZN(new_n12740_));
  NOR2_X1    g12548(.A1(new_n12740_), .A2(new_n12734_), .ZN(new_n12741_));
  AOI22_X1   g12549(.A1(new_n12735_), .A2(\asqrt[29] ), .B1(new_n12733_), .B2(new_n12727_), .ZN(new_n12742_));
  NOR4_X1    g12550(.A1(new_n12657_), .A2(\asqrt[30] ), .A3(new_n12205_), .A4(new_n12210_), .ZN(new_n12743_));
  AOI21_X1   g12551(.A1(new_n12736_), .A2(new_n12478_), .B(new_n7517_), .ZN(new_n12744_));
  NOR2_X1    g12552(.A1(new_n12743_), .A2(new_n12744_), .ZN(new_n12745_));
  NAND2_X1   g12553(.A1(new_n12745_), .A2(new_n7110_), .ZN(new_n12746_));
  INV_X1     g12554(.I(new_n12746_), .ZN(new_n12747_));
  OAI21_X1   g12555(.A1(new_n12742_), .A2(new_n7517_), .B(new_n12747_), .ZN(new_n12748_));
  NAND2_X1   g12556(.A1(new_n12748_), .A2(new_n12741_), .ZN(new_n12749_));
  OAI22_X1   g12557(.A1(new_n12742_), .A2(new_n7517_), .B1(new_n12740_), .B2(new_n12734_), .ZN(new_n12750_));
  NAND2_X1   g12558(.A1(new_n12487_), .A2(\asqrt[31] ), .ZN(new_n12751_));
  NOR4_X1    g12559(.A1(new_n12657_), .A2(\asqrt[31] ), .A3(new_n12213_), .A4(new_n12487_), .ZN(new_n12752_));
  XOR2_X1    g12560(.A1(new_n12752_), .A2(new_n12751_), .Z(new_n12753_));
  NAND2_X1   g12561(.A1(new_n12753_), .A2(new_n6708_), .ZN(new_n12754_));
  AOI21_X1   g12562(.A1(new_n12750_), .A2(\asqrt[31] ), .B(new_n12754_), .ZN(new_n12755_));
  NOR2_X1    g12563(.A1(new_n12755_), .A2(new_n12749_), .ZN(new_n12756_));
  AOI22_X1   g12564(.A1(new_n12750_), .A2(\asqrt[31] ), .B1(new_n12748_), .B2(new_n12741_), .ZN(new_n12757_));
  NOR4_X1    g12565(.A1(new_n12657_), .A2(\asqrt[32] ), .A3(new_n12220_), .A4(new_n12225_), .ZN(new_n12758_));
  AOI21_X1   g12566(.A1(new_n12751_), .A2(new_n12486_), .B(new_n6708_), .ZN(new_n12759_));
  NOR2_X1    g12567(.A1(new_n12758_), .A2(new_n12759_), .ZN(new_n12760_));
  NAND2_X1   g12568(.A1(new_n12760_), .A2(new_n6365_), .ZN(new_n12761_));
  INV_X1     g12569(.I(new_n12761_), .ZN(new_n12762_));
  OAI21_X1   g12570(.A1(new_n12757_), .A2(new_n6708_), .B(new_n12762_), .ZN(new_n12763_));
  NAND2_X1   g12571(.A1(new_n12763_), .A2(new_n12756_), .ZN(new_n12764_));
  OAI22_X1   g12572(.A1(new_n12757_), .A2(new_n6708_), .B1(new_n12755_), .B2(new_n12749_), .ZN(new_n12765_));
  NAND2_X1   g12573(.A1(new_n12494_), .A2(\asqrt[33] ), .ZN(new_n12766_));
  NOR4_X1    g12574(.A1(new_n12657_), .A2(\asqrt[33] ), .A3(new_n12228_), .A4(new_n12494_), .ZN(new_n12767_));
  XOR2_X1    g12575(.A1(new_n12767_), .A2(new_n12766_), .Z(new_n12768_));
  NAND2_X1   g12576(.A1(new_n12768_), .A2(new_n5991_), .ZN(new_n12769_));
  AOI21_X1   g12577(.A1(new_n12765_), .A2(\asqrt[33] ), .B(new_n12769_), .ZN(new_n12770_));
  NOR2_X1    g12578(.A1(new_n12770_), .A2(new_n12764_), .ZN(new_n12771_));
  AOI22_X1   g12579(.A1(new_n12765_), .A2(\asqrt[33] ), .B1(new_n12763_), .B2(new_n12756_), .ZN(new_n12772_));
  NOR4_X1    g12580(.A1(new_n12657_), .A2(\asqrt[34] ), .A3(new_n12235_), .A4(new_n12240_), .ZN(new_n12773_));
  AOI21_X1   g12581(.A1(new_n12766_), .A2(new_n12493_), .B(new_n5991_), .ZN(new_n12774_));
  NOR2_X1    g12582(.A1(new_n12773_), .A2(new_n12774_), .ZN(new_n12775_));
  NAND2_X1   g12583(.A1(new_n12775_), .A2(new_n5626_), .ZN(new_n12776_));
  INV_X1     g12584(.I(new_n12776_), .ZN(new_n12777_));
  OAI21_X1   g12585(.A1(new_n12772_), .A2(new_n5991_), .B(new_n12777_), .ZN(new_n12778_));
  NAND2_X1   g12586(.A1(new_n12778_), .A2(new_n12771_), .ZN(new_n12779_));
  OAI22_X1   g12587(.A1(new_n12772_), .A2(new_n5991_), .B1(new_n12770_), .B2(new_n12764_), .ZN(new_n12780_));
  NAND2_X1   g12588(.A1(new_n12501_), .A2(\asqrt[35] ), .ZN(new_n12781_));
  NOR4_X1    g12589(.A1(new_n12657_), .A2(\asqrt[35] ), .A3(new_n12243_), .A4(new_n12501_), .ZN(new_n12782_));
  XOR2_X1    g12590(.A1(new_n12782_), .A2(new_n12781_), .Z(new_n12783_));
  NAND2_X1   g12591(.A1(new_n12783_), .A2(new_n5273_), .ZN(new_n12784_));
  AOI21_X1   g12592(.A1(new_n12780_), .A2(\asqrt[35] ), .B(new_n12784_), .ZN(new_n12785_));
  NOR2_X1    g12593(.A1(new_n12785_), .A2(new_n12779_), .ZN(new_n12786_));
  AOI22_X1   g12594(.A1(new_n12780_), .A2(\asqrt[35] ), .B1(new_n12778_), .B2(new_n12771_), .ZN(new_n12787_));
  NOR4_X1    g12595(.A1(new_n12657_), .A2(\asqrt[36] ), .A3(new_n12250_), .A4(new_n12255_), .ZN(new_n12788_));
  AOI21_X1   g12596(.A1(new_n12781_), .A2(new_n12500_), .B(new_n5273_), .ZN(new_n12789_));
  NOR2_X1    g12597(.A1(new_n12788_), .A2(new_n12789_), .ZN(new_n12790_));
  NAND2_X1   g12598(.A1(new_n12790_), .A2(new_n4973_), .ZN(new_n12791_));
  INV_X1     g12599(.I(new_n12791_), .ZN(new_n12792_));
  OAI21_X1   g12600(.A1(new_n12787_), .A2(new_n5273_), .B(new_n12792_), .ZN(new_n12793_));
  NAND2_X1   g12601(.A1(new_n12793_), .A2(new_n12786_), .ZN(new_n12794_));
  OAI22_X1   g12602(.A1(new_n12787_), .A2(new_n5273_), .B1(new_n12785_), .B2(new_n12779_), .ZN(new_n12795_));
  NAND2_X1   g12603(.A1(new_n12508_), .A2(\asqrt[37] ), .ZN(new_n12796_));
  NOR4_X1    g12604(.A1(new_n12657_), .A2(\asqrt[37] ), .A3(new_n12258_), .A4(new_n12508_), .ZN(new_n12797_));
  XOR2_X1    g12605(.A1(new_n12797_), .A2(new_n12796_), .Z(new_n12798_));
  NAND2_X1   g12606(.A1(new_n12798_), .A2(new_n4645_), .ZN(new_n12799_));
  AOI21_X1   g12607(.A1(new_n12795_), .A2(\asqrt[37] ), .B(new_n12799_), .ZN(new_n12800_));
  NOR2_X1    g12608(.A1(new_n12800_), .A2(new_n12794_), .ZN(new_n12801_));
  AOI22_X1   g12609(.A1(new_n12795_), .A2(\asqrt[37] ), .B1(new_n12793_), .B2(new_n12786_), .ZN(new_n12802_));
  NOR4_X1    g12610(.A1(new_n12657_), .A2(\asqrt[38] ), .A3(new_n12265_), .A4(new_n12270_), .ZN(new_n12803_));
  AOI21_X1   g12611(.A1(new_n12796_), .A2(new_n12507_), .B(new_n4645_), .ZN(new_n12804_));
  NOR2_X1    g12612(.A1(new_n12803_), .A2(new_n12804_), .ZN(new_n12805_));
  NAND2_X1   g12613(.A1(new_n12805_), .A2(new_n4330_), .ZN(new_n12806_));
  INV_X1     g12614(.I(new_n12806_), .ZN(new_n12807_));
  OAI21_X1   g12615(.A1(new_n12802_), .A2(new_n4645_), .B(new_n12807_), .ZN(new_n12808_));
  NAND2_X1   g12616(.A1(new_n12808_), .A2(new_n12801_), .ZN(new_n12809_));
  OAI22_X1   g12617(.A1(new_n12802_), .A2(new_n4645_), .B1(new_n12800_), .B2(new_n12794_), .ZN(new_n12810_));
  NAND2_X1   g12618(.A1(new_n12515_), .A2(\asqrt[39] ), .ZN(new_n12811_));
  NOR4_X1    g12619(.A1(new_n12657_), .A2(\asqrt[39] ), .A3(new_n12273_), .A4(new_n12515_), .ZN(new_n12812_));
  XOR2_X1    g12620(.A1(new_n12812_), .A2(new_n12811_), .Z(new_n12813_));
  NAND2_X1   g12621(.A1(new_n12813_), .A2(new_n4018_), .ZN(new_n12814_));
  AOI21_X1   g12622(.A1(new_n12810_), .A2(\asqrt[39] ), .B(new_n12814_), .ZN(new_n12815_));
  NOR2_X1    g12623(.A1(new_n12815_), .A2(new_n12809_), .ZN(new_n12816_));
  AOI22_X1   g12624(.A1(new_n12810_), .A2(\asqrt[39] ), .B1(new_n12808_), .B2(new_n12801_), .ZN(new_n12817_));
  NAND2_X1   g12625(.A1(new_n12285_), .A2(\asqrt[40] ), .ZN(new_n12818_));
  NOR4_X1    g12626(.A1(new_n12657_), .A2(\asqrt[40] ), .A3(new_n12280_), .A4(new_n12285_), .ZN(new_n12819_));
  XOR2_X1    g12627(.A1(new_n12819_), .A2(new_n12818_), .Z(new_n12820_));
  NAND2_X1   g12628(.A1(new_n12820_), .A2(new_n3760_), .ZN(new_n12821_));
  INV_X1     g12629(.I(new_n12821_), .ZN(new_n12822_));
  OAI21_X1   g12630(.A1(new_n12817_), .A2(new_n4018_), .B(new_n12822_), .ZN(new_n12823_));
  NAND2_X1   g12631(.A1(new_n12823_), .A2(new_n12816_), .ZN(new_n12824_));
  OAI22_X1   g12632(.A1(new_n12817_), .A2(new_n4018_), .B1(new_n12815_), .B2(new_n12809_), .ZN(new_n12825_));
  NOR4_X1    g12633(.A1(new_n12657_), .A2(\asqrt[41] ), .A3(new_n12288_), .A4(new_n12522_), .ZN(new_n12826_));
  AOI21_X1   g12634(.A1(new_n12818_), .A2(new_n12284_), .B(new_n3760_), .ZN(new_n12827_));
  NOR2_X1    g12635(.A1(new_n12826_), .A2(new_n12827_), .ZN(new_n12828_));
  NAND2_X1   g12636(.A1(new_n12828_), .A2(new_n3481_), .ZN(new_n12829_));
  AOI21_X1   g12637(.A1(new_n12825_), .A2(\asqrt[41] ), .B(new_n12829_), .ZN(new_n12830_));
  NOR2_X1    g12638(.A1(new_n12830_), .A2(new_n12824_), .ZN(new_n12831_));
  AOI22_X1   g12639(.A1(new_n12825_), .A2(\asqrt[41] ), .B1(new_n12823_), .B2(new_n12816_), .ZN(new_n12832_));
  NAND2_X1   g12640(.A1(new_n12300_), .A2(\asqrt[42] ), .ZN(new_n12833_));
  NOR4_X1    g12641(.A1(new_n12657_), .A2(\asqrt[42] ), .A3(new_n12295_), .A4(new_n12300_), .ZN(new_n12834_));
  XOR2_X1    g12642(.A1(new_n12834_), .A2(new_n12833_), .Z(new_n12835_));
  NAND2_X1   g12643(.A1(new_n12835_), .A2(new_n3208_), .ZN(new_n12836_));
  INV_X1     g12644(.I(new_n12836_), .ZN(new_n12837_));
  OAI21_X1   g12645(.A1(new_n12832_), .A2(new_n3481_), .B(new_n12837_), .ZN(new_n12838_));
  NAND2_X1   g12646(.A1(new_n12838_), .A2(new_n12831_), .ZN(new_n12839_));
  OAI22_X1   g12647(.A1(new_n12832_), .A2(new_n3481_), .B1(new_n12830_), .B2(new_n12824_), .ZN(new_n12840_));
  NOR4_X1    g12648(.A1(new_n12657_), .A2(\asqrt[43] ), .A3(new_n12303_), .A4(new_n12529_), .ZN(new_n12841_));
  AOI21_X1   g12649(.A1(new_n12833_), .A2(new_n12299_), .B(new_n3208_), .ZN(new_n12842_));
  NOR2_X1    g12650(.A1(new_n12841_), .A2(new_n12842_), .ZN(new_n12843_));
  NAND2_X1   g12651(.A1(new_n12843_), .A2(new_n2941_), .ZN(new_n12844_));
  AOI21_X1   g12652(.A1(new_n12840_), .A2(\asqrt[43] ), .B(new_n12844_), .ZN(new_n12845_));
  NOR2_X1    g12653(.A1(new_n12845_), .A2(new_n12839_), .ZN(new_n12846_));
  AOI22_X1   g12654(.A1(new_n12840_), .A2(\asqrt[43] ), .B1(new_n12838_), .B2(new_n12831_), .ZN(new_n12847_));
  NAND2_X1   g12655(.A1(new_n12315_), .A2(\asqrt[44] ), .ZN(new_n12848_));
  NOR4_X1    g12656(.A1(new_n12657_), .A2(\asqrt[44] ), .A3(new_n12310_), .A4(new_n12315_), .ZN(new_n12849_));
  XOR2_X1    g12657(.A1(new_n12849_), .A2(new_n12848_), .Z(new_n12850_));
  NAND2_X1   g12658(.A1(new_n12850_), .A2(new_n2728_), .ZN(new_n12851_));
  INV_X1     g12659(.I(new_n12851_), .ZN(new_n12852_));
  OAI21_X1   g12660(.A1(new_n12847_), .A2(new_n2941_), .B(new_n12852_), .ZN(new_n12853_));
  NAND2_X1   g12661(.A1(new_n12853_), .A2(new_n12846_), .ZN(new_n12854_));
  OAI22_X1   g12662(.A1(new_n12847_), .A2(new_n2941_), .B1(new_n12845_), .B2(new_n12839_), .ZN(new_n12855_));
  NAND2_X1   g12663(.A1(new_n12536_), .A2(\asqrt[45] ), .ZN(new_n12856_));
  NOR4_X1    g12664(.A1(new_n12657_), .A2(\asqrt[45] ), .A3(new_n12318_), .A4(new_n12536_), .ZN(new_n12857_));
  XOR2_X1    g12665(.A1(new_n12857_), .A2(new_n12856_), .Z(new_n12858_));
  NAND2_X1   g12666(.A1(new_n12858_), .A2(new_n2488_), .ZN(new_n12859_));
  AOI21_X1   g12667(.A1(new_n12855_), .A2(\asqrt[45] ), .B(new_n12859_), .ZN(new_n12860_));
  NOR2_X1    g12668(.A1(new_n12860_), .A2(new_n12854_), .ZN(new_n12861_));
  AOI22_X1   g12669(.A1(new_n12855_), .A2(\asqrt[45] ), .B1(new_n12853_), .B2(new_n12846_), .ZN(new_n12862_));
  NOR4_X1    g12670(.A1(new_n12657_), .A2(\asqrt[46] ), .A3(new_n12325_), .A4(new_n12330_), .ZN(new_n12863_));
  AOI21_X1   g12671(.A1(new_n12856_), .A2(new_n12535_), .B(new_n2488_), .ZN(new_n12864_));
  NOR2_X1    g12672(.A1(new_n12863_), .A2(new_n12864_), .ZN(new_n12865_));
  NAND2_X1   g12673(.A1(new_n12865_), .A2(new_n2253_), .ZN(new_n12866_));
  INV_X1     g12674(.I(new_n12866_), .ZN(new_n12867_));
  OAI21_X1   g12675(.A1(new_n12862_), .A2(new_n2488_), .B(new_n12867_), .ZN(new_n12868_));
  NAND2_X1   g12676(.A1(new_n12868_), .A2(new_n12861_), .ZN(new_n12869_));
  OAI22_X1   g12677(.A1(new_n12862_), .A2(new_n2488_), .B1(new_n12860_), .B2(new_n12854_), .ZN(new_n12870_));
  NAND2_X1   g12678(.A1(new_n12543_), .A2(\asqrt[47] ), .ZN(new_n12871_));
  NOR4_X1    g12679(.A1(new_n12657_), .A2(\asqrt[47] ), .A3(new_n12333_), .A4(new_n12543_), .ZN(new_n12872_));
  XOR2_X1    g12680(.A1(new_n12872_), .A2(new_n12871_), .Z(new_n12873_));
  NAND2_X1   g12681(.A1(new_n12873_), .A2(new_n2046_), .ZN(new_n12874_));
  AOI21_X1   g12682(.A1(new_n12870_), .A2(\asqrt[47] ), .B(new_n12874_), .ZN(new_n12875_));
  NOR2_X1    g12683(.A1(new_n12875_), .A2(new_n12869_), .ZN(new_n12876_));
  AOI22_X1   g12684(.A1(new_n12870_), .A2(\asqrt[47] ), .B1(new_n12868_), .B2(new_n12861_), .ZN(new_n12877_));
  NOR4_X1    g12685(.A1(new_n12657_), .A2(\asqrt[48] ), .A3(new_n12340_), .A4(new_n12345_), .ZN(new_n12878_));
  AOI21_X1   g12686(.A1(new_n12871_), .A2(new_n12542_), .B(new_n2046_), .ZN(new_n12879_));
  NOR2_X1    g12687(.A1(new_n12878_), .A2(new_n12879_), .ZN(new_n12880_));
  NAND2_X1   g12688(.A1(new_n12880_), .A2(new_n1854_), .ZN(new_n12881_));
  INV_X1     g12689(.I(new_n12881_), .ZN(new_n12882_));
  OAI21_X1   g12690(.A1(new_n12877_), .A2(new_n2046_), .B(new_n12882_), .ZN(new_n12883_));
  NAND2_X1   g12691(.A1(new_n12883_), .A2(new_n12876_), .ZN(new_n12884_));
  OAI22_X1   g12692(.A1(new_n12877_), .A2(new_n2046_), .B1(new_n12875_), .B2(new_n12869_), .ZN(new_n12885_));
  NAND2_X1   g12693(.A1(new_n12550_), .A2(\asqrt[49] ), .ZN(new_n12886_));
  NOR4_X1    g12694(.A1(new_n12657_), .A2(\asqrt[49] ), .A3(new_n12348_), .A4(new_n12550_), .ZN(new_n12887_));
  XOR2_X1    g12695(.A1(new_n12887_), .A2(new_n12886_), .Z(new_n12888_));
  NAND2_X1   g12696(.A1(new_n12888_), .A2(new_n1595_), .ZN(new_n12889_));
  AOI21_X1   g12697(.A1(new_n12885_), .A2(\asqrt[49] ), .B(new_n12889_), .ZN(new_n12890_));
  NOR2_X1    g12698(.A1(new_n12890_), .A2(new_n12884_), .ZN(new_n12891_));
  AOI22_X1   g12699(.A1(new_n12885_), .A2(\asqrt[49] ), .B1(new_n12883_), .B2(new_n12876_), .ZN(new_n12892_));
  NOR4_X1    g12700(.A1(new_n12657_), .A2(\asqrt[50] ), .A3(new_n12355_), .A4(new_n12360_), .ZN(new_n12893_));
  AOI21_X1   g12701(.A1(new_n12886_), .A2(new_n12549_), .B(new_n1595_), .ZN(new_n12894_));
  NOR2_X1    g12702(.A1(new_n12893_), .A2(new_n12894_), .ZN(new_n12895_));
  NAND2_X1   g12703(.A1(new_n12895_), .A2(new_n1436_), .ZN(new_n12896_));
  INV_X1     g12704(.I(new_n12896_), .ZN(new_n12897_));
  OAI21_X1   g12705(.A1(new_n12892_), .A2(new_n1595_), .B(new_n12897_), .ZN(new_n12898_));
  NAND2_X1   g12706(.A1(new_n12898_), .A2(new_n12891_), .ZN(new_n12899_));
  OAI22_X1   g12707(.A1(new_n12892_), .A2(new_n1595_), .B1(new_n12890_), .B2(new_n12884_), .ZN(new_n12900_));
  NAND2_X1   g12708(.A1(new_n12557_), .A2(\asqrt[51] ), .ZN(new_n12901_));
  NOR4_X1    g12709(.A1(new_n12657_), .A2(\asqrt[51] ), .A3(new_n12363_), .A4(new_n12557_), .ZN(new_n12902_));
  XOR2_X1    g12710(.A1(new_n12902_), .A2(new_n12901_), .Z(new_n12903_));
  NAND2_X1   g12711(.A1(new_n12903_), .A2(new_n1260_), .ZN(new_n12904_));
  AOI21_X1   g12712(.A1(new_n12900_), .A2(\asqrt[51] ), .B(new_n12904_), .ZN(new_n12905_));
  NOR2_X1    g12713(.A1(new_n12905_), .A2(new_n12899_), .ZN(new_n12906_));
  AOI22_X1   g12714(.A1(new_n12900_), .A2(\asqrt[51] ), .B1(new_n12898_), .B2(new_n12891_), .ZN(new_n12907_));
  NAND2_X1   g12715(.A1(new_n12375_), .A2(\asqrt[52] ), .ZN(new_n12908_));
  NOR4_X1    g12716(.A1(new_n12657_), .A2(\asqrt[52] ), .A3(new_n12370_), .A4(new_n12375_), .ZN(new_n12909_));
  XOR2_X1    g12717(.A1(new_n12909_), .A2(new_n12908_), .Z(new_n12910_));
  NAND2_X1   g12718(.A1(new_n12910_), .A2(new_n1096_), .ZN(new_n12911_));
  INV_X1     g12719(.I(new_n12911_), .ZN(new_n12912_));
  OAI21_X1   g12720(.A1(new_n12907_), .A2(new_n1260_), .B(new_n12912_), .ZN(new_n12913_));
  NAND2_X1   g12721(.A1(new_n12913_), .A2(new_n12906_), .ZN(new_n12914_));
  OAI22_X1   g12722(.A1(new_n12907_), .A2(new_n1260_), .B1(new_n12905_), .B2(new_n12899_), .ZN(new_n12915_));
  NOR4_X1    g12723(.A1(new_n12657_), .A2(\asqrt[53] ), .A3(new_n12378_), .A4(new_n12564_), .ZN(new_n12916_));
  XOR2_X1    g12724(.A1(new_n12916_), .A2(new_n12578_), .Z(new_n12917_));
  NAND2_X1   g12725(.A1(new_n12917_), .A2(new_n970_), .ZN(new_n12918_));
  AOI21_X1   g12726(.A1(new_n12915_), .A2(\asqrt[53] ), .B(new_n12918_), .ZN(new_n12919_));
  NOR2_X1    g12727(.A1(new_n12919_), .A2(new_n12914_), .ZN(new_n12920_));
  AOI22_X1   g12728(.A1(new_n12915_), .A2(\asqrt[53] ), .B1(new_n12913_), .B2(new_n12906_), .ZN(new_n12921_));
  NOR4_X1    g12729(.A1(new_n12657_), .A2(\asqrt[54] ), .A3(new_n12385_), .A4(new_n12390_), .ZN(new_n12922_));
  XOR2_X1    g12730(.A1(new_n12922_), .A2(new_n12428_), .Z(new_n12923_));
  NAND2_X1   g12731(.A1(new_n12923_), .A2(new_n825_), .ZN(new_n12924_));
  INV_X1     g12732(.I(new_n12924_), .ZN(new_n12925_));
  OAI21_X1   g12733(.A1(new_n12921_), .A2(new_n970_), .B(new_n12925_), .ZN(new_n12926_));
  NAND2_X1   g12734(.A1(new_n12926_), .A2(new_n12920_), .ZN(new_n12927_));
  OAI22_X1   g12735(.A1(new_n12921_), .A2(new_n970_), .B1(new_n12919_), .B2(new_n12914_), .ZN(new_n12928_));
  NOR4_X1    g12736(.A1(new_n12657_), .A2(\asqrt[55] ), .A3(new_n12392_), .A4(new_n12571_), .ZN(new_n12929_));
  XOR2_X1    g12737(.A1(new_n12929_), .A2(new_n12580_), .Z(new_n12930_));
  NAND2_X1   g12738(.A1(new_n12930_), .A2(new_n724_), .ZN(new_n12931_));
  AOI21_X1   g12739(.A1(new_n12928_), .A2(\asqrt[55] ), .B(new_n12931_), .ZN(new_n12932_));
  NOR2_X1    g12740(.A1(new_n12932_), .A2(new_n12927_), .ZN(new_n12933_));
  AOI22_X1   g12741(.A1(new_n12928_), .A2(\asqrt[55] ), .B1(new_n12926_), .B2(new_n12920_), .ZN(new_n12934_));
  NOR4_X1    g12742(.A1(new_n12657_), .A2(\asqrt[56] ), .A3(new_n12398_), .A4(new_n12403_), .ZN(new_n12935_));
  XOR2_X1    g12743(.A1(new_n12935_), .A2(new_n12430_), .Z(new_n12936_));
  NAND2_X1   g12744(.A1(new_n12936_), .A2(new_n587_), .ZN(new_n12937_));
  INV_X1     g12745(.I(new_n12937_), .ZN(new_n12938_));
  OAI21_X1   g12746(.A1(new_n12934_), .A2(new_n724_), .B(new_n12938_), .ZN(new_n12939_));
  NAND2_X1   g12747(.A1(new_n12939_), .A2(new_n12933_), .ZN(new_n12940_));
  OAI22_X1   g12748(.A1(new_n12934_), .A2(new_n724_), .B1(new_n12932_), .B2(new_n12927_), .ZN(new_n12941_));
  NOR4_X1    g12749(.A1(new_n12657_), .A2(\asqrt[57] ), .A3(new_n12405_), .A4(new_n12584_), .ZN(new_n12942_));
  XOR2_X1    g12750(.A1(new_n12942_), .A2(new_n12582_), .Z(new_n12943_));
  NAND2_X1   g12751(.A1(new_n12943_), .A2(new_n504_), .ZN(new_n12944_));
  AOI21_X1   g12752(.A1(new_n12941_), .A2(\asqrt[57] ), .B(new_n12944_), .ZN(new_n12945_));
  NOR2_X1    g12753(.A1(new_n12945_), .A2(new_n12940_), .ZN(new_n12946_));
  AOI22_X1   g12754(.A1(new_n12941_), .A2(\asqrt[57] ), .B1(new_n12939_), .B2(new_n12933_), .ZN(new_n12947_));
  NOR4_X1    g12755(.A1(new_n12657_), .A2(\asqrt[58] ), .A3(new_n12411_), .A4(new_n12416_), .ZN(new_n12948_));
  XOR2_X1    g12756(.A1(new_n12948_), .A2(new_n12432_), .Z(new_n12949_));
  NAND2_X1   g12757(.A1(new_n12949_), .A2(new_n376_), .ZN(new_n12950_));
  INV_X1     g12758(.I(new_n12950_), .ZN(new_n12951_));
  OAI21_X1   g12759(.A1(new_n12947_), .A2(new_n504_), .B(new_n12951_), .ZN(new_n12952_));
  NAND2_X1   g12760(.A1(new_n12952_), .A2(new_n12946_), .ZN(new_n12953_));
  OAI22_X1   g12761(.A1(new_n12947_), .A2(new_n504_), .B1(new_n12945_), .B2(new_n12940_), .ZN(new_n12954_));
  NOR4_X1    g12762(.A1(new_n12657_), .A2(\asqrt[59] ), .A3(new_n12418_), .A4(new_n12592_), .ZN(new_n12955_));
  XOR2_X1    g12763(.A1(new_n12955_), .A2(new_n12590_), .Z(new_n12956_));
  NAND2_X1   g12764(.A1(new_n12956_), .A2(new_n275_), .ZN(new_n12957_));
  AOI21_X1   g12765(.A1(new_n12954_), .A2(\asqrt[59] ), .B(new_n12957_), .ZN(new_n12958_));
  NOR2_X1    g12766(.A1(new_n12958_), .A2(new_n12953_), .ZN(new_n12959_));
  AOI22_X1   g12767(.A1(new_n12954_), .A2(\asqrt[59] ), .B1(new_n12952_), .B2(new_n12946_), .ZN(new_n12960_));
  OAI22_X1   g12768(.A1(new_n12960_), .A2(new_n275_), .B1(new_n12958_), .B2(new_n12953_), .ZN(new_n12961_));
  NOR4_X1    g12769(.A1(new_n12657_), .A2(\asqrt[60] ), .A3(new_n12424_), .A4(new_n12613_), .ZN(new_n12962_));
  XOR2_X1    g12770(.A1(new_n12962_), .A2(new_n12434_), .Z(new_n12963_));
  NAND2_X1   g12771(.A1(new_n12963_), .A2(new_n229_), .ZN(new_n12964_));
  INV_X1     g12772(.I(new_n12964_), .ZN(new_n12965_));
  OAI21_X1   g12773(.A1(new_n12960_), .A2(new_n275_), .B(new_n12965_), .ZN(new_n12966_));
  AOI22_X1   g12774(.A1(new_n12961_), .A2(\asqrt[61] ), .B1(new_n12966_), .B2(new_n12959_), .ZN(new_n12967_));
  NOR2_X1    g12775(.A1(new_n12967_), .A2(new_n196_), .ZN(new_n12968_));
  INV_X1     g12776(.I(new_n12634_), .ZN(new_n12969_));
  AOI21_X1   g12777(.A1(new_n12648_), .A2(new_n12969_), .B(new_n12636_), .ZN(new_n12970_));
  NOR3_X1    g12778(.A1(new_n12633_), .A2(new_n12626_), .A3(new_n12631_), .ZN(new_n12971_));
  NOR2_X1    g12779(.A1(new_n12971_), .A2(new_n12970_), .ZN(new_n12972_));
  NOR3_X1    g12780(.A1(new_n12671_), .A2(new_n11575_), .A3(\asqrt[19] ), .ZN(new_n12973_));
  AOI21_X1   g12781(.A1(new_n12665_), .A2(new_n11574_), .B(new_n12657_), .ZN(new_n12974_));
  NOR4_X1    g12782(.A1(new_n12974_), .A2(new_n12973_), .A3(\asqrt[21] ), .A4(new_n12655_), .ZN(new_n12975_));
  NOR2_X1    g12783(.A1(new_n12975_), .A2(new_n12972_), .ZN(new_n12976_));
  NOR3_X1    g12784(.A1(new_n12971_), .A2(new_n12970_), .A3(new_n12655_), .ZN(new_n12977_));
  NOR3_X1    g12785(.A1(new_n12657_), .A2(new_n12099_), .A3(new_n12682_), .ZN(new_n12978_));
  AOI21_X1   g12786(.A1(\asqrt[19] ), .A2(new_n12680_), .B(new_n12100_), .ZN(new_n12979_));
  NOR3_X1    g12787(.A1(new_n12979_), .A2(new_n12978_), .A3(\asqrt[22] ), .ZN(new_n12980_));
  OAI21_X1   g12788(.A1(new_n12977_), .A2(new_n11631_), .B(new_n12980_), .ZN(new_n12981_));
  NAND2_X1   g12789(.A1(new_n12976_), .A2(new_n12981_), .ZN(new_n12982_));
  OAI22_X1   g12790(.A1(new_n12975_), .A2(new_n12972_), .B1(new_n11631_), .B2(new_n12977_), .ZN(new_n12983_));
  INV_X1     g12791(.I(new_n12691_), .ZN(new_n12984_));
  AOI21_X1   g12792(.A1(new_n12983_), .A2(\asqrt[22] ), .B(new_n12984_), .ZN(new_n12985_));
  NOR2_X1    g12793(.A1(new_n12985_), .A2(new_n12982_), .ZN(new_n12986_));
  AOI22_X1   g12794(.A1(new_n12983_), .A2(\asqrt[22] ), .B1(new_n12976_), .B2(new_n12981_), .ZN(new_n12987_));
  INV_X1     g12795(.I(new_n12698_), .ZN(new_n12988_));
  OAI21_X1   g12796(.A1(new_n12987_), .A2(new_n10614_), .B(new_n12988_), .ZN(new_n12989_));
  NAND2_X1   g12797(.A1(new_n12989_), .A2(new_n12986_), .ZN(new_n12990_));
  OAI22_X1   g12798(.A1(new_n12987_), .A2(new_n10614_), .B1(new_n12985_), .B2(new_n12982_), .ZN(new_n12991_));
  AOI21_X1   g12799(.A1(new_n12991_), .A2(\asqrt[24] ), .B(new_n12705_), .ZN(new_n12992_));
  NOR2_X1    g12800(.A1(new_n12992_), .A2(new_n12990_), .ZN(new_n12993_));
  AOI22_X1   g12801(.A1(new_n12991_), .A2(\asqrt[24] ), .B1(new_n12989_), .B2(new_n12986_), .ZN(new_n12994_));
  INV_X1     g12802(.I(new_n12712_), .ZN(new_n12995_));
  OAI21_X1   g12803(.A1(new_n12994_), .A2(new_n9672_), .B(new_n12995_), .ZN(new_n12996_));
  NAND2_X1   g12804(.A1(new_n12996_), .A2(new_n12993_), .ZN(new_n12997_));
  OAI22_X1   g12805(.A1(new_n12994_), .A2(new_n9672_), .B1(new_n12992_), .B2(new_n12990_), .ZN(new_n12998_));
  AOI21_X1   g12806(.A1(new_n12998_), .A2(\asqrt[26] ), .B(new_n12718_), .ZN(new_n12999_));
  NOR2_X1    g12807(.A1(new_n12999_), .A2(new_n12997_), .ZN(new_n13000_));
  AOI22_X1   g12808(.A1(new_n12998_), .A2(\asqrt[26] ), .B1(new_n12996_), .B2(new_n12993_), .ZN(new_n13001_));
  INV_X1     g12809(.I(new_n12725_), .ZN(new_n13002_));
  OAI21_X1   g12810(.A1(new_n13001_), .A2(new_n8763_), .B(new_n13002_), .ZN(new_n13003_));
  NAND2_X1   g12811(.A1(new_n13003_), .A2(new_n13000_), .ZN(new_n13004_));
  OAI22_X1   g12812(.A1(new_n13001_), .A2(new_n8763_), .B1(new_n12999_), .B2(new_n12997_), .ZN(new_n13005_));
  AOI21_X1   g12813(.A1(new_n13005_), .A2(\asqrt[28] ), .B(new_n12731_), .ZN(new_n13006_));
  NOR2_X1    g12814(.A1(new_n13006_), .A2(new_n13004_), .ZN(new_n13007_));
  AOI22_X1   g12815(.A1(new_n13005_), .A2(\asqrt[28] ), .B1(new_n13003_), .B2(new_n13000_), .ZN(new_n13008_));
  INV_X1     g12816(.I(new_n12739_), .ZN(new_n13009_));
  OAI21_X1   g12817(.A1(new_n13008_), .A2(new_n7931_), .B(new_n13009_), .ZN(new_n13010_));
  NAND2_X1   g12818(.A1(new_n13010_), .A2(new_n13007_), .ZN(new_n13011_));
  OAI22_X1   g12819(.A1(new_n13008_), .A2(new_n7931_), .B1(new_n13006_), .B2(new_n13004_), .ZN(new_n13012_));
  AOI21_X1   g12820(.A1(new_n13012_), .A2(\asqrt[30] ), .B(new_n12746_), .ZN(new_n13013_));
  NOR2_X1    g12821(.A1(new_n13013_), .A2(new_n13011_), .ZN(new_n13014_));
  AOI22_X1   g12822(.A1(new_n13012_), .A2(\asqrt[30] ), .B1(new_n13010_), .B2(new_n13007_), .ZN(new_n13015_));
  INV_X1     g12823(.I(new_n12754_), .ZN(new_n13016_));
  OAI21_X1   g12824(.A1(new_n13015_), .A2(new_n7110_), .B(new_n13016_), .ZN(new_n13017_));
  NAND2_X1   g12825(.A1(new_n13017_), .A2(new_n13014_), .ZN(new_n13018_));
  OAI22_X1   g12826(.A1(new_n13015_), .A2(new_n7110_), .B1(new_n13013_), .B2(new_n13011_), .ZN(new_n13019_));
  AOI21_X1   g12827(.A1(new_n13019_), .A2(\asqrt[32] ), .B(new_n12761_), .ZN(new_n13020_));
  NOR2_X1    g12828(.A1(new_n13020_), .A2(new_n13018_), .ZN(new_n13021_));
  AOI22_X1   g12829(.A1(new_n13019_), .A2(\asqrt[32] ), .B1(new_n13017_), .B2(new_n13014_), .ZN(new_n13022_));
  INV_X1     g12830(.I(new_n12769_), .ZN(new_n13023_));
  OAI21_X1   g12831(.A1(new_n13022_), .A2(new_n6365_), .B(new_n13023_), .ZN(new_n13024_));
  NAND2_X1   g12832(.A1(new_n13024_), .A2(new_n13021_), .ZN(new_n13025_));
  OAI22_X1   g12833(.A1(new_n13022_), .A2(new_n6365_), .B1(new_n13020_), .B2(new_n13018_), .ZN(new_n13026_));
  AOI21_X1   g12834(.A1(new_n13026_), .A2(\asqrt[34] ), .B(new_n12776_), .ZN(new_n13027_));
  NOR2_X1    g12835(.A1(new_n13027_), .A2(new_n13025_), .ZN(new_n13028_));
  AOI22_X1   g12836(.A1(new_n13026_), .A2(\asqrt[34] ), .B1(new_n13024_), .B2(new_n13021_), .ZN(new_n13029_));
  INV_X1     g12837(.I(new_n12784_), .ZN(new_n13030_));
  OAI21_X1   g12838(.A1(new_n13029_), .A2(new_n5626_), .B(new_n13030_), .ZN(new_n13031_));
  NAND2_X1   g12839(.A1(new_n13031_), .A2(new_n13028_), .ZN(new_n13032_));
  OAI22_X1   g12840(.A1(new_n13029_), .A2(new_n5626_), .B1(new_n13027_), .B2(new_n13025_), .ZN(new_n13033_));
  AOI21_X1   g12841(.A1(new_n13033_), .A2(\asqrt[36] ), .B(new_n12791_), .ZN(new_n13034_));
  NOR2_X1    g12842(.A1(new_n13034_), .A2(new_n13032_), .ZN(new_n13035_));
  AOI22_X1   g12843(.A1(new_n13033_), .A2(\asqrt[36] ), .B1(new_n13031_), .B2(new_n13028_), .ZN(new_n13036_));
  INV_X1     g12844(.I(new_n12799_), .ZN(new_n13037_));
  OAI21_X1   g12845(.A1(new_n13036_), .A2(new_n4973_), .B(new_n13037_), .ZN(new_n13038_));
  NAND2_X1   g12846(.A1(new_n13038_), .A2(new_n13035_), .ZN(new_n13039_));
  OAI22_X1   g12847(.A1(new_n13036_), .A2(new_n4973_), .B1(new_n13034_), .B2(new_n13032_), .ZN(new_n13040_));
  AOI21_X1   g12848(.A1(new_n13040_), .A2(\asqrt[38] ), .B(new_n12806_), .ZN(new_n13041_));
  NOR2_X1    g12849(.A1(new_n13041_), .A2(new_n13039_), .ZN(new_n13042_));
  AOI22_X1   g12850(.A1(new_n13040_), .A2(\asqrt[38] ), .B1(new_n13038_), .B2(new_n13035_), .ZN(new_n13043_));
  INV_X1     g12851(.I(new_n12814_), .ZN(new_n13044_));
  OAI21_X1   g12852(.A1(new_n13043_), .A2(new_n4330_), .B(new_n13044_), .ZN(new_n13045_));
  NAND2_X1   g12853(.A1(new_n13045_), .A2(new_n13042_), .ZN(new_n13046_));
  OAI22_X1   g12854(.A1(new_n13043_), .A2(new_n4330_), .B1(new_n13041_), .B2(new_n13039_), .ZN(new_n13047_));
  AOI21_X1   g12855(.A1(new_n13047_), .A2(\asqrt[40] ), .B(new_n12821_), .ZN(new_n13048_));
  NOR2_X1    g12856(.A1(new_n13048_), .A2(new_n13046_), .ZN(new_n13049_));
  AOI22_X1   g12857(.A1(new_n13047_), .A2(\asqrt[40] ), .B1(new_n13045_), .B2(new_n13042_), .ZN(new_n13050_));
  INV_X1     g12858(.I(new_n12829_), .ZN(new_n13051_));
  OAI21_X1   g12859(.A1(new_n13050_), .A2(new_n3760_), .B(new_n13051_), .ZN(new_n13052_));
  NAND2_X1   g12860(.A1(new_n13052_), .A2(new_n13049_), .ZN(new_n13053_));
  OAI22_X1   g12861(.A1(new_n13050_), .A2(new_n3760_), .B1(new_n13048_), .B2(new_n13046_), .ZN(new_n13054_));
  AOI21_X1   g12862(.A1(new_n13054_), .A2(\asqrt[42] ), .B(new_n12836_), .ZN(new_n13055_));
  NOR2_X1    g12863(.A1(new_n13055_), .A2(new_n13053_), .ZN(new_n13056_));
  AOI22_X1   g12864(.A1(new_n13054_), .A2(\asqrt[42] ), .B1(new_n13052_), .B2(new_n13049_), .ZN(new_n13057_));
  INV_X1     g12865(.I(new_n12844_), .ZN(new_n13058_));
  OAI21_X1   g12866(.A1(new_n13057_), .A2(new_n3208_), .B(new_n13058_), .ZN(new_n13059_));
  NAND2_X1   g12867(.A1(new_n13059_), .A2(new_n13056_), .ZN(new_n13060_));
  OAI22_X1   g12868(.A1(new_n13057_), .A2(new_n3208_), .B1(new_n13055_), .B2(new_n13053_), .ZN(new_n13061_));
  AOI21_X1   g12869(.A1(new_n13061_), .A2(\asqrt[44] ), .B(new_n12851_), .ZN(new_n13062_));
  NOR2_X1    g12870(.A1(new_n13062_), .A2(new_n13060_), .ZN(new_n13063_));
  AOI22_X1   g12871(.A1(new_n13061_), .A2(\asqrt[44] ), .B1(new_n13059_), .B2(new_n13056_), .ZN(new_n13064_));
  INV_X1     g12872(.I(new_n12859_), .ZN(new_n13065_));
  OAI21_X1   g12873(.A1(new_n13064_), .A2(new_n2728_), .B(new_n13065_), .ZN(new_n13066_));
  NAND2_X1   g12874(.A1(new_n13066_), .A2(new_n13063_), .ZN(new_n13067_));
  OAI22_X1   g12875(.A1(new_n13064_), .A2(new_n2728_), .B1(new_n13062_), .B2(new_n13060_), .ZN(new_n13068_));
  AOI21_X1   g12876(.A1(new_n13068_), .A2(\asqrt[46] ), .B(new_n12866_), .ZN(new_n13069_));
  NOR2_X1    g12877(.A1(new_n13069_), .A2(new_n13067_), .ZN(new_n13070_));
  AOI22_X1   g12878(.A1(new_n13068_), .A2(\asqrt[46] ), .B1(new_n13066_), .B2(new_n13063_), .ZN(new_n13071_));
  INV_X1     g12879(.I(new_n12874_), .ZN(new_n13072_));
  OAI21_X1   g12880(.A1(new_n13071_), .A2(new_n2253_), .B(new_n13072_), .ZN(new_n13073_));
  NAND2_X1   g12881(.A1(new_n13073_), .A2(new_n13070_), .ZN(new_n13074_));
  OAI22_X1   g12882(.A1(new_n13071_), .A2(new_n2253_), .B1(new_n13069_), .B2(new_n13067_), .ZN(new_n13075_));
  AOI21_X1   g12883(.A1(new_n13075_), .A2(\asqrt[48] ), .B(new_n12881_), .ZN(new_n13076_));
  NOR2_X1    g12884(.A1(new_n13076_), .A2(new_n13074_), .ZN(new_n13077_));
  AOI22_X1   g12885(.A1(new_n13075_), .A2(\asqrt[48] ), .B1(new_n13073_), .B2(new_n13070_), .ZN(new_n13078_));
  INV_X1     g12886(.I(new_n12889_), .ZN(new_n13079_));
  OAI21_X1   g12887(.A1(new_n13078_), .A2(new_n1854_), .B(new_n13079_), .ZN(new_n13080_));
  NAND2_X1   g12888(.A1(new_n13080_), .A2(new_n13077_), .ZN(new_n13081_));
  OAI22_X1   g12889(.A1(new_n13078_), .A2(new_n1854_), .B1(new_n13076_), .B2(new_n13074_), .ZN(new_n13082_));
  AOI21_X1   g12890(.A1(new_n13082_), .A2(\asqrt[50] ), .B(new_n12896_), .ZN(new_n13083_));
  NOR2_X1    g12891(.A1(new_n13083_), .A2(new_n13081_), .ZN(new_n13084_));
  AOI22_X1   g12892(.A1(new_n13082_), .A2(\asqrt[50] ), .B1(new_n13080_), .B2(new_n13077_), .ZN(new_n13085_));
  INV_X1     g12893(.I(new_n12904_), .ZN(new_n13086_));
  OAI21_X1   g12894(.A1(new_n13085_), .A2(new_n1436_), .B(new_n13086_), .ZN(new_n13087_));
  NAND2_X1   g12895(.A1(new_n13087_), .A2(new_n13084_), .ZN(new_n13088_));
  OAI22_X1   g12896(.A1(new_n13085_), .A2(new_n1436_), .B1(new_n13083_), .B2(new_n13081_), .ZN(new_n13089_));
  AOI21_X1   g12897(.A1(new_n13089_), .A2(\asqrt[52] ), .B(new_n12911_), .ZN(new_n13090_));
  NOR2_X1    g12898(.A1(new_n13090_), .A2(new_n13088_), .ZN(new_n13091_));
  AOI22_X1   g12899(.A1(new_n13089_), .A2(\asqrt[52] ), .B1(new_n13087_), .B2(new_n13084_), .ZN(new_n13092_));
  INV_X1     g12900(.I(new_n12918_), .ZN(new_n13093_));
  OAI21_X1   g12901(.A1(new_n13092_), .A2(new_n1096_), .B(new_n13093_), .ZN(new_n13094_));
  NAND2_X1   g12902(.A1(new_n13094_), .A2(new_n13091_), .ZN(new_n13095_));
  OAI22_X1   g12903(.A1(new_n13092_), .A2(new_n1096_), .B1(new_n13090_), .B2(new_n13088_), .ZN(new_n13096_));
  AOI21_X1   g12904(.A1(new_n13096_), .A2(\asqrt[54] ), .B(new_n12924_), .ZN(new_n13097_));
  NOR2_X1    g12905(.A1(new_n13097_), .A2(new_n13095_), .ZN(new_n13098_));
  AOI22_X1   g12906(.A1(new_n13096_), .A2(\asqrt[54] ), .B1(new_n13094_), .B2(new_n13091_), .ZN(new_n13099_));
  INV_X1     g12907(.I(new_n12931_), .ZN(new_n13100_));
  OAI21_X1   g12908(.A1(new_n13099_), .A2(new_n825_), .B(new_n13100_), .ZN(new_n13101_));
  NAND2_X1   g12909(.A1(new_n13101_), .A2(new_n13098_), .ZN(new_n13102_));
  OAI22_X1   g12910(.A1(new_n13099_), .A2(new_n825_), .B1(new_n13097_), .B2(new_n13095_), .ZN(new_n13103_));
  AOI21_X1   g12911(.A1(new_n13103_), .A2(\asqrt[56] ), .B(new_n12937_), .ZN(new_n13104_));
  NOR2_X1    g12912(.A1(new_n13104_), .A2(new_n13102_), .ZN(new_n13105_));
  AOI22_X1   g12913(.A1(new_n13103_), .A2(\asqrt[56] ), .B1(new_n13101_), .B2(new_n13098_), .ZN(new_n13106_));
  INV_X1     g12914(.I(new_n12944_), .ZN(new_n13107_));
  OAI21_X1   g12915(.A1(new_n13106_), .A2(new_n587_), .B(new_n13107_), .ZN(new_n13108_));
  NAND2_X1   g12916(.A1(new_n13108_), .A2(new_n13105_), .ZN(new_n13109_));
  OAI22_X1   g12917(.A1(new_n13106_), .A2(new_n587_), .B1(new_n13104_), .B2(new_n13102_), .ZN(new_n13110_));
  AOI21_X1   g12918(.A1(new_n13110_), .A2(\asqrt[58] ), .B(new_n12950_), .ZN(new_n13111_));
  NOR2_X1    g12919(.A1(new_n13111_), .A2(new_n13109_), .ZN(new_n13112_));
  AOI22_X1   g12920(.A1(new_n13110_), .A2(\asqrt[58] ), .B1(new_n13108_), .B2(new_n13105_), .ZN(new_n13113_));
  INV_X1     g12921(.I(new_n12957_), .ZN(new_n13114_));
  OAI21_X1   g12922(.A1(new_n13113_), .A2(new_n376_), .B(new_n13114_), .ZN(new_n13115_));
  NAND2_X1   g12923(.A1(new_n13115_), .A2(new_n13112_), .ZN(new_n13116_));
  OAI22_X1   g12924(.A1(new_n13113_), .A2(new_n376_), .B1(new_n13111_), .B2(new_n13109_), .ZN(new_n13117_));
  AOI22_X1   g12925(.A1(new_n13117_), .A2(\asqrt[60] ), .B1(new_n13115_), .B2(new_n13112_), .ZN(new_n13118_));
  AOI21_X1   g12926(.A1(new_n13117_), .A2(\asqrt[60] ), .B(new_n12964_), .ZN(new_n13119_));
  OAI22_X1   g12927(.A1(new_n13118_), .A2(new_n229_), .B1(new_n13119_), .B2(new_n13116_), .ZN(new_n13120_));
  NOR2_X1    g12928(.A1(new_n13120_), .A2(\asqrt[62] ), .ZN(new_n13121_));
  NAND3_X1   g12929(.A1(new_n12651_), .A2(new_n12441_), .A3(new_n12619_), .ZN(new_n13122_));
  NOR2_X1    g12930(.A1(new_n12660_), .A2(new_n196_), .ZN(new_n13123_));
  INV_X1     g12931(.I(new_n12645_), .ZN(new_n13124_));
  NAND3_X1   g12932(.A1(\asqrt[19] ), .A2(new_n13123_), .A3(new_n13124_), .ZN(new_n13125_));
  OAI21_X1   g12933(.A1(new_n12616_), .A2(\asqrt[62] ), .B(new_n12443_), .ZN(new_n13126_));
  OAI21_X1   g12934(.A1(\asqrt[19] ), .A2(new_n13126_), .B(new_n13123_), .ZN(new_n13127_));
  NAND2_X1   g12935(.A1(new_n13127_), .A2(new_n13125_), .ZN(new_n13128_));
  INV_X1     g12936(.I(new_n13128_), .ZN(new_n13129_));
  NOR2_X1    g12937(.A1(new_n12624_), .A2(new_n196_), .ZN(new_n13130_));
  INV_X1     g12938(.I(new_n13130_), .ZN(new_n13131_));
  NAND2_X1   g12939(.A1(new_n12941_), .A2(\asqrt[57] ), .ZN(new_n13132_));
  AOI21_X1   g12940(.A1(new_n13132_), .A2(new_n12940_), .B(new_n504_), .ZN(new_n13133_));
  OAI21_X1   g12941(.A1(new_n12946_), .A2(new_n13133_), .B(\asqrt[59] ), .ZN(new_n13134_));
  AOI21_X1   g12942(.A1(new_n12953_), .A2(new_n13134_), .B(new_n275_), .ZN(new_n13135_));
  OAI21_X1   g12943(.A1(new_n12959_), .A2(new_n13135_), .B(\asqrt[61] ), .ZN(new_n13136_));
  NOR2_X1    g12944(.A1(new_n12625_), .A2(\asqrt[62] ), .ZN(new_n13137_));
  INV_X1     g12945(.I(new_n13137_), .ZN(new_n13138_));
  NAND3_X1   g12946(.A1(new_n12966_), .A2(new_n12959_), .A3(new_n13138_), .ZN(new_n13139_));
  OAI21_X1   g12947(.A1(new_n13139_), .A2(new_n13136_), .B(new_n13131_), .ZN(new_n13140_));
  NAND3_X1   g12948(.A1(new_n12657_), .A2(new_n12612_), .A3(new_n12661_), .ZN(new_n13141_));
  AOI21_X1   g12949(.A1(new_n13141_), .A2(new_n12604_), .B(\asqrt[63] ), .ZN(new_n13142_));
  INV_X1     g12950(.I(new_n13142_), .ZN(new_n13143_));
  OAI21_X1   g12951(.A1(new_n13140_), .A2(new_n13143_), .B(new_n13129_), .ZN(new_n13144_));
  NOR4_X1    g12952(.A1(new_n13120_), .A2(\asqrt[62] ), .A3(new_n13128_), .A4(new_n12624_), .ZN(new_n13145_));
  NAND2_X1   g12953(.A1(new_n12639_), .A2(new_n12612_), .ZN(new_n13146_));
  XOR2_X1    g12954(.A1(new_n12639_), .A2(\asqrt[63] ), .Z(new_n13147_));
  AOI21_X1   g12955(.A1(\asqrt[19] ), .A2(new_n13146_), .B(new_n13147_), .ZN(new_n13148_));
  NAND2_X1   g12956(.A1(new_n13145_), .A2(new_n13148_), .ZN(new_n13149_));
  NOR3_X1    g12957(.A1(new_n13149_), .A2(new_n13122_), .A3(new_n13144_), .ZN(\asqrt[18] ));
  NAND4_X1   g12958(.A1(\asqrt[18] ), .A2(new_n12625_), .A3(new_n12968_), .A4(new_n13121_), .ZN(new_n13151_));
  OAI21_X1   g12959(.A1(new_n13120_), .A2(\asqrt[62] ), .B(new_n12624_), .ZN(new_n13152_));
  OAI21_X1   g12960(.A1(\asqrt[18] ), .A2(new_n13152_), .B(new_n12968_), .ZN(new_n13153_));
  NAND2_X1   g12961(.A1(new_n13151_), .A2(new_n13153_), .ZN(new_n13154_));
  INV_X1     g12962(.I(new_n13154_), .ZN(new_n13155_));
  NAND2_X1   g12963(.A1(new_n13110_), .A2(\asqrt[58] ), .ZN(new_n13156_));
  AOI21_X1   g12964(.A1(new_n13156_), .A2(new_n13109_), .B(new_n376_), .ZN(new_n13157_));
  OAI21_X1   g12965(.A1(new_n13112_), .A2(new_n13157_), .B(\asqrt[60] ), .ZN(new_n13158_));
  AOI21_X1   g12966(.A1(new_n13116_), .A2(new_n13158_), .B(new_n229_), .ZN(new_n13159_));
  NOR3_X1    g12967(.A1(new_n12961_), .A2(\asqrt[61] ), .A3(new_n12963_), .ZN(new_n13160_));
  NAND2_X1   g12968(.A1(\asqrt[18] ), .A2(new_n13160_), .ZN(new_n13161_));
  XOR2_X1    g12969(.A1(new_n13161_), .A2(new_n13159_), .Z(new_n13162_));
  NOR2_X1    g12970(.A1(new_n13162_), .A2(new_n196_), .ZN(new_n13163_));
  INV_X1     g12971(.I(new_n13163_), .ZN(new_n13164_));
  INV_X1     g12972(.I(\a[36] ), .ZN(new_n13165_));
  NOR2_X1    g12973(.A1(\a[34] ), .A2(\a[35] ), .ZN(new_n13166_));
  INV_X1     g12974(.I(new_n13166_), .ZN(new_n13167_));
  NOR3_X1    g12975(.A1(new_n12663_), .A2(new_n13165_), .A3(new_n13167_), .ZN(new_n13168_));
  NAND2_X1   g12976(.A1(new_n12669_), .A2(new_n13168_), .ZN(new_n13169_));
  XOR2_X1    g12977(.A1(new_n13169_), .A2(\a[37] ), .Z(new_n13170_));
  INV_X1     g12978(.I(\a[37] ), .ZN(new_n13171_));
  NOR4_X1    g12979(.A1(new_n13149_), .A2(new_n13171_), .A3(new_n13122_), .A4(new_n13144_), .ZN(new_n13172_));
  NOR2_X1    g12980(.A1(new_n13171_), .A2(\a[36] ), .ZN(new_n13173_));
  OAI21_X1   g12981(.A1(new_n13172_), .A2(new_n13173_), .B(new_n13170_), .ZN(new_n13174_));
  INV_X1     g12982(.I(new_n13170_), .ZN(new_n13175_));
  INV_X1     g12983(.I(new_n13122_), .ZN(new_n13176_));
  NOR3_X1    g12984(.A1(new_n13119_), .A2(new_n13116_), .A3(new_n13137_), .ZN(new_n13177_));
  AOI21_X1   g12985(.A1(new_n13177_), .A2(new_n13159_), .B(new_n13130_), .ZN(new_n13178_));
  AOI21_X1   g12986(.A1(new_n13178_), .A2(new_n13142_), .B(new_n13128_), .ZN(new_n13179_));
  NAND4_X1   g12987(.A1(new_n12967_), .A2(new_n196_), .A3(new_n13129_), .A4(new_n12625_), .ZN(new_n13180_));
  INV_X1     g12988(.I(new_n13148_), .ZN(new_n13181_));
  NOR2_X1    g12989(.A1(new_n13180_), .A2(new_n13181_), .ZN(new_n13182_));
  NAND4_X1   g12990(.A1(new_n13182_), .A2(\a[37] ), .A3(new_n13179_), .A4(new_n13176_), .ZN(new_n13183_));
  NAND3_X1   g12991(.A1(new_n13183_), .A2(\a[36] ), .A3(new_n13175_), .ZN(new_n13184_));
  NAND2_X1   g12992(.A1(new_n13174_), .A2(new_n13184_), .ZN(new_n13185_));
  NOR2_X1    g12993(.A1(new_n13149_), .A2(new_n13144_), .ZN(new_n13186_));
  NOR4_X1    g12994(.A1(new_n12618_), .A2(new_n12612_), .A3(new_n12659_), .A4(new_n12619_), .ZN(new_n13187_));
  NAND2_X1   g12995(.A1(\asqrt[19] ), .A2(\a[36] ), .ZN(new_n13188_));
  XOR2_X1    g12996(.A1(new_n13188_), .A2(new_n13187_), .Z(new_n13189_));
  NOR2_X1    g12997(.A1(new_n13189_), .A2(new_n13167_), .ZN(new_n13190_));
  INV_X1     g12998(.I(new_n13190_), .ZN(new_n13191_));
  NAND3_X1   g12999(.A1(new_n13182_), .A2(new_n13176_), .A3(new_n13179_), .ZN(new_n13192_));
  NOR2_X1    g13000(.A1(new_n13176_), .A2(new_n13148_), .ZN(new_n13193_));
  INV_X1     g13001(.I(new_n13193_), .ZN(new_n13194_));
  NOR2_X1    g13002(.A1(new_n13194_), .A2(new_n12657_), .ZN(new_n13195_));
  NAND3_X1   g13003(.A1(new_n13144_), .A2(new_n13180_), .A3(new_n13195_), .ZN(new_n13196_));
  NAND2_X1   g13004(.A1(new_n13196_), .A2(new_n12626_), .ZN(new_n13197_));
  NAND3_X1   g13005(.A1(new_n13197_), .A2(new_n12627_), .A3(new_n13192_), .ZN(new_n13198_));
  INV_X1     g13006(.I(new_n13195_), .ZN(new_n13199_));
  NOR3_X1    g13007(.A1(new_n13179_), .A2(new_n13145_), .A3(new_n13199_), .ZN(new_n13200_));
  OAI21_X1   g13008(.A1(new_n13200_), .A2(\a[38] ), .B(new_n12627_), .ZN(new_n13201_));
  NAND2_X1   g13009(.A1(new_n13201_), .A2(\asqrt[18] ), .ZN(new_n13202_));
  NAND4_X1   g13010(.A1(new_n13202_), .A2(new_n12101_), .A3(new_n13198_), .A4(new_n13191_), .ZN(new_n13203_));
  NAND2_X1   g13011(.A1(new_n13203_), .A2(new_n13185_), .ZN(new_n13204_));
  NAND3_X1   g13012(.A1(new_n13174_), .A2(new_n13184_), .A3(new_n13191_), .ZN(new_n13205_));
  AOI21_X1   g13013(.A1(\asqrt[19] ), .A2(new_n12626_), .B(\a[39] ), .ZN(new_n13206_));
  NOR2_X1    g13014(.A1(new_n12648_), .A2(\a[38] ), .ZN(new_n13207_));
  AOI21_X1   g13015(.A1(\asqrt[19] ), .A2(\a[38] ), .B(new_n12630_), .ZN(new_n13208_));
  OAI21_X1   g13016(.A1(new_n13207_), .A2(new_n13206_), .B(new_n13208_), .ZN(new_n13209_));
  INV_X1     g13017(.I(new_n13209_), .ZN(new_n13210_));
  NAND3_X1   g13018(.A1(\asqrt[18] ), .A2(new_n12656_), .A3(new_n13210_), .ZN(new_n13211_));
  OAI21_X1   g13019(.A1(new_n13192_), .A2(new_n13209_), .B(new_n12655_), .ZN(new_n13212_));
  NAND3_X1   g13020(.A1(new_n13211_), .A2(new_n13212_), .A3(new_n11631_), .ZN(new_n13213_));
  AOI21_X1   g13021(.A1(new_n13205_), .A2(\asqrt[20] ), .B(new_n13213_), .ZN(new_n13214_));
  NOR2_X1    g13022(.A1(new_n13204_), .A2(new_n13214_), .ZN(new_n13215_));
  AOI22_X1   g13023(.A1(new_n13203_), .A2(new_n13185_), .B1(\asqrt[20] ), .B2(new_n13205_), .ZN(new_n13216_));
  NOR2_X1    g13024(.A1(new_n12974_), .A2(new_n12973_), .ZN(new_n13217_));
  NOR4_X1    g13025(.A1(new_n13192_), .A2(\asqrt[21] ), .A3(new_n13217_), .A4(new_n12675_), .ZN(new_n13218_));
  AOI21_X1   g13026(.A1(new_n12972_), .A2(new_n12656_), .B(new_n11631_), .ZN(new_n13219_));
  NOR2_X1    g13027(.A1(new_n13218_), .A2(new_n13219_), .ZN(new_n13220_));
  NAND2_X1   g13028(.A1(new_n13220_), .A2(new_n11105_), .ZN(new_n13221_));
  INV_X1     g13029(.I(new_n13221_), .ZN(new_n13222_));
  OAI21_X1   g13030(.A1(new_n13216_), .A2(new_n11631_), .B(new_n13222_), .ZN(new_n13223_));
  NAND2_X1   g13031(.A1(new_n13205_), .A2(\asqrt[20] ), .ZN(new_n13224_));
  AOI21_X1   g13032(.A1(new_n13204_), .A2(new_n13224_), .B(new_n11631_), .ZN(new_n13225_));
  OAI21_X1   g13033(.A1(new_n13225_), .A2(new_n13215_), .B(\asqrt[22] ), .ZN(new_n13226_));
  NOR2_X1    g13034(.A1(new_n12687_), .A2(new_n11105_), .ZN(new_n13227_));
  NAND2_X1   g13035(.A1(new_n12681_), .A2(new_n12683_), .ZN(new_n13228_));
  NAND4_X1   g13036(.A1(\asqrt[18] ), .A2(new_n11105_), .A3(new_n13228_), .A4(new_n12687_), .ZN(new_n13229_));
  XOR2_X1    g13037(.A1(new_n13229_), .A2(new_n13227_), .Z(new_n13230_));
  NAND2_X1   g13038(.A1(new_n13230_), .A2(new_n10614_), .ZN(new_n13231_));
  INV_X1     g13039(.I(new_n13231_), .ZN(new_n13232_));
  NAND2_X1   g13040(.A1(new_n13226_), .A2(new_n13232_), .ZN(new_n13233_));
  NAND3_X1   g13041(.A1(new_n13233_), .A2(new_n13215_), .A3(new_n13223_), .ZN(new_n13234_));
  INV_X1     g13042(.I(new_n13173_), .ZN(new_n13235_));
  AOI21_X1   g13043(.A1(new_n13183_), .A2(new_n13235_), .B(new_n13175_), .ZN(new_n13236_));
  NOR3_X1    g13044(.A1(new_n13172_), .A2(new_n13165_), .A3(new_n13170_), .ZN(new_n13237_));
  NOR2_X1    g13045(.A1(new_n13237_), .A2(new_n13236_), .ZN(new_n13238_));
  NOR2_X1    g13046(.A1(new_n13201_), .A2(\asqrt[18] ), .ZN(new_n13239_));
  AOI21_X1   g13047(.A1(new_n13197_), .A2(new_n12627_), .B(new_n13192_), .ZN(new_n13240_));
  NOR4_X1    g13048(.A1(new_n13239_), .A2(new_n13240_), .A3(\asqrt[20] ), .A4(new_n13190_), .ZN(new_n13241_));
  NOR2_X1    g13049(.A1(new_n13241_), .A2(new_n13238_), .ZN(new_n13242_));
  NOR3_X1    g13050(.A1(new_n13237_), .A2(new_n13236_), .A3(new_n13190_), .ZN(new_n13243_));
  NOR3_X1    g13051(.A1(new_n13192_), .A2(new_n12655_), .A3(new_n13209_), .ZN(new_n13244_));
  AOI21_X1   g13052(.A1(\asqrt[18] ), .A2(new_n13210_), .B(new_n12656_), .ZN(new_n13245_));
  NOR3_X1    g13053(.A1(new_n13245_), .A2(new_n13244_), .A3(\asqrt[21] ), .ZN(new_n13246_));
  OAI21_X1   g13054(.A1(new_n13243_), .A2(new_n12101_), .B(new_n13246_), .ZN(new_n13247_));
  NAND2_X1   g13055(.A1(new_n13242_), .A2(new_n13247_), .ZN(new_n13248_));
  OAI22_X1   g13056(.A1(new_n13241_), .A2(new_n13238_), .B1(new_n12101_), .B2(new_n13243_), .ZN(new_n13249_));
  AOI21_X1   g13057(.A1(new_n13249_), .A2(\asqrt[21] ), .B(new_n13221_), .ZN(new_n13250_));
  AOI22_X1   g13058(.A1(new_n13249_), .A2(\asqrt[21] ), .B1(new_n13242_), .B2(new_n13247_), .ZN(new_n13251_));
  OAI22_X1   g13059(.A1(new_n13251_), .A2(new_n11105_), .B1(new_n13250_), .B2(new_n13248_), .ZN(new_n13252_));
  NAND2_X1   g13060(.A1(new_n12694_), .A2(\asqrt[23] ), .ZN(new_n13253_));
  NOR2_X1    g13061(.A1(new_n12689_), .A2(new_n12690_), .ZN(new_n13254_));
  NOR4_X1    g13062(.A1(new_n13192_), .A2(\asqrt[23] ), .A3(new_n13254_), .A4(new_n12694_), .ZN(new_n13255_));
  XOR2_X1    g13063(.A1(new_n13255_), .A2(new_n13253_), .Z(new_n13256_));
  NAND2_X1   g13064(.A1(new_n13256_), .A2(new_n10104_), .ZN(new_n13257_));
  AOI21_X1   g13065(.A1(new_n13252_), .A2(\asqrt[23] ), .B(new_n13257_), .ZN(new_n13258_));
  NOR2_X1    g13066(.A1(new_n13258_), .A2(new_n13234_), .ZN(new_n13259_));
  OAI21_X1   g13067(.A1(new_n13225_), .A2(new_n13221_), .B(new_n13215_), .ZN(new_n13260_));
  AOI21_X1   g13068(.A1(new_n13226_), .A2(new_n13232_), .B(new_n13260_), .ZN(new_n13261_));
  AOI21_X1   g13069(.A1(new_n13260_), .A2(new_n13226_), .B(new_n10614_), .ZN(new_n13262_));
  OAI21_X1   g13070(.A1(new_n13261_), .A2(new_n13262_), .B(\asqrt[24] ), .ZN(new_n13263_));
  NOR4_X1    g13071(.A1(new_n13192_), .A2(\asqrt[24] ), .A3(new_n12697_), .A4(new_n12991_), .ZN(new_n13264_));
  AOI21_X1   g13072(.A1(new_n13253_), .A2(new_n12693_), .B(new_n10104_), .ZN(new_n13265_));
  NOR2_X1    g13073(.A1(new_n13264_), .A2(new_n13265_), .ZN(new_n13266_));
  NAND2_X1   g13074(.A1(new_n13266_), .A2(new_n9672_), .ZN(new_n13267_));
  INV_X1     g13075(.I(new_n13267_), .ZN(new_n13268_));
  NAND2_X1   g13076(.A1(new_n13263_), .A2(new_n13268_), .ZN(new_n13269_));
  NAND2_X1   g13077(.A1(new_n13269_), .A2(new_n13259_), .ZN(new_n13270_));
  NOR2_X1    g13078(.A1(new_n13261_), .A2(new_n13262_), .ZN(new_n13271_));
  OAI22_X1   g13079(.A1(new_n13271_), .A2(new_n10104_), .B1(new_n13258_), .B2(new_n13234_), .ZN(new_n13272_));
  NAND2_X1   g13080(.A1(new_n12709_), .A2(\asqrt[25] ), .ZN(new_n13273_));
  NOR4_X1    g13081(.A1(new_n13192_), .A2(\asqrt[25] ), .A3(new_n12704_), .A4(new_n12709_), .ZN(new_n13274_));
  XOR2_X1    g13082(.A1(new_n13274_), .A2(new_n13273_), .Z(new_n13275_));
  NAND2_X1   g13083(.A1(new_n13275_), .A2(new_n9212_), .ZN(new_n13276_));
  AOI21_X1   g13084(.A1(new_n13272_), .A2(\asqrt[25] ), .B(new_n13276_), .ZN(new_n13277_));
  NOR2_X1    g13085(.A1(new_n13277_), .A2(new_n13270_), .ZN(new_n13278_));
  OAI21_X1   g13086(.A1(new_n13262_), .A2(new_n13257_), .B(new_n13261_), .ZN(new_n13279_));
  AOI21_X1   g13087(.A1(new_n13263_), .A2(new_n13268_), .B(new_n13279_), .ZN(new_n13280_));
  AOI21_X1   g13088(.A1(new_n13279_), .A2(new_n13263_), .B(new_n9672_), .ZN(new_n13281_));
  OAI21_X1   g13089(.A1(new_n13280_), .A2(new_n13281_), .B(\asqrt[26] ), .ZN(new_n13282_));
  NOR4_X1    g13090(.A1(new_n13192_), .A2(\asqrt[26] ), .A3(new_n12711_), .A4(new_n12998_), .ZN(new_n13283_));
  AOI21_X1   g13091(.A1(new_n13273_), .A2(new_n12708_), .B(new_n9212_), .ZN(new_n13284_));
  NOR2_X1    g13092(.A1(new_n13283_), .A2(new_n13284_), .ZN(new_n13285_));
  NAND2_X1   g13093(.A1(new_n13285_), .A2(new_n8763_), .ZN(new_n13286_));
  INV_X1     g13094(.I(new_n13286_), .ZN(new_n13287_));
  NAND2_X1   g13095(.A1(new_n13282_), .A2(new_n13287_), .ZN(new_n13288_));
  NAND2_X1   g13096(.A1(new_n13288_), .A2(new_n13278_), .ZN(new_n13289_));
  AOI22_X1   g13097(.A1(new_n13272_), .A2(\asqrt[25] ), .B1(new_n13269_), .B2(new_n13259_), .ZN(new_n13290_));
  OAI22_X1   g13098(.A1(new_n13290_), .A2(new_n9212_), .B1(new_n13277_), .B2(new_n13270_), .ZN(new_n13291_));
  NAND2_X1   g13099(.A1(new_n12722_), .A2(\asqrt[27] ), .ZN(new_n13292_));
  NOR4_X1    g13100(.A1(new_n13192_), .A2(\asqrt[27] ), .A3(new_n12717_), .A4(new_n12722_), .ZN(new_n13293_));
  XOR2_X1    g13101(.A1(new_n13293_), .A2(new_n13292_), .Z(new_n13294_));
  NAND2_X1   g13102(.A1(new_n13294_), .A2(new_n8319_), .ZN(new_n13295_));
  AOI21_X1   g13103(.A1(new_n13291_), .A2(\asqrt[27] ), .B(new_n13295_), .ZN(new_n13296_));
  NOR2_X1    g13104(.A1(new_n13296_), .A2(new_n13289_), .ZN(new_n13297_));
  AOI22_X1   g13105(.A1(new_n13291_), .A2(\asqrt[27] ), .B1(new_n13288_), .B2(new_n13278_), .ZN(new_n13298_));
  NOR4_X1    g13106(.A1(new_n13192_), .A2(\asqrt[28] ), .A3(new_n12724_), .A4(new_n13005_), .ZN(new_n13299_));
  AOI21_X1   g13107(.A1(new_n13292_), .A2(new_n12721_), .B(new_n8319_), .ZN(new_n13300_));
  NOR2_X1    g13108(.A1(new_n13299_), .A2(new_n13300_), .ZN(new_n13301_));
  NAND2_X1   g13109(.A1(new_n13301_), .A2(new_n7931_), .ZN(new_n13302_));
  INV_X1     g13110(.I(new_n13302_), .ZN(new_n13303_));
  OAI21_X1   g13111(.A1(new_n13298_), .A2(new_n8319_), .B(new_n13303_), .ZN(new_n13304_));
  NAND2_X1   g13112(.A1(new_n13304_), .A2(new_n13297_), .ZN(new_n13305_));
  OAI22_X1   g13113(.A1(new_n13298_), .A2(new_n8319_), .B1(new_n13296_), .B2(new_n13289_), .ZN(new_n13306_));
  NAND2_X1   g13114(.A1(new_n12735_), .A2(\asqrt[29] ), .ZN(new_n13307_));
  NOR4_X1    g13115(.A1(new_n13192_), .A2(\asqrt[29] ), .A3(new_n12730_), .A4(new_n12735_), .ZN(new_n13308_));
  XOR2_X1    g13116(.A1(new_n13308_), .A2(new_n13307_), .Z(new_n13309_));
  NAND2_X1   g13117(.A1(new_n13309_), .A2(new_n7517_), .ZN(new_n13310_));
  AOI21_X1   g13118(.A1(new_n13306_), .A2(\asqrt[29] ), .B(new_n13310_), .ZN(new_n13311_));
  NOR2_X1    g13119(.A1(new_n13311_), .A2(new_n13305_), .ZN(new_n13312_));
  AOI22_X1   g13120(.A1(new_n13306_), .A2(\asqrt[29] ), .B1(new_n13304_), .B2(new_n13297_), .ZN(new_n13313_));
  NAND2_X1   g13121(.A1(new_n13012_), .A2(\asqrt[30] ), .ZN(new_n13314_));
  NOR4_X1    g13122(.A1(new_n13192_), .A2(\asqrt[30] ), .A3(new_n12738_), .A4(new_n13012_), .ZN(new_n13315_));
  XOR2_X1    g13123(.A1(new_n13315_), .A2(new_n13314_), .Z(new_n13316_));
  NAND2_X1   g13124(.A1(new_n13316_), .A2(new_n7110_), .ZN(new_n13317_));
  INV_X1     g13125(.I(new_n13317_), .ZN(new_n13318_));
  OAI21_X1   g13126(.A1(new_n13313_), .A2(new_n7517_), .B(new_n13318_), .ZN(new_n13319_));
  NAND2_X1   g13127(.A1(new_n13319_), .A2(new_n13312_), .ZN(new_n13320_));
  OAI22_X1   g13128(.A1(new_n13313_), .A2(new_n7517_), .B1(new_n13311_), .B2(new_n13305_), .ZN(new_n13321_));
  NOR4_X1    g13129(.A1(new_n13192_), .A2(\asqrt[31] ), .A3(new_n12745_), .A4(new_n12750_), .ZN(new_n13322_));
  AOI21_X1   g13130(.A1(new_n13314_), .A2(new_n13011_), .B(new_n7110_), .ZN(new_n13323_));
  NOR2_X1    g13131(.A1(new_n13322_), .A2(new_n13323_), .ZN(new_n13324_));
  NAND2_X1   g13132(.A1(new_n13324_), .A2(new_n6708_), .ZN(new_n13325_));
  AOI21_X1   g13133(.A1(new_n13321_), .A2(\asqrt[31] ), .B(new_n13325_), .ZN(new_n13326_));
  NOR2_X1    g13134(.A1(new_n13326_), .A2(new_n13320_), .ZN(new_n13327_));
  AOI22_X1   g13135(.A1(new_n13321_), .A2(\asqrt[31] ), .B1(new_n13319_), .B2(new_n13312_), .ZN(new_n13328_));
  NAND2_X1   g13136(.A1(new_n13019_), .A2(\asqrt[32] ), .ZN(new_n13329_));
  NOR4_X1    g13137(.A1(new_n13192_), .A2(\asqrt[32] ), .A3(new_n12753_), .A4(new_n13019_), .ZN(new_n13330_));
  XOR2_X1    g13138(.A1(new_n13330_), .A2(new_n13329_), .Z(new_n13331_));
  NAND2_X1   g13139(.A1(new_n13331_), .A2(new_n6365_), .ZN(new_n13332_));
  INV_X1     g13140(.I(new_n13332_), .ZN(new_n13333_));
  OAI21_X1   g13141(.A1(new_n13328_), .A2(new_n6708_), .B(new_n13333_), .ZN(new_n13334_));
  NAND2_X1   g13142(.A1(new_n13334_), .A2(new_n13327_), .ZN(new_n13335_));
  OAI22_X1   g13143(.A1(new_n13328_), .A2(new_n6708_), .B1(new_n13326_), .B2(new_n13320_), .ZN(new_n13336_));
  NOR4_X1    g13144(.A1(new_n13192_), .A2(\asqrt[33] ), .A3(new_n12760_), .A4(new_n12765_), .ZN(new_n13337_));
  AOI21_X1   g13145(.A1(new_n13329_), .A2(new_n13018_), .B(new_n6365_), .ZN(new_n13338_));
  NOR2_X1    g13146(.A1(new_n13337_), .A2(new_n13338_), .ZN(new_n13339_));
  NAND2_X1   g13147(.A1(new_n13339_), .A2(new_n5991_), .ZN(new_n13340_));
  AOI21_X1   g13148(.A1(new_n13336_), .A2(\asqrt[33] ), .B(new_n13340_), .ZN(new_n13341_));
  NOR2_X1    g13149(.A1(new_n13341_), .A2(new_n13335_), .ZN(new_n13342_));
  AOI22_X1   g13150(.A1(new_n13336_), .A2(\asqrt[33] ), .B1(new_n13334_), .B2(new_n13327_), .ZN(new_n13343_));
  NAND2_X1   g13151(.A1(new_n13026_), .A2(\asqrt[34] ), .ZN(new_n13344_));
  NOR4_X1    g13152(.A1(new_n13192_), .A2(\asqrt[34] ), .A3(new_n12768_), .A4(new_n13026_), .ZN(new_n13345_));
  XOR2_X1    g13153(.A1(new_n13345_), .A2(new_n13344_), .Z(new_n13346_));
  NAND2_X1   g13154(.A1(new_n13346_), .A2(new_n5626_), .ZN(new_n13347_));
  INV_X1     g13155(.I(new_n13347_), .ZN(new_n13348_));
  OAI21_X1   g13156(.A1(new_n13343_), .A2(new_n5991_), .B(new_n13348_), .ZN(new_n13349_));
  NAND2_X1   g13157(.A1(new_n13349_), .A2(new_n13342_), .ZN(new_n13350_));
  OAI22_X1   g13158(.A1(new_n13343_), .A2(new_n5991_), .B1(new_n13341_), .B2(new_n13335_), .ZN(new_n13351_));
  NOR4_X1    g13159(.A1(new_n13192_), .A2(\asqrt[35] ), .A3(new_n12775_), .A4(new_n12780_), .ZN(new_n13352_));
  AOI21_X1   g13160(.A1(new_n13344_), .A2(new_n13025_), .B(new_n5626_), .ZN(new_n13353_));
  NOR2_X1    g13161(.A1(new_n13352_), .A2(new_n13353_), .ZN(new_n13354_));
  NAND2_X1   g13162(.A1(new_n13354_), .A2(new_n5273_), .ZN(new_n13355_));
  AOI21_X1   g13163(.A1(new_n13351_), .A2(\asqrt[35] ), .B(new_n13355_), .ZN(new_n13356_));
  NOR2_X1    g13164(.A1(new_n13356_), .A2(new_n13350_), .ZN(new_n13357_));
  AOI22_X1   g13165(.A1(new_n13351_), .A2(\asqrt[35] ), .B1(new_n13349_), .B2(new_n13342_), .ZN(new_n13358_));
  NAND2_X1   g13166(.A1(new_n13033_), .A2(\asqrt[36] ), .ZN(new_n13359_));
  NOR4_X1    g13167(.A1(new_n13192_), .A2(\asqrt[36] ), .A3(new_n12783_), .A4(new_n13033_), .ZN(new_n13360_));
  XOR2_X1    g13168(.A1(new_n13360_), .A2(new_n13359_), .Z(new_n13361_));
  NAND2_X1   g13169(.A1(new_n13361_), .A2(new_n4973_), .ZN(new_n13362_));
  INV_X1     g13170(.I(new_n13362_), .ZN(new_n13363_));
  OAI21_X1   g13171(.A1(new_n13358_), .A2(new_n5273_), .B(new_n13363_), .ZN(new_n13364_));
  NAND2_X1   g13172(.A1(new_n13364_), .A2(new_n13357_), .ZN(new_n13365_));
  OAI22_X1   g13173(.A1(new_n13358_), .A2(new_n5273_), .B1(new_n13356_), .B2(new_n13350_), .ZN(new_n13366_));
  NOR4_X1    g13174(.A1(new_n13192_), .A2(\asqrt[37] ), .A3(new_n12790_), .A4(new_n12795_), .ZN(new_n13367_));
  AOI21_X1   g13175(.A1(new_n13359_), .A2(new_n13032_), .B(new_n4973_), .ZN(new_n13368_));
  NOR2_X1    g13176(.A1(new_n13367_), .A2(new_n13368_), .ZN(new_n13369_));
  NAND2_X1   g13177(.A1(new_n13369_), .A2(new_n4645_), .ZN(new_n13370_));
  AOI21_X1   g13178(.A1(new_n13366_), .A2(\asqrt[37] ), .B(new_n13370_), .ZN(new_n13371_));
  NOR2_X1    g13179(.A1(new_n13371_), .A2(new_n13365_), .ZN(new_n13372_));
  AOI22_X1   g13180(.A1(new_n13366_), .A2(\asqrt[37] ), .B1(new_n13364_), .B2(new_n13357_), .ZN(new_n13373_));
  NAND2_X1   g13181(.A1(new_n13040_), .A2(\asqrt[38] ), .ZN(new_n13374_));
  NOR4_X1    g13182(.A1(new_n13192_), .A2(\asqrt[38] ), .A3(new_n12798_), .A4(new_n13040_), .ZN(new_n13375_));
  XOR2_X1    g13183(.A1(new_n13375_), .A2(new_n13374_), .Z(new_n13376_));
  NAND2_X1   g13184(.A1(new_n13376_), .A2(new_n4330_), .ZN(new_n13377_));
  INV_X1     g13185(.I(new_n13377_), .ZN(new_n13378_));
  OAI21_X1   g13186(.A1(new_n13373_), .A2(new_n4645_), .B(new_n13378_), .ZN(new_n13379_));
  NAND2_X1   g13187(.A1(new_n13379_), .A2(new_n13372_), .ZN(new_n13380_));
  OAI22_X1   g13188(.A1(new_n13373_), .A2(new_n4645_), .B1(new_n13371_), .B2(new_n13365_), .ZN(new_n13381_));
  NAND2_X1   g13189(.A1(new_n12810_), .A2(\asqrt[39] ), .ZN(new_n13382_));
  NOR4_X1    g13190(.A1(new_n13192_), .A2(\asqrt[39] ), .A3(new_n12805_), .A4(new_n12810_), .ZN(new_n13383_));
  XOR2_X1    g13191(.A1(new_n13383_), .A2(new_n13382_), .Z(new_n13384_));
  NAND2_X1   g13192(.A1(new_n13384_), .A2(new_n4018_), .ZN(new_n13385_));
  AOI21_X1   g13193(.A1(new_n13381_), .A2(\asqrt[39] ), .B(new_n13385_), .ZN(new_n13386_));
  NOR2_X1    g13194(.A1(new_n13386_), .A2(new_n13380_), .ZN(new_n13387_));
  AOI22_X1   g13195(.A1(new_n13381_), .A2(\asqrt[39] ), .B1(new_n13379_), .B2(new_n13372_), .ZN(new_n13388_));
  NOR4_X1    g13196(.A1(new_n13192_), .A2(\asqrt[40] ), .A3(new_n12813_), .A4(new_n13047_), .ZN(new_n13389_));
  AOI21_X1   g13197(.A1(new_n13382_), .A2(new_n12809_), .B(new_n4018_), .ZN(new_n13390_));
  NOR2_X1    g13198(.A1(new_n13389_), .A2(new_n13390_), .ZN(new_n13391_));
  NAND2_X1   g13199(.A1(new_n13391_), .A2(new_n3760_), .ZN(new_n13392_));
  INV_X1     g13200(.I(new_n13392_), .ZN(new_n13393_));
  OAI21_X1   g13201(.A1(new_n13388_), .A2(new_n4018_), .B(new_n13393_), .ZN(new_n13394_));
  NAND2_X1   g13202(.A1(new_n13394_), .A2(new_n13387_), .ZN(new_n13395_));
  OAI22_X1   g13203(.A1(new_n13388_), .A2(new_n4018_), .B1(new_n13386_), .B2(new_n13380_), .ZN(new_n13396_));
  NAND2_X1   g13204(.A1(new_n12825_), .A2(\asqrt[41] ), .ZN(new_n13397_));
  NOR4_X1    g13205(.A1(new_n13192_), .A2(\asqrt[41] ), .A3(new_n12820_), .A4(new_n12825_), .ZN(new_n13398_));
  XOR2_X1    g13206(.A1(new_n13398_), .A2(new_n13397_), .Z(new_n13399_));
  NAND2_X1   g13207(.A1(new_n13399_), .A2(new_n3481_), .ZN(new_n13400_));
  AOI21_X1   g13208(.A1(new_n13396_), .A2(\asqrt[41] ), .B(new_n13400_), .ZN(new_n13401_));
  NOR2_X1    g13209(.A1(new_n13401_), .A2(new_n13395_), .ZN(new_n13402_));
  AOI22_X1   g13210(.A1(new_n13396_), .A2(\asqrt[41] ), .B1(new_n13394_), .B2(new_n13387_), .ZN(new_n13403_));
  NOR4_X1    g13211(.A1(new_n13192_), .A2(\asqrt[42] ), .A3(new_n12828_), .A4(new_n13054_), .ZN(new_n13404_));
  AOI21_X1   g13212(.A1(new_n13397_), .A2(new_n12824_), .B(new_n3481_), .ZN(new_n13405_));
  NOR2_X1    g13213(.A1(new_n13404_), .A2(new_n13405_), .ZN(new_n13406_));
  NAND2_X1   g13214(.A1(new_n13406_), .A2(new_n3208_), .ZN(new_n13407_));
  INV_X1     g13215(.I(new_n13407_), .ZN(new_n13408_));
  OAI21_X1   g13216(.A1(new_n13403_), .A2(new_n3481_), .B(new_n13408_), .ZN(new_n13409_));
  NAND2_X1   g13217(.A1(new_n13409_), .A2(new_n13402_), .ZN(new_n13410_));
  OAI22_X1   g13218(.A1(new_n13403_), .A2(new_n3481_), .B1(new_n13401_), .B2(new_n13395_), .ZN(new_n13411_));
  NAND2_X1   g13219(.A1(new_n12840_), .A2(\asqrt[43] ), .ZN(new_n13412_));
  NOR4_X1    g13220(.A1(new_n13192_), .A2(\asqrt[43] ), .A3(new_n12835_), .A4(new_n12840_), .ZN(new_n13413_));
  XOR2_X1    g13221(.A1(new_n13413_), .A2(new_n13412_), .Z(new_n13414_));
  NAND2_X1   g13222(.A1(new_n13414_), .A2(new_n2941_), .ZN(new_n13415_));
  AOI21_X1   g13223(.A1(new_n13411_), .A2(\asqrt[43] ), .B(new_n13415_), .ZN(new_n13416_));
  NOR2_X1    g13224(.A1(new_n13416_), .A2(new_n13410_), .ZN(new_n13417_));
  AOI22_X1   g13225(.A1(new_n13411_), .A2(\asqrt[43] ), .B1(new_n13409_), .B2(new_n13402_), .ZN(new_n13418_));
  NAND2_X1   g13226(.A1(new_n13061_), .A2(\asqrt[44] ), .ZN(new_n13419_));
  NOR4_X1    g13227(.A1(new_n13192_), .A2(\asqrt[44] ), .A3(new_n12843_), .A4(new_n13061_), .ZN(new_n13420_));
  XOR2_X1    g13228(.A1(new_n13420_), .A2(new_n13419_), .Z(new_n13421_));
  NAND2_X1   g13229(.A1(new_n13421_), .A2(new_n2728_), .ZN(new_n13422_));
  INV_X1     g13230(.I(new_n13422_), .ZN(new_n13423_));
  OAI21_X1   g13231(.A1(new_n13418_), .A2(new_n2941_), .B(new_n13423_), .ZN(new_n13424_));
  NAND2_X1   g13232(.A1(new_n13424_), .A2(new_n13417_), .ZN(new_n13425_));
  OAI22_X1   g13233(.A1(new_n13418_), .A2(new_n2941_), .B1(new_n13416_), .B2(new_n13410_), .ZN(new_n13426_));
  NOR4_X1    g13234(.A1(new_n13192_), .A2(\asqrt[45] ), .A3(new_n12850_), .A4(new_n12855_), .ZN(new_n13427_));
  AOI21_X1   g13235(.A1(new_n13419_), .A2(new_n13060_), .B(new_n2728_), .ZN(new_n13428_));
  NOR2_X1    g13236(.A1(new_n13427_), .A2(new_n13428_), .ZN(new_n13429_));
  NAND2_X1   g13237(.A1(new_n13429_), .A2(new_n2488_), .ZN(new_n13430_));
  AOI21_X1   g13238(.A1(new_n13426_), .A2(\asqrt[45] ), .B(new_n13430_), .ZN(new_n13431_));
  NOR2_X1    g13239(.A1(new_n13431_), .A2(new_n13425_), .ZN(new_n13432_));
  AOI22_X1   g13240(.A1(new_n13426_), .A2(\asqrt[45] ), .B1(new_n13424_), .B2(new_n13417_), .ZN(new_n13433_));
  NAND2_X1   g13241(.A1(new_n13068_), .A2(\asqrt[46] ), .ZN(new_n13434_));
  NOR4_X1    g13242(.A1(new_n13192_), .A2(\asqrt[46] ), .A3(new_n12858_), .A4(new_n13068_), .ZN(new_n13435_));
  XOR2_X1    g13243(.A1(new_n13435_), .A2(new_n13434_), .Z(new_n13436_));
  NAND2_X1   g13244(.A1(new_n13436_), .A2(new_n2253_), .ZN(new_n13437_));
  INV_X1     g13245(.I(new_n13437_), .ZN(new_n13438_));
  OAI21_X1   g13246(.A1(new_n13433_), .A2(new_n2488_), .B(new_n13438_), .ZN(new_n13439_));
  NAND2_X1   g13247(.A1(new_n13439_), .A2(new_n13432_), .ZN(new_n13440_));
  OAI22_X1   g13248(.A1(new_n13433_), .A2(new_n2488_), .B1(new_n13431_), .B2(new_n13425_), .ZN(new_n13441_));
  NOR4_X1    g13249(.A1(new_n13192_), .A2(\asqrt[47] ), .A3(new_n12865_), .A4(new_n12870_), .ZN(new_n13442_));
  AOI21_X1   g13250(.A1(new_n13434_), .A2(new_n13067_), .B(new_n2253_), .ZN(new_n13443_));
  NOR2_X1    g13251(.A1(new_n13442_), .A2(new_n13443_), .ZN(new_n13444_));
  NAND2_X1   g13252(.A1(new_n13444_), .A2(new_n2046_), .ZN(new_n13445_));
  AOI21_X1   g13253(.A1(new_n13441_), .A2(\asqrt[47] ), .B(new_n13445_), .ZN(new_n13446_));
  NOR2_X1    g13254(.A1(new_n13446_), .A2(new_n13440_), .ZN(new_n13447_));
  AOI22_X1   g13255(.A1(new_n13441_), .A2(\asqrt[47] ), .B1(new_n13439_), .B2(new_n13432_), .ZN(new_n13448_));
  NAND2_X1   g13256(.A1(new_n13075_), .A2(\asqrt[48] ), .ZN(new_n13449_));
  NOR4_X1    g13257(.A1(new_n13192_), .A2(\asqrt[48] ), .A3(new_n12873_), .A4(new_n13075_), .ZN(new_n13450_));
  XOR2_X1    g13258(.A1(new_n13450_), .A2(new_n13449_), .Z(new_n13451_));
  NAND2_X1   g13259(.A1(new_n13451_), .A2(new_n1854_), .ZN(new_n13452_));
  INV_X1     g13260(.I(new_n13452_), .ZN(new_n13453_));
  OAI21_X1   g13261(.A1(new_n13448_), .A2(new_n2046_), .B(new_n13453_), .ZN(new_n13454_));
  NAND2_X1   g13262(.A1(new_n13454_), .A2(new_n13447_), .ZN(new_n13455_));
  OAI22_X1   g13263(.A1(new_n13448_), .A2(new_n2046_), .B1(new_n13446_), .B2(new_n13440_), .ZN(new_n13456_));
  NOR4_X1    g13264(.A1(new_n13192_), .A2(\asqrt[49] ), .A3(new_n12880_), .A4(new_n12885_), .ZN(new_n13457_));
  AOI21_X1   g13265(.A1(new_n13449_), .A2(new_n13074_), .B(new_n1854_), .ZN(new_n13458_));
  NOR2_X1    g13266(.A1(new_n13457_), .A2(new_n13458_), .ZN(new_n13459_));
  NAND2_X1   g13267(.A1(new_n13459_), .A2(new_n1595_), .ZN(new_n13460_));
  AOI21_X1   g13268(.A1(new_n13456_), .A2(\asqrt[49] ), .B(new_n13460_), .ZN(new_n13461_));
  NOR2_X1    g13269(.A1(new_n13461_), .A2(new_n13455_), .ZN(new_n13462_));
  AOI22_X1   g13270(.A1(new_n13456_), .A2(\asqrt[49] ), .B1(new_n13454_), .B2(new_n13447_), .ZN(new_n13463_));
  NAND2_X1   g13271(.A1(new_n13082_), .A2(\asqrt[50] ), .ZN(new_n13464_));
  NOR4_X1    g13272(.A1(new_n13192_), .A2(\asqrt[50] ), .A3(new_n12888_), .A4(new_n13082_), .ZN(new_n13465_));
  XOR2_X1    g13273(.A1(new_n13465_), .A2(new_n13464_), .Z(new_n13466_));
  NAND2_X1   g13274(.A1(new_n13466_), .A2(new_n1436_), .ZN(new_n13467_));
  INV_X1     g13275(.I(new_n13467_), .ZN(new_n13468_));
  OAI21_X1   g13276(.A1(new_n13463_), .A2(new_n1595_), .B(new_n13468_), .ZN(new_n13469_));
  NAND2_X1   g13277(.A1(new_n13469_), .A2(new_n13462_), .ZN(new_n13470_));
  OAI22_X1   g13278(.A1(new_n13463_), .A2(new_n1595_), .B1(new_n13461_), .B2(new_n13455_), .ZN(new_n13471_));
  NAND2_X1   g13279(.A1(new_n12900_), .A2(\asqrt[51] ), .ZN(new_n13472_));
  NOR4_X1    g13280(.A1(new_n13192_), .A2(\asqrt[51] ), .A3(new_n12895_), .A4(new_n12900_), .ZN(new_n13473_));
  XOR2_X1    g13281(.A1(new_n13473_), .A2(new_n13472_), .Z(new_n13474_));
  NAND2_X1   g13282(.A1(new_n13474_), .A2(new_n1260_), .ZN(new_n13475_));
  AOI21_X1   g13283(.A1(new_n13471_), .A2(\asqrt[51] ), .B(new_n13475_), .ZN(new_n13476_));
  NOR2_X1    g13284(.A1(new_n13476_), .A2(new_n13470_), .ZN(new_n13477_));
  AOI22_X1   g13285(.A1(new_n13471_), .A2(\asqrt[51] ), .B1(new_n13469_), .B2(new_n13462_), .ZN(new_n13478_));
  NOR4_X1    g13286(.A1(new_n13192_), .A2(\asqrt[52] ), .A3(new_n12903_), .A4(new_n13089_), .ZN(new_n13479_));
  AOI21_X1   g13287(.A1(new_n13472_), .A2(new_n12899_), .B(new_n1260_), .ZN(new_n13480_));
  NOR2_X1    g13288(.A1(new_n13479_), .A2(new_n13480_), .ZN(new_n13481_));
  NAND2_X1   g13289(.A1(new_n13481_), .A2(new_n1096_), .ZN(new_n13482_));
  INV_X1     g13290(.I(new_n13482_), .ZN(new_n13483_));
  OAI21_X1   g13291(.A1(new_n13478_), .A2(new_n1260_), .B(new_n13483_), .ZN(new_n13484_));
  NAND2_X1   g13292(.A1(new_n13484_), .A2(new_n13477_), .ZN(new_n13485_));
  OAI22_X1   g13293(.A1(new_n13478_), .A2(new_n1260_), .B1(new_n13476_), .B2(new_n13470_), .ZN(new_n13486_));
  NAND2_X1   g13294(.A1(new_n12915_), .A2(\asqrt[53] ), .ZN(new_n13487_));
  NOR4_X1    g13295(.A1(new_n13192_), .A2(\asqrt[53] ), .A3(new_n12910_), .A4(new_n12915_), .ZN(new_n13488_));
  XOR2_X1    g13296(.A1(new_n13488_), .A2(new_n13487_), .Z(new_n13489_));
  NAND2_X1   g13297(.A1(new_n13489_), .A2(new_n970_), .ZN(new_n13490_));
  AOI21_X1   g13298(.A1(new_n13486_), .A2(\asqrt[53] ), .B(new_n13490_), .ZN(new_n13491_));
  NOR2_X1    g13299(.A1(new_n13491_), .A2(new_n13485_), .ZN(new_n13492_));
  AOI22_X1   g13300(.A1(new_n13486_), .A2(\asqrt[53] ), .B1(new_n13484_), .B2(new_n13477_), .ZN(new_n13493_));
  NOR4_X1    g13301(.A1(new_n13192_), .A2(\asqrt[54] ), .A3(new_n12917_), .A4(new_n13096_), .ZN(new_n13494_));
  AOI21_X1   g13302(.A1(new_n13487_), .A2(new_n12914_), .B(new_n970_), .ZN(new_n13495_));
  NOR2_X1    g13303(.A1(new_n13494_), .A2(new_n13495_), .ZN(new_n13496_));
  NAND2_X1   g13304(.A1(new_n13496_), .A2(new_n825_), .ZN(new_n13497_));
  INV_X1     g13305(.I(new_n13497_), .ZN(new_n13498_));
  OAI21_X1   g13306(.A1(new_n13493_), .A2(new_n970_), .B(new_n13498_), .ZN(new_n13499_));
  NAND2_X1   g13307(.A1(new_n13499_), .A2(new_n13492_), .ZN(new_n13500_));
  OAI22_X1   g13308(.A1(new_n13493_), .A2(new_n970_), .B1(new_n13491_), .B2(new_n13485_), .ZN(new_n13501_));
  NAND2_X1   g13309(.A1(new_n12928_), .A2(\asqrt[55] ), .ZN(new_n13502_));
  NOR4_X1    g13310(.A1(new_n13192_), .A2(\asqrt[55] ), .A3(new_n12923_), .A4(new_n12928_), .ZN(new_n13503_));
  XOR2_X1    g13311(.A1(new_n13503_), .A2(new_n13502_), .Z(new_n13504_));
  NAND2_X1   g13312(.A1(new_n13504_), .A2(new_n724_), .ZN(new_n13505_));
  AOI21_X1   g13313(.A1(new_n13501_), .A2(\asqrt[55] ), .B(new_n13505_), .ZN(new_n13506_));
  NOR2_X1    g13314(.A1(new_n13506_), .A2(new_n13500_), .ZN(new_n13507_));
  AOI22_X1   g13315(.A1(new_n13501_), .A2(\asqrt[55] ), .B1(new_n13499_), .B2(new_n13492_), .ZN(new_n13508_));
  NOR4_X1    g13316(.A1(new_n13192_), .A2(\asqrt[56] ), .A3(new_n12930_), .A4(new_n13103_), .ZN(new_n13509_));
  AOI21_X1   g13317(.A1(new_n13502_), .A2(new_n12927_), .B(new_n724_), .ZN(new_n13510_));
  NOR2_X1    g13318(.A1(new_n13509_), .A2(new_n13510_), .ZN(new_n13511_));
  NAND2_X1   g13319(.A1(new_n13511_), .A2(new_n587_), .ZN(new_n13512_));
  INV_X1     g13320(.I(new_n13512_), .ZN(new_n13513_));
  OAI21_X1   g13321(.A1(new_n13508_), .A2(new_n724_), .B(new_n13513_), .ZN(new_n13514_));
  NAND2_X1   g13322(.A1(new_n13514_), .A2(new_n13507_), .ZN(new_n13515_));
  OAI22_X1   g13323(.A1(new_n13216_), .A2(new_n11631_), .B1(new_n13204_), .B2(new_n13214_), .ZN(new_n13516_));
  AOI22_X1   g13324(.A1(new_n13516_), .A2(\asqrt[22] ), .B1(new_n13223_), .B2(new_n13215_), .ZN(new_n13517_));
  INV_X1     g13325(.I(new_n13257_), .ZN(new_n13518_));
  OAI21_X1   g13326(.A1(new_n13517_), .A2(new_n10614_), .B(new_n13518_), .ZN(new_n13519_));
  AOI21_X1   g13327(.A1(new_n13516_), .A2(\asqrt[22] ), .B(new_n13231_), .ZN(new_n13520_));
  OAI22_X1   g13328(.A1(new_n13517_), .A2(new_n10614_), .B1(new_n13520_), .B2(new_n13260_), .ZN(new_n13521_));
  AOI22_X1   g13329(.A1(new_n13521_), .A2(\asqrt[24] ), .B1(new_n13519_), .B2(new_n13261_), .ZN(new_n13522_));
  INV_X1     g13330(.I(new_n13276_), .ZN(new_n13523_));
  OAI21_X1   g13331(.A1(new_n13522_), .A2(new_n9672_), .B(new_n13523_), .ZN(new_n13524_));
  NAND2_X1   g13332(.A1(new_n13524_), .A2(new_n13280_), .ZN(new_n13525_));
  AOI21_X1   g13333(.A1(new_n13521_), .A2(\asqrt[24] ), .B(new_n13267_), .ZN(new_n13526_));
  OAI22_X1   g13334(.A1(new_n13522_), .A2(new_n9672_), .B1(new_n13526_), .B2(new_n13279_), .ZN(new_n13527_));
  AOI21_X1   g13335(.A1(new_n13527_), .A2(\asqrt[26] ), .B(new_n13286_), .ZN(new_n13528_));
  NOR2_X1    g13336(.A1(new_n13528_), .A2(new_n13525_), .ZN(new_n13529_));
  AOI22_X1   g13337(.A1(new_n13527_), .A2(\asqrt[26] ), .B1(new_n13524_), .B2(new_n13280_), .ZN(new_n13530_));
  INV_X1     g13338(.I(new_n13295_), .ZN(new_n13531_));
  OAI21_X1   g13339(.A1(new_n13530_), .A2(new_n8763_), .B(new_n13531_), .ZN(new_n13532_));
  NAND2_X1   g13340(.A1(new_n13532_), .A2(new_n13529_), .ZN(new_n13533_));
  OAI22_X1   g13341(.A1(new_n13530_), .A2(new_n8763_), .B1(new_n13528_), .B2(new_n13525_), .ZN(new_n13534_));
  AOI21_X1   g13342(.A1(new_n13534_), .A2(\asqrt[28] ), .B(new_n13302_), .ZN(new_n13535_));
  NOR2_X1    g13343(.A1(new_n13535_), .A2(new_n13533_), .ZN(new_n13536_));
  AOI22_X1   g13344(.A1(new_n13534_), .A2(\asqrt[28] ), .B1(new_n13532_), .B2(new_n13529_), .ZN(new_n13537_));
  INV_X1     g13345(.I(new_n13310_), .ZN(new_n13538_));
  OAI21_X1   g13346(.A1(new_n13537_), .A2(new_n7931_), .B(new_n13538_), .ZN(new_n13539_));
  NAND2_X1   g13347(.A1(new_n13539_), .A2(new_n13536_), .ZN(new_n13540_));
  OAI22_X1   g13348(.A1(new_n13537_), .A2(new_n7931_), .B1(new_n13535_), .B2(new_n13533_), .ZN(new_n13541_));
  AOI21_X1   g13349(.A1(new_n13541_), .A2(\asqrt[30] ), .B(new_n13317_), .ZN(new_n13542_));
  NOR2_X1    g13350(.A1(new_n13542_), .A2(new_n13540_), .ZN(new_n13543_));
  AOI22_X1   g13351(.A1(new_n13541_), .A2(\asqrt[30] ), .B1(new_n13539_), .B2(new_n13536_), .ZN(new_n13544_));
  INV_X1     g13352(.I(new_n13325_), .ZN(new_n13545_));
  OAI21_X1   g13353(.A1(new_n13544_), .A2(new_n7110_), .B(new_n13545_), .ZN(new_n13546_));
  NAND2_X1   g13354(.A1(new_n13546_), .A2(new_n13543_), .ZN(new_n13547_));
  OAI22_X1   g13355(.A1(new_n13544_), .A2(new_n7110_), .B1(new_n13542_), .B2(new_n13540_), .ZN(new_n13548_));
  AOI21_X1   g13356(.A1(new_n13548_), .A2(\asqrt[32] ), .B(new_n13332_), .ZN(new_n13549_));
  NOR2_X1    g13357(.A1(new_n13549_), .A2(new_n13547_), .ZN(new_n13550_));
  AOI22_X1   g13358(.A1(new_n13548_), .A2(\asqrt[32] ), .B1(new_n13546_), .B2(new_n13543_), .ZN(new_n13551_));
  INV_X1     g13359(.I(new_n13340_), .ZN(new_n13552_));
  OAI21_X1   g13360(.A1(new_n13551_), .A2(new_n6365_), .B(new_n13552_), .ZN(new_n13553_));
  NAND2_X1   g13361(.A1(new_n13553_), .A2(new_n13550_), .ZN(new_n13554_));
  OAI22_X1   g13362(.A1(new_n13551_), .A2(new_n6365_), .B1(new_n13549_), .B2(new_n13547_), .ZN(new_n13555_));
  AOI21_X1   g13363(.A1(new_n13555_), .A2(\asqrt[34] ), .B(new_n13347_), .ZN(new_n13556_));
  NOR2_X1    g13364(.A1(new_n13556_), .A2(new_n13554_), .ZN(new_n13557_));
  AOI22_X1   g13365(.A1(new_n13555_), .A2(\asqrt[34] ), .B1(new_n13553_), .B2(new_n13550_), .ZN(new_n13558_));
  INV_X1     g13366(.I(new_n13355_), .ZN(new_n13559_));
  OAI21_X1   g13367(.A1(new_n13558_), .A2(new_n5626_), .B(new_n13559_), .ZN(new_n13560_));
  NAND2_X1   g13368(.A1(new_n13560_), .A2(new_n13557_), .ZN(new_n13561_));
  OAI22_X1   g13369(.A1(new_n13558_), .A2(new_n5626_), .B1(new_n13556_), .B2(new_n13554_), .ZN(new_n13562_));
  AOI21_X1   g13370(.A1(new_n13562_), .A2(\asqrt[36] ), .B(new_n13362_), .ZN(new_n13563_));
  NOR2_X1    g13371(.A1(new_n13563_), .A2(new_n13561_), .ZN(new_n13564_));
  AOI22_X1   g13372(.A1(new_n13562_), .A2(\asqrt[36] ), .B1(new_n13560_), .B2(new_n13557_), .ZN(new_n13565_));
  INV_X1     g13373(.I(new_n13370_), .ZN(new_n13566_));
  OAI21_X1   g13374(.A1(new_n13565_), .A2(new_n4973_), .B(new_n13566_), .ZN(new_n13567_));
  NAND2_X1   g13375(.A1(new_n13567_), .A2(new_n13564_), .ZN(new_n13568_));
  OAI22_X1   g13376(.A1(new_n13565_), .A2(new_n4973_), .B1(new_n13563_), .B2(new_n13561_), .ZN(new_n13569_));
  AOI21_X1   g13377(.A1(new_n13569_), .A2(\asqrt[38] ), .B(new_n13377_), .ZN(new_n13570_));
  NOR2_X1    g13378(.A1(new_n13570_), .A2(new_n13568_), .ZN(new_n13571_));
  AOI22_X1   g13379(.A1(new_n13569_), .A2(\asqrt[38] ), .B1(new_n13567_), .B2(new_n13564_), .ZN(new_n13572_));
  INV_X1     g13380(.I(new_n13385_), .ZN(new_n13573_));
  OAI21_X1   g13381(.A1(new_n13572_), .A2(new_n4330_), .B(new_n13573_), .ZN(new_n13574_));
  NAND2_X1   g13382(.A1(new_n13574_), .A2(new_n13571_), .ZN(new_n13575_));
  OAI22_X1   g13383(.A1(new_n13572_), .A2(new_n4330_), .B1(new_n13570_), .B2(new_n13568_), .ZN(new_n13576_));
  AOI21_X1   g13384(.A1(new_n13576_), .A2(\asqrt[40] ), .B(new_n13392_), .ZN(new_n13577_));
  NOR2_X1    g13385(.A1(new_n13577_), .A2(new_n13575_), .ZN(new_n13578_));
  AOI22_X1   g13386(.A1(new_n13576_), .A2(\asqrt[40] ), .B1(new_n13574_), .B2(new_n13571_), .ZN(new_n13579_));
  INV_X1     g13387(.I(new_n13400_), .ZN(new_n13580_));
  OAI21_X1   g13388(.A1(new_n13579_), .A2(new_n3760_), .B(new_n13580_), .ZN(new_n13581_));
  NAND2_X1   g13389(.A1(new_n13581_), .A2(new_n13578_), .ZN(new_n13582_));
  OAI22_X1   g13390(.A1(new_n13579_), .A2(new_n3760_), .B1(new_n13577_), .B2(new_n13575_), .ZN(new_n13583_));
  AOI21_X1   g13391(.A1(new_n13583_), .A2(\asqrt[42] ), .B(new_n13407_), .ZN(new_n13584_));
  NOR2_X1    g13392(.A1(new_n13584_), .A2(new_n13582_), .ZN(new_n13585_));
  AOI22_X1   g13393(.A1(new_n13583_), .A2(\asqrt[42] ), .B1(new_n13581_), .B2(new_n13578_), .ZN(new_n13586_));
  INV_X1     g13394(.I(new_n13415_), .ZN(new_n13587_));
  OAI21_X1   g13395(.A1(new_n13586_), .A2(new_n3208_), .B(new_n13587_), .ZN(new_n13588_));
  NAND2_X1   g13396(.A1(new_n13588_), .A2(new_n13585_), .ZN(new_n13589_));
  OAI22_X1   g13397(.A1(new_n13586_), .A2(new_n3208_), .B1(new_n13584_), .B2(new_n13582_), .ZN(new_n13590_));
  AOI21_X1   g13398(.A1(new_n13590_), .A2(\asqrt[44] ), .B(new_n13422_), .ZN(new_n13591_));
  NOR2_X1    g13399(.A1(new_n13591_), .A2(new_n13589_), .ZN(new_n13592_));
  AOI22_X1   g13400(.A1(new_n13590_), .A2(\asqrt[44] ), .B1(new_n13588_), .B2(new_n13585_), .ZN(new_n13593_));
  INV_X1     g13401(.I(new_n13430_), .ZN(new_n13594_));
  OAI21_X1   g13402(.A1(new_n13593_), .A2(new_n2728_), .B(new_n13594_), .ZN(new_n13595_));
  NAND2_X1   g13403(.A1(new_n13595_), .A2(new_n13592_), .ZN(new_n13596_));
  OAI22_X1   g13404(.A1(new_n13593_), .A2(new_n2728_), .B1(new_n13591_), .B2(new_n13589_), .ZN(new_n13597_));
  AOI21_X1   g13405(.A1(new_n13597_), .A2(\asqrt[46] ), .B(new_n13437_), .ZN(new_n13598_));
  NOR2_X1    g13406(.A1(new_n13598_), .A2(new_n13596_), .ZN(new_n13599_));
  AOI22_X1   g13407(.A1(new_n13597_), .A2(\asqrt[46] ), .B1(new_n13595_), .B2(new_n13592_), .ZN(new_n13600_));
  INV_X1     g13408(.I(new_n13445_), .ZN(new_n13601_));
  OAI21_X1   g13409(.A1(new_n13600_), .A2(new_n2253_), .B(new_n13601_), .ZN(new_n13602_));
  NAND2_X1   g13410(.A1(new_n13602_), .A2(new_n13599_), .ZN(new_n13603_));
  OAI22_X1   g13411(.A1(new_n13600_), .A2(new_n2253_), .B1(new_n13598_), .B2(new_n13596_), .ZN(new_n13604_));
  AOI21_X1   g13412(.A1(new_n13604_), .A2(\asqrt[48] ), .B(new_n13452_), .ZN(new_n13605_));
  NOR2_X1    g13413(.A1(new_n13605_), .A2(new_n13603_), .ZN(new_n13606_));
  AOI22_X1   g13414(.A1(new_n13604_), .A2(\asqrt[48] ), .B1(new_n13602_), .B2(new_n13599_), .ZN(new_n13607_));
  INV_X1     g13415(.I(new_n13460_), .ZN(new_n13608_));
  OAI21_X1   g13416(.A1(new_n13607_), .A2(new_n1854_), .B(new_n13608_), .ZN(new_n13609_));
  NAND2_X1   g13417(.A1(new_n13609_), .A2(new_n13606_), .ZN(new_n13610_));
  OAI22_X1   g13418(.A1(new_n13607_), .A2(new_n1854_), .B1(new_n13605_), .B2(new_n13603_), .ZN(new_n13611_));
  AOI21_X1   g13419(.A1(new_n13611_), .A2(\asqrt[50] ), .B(new_n13467_), .ZN(new_n13612_));
  NOR2_X1    g13420(.A1(new_n13612_), .A2(new_n13610_), .ZN(new_n13613_));
  AOI22_X1   g13421(.A1(new_n13611_), .A2(\asqrt[50] ), .B1(new_n13609_), .B2(new_n13606_), .ZN(new_n13614_));
  INV_X1     g13422(.I(new_n13475_), .ZN(new_n13615_));
  OAI21_X1   g13423(.A1(new_n13614_), .A2(new_n1436_), .B(new_n13615_), .ZN(new_n13616_));
  NAND2_X1   g13424(.A1(new_n13616_), .A2(new_n13613_), .ZN(new_n13617_));
  OAI22_X1   g13425(.A1(new_n13614_), .A2(new_n1436_), .B1(new_n13612_), .B2(new_n13610_), .ZN(new_n13618_));
  AOI21_X1   g13426(.A1(new_n13618_), .A2(\asqrt[52] ), .B(new_n13482_), .ZN(new_n13619_));
  NOR2_X1    g13427(.A1(new_n13619_), .A2(new_n13617_), .ZN(new_n13620_));
  AOI22_X1   g13428(.A1(new_n13618_), .A2(\asqrt[52] ), .B1(new_n13616_), .B2(new_n13613_), .ZN(new_n13621_));
  INV_X1     g13429(.I(new_n13490_), .ZN(new_n13622_));
  OAI21_X1   g13430(.A1(new_n13621_), .A2(new_n1096_), .B(new_n13622_), .ZN(new_n13623_));
  NAND2_X1   g13431(.A1(new_n13623_), .A2(new_n13620_), .ZN(new_n13624_));
  OAI22_X1   g13432(.A1(new_n13621_), .A2(new_n1096_), .B1(new_n13619_), .B2(new_n13617_), .ZN(new_n13625_));
  AOI21_X1   g13433(.A1(new_n13625_), .A2(\asqrt[54] ), .B(new_n13497_), .ZN(new_n13626_));
  NOR2_X1    g13434(.A1(new_n13626_), .A2(new_n13624_), .ZN(new_n13627_));
  NAND2_X1   g13435(.A1(new_n13618_), .A2(\asqrt[52] ), .ZN(new_n13628_));
  AOI21_X1   g13436(.A1(new_n13628_), .A2(new_n13617_), .B(new_n1096_), .ZN(new_n13629_));
  OAI21_X1   g13437(.A1(new_n13620_), .A2(new_n13629_), .B(\asqrt[54] ), .ZN(new_n13630_));
  AOI21_X1   g13438(.A1(new_n13624_), .A2(new_n13630_), .B(new_n825_), .ZN(new_n13631_));
  OAI21_X1   g13439(.A1(new_n13627_), .A2(new_n13631_), .B(\asqrt[56] ), .ZN(new_n13632_));
  INV_X1     g13440(.I(new_n13632_), .ZN(new_n13633_));
  OAI21_X1   g13441(.A1(new_n13633_), .A2(new_n13507_), .B(\asqrt[57] ), .ZN(new_n13634_));
  NOR4_X1    g13442(.A1(new_n13192_), .A2(\asqrt[57] ), .A3(new_n12936_), .A4(new_n12941_), .ZN(new_n13635_));
  XOR2_X1    g13443(.A1(new_n13635_), .A2(new_n13132_), .Z(new_n13636_));
  AND2_X2    g13444(.A1(new_n13636_), .A2(new_n504_), .Z(new_n13637_));
  AOI21_X1   g13445(.A1(new_n13634_), .A2(new_n13637_), .B(new_n13515_), .ZN(new_n13638_));
  OAI22_X1   g13446(.A1(new_n13508_), .A2(new_n724_), .B1(new_n13506_), .B2(new_n13500_), .ZN(new_n13639_));
  AOI22_X1   g13447(.A1(new_n13639_), .A2(\asqrt[57] ), .B1(new_n13514_), .B2(new_n13507_), .ZN(new_n13640_));
  NOR4_X1    g13448(.A1(new_n13192_), .A2(\asqrt[58] ), .A3(new_n12943_), .A4(new_n13110_), .ZN(new_n13641_));
  XOR2_X1    g13449(.A1(new_n13641_), .A2(new_n13156_), .Z(new_n13642_));
  NAND2_X1   g13450(.A1(new_n13642_), .A2(new_n376_), .ZN(new_n13643_));
  INV_X1     g13451(.I(new_n13643_), .ZN(new_n13644_));
  OAI21_X1   g13452(.A1(new_n13640_), .A2(new_n504_), .B(new_n13644_), .ZN(new_n13645_));
  NAND2_X1   g13453(.A1(new_n13645_), .A2(new_n13638_), .ZN(new_n13646_));
  AOI21_X1   g13454(.A1(new_n13634_), .A2(new_n13515_), .B(new_n504_), .ZN(new_n13647_));
  OAI21_X1   g13455(.A1(new_n13638_), .A2(new_n13647_), .B(\asqrt[59] ), .ZN(new_n13648_));
  NOR4_X1    g13456(.A1(new_n13192_), .A2(\asqrt[59] ), .A3(new_n12949_), .A4(new_n12954_), .ZN(new_n13649_));
  XOR2_X1    g13457(.A1(new_n13649_), .A2(new_n13134_), .Z(new_n13650_));
  AND2_X2    g13458(.A1(new_n13650_), .A2(new_n275_), .Z(new_n13651_));
  AOI21_X1   g13459(.A1(new_n13648_), .A2(new_n13651_), .B(new_n13646_), .ZN(new_n13652_));
  AOI22_X1   g13460(.A1(new_n13625_), .A2(\asqrt[54] ), .B1(new_n13623_), .B2(new_n13620_), .ZN(new_n13653_));
  INV_X1     g13461(.I(new_n13505_), .ZN(new_n13654_));
  OAI21_X1   g13462(.A1(new_n13653_), .A2(new_n825_), .B(new_n13654_), .ZN(new_n13655_));
  NAND2_X1   g13463(.A1(new_n13655_), .A2(new_n13627_), .ZN(new_n13656_));
  OAI22_X1   g13464(.A1(new_n13653_), .A2(new_n825_), .B1(new_n13626_), .B2(new_n13624_), .ZN(new_n13657_));
  AOI21_X1   g13465(.A1(new_n13657_), .A2(\asqrt[56] ), .B(new_n13512_), .ZN(new_n13658_));
  NOR2_X1    g13466(.A1(new_n13658_), .A2(new_n13656_), .ZN(new_n13659_));
  AOI22_X1   g13467(.A1(new_n13657_), .A2(\asqrt[56] ), .B1(new_n13655_), .B2(new_n13627_), .ZN(new_n13660_));
  OAI21_X1   g13468(.A1(new_n13660_), .A2(new_n587_), .B(new_n13637_), .ZN(new_n13661_));
  NAND2_X1   g13469(.A1(new_n13661_), .A2(new_n13659_), .ZN(new_n13662_));
  AOI21_X1   g13470(.A1(new_n13656_), .A2(new_n13632_), .B(new_n587_), .ZN(new_n13663_));
  OAI21_X1   g13471(.A1(new_n13659_), .A2(new_n13663_), .B(\asqrt[58] ), .ZN(new_n13664_));
  NAND2_X1   g13472(.A1(new_n13662_), .A2(new_n13664_), .ZN(new_n13665_));
  AOI22_X1   g13473(.A1(new_n13665_), .A2(\asqrt[59] ), .B1(new_n13645_), .B2(new_n13638_), .ZN(new_n13666_));
  NOR4_X1    g13474(.A1(new_n13192_), .A2(\asqrt[60] ), .A3(new_n12956_), .A4(new_n13117_), .ZN(new_n13667_));
  XOR2_X1    g13475(.A1(new_n13667_), .A2(new_n13158_), .Z(new_n13668_));
  NAND2_X1   g13476(.A1(new_n13668_), .A2(new_n229_), .ZN(new_n13669_));
  INV_X1     g13477(.I(new_n13669_), .ZN(new_n13670_));
  OAI21_X1   g13478(.A1(new_n13666_), .A2(new_n275_), .B(new_n13670_), .ZN(new_n13671_));
  OAI22_X1   g13479(.A1(new_n13660_), .A2(new_n587_), .B1(new_n13658_), .B2(new_n13656_), .ZN(new_n13672_));
  AOI21_X1   g13480(.A1(new_n13672_), .A2(\asqrt[58] ), .B(new_n13643_), .ZN(new_n13673_));
  NOR2_X1    g13481(.A1(new_n13673_), .A2(new_n13662_), .ZN(new_n13674_));
  AOI22_X1   g13482(.A1(new_n13672_), .A2(\asqrt[58] ), .B1(new_n13661_), .B2(new_n13659_), .ZN(new_n13675_));
  OAI21_X1   g13483(.A1(new_n13675_), .A2(new_n376_), .B(new_n13651_), .ZN(new_n13676_));
  NAND2_X1   g13484(.A1(new_n13676_), .A2(new_n13674_), .ZN(new_n13677_));
  AOI21_X1   g13485(.A1(new_n13662_), .A2(new_n13664_), .B(new_n376_), .ZN(new_n13678_));
  OAI21_X1   g13486(.A1(new_n13674_), .A2(new_n13678_), .B(\asqrt[60] ), .ZN(new_n13679_));
  AOI21_X1   g13487(.A1(new_n13677_), .A2(new_n13679_), .B(new_n229_), .ZN(new_n13680_));
  INV_X1     g13488(.I(new_n13162_), .ZN(new_n13681_));
  NOR2_X1    g13489(.A1(new_n13681_), .A2(\asqrt[62] ), .ZN(new_n13682_));
  INV_X1     g13490(.I(new_n13682_), .ZN(new_n13683_));
  NAND4_X1   g13491(.A1(new_n13680_), .A2(new_n13652_), .A3(new_n13671_), .A4(new_n13683_), .ZN(new_n13684_));
  NAND3_X1   g13492(.A1(new_n13192_), .A2(new_n13128_), .A3(new_n13180_), .ZN(new_n13685_));
  AOI21_X1   g13493(.A1(new_n13685_), .A2(new_n13140_), .B(\asqrt[63] ), .ZN(new_n13686_));
  NAND3_X1   g13494(.A1(new_n13684_), .A2(new_n13164_), .A3(new_n13686_), .ZN(new_n13687_));
  OAI22_X1   g13495(.A1(new_n13675_), .A2(new_n376_), .B1(new_n13673_), .B2(new_n13662_), .ZN(new_n13688_));
  AOI21_X1   g13496(.A1(new_n13688_), .A2(\asqrt[60] ), .B(new_n13669_), .ZN(new_n13689_));
  AOI22_X1   g13497(.A1(new_n13688_), .A2(\asqrt[60] ), .B1(new_n13676_), .B2(new_n13674_), .ZN(new_n13690_));
  OAI22_X1   g13498(.A1(new_n13690_), .A2(new_n229_), .B1(new_n13689_), .B2(new_n13677_), .ZN(new_n13691_));
  NOR4_X1    g13499(.A1(new_n13691_), .A2(\asqrt[62] ), .A3(new_n13154_), .A4(new_n13162_), .ZN(new_n13692_));
  AOI21_X1   g13500(.A1(new_n13155_), .A2(new_n13687_), .B(new_n13692_), .ZN(new_n13693_));
  INV_X1     g13501(.I(\a[32] ), .ZN(new_n13694_));
  OAI21_X1   g13502(.A1(new_n13129_), .A2(new_n13140_), .B(\asqrt[18] ), .ZN(new_n13695_));
  XOR2_X1    g13503(.A1(new_n13140_), .A2(\asqrt[63] ), .Z(new_n13696_));
  NAND2_X1   g13504(.A1(new_n13695_), .A2(new_n13696_), .ZN(new_n13697_));
  INV_X1     g13505(.I(new_n13697_), .ZN(new_n13698_));
  NAND3_X1   g13506(.A1(new_n13186_), .A2(new_n13122_), .A3(new_n13129_), .ZN(new_n13699_));
  INV_X1     g13507(.I(new_n13699_), .ZN(new_n13700_));
  NOR2_X1    g13508(.A1(new_n13698_), .A2(new_n13700_), .ZN(new_n13701_));
  NOR2_X1    g13509(.A1(\a[30] ), .A2(\a[31] ), .ZN(new_n13702_));
  INV_X1     g13510(.I(new_n13702_), .ZN(new_n13703_));
  NOR3_X1    g13511(.A1(new_n13701_), .A2(new_n13694_), .A3(new_n13703_), .ZN(new_n13704_));
  NAND2_X1   g13512(.A1(new_n13693_), .A2(new_n13704_), .ZN(new_n13705_));
  XOR2_X1    g13513(.A1(new_n13705_), .A2(\a[33] ), .Z(new_n13706_));
  INV_X1     g13514(.I(\a[33] ), .ZN(new_n13707_));
  NAND2_X1   g13515(.A1(new_n13671_), .A2(new_n13652_), .ZN(new_n13708_));
  NAND2_X1   g13516(.A1(new_n13680_), .A2(new_n13683_), .ZN(new_n13709_));
  OAI21_X1   g13517(.A1(new_n13709_), .A2(new_n13708_), .B(new_n13164_), .ZN(new_n13710_));
  INV_X1     g13518(.I(new_n13686_), .ZN(new_n13711_));
  OAI21_X1   g13519(.A1(new_n13710_), .A2(new_n13711_), .B(new_n13155_), .ZN(new_n13712_));
  NAND2_X1   g13520(.A1(new_n13692_), .A2(new_n13698_), .ZN(new_n13713_));
  NOR2_X1    g13521(.A1(new_n13713_), .A2(new_n13712_), .ZN(new_n13714_));
  NAND3_X1   g13522(.A1(new_n13714_), .A2(new_n13155_), .A3(new_n13699_), .ZN(new_n13715_));
  NAND2_X1   g13523(.A1(new_n13677_), .A2(new_n13679_), .ZN(new_n13716_));
  AOI22_X1   g13524(.A1(new_n13716_), .A2(\asqrt[61] ), .B1(new_n13671_), .B2(new_n13652_), .ZN(new_n13717_));
  NOR2_X1    g13525(.A1(new_n13717_), .A2(new_n196_), .ZN(new_n13718_));
  AOI21_X1   g13526(.A1(new_n13646_), .A2(new_n13648_), .B(new_n275_), .ZN(new_n13719_));
  OAI21_X1   g13527(.A1(new_n13652_), .A2(new_n13719_), .B(\asqrt[61] ), .ZN(new_n13720_));
  NAND4_X1   g13528(.A1(new_n13708_), .A2(new_n196_), .A3(new_n13720_), .A4(new_n13681_), .ZN(new_n13721_));
  INV_X1     g13529(.I(new_n13721_), .ZN(new_n13722_));
  NOR3_X1    g13530(.A1(new_n13713_), .A2(new_n13712_), .A3(new_n13699_), .ZN(\asqrt[17] ));
  NAND3_X1   g13531(.A1(\asqrt[17] ), .A2(new_n13718_), .A3(new_n13722_), .ZN(new_n13724_));
  OAI21_X1   g13532(.A1(new_n13691_), .A2(\asqrt[62] ), .B(new_n13162_), .ZN(new_n13725_));
  OAI21_X1   g13533(.A1(\asqrt[17] ), .A2(new_n13725_), .B(new_n13718_), .ZN(new_n13726_));
  NAND2_X1   g13534(.A1(new_n13726_), .A2(new_n13724_), .ZN(new_n13727_));
  INV_X1     g13535(.I(new_n13727_), .ZN(new_n13728_));
  NOR3_X1    g13536(.A1(new_n13716_), .A2(\asqrt[61] ), .A3(new_n13668_), .ZN(new_n13729_));
  NAND2_X1   g13537(.A1(\asqrt[17] ), .A2(new_n13729_), .ZN(new_n13730_));
  XOR2_X1    g13538(.A1(new_n13730_), .A2(new_n13680_), .Z(new_n13731_));
  NOR2_X1    g13539(.A1(new_n13731_), .A2(new_n196_), .ZN(new_n13732_));
  INV_X1     g13540(.I(new_n13732_), .ZN(new_n13733_));
  INV_X1     g13541(.I(\a[34] ), .ZN(new_n13734_));
  NOR2_X1    g13542(.A1(\a[32] ), .A2(\a[33] ), .ZN(new_n13735_));
  INV_X1     g13543(.I(new_n13735_), .ZN(new_n13736_));
  NOR2_X1    g13544(.A1(new_n13736_), .A2(new_n13734_), .ZN(new_n13737_));
  NAND4_X1   g13545(.A1(new_n13144_), .A2(new_n13180_), .A3(new_n13194_), .A4(new_n13737_), .ZN(new_n13738_));
  XOR2_X1    g13546(.A1(new_n13738_), .A2(\a[35] ), .Z(new_n13739_));
  INV_X1     g13547(.I(\a[35] ), .ZN(new_n13740_));
  NOR4_X1    g13548(.A1(new_n13713_), .A2(new_n13712_), .A3(new_n13740_), .A4(new_n13699_), .ZN(new_n13741_));
  NOR2_X1    g13549(.A1(new_n13739_), .A2(\a[34] ), .ZN(new_n13742_));
  OAI21_X1   g13550(.A1(new_n13741_), .A2(new_n13742_), .B(new_n13739_), .ZN(new_n13743_));
  INV_X1     g13551(.I(new_n13739_), .ZN(new_n13744_));
  NOR2_X1    g13552(.A1(new_n13689_), .A2(new_n13677_), .ZN(new_n13745_));
  NOR3_X1    g13553(.A1(new_n13690_), .A2(new_n229_), .A3(new_n13682_), .ZN(new_n13746_));
  AOI21_X1   g13554(.A1(new_n13746_), .A2(new_n13745_), .B(new_n13163_), .ZN(new_n13747_));
  AOI21_X1   g13555(.A1(new_n13747_), .A2(new_n13686_), .B(new_n13154_), .ZN(new_n13748_));
  AOI21_X1   g13556(.A1(new_n13691_), .A2(\asqrt[62] ), .B(new_n13155_), .ZN(new_n13749_));
  NOR3_X1    g13557(.A1(new_n13749_), .A2(new_n13721_), .A3(new_n13697_), .ZN(new_n13750_));
  NAND4_X1   g13558(.A1(new_n13750_), .A2(\a[35] ), .A3(new_n13748_), .A4(new_n13700_), .ZN(new_n13751_));
  NAND3_X1   g13559(.A1(new_n13751_), .A2(\a[34] ), .A3(new_n13744_), .ZN(new_n13752_));
  NAND2_X1   g13560(.A1(new_n13743_), .A2(new_n13752_), .ZN(new_n13753_));
  NAND2_X1   g13561(.A1(new_n13178_), .A2(new_n13142_), .ZN(new_n13754_));
  NAND4_X1   g13562(.A1(new_n13182_), .A2(new_n13176_), .A3(new_n13129_), .A4(new_n13754_), .ZN(new_n13755_));
  NOR2_X1    g13563(.A1(new_n13192_), .A2(new_n13734_), .ZN(new_n13756_));
  XOR2_X1    g13564(.A1(new_n13756_), .A2(new_n13755_), .Z(new_n13757_));
  NOR2_X1    g13565(.A1(new_n13757_), .A2(new_n13736_), .ZN(new_n13758_));
  INV_X1     g13566(.I(new_n13758_), .ZN(new_n13759_));
  NAND3_X1   g13567(.A1(new_n13750_), .A2(new_n13748_), .A3(new_n13700_), .ZN(new_n13760_));
  NOR4_X1    g13568(.A1(new_n13720_), .A2(new_n13677_), .A3(new_n13689_), .A4(new_n13682_), .ZN(new_n13761_));
  NOR3_X1    g13569(.A1(new_n13761_), .A2(new_n13163_), .A3(new_n13711_), .ZN(new_n13762_));
  NAND4_X1   g13570(.A1(new_n13717_), .A2(new_n196_), .A3(new_n13155_), .A4(new_n13681_), .ZN(new_n13763_));
  OAI21_X1   g13571(.A1(new_n13762_), .A2(new_n13154_), .B(new_n13763_), .ZN(new_n13764_));
  NAND2_X1   g13572(.A1(new_n13701_), .A2(\asqrt[18] ), .ZN(new_n13765_));
  OAI21_X1   g13573(.A1(new_n13764_), .A2(new_n13765_), .B(new_n13165_), .ZN(new_n13766_));
  NAND3_X1   g13574(.A1(new_n13766_), .A2(new_n13166_), .A3(new_n13760_), .ZN(new_n13767_));
  INV_X1     g13575(.I(new_n13765_), .ZN(new_n13768_));
  AOI21_X1   g13576(.A1(new_n13693_), .A2(new_n13768_), .B(\a[36] ), .ZN(new_n13769_));
  OAI21_X1   g13577(.A1(new_n13769_), .A2(new_n13167_), .B(\asqrt[17] ), .ZN(new_n13770_));
  NAND4_X1   g13578(.A1(new_n13767_), .A2(new_n13770_), .A3(new_n12657_), .A4(new_n13759_), .ZN(new_n13771_));
  NAND2_X1   g13579(.A1(new_n13771_), .A2(new_n13753_), .ZN(new_n13772_));
  NAND3_X1   g13580(.A1(new_n13743_), .A2(new_n13752_), .A3(new_n13759_), .ZN(new_n13773_));
  AOI21_X1   g13581(.A1(\asqrt[18] ), .A2(new_n13165_), .B(\a[37] ), .ZN(new_n13774_));
  NOR2_X1    g13582(.A1(new_n13183_), .A2(\a[36] ), .ZN(new_n13775_));
  AOI21_X1   g13583(.A1(\asqrt[18] ), .A2(\a[36] ), .B(new_n13169_), .ZN(new_n13776_));
  OAI21_X1   g13584(.A1(new_n13775_), .A2(new_n13774_), .B(new_n13776_), .ZN(new_n13777_));
  INV_X1     g13585(.I(new_n13777_), .ZN(new_n13778_));
  NAND3_X1   g13586(.A1(\asqrt[17] ), .A2(new_n13191_), .A3(new_n13778_), .ZN(new_n13779_));
  OAI21_X1   g13587(.A1(new_n13760_), .A2(new_n13777_), .B(new_n13190_), .ZN(new_n13780_));
  NAND3_X1   g13588(.A1(new_n13779_), .A2(new_n13780_), .A3(new_n12101_), .ZN(new_n13781_));
  AOI21_X1   g13589(.A1(new_n13773_), .A2(\asqrt[19] ), .B(new_n13781_), .ZN(new_n13782_));
  NOR2_X1    g13590(.A1(new_n13772_), .A2(new_n13782_), .ZN(new_n13783_));
  AOI22_X1   g13591(.A1(new_n13771_), .A2(new_n13753_), .B1(\asqrt[19] ), .B2(new_n13773_), .ZN(new_n13784_));
  AOI21_X1   g13592(.A1(new_n13202_), .A2(new_n13198_), .B(\asqrt[20] ), .ZN(new_n13785_));
  AND4_X2    g13593(.A1(new_n13243_), .A2(\asqrt[17] ), .A3(new_n13224_), .A4(new_n13785_), .Z(new_n13786_));
  NOR2_X1    g13594(.A1(new_n13243_), .A2(new_n12101_), .ZN(new_n13787_));
  NOR3_X1    g13595(.A1(new_n13786_), .A2(\asqrt[21] ), .A3(new_n13787_), .ZN(new_n13788_));
  OAI21_X1   g13596(.A1(new_n13784_), .A2(new_n12101_), .B(new_n13788_), .ZN(new_n13789_));
  NAND2_X1   g13597(.A1(new_n13789_), .A2(new_n13783_), .ZN(new_n13790_));
  OAI22_X1   g13598(.A1(new_n13784_), .A2(new_n12101_), .B1(new_n13772_), .B2(new_n13782_), .ZN(new_n13791_));
  NAND2_X1   g13599(.A1(new_n13211_), .A2(new_n13212_), .ZN(new_n13792_));
  NAND4_X1   g13600(.A1(\asqrt[17] ), .A2(new_n11631_), .A3(new_n13792_), .A4(new_n13216_), .ZN(new_n13793_));
  XOR2_X1    g13601(.A1(new_n13793_), .A2(new_n13225_), .Z(new_n13794_));
  NAND2_X1   g13602(.A1(new_n13794_), .A2(new_n11105_), .ZN(new_n13795_));
  AOI21_X1   g13603(.A1(new_n13791_), .A2(\asqrt[21] ), .B(new_n13795_), .ZN(new_n13796_));
  NOR2_X1    g13604(.A1(new_n13796_), .A2(new_n13790_), .ZN(new_n13797_));
  AOI22_X1   g13605(.A1(new_n13791_), .A2(\asqrt[21] ), .B1(new_n13789_), .B2(new_n13783_), .ZN(new_n13798_));
  NOR4_X1    g13606(.A1(new_n13760_), .A2(\asqrt[22] ), .A3(new_n13220_), .A4(new_n13516_), .ZN(new_n13799_));
  XOR2_X1    g13607(.A1(new_n13799_), .A2(new_n13226_), .Z(new_n13800_));
  NAND2_X1   g13608(.A1(new_n13800_), .A2(new_n10614_), .ZN(new_n13801_));
  INV_X1     g13609(.I(new_n13801_), .ZN(new_n13802_));
  OAI21_X1   g13610(.A1(new_n13798_), .A2(new_n11105_), .B(new_n13802_), .ZN(new_n13803_));
  NAND2_X1   g13611(.A1(new_n13803_), .A2(new_n13797_), .ZN(new_n13804_));
  OAI22_X1   g13612(.A1(new_n13798_), .A2(new_n11105_), .B1(new_n13796_), .B2(new_n13790_), .ZN(new_n13805_));
  NOR4_X1    g13613(.A1(new_n13760_), .A2(\asqrt[23] ), .A3(new_n13230_), .A4(new_n13252_), .ZN(new_n13806_));
  XNOR2_X1   g13614(.A1(new_n13806_), .A2(new_n13262_), .ZN(new_n13807_));
  NAND2_X1   g13615(.A1(new_n13807_), .A2(new_n10104_), .ZN(new_n13808_));
  AOI21_X1   g13616(.A1(new_n13805_), .A2(\asqrt[23] ), .B(new_n13808_), .ZN(new_n13809_));
  NOR2_X1    g13617(.A1(new_n13809_), .A2(new_n13804_), .ZN(new_n13810_));
  AOI22_X1   g13618(.A1(new_n13805_), .A2(\asqrt[23] ), .B1(new_n13803_), .B2(new_n13797_), .ZN(new_n13811_));
  NOR4_X1    g13619(.A1(new_n13760_), .A2(\asqrt[24] ), .A3(new_n13256_), .A4(new_n13521_), .ZN(new_n13812_));
  XOR2_X1    g13620(.A1(new_n13812_), .A2(new_n13263_), .Z(new_n13813_));
  NAND2_X1   g13621(.A1(new_n13813_), .A2(new_n9672_), .ZN(new_n13814_));
  INV_X1     g13622(.I(new_n13814_), .ZN(new_n13815_));
  OAI21_X1   g13623(.A1(new_n13811_), .A2(new_n10104_), .B(new_n13815_), .ZN(new_n13816_));
  NAND2_X1   g13624(.A1(new_n13816_), .A2(new_n13810_), .ZN(new_n13817_));
  OAI22_X1   g13625(.A1(new_n13811_), .A2(new_n10104_), .B1(new_n13809_), .B2(new_n13804_), .ZN(new_n13818_));
  NOR4_X1    g13626(.A1(new_n13760_), .A2(\asqrt[25] ), .A3(new_n13266_), .A4(new_n13272_), .ZN(new_n13819_));
  XNOR2_X1   g13627(.A1(new_n13819_), .A2(new_n13281_), .ZN(new_n13820_));
  NAND2_X1   g13628(.A1(new_n13820_), .A2(new_n9212_), .ZN(new_n13821_));
  AOI21_X1   g13629(.A1(new_n13818_), .A2(\asqrt[25] ), .B(new_n13821_), .ZN(new_n13822_));
  NOR2_X1    g13630(.A1(new_n13822_), .A2(new_n13817_), .ZN(new_n13823_));
  AOI22_X1   g13631(.A1(new_n13818_), .A2(\asqrt[25] ), .B1(new_n13816_), .B2(new_n13810_), .ZN(new_n13824_));
  NOR4_X1    g13632(.A1(new_n13760_), .A2(\asqrt[26] ), .A3(new_n13275_), .A4(new_n13527_), .ZN(new_n13825_));
  XOR2_X1    g13633(.A1(new_n13825_), .A2(new_n13282_), .Z(new_n13826_));
  NAND2_X1   g13634(.A1(new_n13826_), .A2(new_n8763_), .ZN(new_n13827_));
  INV_X1     g13635(.I(new_n13827_), .ZN(new_n13828_));
  OAI21_X1   g13636(.A1(new_n13824_), .A2(new_n9212_), .B(new_n13828_), .ZN(new_n13829_));
  NAND2_X1   g13637(.A1(new_n13829_), .A2(new_n13823_), .ZN(new_n13830_));
  OAI22_X1   g13638(.A1(new_n13824_), .A2(new_n9212_), .B1(new_n13822_), .B2(new_n13817_), .ZN(new_n13831_));
  NAND2_X1   g13639(.A1(new_n13291_), .A2(\asqrt[27] ), .ZN(new_n13832_));
  NOR4_X1    g13640(.A1(new_n13760_), .A2(\asqrt[27] ), .A3(new_n13285_), .A4(new_n13291_), .ZN(new_n13833_));
  XOR2_X1    g13641(.A1(new_n13833_), .A2(new_n13832_), .Z(new_n13834_));
  NAND2_X1   g13642(.A1(new_n13834_), .A2(new_n8319_), .ZN(new_n13835_));
  AOI21_X1   g13643(.A1(new_n13831_), .A2(\asqrt[27] ), .B(new_n13835_), .ZN(new_n13836_));
  NOR2_X1    g13644(.A1(new_n13836_), .A2(new_n13830_), .ZN(new_n13837_));
  AOI22_X1   g13645(.A1(new_n13831_), .A2(\asqrt[27] ), .B1(new_n13829_), .B2(new_n13823_), .ZN(new_n13838_));
  NOR4_X1    g13646(.A1(new_n13760_), .A2(\asqrt[28] ), .A3(new_n13294_), .A4(new_n13534_), .ZN(new_n13839_));
  AOI21_X1   g13647(.A1(new_n13832_), .A2(new_n13289_), .B(new_n8319_), .ZN(new_n13840_));
  NOR2_X1    g13648(.A1(new_n13839_), .A2(new_n13840_), .ZN(new_n13841_));
  NAND2_X1   g13649(.A1(new_n13841_), .A2(new_n7931_), .ZN(new_n13842_));
  INV_X1     g13650(.I(new_n13842_), .ZN(new_n13843_));
  OAI21_X1   g13651(.A1(new_n13838_), .A2(new_n8319_), .B(new_n13843_), .ZN(new_n13844_));
  NAND2_X1   g13652(.A1(new_n13844_), .A2(new_n13837_), .ZN(new_n13845_));
  OAI22_X1   g13653(.A1(new_n13838_), .A2(new_n8319_), .B1(new_n13836_), .B2(new_n13830_), .ZN(new_n13846_));
  NAND2_X1   g13654(.A1(new_n13306_), .A2(\asqrt[29] ), .ZN(new_n13847_));
  NOR4_X1    g13655(.A1(new_n13760_), .A2(\asqrt[29] ), .A3(new_n13301_), .A4(new_n13306_), .ZN(new_n13848_));
  XOR2_X1    g13656(.A1(new_n13848_), .A2(new_n13847_), .Z(new_n13849_));
  NAND2_X1   g13657(.A1(new_n13849_), .A2(new_n7517_), .ZN(new_n13850_));
  AOI21_X1   g13658(.A1(new_n13846_), .A2(\asqrt[29] ), .B(new_n13850_), .ZN(new_n13851_));
  NOR2_X1    g13659(.A1(new_n13851_), .A2(new_n13845_), .ZN(new_n13852_));
  AOI22_X1   g13660(.A1(new_n13846_), .A2(\asqrt[29] ), .B1(new_n13844_), .B2(new_n13837_), .ZN(new_n13853_));
  NOR4_X1    g13661(.A1(new_n13760_), .A2(\asqrt[30] ), .A3(new_n13309_), .A4(new_n13541_), .ZN(new_n13854_));
  AOI21_X1   g13662(.A1(new_n13847_), .A2(new_n13305_), .B(new_n7517_), .ZN(new_n13855_));
  NOR2_X1    g13663(.A1(new_n13854_), .A2(new_n13855_), .ZN(new_n13856_));
  NAND2_X1   g13664(.A1(new_n13856_), .A2(new_n7110_), .ZN(new_n13857_));
  INV_X1     g13665(.I(new_n13857_), .ZN(new_n13858_));
  OAI21_X1   g13666(.A1(new_n13853_), .A2(new_n7517_), .B(new_n13858_), .ZN(new_n13859_));
  NAND2_X1   g13667(.A1(new_n13859_), .A2(new_n13852_), .ZN(new_n13860_));
  OAI22_X1   g13668(.A1(new_n13853_), .A2(new_n7517_), .B1(new_n13851_), .B2(new_n13845_), .ZN(new_n13861_));
  NAND2_X1   g13669(.A1(new_n13321_), .A2(\asqrt[31] ), .ZN(new_n13862_));
  NOR4_X1    g13670(.A1(new_n13760_), .A2(\asqrt[31] ), .A3(new_n13316_), .A4(new_n13321_), .ZN(new_n13863_));
  XOR2_X1    g13671(.A1(new_n13863_), .A2(new_n13862_), .Z(new_n13864_));
  NAND2_X1   g13672(.A1(new_n13864_), .A2(new_n6708_), .ZN(new_n13865_));
  AOI21_X1   g13673(.A1(new_n13861_), .A2(\asqrt[31] ), .B(new_n13865_), .ZN(new_n13866_));
  NOR2_X1    g13674(.A1(new_n13866_), .A2(new_n13860_), .ZN(new_n13867_));
  AOI22_X1   g13675(.A1(new_n13861_), .A2(\asqrt[31] ), .B1(new_n13859_), .B2(new_n13852_), .ZN(new_n13868_));
  NOR4_X1    g13676(.A1(new_n13760_), .A2(\asqrt[32] ), .A3(new_n13324_), .A4(new_n13548_), .ZN(new_n13869_));
  AOI21_X1   g13677(.A1(new_n13862_), .A2(new_n13320_), .B(new_n6708_), .ZN(new_n13870_));
  NOR2_X1    g13678(.A1(new_n13869_), .A2(new_n13870_), .ZN(new_n13871_));
  NAND2_X1   g13679(.A1(new_n13871_), .A2(new_n6365_), .ZN(new_n13872_));
  INV_X1     g13680(.I(new_n13872_), .ZN(new_n13873_));
  OAI21_X1   g13681(.A1(new_n13868_), .A2(new_n6708_), .B(new_n13873_), .ZN(new_n13874_));
  NAND2_X1   g13682(.A1(new_n13874_), .A2(new_n13867_), .ZN(new_n13875_));
  OAI22_X1   g13683(.A1(new_n13868_), .A2(new_n6708_), .B1(new_n13866_), .B2(new_n13860_), .ZN(new_n13876_));
  NAND2_X1   g13684(.A1(new_n13336_), .A2(\asqrt[33] ), .ZN(new_n13877_));
  NOR4_X1    g13685(.A1(new_n13760_), .A2(\asqrt[33] ), .A3(new_n13331_), .A4(new_n13336_), .ZN(new_n13878_));
  XOR2_X1    g13686(.A1(new_n13878_), .A2(new_n13877_), .Z(new_n13879_));
  NAND2_X1   g13687(.A1(new_n13879_), .A2(new_n5991_), .ZN(new_n13880_));
  AOI21_X1   g13688(.A1(new_n13876_), .A2(\asqrt[33] ), .B(new_n13880_), .ZN(new_n13881_));
  NOR2_X1    g13689(.A1(new_n13881_), .A2(new_n13875_), .ZN(new_n13882_));
  AOI22_X1   g13690(.A1(new_n13876_), .A2(\asqrt[33] ), .B1(new_n13874_), .B2(new_n13867_), .ZN(new_n13883_));
  NOR4_X1    g13691(.A1(new_n13760_), .A2(\asqrt[34] ), .A3(new_n13339_), .A4(new_n13555_), .ZN(new_n13884_));
  AOI21_X1   g13692(.A1(new_n13877_), .A2(new_n13335_), .B(new_n5991_), .ZN(new_n13885_));
  NOR2_X1    g13693(.A1(new_n13884_), .A2(new_n13885_), .ZN(new_n13886_));
  NAND2_X1   g13694(.A1(new_n13886_), .A2(new_n5626_), .ZN(new_n13887_));
  INV_X1     g13695(.I(new_n13887_), .ZN(new_n13888_));
  OAI21_X1   g13696(.A1(new_n13883_), .A2(new_n5991_), .B(new_n13888_), .ZN(new_n13889_));
  NAND2_X1   g13697(.A1(new_n13889_), .A2(new_n13882_), .ZN(new_n13890_));
  OAI22_X1   g13698(.A1(new_n13883_), .A2(new_n5991_), .B1(new_n13881_), .B2(new_n13875_), .ZN(new_n13891_));
  NAND2_X1   g13699(.A1(new_n13351_), .A2(\asqrt[35] ), .ZN(new_n13892_));
  NOR4_X1    g13700(.A1(new_n13760_), .A2(\asqrt[35] ), .A3(new_n13346_), .A4(new_n13351_), .ZN(new_n13893_));
  XOR2_X1    g13701(.A1(new_n13893_), .A2(new_n13892_), .Z(new_n13894_));
  NAND2_X1   g13702(.A1(new_n13894_), .A2(new_n5273_), .ZN(new_n13895_));
  AOI21_X1   g13703(.A1(new_n13891_), .A2(\asqrt[35] ), .B(new_n13895_), .ZN(new_n13896_));
  NOR2_X1    g13704(.A1(new_n13896_), .A2(new_n13890_), .ZN(new_n13897_));
  AOI22_X1   g13705(.A1(new_n13891_), .A2(\asqrt[35] ), .B1(new_n13889_), .B2(new_n13882_), .ZN(new_n13898_));
  NOR4_X1    g13706(.A1(new_n13760_), .A2(\asqrt[36] ), .A3(new_n13354_), .A4(new_n13562_), .ZN(new_n13899_));
  AOI21_X1   g13707(.A1(new_n13892_), .A2(new_n13350_), .B(new_n5273_), .ZN(new_n13900_));
  NOR2_X1    g13708(.A1(new_n13899_), .A2(new_n13900_), .ZN(new_n13901_));
  NAND2_X1   g13709(.A1(new_n13901_), .A2(new_n4973_), .ZN(new_n13902_));
  INV_X1     g13710(.I(new_n13902_), .ZN(new_n13903_));
  OAI21_X1   g13711(.A1(new_n13898_), .A2(new_n5273_), .B(new_n13903_), .ZN(new_n13904_));
  NAND2_X1   g13712(.A1(new_n13904_), .A2(new_n13897_), .ZN(new_n13905_));
  OAI22_X1   g13713(.A1(new_n13898_), .A2(new_n5273_), .B1(new_n13896_), .B2(new_n13890_), .ZN(new_n13906_));
  NAND2_X1   g13714(.A1(new_n13366_), .A2(\asqrt[37] ), .ZN(new_n13907_));
  NOR4_X1    g13715(.A1(new_n13760_), .A2(\asqrt[37] ), .A3(new_n13361_), .A4(new_n13366_), .ZN(new_n13908_));
  XOR2_X1    g13716(.A1(new_n13908_), .A2(new_n13907_), .Z(new_n13909_));
  NAND2_X1   g13717(.A1(new_n13909_), .A2(new_n4645_), .ZN(new_n13910_));
  AOI21_X1   g13718(.A1(new_n13906_), .A2(\asqrt[37] ), .B(new_n13910_), .ZN(new_n13911_));
  NOR2_X1    g13719(.A1(new_n13911_), .A2(new_n13905_), .ZN(new_n13912_));
  AOI22_X1   g13720(.A1(new_n13906_), .A2(\asqrt[37] ), .B1(new_n13904_), .B2(new_n13897_), .ZN(new_n13913_));
  NAND2_X1   g13721(.A1(new_n13569_), .A2(\asqrt[38] ), .ZN(new_n13914_));
  NOR4_X1    g13722(.A1(new_n13760_), .A2(\asqrt[38] ), .A3(new_n13369_), .A4(new_n13569_), .ZN(new_n13915_));
  XOR2_X1    g13723(.A1(new_n13915_), .A2(new_n13914_), .Z(new_n13916_));
  NAND2_X1   g13724(.A1(new_n13916_), .A2(new_n4330_), .ZN(new_n13917_));
  INV_X1     g13725(.I(new_n13917_), .ZN(new_n13918_));
  OAI21_X1   g13726(.A1(new_n13913_), .A2(new_n4645_), .B(new_n13918_), .ZN(new_n13919_));
  NAND2_X1   g13727(.A1(new_n13919_), .A2(new_n13912_), .ZN(new_n13920_));
  OAI22_X1   g13728(.A1(new_n13913_), .A2(new_n4645_), .B1(new_n13911_), .B2(new_n13905_), .ZN(new_n13921_));
  NOR4_X1    g13729(.A1(new_n13760_), .A2(\asqrt[39] ), .A3(new_n13376_), .A4(new_n13381_), .ZN(new_n13922_));
  AOI21_X1   g13730(.A1(new_n13914_), .A2(new_n13568_), .B(new_n4330_), .ZN(new_n13923_));
  NOR2_X1    g13731(.A1(new_n13922_), .A2(new_n13923_), .ZN(new_n13924_));
  NAND2_X1   g13732(.A1(new_n13924_), .A2(new_n4018_), .ZN(new_n13925_));
  AOI21_X1   g13733(.A1(new_n13921_), .A2(\asqrt[39] ), .B(new_n13925_), .ZN(new_n13926_));
  NOR2_X1    g13734(.A1(new_n13926_), .A2(new_n13920_), .ZN(new_n13927_));
  AOI22_X1   g13735(.A1(new_n13921_), .A2(\asqrt[39] ), .B1(new_n13919_), .B2(new_n13912_), .ZN(new_n13928_));
  NAND2_X1   g13736(.A1(new_n13576_), .A2(\asqrt[40] ), .ZN(new_n13929_));
  NOR4_X1    g13737(.A1(new_n13760_), .A2(\asqrt[40] ), .A3(new_n13384_), .A4(new_n13576_), .ZN(new_n13930_));
  XOR2_X1    g13738(.A1(new_n13930_), .A2(new_n13929_), .Z(new_n13931_));
  NAND2_X1   g13739(.A1(new_n13931_), .A2(new_n3760_), .ZN(new_n13932_));
  INV_X1     g13740(.I(new_n13932_), .ZN(new_n13933_));
  OAI21_X1   g13741(.A1(new_n13928_), .A2(new_n4018_), .B(new_n13933_), .ZN(new_n13934_));
  NAND2_X1   g13742(.A1(new_n13934_), .A2(new_n13927_), .ZN(new_n13935_));
  OAI22_X1   g13743(.A1(new_n13928_), .A2(new_n4018_), .B1(new_n13926_), .B2(new_n13920_), .ZN(new_n13936_));
  NOR4_X1    g13744(.A1(new_n13760_), .A2(\asqrt[41] ), .A3(new_n13391_), .A4(new_n13396_), .ZN(new_n13937_));
  AOI21_X1   g13745(.A1(new_n13929_), .A2(new_n13575_), .B(new_n3760_), .ZN(new_n13938_));
  NOR2_X1    g13746(.A1(new_n13937_), .A2(new_n13938_), .ZN(new_n13939_));
  NAND2_X1   g13747(.A1(new_n13939_), .A2(new_n3481_), .ZN(new_n13940_));
  AOI21_X1   g13748(.A1(new_n13936_), .A2(\asqrt[41] ), .B(new_n13940_), .ZN(new_n13941_));
  NOR2_X1    g13749(.A1(new_n13941_), .A2(new_n13935_), .ZN(new_n13942_));
  AOI22_X1   g13750(.A1(new_n13936_), .A2(\asqrt[41] ), .B1(new_n13934_), .B2(new_n13927_), .ZN(new_n13943_));
  NAND2_X1   g13751(.A1(new_n13583_), .A2(\asqrt[42] ), .ZN(new_n13944_));
  NOR4_X1    g13752(.A1(new_n13760_), .A2(\asqrt[42] ), .A3(new_n13399_), .A4(new_n13583_), .ZN(new_n13945_));
  XOR2_X1    g13753(.A1(new_n13945_), .A2(new_n13944_), .Z(new_n13946_));
  NAND2_X1   g13754(.A1(new_n13946_), .A2(new_n3208_), .ZN(new_n13947_));
  INV_X1     g13755(.I(new_n13947_), .ZN(new_n13948_));
  OAI21_X1   g13756(.A1(new_n13943_), .A2(new_n3481_), .B(new_n13948_), .ZN(new_n13949_));
  NAND2_X1   g13757(.A1(new_n13949_), .A2(new_n13942_), .ZN(new_n13950_));
  OAI22_X1   g13758(.A1(new_n13943_), .A2(new_n3481_), .B1(new_n13941_), .B2(new_n13935_), .ZN(new_n13951_));
  NAND2_X1   g13759(.A1(new_n13411_), .A2(\asqrt[43] ), .ZN(new_n13952_));
  NOR4_X1    g13760(.A1(new_n13760_), .A2(\asqrt[43] ), .A3(new_n13406_), .A4(new_n13411_), .ZN(new_n13953_));
  XOR2_X1    g13761(.A1(new_n13953_), .A2(new_n13952_), .Z(new_n13954_));
  NAND2_X1   g13762(.A1(new_n13954_), .A2(new_n2941_), .ZN(new_n13955_));
  AOI21_X1   g13763(.A1(new_n13951_), .A2(\asqrt[43] ), .B(new_n13955_), .ZN(new_n13956_));
  NOR2_X1    g13764(.A1(new_n13956_), .A2(new_n13950_), .ZN(new_n13957_));
  AOI22_X1   g13765(.A1(new_n13951_), .A2(\asqrt[43] ), .B1(new_n13949_), .B2(new_n13942_), .ZN(new_n13958_));
  NOR4_X1    g13766(.A1(new_n13760_), .A2(\asqrt[44] ), .A3(new_n13414_), .A4(new_n13590_), .ZN(new_n13959_));
  AOI21_X1   g13767(.A1(new_n13952_), .A2(new_n13410_), .B(new_n2941_), .ZN(new_n13960_));
  NOR2_X1    g13768(.A1(new_n13959_), .A2(new_n13960_), .ZN(new_n13961_));
  NAND2_X1   g13769(.A1(new_n13961_), .A2(new_n2728_), .ZN(new_n13962_));
  INV_X1     g13770(.I(new_n13962_), .ZN(new_n13963_));
  OAI21_X1   g13771(.A1(new_n13958_), .A2(new_n2941_), .B(new_n13963_), .ZN(new_n13964_));
  NAND2_X1   g13772(.A1(new_n13964_), .A2(new_n13957_), .ZN(new_n13965_));
  OAI22_X1   g13773(.A1(new_n13958_), .A2(new_n2941_), .B1(new_n13956_), .B2(new_n13950_), .ZN(new_n13966_));
  NAND2_X1   g13774(.A1(new_n13426_), .A2(\asqrt[45] ), .ZN(new_n13967_));
  NOR4_X1    g13775(.A1(new_n13760_), .A2(\asqrt[45] ), .A3(new_n13421_), .A4(new_n13426_), .ZN(new_n13968_));
  XOR2_X1    g13776(.A1(new_n13968_), .A2(new_n13967_), .Z(new_n13969_));
  NAND2_X1   g13777(.A1(new_n13969_), .A2(new_n2488_), .ZN(new_n13970_));
  AOI21_X1   g13778(.A1(new_n13966_), .A2(\asqrt[45] ), .B(new_n13970_), .ZN(new_n13971_));
  NOR2_X1    g13779(.A1(new_n13971_), .A2(new_n13965_), .ZN(new_n13972_));
  AOI22_X1   g13780(.A1(new_n13966_), .A2(\asqrt[45] ), .B1(new_n13964_), .B2(new_n13957_), .ZN(new_n13973_));
  NOR4_X1    g13781(.A1(new_n13760_), .A2(\asqrt[46] ), .A3(new_n13429_), .A4(new_n13597_), .ZN(new_n13974_));
  AOI21_X1   g13782(.A1(new_n13967_), .A2(new_n13425_), .B(new_n2488_), .ZN(new_n13975_));
  NOR2_X1    g13783(.A1(new_n13974_), .A2(new_n13975_), .ZN(new_n13976_));
  NAND2_X1   g13784(.A1(new_n13976_), .A2(new_n2253_), .ZN(new_n13977_));
  INV_X1     g13785(.I(new_n13977_), .ZN(new_n13978_));
  OAI21_X1   g13786(.A1(new_n13973_), .A2(new_n2488_), .B(new_n13978_), .ZN(new_n13979_));
  NAND2_X1   g13787(.A1(new_n13979_), .A2(new_n13972_), .ZN(new_n13980_));
  OAI22_X1   g13788(.A1(new_n13973_), .A2(new_n2488_), .B1(new_n13971_), .B2(new_n13965_), .ZN(new_n13981_));
  NAND2_X1   g13789(.A1(new_n13441_), .A2(\asqrt[47] ), .ZN(new_n13982_));
  NOR4_X1    g13790(.A1(new_n13760_), .A2(\asqrt[47] ), .A3(new_n13436_), .A4(new_n13441_), .ZN(new_n13983_));
  XOR2_X1    g13791(.A1(new_n13983_), .A2(new_n13982_), .Z(new_n13984_));
  NAND2_X1   g13792(.A1(new_n13984_), .A2(new_n2046_), .ZN(new_n13985_));
  AOI21_X1   g13793(.A1(new_n13981_), .A2(\asqrt[47] ), .B(new_n13985_), .ZN(new_n13986_));
  NOR2_X1    g13794(.A1(new_n13986_), .A2(new_n13980_), .ZN(new_n13987_));
  AOI22_X1   g13795(.A1(new_n13981_), .A2(\asqrt[47] ), .B1(new_n13979_), .B2(new_n13972_), .ZN(new_n13988_));
  NOR4_X1    g13796(.A1(new_n13760_), .A2(\asqrt[48] ), .A3(new_n13444_), .A4(new_n13604_), .ZN(new_n13989_));
  AOI21_X1   g13797(.A1(new_n13982_), .A2(new_n13440_), .B(new_n2046_), .ZN(new_n13990_));
  NOR2_X1    g13798(.A1(new_n13989_), .A2(new_n13990_), .ZN(new_n13991_));
  NAND2_X1   g13799(.A1(new_n13991_), .A2(new_n1854_), .ZN(new_n13992_));
  INV_X1     g13800(.I(new_n13992_), .ZN(new_n13993_));
  OAI21_X1   g13801(.A1(new_n13988_), .A2(new_n2046_), .B(new_n13993_), .ZN(new_n13994_));
  NAND2_X1   g13802(.A1(new_n13994_), .A2(new_n13987_), .ZN(new_n13995_));
  OAI22_X1   g13803(.A1(new_n13988_), .A2(new_n2046_), .B1(new_n13986_), .B2(new_n13980_), .ZN(new_n13996_));
  NAND2_X1   g13804(.A1(new_n13456_), .A2(\asqrt[49] ), .ZN(new_n13997_));
  NOR4_X1    g13805(.A1(new_n13760_), .A2(\asqrt[49] ), .A3(new_n13451_), .A4(new_n13456_), .ZN(new_n13998_));
  XOR2_X1    g13806(.A1(new_n13998_), .A2(new_n13997_), .Z(new_n13999_));
  NAND2_X1   g13807(.A1(new_n13999_), .A2(new_n1595_), .ZN(new_n14000_));
  AOI21_X1   g13808(.A1(new_n13996_), .A2(\asqrt[49] ), .B(new_n14000_), .ZN(new_n14001_));
  NOR2_X1    g13809(.A1(new_n14001_), .A2(new_n13995_), .ZN(new_n14002_));
  AOI22_X1   g13810(.A1(new_n13996_), .A2(\asqrt[49] ), .B1(new_n13994_), .B2(new_n13987_), .ZN(new_n14003_));
  NAND2_X1   g13811(.A1(new_n13611_), .A2(\asqrt[50] ), .ZN(new_n14004_));
  NOR4_X1    g13812(.A1(new_n13760_), .A2(\asqrt[50] ), .A3(new_n13459_), .A4(new_n13611_), .ZN(new_n14005_));
  XOR2_X1    g13813(.A1(new_n14005_), .A2(new_n14004_), .Z(new_n14006_));
  NAND2_X1   g13814(.A1(new_n14006_), .A2(new_n1436_), .ZN(new_n14007_));
  INV_X1     g13815(.I(new_n14007_), .ZN(new_n14008_));
  OAI21_X1   g13816(.A1(new_n14003_), .A2(new_n1595_), .B(new_n14008_), .ZN(new_n14009_));
  NAND2_X1   g13817(.A1(new_n14009_), .A2(new_n14002_), .ZN(new_n14010_));
  OAI22_X1   g13818(.A1(new_n14003_), .A2(new_n1595_), .B1(new_n14001_), .B2(new_n13995_), .ZN(new_n14011_));
  NOR4_X1    g13819(.A1(new_n13760_), .A2(\asqrt[51] ), .A3(new_n13466_), .A4(new_n13471_), .ZN(new_n14012_));
  AOI21_X1   g13820(.A1(new_n14004_), .A2(new_n13610_), .B(new_n1436_), .ZN(new_n14013_));
  NOR2_X1    g13821(.A1(new_n14012_), .A2(new_n14013_), .ZN(new_n14014_));
  NAND2_X1   g13822(.A1(new_n14014_), .A2(new_n1260_), .ZN(new_n14015_));
  AOI21_X1   g13823(.A1(new_n14011_), .A2(\asqrt[51] ), .B(new_n14015_), .ZN(new_n14016_));
  NOR2_X1    g13824(.A1(new_n14016_), .A2(new_n14010_), .ZN(new_n14017_));
  AOI22_X1   g13825(.A1(new_n14011_), .A2(\asqrt[51] ), .B1(new_n14009_), .B2(new_n14002_), .ZN(new_n14018_));
  NOR4_X1    g13826(.A1(new_n13760_), .A2(\asqrt[52] ), .A3(new_n13474_), .A4(new_n13618_), .ZN(new_n14019_));
  XOR2_X1    g13827(.A1(new_n14019_), .A2(new_n13628_), .Z(new_n14020_));
  NAND2_X1   g13828(.A1(new_n14020_), .A2(new_n1096_), .ZN(new_n14021_));
  INV_X1     g13829(.I(new_n14021_), .ZN(new_n14022_));
  OAI21_X1   g13830(.A1(new_n14018_), .A2(new_n1260_), .B(new_n14022_), .ZN(new_n14023_));
  NAND2_X1   g13831(.A1(new_n14023_), .A2(new_n14017_), .ZN(new_n14024_));
  OAI22_X1   g13832(.A1(new_n14018_), .A2(new_n1260_), .B1(new_n14016_), .B2(new_n14010_), .ZN(new_n14025_));
  NOR4_X1    g13833(.A1(new_n13760_), .A2(\asqrt[53] ), .A3(new_n13481_), .A4(new_n13486_), .ZN(new_n14026_));
  XNOR2_X1   g13834(.A1(new_n14026_), .A2(new_n13629_), .ZN(new_n14027_));
  NAND2_X1   g13835(.A1(new_n14027_), .A2(new_n970_), .ZN(new_n14028_));
  AOI21_X1   g13836(.A1(new_n14025_), .A2(\asqrt[53] ), .B(new_n14028_), .ZN(new_n14029_));
  NOR2_X1    g13837(.A1(new_n14029_), .A2(new_n14024_), .ZN(new_n14030_));
  AOI22_X1   g13838(.A1(new_n14025_), .A2(\asqrt[53] ), .B1(new_n14023_), .B2(new_n14017_), .ZN(new_n14031_));
  NOR4_X1    g13839(.A1(new_n13760_), .A2(\asqrt[54] ), .A3(new_n13489_), .A4(new_n13625_), .ZN(new_n14032_));
  XOR2_X1    g13840(.A1(new_n14032_), .A2(new_n13630_), .Z(new_n14033_));
  NAND2_X1   g13841(.A1(new_n14033_), .A2(new_n825_), .ZN(new_n14034_));
  INV_X1     g13842(.I(new_n14034_), .ZN(new_n14035_));
  OAI21_X1   g13843(.A1(new_n14031_), .A2(new_n970_), .B(new_n14035_), .ZN(new_n14036_));
  NAND2_X1   g13844(.A1(new_n14036_), .A2(new_n14030_), .ZN(new_n14037_));
  OAI22_X1   g13845(.A1(new_n14031_), .A2(new_n970_), .B1(new_n14029_), .B2(new_n14024_), .ZN(new_n14038_));
  NOR4_X1    g13846(.A1(new_n13760_), .A2(\asqrt[55] ), .A3(new_n13496_), .A4(new_n13501_), .ZN(new_n14039_));
  XNOR2_X1   g13847(.A1(new_n14039_), .A2(new_n13631_), .ZN(new_n14040_));
  NAND2_X1   g13848(.A1(new_n14040_), .A2(new_n724_), .ZN(new_n14041_));
  AOI21_X1   g13849(.A1(new_n14038_), .A2(\asqrt[55] ), .B(new_n14041_), .ZN(new_n14042_));
  NOR2_X1    g13850(.A1(new_n14042_), .A2(new_n14037_), .ZN(new_n14043_));
  AOI22_X1   g13851(.A1(new_n14038_), .A2(\asqrt[55] ), .B1(new_n14036_), .B2(new_n14030_), .ZN(new_n14044_));
  NOR4_X1    g13852(.A1(new_n13760_), .A2(\asqrt[56] ), .A3(new_n13504_), .A4(new_n13657_), .ZN(new_n14045_));
  XOR2_X1    g13853(.A1(new_n14045_), .A2(new_n13632_), .Z(new_n14046_));
  NAND2_X1   g13854(.A1(new_n14046_), .A2(new_n587_), .ZN(new_n14047_));
  INV_X1     g13855(.I(new_n14047_), .ZN(new_n14048_));
  OAI21_X1   g13856(.A1(new_n14044_), .A2(new_n724_), .B(new_n14048_), .ZN(new_n14049_));
  NAND2_X1   g13857(.A1(new_n14049_), .A2(new_n14043_), .ZN(new_n14050_));
  OAI22_X1   g13858(.A1(new_n14044_), .A2(new_n724_), .B1(new_n14042_), .B2(new_n14037_), .ZN(new_n14051_));
  NOR4_X1    g13859(.A1(new_n13760_), .A2(\asqrt[57] ), .A3(new_n13511_), .A4(new_n13639_), .ZN(new_n14052_));
  XOR2_X1    g13860(.A1(new_n14052_), .A2(new_n13634_), .Z(new_n14053_));
  NAND2_X1   g13861(.A1(new_n14053_), .A2(new_n504_), .ZN(new_n14054_));
  AOI21_X1   g13862(.A1(new_n14051_), .A2(\asqrt[57] ), .B(new_n14054_), .ZN(new_n14055_));
  NOR2_X1    g13863(.A1(new_n14055_), .A2(new_n14050_), .ZN(new_n14056_));
  AOI22_X1   g13864(.A1(new_n14051_), .A2(\asqrt[57] ), .B1(new_n14049_), .B2(new_n14043_), .ZN(new_n14057_));
  NOR4_X1    g13865(.A1(new_n13760_), .A2(\asqrt[58] ), .A3(new_n13636_), .A4(new_n13672_), .ZN(new_n14058_));
  XOR2_X1    g13866(.A1(new_n14058_), .A2(new_n13664_), .Z(new_n14059_));
  NAND2_X1   g13867(.A1(new_n14059_), .A2(new_n376_), .ZN(new_n14060_));
  INV_X1     g13868(.I(new_n14060_), .ZN(new_n14061_));
  OAI21_X1   g13869(.A1(new_n14057_), .A2(new_n504_), .B(new_n14061_), .ZN(new_n14062_));
  NAND2_X1   g13870(.A1(new_n14062_), .A2(new_n14056_), .ZN(new_n14063_));
  OAI22_X1   g13871(.A1(new_n14057_), .A2(new_n504_), .B1(new_n14055_), .B2(new_n14050_), .ZN(new_n14064_));
  NOR4_X1    g13872(.A1(new_n13760_), .A2(\asqrt[59] ), .A3(new_n13642_), .A4(new_n13665_), .ZN(new_n14065_));
  XOR2_X1    g13873(.A1(new_n14065_), .A2(new_n13648_), .Z(new_n14066_));
  NAND2_X1   g13874(.A1(new_n14066_), .A2(new_n275_), .ZN(new_n14067_));
  AOI21_X1   g13875(.A1(new_n14064_), .A2(\asqrt[59] ), .B(new_n14067_), .ZN(new_n14068_));
  NOR2_X1    g13876(.A1(new_n14068_), .A2(new_n14063_), .ZN(new_n14069_));
  AOI22_X1   g13877(.A1(new_n14064_), .A2(\asqrt[59] ), .B1(new_n14062_), .B2(new_n14056_), .ZN(new_n14070_));
  NOR4_X1    g13878(.A1(new_n13760_), .A2(\asqrt[60] ), .A3(new_n13650_), .A4(new_n13688_), .ZN(new_n14071_));
  XOR2_X1    g13879(.A1(new_n14071_), .A2(new_n13679_), .Z(new_n14072_));
  NAND2_X1   g13880(.A1(new_n14072_), .A2(new_n229_), .ZN(new_n14073_));
  INV_X1     g13881(.I(new_n14073_), .ZN(new_n14074_));
  OAI21_X1   g13882(.A1(new_n14070_), .A2(new_n275_), .B(new_n14074_), .ZN(new_n14075_));
  NAND2_X1   g13883(.A1(new_n14075_), .A2(new_n14069_), .ZN(new_n14076_));
  OAI22_X1   g13884(.A1(new_n14070_), .A2(new_n275_), .B1(new_n14068_), .B2(new_n14063_), .ZN(new_n14077_));
  INV_X1     g13885(.I(new_n13731_), .ZN(new_n14078_));
  NOR2_X1    g13886(.A1(new_n14078_), .A2(\asqrt[62] ), .ZN(new_n14079_));
  INV_X1     g13887(.I(new_n14079_), .ZN(new_n14080_));
  NAND3_X1   g13888(.A1(new_n14077_), .A2(\asqrt[61] ), .A3(new_n14080_), .ZN(new_n14081_));
  OAI21_X1   g13889(.A1(new_n14081_), .A2(new_n14076_), .B(new_n13733_), .ZN(new_n14082_));
  NAND3_X1   g13890(.A1(new_n13760_), .A2(new_n13154_), .A3(new_n13763_), .ZN(new_n14083_));
  AOI21_X1   g13891(.A1(new_n14083_), .A2(new_n13710_), .B(\asqrt[63] ), .ZN(new_n14084_));
  INV_X1     g13892(.I(new_n14084_), .ZN(new_n14085_));
  OAI21_X1   g13893(.A1(new_n14082_), .A2(new_n14085_), .B(new_n13728_), .ZN(new_n14086_));
  INV_X1     g13894(.I(new_n13742_), .ZN(new_n14087_));
  AOI21_X1   g13895(.A1(new_n13751_), .A2(new_n14087_), .B(new_n13744_), .ZN(new_n14088_));
  NOR3_X1    g13896(.A1(new_n13741_), .A2(new_n13734_), .A3(new_n13739_), .ZN(new_n14089_));
  NOR2_X1    g13897(.A1(new_n14089_), .A2(new_n14088_), .ZN(new_n14090_));
  NOR3_X1    g13898(.A1(new_n13769_), .A2(new_n13167_), .A3(\asqrt[17] ), .ZN(new_n14091_));
  AOI21_X1   g13899(.A1(new_n13766_), .A2(new_n13166_), .B(new_n13760_), .ZN(new_n14092_));
  NOR4_X1    g13900(.A1(new_n14092_), .A2(new_n14091_), .A3(\asqrt[19] ), .A4(new_n13758_), .ZN(new_n14093_));
  NOR2_X1    g13901(.A1(new_n14093_), .A2(new_n14090_), .ZN(new_n14094_));
  NOR3_X1    g13902(.A1(new_n14089_), .A2(new_n14088_), .A3(new_n13758_), .ZN(new_n14095_));
  NOR3_X1    g13903(.A1(new_n13760_), .A2(new_n13190_), .A3(new_n13777_), .ZN(new_n14096_));
  AOI21_X1   g13904(.A1(\asqrt[17] ), .A2(new_n13778_), .B(new_n13191_), .ZN(new_n14097_));
  NOR3_X1    g13905(.A1(new_n14097_), .A2(new_n14096_), .A3(\asqrt[20] ), .ZN(new_n14098_));
  OAI21_X1   g13906(.A1(new_n14095_), .A2(new_n12657_), .B(new_n14098_), .ZN(new_n14099_));
  NAND2_X1   g13907(.A1(new_n14094_), .A2(new_n14099_), .ZN(new_n14100_));
  OAI22_X1   g13908(.A1(new_n14093_), .A2(new_n14090_), .B1(new_n12657_), .B2(new_n14095_), .ZN(new_n14101_));
  INV_X1     g13909(.I(new_n13788_), .ZN(new_n14102_));
  AOI21_X1   g13910(.A1(new_n14101_), .A2(\asqrt[20] ), .B(new_n14102_), .ZN(new_n14103_));
  NOR2_X1    g13911(.A1(new_n14103_), .A2(new_n14100_), .ZN(new_n14104_));
  AOI22_X1   g13912(.A1(new_n14101_), .A2(\asqrt[20] ), .B1(new_n14094_), .B2(new_n14099_), .ZN(new_n14105_));
  INV_X1     g13913(.I(new_n13795_), .ZN(new_n14106_));
  OAI21_X1   g13914(.A1(new_n14105_), .A2(new_n11631_), .B(new_n14106_), .ZN(new_n14107_));
  NAND2_X1   g13915(.A1(new_n14107_), .A2(new_n14104_), .ZN(new_n14108_));
  OAI22_X1   g13916(.A1(new_n14105_), .A2(new_n11631_), .B1(new_n14103_), .B2(new_n14100_), .ZN(new_n14109_));
  AOI21_X1   g13917(.A1(new_n14109_), .A2(\asqrt[22] ), .B(new_n13801_), .ZN(new_n14110_));
  NOR2_X1    g13918(.A1(new_n14110_), .A2(new_n14108_), .ZN(new_n14111_));
  AOI22_X1   g13919(.A1(new_n14109_), .A2(\asqrt[22] ), .B1(new_n14107_), .B2(new_n14104_), .ZN(new_n14112_));
  INV_X1     g13920(.I(new_n13808_), .ZN(new_n14113_));
  OAI21_X1   g13921(.A1(new_n14112_), .A2(new_n10614_), .B(new_n14113_), .ZN(new_n14114_));
  NAND2_X1   g13922(.A1(new_n14114_), .A2(new_n14111_), .ZN(new_n14115_));
  OAI22_X1   g13923(.A1(new_n14112_), .A2(new_n10614_), .B1(new_n14110_), .B2(new_n14108_), .ZN(new_n14116_));
  AOI21_X1   g13924(.A1(new_n14116_), .A2(\asqrt[24] ), .B(new_n13814_), .ZN(new_n14117_));
  NOR2_X1    g13925(.A1(new_n14117_), .A2(new_n14115_), .ZN(new_n14118_));
  AOI22_X1   g13926(.A1(new_n14116_), .A2(\asqrt[24] ), .B1(new_n14114_), .B2(new_n14111_), .ZN(new_n14119_));
  INV_X1     g13927(.I(new_n13821_), .ZN(new_n14120_));
  OAI21_X1   g13928(.A1(new_n14119_), .A2(new_n9672_), .B(new_n14120_), .ZN(new_n14121_));
  NAND2_X1   g13929(.A1(new_n14121_), .A2(new_n14118_), .ZN(new_n14122_));
  OAI22_X1   g13930(.A1(new_n14119_), .A2(new_n9672_), .B1(new_n14117_), .B2(new_n14115_), .ZN(new_n14123_));
  AOI21_X1   g13931(.A1(new_n14123_), .A2(\asqrt[26] ), .B(new_n13827_), .ZN(new_n14124_));
  NOR2_X1    g13932(.A1(new_n14124_), .A2(new_n14122_), .ZN(new_n14125_));
  AOI22_X1   g13933(.A1(new_n14123_), .A2(\asqrt[26] ), .B1(new_n14121_), .B2(new_n14118_), .ZN(new_n14126_));
  INV_X1     g13934(.I(new_n13835_), .ZN(new_n14127_));
  OAI21_X1   g13935(.A1(new_n14126_), .A2(new_n8763_), .B(new_n14127_), .ZN(new_n14128_));
  NAND2_X1   g13936(.A1(new_n14128_), .A2(new_n14125_), .ZN(new_n14129_));
  OAI22_X1   g13937(.A1(new_n14126_), .A2(new_n8763_), .B1(new_n14124_), .B2(new_n14122_), .ZN(new_n14130_));
  AOI21_X1   g13938(.A1(new_n14130_), .A2(\asqrt[28] ), .B(new_n13842_), .ZN(new_n14131_));
  NOR2_X1    g13939(.A1(new_n14131_), .A2(new_n14129_), .ZN(new_n14132_));
  AOI22_X1   g13940(.A1(new_n14130_), .A2(\asqrt[28] ), .B1(new_n14128_), .B2(new_n14125_), .ZN(new_n14133_));
  INV_X1     g13941(.I(new_n13850_), .ZN(new_n14134_));
  OAI21_X1   g13942(.A1(new_n14133_), .A2(new_n7931_), .B(new_n14134_), .ZN(new_n14135_));
  NAND2_X1   g13943(.A1(new_n14135_), .A2(new_n14132_), .ZN(new_n14136_));
  OAI22_X1   g13944(.A1(new_n14133_), .A2(new_n7931_), .B1(new_n14131_), .B2(new_n14129_), .ZN(new_n14137_));
  AOI21_X1   g13945(.A1(new_n14137_), .A2(\asqrt[30] ), .B(new_n13857_), .ZN(new_n14138_));
  NOR2_X1    g13946(.A1(new_n14138_), .A2(new_n14136_), .ZN(new_n14139_));
  AOI22_X1   g13947(.A1(new_n14137_), .A2(\asqrt[30] ), .B1(new_n14135_), .B2(new_n14132_), .ZN(new_n14140_));
  INV_X1     g13948(.I(new_n13865_), .ZN(new_n14141_));
  OAI21_X1   g13949(.A1(new_n14140_), .A2(new_n7110_), .B(new_n14141_), .ZN(new_n14142_));
  NAND2_X1   g13950(.A1(new_n14142_), .A2(new_n14139_), .ZN(new_n14143_));
  OAI22_X1   g13951(.A1(new_n14140_), .A2(new_n7110_), .B1(new_n14138_), .B2(new_n14136_), .ZN(new_n14144_));
  AOI21_X1   g13952(.A1(new_n14144_), .A2(\asqrt[32] ), .B(new_n13872_), .ZN(new_n14145_));
  NOR2_X1    g13953(.A1(new_n14145_), .A2(new_n14143_), .ZN(new_n14146_));
  AOI22_X1   g13954(.A1(new_n14144_), .A2(\asqrt[32] ), .B1(new_n14142_), .B2(new_n14139_), .ZN(new_n14147_));
  INV_X1     g13955(.I(new_n13880_), .ZN(new_n14148_));
  OAI21_X1   g13956(.A1(new_n14147_), .A2(new_n6365_), .B(new_n14148_), .ZN(new_n14149_));
  NAND2_X1   g13957(.A1(new_n14149_), .A2(new_n14146_), .ZN(new_n14150_));
  OAI22_X1   g13958(.A1(new_n14147_), .A2(new_n6365_), .B1(new_n14145_), .B2(new_n14143_), .ZN(new_n14151_));
  AOI21_X1   g13959(.A1(new_n14151_), .A2(\asqrt[34] ), .B(new_n13887_), .ZN(new_n14152_));
  NOR2_X1    g13960(.A1(new_n14152_), .A2(new_n14150_), .ZN(new_n14153_));
  AOI22_X1   g13961(.A1(new_n14151_), .A2(\asqrt[34] ), .B1(new_n14149_), .B2(new_n14146_), .ZN(new_n14154_));
  INV_X1     g13962(.I(new_n13895_), .ZN(new_n14155_));
  OAI21_X1   g13963(.A1(new_n14154_), .A2(new_n5626_), .B(new_n14155_), .ZN(new_n14156_));
  NAND2_X1   g13964(.A1(new_n14156_), .A2(new_n14153_), .ZN(new_n14157_));
  OAI22_X1   g13965(.A1(new_n14154_), .A2(new_n5626_), .B1(new_n14152_), .B2(new_n14150_), .ZN(new_n14158_));
  AOI21_X1   g13966(.A1(new_n14158_), .A2(\asqrt[36] ), .B(new_n13902_), .ZN(new_n14159_));
  NOR2_X1    g13967(.A1(new_n14159_), .A2(new_n14157_), .ZN(new_n14160_));
  AOI22_X1   g13968(.A1(new_n14158_), .A2(\asqrt[36] ), .B1(new_n14156_), .B2(new_n14153_), .ZN(new_n14161_));
  INV_X1     g13969(.I(new_n13910_), .ZN(new_n14162_));
  OAI21_X1   g13970(.A1(new_n14161_), .A2(new_n4973_), .B(new_n14162_), .ZN(new_n14163_));
  NAND2_X1   g13971(.A1(new_n14163_), .A2(new_n14160_), .ZN(new_n14164_));
  OAI22_X1   g13972(.A1(new_n14161_), .A2(new_n4973_), .B1(new_n14159_), .B2(new_n14157_), .ZN(new_n14165_));
  AOI21_X1   g13973(.A1(new_n14165_), .A2(\asqrt[38] ), .B(new_n13917_), .ZN(new_n14166_));
  NOR2_X1    g13974(.A1(new_n14166_), .A2(new_n14164_), .ZN(new_n14167_));
  AOI22_X1   g13975(.A1(new_n14165_), .A2(\asqrt[38] ), .B1(new_n14163_), .B2(new_n14160_), .ZN(new_n14168_));
  INV_X1     g13976(.I(new_n13925_), .ZN(new_n14169_));
  OAI21_X1   g13977(.A1(new_n14168_), .A2(new_n4330_), .B(new_n14169_), .ZN(new_n14170_));
  NAND2_X1   g13978(.A1(new_n14170_), .A2(new_n14167_), .ZN(new_n14171_));
  OAI22_X1   g13979(.A1(new_n14168_), .A2(new_n4330_), .B1(new_n14166_), .B2(new_n14164_), .ZN(new_n14172_));
  AOI21_X1   g13980(.A1(new_n14172_), .A2(\asqrt[40] ), .B(new_n13932_), .ZN(new_n14173_));
  NOR2_X1    g13981(.A1(new_n14173_), .A2(new_n14171_), .ZN(new_n14174_));
  AOI22_X1   g13982(.A1(new_n14172_), .A2(\asqrt[40] ), .B1(new_n14170_), .B2(new_n14167_), .ZN(new_n14175_));
  INV_X1     g13983(.I(new_n13940_), .ZN(new_n14176_));
  OAI21_X1   g13984(.A1(new_n14175_), .A2(new_n3760_), .B(new_n14176_), .ZN(new_n14177_));
  NAND2_X1   g13985(.A1(new_n14177_), .A2(new_n14174_), .ZN(new_n14178_));
  OAI22_X1   g13986(.A1(new_n14175_), .A2(new_n3760_), .B1(new_n14173_), .B2(new_n14171_), .ZN(new_n14179_));
  AOI21_X1   g13987(.A1(new_n14179_), .A2(\asqrt[42] ), .B(new_n13947_), .ZN(new_n14180_));
  NOR2_X1    g13988(.A1(new_n14180_), .A2(new_n14178_), .ZN(new_n14181_));
  AOI22_X1   g13989(.A1(new_n14179_), .A2(\asqrt[42] ), .B1(new_n14177_), .B2(new_n14174_), .ZN(new_n14182_));
  INV_X1     g13990(.I(new_n13955_), .ZN(new_n14183_));
  OAI21_X1   g13991(.A1(new_n14182_), .A2(new_n3208_), .B(new_n14183_), .ZN(new_n14184_));
  NAND2_X1   g13992(.A1(new_n14184_), .A2(new_n14181_), .ZN(new_n14185_));
  OAI22_X1   g13993(.A1(new_n14182_), .A2(new_n3208_), .B1(new_n14180_), .B2(new_n14178_), .ZN(new_n14186_));
  AOI21_X1   g13994(.A1(new_n14186_), .A2(\asqrt[44] ), .B(new_n13962_), .ZN(new_n14187_));
  NOR2_X1    g13995(.A1(new_n14187_), .A2(new_n14185_), .ZN(new_n14188_));
  AOI22_X1   g13996(.A1(new_n14186_), .A2(\asqrt[44] ), .B1(new_n14184_), .B2(new_n14181_), .ZN(new_n14189_));
  INV_X1     g13997(.I(new_n13970_), .ZN(new_n14190_));
  OAI21_X1   g13998(.A1(new_n14189_), .A2(new_n2728_), .B(new_n14190_), .ZN(new_n14191_));
  NAND2_X1   g13999(.A1(new_n14191_), .A2(new_n14188_), .ZN(new_n14192_));
  OAI22_X1   g14000(.A1(new_n14189_), .A2(new_n2728_), .B1(new_n14187_), .B2(new_n14185_), .ZN(new_n14193_));
  AOI21_X1   g14001(.A1(new_n14193_), .A2(\asqrt[46] ), .B(new_n13977_), .ZN(new_n14194_));
  NOR2_X1    g14002(.A1(new_n14194_), .A2(new_n14192_), .ZN(new_n14195_));
  AOI22_X1   g14003(.A1(new_n14193_), .A2(\asqrt[46] ), .B1(new_n14191_), .B2(new_n14188_), .ZN(new_n14196_));
  INV_X1     g14004(.I(new_n13985_), .ZN(new_n14197_));
  OAI21_X1   g14005(.A1(new_n14196_), .A2(new_n2253_), .B(new_n14197_), .ZN(new_n14198_));
  NAND2_X1   g14006(.A1(new_n14198_), .A2(new_n14195_), .ZN(new_n14199_));
  OAI22_X1   g14007(.A1(new_n14196_), .A2(new_n2253_), .B1(new_n14194_), .B2(new_n14192_), .ZN(new_n14200_));
  AOI21_X1   g14008(.A1(new_n14200_), .A2(\asqrt[48] ), .B(new_n13992_), .ZN(new_n14201_));
  NOR2_X1    g14009(.A1(new_n14201_), .A2(new_n14199_), .ZN(new_n14202_));
  AOI22_X1   g14010(.A1(new_n14200_), .A2(\asqrt[48] ), .B1(new_n14198_), .B2(new_n14195_), .ZN(new_n14203_));
  INV_X1     g14011(.I(new_n14000_), .ZN(new_n14204_));
  OAI21_X1   g14012(.A1(new_n14203_), .A2(new_n1854_), .B(new_n14204_), .ZN(new_n14205_));
  NAND2_X1   g14013(.A1(new_n14205_), .A2(new_n14202_), .ZN(new_n14206_));
  OAI22_X1   g14014(.A1(new_n14203_), .A2(new_n1854_), .B1(new_n14201_), .B2(new_n14199_), .ZN(new_n14207_));
  AOI21_X1   g14015(.A1(new_n14207_), .A2(\asqrt[50] ), .B(new_n14007_), .ZN(new_n14208_));
  NOR2_X1    g14016(.A1(new_n14208_), .A2(new_n14206_), .ZN(new_n14209_));
  AOI22_X1   g14017(.A1(new_n14207_), .A2(\asqrt[50] ), .B1(new_n14205_), .B2(new_n14202_), .ZN(new_n14210_));
  INV_X1     g14018(.I(new_n14015_), .ZN(new_n14211_));
  OAI21_X1   g14019(.A1(new_n14210_), .A2(new_n1436_), .B(new_n14211_), .ZN(new_n14212_));
  NAND2_X1   g14020(.A1(new_n14212_), .A2(new_n14209_), .ZN(new_n14213_));
  OAI22_X1   g14021(.A1(new_n14210_), .A2(new_n1436_), .B1(new_n14208_), .B2(new_n14206_), .ZN(new_n14214_));
  AOI21_X1   g14022(.A1(new_n14214_), .A2(\asqrt[52] ), .B(new_n14021_), .ZN(new_n14215_));
  NOR2_X1    g14023(.A1(new_n14215_), .A2(new_n14213_), .ZN(new_n14216_));
  AOI22_X1   g14024(.A1(new_n14214_), .A2(\asqrt[52] ), .B1(new_n14212_), .B2(new_n14209_), .ZN(new_n14217_));
  INV_X1     g14025(.I(new_n14028_), .ZN(new_n14218_));
  OAI21_X1   g14026(.A1(new_n14217_), .A2(new_n1096_), .B(new_n14218_), .ZN(new_n14219_));
  NAND2_X1   g14027(.A1(new_n14219_), .A2(new_n14216_), .ZN(new_n14220_));
  OAI22_X1   g14028(.A1(new_n14217_), .A2(new_n1096_), .B1(new_n14215_), .B2(new_n14213_), .ZN(new_n14221_));
  AOI21_X1   g14029(.A1(new_n14221_), .A2(\asqrt[54] ), .B(new_n14034_), .ZN(new_n14222_));
  NOR2_X1    g14030(.A1(new_n14222_), .A2(new_n14220_), .ZN(new_n14223_));
  AOI22_X1   g14031(.A1(new_n14221_), .A2(\asqrt[54] ), .B1(new_n14219_), .B2(new_n14216_), .ZN(new_n14224_));
  INV_X1     g14032(.I(new_n14041_), .ZN(new_n14225_));
  OAI21_X1   g14033(.A1(new_n14224_), .A2(new_n825_), .B(new_n14225_), .ZN(new_n14226_));
  NAND2_X1   g14034(.A1(new_n14226_), .A2(new_n14223_), .ZN(new_n14227_));
  OAI22_X1   g14035(.A1(new_n14224_), .A2(new_n825_), .B1(new_n14222_), .B2(new_n14220_), .ZN(new_n14228_));
  AOI21_X1   g14036(.A1(new_n14228_), .A2(\asqrt[56] ), .B(new_n14047_), .ZN(new_n14229_));
  NOR2_X1    g14037(.A1(new_n14229_), .A2(new_n14227_), .ZN(new_n14230_));
  AOI22_X1   g14038(.A1(new_n14228_), .A2(\asqrt[56] ), .B1(new_n14226_), .B2(new_n14223_), .ZN(new_n14231_));
  INV_X1     g14039(.I(new_n14054_), .ZN(new_n14232_));
  OAI21_X1   g14040(.A1(new_n14231_), .A2(new_n587_), .B(new_n14232_), .ZN(new_n14233_));
  NAND2_X1   g14041(.A1(new_n14233_), .A2(new_n14230_), .ZN(new_n14234_));
  OAI22_X1   g14042(.A1(new_n14231_), .A2(new_n587_), .B1(new_n14229_), .B2(new_n14227_), .ZN(new_n14235_));
  AOI21_X1   g14043(.A1(new_n14235_), .A2(\asqrt[58] ), .B(new_n14060_), .ZN(new_n14236_));
  NOR2_X1    g14044(.A1(new_n14236_), .A2(new_n14234_), .ZN(new_n14237_));
  AOI22_X1   g14045(.A1(new_n14235_), .A2(\asqrt[58] ), .B1(new_n14233_), .B2(new_n14230_), .ZN(new_n14238_));
  INV_X1     g14046(.I(new_n14067_), .ZN(new_n14239_));
  OAI21_X1   g14047(.A1(new_n14238_), .A2(new_n376_), .B(new_n14239_), .ZN(new_n14240_));
  NAND2_X1   g14048(.A1(new_n14240_), .A2(new_n14237_), .ZN(new_n14241_));
  OAI22_X1   g14049(.A1(new_n14238_), .A2(new_n376_), .B1(new_n14236_), .B2(new_n14234_), .ZN(new_n14242_));
  AOI21_X1   g14050(.A1(new_n14242_), .A2(\asqrt[60] ), .B(new_n14073_), .ZN(new_n14243_));
  AOI22_X1   g14051(.A1(new_n14242_), .A2(\asqrt[60] ), .B1(new_n14240_), .B2(new_n14237_), .ZN(new_n14244_));
  OAI22_X1   g14052(.A1(new_n14244_), .A2(new_n229_), .B1(new_n14243_), .B2(new_n14241_), .ZN(new_n14245_));
  NOR4_X1    g14053(.A1(new_n14245_), .A2(\asqrt[62] ), .A3(new_n13727_), .A4(new_n13731_), .ZN(new_n14246_));
  NAND2_X1   g14054(.A1(new_n13747_), .A2(new_n13154_), .ZN(new_n14247_));
  XOR2_X1    g14055(.A1(new_n13747_), .A2(\asqrt[63] ), .Z(new_n14248_));
  AOI21_X1   g14056(.A1(\asqrt[17] ), .A2(new_n14247_), .B(new_n14248_), .ZN(new_n14249_));
  NAND2_X1   g14057(.A1(new_n14246_), .A2(new_n14249_), .ZN(new_n14250_));
  NOR4_X1    g14058(.A1(new_n14250_), .A2(new_n13707_), .A3(new_n14086_), .A4(new_n13715_), .ZN(new_n14251_));
  NOR2_X1    g14059(.A1(new_n13707_), .A2(\a[32] ), .ZN(new_n14252_));
  OAI21_X1   g14060(.A1(new_n14251_), .A2(new_n14252_), .B(new_n13706_), .ZN(new_n14253_));
  INV_X1     g14061(.I(new_n13706_), .ZN(new_n14254_));
  INV_X1     g14062(.I(new_n13715_), .ZN(new_n14255_));
  NOR2_X1    g14063(.A1(new_n14243_), .A2(new_n14241_), .ZN(new_n14256_));
  NOR3_X1    g14064(.A1(new_n14244_), .A2(new_n229_), .A3(new_n14079_), .ZN(new_n14257_));
  AOI21_X1   g14065(.A1(new_n14257_), .A2(new_n14256_), .B(new_n13732_), .ZN(new_n14258_));
  AOI21_X1   g14066(.A1(new_n14258_), .A2(new_n14084_), .B(new_n13727_), .ZN(new_n14259_));
  AOI22_X1   g14067(.A1(new_n14077_), .A2(\asqrt[61] ), .B1(new_n14075_), .B2(new_n14069_), .ZN(new_n14260_));
  NAND4_X1   g14068(.A1(new_n14260_), .A2(new_n196_), .A3(new_n13728_), .A4(new_n14078_), .ZN(new_n14261_));
  INV_X1     g14069(.I(new_n14249_), .ZN(new_n14262_));
  NOR2_X1    g14070(.A1(new_n14261_), .A2(new_n14262_), .ZN(new_n14263_));
  NAND4_X1   g14071(.A1(new_n14263_), .A2(new_n14259_), .A3(\a[33] ), .A4(new_n14255_), .ZN(new_n14264_));
  NAND3_X1   g14072(.A1(new_n14264_), .A2(\a[32] ), .A3(new_n14254_), .ZN(new_n14265_));
  NAND2_X1   g14073(.A1(new_n14253_), .A2(new_n14265_), .ZN(new_n14266_));
  NOR2_X1    g14074(.A1(new_n14250_), .A2(new_n14086_), .ZN(new_n14267_));
  NOR4_X1    g14075(.A1(new_n13713_), .A2(new_n13154_), .A3(new_n13762_), .A4(new_n13699_), .ZN(new_n14268_));
  NAND2_X1   g14076(.A1(\asqrt[17] ), .A2(\a[32] ), .ZN(new_n14269_));
  XOR2_X1    g14077(.A1(new_n14269_), .A2(new_n14268_), .Z(new_n14270_));
  NOR2_X1    g14078(.A1(new_n14270_), .A2(new_n13703_), .ZN(new_n14271_));
  INV_X1     g14079(.I(new_n14271_), .ZN(new_n14272_));
  NAND3_X1   g14080(.A1(new_n14263_), .A2(new_n14259_), .A3(new_n14255_), .ZN(new_n14273_));
  NAND2_X1   g14081(.A1(new_n14038_), .A2(\asqrt[55] ), .ZN(new_n14274_));
  AOI21_X1   g14082(.A1(new_n14274_), .A2(new_n14037_), .B(new_n724_), .ZN(new_n14275_));
  OAI21_X1   g14083(.A1(new_n14043_), .A2(new_n14275_), .B(\asqrt[57] ), .ZN(new_n14276_));
  AOI21_X1   g14084(.A1(new_n14050_), .A2(new_n14276_), .B(new_n504_), .ZN(new_n14277_));
  OAI21_X1   g14085(.A1(new_n14056_), .A2(new_n14277_), .B(\asqrt[59] ), .ZN(new_n14278_));
  AOI21_X1   g14086(.A1(new_n14063_), .A2(new_n14278_), .B(new_n275_), .ZN(new_n14279_));
  OAI21_X1   g14087(.A1(new_n14069_), .A2(new_n14279_), .B(\asqrt[61] ), .ZN(new_n14280_));
  NOR3_X1    g14088(.A1(new_n14076_), .A2(new_n14280_), .A3(new_n14079_), .ZN(new_n14281_));
  NOR3_X1    g14089(.A1(new_n14281_), .A2(new_n13732_), .A3(new_n14085_), .ZN(new_n14282_));
  OAI21_X1   g14090(.A1(new_n14282_), .A2(new_n13727_), .B(new_n14261_), .ZN(new_n14283_));
  NOR2_X1    g14091(.A1(new_n14255_), .A2(new_n14249_), .ZN(new_n14284_));
  NAND2_X1   g14092(.A1(new_n14284_), .A2(\asqrt[17] ), .ZN(new_n14285_));
  OAI21_X1   g14093(.A1(new_n14283_), .A2(new_n14285_), .B(new_n13734_), .ZN(new_n14286_));
  NAND3_X1   g14094(.A1(new_n14286_), .A2(new_n13735_), .A3(new_n14273_), .ZN(new_n14287_));
  NOR3_X1    g14095(.A1(new_n14250_), .A2(new_n13715_), .A3(new_n14086_), .ZN(\asqrt[16] ));
  NAND2_X1   g14096(.A1(new_n14228_), .A2(\asqrt[56] ), .ZN(new_n14289_));
  AOI21_X1   g14097(.A1(new_n14289_), .A2(new_n14227_), .B(new_n587_), .ZN(new_n14290_));
  OAI21_X1   g14098(.A1(new_n14230_), .A2(new_n14290_), .B(\asqrt[58] ), .ZN(new_n14291_));
  AOI21_X1   g14099(.A1(new_n14234_), .A2(new_n14291_), .B(new_n376_), .ZN(new_n14292_));
  OAI21_X1   g14100(.A1(new_n14237_), .A2(new_n14292_), .B(\asqrt[60] ), .ZN(new_n14293_));
  AOI21_X1   g14101(.A1(new_n14241_), .A2(new_n14293_), .B(new_n229_), .ZN(new_n14294_));
  NAND4_X1   g14102(.A1(new_n14294_), .A2(new_n14069_), .A3(new_n14075_), .A4(new_n14080_), .ZN(new_n14295_));
  NAND3_X1   g14103(.A1(new_n14295_), .A2(new_n13733_), .A3(new_n14084_), .ZN(new_n14296_));
  AOI21_X1   g14104(.A1(new_n13728_), .A2(new_n14296_), .B(new_n14246_), .ZN(new_n14297_));
  INV_X1     g14105(.I(new_n14285_), .ZN(new_n14298_));
  AOI21_X1   g14106(.A1(new_n14297_), .A2(new_n14298_), .B(\a[34] ), .ZN(new_n14299_));
  OAI21_X1   g14107(.A1(new_n14299_), .A2(new_n13736_), .B(\asqrt[16] ), .ZN(new_n14300_));
  NAND4_X1   g14108(.A1(new_n14300_), .A2(new_n14287_), .A3(new_n13192_), .A4(new_n14272_), .ZN(new_n14301_));
  NAND2_X1   g14109(.A1(new_n14301_), .A2(new_n14266_), .ZN(new_n14302_));
  NAND3_X1   g14110(.A1(new_n14253_), .A2(new_n14265_), .A3(new_n14272_), .ZN(new_n14303_));
  AOI21_X1   g14111(.A1(\asqrt[17] ), .A2(new_n13734_), .B(\a[35] ), .ZN(new_n14304_));
  NOR2_X1    g14112(.A1(new_n13751_), .A2(\a[34] ), .ZN(new_n14305_));
  AOI21_X1   g14113(.A1(\asqrt[17] ), .A2(\a[34] ), .B(new_n13738_), .ZN(new_n14306_));
  OAI21_X1   g14114(.A1(new_n14305_), .A2(new_n14304_), .B(new_n14306_), .ZN(new_n14307_));
  INV_X1     g14115(.I(new_n14307_), .ZN(new_n14308_));
  NAND3_X1   g14116(.A1(\asqrt[16] ), .A2(new_n13759_), .A3(new_n14308_), .ZN(new_n14309_));
  OAI21_X1   g14117(.A1(new_n14273_), .A2(new_n14307_), .B(new_n13758_), .ZN(new_n14310_));
  NAND3_X1   g14118(.A1(new_n14309_), .A2(new_n14310_), .A3(new_n12657_), .ZN(new_n14311_));
  AOI21_X1   g14119(.A1(new_n14303_), .A2(\asqrt[18] ), .B(new_n14311_), .ZN(new_n14312_));
  NOR2_X1    g14120(.A1(new_n14302_), .A2(new_n14312_), .ZN(new_n14313_));
  NAND2_X1   g14121(.A1(new_n14303_), .A2(\asqrt[18] ), .ZN(new_n14314_));
  AOI21_X1   g14122(.A1(new_n14302_), .A2(new_n14314_), .B(new_n12657_), .ZN(new_n14315_));
  NAND2_X1   g14123(.A1(new_n13773_), .A2(\asqrt[19] ), .ZN(new_n14316_));
  INV_X1     g14124(.I(new_n14316_), .ZN(new_n14317_));
  NAND2_X1   g14125(.A1(new_n13767_), .A2(new_n13770_), .ZN(new_n14318_));
  NAND3_X1   g14126(.A1(new_n14318_), .A2(new_n14095_), .A3(new_n12657_), .ZN(new_n14319_));
  NOR3_X1    g14127(.A1(new_n14273_), .A2(new_n14317_), .A3(new_n14319_), .ZN(new_n14320_));
  NOR2_X1    g14128(.A1(new_n14273_), .A2(new_n14319_), .ZN(new_n14321_));
  NOR2_X1    g14129(.A1(new_n14321_), .A2(new_n14316_), .ZN(new_n14322_));
  NOR3_X1    g14130(.A1(new_n14322_), .A2(\asqrt[20] ), .A3(new_n14320_), .ZN(new_n14323_));
  INV_X1     g14131(.I(new_n14323_), .ZN(new_n14324_));
  OAI21_X1   g14132(.A1(new_n14315_), .A2(new_n14324_), .B(new_n14313_), .ZN(new_n14325_));
  OAI21_X1   g14133(.A1(new_n14315_), .A2(new_n14313_), .B(\asqrt[20] ), .ZN(new_n14326_));
  NAND2_X1   g14134(.A1(new_n14101_), .A2(\asqrt[20] ), .ZN(new_n14327_));
  NOR2_X1    g14135(.A1(new_n14097_), .A2(new_n14096_), .ZN(new_n14328_));
  NOR4_X1    g14136(.A1(new_n14273_), .A2(\asqrt[20] ), .A3(new_n14328_), .A4(new_n14101_), .ZN(new_n14329_));
  XOR2_X1    g14137(.A1(new_n14329_), .A2(new_n14327_), .Z(new_n14330_));
  NAND2_X1   g14138(.A1(new_n14330_), .A2(new_n11631_), .ZN(new_n14331_));
  INV_X1     g14139(.I(new_n14331_), .ZN(new_n14332_));
  AOI21_X1   g14140(.A1(new_n14326_), .A2(new_n14332_), .B(new_n14325_), .ZN(new_n14333_));
  AOI21_X1   g14141(.A1(new_n14325_), .A2(new_n14326_), .B(new_n11631_), .ZN(new_n14334_));
  NAND2_X1   g14142(.A1(new_n13791_), .A2(\asqrt[21] ), .ZN(new_n14335_));
  NOR2_X1    g14143(.A1(new_n13786_), .A2(new_n13787_), .ZN(new_n14336_));
  NOR4_X1    g14144(.A1(new_n14273_), .A2(\asqrt[21] ), .A3(new_n14336_), .A4(new_n13791_), .ZN(new_n14337_));
  XOR2_X1    g14145(.A1(new_n14337_), .A2(new_n14335_), .Z(new_n14338_));
  NAND2_X1   g14146(.A1(new_n14338_), .A2(new_n11105_), .ZN(new_n14339_));
  OAI21_X1   g14147(.A1(new_n14334_), .A2(new_n14339_), .B(new_n14333_), .ZN(new_n14340_));
  OAI21_X1   g14148(.A1(new_n14333_), .A2(new_n14334_), .B(\asqrt[22] ), .ZN(new_n14341_));
  NOR4_X1    g14149(.A1(new_n14273_), .A2(\asqrt[22] ), .A3(new_n13794_), .A4(new_n14109_), .ZN(new_n14342_));
  AOI21_X1   g14150(.A1(new_n14335_), .A2(new_n13790_), .B(new_n11105_), .ZN(new_n14343_));
  NOR2_X1    g14151(.A1(new_n14342_), .A2(new_n14343_), .ZN(new_n14344_));
  NAND2_X1   g14152(.A1(new_n14344_), .A2(new_n10614_), .ZN(new_n14345_));
  INV_X1     g14153(.I(new_n14345_), .ZN(new_n14346_));
  AOI21_X1   g14154(.A1(new_n14341_), .A2(new_n14346_), .B(new_n14340_), .ZN(new_n14347_));
  AOI22_X1   g14155(.A1(new_n14301_), .A2(new_n14266_), .B1(\asqrt[18] ), .B2(new_n14303_), .ZN(new_n14348_));
  OAI21_X1   g14156(.A1(new_n14348_), .A2(new_n12657_), .B(new_n14323_), .ZN(new_n14349_));
  OAI22_X1   g14157(.A1(new_n14348_), .A2(new_n12657_), .B1(new_n14302_), .B2(new_n14312_), .ZN(new_n14350_));
  AOI22_X1   g14158(.A1(new_n14350_), .A2(\asqrt[20] ), .B1(new_n14349_), .B2(new_n14313_), .ZN(new_n14351_));
  INV_X1     g14159(.I(new_n14339_), .ZN(new_n14352_));
  OAI21_X1   g14160(.A1(new_n14351_), .A2(new_n11631_), .B(new_n14352_), .ZN(new_n14353_));
  AOI21_X1   g14161(.A1(new_n14350_), .A2(\asqrt[20] ), .B(new_n14331_), .ZN(new_n14354_));
  OAI22_X1   g14162(.A1(new_n14351_), .A2(new_n11631_), .B1(new_n14354_), .B2(new_n14325_), .ZN(new_n14355_));
  AOI22_X1   g14163(.A1(new_n14355_), .A2(\asqrt[22] ), .B1(new_n14353_), .B2(new_n14333_), .ZN(new_n14356_));
  NAND2_X1   g14164(.A1(new_n13805_), .A2(\asqrt[23] ), .ZN(new_n14357_));
  NOR4_X1    g14165(.A1(new_n14273_), .A2(\asqrt[23] ), .A3(new_n13800_), .A4(new_n13805_), .ZN(new_n14358_));
  XOR2_X1    g14166(.A1(new_n14358_), .A2(new_n14357_), .Z(new_n14359_));
  NAND2_X1   g14167(.A1(new_n14359_), .A2(new_n10104_), .ZN(new_n14360_));
  INV_X1     g14168(.I(new_n14360_), .ZN(new_n14361_));
  OAI21_X1   g14169(.A1(new_n14356_), .A2(new_n10614_), .B(new_n14361_), .ZN(new_n14362_));
  NAND2_X1   g14170(.A1(new_n14362_), .A2(new_n14347_), .ZN(new_n14363_));
  AOI21_X1   g14171(.A1(new_n14355_), .A2(\asqrt[22] ), .B(new_n14345_), .ZN(new_n14364_));
  OAI22_X1   g14172(.A1(new_n14356_), .A2(new_n10614_), .B1(new_n14364_), .B2(new_n14340_), .ZN(new_n14365_));
  NOR4_X1    g14173(.A1(new_n14273_), .A2(\asqrt[24] ), .A3(new_n13807_), .A4(new_n14116_), .ZN(new_n14366_));
  AOI21_X1   g14174(.A1(new_n14357_), .A2(new_n13804_), .B(new_n10104_), .ZN(new_n14367_));
  NOR2_X1    g14175(.A1(new_n14366_), .A2(new_n14367_), .ZN(new_n14368_));
  NAND2_X1   g14176(.A1(new_n14368_), .A2(new_n9672_), .ZN(new_n14369_));
  AOI21_X1   g14177(.A1(new_n14365_), .A2(\asqrt[24] ), .B(new_n14369_), .ZN(new_n14370_));
  NOR2_X1    g14178(.A1(new_n14370_), .A2(new_n14363_), .ZN(new_n14371_));
  AOI22_X1   g14179(.A1(new_n14365_), .A2(\asqrt[24] ), .B1(new_n14362_), .B2(new_n14347_), .ZN(new_n14372_));
  NAND2_X1   g14180(.A1(new_n13818_), .A2(\asqrt[25] ), .ZN(new_n14373_));
  NOR4_X1    g14181(.A1(new_n14273_), .A2(\asqrt[25] ), .A3(new_n13813_), .A4(new_n13818_), .ZN(new_n14374_));
  XOR2_X1    g14182(.A1(new_n14374_), .A2(new_n14373_), .Z(new_n14375_));
  NAND2_X1   g14183(.A1(new_n14375_), .A2(new_n9212_), .ZN(new_n14376_));
  INV_X1     g14184(.I(new_n14376_), .ZN(new_n14377_));
  OAI21_X1   g14185(.A1(new_n14372_), .A2(new_n9672_), .B(new_n14377_), .ZN(new_n14378_));
  NAND2_X1   g14186(.A1(new_n14378_), .A2(new_n14371_), .ZN(new_n14379_));
  OAI22_X1   g14187(.A1(new_n14372_), .A2(new_n9672_), .B1(new_n14370_), .B2(new_n14363_), .ZN(new_n14380_));
  NOR4_X1    g14188(.A1(new_n14273_), .A2(\asqrt[26] ), .A3(new_n13820_), .A4(new_n14123_), .ZN(new_n14381_));
  AOI21_X1   g14189(.A1(new_n14373_), .A2(new_n13817_), .B(new_n9212_), .ZN(new_n14382_));
  NOR2_X1    g14190(.A1(new_n14381_), .A2(new_n14382_), .ZN(new_n14383_));
  NAND2_X1   g14191(.A1(new_n14383_), .A2(new_n8763_), .ZN(new_n14384_));
  AOI21_X1   g14192(.A1(new_n14380_), .A2(\asqrt[26] ), .B(new_n14384_), .ZN(new_n14385_));
  NOR2_X1    g14193(.A1(new_n14385_), .A2(new_n14379_), .ZN(new_n14386_));
  AOI22_X1   g14194(.A1(new_n14380_), .A2(\asqrt[26] ), .B1(new_n14378_), .B2(new_n14371_), .ZN(new_n14387_));
  NAND2_X1   g14195(.A1(new_n13831_), .A2(\asqrt[27] ), .ZN(new_n14388_));
  NOR4_X1    g14196(.A1(new_n14273_), .A2(\asqrt[27] ), .A3(new_n13826_), .A4(new_n13831_), .ZN(new_n14389_));
  XOR2_X1    g14197(.A1(new_n14389_), .A2(new_n14388_), .Z(new_n14390_));
  NAND2_X1   g14198(.A1(new_n14390_), .A2(new_n8319_), .ZN(new_n14391_));
  INV_X1     g14199(.I(new_n14391_), .ZN(new_n14392_));
  OAI21_X1   g14200(.A1(new_n14387_), .A2(new_n8763_), .B(new_n14392_), .ZN(new_n14393_));
  NAND2_X1   g14201(.A1(new_n14393_), .A2(new_n14386_), .ZN(new_n14394_));
  OAI22_X1   g14202(.A1(new_n14387_), .A2(new_n8763_), .B1(new_n14385_), .B2(new_n14379_), .ZN(new_n14395_));
  NAND2_X1   g14203(.A1(new_n14130_), .A2(\asqrt[28] ), .ZN(new_n14396_));
  NOR4_X1    g14204(.A1(new_n14273_), .A2(\asqrt[28] ), .A3(new_n13834_), .A4(new_n14130_), .ZN(new_n14397_));
  XOR2_X1    g14205(.A1(new_n14397_), .A2(new_n14396_), .Z(new_n14398_));
  NAND2_X1   g14206(.A1(new_n14398_), .A2(new_n7931_), .ZN(new_n14399_));
  AOI21_X1   g14207(.A1(new_n14395_), .A2(\asqrt[28] ), .B(new_n14399_), .ZN(new_n14400_));
  NOR2_X1    g14208(.A1(new_n14400_), .A2(new_n14394_), .ZN(new_n14401_));
  AOI22_X1   g14209(.A1(new_n14395_), .A2(\asqrt[28] ), .B1(new_n14393_), .B2(new_n14386_), .ZN(new_n14402_));
  NOR4_X1    g14210(.A1(new_n14273_), .A2(\asqrt[29] ), .A3(new_n13841_), .A4(new_n13846_), .ZN(new_n14403_));
  AOI21_X1   g14211(.A1(new_n14396_), .A2(new_n14129_), .B(new_n7931_), .ZN(new_n14404_));
  NOR2_X1    g14212(.A1(new_n14403_), .A2(new_n14404_), .ZN(new_n14405_));
  NAND2_X1   g14213(.A1(new_n14405_), .A2(new_n7517_), .ZN(new_n14406_));
  INV_X1     g14214(.I(new_n14406_), .ZN(new_n14407_));
  OAI21_X1   g14215(.A1(new_n14402_), .A2(new_n7931_), .B(new_n14407_), .ZN(new_n14408_));
  NAND2_X1   g14216(.A1(new_n14408_), .A2(new_n14401_), .ZN(new_n14409_));
  OAI22_X1   g14217(.A1(new_n14402_), .A2(new_n7931_), .B1(new_n14400_), .B2(new_n14394_), .ZN(new_n14410_));
  NAND2_X1   g14218(.A1(new_n14137_), .A2(\asqrt[30] ), .ZN(new_n14411_));
  NOR4_X1    g14219(.A1(new_n14273_), .A2(\asqrt[30] ), .A3(new_n13849_), .A4(new_n14137_), .ZN(new_n14412_));
  XOR2_X1    g14220(.A1(new_n14412_), .A2(new_n14411_), .Z(new_n14413_));
  NAND2_X1   g14221(.A1(new_n14413_), .A2(new_n7110_), .ZN(new_n14414_));
  AOI21_X1   g14222(.A1(new_n14410_), .A2(\asqrt[30] ), .B(new_n14414_), .ZN(new_n14415_));
  NOR2_X1    g14223(.A1(new_n14415_), .A2(new_n14409_), .ZN(new_n14416_));
  AOI22_X1   g14224(.A1(new_n14410_), .A2(\asqrt[30] ), .B1(new_n14408_), .B2(new_n14401_), .ZN(new_n14417_));
  NOR4_X1    g14225(.A1(new_n14273_), .A2(\asqrt[31] ), .A3(new_n13856_), .A4(new_n13861_), .ZN(new_n14418_));
  AOI21_X1   g14226(.A1(new_n14411_), .A2(new_n14136_), .B(new_n7110_), .ZN(new_n14419_));
  NOR2_X1    g14227(.A1(new_n14418_), .A2(new_n14419_), .ZN(new_n14420_));
  NAND2_X1   g14228(.A1(new_n14420_), .A2(new_n6708_), .ZN(new_n14421_));
  INV_X1     g14229(.I(new_n14421_), .ZN(new_n14422_));
  OAI21_X1   g14230(.A1(new_n14417_), .A2(new_n7110_), .B(new_n14422_), .ZN(new_n14423_));
  NAND2_X1   g14231(.A1(new_n14423_), .A2(new_n14416_), .ZN(new_n14424_));
  OAI22_X1   g14232(.A1(new_n14417_), .A2(new_n7110_), .B1(new_n14415_), .B2(new_n14409_), .ZN(new_n14425_));
  NAND2_X1   g14233(.A1(new_n14144_), .A2(\asqrt[32] ), .ZN(new_n14426_));
  NOR4_X1    g14234(.A1(new_n14273_), .A2(\asqrt[32] ), .A3(new_n13864_), .A4(new_n14144_), .ZN(new_n14427_));
  XOR2_X1    g14235(.A1(new_n14427_), .A2(new_n14426_), .Z(new_n14428_));
  NAND2_X1   g14236(.A1(new_n14428_), .A2(new_n6365_), .ZN(new_n14429_));
  AOI21_X1   g14237(.A1(new_n14425_), .A2(\asqrt[32] ), .B(new_n14429_), .ZN(new_n14430_));
  NOR2_X1    g14238(.A1(new_n14430_), .A2(new_n14424_), .ZN(new_n14431_));
  AOI22_X1   g14239(.A1(new_n14425_), .A2(\asqrt[32] ), .B1(new_n14423_), .B2(new_n14416_), .ZN(new_n14432_));
  NOR4_X1    g14240(.A1(new_n14273_), .A2(\asqrt[33] ), .A3(new_n13871_), .A4(new_n13876_), .ZN(new_n14433_));
  AOI21_X1   g14241(.A1(new_n14426_), .A2(new_n14143_), .B(new_n6365_), .ZN(new_n14434_));
  NOR2_X1    g14242(.A1(new_n14433_), .A2(new_n14434_), .ZN(new_n14435_));
  NAND2_X1   g14243(.A1(new_n14435_), .A2(new_n5991_), .ZN(new_n14436_));
  INV_X1     g14244(.I(new_n14436_), .ZN(new_n14437_));
  OAI21_X1   g14245(.A1(new_n14432_), .A2(new_n6365_), .B(new_n14437_), .ZN(new_n14438_));
  NAND2_X1   g14246(.A1(new_n14438_), .A2(new_n14431_), .ZN(new_n14439_));
  OAI22_X1   g14247(.A1(new_n14432_), .A2(new_n6365_), .B1(new_n14430_), .B2(new_n14424_), .ZN(new_n14440_));
  NAND2_X1   g14248(.A1(new_n14151_), .A2(\asqrt[34] ), .ZN(new_n14441_));
  NOR4_X1    g14249(.A1(new_n14273_), .A2(\asqrt[34] ), .A3(new_n13879_), .A4(new_n14151_), .ZN(new_n14442_));
  XOR2_X1    g14250(.A1(new_n14442_), .A2(new_n14441_), .Z(new_n14443_));
  NAND2_X1   g14251(.A1(new_n14443_), .A2(new_n5626_), .ZN(new_n14444_));
  AOI21_X1   g14252(.A1(new_n14440_), .A2(\asqrt[34] ), .B(new_n14444_), .ZN(new_n14445_));
  NOR2_X1    g14253(.A1(new_n14445_), .A2(new_n14439_), .ZN(new_n14446_));
  AOI22_X1   g14254(.A1(new_n14440_), .A2(\asqrt[34] ), .B1(new_n14438_), .B2(new_n14431_), .ZN(new_n14447_));
  NOR4_X1    g14255(.A1(new_n14273_), .A2(\asqrt[35] ), .A3(new_n13886_), .A4(new_n13891_), .ZN(new_n14448_));
  AOI21_X1   g14256(.A1(new_n14441_), .A2(new_n14150_), .B(new_n5626_), .ZN(new_n14449_));
  NOR2_X1    g14257(.A1(new_n14448_), .A2(new_n14449_), .ZN(new_n14450_));
  NAND2_X1   g14258(.A1(new_n14450_), .A2(new_n5273_), .ZN(new_n14451_));
  INV_X1     g14259(.I(new_n14451_), .ZN(new_n14452_));
  OAI21_X1   g14260(.A1(new_n14447_), .A2(new_n5626_), .B(new_n14452_), .ZN(new_n14453_));
  NAND2_X1   g14261(.A1(new_n14453_), .A2(new_n14446_), .ZN(new_n14454_));
  OAI22_X1   g14262(.A1(new_n14447_), .A2(new_n5626_), .B1(new_n14445_), .B2(new_n14439_), .ZN(new_n14455_));
  NAND2_X1   g14263(.A1(new_n14158_), .A2(\asqrt[36] ), .ZN(new_n14456_));
  NOR4_X1    g14264(.A1(new_n14273_), .A2(\asqrt[36] ), .A3(new_n13894_), .A4(new_n14158_), .ZN(new_n14457_));
  XOR2_X1    g14265(.A1(new_n14457_), .A2(new_n14456_), .Z(new_n14458_));
  NAND2_X1   g14266(.A1(new_n14458_), .A2(new_n4973_), .ZN(new_n14459_));
  AOI21_X1   g14267(.A1(new_n14455_), .A2(\asqrt[36] ), .B(new_n14459_), .ZN(new_n14460_));
  NOR2_X1    g14268(.A1(new_n14460_), .A2(new_n14454_), .ZN(new_n14461_));
  AOI22_X1   g14269(.A1(new_n14455_), .A2(\asqrt[36] ), .B1(new_n14453_), .B2(new_n14446_), .ZN(new_n14462_));
  NAND2_X1   g14270(.A1(new_n13906_), .A2(\asqrt[37] ), .ZN(new_n14463_));
  NOR4_X1    g14271(.A1(new_n14273_), .A2(\asqrt[37] ), .A3(new_n13901_), .A4(new_n13906_), .ZN(new_n14464_));
  XOR2_X1    g14272(.A1(new_n14464_), .A2(new_n14463_), .Z(new_n14465_));
  NAND2_X1   g14273(.A1(new_n14465_), .A2(new_n4645_), .ZN(new_n14466_));
  INV_X1     g14274(.I(new_n14466_), .ZN(new_n14467_));
  OAI21_X1   g14275(.A1(new_n14462_), .A2(new_n4973_), .B(new_n14467_), .ZN(new_n14468_));
  NAND2_X1   g14276(.A1(new_n14468_), .A2(new_n14461_), .ZN(new_n14469_));
  OAI22_X1   g14277(.A1(new_n14462_), .A2(new_n4973_), .B1(new_n14460_), .B2(new_n14454_), .ZN(new_n14470_));
  NOR4_X1    g14278(.A1(new_n14273_), .A2(\asqrt[38] ), .A3(new_n13909_), .A4(new_n14165_), .ZN(new_n14471_));
  AOI21_X1   g14279(.A1(new_n14463_), .A2(new_n13905_), .B(new_n4645_), .ZN(new_n14472_));
  NOR2_X1    g14280(.A1(new_n14471_), .A2(new_n14472_), .ZN(new_n14473_));
  NAND2_X1   g14281(.A1(new_n14473_), .A2(new_n4330_), .ZN(new_n14474_));
  AOI21_X1   g14282(.A1(new_n14470_), .A2(\asqrt[38] ), .B(new_n14474_), .ZN(new_n14475_));
  NOR2_X1    g14283(.A1(new_n14475_), .A2(new_n14469_), .ZN(new_n14476_));
  AOI22_X1   g14284(.A1(new_n14470_), .A2(\asqrt[38] ), .B1(new_n14468_), .B2(new_n14461_), .ZN(new_n14477_));
  NAND2_X1   g14285(.A1(new_n13921_), .A2(\asqrt[39] ), .ZN(new_n14478_));
  NOR4_X1    g14286(.A1(new_n14273_), .A2(\asqrt[39] ), .A3(new_n13916_), .A4(new_n13921_), .ZN(new_n14479_));
  XOR2_X1    g14287(.A1(new_n14479_), .A2(new_n14478_), .Z(new_n14480_));
  NAND2_X1   g14288(.A1(new_n14480_), .A2(new_n4018_), .ZN(new_n14481_));
  INV_X1     g14289(.I(new_n14481_), .ZN(new_n14482_));
  OAI21_X1   g14290(.A1(new_n14477_), .A2(new_n4330_), .B(new_n14482_), .ZN(new_n14483_));
  NAND2_X1   g14291(.A1(new_n14483_), .A2(new_n14476_), .ZN(new_n14484_));
  OAI22_X1   g14292(.A1(new_n14477_), .A2(new_n4330_), .B1(new_n14475_), .B2(new_n14469_), .ZN(new_n14485_));
  NOR4_X1    g14293(.A1(new_n14273_), .A2(\asqrt[40] ), .A3(new_n13924_), .A4(new_n14172_), .ZN(new_n14486_));
  AOI21_X1   g14294(.A1(new_n14478_), .A2(new_n13920_), .B(new_n4018_), .ZN(new_n14487_));
  NOR2_X1    g14295(.A1(new_n14486_), .A2(new_n14487_), .ZN(new_n14488_));
  NAND2_X1   g14296(.A1(new_n14488_), .A2(new_n3760_), .ZN(new_n14489_));
  AOI21_X1   g14297(.A1(new_n14485_), .A2(\asqrt[40] ), .B(new_n14489_), .ZN(new_n14490_));
  NOR2_X1    g14298(.A1(new_n14490_), .A2(new_n14484_), .ZN(new_n14491_));
  AOI22_X1   g14299(.A1(new_n14485_), .A2(\asqrt[40] ), .B1(new_n14483_), .B2(new_n14476_), .ZN(new_n14492_));
  NAND2_X1   g14300(.A1(new_n13936_), .A2(\asqrt[41] ), .ZN(new_n14493_));
  NOR4_X1    g14301(.A1(new_n14273_), .A2(\asqrt[41] ), .A3(new_n13931_), .A4(new_n13936_), .ZN(new_n14494_));
  XOR2_X1    g14302(.A1(new_n14494_), .A2(new_n14493_), .Z(new_n14495_));
  NAND2_X1   g14303(.A1(new_n14495_), .A2(new_n3481_), .ZN(new_n14496_));
  INV_X1     g14304(.I(new_n14496_), .ZN(new_n14497_));
  OAI21_X1   g14305(.A1(new_n14492_), .A2(new_n3760_), .B(new_n14497_), .ZN(new_n14498_));
  NAND2_X1   g14306(.A1(new_n14498_), .A2(new_n14491_), .ZN(new_n14499_));
  OAI22_X1   g14307(.A1(new_n14492_), .A2(new_n3760_), .B1(new_n14490_), .B2(new_n14484_), .ZN(new_n14500_));
  NOR4_X1    g14308(.A1(new_n14273_), .A2(\asqrt[42] ), .A3(new_n13939_), .A4(new_n14179_), .ZN(new_n14501_));
  AOI21_X1   g14309(.A1(new_n14493_), .A2(new_n13935_), .B(new_n3481_), .ZN(new_n14502_));
  NOR2_X1    g14310(.A1(new_n14501_), .A2(new_n14502_), .ZN(new_n14503_));
  NAND2_X1   g14311(.A1(new_n14503_), .A2(new_n3208_), .ZN(new_n14504_));
  AOI21_X1   g14312(.A1(new_n14500_), .A2(\asqrt[42] ), .B(new_n14504_), .ZN(new_n14505_));
  NOR2_X1    g14313(.A1(new_n14505_), .A2(new_n14499_), .ZN(new_n14506_));
  AOI22_X1   g14314(.A1(new_n14500_), .A2(\asqrt[42] ), .B1(new_n14498_), .B2(new_n14491_), .ZN(new_n14507_));
  NAND2_X1   g14315(.A1(new_n13951_), .A2(\asqrt[43] ), .ZN(new_n14508_));
  NOR4_X1    g14316(.A1(new_n14273_), .A2(\asqrt[43] ), .A3(new_n13946_), .A4(new_n13951_), .ZN(new_n14509_));
  XOR2_X1    g14317(.A1(new_n14509_), .A2(new_n14508_), .Z(new_n14510_));
  NAND2_X1   g14318(.A1(new_n14510_), .A2(new_n2941_), .ZN(new_n14511_));
  INV_X1     g14319(.I(new_n14511_), .ZN(new_n14512_));
  OAI21_X1   g14320(.A1(new_n14507_), .A2(new_n3208_), .B(new_n14512_), .ZN(new_n14513_));
  NAND2_X1   g14321(.A1(new_n14513_), .A2(new_n14506_), .ZN(new_n14514_));
  OAI22_X1   g14322(.A1(new_n14507_), .A2(new_n3208_), .B1(new_n14505_), .B2(new_n14499_), .ZN(new_n14515_));
  NAND2_X1   g14323(.A1(new_n14186_), .A2(\asqrt[44] ), .ZN(new_n14516_));
  NOR4_X1    g14324(.A1(new_n14273_), .A2(\asqrt[44] ), .A3(new_n13954_), .A4(new_n14186_), .ZN(new_n14517_));
  XOR2_X1    g14325(.A1(new_n14517_), .A2(new_n14516_), .Z(new_n14518_));
  NAND2_X1   g14326(.A1(new_n14518_), .A2(new_n2728_), .ZN(new_n14519_));
  AOI21_X1   g14327(.A1(new_n14515_), .A2(\asqrt[44] ), .B(new_n14519_), .ZN(new_n14520_));
  NOR2_X1    g14328(.A1(new_n14520_), .A2(new_n14514_), .ZN(new_n14521_));
  AOI22_X1   g14329(.A1(new_n14515_), .A2(\asqrt[44] ), .B1(new_n14513_), .B2(new_n14506_), .ZN(new_n14522_));
  NOR4_X1    g14330(.A1(new_n14273_), .A2(\asqrt[45] ), .A3(new_n13961_), .A4(new_n13966_), .ZN(new_n14523_));
  AOI21_X1   g14331(.A1(new_n14516_), .A2(new_n14185_), .B(new_n2728_), .ZN(new_n14524_));
  NOR2_X1    g14332(.A1(new_n14523_), .A2(new_n14524_), .ZN(new_n14525_));
  NAND2_X1   g14333(.A1(new_n14525_), .A2(new_n2488_), .ZN(new_n14526_));
  INV_X1     g14334(.I(new_n14526_), .ZN(new_n14527_));
  OAI21_X1   g14335(.A1(new_n14522_), .A2(new_n2728_), .B(new_n14527_), .ZN(new_n14528_));
  NAND2_X1   g14336(.A1(new_n14528_), .A2(new_n14521_), .ZN(new_n14529_));
  OAI22_X1   g14337(.A1(new_n14522_), .A2(new_n2728_), .B1(new_n14520_), .B2(new_n14514_), .ZN(new_n14530_));
  NAND2_X1   g14338(.A1(new_n14193_), .A2(\asqrt[46] ), .ZN(new_n14531_));
  NOR4_X1    g14339(.A1(new_n14273_), .A2(\asqrt[46] ), .A3(new_n13969_), .A4(new_n14193_), .ZN(new_n14532_));
  XOR2_X1    g14340(.A1(new_n14532_), .A2(new_n14531_), .Z(new_n14533_));
  NAND2_X1   g14341(.A1(new_n14533_), .A2(new_n2253_), .ZN(new_n14534_));
  AOI21_X1   g14342(.A1(new_n14530_), .A2(\asqrt[46] ), .B(new_n14534_), .ZN(new_n14535_));
  NOR2_X1    g14343(.A1(new_n14535_), .A2(new_n14529_), .ZN(new_n14536_));
  AOI22_X1   g14344(.A1(new_n14530_), .A2(\asqrt[46] ), .B1(new_n14528_), .B2(new_n14521_), .ZN(new_n14537_));
  NOR4_X1    g14345(.A1(new_n14273_), .A2(\asqrt[47] ), .A3(new_n13976_), .A4(new_n13981_), .ZN(new_n14538_));
  AOI21_X1   g14346(.A1(new_n14531_), .A2(new_n14192_), .B(new_n2253_), .ZN(new_n14539_));
  NOR2_X1    g14347(.A1(new_n14538_), .A2(new_n14539_), .ZN(new_n14540_));
  NAND2_X1   g14348(.A1(new_n14540_), .A2(new_n2046_), .ZN(new_n14541_));
  INV_X1     g14349(.I(new_n14541_), .ZN(new_n14542_));
  OAI21_X1   g14350(.A1(new_n14537_), .A2(new_n2253_), .B(new_n14542_), .ZN(new_n14543_));
  NAND2_X1   g14351(.A1(new_n14543_), .A2(new_n14536_), .ZN(new_n14544_));
  OAI22_X1   g14352(.A1(new_n14537_), .A2(new_n2253_), .B1(new_n14535_), .B2(new_n14529_), .ZN(new_n14545_));
  NAND2_X1   g14353(.A1(new_n14200_), .A2(\asqrt[48] ), .ZN(new_n14546_));
  NOR4_X1    g14354(.A1(new_n14273_), .A2(\asqrt[48] ), .A3(new_n13984_), .A4(new_n14200_), .ZN(new_n14547_));
  XOR2_X1    g14355(.A1(new_n14547_), .A2(new_n14546_), .Z(new_n14548_));
  NAND2_X1   g14356(.A1(new_n14548_), .A2(new_n1854_), .ZN(new_n14549_));
  AOI21_X1   g14357(.A1(new_n14545_), .A2(\asqrt[48] ), .B(new_n14549_), .ZN(new_n14550_));
  NOR2_X1    g14358(.A1(new_n14550_), .A2(new_n14544_), .ZN(new_n14551_));
  AOI22_X1   g14359(.A1(new_n14545_), .A2(\asqrt[48] ), .B1(new_n14543_), .B2(new_n14536_), .ZN(new_n14552_));
  NAND2_X1   g14360(.A1(new_n13996_), .A2(\asqrt[49] ), .ZN(new_n14553_));
  NOR4_X1    g14361(.A1(new_n14273_), .A2(\asqrt[49] ), .A3(new_n13991_), .A4(new_n13996_), .ZN(new_n14554_));
  XOR2_X1    g14362(.A1(new_n14554_), .A2(new_n14553_), .Z(new_n14555_));
  NAND2_X1   g14363(.A1(new_n14555_), .A2(new_n1595_), .ZN(new_n14556_));
  INV_X1     g14364(.I(new_n14556_), .ZN(new_n14557_));
  OAI21_X1   g14365(.A1(new_n14552_), .A2(new_n1854_), .B(new_n14557_), .ZN(new_n14558_));
  NAND2_X1   g14366(.A1(new_n14558_), .A2(new_n14551_), .ZN(new_n14559_));
  OAI22_X1   g14367(.A1(new_n14552_), .A2(new_n1854_), .B1(new_n14550_), .B2(new_n14544_), .ZN(new_n14560_));
  NOR4_X1    g14368(.A1(new_n14273_), .A2(\asqrt[50] ), .A3(new_n13999_), .A4(new_n14207_), .ZN(new_n14561_));
  AOI21_X1   g14369(.A1(new_n14553_), .A2(new_n13995_), .B(new_n1595_), .ZN(new_n14562_));
  NOR2_X1    g14370(.A1(new_n14561_), .A2(new_n14562_), .ZN(new_n14563_));
  NAND2_X1   g14371(.A1(new_n14563_), .A2(new_n1436_), .ZN(new_n14564_));
  AOI21_X1   g14372(.A1(new_n14560_), .A2(\asqrt[50] ), .B(new_n14564_), .ZN(new_n14565_));
  NOR2_X1    g14373(.A1(new_n14565_), .A2(new_n14559_), .ZN(new_n14566_));
  AOI22_X1   g14374(.A1(new_n14560_), .A2(\asqrt[50] ), .B1(new_n14558_), .B2(new_n14551_), .ZN(new_n14567_));
  NAND2_X1   g14375(.A1(new_n14011_), .A2(\asqrt[51] ), .ZN(new_n14568_));
  NOR4_X1    g14376(.A1(new_n14273_), .A2(\asqrt[51] ), .A3(new_n14006_), .A4(new_n14011_), .ZN(new_n14569_));
  XOR2_X1    g14377(.A1(new_n14569_), .A2(new_n14568_), .Z(new_n14570_));
  NAND2_X1   g14378(.A1(new_n14570_), .A2(new_n1260_), .ZN(new_n14571_));
  INV_X1     g14379(.I(new_n14571_), .ZN(new_n14572_));
  OAI21_X1   g14380(.A1(new_n14567_), .A2(new_n1436_), .B(new_n14572_), .ZN(new_n14573_));
  NAND2_X1   g14381(.A1(new_n14573_), .A2(new_n14566_), .ZN(new_n14574_));
  OAI22_X1   g14382(.A1(new_n14567_), .A2(new_n1436_), .B1(new_n14565_), .B2(new_n14559_), .ZN(new_n14575_));
  NOR4_X1    g14383(.A1(new_n14273_), .A2(\asqrt[52] ), .A3(new_n14014_), .A4(new_n14214_), .ZN(new_n14576_));
  AOI21_X1   g14384(.A1(new_n14568_), .A2(new_n14010_), .B(new_n1260_), .ZN(new_n14577_));
  NOR2_X1    g14385(.A1(new_n14576_), .A2(new_n14577_), .ZN(new_n14578_));
  NAND2_X1   g14386(.A1(new_n14578_), .A2(new_n1096_), .ZN(new_n14579_));
  AOI21_X1   g14387(.A1(new_n14575_), .A2(\asqrt[52] ), .B(new_n14579_), .ZN(new_n14580_));
  NOR2_X1    g14388(.A1(new_n14580_), .A2(new_n14574_), .ZN(new_n14581_));
  AOI22_X1   g14389(.A1(new_n14575_), .A2(\asqrt[52] ), .B1(new_n14573_), .B2(new_n14566_), .ZN(new_n14582_));
  NAND2_X1   g14390(.A1(new_n14025_), .A2(\asqrt[53] ), .ZN(new_n14583_));
  NOR4_X1    g14391(.A1(new_n14273_), .A2(\asqrt[53] ), .A3(new_n14020_), .A4(new_n14025_), .ZN(new_n14584_));
  XOR2_X1    g14392(.A1(new_n14584_), .A2(new_n14583_), .Z(new_n14585_));
  NAND2_X1   g14393(.A1(new_n14585_), .A2(new_n970_), .ZN(new_n14586_));
  INV_X1     g14394(.I(new_n14586_), .ZN(new_n14587_));
  OAI21_X1   g14395(.A1(new_n14582_), .A2(new_n1096_), .B(new_n14587_), .ZN(new_n14588_));
  NAND2_X1   g14396(.A1(new_n14588_), .A2(new_n14581_), .ZN(new_n14589_));
  OAI22_X1   g14397(.A1(new_n14582_), .A2(new_n1096_), .B1(new_n14580_), .B2(new_n14574_), .ZN(new_n14590_));
  NOR2_X1    g14398(.A1(new_n14031_), .A2(new_n970_), .ZN(new_n14591_));
  NOR4_X1    g14399(.A1(new_n14273_), .A2(\asqrt[54] ), .A3(new_n14027_), .A4(new_n14221_), .ZN(new_n14592_));
  XNOR2_X1   g14400(.A1(new_n14592_), .A2(new_n14591_), .ZN(new_n14593_));
  NAND2_X1   g14401(.A1(new_n14593_), .A2(new_n825_), .ZN(new_n14594_));
  AOI21_X1   g14402(.A1(new_n14590_), .A2(\asqrt[54] ), .B(new_n14594_), .ZN(new_n14595_));
  NOR2_X1    g14403(.A1(new_n14595_), .A2(new_n14589_), .ZN(new_n14596_));
  AOI22_X1   g14404(.A1(new_n14590_), .A2(\asqrt[54] ), .B1(new_n14588_), .B2(new_n14581_), .ZN(new_n14597_));
  NOR4_X1    g14405(.A1(new_n14273_), .A2(\asqrt[55] ), .A3(new_n14033_), .A4(new_n14038_), .ZN(new_n14598_));
  XOR2_X1    g14406(.A1(new_n14598_), .A2(new_n14274_), .Z(new_n14599_));
  NAND2_X1   g14407(.A1(new_n14599_), .A2(new_n724_), .ZN(new_n14600_));
  INV_X1     g14408(.I(new_n14600_), .ZN(new_n14601_));
  OAI21_X1   g14409(.A1(new_n14597_), .A2(new_n825_), .B(new_n14601_), .ZN(new_n14602_));
  NAND2_X1   g14410(.A1(new_n14602_), .A2(new_n14596_), .ZN(new_n14603_));
  OAI22_X1   g14411(.A1(new_n14597_), .A2(new_n825_), .B1(new_n14595_), .B2(new_n14589_), .ZN(new_n14604_));
  NOR4_X1    g14412(.A1(new_n14273_), .A2(\asqrt[56] ), .A3(new_n14040_), .A4(new_n14228_), .ZN(new_n14605_));
  XOR2_X1    g14413(.A1(new_n14605_), .A2(new_n14289_), .Z(new_n14606_));
  NAND2_X1   g14414(.A1(new_n14606_), .A2(new_n587_), .ZN(new_n14607_));
  AOI21_X1   g14415(.A1(new_n14604_), .A2(\asqrt[56] ), .B(new_n14607_), .ZN(new_n14608_));
  NOR2_X1    g14416(.A1(new_n14608_), .A2(new_n14603_), .ZN(new_n14609_));
  AOI22_X1   g14417(.A1(new_n14604_), .A2(\asqrt[56] ), .B1(new_n14602_), .B2(new_n14596_), .ZN(new_n14610_));
  NOR4_X1    g14418(.A1(new_n14273_), .A2(\asqrt[57] ), .A3(new_n14046_), .A4(new_n14051_), .ZN(new_n14611_));
  XOR2_X1    g14419(.A1(new_n14611_), .A2(new_n14276_), .Z(new_n14612_));
  AND2_X2    g14420(.A1(new_n14612_), .A2(new_n504_), .Z(new_n14613_));
  OAI21_X1   g14421(.A1(new_n14610_), .A2(new_n587_), .B(new_n14613_), .ZN(new_n14614_));
  NAND2_X1   g14422(.A1(new_n14614_), .A2(new_n14609_), .ZN(new_n14615_));
  OAI22_X1   g14423(.A1(new_n14610_), .A2(new_n587_), .B1(new_n14608_), .B2(new_n14603_), .ZN(new_n14616_));
  NOR4_X1    g14424(.A1(new_n14273_), .A2(\asqrt[58] ), .A3(new_n14053_), .A4(new_n14235_), .ZN(new_n14617_));
  XOR2_X1    g14425(.A1(new_n14617_), .A2(new_n14291_), .Z(new_n14618_));
  NAND2_X1   g14426(.A1(new_n14618_), .A2(new_n376_), .ZN(new_n14619_));
  AOI21_X1   g14427(.A1(new_n14616_), .A2(\asqrt[58] ), .B(new_n14619_), .ZN(new_n14620_));
  NOR2_X1    g14428(.A1(new_n14620_), .A2(new_n14615_), .ZN(new_n14621_));
  AOI22_X1   g14429(.A1(new_n14616_), .A2(\asqrt[58] ), .B1(new_n14614_), .B2(new_n14609_), .ZN(new_n14622_));
  NOR4_X1    g14430(.A1(new_n14273_), .A2(\asqrt[59] ), .A3(new_n14059_), .A4(new_n14064_), .ZN(new_n14623_));
  XOR2_X1    g14431(.A1(new_n14623_), .A2(new_n14278_), .Z(new_n14624_));
  AND2_X2    g14432(.A1(new_n14624_), .A2(new_n275_), .Z(new_n14625_));
  OAI21_X1   g14433(.A1(new_n14622_), .A2(new_n376_), .B(new_n14625_), .ZN(new_n14626_));
  NAND2_X1   g14434(.A1(new_n14626_), .A2(new_n14621_), .ZN(new_n14627_));
  NAND2_X1   g14435(.A1(new_n14575_), .A2(\asqrt[52] ), .ZN(new_n14628_));
  AOI21_X1   g14436(.A1(new_n14628_), .A2(new_n14574_), .B(new_n1096_), .ZN(new_n14629_));
  OAI21_X1   g14437(.A1(new_n14581_), .A2(new_n14629_), .B(\asqrt[54] ), .ZN(new_n14630_));
  AOI21_X1   g14438(.A1(new_n14589_), .A2(new_n14630_), .B(new_n825_), .ZN(new_n14631_));
  OAI21_X1   g14439(.A1(new_n14596_), .A2(new_n14631_), .B(\asqrt[56] ), .ZN(new_n14632_));
  AOI21_X1   g14440(.A1(new_n14603_), .A2(new_n14632_), .B(new_n587_), .ZN(new_n14633_));
  OAI21_X1   g14441(.A1(new_n14609_), .A2(new_n14633_), .B(\asqrt[58] ), .ZN(new_n14634_));
  AOI21_X1   g14442(.A1(new_n14615_), .A2(new_n14634_), .B(new_n376_), .ZN(new_n14635_));
  OAI21_X1   g14443(.A1(new_n14621_), .A2(new_n14635_), .B(\asqrt[60] ), .ZN(new_n14636_));
  AOI21_X1   g14444(.A1(new_n14627_), .A2(new_n14636_), .B(new_n229_), .ZN(new_n14637_));
  NOR2_X1    g14445(.A1(new_n14260_), .A2(new_n196_), .ZN(new_n14638_));
  NOR2_X1    g14446(.A1(new_n14245_), .A2(\asqrt[62] ), .ZN(new_n14639_));
  NAND3_X1   g14447(.A1(new_n14639_), .A2(new_n14638_), .A3(new_n14078_), .ZN(new_n14640_));
  NOR2_X1    g14448(.A1(new_n14273_), .A2(new_n14640_), .ZN(new_n14641_));
  OR3_X2     g14449(.A1(\asqrt[16] ), .A2(new_n14078_), .A3(new_n14639_), .Z(new_n14642_));
  AOI21_X1   g14450(.A1(new_n14642_), .A2(new_n14638_), .B(new_n14641_), .ZN(new_n14643_));
  NOR4_X1    g14451(.A1(new_n14273_), .A2(\asqrt[61] ), .A3(new_n14072_), .A4(new_n14077_), .ZN(new_n14644_));
  XOR2_X1    g14452(.A1(new_n14644_), .A2(new_n14280_), .Z(new_n14645_));
  NOR2_X1    g14453(.A1(new_n14645_), .A2(new_n196_), .ZN(new_n14646_));
  INV_X1     g14454(.I(new_n14646_), .ZN(new_n14647_));
  NAND2_X1   g14455(.A1(new_n14326_), .A2(new_n14332_), .ZN(new_n14648_));
  NAND3_X1   g14456(.A1(new_n14648_), .A2(new_n14313_), .A3(new_n14349_), .ZN(new_n14649_));
  INV_X1     g14457(.I(new_n14252_), .ZN(new_n14650_));
  AOI21_X1   g14458(.A1(new_n14264_), .A2(new_n14650_), .B(new_n14254_), .ZN(new_n14651_));
  NOR3_X1    g14459(.A1(new_n14251_), .A2(new_n13694_), .A3(new_n13706_), .ZN(new_n14652_));
  NOR2_X1    g14460(.A1(new_n14652_), .A2(new_n14651_), .ZN(new_n14653_));
  NOR3_X1    g14461(.A1(new_n14299_), .A2(new_n13736_), .A3(\asqrt[16] ), .ZN(new_n14654_));
  AOI21_X1   g14462(.A1(new_n14286_), .A2(new_n13735_), .B(new_n14273_), .ZN(new_n14655_));
  NOR4_X1    g14463(.A1(new_n14654_), .A2(new_n14655_), .A3(\asqrt[18] ), .A4(new_n14271_), .ZN(new_n14656_));
  NOR2_X1    g14464(.A1(new_n14656_), .A2(new_n14653_), .ZN(new_n14657_));
  NOR3_X1    g14465(.A1(new_n14652_), .A2(new_n14651_), .A3(new_n14271_), .ZN(new_n14658_));
  NOR3_X1    g14466(.A1(new_n14273_), .A2(new_n13758_), .A3(new_n14307_), .ZN(new_n14659_));
  AOI21_X1   g14467(.A1(\asqrt[16] ), .A2(new_n14308_), .B(new_n13759_), .ZN(new_n14660_));
  NOR3_X1    g14468(.A1(new_n14660_), .A2(new_n14659_), .A3(\asqrt[19] ), .ZN(new_n14661_));
  OAI21_X1   g14469(.A1(new_n14658_), .A2(new_n13192_), .B(new_n14661_), .ZN(new_n14662_));
  NAND2_X1   g14470(.A1(new_n14657_), .A2(new_n14662_), .ZN(new_n14663_));
  OAI22_X1   g14471(.A1(new_n14656_), .A2(new_n14653_), .B1(new_n13192_), .B2(new_n14658_), .ZN(new_n14664_));
  AOI21_X1   g14472(.A1(new_n14664_), .A2(\asqrt[19] ), .B(new_n14324_), .ZN(new_n14665_));
  AOI22_X1   g14473(.A1(new_n14664_), .A2(\asqrt[19] ), .B1(new_n14657_), .B2(new_n14662_), .ZN(new_n14666_));
  OAI22_X1   g14474(.A1(new_n14666_), .A2(new_n12101_), .B1(new_n14665_), .B2(new_n14663_), .ZN(new_n14667_));
  AOI21_X1   g14475(.A1(new_n14667_), .A2(\asqrt[21] ), .B(new_n14339_), .ZN(new_n14668_));
  NOR2_X1    g14476(.A1(new_n14668_), .A2(new_n14649_), .ZN(new_n14669_));
  NAND2_X1   g14477(.A1(new_n14341_), .A2(new_n14346_), .ZN(new_n14670_));
  NAND2_X1   g14478(.A1(new_n14670_), .A2(new_n14669_), .ZN(new_n14671_));
  NOR2_X1    g14479(.A1(new_n14333_), .A2(new_n14334_), .ZN(new_n14672_));
  OAI22_X1   g14480(.A1(new_n14672_), .A2(new_n11105_), .B1(new_n14668_), .B2(new_n14649_), .ZN(new_n14673_));
  AOI21_X1   g14481(.A1(new_n14673_), .A2(\asqrt[23] ), .B(new_n14360_), .ZN(new_n14674_));
  NOR2_X1    g14482(.A1(new_n14674_), .A2(new_n14671_), .ZN(new_n14675_));
  AOI21_X1   g14483(.A1(new_n14340_), .A2(new_n14341_), .B(new_n10614_), .ZN(new_n14676_));
  OAI21_X1   g14484(.A1(new_n14347_), .A2(new_n14676_), .B(\asqrt[24] ), .ZN(new_n14677_));
  INV_X1     g14485(.I(new_n14369_), .ZN(new_n14678_));
  NAND2_X1   g14486(.A1(new_n14677_), .A2(new_n14678_), .ZN(new_n14679_));
  NAND2_X1   g14487(.A1(new_n14679_), .A2(new_n14675_), .ZN(new_n14680_));
  AOI22_X1   g14488(.A1(new_n14673_), .A2(\asqrt[23] ), .B1(new_n14670_), .B2(new_n14669_), .ZN(new_n14681_));
  OAI22_X1   g14489(.A1(new_n14681_), .A2(new_n10104_), .B1(new_n14674_), .B2(new_n14671_), .ZN(new_n14682_));
  AOI21_X1   g14490(.A1(new_n14682_), .A2(\asqrt[25] ), .B(new_n14376_), .ZN(new_n14683_));
  NOR2_X1    g14491(.A1(new_n14683_), .A2(new_n14680_), .ZN(new_n14684_));
  AOI22_X1   g14492(.A1(new_n14682_), .A2(\asqrt[25] ), .B1(new_n14679_), .B2(new_n14675_), .ZN(new_n14685_));
  INV_X1     g14493(.I(new_n14384_), .ZN(new_n14686_));
  OAI21_X1   g14494(.A1(new_n14685_), .A2(new_n9212_), .B(new_n14686_), .ZN(new_n14687_));
  NAND2_X1   g14495(.A1(new_n14687_), .A2(new_n14684_), .ZN(new_n14688_));
  OAI22_X1   g14496(.A1(new_n14685_), .A2(new_n9212_), .B1(new_n14683_), .B2(new_n14680_), .ZN(new_n14689_));
  AOI21_X1   g14497(.A1(new_n14689_), .A2(\asqrt[27] ), .B(new_n14391_), .ZN(new_n14690_));
  NOR2_X1    g14498(.A1(new_n14690_), .A2(new_n14688_), .ZN(new_n14691_));
  AOI22_X1   g14499(.A1(new_n14689_), .A2(\asqrt[27] ), .B1(new_n14687_), .B2(new_n14684_), .ZN(new_n14692_));
  INV_X1     g14500(.I(new_n14399_), .ZN(new_n14693_));
  OAI21_X1   g14501(.A1(new_n14692_), .A2(new_n8319_), .B(new_n14693_), .ZN(new_n14694_));
  NAND2_X1   g14502(.A1(new_n14694_), .A2(new_n14691_), .ZN(new_n14695_));
  OAI22_X1   g14503(.A1(new_n14692_), .A2(new_n8319_), .B1(new_n14690_), .B2(new_n14688_), .ZN(new_n14696_));
  AOI21_X1   g14504(.A1(new_n14696_), .A2(\asqrt[29] ), .B(new_n14406_), .ZN(new_n14697_));
  NOR2_X1    g14505(.A1(new_n14697_), .A2(new_n14695_), .ZN(new_n14698_));
  AOI22_X1   g14506(.A1(new_n14696_), .A2(\asqrt[29] ), .B1(new_n14694_), .B2(new_n14691_), .ZN(new_n14699_));
  INV_X1     g14507(.I(new_n14414_), .ZN(new_n14700_));
  OAI21_X1   g14508(.A1(new_n14699_), .A2(new_n7517_), .B(new_n14700_), .ZN(new_n14701_));
  NAND2_X1   g14509(.A1(new_n14701_), .A2(new_n14698_), .ZN(new_n14702_));
  OAI22_X1   g14510(.A1(new_n14699_), .A2(new_n7517_), .B1(new_n14697_), .B2(new_n14695_), .ZN(new_n14703_));
  AOI21_X1   g14511(.A1(new_n14703_), .A2(\asqrt[31] ), .B(new_n14421_), .ZN(new_n14704_));
  NOR2_X1    g14512(.A1(new_n14704_), .A2(new_n14702_), .ZN(new_n14705_));
  AOI22_X1   g14513(.A1(new_n14703_), .A2(\asqrt[31] ), .B1(new_n14701_), .B2(new_n14698_), .ZN(new_n14706_));
  INV_X1     g14514(.I(new_n14429_), .ZN(new_n14707_));
  OAI21_X1   g14515(.A1(new_n14706_), .A2(new_n6708_), .B(new_n14707_), .ZN(new_n14708_));
  NAND2_X1   g14516(.A1(new_n14708_), .A2(new_n14705_), .ZN(new_n14709_));
  OAI22_X1   g14517(.A1(new_n14706_), .A2(new_n6708_), .B1(new_n14704_), .B2(new_n14702_), .ZN(new_n14710_));
  AOI21_X1   g14518(.A1(new_n14710_), .A2(\asqrt[33] ), .B(new_n14436_), .ZN(new_n14711_));
  NOR2_X1    g14519(.A1(new_n14711_), .A2(new_n14709_), .ZN(new_n14712_));
  AOI22_X1   g14520(.A1(new_n14710_), .A2(\asqrt[33] ), .B1(new_n14708_), .B2(new_n14705_), .ZN(new_n14713_));
  INV_X1     g14521(.I(new_n14444_), .ZN(new_n14714_));
  OAI21_X1   g14522(.A1(new_n14713_), .A2(new_n5991_), .B(new_n14714_), .ZN(new_n14715_));
  NAND2_X1   g14523(.A1(new_n14715_), .A2(new_n14712_), .ZN(new_n14716_));
  OAI22_X1   g14524(.A1(new_n14713_), .A2(new_n5991_), .B1(new_n14711_), .B2(new_n14709_), .ZN(new_n14717_));
  AOI21_X1   g14525(.A1(new_n14717_), .A2(\asqrt[35] ), .B(new_n14451_), .ZN(new_n14718_));
  NOR2_X1    g14526(.A1(new_n14718_), .A2(new_n14716_), .ZN(new_n14719_));
  AOI22_X1   g14527(.A1(new_n14717_), .A2(\asqrt[35] ), .B1(new_n14715_), .B2(new_n14712_), .ZN(new_n14720_));
  INV_X1     g14528(.I(new_n14459_), .ZN(new_n14721_));
  OAI21_X1   g14529(.A1(new_n14720_), .A2(new_n5273_), .B(new_n14721_), .ZN(new_n14722_));
  NAND2_X1   g14530(.A1(new_n14722_), .A2(new_n14719_), .ZN(new_n14723_));
  OAI22_X1   g14531(.A1(new_n14720_), .A2(new_n5273_), .B1(new_n14718_), .B2(new_n14716_), .ZN(new_n14724_));
  AOI21_X1   g14532(.A1(new_n14724_), .A2(\asqrt[37] ), .B(new_n14466_), .ZN(new_n14725_));
  NOR2_X1    g14533(.A1(new_n14725_), .A2(new_n14723_), .ZN(new_n14726_));
  AOI22_X1   g14534(.A1(new_n14724_), .A2(\asqrt[37] ), .B1(new_n14722_), .B2(new_n14719_), .ZN(new_n14727_));
  INV_X1     g14535(.I(new_n14474_), .ZN(new_n14728_));
  OAI21_X1   g14536(.A1(new_n14727_), .A2(new_n4645_), .B(new_n14728_), .ZN(new_n14729_));
  NAND2_X1   g14537(.A1(new_n14729_), .A2(new_n14726_), .ZN(new_n14730_));
  OAI22_X1   g14538(.A1(new_n14727_), .A2(new_n4645_), .B1(new_n14725_), .B2(new_n14723_), .ZN(new_n14731_));
  AOI21_X1   g14539(.A1(new_n14731_), .A2(\asqrt[39] ), .B(new_n14481_), .ZN(new_n14732_));
  NOR2_X1    g14540(.A1(new_n14732_), .A2(new_n14730_), .ZN(new_n14733_));
  AOI22_X1   g14541(.A1(new_n14731_), .A2(\asqrt[39] ), .B1(new_n14729_), .B2(new_n14726_), .ZN(new_n14734_));
  INV_X1     g14542(.I(new_n14489_), .ZN(new_n14735_));
  OAI21_X1   g14543(.A1(new_n14734_), .A2(new_n4018_), .B(new_n14735_), .ZN(new_n14736_));
  NAND2_X1   g14544(.A1(new_n14736_), .A2(new_n14733_), .ZN(new_n14737_));
  OAI22_X1   g14545(.A1(new_n14734_), .A2(new_n4018_), .B1(new_n14732_), .B2(new_n14730_), .ZN(new_n14738_));
  AOI21_X1   g14546(.A1(new_n14738_), .A2(\asqrt[41] ), .B(new_n14496_), .ZN(new_n14739_));
  NOR2_X1    g14547(.A1(new_n14739_), .A2(new_n14737_), .ZN(new_n14740_));
  AOI22_X1   g14548(.A1(new_n14738_), .A2(\asqrt[41] ), .B1(new_n14736_), .B2(new_n14733_), .ZN(new_n14741_));
  INV_X1     g14549(.I(new_n14504_), .ZN(new_n14742_));
  OAI21_X1   g14550(.A1(new_n14741_), .A2(new_n3481_), .B(new_n14742_), .ZN(new_n14743_));
  NAND2_X1   g14551(.A1(new_n14743_), .A2(new_n14740_), .ZN(new_n14744_));
  OAI22_X1   g14552(.A1(new_n14741_), .A2(new_n3481_), .B1(new_n14739_), .B2(new_n14737_), .ZN(new_n14745_));
  AOI21_X1   g14553(.A1(new_n14745_), .A2(\asqrt[43] ), .B(new_n14511_), .ZN(new_n14746_));
  NOR2_X1    g14554(.A1(new_n14746_), .A2(new_n14744_), .ZN(new_n14747_));
  AOI22_X1   g14555(.A1(new_n14745_), .A2(\asqrt[43] ), .B1(new_n14743_), .B2(new_n14740_), .ZN(new_n14748_));
  INV_X1     g14556(.I(new_n14519_), .ZN(new_n14749_));
  OAI21_X1   g14557(.A1(new_n14748_), .A2(new_n2941_), .B(new_n14749_), .ZN(new_n14750_));
  NAND2_X1   g14558(.A1(new_n14750_), .A2(new_n14747_), .ZN(new_n14751_));
  OAI22_X1   g14559(.A1(new_n14748_), .A2(new_n2941_), .B1(new_n14746_), .B2(new_n14744_), .ZN(new_n14752_));
  AOI21_X1   g14560(.A1(new_n14752_), .A2(\asqrt[45] ), .B(new_n14526_), .ZN(new_n14753_));
  NOR2_X1    g14561(.A1(new_n14753_), .A2(new_n14751_), .ZN(new_n14754_));
  AOI22_X1   g14562(.A1(new_n14752_), .A2(\asqrt[45] ), .B1(new_n14750_), .B2(new_n14747_), .ZN(new_n14755_));
  INV_X1     g14563(.I(new_n14534_), .ZN(new_n14756_));
  OAI21_X1   g14564(.A1(new_n14755_), .A2(new_n2488_), .B(new_n14756_), .ZN(new_n14757_));
  NAND2_X1   g14565(.A1(new_n14757_), .A2(new_n14754_), .ZN(new_n14758_));
  OAI22_X1   g14566(.A1(new_n14755_), .A2(new_n2488_), .B1(new_n14753_), .B2(new_n14751_), .ZN(new_n14759_));
  AOI21_X1   g14567(.A1(new_n14759_), .A2(\asqrt[47] ), .B(new_n14541_), .ZN(new_n14760_));
  NOR2_X1    g14568(.A1(new_n14760_), .A2(new_n14758_), .ZN(new_n14761_));
  AOI22_X1   g14569(.A1(new_n14759_), .A2(\asqrt[47] ), .B1(new_n14757_), .B2(new_n14754_), .ZN(new_n14762_));
  INV_X1     g14570(.I(new_n14549_), .ZN(new_n14763_));
  OAI21_X1   g14571(.A1(new_n14762_), .A2(new_n2046_), .B(new_n14763_), .ZN(new_n14764_));
  NAND2_X1   g14572(.A1(new_n14764_), .A2(new_n14761_), .ZN(new_n14765_));
  OAI22_X1   g14573(.A1(new_n14762_), .A2(new_n2046_), .B1(new_n14760_), .B2(new_n14758_), .ZN(new_n14766_));
  AOI21_X1   g14574(.A1(new_n14766_), .A2(\asqrt[49] ), .B(new_n14556_), .ZN(new_n14767_));
  NOR2_X1    g14575(.A1(new_n14767_), .A2(new_n14765_), .ZN(new_n14768_));
  AOI22_X1   g14576(.A1(new_n14766_), .A2(\asqrt[49] ), .B1(new_n14764_), .B2(new_n14761_), .ZN(new_n14769_));
  INV_X1     g14577(.I(new_n14564_), .ZN(new_n14770_));
  OAI21_X1   g14578(.A1(new_n14769_), .A2(new_n1595_), .B(new_n14770_), .ZN(new_n14771_));
  NAND2_X1   g14579(.A1(new_n14771_), .A2(new_n14768_), .ZN(new_n14772_));
  OAI22_X1   g14580(.A1(new_n14769_), .A2(new_n1595_), .B1(new_n14767_), .B2(new_n14765_), .ZN(new_n14773_));
  AOI21_X1   g14581(.A1(new_n14773_), .A2(\asqrt[51] ), .B(new_n14571_), .ZN(new_n14774_));
  NOR2_X1    g14582(.A1(new_n14774_), .A2(new_n14772_), .ZN(new_n14775_));
  AOI22_X1   g14583(.A1(new_n14773_), .A2(\asqrt[51] ), .B1(new_n14771_), .B2(new_n14768_), .ZN(new_n14776_));
  INV_X1     g14584(.I(new_n14579_), .ZN(new_n14777_));
  OAI21_X1   g14585(.A1(new_n14776_), .A2(new_n1260_), .B(new_n14777_), .ZN(new_n14778_));
  NAND2_X1   g14586(.A1(new_n14778_), .A2(new_n14775_), .ZN(new_n14779_));
  OAI22_X1   g14587(.A1(new_n14776_), .A2(new_n1260_), .B1(new_n14774_), .B2(new_n14772_), .ZN(new_n14780_));
  AOI21_X1   g14588(.A1(new_n14780_), .A2(\asqrt[53] ), .B(new_n14586_), .ZN(new_n14781_));
  NOR2_X1    g14589(.A1(new_n14781_), .A2(new_n14779_), .ZN(new_n14782_));
  AOI22_X1   g14590(.A1(new_n14780_), .A2(\asqrt[53] ), .B1(new_n14778_), .B2(new_n14775_), .ZN(new_n14783_));
  INV_X1     g14591(.I(new_n14594_), .ZN(new_n14784_));
  OAI21_X1   g14592(.A1(new_n14783_), .A2(new_n970_), .B(new_n14784_), .ZN(new_n14785_));
  NAND2_X1   g14593(.A1(new_n14785_), .A2(new_n14782_), .ZN(new_n14786_));
  OAI22_X1   g14594(.A1(new_n14783_), .A2(new_n970_), .B1(new_n14781_), .B2(new_n14779_), .ZN(new_n14787_));
  AOI21_X1   g14595(.A1(new_n14787_), .A2(\asqrt[55] ), .B(new_n14600_), .ZN(new_n14788_));
  NOR2_X1    g14596(.A1(new_n14788_), .A2(new_n14786_), .ZN(new_n14789_));
  AOI22_X1   g14597(.A1(new_n14787_), .A2(\asqrt[55] ), .B1(new_n14785_), .B2(new_n14782_), .ZN(new_n14790_));
  INV_X1     g14598(.I(new_n14607_), .ZN(new_n14791_));
  OAI21_X1   g14599(.A1(new_n14790_), .A2(new_n724_), .B(new_n14791_), .ZN(new_n14792_));
  NAND2_X1   g14600(.A1(new_n14792_), .A2(new_n14789_), .ZN(new_n14793_));
  NAND2_X1   g14601(.A1(new_n14787_), .A2(\asqrt[55] ), .ZN(new_n14794_));
  AOI21_X1   g14602(.A1(new_n14794_), .A2(new_n14786_), .B(new_n724_), .ZN(new_n14795_));
  OAI21_X1   g14603(.A1(new_n14789_), .A2(new_n14795_), .B(\asqrt[57] ), .ZN(new_n14796_));
  AOI21_X1   g14604(.A1(new_n14796_), .A2(new_n14613_), .B(new_n14793_), .ZN(new_n14797_));
  OAI22_X1   g14605(.A1(new_n14790_), .A2(new_n724_), .B1(new_n14788_), .B2(new_n14786_), .ZN(new_n14798_));
  AOI22_X1   g14606(.A1(new_n14798_), .A2(\asqrt[57] ), .B1(new_n14792_), .B2(new_n14789_), .ZN(new_n14799_));
  INV_X1     g14607(.I(new_n14619_), .ZN(new_n14800_));
  OAI21_X1   g14608(.A1(new_n14799_), .A2(new_n504_), .B(new_n14800_), .ZN(new_n14801_));
  NAND2_X1   g14609(.A1(new_n14801_), .A2(new_n14797_), .ZN(new_n14802_));
  AOI21_X1   g14610(.A1(new_n14793_), .A2(new_n14796_), .B(new_n504_), .ZN(new_n14803_));
  OAI21_X1   g14611(.A1(new_n14797_), .A2(new_n14803_), .B(\asqrt[59] ), .ZN(new_n14804_));
  AOI21_X1   g14612(.A1(new_n14804_), .A2(new_n14625_), .B(new_n14802_), .ZN(new_n14805_));
  NAND2_X1   g14613(.A1(new_n14615_), .A2(new_n14634_), .ZN(new_n14806_));
  AOI22_X1   g14614(.A1(new_n14806_), .A2(\asqrt[59] ), .B1(new_n14801_), .B2(new_n14797_), .ZN(new_n14807_));
  NOR4_X1    g14615(.A1(new_n14273_), .A2(\asqrt[60] ), .A3(new_n14066_), .A4(new_n14242_), .ZN(new_n14808_));
  XOR2_X1    g14616(.A1(new_n14808_), .A2(new_n14293_), .Z(new_n14809_));
  NAND2_X1   g14617(.A1(new_n14809_), .A2(new_n229_), .ZN(new_n14810_));
  INV_X1     g14618(.I(new_n14810_), .ZN(new_n14811_));
  OAI21_X1   g14619(.A1(new_n14807_), .A2(new_n275_), .B(new_n14811_), .ZN(new_n14812_));
  NAND2_X1   g14620(.A1(new_n14812_), .A2(new_n14805_), .ZN(new_n14813_));
  INV_X1     g14621(.I(new_n14645_), .ZN(new_n14814_));
  NOR2_X1    g14622(.A1(new_n14814_), .A2(\asqrt[62] ), .ZN(new_n14815_));
  INV_X1     g14623(.I(new_n14815_), .ZN(new_n14816_));
  NAND2_X1   g14624(.A1(new_n14637_), .A2(new_n14816_), .ZN(new_n14817_));
  OAI21_X1   g14625(.A1(new_n14817_), .A2(new_n14813_), .B(new_n14647_), .ZN(new_n14818_));
  NOR3_X1    g14626(.A1(\asqrt[16] ), .A2(new_n13728_), .A3(new_n14246_), .ZN(new_n14819_));
  OAI21_X1   g14627(.A1(new_n14819_), .A2(new_n14258_), .B(new_n231_), .ZN(new_n14820_));
  OAI21_X1   g14628(.A1(new_n14818_), .A2(new_n14820_), .B(new_n14643_), .ZN(new_n14821_));
  OAI21_X1   g14629(.A1(new_n13728_), .A2(new_n14082_), .B(\asqrt[16] ), .ZN(new_n14822_));
  XOR2_X1    g14630(.A1(new_n14082_), .A2(\asqrt[63] ), .Z(new_n14823_));
  NAND2_X1   g14631(.A1(new_n14822_), .A2(new_n14823_), .ZN(new_n14824_));
  INV_X1     g14632(.I(new_n14824_), .ZN(new_n14825_));
  INV_X1     g14633(.I(new_n14643_), .ZN(new_n14826_));
  OAI22_X1   g14634(.A1(new_n14622_), .A2(new_n376_), .B1(new_n14620_), .B2(new_n14615_), .ZN(new_n14827_));
  AOI21_X1   g14635(.A1(new_n14827_), .A2(\asqrt[60] ), .B(new_n14810_), .ZN(new_n14828_));
  AOI22_X1   g14636(.A1(new_n14827_), .A2(\asqrt[60] ), .B1(new_n14626_), .B2(new_n14621_), .ZN(new_n14829_));
  OAI22_X1   g14637(.A1(new_n14829_), .A2(new_n229_), .B1(new_n14828_), .B2(new_n14627_), .ZN(new_n14830_));
  NOR4_X1    g14638(.A1(new_n14830_), .A2(\asqrt[62] ), .A3(new_n14826_), .A4(new_n14645_), .ZN(new_n14831_));
  NAND2_X1   g14639(.A1(new_n14831_), .A2(new_n14825_), .ZN(new_n14832_));
  NAND3_X1   g14640(.A1(new_n14267_), .A2(new_n13715_), .A3(new_n13728_), .ZN(new_n14833_));
  NOR3_X1    g14641(.A1(new_n14832_), .A2(new_n14821_), .A3(new_n14833_), .ZN(\asqrt[15] ));
  NAND2_X1   g14642(.A1(new_n14627_), .A2(new_n14636_), .ZN(new_n14835_));
  NOR3_X1    g14643(.A1(new_n14835_), .A2(\asqrt[61] ), .A3(new_n14809_), .ZN(new_n14836_));
  NAND2_X1   g14644(.A1(\asqrt[15] ), .A2(new_n14836_), .ZN(new_n14837_));
  XOR2_X1    g14645(.A1(new_n14837_), .A2(new_n14637_), .Z(new_n14838_));
  INV_X1     g14646(.I(new_n14838_), .ZN(new_n14839_));
  INV_X1     g14647(.I(\a[30] ), .ZN(new_n14840_));
  NOR2_X1    g14648(.A1(\a[28] ), .A2(\a[29] ), .ZN(new_n14841_));
  INV_X1     g14649(.I(new_n14841_), .ZN(new_n14842_));
  NOR3_X1    g14650(.A1(new_n14284_), .A2(new_n14840_), .A3(new_n14842_), .ZN(new_n14843_));
  NAND2_X1   g14651(.A1(new_n14297_), .A2(new_n14843_), .ZN(new_n14844_));
  XOR2_X1    g14652(.A1(new_n14844_), .A2(\a[31] ), .Z(new_n14845_));
  INV_X1     g14653(.I(\a[31] ), .ZN(new_n14846_));
  NOR4_X1    g14654(.A1(new_n14832_), .A2(new_n14821_), .A3(new_n14846_), .A4(new_n14833_), .ZN(new_n14847_));
  NOR2_X1    g14655(.A1(new_n14846_), .A2(\a[30] ), .ZN(new_n14848_));
  OAI21_X1   g14656(.A1(new_n14847_), .A2(new_n14848_), .B(new_n14845_), .ZN(new_n14849_));
  INV_X1     g14657(.I(new_n14845_), .ZN(new_n14850_));
  NOR2_X1    g14658(.A1(new_n14828_), .A2(new_n14627_), .ZN(new_n14851_));
  NOR3_X1    g14659(.A1(new_n14829_), .A2(new_n229_), .A3(new_n14815_), .ZN(new_n14852_));
  AOI21_X1   g14660(.A1(new_n14852_), .A2(new_n14851_), .B(new_n14646_), .ZN(new_n14853_));
  INV_X1     g14661(.I(new_n14820_), .ZN(new_n14854_));
  AOI21_X1   g14662(.A1(new_n14853_), .A2(new_n14854_), .B(new_n14826_), .ZN(new_n14855_));
  AOI21_X1   g14663(.A1(new_n14830_), .A2(\asqrt[62] ), .B(new_n14643_), .ZN(new_n14856_));
  AOI21_X1   g14664(.A1(new_n14802_), .A2(new_n14804_), .B(new_n275_), .ZN(new_n14857_));
  OAI21_X1   g14665(.A1(new_n14805_), .A2(new_n14857_), .B(\asqrt[61] ), .ZN(new_n14858_));
  NAND4_X1   g14666(.A1(new_n14813_), .A2(new_n196_), .A3(new_n14858_), .A4(new_n14814_), .ZN(new_n14859_));
  NOR3_X1    g14667(.A1(new_n14856_), .A2(new_n14824_), .A3(new_n14859_), .ZN(new_n14860_));
  INV_X1     g14668(.I(new_n14833_), .ZN(new_n14861_));
  NAND4_X1   g14669(.A1(new_n14860_), .A2(\a[31] ), .A3(new_n14855_), .A4(new_n14861_), .ZN(new_n14862_));
  NAND3_X1   g14670(.A1(new_n14862_), .A2(\a[30] ), .A3(new_n14850_), .ZN(new_n14863_));
  NAND2_X1   g14671(.A1(new_n14849_), .A2(new_n14863_), .ZN(new_n14864_));
  NOR2_X1    g14672(.A1(new_n14832_), .A2(new_n14821_), .ZN(new_n14865_));
  NAND4_X1   g14673(.A1(new_n14263_), .A2(new_n14255_), .A3(new_n13728_), .A4(new_n14296_), .ZN(new_n14866_));
  NOR2_X1    g14674(.A1(new_n14273_), .A2(new_n14840_), .ZN(new_n14867_));
  XOR2_X1    g14675(.A1(new_n14867_), .A2(new_n14866_), .Z(new_n14868_));
  NOR2_X1    g14676(.A1(new_n14868_), .A2(new_n14842_), .ZN(new_n14869_));
  INV_X1     g14677(.I(new_n14869_), .ZN(new_n14870_));
  NAND3_X1   g14678(.A1(new_n14860_), .A2(new_n14855_), .A3(new_n14861_), .ZN(new_n14871_));
  NOR4_X1    g14679(.A1(new_n14858_), .A2(new_n14627_), .A3(new_n14828_), .A4(new_n14815_), .ZN(new_n14872_));
  NOR3_X1    g14680(.A1(new_n14872_), .A2(new_n14646_), .A3(new_n14820_), .ZN(new_n14873_));
  AOI22_X1   g14681(.A1(new_n14835_), .A2(\asqrt[61] ), .B1(new_n14812_), .B2(new_n14805_), .ZN(new_n14874_));
  NAND4_X1   g14682(.A1(new_n14874_), .A2(new_n196_), .A3(new_n14643_), .A4(new_n14814_), .ZN(new_n14875_));
  OAI21_X1   g14683(.A1(new_n14873_), .A2(new_n14826_), .B(new_n14875_), .ZN(new_n14876_));
  NOR2_X1    g14684(.A1(new_n14825_), .A2(new_n14861_), .ZN(new_n14877_));
  NAND2_X1   g14685(.A1(new_n14877_), .A2(\asqrt[16] ), .ZN(new_n14878_));
  OAI21_X1   g14686(.A1(new_n14876_), .A2(new_n14878_), .B(new_n13694_), .ZN(new_n14879_));
  NAND3_X1   g14687(.A1(new_n14879_), .A2(new_n13702_), .A3(new_n14871_), .ZN(new_n14880_));
  NAND4_X1   g14688(.A1(new_n14637_), .A2(new_n14805_), .A3(new_n14812_), .A4(new_n14816_), .ZN(new_n14881_));
  NAND3_X1   g14689(.A1(new_n14881_), .A2(new_n14647_), .A3(new_n14854_), .ZN(new_n14882_));
  AOI21_X1   g14690(.A1(new_n14643_), .A2(new_n14882_), .B(new_n14831_), .ZN(new_n14883_));
  INV_X1     g14691(.I(new_n14878_), .ZN(new_n14884_));
  AOI21_X1   g14692(.A1(new_n14883_), .A2(new_n14884_), .B(\a[32] ), .ZN(new_n14885_));
  OAI21_X1   g14693(.A1(new_n14885_), .A2(new_n13703_), .B(\asqrt[15] ), .ZN(new_n14886_));
  NAND4_X1   g14694(.A1(new_n14880_), .A2(new_n14886_), .A3(new_n13760_), .A4(new_n14870_), .ZN(new_n14887_));
  NAND2_X1   g14695(.A1(new_n14887_), .A2(new_n14864_), .ZN(new_n14888_));
  NAND3_X1   g14696(.A1(new_n14849_), .A2(new_n14863_), .A3(new_n14870_), .ZN(new_n14889_));
  INV_X1     g14697(.I(new_n13705_), .ZN(new_n14890_));
  NOR2_X1    g14698(.A1(new_n14273_), .A2(\a[32] ), .ZN(new_n14891_));
  OAI22_X1   g14699(.A1(new_n14891_), .A2(\a[33] ), .B1(\a[32] ), .B2(new_n14264_), .ZN(new_n14892_));
  NAND2_X1   g14700(.A1(\asqrt[16] ), .A2(\a[32] ), .ZN(new_n14893_));
  AND3_X2    g14701(.A1(new_n14892_), .A2(new_n14890_), .A3(new_n14893_), .Z(new_n14894_));
  NAND3_X1   g14702(.A1(\asqrt[15] ), .A2(new_n14272_), .A3(new_n14894_), .ZN(new_n14895_));
  INV_X1     g14703(.I(new_n14894_), .ZN(new_n14896_));
  OAI21_X1   g14704(.A1(new_n14871_), .A2(new_n14896_), .B(new_n14271_), .ZN(new_n14897_));
  NAND3_X1   g14705(.A1(new_n14895_), .A2(new_n14897_), .A3(new_n13192_), .ZN(new_n14898_));
  AOI21_X1   g14706(.A1(new_n14889_), .A2(\asqrt[17] ), .B(new_n14898_), .ZN(new_n14899_));
  NOR2_X1    g14707(.A1(new_n14888_), .A2(new_n14899_), .ZN(new_n14900_));
  AOI22_X1   g14708(.A1(new_n14887_), .A2(new_n14864_), .B1(\asqrt[17] ), .B2(new_n14889_), .ZN(new_n14901_));
  AOI21_X1   g14709(.A1(new_n14300_), .A2(new_n14287_), .B(\asqrt[18] ), .ZN(new_n14902_));
  AND4_X2    g14710(.A1(new_n14658_), .A2(\asqrt[15] ), .A3(new_n14314_), .A4(new_n14902_), .Z(new_n14903_));
  NOR2_X1    g14711(.A1(new_n14658_), .A2(new_n13192_), .ZN(new_n14904_));
  NOR3_X1    g14712(.A1(new_n14903_), .A2(\asqrt[19] ), .A3(new_n14904_), .ZN(new_n14905_));
  OAI21_X1   g14713(.A1(new_n14901_), .A2(new_n13192_), .B(new_n14905_), .ZN(new_n14906_));
  NAND2_X1   g14714(.A1(new_n14906_), .A2(new_n14900_), .ZN(new_n14907_));
  OAI22_X1   g14715(.A1(new_n14901_), .A2(new_n13192_), .B1(new_n14888_), .B2(new_n14899_), .ZN(new_n14908_));
  NAND2_X1   g14716(.A1(new_n14309_), .A2(new_n14310_), .ZN(new_n14909_));
  NAND4_X1   g14717(.A1(\asqrt[15] ), .A2(new_n12657_), .A3(new_n14909_), .A4(new_n14348_), .ZN(new_n14910_));
  XOR2_X1    g14718(.A1(new_n14910_), .A2(new_n14315_), .Z(new_n14911_));
  NAND2_X1   g14719(.A1(new_n14911_), .A2(new_n12101_), .ZN(new_n14912_));
  AOI21_X1   g14720(.A1(new_n14908_), .A2(\asqrt[19] ), .B(new_n14912_), .ZN(new_n14913_));
  NOR2_X1    g14721(.A1(new_n14913_), .A2(new_n14907_), .ZN(new_n14914_));
  AOI22_X1   g14722(.A1(new_n14908_), .A2(\asqrt[19] ), .B1(new_n14906_), .B2(new_n14900_), .ZN(new_n14915_));
  NOR2_X1    g14723(.A1(new_n14322_), .A2(new_n14320_), .ZN(new_n14916_));
  NOR4_X1    g14724(.A1(new_n14871_), .A2(\asqrt[20] ), .A3(new_n14916_), .A4(new_n14350_), .ZN(new_n14917_));
  XOR2_X1    g14725(.A1(new_n14917_), .A2(new_n14326_), .Z(new_n14918_));
  NAND2_X1   g14726(.A1(new_n14918_), .A2(new_n11631_), .ZN(new_n14919_));
  INV_X1     g14727(.I(new_n14919_), .ZN(new_n14920_));
  OAI21_X1   g14728(.A1(new_n14915_), .A2(new_n12101_), .B(new_n14920_), .ZN(new_n14921_));
  NAND2_X1   g14729(.A1(new_n14921_), .A2(new_n14914_), .ZN(new_n14922_));
  OAI22_X1   g14730(.A1(new_n14915_), .A2(new_n12101_), .B1(new_n14913_), .B2(new_n14907_), .ZN(new_n14923_));
  NOR4_X1    g14731(.A1(new_n14871_), .A2(\asqrt[21] ), .A3(new_n14330_), .A4(new_n14667_), .ZN(new_n14924_));
  XNOR2_X1   g14732(.A1(new_n14924_), .A2(new_n14334_), .ZN(new_n14925_));
  NAND2_X1   g14733(.A1(new_n14925_), .A2(new_n11105_), .ZN(new_n14926_));
  AOI21_X1   g14734(.A1(new_n14923_), .A2(\asqrt[21] ), .B(new_n14926_), .ZN(new_n14927_));
  NOR2_X1    g14735(.A1(new_n14927_), .A2(new_n14922_), .ZN(new_n14928_));
  AOI22_X1   g14736(.A1(new_n14923_), .A2(\asqrt[21] ), .B1(new_n14921_), .B2(new_n14914_), .ZN(new_n14929_));
  NOR4_X1    g14737(.A1(new_n14871_), .A2(\asqrt[22] ), .A3(new_n14338_), .A4(new_n14355_), .ZN(new_n14930_));
  XOR2_X1    g14738(.A1(new_n14930_), .A2(new_n14341_), .Z(new_n14931_));
  NAND2_X1   g14739(.A1(new_n14931_), .A2(new_n10614_), .ZN(new_n14932_));
  INV_X1     g14740(.I(new_n14932_), .ZN(new_n14933_));
  OAI21_X1   g14741(.A1(new_n14929_), .A2(new_n11105_), .B(new_n14933_), .ZN(new_n14934_));
  NAND2_X1   g14742(.A1(new_n14934_), .A2(new_n14928_), .ZN(new_n14935_));
  OAI22_X1   g14743(.A1(new_n14929_), .A2(new_n11105_), .B1(new_n14927_), .B2(new_n14922_), .ZN(new_n14936_));
  NOR4_X1    g14744(.A1(new_n14871_), .A2(\asqrt[23] ), .A3(new_n14344_), .A4(new_n14673_), .ZN(new_n14937_));
  XNOR2_X1   g14745(.A1(new_n14937_), .A2(new_n14676_), .ZN(new_n14938_));
  NAND2_X1   g14746(.A1(new_n14938_), .A2(new_n10104_), .ZN(new_n14939_));
  AOI21_X1   g14747(.A1(new_n14936_), .A2(\asqrt[23] ), .B(new_n14939_), .ZN(new_n14940_));
  NOR2_X1    g14748(.A1(new_n14940_), .A2(new_n14935_), .ZN(new_n14941_));
  AOI22_X1   g14749(.A1(new_n14936_), .A2(\asqrt[23] ), .B1(new_n14934_), .B2(new_n14928_), .ZN(new_n14942_));
  NOR4_X1    g14750(.A1(new_n14871_), .A2(\asqrt[24] ), .A3(new_n14359_), .A4(new_n14365_), .ZN(new_n14943_));
  XOR2_X1    g14751(.A1(new_n14943_), .A2(new_n14677_), .Z(new_n14944_));
  NAND2_X1   g14752(.A1(new_n14944_), .A2(new_n9672_), .ZN(new_n14945_));
  INV_X1     g14753(.I(new_n14945_), .ZN(new_n14946_));
  OAI21_X1   g14754(.A1(new_n14942_), .A2(new_n10104_), .B(new_n14946_), .ZN(new_n14947_));
  NAND2_X1   g14755(.A1(new_n14947_), .A2(new_n14941_), .ZN(new_n14948_));
  OAI22_X1   g14756(.A1(new_n14942_), .A2(new_n10104_), .B1(new_n14940_), .B2(new_n14935_), .ZN(new_n14949_));
  NAND2_X1   g14757(.A1(new_n14682_), .A2(\asqrt[25] ), .ZN(new_n14950_));
  NOR4_X1    g14758(.A1(new_n14871_), .A2(\asqrt[25] ), .A3(new_n14368_), .A4(new_n14682_), .ZN(new_n14951_));
  XOR2_X1    g14759(.A1(new_n14951_), .A2(new_n14950_), .Z(new_n14952_));
  NAND2_X1   g14760(.A1(new_n14952_), .A2(new_n9212_), .ZN(new_n14953_));
  AOI21_X1   g14761(.A1(new_n14949_), .A2(\asqrt[25] ), .B(new_n14953_), .ZN(new_n14954_));
  NOR2_X1    g14762(.A1(new_n14954_), .A2(new_n14948_), .ZN(new_n14955_));
  AOI22_X1   g14763(.A1(new_n14949_), .A2(\asqrt[25] ), .B1(new_n14947_), .B2(new_n14941_), .ZN(new_n14956_));
  NOR4_X1    g14764(.A1(new_n14871_), .A2(\asqrt[26] ), .A3(new_n14375_), .A4(new_n14380_), .ZN(new_n14957_));
  AOI21_X1   g14765(.A1(new_n14950_), .A2(new_n14680_), .B(new_n9212_), .ZN(new_n14958_));
  NOR2_X1    g14766(.A1(new_n14957_), .A2(new_n14958_), .ZN(new_n14959_));
  NAND2_X1   g14767(.A1(new_n14959_), .A2(new_n8763_), .ZN(new_n14960_));
  INV_X1     g14768(.I(new_n14960_), .ZN(new_n14961_));
  OAI21_X1   g14769(.A1(new_n14956_), .A2(new_n9212_), .B(new_n14961_), .ZN(new_n14962_));
  NAND2_X1   g14770(.A1(new_n14962_), .A2(new_n14955_), .ZN(new_n14963_));
  OAI22_X1   g14771(.A1(new_n14956_), .A2(new_n9212_), .B1(new_n14954_), .B2(new_n14948_), .ZN(new_n14964_));
  NAND2_X1   g14772(.A1(new_n14689_), .A2(\asqrt[27] ), .ZN(new_n14965_));
  NOR4_X1    g14773(.A1(new_n14871_), .A2(\asqrt[27] ), .A3(new_n14383_), .A4(new_n14689_), .ZN(new_n14966_));
  XOR2_X1    g14774(.A1(new_n14966_), .A2(new_n14965_), .Z(new_n14967_));
  NAND2_X1   g14775(.A1(new_n14967_), .A2(new_n8319_), .ZN(new_n14968_));
  AOI21_X1   g14776(.A1(new_n14964_), .A2(\asqrt[27] ), .B(new_n14968_), .ZN(new_n14969_));
  NOR2_X1    g14777(.A1(new_n14969_), .A2(new_n14963_), .ZN(new_n14970_));
  AOI22_X1   g14778(.A1(new_n14964_), .A2(\asqrt[27] ), .B1(new_n14962_), .B2(new_n14955_), .ZN(new_n14971_));
  NOR4_X1    g14779(.A1(new_n14871_), .A2(\asqrt[28] ), .A3(new_n14390_), .A4(new_n14395_), .ZN(new_n14972_));
  AOI21_X1   g14780(.A1(new_n14965_), .A2(new_n14688_), .B(new_n8319_), .ZN(new_n14973_));
  NOR2_X1    g14781(.A1(new_n14972_), .A2(new_n14973_), .ZN(new_n14974_));
  NAND2_X1   g14782(.A1(new_n14974_), .A2(new_n7931_), .ZN(new_n14975_));
  INV_X1     g14783(.I(new_n14975_), .ZN(new_n14976_));
  OAI21_X1   g14784(.A1(new_n14971_), .A2(new_n8319_), .B(new_n14976_), .ZN(new_n14977_));
  NAND2_X1   g14785(.A1(new_n14977_), .A2(new_n14970_), .ZN(new_n14978_));
  OAI22_X1   g14786(.A1(new_n14971_), .A2(new_n8319_), .B1(new_n14969_), .B2(new_n14963_), .ZN(new_n14979_));
  NAND2_X1   g14787(.A1(new_n14696_), .A2(\asqrt[29] ), .ZN(new_n14980_));
  NOR4_X1    g14788(.A1(new_n14871_), .A2(\asqrt[29] ), .A3(new_n14398_), .A4(new_n14696_), .ZN(new_n14981_));
  XOR2_X1    g14789(.A1(new_n14981_), .A2(new_n14980_), .Z(new_n14982_));
  NAND2_X1   g14790(.A1(new_n14982_), .A2(new_n7517_), .ZN(new_n14983_));
  AOI21_X1   g14791(.A1(new_n14979_), .A2(\asqrt[29] ), .B(new_n14983_), .ZN(new_n14984_));
  NOR2_X1    g14792(.A1(new_n14984_), .A2(new_n14978_), .ZN(new_n14985_));
  AOI22_X1   g14793(.A1(new_n14979_), .A2(\asqrt[29] ), .B1(new_n14977_), .B2(new_n14970_), .ZN(new_n14986_));
  NOR4_X1    g14794(.A1(new_n14871_), .A2(\asqrt[30] ), .A3(new_n14405_), .A4(new_n14410_), .ZN(new_n14987_));
  AOI21_X1   g14795(.A1(new_n14980_), .A2(new_n14695_), .B(new_n7517_), .ZN(new_n14988_));
  NOR2_X1    g14796(.A1(new_n14987_), .A2(new_n14988_), .ZN(new_n14989_));
  NAND2_X1   g14797(.A1(new_n14989_), .A2(new_n7110_), .ZN(new_n14990_));
  INV_X1     g14798(.I(new_n14990_), .ZN(new_n14991_));
  OAI21_X1   g14799(.A1(new_n14986_), .A2(new_n7517_), .B(new_n14991_), .ZN(new_n14992_));
  NAND2_X1   g14800(.A1(new_n14992_), .A2(new_n14985_), .ZN(new_n14993_));
  OAI22_X1   g14801(.A1(new_n14986_), .A2(new_n7517_), .B1(new_n14984_), .B2(new_n14978_), .ZN(new_n14994_));
  NAND2_X1   g14802(.A1(new_n14703_), .A2(\asqrt[31] ), .ZN(new_n14995_));
  NOR4_X1    g14803(.A1(new_n14871_), .A2(\asqrt[31] ), .A3(new_n14413_), .A4(new_n14703_), .ZN(new_n14996_));
  XOR2_X1    g14804(.A1(new_n14996_), .A2(new_n14995_), .Z(new_n14997_));
  NAND2_X1   g14805(.A1(new_n14997_), .A2(new_n6708_), .ZN(new_n14998_));
  AOI21_X1   g14806(.A1(new_n14994_), .A2(\asqrt[31] ), .B(new_n14998_), .ZN(new_n14999_));
  NOR2_X1    g14807(.A1(new_n14999_), .A2(new_n14993_), .ZN(new_n15000_));
  AOI22_X1   g14808(.A1(new_n14994_), .A2(\asqrt[31] ), .B1(new_n14992_), .B2(new_n14985_), .ZN(new_n15001_));
  NOR4_X1    g14809(.A1(new_n14871_), .A2(\asqrt[32] ), .A3(new_n14420_), .A4(new_n14425_), .ZN(new_n15002_));
  AOI21_X1   g14810(.A1(new_n14995_), .A2(new_n14702_), .B(new_n6708_), .ZN(new_n15003_));
  NOR2_X1    g14811(.A1(new_n15002_), .A2(new_n15003_), .ZN(new_n15004_));
  NAND2_X1   g14812(.A1(new_n15004_), .A2(new_n6365_), .ZN(new_n15005_));
  INV_X1     g14813(.I(new_n15005_), .ZN(new_n15006_));
  OAI21_X1   g14814(.A1(new_n15001_), .A2(new_n6708_), .B(new_n15006_), .ZN(new_n15007_));
  NAND2_X1   g14815(.A1(new_n15007_), .A2(new_n15000_), .ZN(new_n15008_));
  OAI22_X1   g14816(.A1(new_n15001_), .A2(new_n6708_), .B1(new_n14999_), .B2(new_n14993_), .ZN(new_n15009_));
  NAND2_X1   g14817(.A1(new_n14710_), .A2(\asqrt[33] ), .ZN(new_n15010_));
  NOR4_X1    g14818(.A1(new_n14871_), .A2(\asqrt[33] ), .A3(new_n14428_), .A4(new_n14710_), .ZN(new_n15011_));
  XOR2_X1    g14819(.A1(new_n15011_), .A2(new_n15010_), .Z(new_n15012_));
  NAND2_X1   g14820(.A1(new_n15012_), .A2(new_n5991_), .ZN(new_n15013_));
  AOI21_X1   g14821(.A1(new_n15009_), .A2(\asqrt[33] ), .B(new_n15013_), .ZN(new_n15014_));
  NOR2_X1    g14822(.A1(new_n15014_), .A2(new_n15008_), .ZN(new_n15015_));
  AOI22_X1   g14823(.A1(new_n15009_), .A2(\asqrt[33] ), .B1(new_n15007_), .B2(new_n15000_), .ZN(new_n15016_));
  NOR4_X1    g14824(.A1(new_n14871_), .A2(\asqrt[34] ), .A3(new_n14435_), .A4(new_n14440_), .ZN(new_n15017_));
  AOI21_X1   g14825(.A1(new_n15010_), .A2(new_n14709_), .B(new_n5991_), .ZN(new_n15018_));
  NOR2_X1    g14826(.A1(new_n15017_), .A2(new_n15018_), .ZN(new_n15019_));
  NAND2_X1   g14827(.A1(new_n15019_), .A2(new_n5626_), .ZN(new_n15020_));
  INV_X1     g14828(.I(new_n15020_), .ZN(new_n15021_));
  OAI21_X1   g14829(.A1(new_n15016_), .A2(new_n5991_), .B(new_n15021_), .ZN(new_n15022_));
  NAND2_X1   g14830(.A1(new_n15022_), .A2(new_n15015_), .ZN(new_n15023_));
  OAI22_X1   g14831(.A1(new_n15016_), .A2(new_n5991_), .B1(new_n15014_), .B2(new_n15008_), .ZN(new_n15024_));
  NAND2_X1   g14832(.A1(new_n14717_), .A2(\asqrt[35] ), .ZN(new_n15025_));
  NOR4_X1    g14833(.A1(new_n14871_), .A2(\asqrt[35] ), .A3(new_n14443_), .A4(new_n14717_), .ZN(new_n15026_));
  XOR2_X1    g14834(.A1(new_n15026_), .A2(new_n15025_), .Z(new_n15027_));
  NAND2_X1   g14835(.A1(new_n15027_), .A2(new_n5273_), .ZN(new_n15028_));
  AOI21_X1   g14836(.A1(new_n15024_), .A2(\asqrt[35] ), .B(new_n15028_), .ZN(new_n15029_));
  NOR2_X1    g14837(.A1(new_n15029_), .A2(new_n15023_), .ZN(new_n15030_));
  AOI22_X1   g14838(.A1(new_n15024_), .A2(\asqrt[35] ), .B1(new_n15022_), .B2(new_n15015_), .ZN(new_n15031_));
  NAND2_X1   g14839(.A1(new_n14455_), .A2(\asqrt[36] ), .ZN(new_n15032_));
  NOR4_X1    g14840(.A1(new_n14871_), .A2(\asqrt[36] ), .A3(new_n14450_), .A4(new_n14455_), .ZN(new_n15033_));
  XOR2_X1    g14841(.A1(new_n15033_), .A2(new_n15032_), .Z(new_n15034_));
  NAND2_X1   g14842(.A1(new_n15034_), .A2(new_n4973_), .ZN(new_n15035_));
  INV_X1     g14843(.I(new_n15035_), .ZN(new_n15036_));
  OAI21_X1   g14844(.A1(new_n15031_), .A2(new_n5273_), .B(new_n15036_), .ZN(new_n15037_));
  NAND2_X1   g14845(.A1(new_n15037_), .A2(new_n15030_), .ZN(new_n15038_));
  OAI22_X1   g14846(.A1(new_n15031_), .A2(new_n5273_), .B1(new_n15029_), .B2(new_n15023_), .ZN(new_n15039_));
  NOR4_X1    g14847(.A1(new_n14871_), .A2(\asqrt[37] ), .A3(new_n14458_), .A4(new_n14724_), .ZN(new_n15040_));
  AOI21_X1   g14848(.A1(new_n15032_), .A2(new_n14454_), .B(new_n4973_), .ZN(new_n15041_));
  NOR2_X1    g14849(.A1(new_n15040_), .A2(new_n15041_), .ZN(new_n15042_));
  NAND2_X1   g14850(.A1(new_n15042_), .A2(new_n4645_), .ZN(new_n15043_));
  AOI21_X1   g14851(.A1(new_n15039_), .A2(\asqrt[37] ), .B(new_n15043_), .ZN(new_n15044_));
  NOR2_X1    g14852(.A1(new_n15044_), .A2(new_n15038_), .ZN(new_n15045_));
  AOI22_X1   g14853(.A1(new_n15039_), .A2(\asqrt[37] ), .B1(new_n15037_), .B2(new_n15030_), .ZN(new_n15046_));
  NAND2_X1   g14854(.A1(new_n14470_), .A2(\asqrt[38] ), .ZN(new_n15047_));
  NOR4_X1    g14855(.A1(new_n14871_), .A2(\asqrt[38] ), .A3(new_n14465_), .A4(new_n14470_), .ZN(new_n15048_));
  XOR2_X1    g14856(.A1(new_n15048_), .A2(new_n15047_), .Z(new_n15049_));
  NAND2_X1   g14857(.A1(new_n15049_), .A2(new_n4330_), .ZN(new_n15050_));
  INV_X1     g14858(.I(new_n15050_), .ZN(new_n15051_));
  OAI21_X1   g14859(.A1(new_n15046_), .A2(new_n4645_), .B(new_n15051_), .ZN(new_n15052_));
  NAND2_X1   g14860(.A1(new_n15052_), .A2(new_n15045_), .ZN(new_n15053_));
  OAI22_X1   g14861(.A1(new_n15046_), .A2(new_n4645_), .B1(new_n15044_), .B2(new_n15038_), .ZN(new_n15054_));
  NOR4_X1    g14862(.A1(new_n14871_), .A2(\asqrt[39] ), .A3(new_n14473_), .A4(new_n14731_), .ZN(new_n15055_));
  AOI21_X1   g14863(.A1(new_n15047_), .A2(new_n14469_), .B(new_n4330_), .ZN(new_n15056_));
  NOR2_X1    g14864(.A1(new_n15055_), .A2(new_n15056_), .ZN(new_n15057_));
  NAND2_X1   g14865(.A1(new_n15057_), .A2(new_n4018_), .ZN(new_n15058_));
  AOI21_X1   g14866(.A1(new_n15054_), .A2(\asqrt[39] ), .B(new_n15058_), .ZN(new_n15059_));
  NOR2_X1    g14867(.A1(new_n15059_), .A2(new_n15053_), .ZN(new_n15060_));
  AOI22_X1   g14868(.A1(new_n15054_), .A2(\asqrt[39] ), .B1(new_n15052_), .B2(new_n15045_), .ZN(new_n15061_));
  NAND2_X1   g14869(.A1(new_n14485_), .A2(\asqrt[40] ), .ZN(new_n15062_));
  NOR4_X1    g14870(.A1(new_n14871_), .A2(\asqrt[40] ), .A3(new_n14480_), .A4(new_n14485_), .ZN(new_n15063_));
  XOR2_X1    g14871(.A1(new_n15063_), .A2(new_n15062_), .Z(new_n15064_));
  NAND2_X1   g14872(.A1(new_n15064_), .A2(new_n3760_), .ZN(new_n15065_));
  INV_X1     g14873(.I(new_n15065_), .ZN(new_n15066_));
  OAI21_X1   g14874(.A1(new_n15061_), .A2(new_n4018_), .B(new_n15066_), .ZN(new_n15067_));
  NAND2_X1   g14875(.A1(new_n15067_), .A2(new_n15060_), .ZN(new_n15068_));
  OAI22_X1   g14876(.A1(new_n15061_), .A2(new_n4018_), .B1(new_n15059_), .B2(new_n15053_), .ZN(new_n15069_));
  NAND2_X1   g14877(.A1(new_n14738_), .A2(\asqrt[41] ), .ZN(new_n15070_));
  NOR4_X1    g14878(.A1(new_n14871_), .A2(\asqrt[41] ), .A3(new_n14488_), .A4(new_n14738_), .ZN(new_n15071_));
  XOR2_X1    g14879(.A1(new_n15071_), .A2(new_n15070_), .Z(new_n15072_));
  NAND2_X1   g14880(.A1(new_n15072_), .A2(new_n3481_), .ZN(new_n15073_));
  AOI21_X1   g14881(.A1(new_n15069_), .A2(\asqrt[41] ), .B(new_n15073_), .ZN(new_n15074_));
  NOR2_X1    g14882(.A1(new_n15074_), .A2(new_n15068_), .ZN(new_n15075_));
  AOI22_X1   g14883(.A1(new_n15069_), .A2(\asqrt[41] ), .B1(new_n15067_), .B2(new_n15060_), .ZN(new_n15076_));
  NOR4_X1    g14884(.A1(new_n14871_), .A2(\asqrt[42] ), .A3(new_n14495_), .A4(new_n14500_), .ZN(new_n15077_));
  AOI21_X1   g14885(.A1(new_n15070_), .A2(new_n14737_), .B(new_n3481_), .ZN(new_n15078_));
  NOR2_X1    g14886(.A1(new_n15077_), .A2(new_n15078_), .ZN(new_n15079_));
  NAND2_X1   g14887(.A1(new_n15079_), .A2(new_n3208_), .ZN(new_n15080_));
  INV_X1     g14888(.I(new_n15080_), .ZN(new_n15081_));
  OAI21_X1   g14889(.A1(new_n15076_), .A2(new_n3481_), .B(new_n15081_), .ZN(new_n15082_));
  NAND2_X1   g14890(.A1(new_n15082_), .A2(new_n15075_), .ZN(new_n15083_));
  OAI22_X1   g14891(.A1(new_n15076_), .A2(new_n3481_), .B1(new_n15074_), .B2(new_n15068_), .ZN(new_n15084_));
  NAND2_X1   g14892(.A1(new_n14745_), .A2(\asqrt[43] ), .ZN(new_n15085_));
  NOR4_X1    g14893(.A1(new_n14871_), .A2(\asqrt[43] ), .A3(new_n14503_), .A4(new_n14745_), .ZN(new_n15086_));
  XOR2_X1    g14894(.A1(new_n15086_), .A2(new_n15085_), .Z(new_n15087_));
  NAND2_X1   g14895(.A1(new_n15087_), .A2(new_n2941_), .ZN(new_n15088_));
  AOI21_X1   g14896(.A1(new_n15084_), .A2(\asqrt[43] ), .B(new_n15088_), .ZN(new_n15089_));
  NOR2_X1    g14897(.A1(new_n15089_), .A2(new_n15083_), .ZN(new_n15090_));
  AOI22_X1   g14898(.A1(new_n15084_), .A2(\asqrt[43] ), .B1(new_n15082_), .B2(new_n15075_), .ZN(new_n15091_));
  NOR4_X1    g14899(.A1(new_n14871_), .A2(\asqrt[44] ), .A3(new_n14510_), .A4(new_n14515_), .ZN(new_n15092_));
  AOI21_X1   g14900(.A1(new_n15085_), .A2(new_n14744_), .B(new_n2941_), .ZN(new_n15093_));
  NOR2_X1    g14901(.A1(new_n15092_), .A2(new_n15093_), .ZN(new_n15094_));
  NAND2_X1   g14902(.A1(new_n15094_), .A2(new_n2728_), .ZN(new_n15095_));
  INV_X1     g14903(.I(new_n15095_), .ZN(new_n15096_));
  OAI21_X1   g14904(.A1(new_n15091_), .A2(new_n2941_), .B(new_n15096_), .ZN(new_n15097_));
  NAND2_X1   g14905(.A1(new_n15097_), .A2(new_n15090_), .ZN(new_n15098_));
  OAI22_X1   g14906(.A1(new_n15091_), .A2(new_n2941_), .B1(new_n15089_), .B2(new_n15083_), .ZN(new_n15099_));
  NAND2_X1   g14907(.A1(new_n14752_), .A2(\asqrt[45] ), .ZN(new_n15100_));
  NOR4_X1    g14908(.A1(new_n14871_), .A2(\asqrt[45] ), .A3(new_n14518_), .A4(new_n14752_), .ZN(new_n15101_));
  XOR2_X1    g14909(.A1(new_n15101_), .A2(new_n15100_), .Z(new_n15102_));
  NAND2_X1   g14910(.A1(new_n15102_), .A2(new_n2488_), .ZN(new_n15103_));
  AOI21_X1   g14911(.A1(new_n15099_), .A2(\asqrt[45] ), .B(new_n15103_), .ZN(new_n15104_));
  NOR2_X1    g14912(.A1(new_n15104_), .A2(new_n15098_), .ZN(new_n15105_));
  AOI22_X1   g14913(.A1(new_n15099_), .A2(\asqrt[45] ), .B1(new_n15097_), .B2(new_n15090_), .ZN(new_n15106_));
  NOR4_X1    g14914(.A1(new_n14871_), .A2(\asqrt[46] ), .A3(new_n14525_), .A4(new_n14530_), .ZN(new_n15107_));
  AOI21_X1   g14915(.A1(new_n15100_), .A2(new_n14751_), .B(new_n2488_), .ZN(new_n15108_));
  NOR2_X1    g14916(.A1(new_n15107_), .A2(new_n15108_), .ZN(new_n15109_));
  NAND2_X1   g14917(.A1(new_n15109_), .A2(new_n2253_), .ZN(new_n15110_));
  INV_X1     g14918(.I(new_n15110_), .ZN(new_n15111_));
  OAI21_X1   g14919(.A1(new_n15106_), .A2(new_n2488_), .B(new_n15111_), .ZN(new_n15112_));
  NAND2_X1   g14920(.A1(new_n15112_), .A2(new_n15105_), .ZN(new_n15113_));
  OAI22_X1   g14921(.A1(new_n15106_), .A2(new_n2488_), .B1(new_n15104_), .B2(new_n15098_), .ZN(new_n15114_));
  NAND2_X1   g14922(.A1(new_n14759_), .A2(\asqrt[47] ), .ZN(new_n15115_));
  NOR4_X1    g14923(.A1(new_n14871_), .A2(\asqrt[47] ), .A3(new_n14533_), .A4(new_n14759_), .ZN(new_n15116_));
  XOR2_X1    g14924(.A1(new_n15116_), .A2(new_n15115_), .Z(new_n15117_));
  NAND2_X1   g14925(.A1(new_n15117_), .A2(new_n2046_), .ZN(new_n15118_));
  AOI21_X1   g14926(.A1(new_n15114_), .A2(\asqrt[47] ), .B(new_n15118_), .ZN(new_n15119_));
  NOR2_X1    g14927(.A1(new_n15119_), .A2(new_n15113_), .ZN(new_n15120_));
  AOI22_X1   g14928(.A1(new_n15114_), .A2(\asqrt[47] ), .B1(new_n15112_), .B2(new_n15105_), .ZN(new_n15121_));
  NAND2_X1   g14929(.A1(new_n14545_), .A2(\asqrt[48] ), .ZN(new_n15122_));
  NOR4_X1    g14930(.A1(new_n14871_), .A2(\asqrt[48] ), .A3(new_n14540_), .A4(new_n14545_), .ZN(new_n15123_));
  XOR2_X1    g14931(.A1(new_n15123_), .A2(new_n15122_), .Z(new_n15124_));
  NAND2_X1   g14932(.A1(new_n15124_), .A2(new_n1854_), .ZN(new_n15125_));
  INV_X1     g14933(.I(new_n15125_), .ZN(new_n15126_));
  OAI21_X1   g14934(.A1(new_n15121_), .A2(new_n2046_), .B(new_n15126_), .ZN(new_n15127_));
  NAND2_X1   g14935(.A1(new_n15127_), .A2(new_n15120_), .ZN(new_n15128_));
  OAI22_X1   g14936(.A1(new_n15121_), .A2(new_n2046_), .B1(new_n15119_), .B2(new_n15113_), .ZN(new_n15129_));
  NOR4_X1    g14937(.A1(new_n14871_), .A2(\asqrt[49] ), .A3(new_n14548_), .A4(new_n14766_), .ZN(new_n15130_));
  AOI21_X1   g14938(.A1(new_n15122_), .A2(new_n14544_), .B(new_n1854_), .ZN(new_n15131_));
  NOR2_X1    g14939(.A1(new_n15130_), .A2(new_n15131_), .ZN(new_n15132_));
  NAND2_X1   g14940(.A1(new_n15132_), .A2(new_n1595_), .ZN(new_n15133_));
  AOI21_X1   g14941(.A1(new_n15129_), .A2(\asqrt[49] ), .B(new_n15133_), .ZN(new_n15134_));
  NOR2_X1    g14942(.A1(new_n15134_), .A2(new_n15128_), .ZN(new_n15135_));
  AOI22_X1   g14943(.A1(new_n15129_), .A2(\asqrt[49] ), .B1(new_n15127_), .B2(new_n15120_), .ZN(new_n15136_));
  NAND2_X1   g14944(.A1(new_n14560_), .A2(\asqrt[50] ), .ZN(new_n15137_));
  NOR4_X1    g14945(.A1(new_n14871_), .A2(\asqrt[50] ), .A3(new_n14555_), .A4(new_n14560_), .ZN(new_n15138_));
  XOR2_X1    g14946(.A1(new_n15138_), .A2(new_n15137_), .Z(new_n15139_));
  NAND2_X1   g14947(.A1(new_n15139_), .A2(new_n1436_), .ZN(new_n15140_));
  INV_X1     g14948(.I(new_n15140_), .ZN(new_n15141_));
  OAI21_X1   g14949(.A1(new_n15136_), .A2(new_n1595_), .B(new_n15141_), .ZN(new_n15142_));
  NAND2_X1   g14950(.A1(new_n15142_), .A2(new_n15135_), .ZN(new_n15143_));
  OAI22_X1   g14951(.A1(new_n15136_), .A2(new_n1595_), .B1(new_n15134_), .B2(new_n15128_), .ZN(new_n15144_));
  NOR2_X1    g14952(.A1(new_n14567_), .A2(new_n1436_), .ZN(new_n15145_));
  NOR4_X1    g14953(.A1(new_n14871_), .A2(\asqrt[51] ), .A3(new_n14563_), .A4(new_n14773_), .ZN(new_n15146_));
  XNOR2_X1   g14954(.A1(new_n15146_), .A2(new_n15145_), .ZN(new_n15147_));
  NAND2_X1   g14955(.A1(new_n15147_), .A2(new_n1260_), .ZN(new_n15148_));
  AOI21_X1   g14956(.A1(new_n15144_), .A2(\asqrt[51] ), .B(new_n15148_), .ZN(new_n15149_));
  NOR2_X1    g14957(.A1(new_n15149_), .A2(new_n15143_), .ZN(new_n15150_));
  AOI22_X1   g14958(.A1(new_n15144_), .A2(\asqrt[51] ), .B1(new_n15142_), .B2(new_n15135_), .ZN(new_n15151_));
  NOR4_X1    g14959(.A1(new_n14871_), .A2(\asqrt[52] ), .A3(new_n14570_), .A4(new_n14575_), .ZN(new_n15152_));
  XOR2_X1    g14960(.A1(new_n15152_), .A2(new_n14628_), .Z(new_n15153_));
  NAND2_X1   g14961(.A1(new_n15153_), .A2(new_n1096_), .ZN(new_n15154_));
  INV_X1     g14962(.I(new_n15154_), .ZN(new_n15155_));
  OAI21_X1   g14963(.A1(new_n15151_), .A2(new_n1260_), .B(new_n15155_), .ZN(new_n15156_));
  NAND2_X1   g14964(.A1(new_n15156_), .A2(new_n15150_), .ZN(new_n15157_));
  OAI22_X1   g14965(.A1(new_n15151_), .A2(new_n1260_), .B1(new_n15149_), .B2(new_n15143_), .ZN(new_n15158_));
  NOR4_X1    g14966(.A1(new_n14871_), .A2(\asqrt[53] ), .A3(new_n14578_), .A4(new_n14780_), .ZN(new_n15159_));
  XNOR2_X1   g14967(.A1(new_n15159_), .A2(new_n14629_), .ZN(new_n15160_));
  NAND2_X1   g14968(.A1(new_n15160_), .A2(new_n970_), .ZN(new_n15161_));
  AOI21_X1   g14969(.A1(new_n15158_), .A2(\asqrt[53] ), .B(new_n15161_), .ZN(new_n15162_));
  NOR2_X1    g14970(.A1(new_n15162_), .A2(new_n15157_), .ZN(new_n15163_));
  AOI22_X1   g14971(.A1(new_n15158_), .A2(\asqrt[53] ), .B1(new_n15156_), .B2(new_n15150_), .ZN(new_n15164_));
  NOR4_X1    g14972(.A1(new_n14871_), .A2(\asqrt[54] ), .A3(new_n14585_), .A4(new_n14590_), .ZN(new_n15165_));
  XOR2_X1    g14973(.A1(new_n15165_), .A2(new_n14630_), .Z(new_n15166_));
  NAND2_X1   g14974(.A1(new_n15166_), .A2(new_n825_), .ZN(new_n15167_));
  INV_X1     g14975(.I(new_n15167_), .ZN(new_n15168_));
  OAI21_X1   g14976(.A1(new_n15164_), .A2(new_n970_), .B(new_n15168_), .ZN(new_n15169_));
  NAND2_X1   g14977(.A1(new_n15169_), .A2(new_n15163_), .ZN(new_n15170_));
  OAI22_X1   g14978(.A1(new_n15164_), .A2(new_n970_), .B1(new_n15162_), .B2(new_n15157_), .ZN(new_n15171_));
  NOR4_X1    g14979(.A1(new_n14871_), .A2(\asqrt[55] ), .A3(new_n14593_), .A4(new_n14787_), .ZN(new_n15172_));
  XOR2_X1    g14980(.A1(new_n15172_), .A2(new_n14794_), .Z(new_n15173_));
  NAND2_X1   g14981(.A1(new_n15173_), .A2(new_n724_), .ZN(new_n15174_));
  AOI21_X1   g14982(.A1(new_n15171_), .A2(\asqrt[55] ), .B(new_n15174_), .ZN(new_n15175_));
  NOR2_X1    g14983(.A1(new_n15175_), .A2(new_n15170_), .ZN(new_n15176_));
  AOI22_X1   g14984(.A1(new_n15171_), .A2(\asqrt[55] ), .B1(new_n15169_), .B2(new_n15163_), .ZN(new_n15177_));
  NOR4_X1    g14985(.A1(new_n14871_), .A2(\asqrt[56] ), .A3(new_n14599_), .A4(new_n14604_), .ZN(new_n15178_));
  XOR2_X1    g14986(.A1(new_n15178_), .A2(new_n14632_), .Z(new_n15179_));
  NAND2_X1   g14987(.A1(new_n15179_), .A2(new_n587_), .ZN(new_n15180_));
  INV_X1     g14988(.I(new_n15180_), .ZN(new_n15181_));
  OAI21_X1   g14989(.A1(new_n15177_), .A2(new_n724_), .B(new_n15181_), .ZN(new_n15182_));
  NAND2_X1   g14990(.A1(new_n15182_), .A2(new_n15176_), .ZN(new_n15183_));
  OAI22_X1   g14991(.A1(new_n15177_), .A2(new_n724_), .B1(new_n15175_), .B2(new_n15170_), .ZN(new_n15184_));
  NOR4_X1    g14992(.A1(new_n14871_), .A2(\asqrt[57] ), .A3(new_n14606_), .A4(new_n14798_), .ZN(new_n15185_));
  XOR2_X1    g14993(.A1(new_n15185_), .A2(new_n14796_), .Z(new_n15186_));
  NAND2_X1   g14994(.A1(new_n15186_), .A2(new_n504_), .ZN(new_n15187_));
  AOI21_X1   g14995(.A1(new_n15184_), .A2(\asqrt[57] ), .B(new_n15187_), .ZN(new_n15188_));
  NOR2_X1    g14996(.A1(new_n15188_), .A2(new_n15183_), .ZN(new_n15189_));
  AOI22_X1   g14997(.A1(new_n15184_), .A2(\asqrt[57] ), .B1(new_n15182_), .B2(new_n15176_), .ZN(new_n15190_));
  NOR4_X1    g14998(.A1(new_n14871_), .A2(\asqrt[58] ), .A3(new_n14612_), .A4(new_n14616_), .ZN(new_n15191_));
  XOR2_X1    g14999(.A1(new_n15191_), .A2(new_n14634_), .Z(new_n15192_));
  NAND2_X1   g15000(.A1(new_n15192_), .A2(new_n376_), .ZN(new_n15193_));
  INV_X1     g15001(.I(new_n15193_), .ZN(new_n15194_));
  OAI21_X1   g15002(.A1(new_n15190_), .A2(new_n504_), .B(new_n15194_), .ZN(new_n15195_));
  NAND2_X1   g15003(.A1(new_n15195_), .A2(new_n15189_), .ZN(new_n15196_));
  OAI22_X1   g15004(.A1(new_n15190_), .A2(new_n504_), .B1(new_n15188_), .B2(new_n15183_), .ZN(new_n15197_));
  NOR4_X1    g15005(.A1(new_n14871_), .A2(\asqrt[59] ), .A3(new_n14618_), .A4(new_n14806_), .ZN(new_n15198_));
  XOR2_X1    g15006(.A1(new_n15198_), .A2(new_n14804_), .Z(new_n15199_));
  NAND2_X1   g15007(.A1(new_n15199_), .A2(new_n275_), .ZN(new_n15200_));
  AOI21_X1   g15008(.A1(new_n15197_), .A2(\asqrt[59] ), .B(new_n15200_), .ZN(new_n15201_));
  NOR2_X1    g15009(.A1(new_n15201_), .A2(new_n15196_), .ZN(new_n15202_));
  AOI22_X1   g15010(.A1(new_n15197_), .A2(\asqrt[59] ), .B1(new_n15195_), .B2(new_n15189_), .ZN(new_n15203_));
  OAI22_X1   g15011(.A1(new_n15203_), .A2(new_n275_), .B1(new_n15201_), .B2(new_n15196_), .ZN(new_n15204_));
  NOR4_X1    g15012(.A1(new_n14871_), .A2(\asqrt[60] ), .A3(new_n14624_), .A4(new_n14827_), .ZN(new_n15205_));
  XOR2_X1    g15013(.A1(new_n15205_), .A2(new_n14636_), .Z(new_n15206_));
  NAND2_X1   g15014(.A1(new_n15206_), .A2(new_n229_), .ZN(new_n15207_));
  INV_X1     g15015(.I(new_n15207_), .ZN(new_n15208_));
  OAI21_X1   g15016(.A1(new_n15203_), .A2(new_n275_), .B(new_n15208_), .ZN(new_n15209_));
  AOI22_X1   g15017(.A1(new_n15204_), .A2(\asqrt[61] ), .B1(new_n15209_), .B2(new_n15202_), .ZN(new_n15210_));
  NOR2_X1    g15018(.A1(new_n15210_), .A2(new_n196_), .ZN(new_n15211_));
  INV_X1     g15019(.I(new_n14848_), .ZN(new_n15212_));
  AOI21_X1   g15020(.A1(new_n14862_), .A2(new_n15212_), .B(new_n14850_), .ZN(new_n15213_));
  NOR3_X1    g15021(.A1(new_n14847_), .A2(new_n14840_), .A3(new_n14845_), .ZN(new_n15214_));
  NOR2_X1    g15022(.A1(new_n15214_), .A2(new_n15213_), .ZN(new_n15215_));
  NOR3_X1    g15023(.A1(new_n14885_), .A2(new_n13703_), .A3(\asqrt[15] ), .ZN(new_n15216_));
  AOI21_X1   g15024(.A1(new_n14879_), .A2(new_n13702_), .B(new_n14871_), .ZN(new_n15217_));
  NOR4_X1    g15025(.A1(new_n15217_), .A2(new_n15216_), .A3(\asqrt[17] ), .A4(new_n14869_), .ZN(new_n15218_));
  NOR2_X1    g15026(.A1(new_n15218_), .A2(new_n15215_), .ZN(new_n15219_));
  NOR3_X1    g15027(.A1(new_n15214_), .A2(new_n15213_), .A3(new_n14869_), .ZN(new_n15220_));
  NOR3_X1    g15028(.A1(new_n14871_), .A2(new_n14271_), .A3(new_n14896_), .ZN(new_n15221_));
  AOI21_X1   g15029(.A1(\asqrt[15] ), .A2(new_n14894_), .B(new_n14272_), .ZN(new_n15222_));
  NOR3_X1    g15030(.A1(new_n15222_), .A2(new_n15221_), .A3(\asqrt[18] ), .ZN(new_n15223_));
  OAI21_X1   g15031(.A1(new_n15220_), .A2(new_n13760_), .B(new_n15223_), .ZN(new_n15224_));
  NAND2_X1   g15032(.A1(new_n15219_), .A2(new_n15224_), .ZN(new_n15225_));
  OAI22_X1   g15033(.A1(new_n15218_), .A2(new_n15215_), .B1(new_n13760_), .B2(new_n15220_), .ZN(new_n15226_));
  INV_X1     g15034(.I(new_n14905_), .ZN(new_n15227_));
  AOI21_X1   g15035(.A1(new_n15226_), .A2(\asqrt[18] ), .B(new_n15227_), .ZN(new_n15228_));
  NOR2_X1    g15036(.A1(new_n15228_), .A2(new_n15225_), .ZN(new_n15229_));
  AOI22_X1   g15037(.A1(new_n15226_), .A2(\asqrt[18] ), .B1(new_n15219_), .B2(new_n15224_), .ZN(new_n15230_));
  INV_X1     g15038(.I(new_n14912_), .ZN(new_n15231_));
  OAI21_X1   g15039(.A1(new_n15230_), .A2(new_n12657_), .B(new_n15231_), .ZN(new_n15232_));
  NAND2_X1   g15040(.A1(new_n15232_), .A2(new_n15229_), .ZN(new_n15233_));
  OAI22_X1   g15041(.A1(new_n15230_), .A2(new_n12657_), .B1(new_n15228_), .B2(new_n15225_), .ZN(new_n15234_));
  AOI21_X1   g15042(.A1(new_n15234_), .A2(\asqrt[20] ), .B(new_n14919_), .ZN(new_n15235_));
  NOR2_X1    g15043(.A1(new_n15235_), .A2(new_n15233_), .ZN(new_n15236_));
  AOI22_X1   g15044(.A1(new_n15234_), .A2(\asqrt[20] ), .B1(new_n15232_), .B2(new_n15229_), .ZN(new_n15237_));
  INV_X1     g15045(.I(new_n14926_), .ZN(new_n15238_));
  OAI21_X1   g15046(.A1(new_n15237_), .A2(new_n11631_), .B(new_n15238_), .ZN(new_n15239_));
  NAND2_X1   g15047(.A1(new_n15239_), .A2(new_n15236_), .ZN(new_n15240_));
  OAI22_X1   g15048(.A1(new_n15237_), .A2(new_n11631_), .B1(new_n15235_), .B2(new_n15233_), .ZN(new_n15241_));
  AOI21_X1   g15049(.A1(new_n15241_), .A2(\asqrt[22] ), .B(new_n14932_), .ZN(new_n15242_));
  NOR2_X1    g15050(.A1(new_n15242_), .A2(new_n15240_), .ZN(new_n15243_));
  AOI22_X1   g15051(.A1(new_n15241_), .A2(\asqrt[22] ), .B1(new_n15239_), .B2(new_n15236_), .ZN(new_n15244_));
  INV_X1     g15052(.I(new_n14939_), .ZN(new_n15245_));
  OAI21_X1   g15053(.A1(new_n15244_), .A2(new_n10614_), .B(new_n15245_), .ZN(new_n15246_));
  NAND2_X1   g15054(.A1(new_n15246_), .A2(new_n15243_), .ZN(new_n15247_));
  OAI22_X1   g15055(.A1(new_n15244_), .A2(new_n10614_), .B1(new_n15242_), .B2(new_n15240_), .ZN(new_n15248_));
  AOI21_X1   g15056(.A1(new_n15248_), .A2(\asqrt[24] ), .B(new_n14945_), .ZN(new_n15249_));
  NOR2_X1    g15057(.A1(new_n15249_), .A2(new_n15247_), .ZN(new_n15250_));
  AOI22_X1   g15058(.A1(new_n15248_), .A2(\asqrt[24] ), .B1(new_n15246_), .B2(new_n15243_), .ZN(new_n15251_));
  INV_X1     g15059(.I(new_n14953_), .ZN(new_n15252_));
  OAI21_X1   g15060(.A1(new_n15251_), .A2(new_n9672_), .B(new_n15252_), .ZN(new_n15253_));
  NAND2_X1   g15061(.A1(new_n15253_), .A2(new_n15250_), .ZN(new_n15254_));
  OAI22_X1   g15062(.A1(new_n15251_), .A2(new_n9672_), .B1(new_n15249_), .B2(new_n15247_), .ZN(new_n15255_));
  AOI21_X1   g15063(.A1(new_n15255_), .A2(\asqrt[26] ), .B(new_n14960_), .ZN(new_n15256_));
  NOR2_X1    g15064(.A1(new_n15256_), .A2(new_n15254_), .ZN(new_n15257_));
  AOI22_X1   g15065(.A1(new_n15255_), .A2(\asqrt[26] ), .B1(new_n15253_), .B2(new_n15250_), .ZN(new_n15258_));
  INV_X1     g15066(.I(new_n14968_), .ZN(new_n15259_));
  OAI21_X1   g15067(.A1(new_n15258_), .A2(new_n8763_), .B(new_n15259_), .ZN(new_n15260_));
  NAND2_X1   g15068(.A1(new_n15260_), .A2(new_n15257_), .ZN(new_n15261_));
  OAI22_X1   g15069(.A1(new_n15258_), .A2(new_n8763_), .B1(new_n15256_), .B2(new_n15254_), .ZN(new_n15262_));
  AOI21_X1   g15070(.A1(new_n15262_), .A2(\asqrt[28] ), .B(new_n14975_), .ZN(new_n15263_));
  NOR2_X1    g15071(.A1(new_n15263_), .A2(new_n15261_), .ZN(new_n15264_));
  AOI22_X1   g15072(.A1(new_n15262_), .A2(\asqrt[28] ), .B1(new_n15260_), .B2(new_n15257_), .ZN(new_n15265_));
  INV_X1     g15073(.I(new_n14983_), .ZN(new_n15266_));
  OAI21_X1   g15074(.A1(new_n15265_), .A2(new_n7931_), .B(new_n15266_), .ZN(new_n15267_));
  NAND2_X1   g15075(.A1(new_n15267_), .A2(new_n15264_), .ZN(new_n15268_));
  OAI22_X1   g15076(.A1(new_n15265_), .A2(new_n7931_), .B1(new_n15263_), .B2(new_n15261_), .ZN(new_n15269_));
  AOI21_X1   g15077(.A1(new_n15269_), .A2(\asqrt[30] ), .B(new_n14990_), .ZN(new_n15270_));
  NOR2_X1    g15078(.A1(new_n15270_), .A2(new_n15268_), .ZN(new_n15271_));
  AOI22_X1   g15079(.A1(new_n15269_), .A2(\asqrt[30] ), .B1(new_n15267_), .B2(new_n15264_), .ZN(new_n15272_));
  INV_X1     g15080(.I(new_n14998_), .ZN(new_n15273_));
  OAI21_X1   g15081(.A1(new_n15272_), .A2(new_n7110_), .B(new_n15273_), .ZN(new_n15274_));
  NAND2_X1   g15082(.A1(new_n15274_), .A2(new_n15271_), .ZN(new_n15275_));
  OAI22_X1   g15083(.A1(new_n15272_), .A2(new_n7110_), .B1(new_n15270_), .B2(new_n15268_), .ZN(new_n15276_));
  AOI21_X1   g15084(.A1(new_n15276_), .A2(\asqrt[32] ), .B(new_n15005_), .ZN(new_n15277_));
  NOR2_X1    g15085(.A1(new_n15277_), .A2(new_n15275_), .ZN(new_n15278_));
  AOI22_X1   g15086(.A1(new_n15276_), .A2(\asqrt[32] ), .B1(new_n15274_), .B2(new_n15271_), .ZN(new_n15279_));
  INV_X1     g15087(.I(new_n15013_), .ZN(new_n15280_));
  OAI21_X1   g15088(.A1(new_n15279_), .A2(new_n6365_), .B(new_n15280_), .ZN(new_n15281_));
  NAND2_X1   g15089(.A1(new_n15281_), .A2(new_n15278_), .ZN(new_n15282_));
  OAI22_X1   g15090(.A1(new_n15279_), .A2(new_n6365_), .B1(new_n15277_), .B2(new_n15275_), .ZN(new_n15283_));
  AOI21_X1   g15091(.A1(new_n15283_), .A2(\asqrt[34] ), .B(new_n15020_), .ZN(new_n15284_));
  NOR2_X1    g15092(.A1(new_n15284_), .A2(new_n15282_), .ZN(new_n15285_));
  AOI22_X1   g15093(.A1(new_n15283_), .A2(\asqrt[34] ), .B1(new_n15281_), .B2(new_n15278_), .ZN(new_n15286_));
  INV_X1     g15094(.I(new_n15028_), .ZN(new_n15287_));
  OAI21_X1   g15095(.A1(new_n15286_), .A2(new_n5626_), .B(new_n15287_), .ZN(new_n15288_));
  NAND2_X1   g15096(.A1(new_n15288_), .A2(new_n15285_), .ZN(new_n15289_));
  OAI22_X1   g15097(.A1(new_n15286_), .A2(new_n5626_), .B1(new_n15284_), .B2(new_n15282_), .ZN(new_n15290_));
  AOI21_X1   g15098(.A1(new_n15290_), .A2(\asqrt[36] ), .B(new_n15035_), .ZN(new_n15291_));
  NOR2_X1    g15099(.A1(new_n15291_), .A2(new_n15289_), .ZN(new_n15292_));
  AOI22_X1   g15100(.A1(new_n15290_), .A2(\asqrt[36] ), .B1(new_n15288_), .B2(new_n15285_), .ZN(new_n15293_));
  INV_X1     g15101(.I(new_n15043_), .ZN(new_n15294_));
  OAI21_X1   g15102(.A1(new_n15293_), .A2(new_n4973_), .B(new_n15294_), .ZN(new_n15295_));
  NAND2_X1   g15103(.A1(new_n15295_), .A2(new_n15292_), .ZN(new_n15296_));
  OAI22_X1   g15104(.A1(new_n15293_), .A2(new_n4973_), .B1(new_n15291_), .B2(new_n15289_), .ZN(new_n15297_));
  AOI21_X1   g15105(.A1(new_n15297_), .A2(\asqrt[38] ), .B(new_n15050_), .ZN(new_n15298_));
  NOR2_X1    g15106(.A1(new_n15298_), .A2(new_n15296_), .ZN(new_n15299_));
  AOI22_X1   g15107(.A1(new_n15297_), .A2(\asqrt[38] ), .B1(new_n15295_), .B2(new_n15292_), .ZN(new_n15300_));
  INV_X1     g15108(.I(new_n15058_), .ZN(new_n15301_));
  OAI21_X1   g15109(.A1(new_n15300_), .A2(new_n4330_), .B(new_n15301_), .ZN(new_n15302_));
  NAND2_X1   g15110(.A1(new_n15302_), .A2(new_n15299_), .ZN(new_n15303_));
  OAI22_X1   g15111(.A1(new_n15300_), .A2(new_n4330_), .B1(new_n15298_), .B2(new_n15296_), .ZN(new_n15304_));
  AOI21_X1   g15112(.A1(new_n15304_), .A2(\asqrt[40] ), .B(new_n15065_), .ZN(new_n15305_));
  NOR2_X1    g15113(.A1(new_n15305_), .A2(new_n15303_), .ZN(new_n15306_));
  AOI22_X1   g15114(.A1(new_n15304_), .A2(\asqrt[40] ), .B1(new_n15302_), .B2(new_n15299_), .ZN(new_n15307_));
  INV_X1     g15115(.I(new_n15073_), .ZN(new_n15308_));
  OAI21_X1   g15116(.A1(new_n15307_), .A2(new_n3760_), .B(new_n15308_), .ZN(new_n15309_));
  NAND2_X1   g15117(.A1(new_n15309_), .A2(new_n15306_), .ZN(new_n15310_));
  OAI22_X1   g15118(.A1(new_n15307_), .A2(new_n3760_), .B1(new_n15305_), .B2(new_n15303_), .ZN(new_n15311_));
  AOI21_X1   g15119(.A1(new_n15311_), .A2(\asqrt[42] ), .B(new_n15080_), .ZN(new_n15312_));
  NOR2_X1    g15120(.A1(new_n15312_), .A2(new_n15310_), .ZN(new_n15313_));
  AOI22_X1   g15121(.A1(new_n15311_), .A2(\asqrt[42] ), .B1(new_n15309_), .B2(new_n15306_), .ZN(new_n15314_));
  INV_X1     g15122(.I(new_n15088_), .ZN(new_n15315_));
  OAI21_X1   g15123(.A1(new_n15314_), .A2(new_n3208_), .B(new_n15315_), .ZN(new_n15316_));
  NAND2_X1   g15124(.A1(new_n15316_), .A2(new_n15313_), .ZN(new_n15317_));
  OAI22_X1   g15125(.A1(new_n15314_), .A2(new_n3208_), .B1(new_n15312_), .B2(new_n15310_), .ZN(new_n15318_));
  AOI21_X1   g15126(.A1(new_n15318_), .A2(\asqrt[44] ), .B(new_n15095_), .ZN(new_n15319_));
  NOR2_X1    g15127(.A1(new_n15319_), .A2(new_n15317_), .ZN(new_n15320_));
  AOI22_X1   g15128(.A1(new_n15318_), .A2(\asqrt[44] ), .B1(new_n15316_), .B2(new_n15313_), .ZN(new_n15321_));
  INV_X1     g15129(.I(new_n15103_), .ZN(new_n15322_));
  OAI21_X1   g15130(.A1(new_n15321_), .A2(new_n2728_), .B(new_n15322_), .ZN(new_n15323_));
  NAND2_X1   g15131(.A1(new_n15323_), .A2(new_n15320_), .ZN(new_n15324_));
  OAI22_X1   g15132(.A1(new_n15321_), .A2(new_n2728_), .B1(new_n15319_), .B2(new_n15317_), .ZN(new_n15325_));
  AOI21_X1   g15133(.A1(new_n15325_), .A2(\asqrt[46] ), .B(new_n15110_), .ZN(new_n15326_));
  NOR2_X1    g15134(.A1(new_n15326_), .A2(new_n15324_), .ZN(new_n15327_));
  AOI22_X1   g15135(.A1(new_n15325_), .A2(\asqrt[46] ), .B1(new_n15323_), .B2(new_n15320_), .ZN(new_n15328_));
  INV_X1     g15136(.I(new_n15118_), .ZN(new_n15329_));
  OAI21_X1   g15137(.A1(new_n15328_), .A2(new_n2253_), .B(new_n15329_), .ZN(new_n15330_));
  NAND2_X1   g15138(.A1(new_n15330_), .A2(new_n15327_), .ZN(new_n15331_));
  OAI22_X1   g15139(.A1(new_n15328_), .A2(new_n2253_), .B1(new_n15326_), .B2(new_n15324_), .ZN(new_n15332_));
  AOI21_X1   g15140(.A1(new_n15332_), .A2(\asqrt[48] ), .B(new_n15125_), .ZN(new_n15333_));
  NOR2_X1    g15141(.A1(new_n15333_), .A2(new_n15331_), .ZN(new_n15334_));
  AOI22_X1   g15142(.A1(new_n15332_), .A2(\asqrt[48] ), .B1(new_n15330_), .B2(new_n15327_), .ZN(new_n15335_));
  INV_X1     g15143(.I(new_n15133_), .ZN(new_n15336_));
  OAI21_X1   g15144(.A1(new_n15335_), .A2(new_n1854_), .B(new_n15336_), .ZN(new_n15337_));
  NAND2_X1   g15145(.A1(new_n15337_), .A2(new_n15334_), .ZN(new_n15338_));
  OAI22_X1   g15146(.A1(new_n15335_), .A2(new_n1854_), .B1(new_n15333_), .B2(new_n15331_), .ZN(new_n15339_));
  AOI21_X1   g15147(.A1(new_n15339_), .A2(\asqrt[50] ), .B(new_n15140_), .ZN(new_n15340_));
  NOR2_X1    g15148(.A1(new_n15340_), .A2(new_n15338_), .ZN(new_n15341_));
  AOI22_X1   g15149(.A1(new_n15339_), .A2(\asqrt[50] ), .B1(new_n15337_), .B2(new_n15334_), .ZN(new_n15342_));
  INV_X1     g15150(.I(new_n15148_), .ZN(new_n15343_));
  OAI21_X1   g15151(.A1(new_n15342_), .A2(new_n1436_), .B(new_n15343_), .ZN(new_n15344_));
  NAND2_X1   g15152(.A1(new_n15344_), .A2(new_n15341_), .ZN(new_n15345_));
  OAI22_X1   g15153(.A1(new_n15342_), .A2(new_n1436_), .B1(new_n15340_), .B2(new_n15338_), .ZN(new_n15346_));
  AOI21_X1   g15154(.A1(new_n15346_), .A2(\asqrt[52] ), .B(new_n15154_), .ZN(new_n15347_));
  NOR2_X1    g15155(.A1(new_n15347_), .A2(new_n15345_), .ZN(new_n15348_));
  AOI22_X1   g15156(.A1(new_n15346_), .A2(\asqrt[52] ), .B1(new_n15344_), .B2(new_n15341_), .ZN(new_n15349_));
  INV_X1     g15157(.I(new_n15161_), .ZN(new_n15350_));
  OAI21_X1   g15158(.A1(new_n15349_), .A2(new_n1096_), .B(new_n15350_), .ZN(new_n15351_));
  NAND2_X1   g15159(.A1(new_n15351_), .A2(new_n15348_), .ZN(new_n15352_));
  OAI22_X1   g15160(.A1(new_n15349_), .A2(new_n1096_), .B1(new_n15347_), .B2(new_n15345_), .ZN(new_n15353_));
  AOI21_X1   g15161(.A1(new_n15353_), .A2(\asqrt[54] ), .B(new_n15167_), .ZN(new_n15354_));
  NOR2_X1    g15162(.A1(new_n15354_), .A2(new_n15352_), .ZN(new_n15355_));
  AOI22_X1   g15163(.A1(new_n15353_), .A2(\asqrt[54] ), .B1(new_n15351_), .B2(new_n15348_), .ZN(new_n15356_));
  INV_X1     g15164(.I(new_n15174_), .ZN(new_n15357_));
  OAI21_X1   g15165(.A1(new_n15356_), .A2(new_n825_), .B(new_n15357_), .ZN(new_n15358_));
  NAND2_X1   g15166(.A1(new_n15358_), .A2(new_n15355_), .ZN(new_n15359_));
  OAI22_X1   g15167(.A1(new_n15356_), .A2(new_n825_), .B1(new_n15354_), .B2(new_n15352_), .ZN(new_n15360_));
  AOI21_X1   g15168(.A1(new_n15360_), .A2(\asqrt[56] ), .B(new_n15180_), .ZN(new_n15361_));
  NOR2_X1    g15169(.A1(new_n15361_), .A2(new_n15359_), .ZN(new_n15362_));
  AOI22_X1   g15170(.A1(new_n15360_), .A2(\asqrt[56] ), .B1(new_n15358_), .B2(new_n15355_), .ZN(new_n15363_));
  INV_X1     g15171(.I(new_n15187_), .ZN(new_n15364_));
  OAI21_X1   g15172(.A1(new_n15363_), .A2(new_n587_), .B(new_n15364_), .ZN(new_n15365_));
  NAND2_X1   g15173(.A1(new_n15365_), .A2(new_n15362_), .ZN(new_n15366_));
  OAI22_X1   g15174(.A1(new_n15363_), .A2(new_n587_), .B1(new_n15361_), .B2(new_n15359_), .ZN(new_n15367_));
  AOI21_X1   g15175(.A1(new_n15367_), .A2(\asqrt[58] ), .B(new_n15193_), .ZN(new_n15368_));
  NOR2_X1    g15176(.A1(new_n15368_), .A2(new_n15366_), .ZN(new_n15369_));
  AOI22_X1   g15177(.A1(new_n15367_), .A2(\asqrt[58] ), .B1(new_n15365_), .B2(new_n15362_), .ZN(new_n15370_));
  INV_X1     g15178(.I(new_n15200_), .ZN(new_n15371_));
  OAI21_X1   g15179(.A1(new_n15370_), .A2(new_n376_), .B(new_n15371_), .ZN(new_n15372_));
  NAND2_X1   g15180(.A1(new_n15372_), .A2(new_n15369_), .ZN(new_n15373_));
  OAI22_X1   g15181(.A1(new_n15370_), .A2(new_n376_), .B1(new_n15368_), .B2(new_n15366_), .ZN(new_n15374_));
  AOI22_X1   g15182(.A1(new_n15374_), .A2(\asqrt[60] ), .B1(new_n15372_), .B2(new_n15369_), .ZN(new_n15375_));
  AOI21_X1   g15183(.A1(new_n15374_), .A2(\asqrt[60] ), .B(new_n15207_), .ZN(new_n15376_));
  OAI22_X1   g15184(.A1(new_n15375_), .A2(new_n229_), .B1(new_n15376_), .B2(new_n15373_), .ZN(new_n15377_));
  NOR2_X1    g15185(.A1(new_n15377_), .A2(\asqrt[62] ), .ZN(new_n15378_));
  NAND3_X1   g15186(.A1(new_n14865_), .A2(new_n14643_), .A3(new_n14833_), .ZN(new_n15379_));
  NOR2_X1    g15187(.A1(new_n14874_), .A2(new_n196_), .ZN(new_n15380_));
  INV_X1     g15188(.I(new_n14859_), .ZN(new_n15381_));
  NAND3_X1   g15189(.A1(\asqrt[15] ), .A2(new_n15380_), .A3(new_n15381_), .ZN(new_n15382_));
  OAI21_X1   g15190(.A1(new_n14830_), .A2(\asqrt[62] ), .B(new_n14645_), .ZN(new_n15383_));
  OAI21_X1   g15191(.A1(\asqrt[15] ), .A2(new_n15383_), .B(new_n15380_), .ZN(new_n15384_));
  NAND2_X1   g15192(.A1(new_n15384_), .A2(new_n15382_), .ZN(new_n15385_));
  INV_X1     g15193(.I(new_n15385_), .ZN(new_n15386_));
  NOR2_X1    g15194(.A1(new_n14838_), .A2(new_n196_), .ZN(new_n15387_));
  INV_X1     g15195(.I(new_n15387_), .ZN(new_n15388_));
  NAND2_X1   g15196(.A1(new_n15197_), .A2(\asqrt[59] ), .ZN(new_n15389_));
  AOI21_X1   g15197(.A1(new_n15389_), .A2(new_n15196_), .B(new_n275_), .ZN(new_n15390_));
  OAI21_X1   g15198(.A1(new_n15202_), .A2(new_n15390_), .B(\asqrt[61] ), .ZN(new_n15391_));
  NOR2_X1    g15199(.A1(new_n14839_), .A2(\asqrt[62] ), .ZN(new_n15392_));
  INV_X1     g15200(.I(new_n15392_), .ZN(new_n15393_));
  NAND3_X1   g15201(.A1(new_n15209_), .A2(new_n15202_), .A3(new_n15393_), .ZN(new_n15394_));
  OAI21_X1   g15202(.A1(new_n15394_), .A2(new_n15391_), .B(new_n15388_), .ZN(new_n15395_));
  NAND3_X1   g15203(.A1(new_n14871_), .A2(new_n14826_), .A3(new_n14875_), .ZN(new_n15396_));
  AOI21_X1   g15204(.A1(new_n15396_), .A2(new_n14818_), .B(\asqrt[63] ), .ZN(new_n15397_));
  INV_X1     g15205(.I(new_n15397_), .ZN(new_n15398_));
  OAI21_X1   g15206(.A1(new_n15395_), .A2(new_n15398_), .B(new_n15386_), .ZN(new_n15399_));
  NOR4_X1    g15207(.A1(new_n15377_), .A2(\asqrt[62] ), .A3(new_n15385_), .A4(new_n14838_), .ZN(new_n15400_));
  NAND2_X1   g15208(.A1(new_n14853_), .A2(new_n14826_), .ZN(new_n15401_));
  XOR2_X1    g15209(.A1(new_n14853_), .A2(\asqrt[63] ), .Z(new_n15402_));
  AOI21_X1   g15210(.A1(\asqrt[15] ), .A2(new_n15401_), .B(new_n15402_), .ZN(new_n15403_));
  NAND2_X1   g15211(.A1(new_n15400_), .A2(new_n15403_), .ZN(new_n15404_));
  NOR3_X1    g15212(.A1(new_n15404_), .A2(new_n15379_), .A3(new_n15399_), .ZN(\asqrt[14] ));
  NAND4_X1   g15213(.A1(\asqrt[14] ), .A2(new_n14839_), .A3(new_n15211_), .A4(new_n15378_), .ZN(new_n15406_));
  OAI21_X1   g15214(.A1(new_n15377_), .A2(\asqrt[62] ), .B(new_n14838_), .ZN(new_n15407_));
  OAI21_X1   g15215(.A1(\asqrt[14] ), .A2(new_n15407_), .B(new_n15211_), .ZN(new_n15408_));
  NAND2_X1   g15216(.A1(new_n15406_), .A2(new_n15408_), .ZN(new_n15409_));
  INV_X1     g15217(.I(new_n15409_), .ZN(new_n15410_));
  NAND2_X1   g15218(.A1(new_n15367_), .A2(\asqrt[58] ), .ZN(new_n15411_));
  AOI21_X1   g15219(.A1(new_n15411_), .A2(new_n15366_), .B(new_n376_), .ZN(new_n15412_));
  OAI21_X1   g15220(.A1(new_n15369_), .A2(new_n15412_), .B(\asqrt[60] ), .ZN(new_n15413_));
  AOI21_X1   g15221(.A1(new_n15373_), .A2(new_n15413_), .B(new_n229_), .ZN(new_n15414_));
  NOR3_X1    g15222(.A1(new_n15204_), .A2(\asqrt[61] ), .A3(new_n15206_), .ZN(new_n15415_));
  NAND2_X1   g15223(.A1(\asqrt[14] ), .A2(new_n15415_), .ZN(new_n15416_));
  XOR2_X1    g15224(.A1(new_n15416_), .A2(new_n15414_), .Z(new_n15417_));
  NOR2_X1    g15225(.A1(new_n15417_), .A2(new_n196_), .ZN(new_n15418_));
  INV_X1     g15226(.I(new_n15418_), .ZN(new_n15419_));
  INV_X1     g15227(.I(\a[28] ), .ZN(new_n15420_));
  NOR2_X1    g15228(.A1(\a[26] ), .A2(\a[27] ), .ZN(new_n15421_));
  INV_X1     g15229(.I(new_n15421_), .ZN(new_n15422_));
  NOR3_X1    g15230(.A1(new_n14877_), .A2(new_n15420_), .A3(new_n15422_), .ZN(new_n15423_));
  NAND2_X1   g15231(.A1(new_n14883_), .A2(new_n15423_), .ZN(new_n15424_));
  XOR2_X1    g15232(.A1(new_n15424_), .A2(\a[29] ), .Z(new_n15425_));
  INV_X1     g15233(.I(\a[29] ), .ZN(new_n15426_));
  NOR4_X1    g15234(.A1(new_n15404_), .A2(new_n15426_), .A3(new_n15379_), .A4(new_n15399_), .ZN(new_n15427_));
  NOR2_X1    g15235(.A1(new_n15426_), .A2(\a[28] ), .ZN(new_n15428_));
  OAI21_X1   g15236(.A1(new_n15427_), .A2(new_n15428_), .B(new_n15425_), .ZN(new_n15429_));
  INV_X1     g15237(.I(new_n15425_), .ZN(new_n15430_));
  INV_X1     g15238(.I(new_n15379_), .ZN(new_n15431_));
  NOR3_X1    g15239(.A1(new_n15376_), .A2(new_n15373_), .A3(new_n15392_), .ZN(new_n15432_));
  AOI21_X1   g15240(.A1(new_n15432_), .A2(new_n15414_), .B(new_n15387_), .ZN(new_n15433_));
  AOI21_X1   g15241(.A1(new_n15433_), .A2(new_n15397_), .B(new_n15385_), .ZN(new_n15434_));
  NAND4_X1   g15242(.A1(new_n15210_), .A2(new_n196_), .A3(new_n15386_), .A4(new_n14839_), .ZN(new_n15435_));
  INV_X1     g15243(.I(new_n15403_), .ZN(new_n15436_));
  NOR2_X1    g15244(.A1(new_n15435_), .A2(new_n15436_), .ZN(new_n15437_));
  NAND4_X1   g15245(.A1(new_n15437_), .A2(\a[29] ), .A3(new_n15434_), .A4(new_n15431_), .ZN(new_n15438_));
  NAND3_X1   g15246(.A1(new_n15438_), .A2(\a[28] ), .A3(new_n15430_), .ZN(new_n15439_));
  NAND2_X1   g15247(.A1(new_n15429_), .A2(new_n15439_), .ZN(new_n15440_));
  NOR2_X1    g15248(.A1(new_n15404_), .A2(new_n15399_), .ZN(new_n15441_));
  NOR4_X1    g15249(.A1(new_n14832_), .A2(new_n14826_), .A3(new_n14873_), .A4(new_n14833_), .ZN(new_n15442_));
  NAND2_X1   g15250(.A1(\asqrt[15] ), .A2(\a[28] ), .ZN(new_n15443_));
  XOR2_X1    g15251(.A1(new_n15443_), .A2(new_n15442_), .Z(new_n15444_));
  NOR2_X1    g15252(.A1(new_n15444_), .A2(new_n15422_), .ZN(new_n15445_));
  INV_X1     g15253(.I(new_n15445_), .ZN(new_n15446_));
  NAND3_X1   g15254(.A1(new_n15437_), .A2(new_n15431_), .A3(new_n15434_), .ZN(new_n15447_));
  NOR2_X1    g15255(.A1(new_n15431_), .A2(new_n15403_), .ZN(new_n15448_));
  NAND2_X1   g15256(.A1(new_n15448_), .A2(\asqrt[15] ), .ZN(new_n15449_));
  INV_X1     g15257(.I(new_n15449_), .ZN(new_n15450_));
  NAND3_X1   g15258(.A1(new_n15399_), .A2(new_n15435_), .A3(new_n15450_), .ZN(new_n15451_));
  NAND2_X1   g15259(.A1(new_n15451_), .A2(new_n14840_), .ZN(new_n15452_));
  NAND3_X1   g15260(.A1(new_n15452_), .A2(new_n14841_), .A3(new_n15447_), .ZN(new_n15453_));
  NOR3_X1    g15261(.A1(new_n15434_), .A2(new_n15400_), .A3(new_n15449_), .ZN(new_n15454_));
  OAI21_X1   g15262(.A1(new_n15454_), .A2(\a[30] ), .B(new_n14841_), .ZN(new_n15455_));
  NAND2_X1   g15263(.A1(new_n15455_), .A2(\asqrt[14] ), .ZN(new_n15456_));
  NAND4_X1   g15264(.A1(new_n15456_), .A2(new_n14273_), .A3(new_n15453_), .A4(new_n15446_), .ZN(new_n15457_));
  NAND2_X1   g15265(.A1(new_n15457_), .A2(new_n15440_), .ZN(new_n15458_));
  NAND3_X1   g15266(.A1(new_n15429_), .A2(new_n15439_), .A3(new_n15446_), .ZN(new_n15459_));
  AOI21_X1   g15267(.A1(\asqrt[15] ), .A2(new_n14840_), .B(\a[31] ), .ZN(new_n15460_));
  NOR2_X1    g15268(.A1(new_n14862_), .A2(\a[30] ), .ZN(new_n15461_));
  AOI21_X1   g15269(.A1(\asqrt[15] ), .A2(\a[30] ), .B(new_n14844_), .ZN(new_n15462_));
  OAI21_X1   g15270(.A1(new_n15461_), .A2(new_n15460_), .B(new_n15462_), .ZN(new_n15463_));
  INV_X1     g15271(.I(new_n15463_), .ZN(new_n15464_));
  NAND3_X1   g15272(.A1(\asqrt[14] ), .A2(new_n14870_), .A3(new_n15464_), .ZN(new_n15465_));
  OAI21_X1   g15273(.A1(new_n15447_), .A2(new_n15463_), .B(new_n14869_), .ZN(new_n15466_));
  NAND3_X1   g15274(.A1(new_n15465_), .A2(new_n15466_), .A3(new_n13760_), .ZN(new_n15467_));
  AOI21_X1   g15275(.A1(new_n15459_), .A2(\asqrt[16] ), .B(new_n15467_), .ZN(new_n15468_));
  NOR2_X1    g15276(.A1(new_n15458_), .A2(new_n15468_), .ZN(new_n15469_));
  AOI22_X1   g15277(.A1(new_n15457_), .A2(new_n15440_), .B1(\asqrt[16] ), .B2(new_n15459_), .ZN(new_n15470_));
  NOR2_X1    g15278(.A1(new_n15217_), .A2(new_n15216_), .ZN(new_n15471_));
  NOR4_X1    g15279(.A1(new_n15447_), .A2(\asqrt[17] ), .A3(new_n15471_), .A4(new_n14889_), .ZN(new_n15472_));
  AOI21_X1   g15280(.A1(new_n15215_), .A2(new_n14870_), .B(new_n13760_), .ZN(new_n15473_));
  NOR2_X1    g15281(.A1(new_n15472_), .A2(new_n15473_), .ZN(new_n15474_));
  NAND2_X1   g15282(.A1(new_n15474_), .A2(new_n13192_), .ZN(new_n15475_));
  INV_X1     g15283(.I(new_n15475_), .ZN(new_n15476_));
  OAI21_X1   g15284(.A1(new_n15470_), .A2(new_n13760_), .B(new_n15476_), .ZN(new_n15477_));
  NAND2_X1   g15285(.A1(new_n15459_), .A2(\asqrt[16] ), .ZN(new_n15478_));
  AOI21_X1   g15286(.A1(new_n15458_), .A2(new_n15478_), .B(new_n13760_), .ZN(new_n15479_));
  OAI21_X1   g15287(.A1(new_n15479_), .A2(new_n15469_), .B(\asqrt[18] ), .ZN(new_n15480_));
  NOR2_X1    g15288(.A1(new_n14901_), .A2(new_n13192_), .ZN(new_n15481_));
  NAND2_X1   g15289(.A1(new_n14895_), .A2(new_n14897_), .ZN(new_n15482_));
  NAND4_X1   g15290(.A1(\asqrt[14] ), .A2(new_n13192_), .A3(new_n15482_), .A4(new_n14901_), .ZN(new_n15483_));
  XOR2_X1    g15291(.A1(new_n15483_), .A2(new_n15481_), .Z(new_n15484_));
  NAND2_X1   g15292(.A1(new_n15484_), .A2(new_n12657_), .ZN(new_n15485_));
  INV_X1     g15293(.I(new_n15485_), .ZN(new_n15486_));
  NAND2_X1   g15294(.A1(new_n15480_), .A2(new_n15486_), .ZN(new_n15487_));
  NAND3_X1   g15295(.A1(new_n15487_), .A2(new_n15469_), .A3(new_n15477_), .ZN(new_n15488_));
  INV_X1     g15296(.I(new_n15428_), .ZN(new_n15489_));
  AOI21_X1   g15297(.A1(new_n15438_), .A2(new_n15489_), .B(new_n15430_), .ZN(new_n15490_));
  NOR3_X1    g15298(.A1(new_n15427_), .A2(new_n15420_), .A3(new_n15425_), .ZN(new_n15491_));
  NOR2_X1    g15299(.A1(new_n15491_), .A2(new_n15490_), .ZN(new_n15492_));
  NOR2_X1    g15300(.A1(new_n15455_), .A2(\asqrt[14] ), .ZN(new_n15493_));
  AOI21_X1   g15301(.A1(new_n15452_), .A2(new_n14841_), .B(new_n15447_), .ZN(new_n15494_));
  NOR4_X1    g15302(.A1(new_n15493_), .A2(\asqrt[16] ), .A3(new_n15494_), .A4(new_n15445_), .ZN(new_n15495_));
  NOR2_X1    g15303(.A1(new_n15495_), .A2(new_n15492_), .ZN(new_n15496_));
  NOR3_X1    g15304(.A1(new_n15491_), .A2(new_n15490_), .A3(new_n15445_), .ZN(new_n15497_));
  NOR3_X1    g15305(.A1(new_n15447_), .A2(new_n14869_), .A3(new_n15463_), .ZN(new_n15498_));
  AOI21_X1   g15306(.A1(\asqrt[14] ), .A2(new_n15464_), .B(new_n14870_), .ZN(new_n15499_));
  NOR3_X1    g15307(.A1(new_n15499_), .A2(new_n15498_), .A3(\asqrt[17] ), .ZN(new_n15500_));
  OAI21_X1   g15308(.A1(new_n15497_), .A2(new_n14273_), .B(new_n15500_), .ZN(new_n15501_));
  NAND2_X1   g15309(.A1(new_n15496_), .A2(new_n15501_), .ZN(new_n15502_));
  OAI22_X1   g15310(.A1(new_n15495_), .A2(new_n15492_), .B1(new_n14273_), .B2(new_n15497_), .ZN(new_n15503_));
  AOI21_X1   g15311(.A1(new_n15503_), .A2(\asqrt[17] ), .B(new_n15475_), .ZN(new_n15504_));
  AOI22_X1   g15312(.A1(new_n15503_), .A2(\asqrt[17] ), .B1(new_n15496_), .B2(new_n15501_), .ZN(new_n15505_));
  OAI22_X1   g15313(.A1(new_n15505_), .A2(new_n13192_), .B1(new_n15504_), .B2(new_n15502_), .ZN(new_n15506_));
  NAND2_X1   g15314(.A1(new_n14908_), .A2(\asqrt[19] ), .ZN(new_n15507_));
  NOR2_X1    g15315(.A1(new_n14903_), .A2(new_n14904_), .ZN(new_n15508_));
  NOR4_X1    g15316(.A1(new_n15447_), .A2(\asqrt[19] ), .A3(new_n15508_), .A4(new_n14908_), .ZN(new_n15509_));
  XOR2_X1    g15317(.A1(new_n15509_), .A2(new_n15507_), .Z(new_n15510_));
  NAND2_X1   g15318(.A1(new_n15510_), .A2(new_n12101_), .ZN(new_n15511_));
  AOI21_X1   g15319(.A1(new_n15506_), .A2(\asqrt[19] ), .B(new_n15511_), .ZN(new_n15512_));
  NOR2_X1    g15320(.A1(new_n15512_), .A2(new_n15488_), .ZN(new_n15513_));
  OAI21_X1   g15321(.A1(new_n15479_), .A2(new_n15475_), .B(new_n15469_), .ZN(new_n15514_));
  AOI21_X1   g15322(.A1(new_n15480_), .A2(new_n15486_), .B(new_n15514_), .ZN(new_n15515_));
  AOI21_X1   g15323(.A1(new_n15514_), .A2(new_n15480_), .B(new_n12657_), .ZN(new_n15516_));
  OAI21_X1   g15324(.A1(new_n15515_), .A2(new_n15516_), .B(\asqrt[20] ), .ZN(new_n15517_));
  NOR4_X1    g15325(.A1(new_n15447_), .A2(\asqrt[20] ), .A3(new_n14911_), .A4(new_n15234_), .ZN(new_n15518_));
  AOI21_X1   g15326(.A1(new_n15507_), .A2(new_n14907_), .B(new_n12101_), .ZN(new_n15519_));
  NOR2_X1    g15327(.A1(new_n15518_), .A2(new_n15519_), .ZN(new_n15520_));
  NAND2_X1   g15328(.A1(new_n15520_), .A2(new_n11631_), .ZN(new_n15521_));
  INV_X1     g15329(.I(new_n15521_), .ZN(new_n15522_));
  NAND2_X1   g15330(.A1(new_n15517_), .A2(new_n15522_), .ZN(new_n15523_));
  NAND2_X1   g15331(.A1(new_n15523_), .A2(new_n15513_), .ZN(new_n15524_));
  NOR2_X1    g15332(.A1(new_n15515_), .A2(new_n15516_), .ZN(new_n15525_));
  OAI22_X1   g15333(.A1(new_n15525_), .A2(new_n12101_), .B1(new_n15512_), .B2(new_n15488_), .ZN(new_n15526_));
  NAND2_X1   g15334(.A1(new_n14923_), .A2(\asqrt[21] ), .ZN(new_n15527_));
  NOR4_X1    g15335(.A1(new_n15447_), .A2(\asqrt[21] ), .A3(new_n14918_), .A4(new_n14923_), .ZN(new_n15528_));
  XOR2_X1    g15336(.A1(new_n15528_), .A2(new_n15527_), .Z(new_n15529_));
  NAND2_X1   g15337(.A1(new_n15529_), .A2(new_n11105_), .ZN(new_n15530_));
  AOI21_X1   g15338(.A1(new_n15526_), .A2(\asqrt[21] ), .B(new_n15530_), .ZN(new_n15531_));
  NOR2_X1    g15339(.A1(new_n15531_), .A2(new_n15524_), .ZN(new_n15532_));
  OAI21_X1   g15340(.A1(new_n15516_), .A2(new_n15511_), .B(new_n15515_), .ZN(new_n15533_));
  AOI21_X1   g15341(.A1(new_n15517_), .A2(new_n15522_), .B(new_n15533_), .ZN(new_n15534_));
  AOI21_X1   g15342(.A1(new_n15533_), .A2(new_n15517_), .B(new_n11631_), .ZN(new_n15535_));
  OAI21_X1   g15343(.A1(new_n15534_), .A2(new_n15535_), .B(\asqrt[22] ), .ZN(new_n15536_));
  NOR4_X1    g15344(.A1(new_n15447_), .A2(\asqrt[22] ), .A3(new_n14925_), .A4(new_n15241_), .ZN(new_n15537_));
  AOI21_X1   g15345(.A1(new_n15527_), .A2(new_n14922_), .B(new_n11105_), .ZN(new_n15538_));
  NOR2_X1    g15346(.A1(new_n15537_), .A2(new_n15538_), .ZN(new_n15539_));
  NAND2_X1   g15347(.A1(new_n15539_), .A2(new_n10614_), .ZN(new_n15540_));
  INV_X1     g15348(.I(new_n15540_), .ZN(new_n15541_));
  NAND2_X1   g15349(.A1(new_n15536_), .A2(new_n15541_), .ZN(new_n15542_));
  NAND2_X1   g15350(.A1(new_n15542_), .A2(new_n15532_), .ZN(new_n15543_));
  AOI22_X1   g15351(.A1(new_n15526_), .A2(\asqrt[21] ), .B1(new_n15523_), .B2(new_n15513_), .ZN(new_n15544_));
  OAI22_X1   g15352(.A1(new_n15544_), .A2(new_n11105_), .B1(new_n15531_), .B2(new_n15524_), .ZN(new_n15545_));
  NAND2_X1   g15353(.A1(new_n14936_), .A2(\asqrt[23] ), .ZN(new_n15546_));
  NOR4_X1    g15354(.A1(new_n15447_), .A2(\asqrt[23] ), .A3(new_n14931_), .A4(new_n14936_), .ZN(new_n15547_));
  XOR2_X1    g15355(.A1(new_n15547_), .A2(new_n15546_), .Z(new_n15548_));
  NAND2_X1   g15356(.A1(new_n15548_), .A2(new_n10104_), .ZN(new_n15549_));
  AOI21_X1   g15357(.A1(new_n15545_), .A2(\asqrt[23] ), .B(new_n15549_), .ZN(new_n15550_));
  NOR2_X1    g15358(.A1(new_n15550_), .A2(new_n15543_), .ZN(new_n15551_));
  AOI22_X1   g15359(.A1(new_n15545_), .A2(\asqrt[23] ), .B1(new_n15542_), .B2(new_n15532_), .ZN(new_n15552_));
  NOR4_X1    g15360(.A1(new_n15447_), .A2(\asqrt[24] ), .A3(new_n14938_), .A4(new_n15248_), .ZN(new_n15553_));
  AOI21_X1   g15361(.A1(new_n15546_), .A2(new_n14935_), .B(new_n10104_), .ZN(new_n15554_));
  NOR2_X1    g15362(.A1(new_n15553_), .A2(new_n15554_), .ZN(new_n15555_));
  NAND2_X1   g15363(.A1(new_n15555_), .A2(new_n9672_), .ZN(new_n15556_));
  INV_X1     g15364(.I(new_n15556_), .ZN(new_n15557_));
  OAI21_X1   g15365(.A1(new_n15552_), .A2(new_n10104_), .B(new_n15557_), .ZN(new_n15558_));
  NAND2_X1   g15366(.A1(new_n15558_), .A2(new_n15551_), .ZN(new_n15559_));
  OAI22_X1   g15367(.A1(new_n15552_), .A2(new_n10104_), .B1(new_n15550_), .B2(new_n15543_), .ZN(new_n15560_));
  NAND2_X1   g15368(.A1(new_n14949_), .A2(\asqrt[25] ), .ZN(new_n15561_));
  NOR4_X1    g15369(.A1(new_n15447_), .A2(\asqrt[25] ), .A3(new_n14944_), .A4(new_n14949_), .ZN(new_n15562_));
  XOR2_X1    g15370(.A1(new_n15562_), .A2(new_n15561_), .Z(new_n15563_));
  NAND2_X1   g15371(.A1(new_n15563_), .A2(new_n9212_), .ZN(new_n15564_));
  AOI21_X1   g15372(.A1(new_n15560_), .A2(\asqrt[25] ), .B(new_n15564_), .ZN(new_n15565_));
  NOR2_X1    g15373(.A1(new_n15565_), .A2(new_n15559_), .ZN(new_n15566_));
  AOI22_X1   g15374(.A1(new_n15560_), .A2(\asqrt[25] ), .B1(new_n15558_), .B2(new_n15551_), .ZN(new_n15567_));
  NAND2_X1   g15375(.A1(new_n15255_), .A2(\asqrt[26] ), .ZN(new_n15568_));
  NOR4_X1    g15376(.A1(new_n15447_), .A2(\asqrt[26] ), .A3(new_n14952_), .A4(new_n15255_), .ZN(new_n15569_));
  XOR2_X1    g15377(.A1(new_n15569_), .A2(new_n15568_), .Z(new_n15570_));
  NAND2_X1   g15378(.A1(new_n15570_), .A2(new_n8763_), .ZN(new_n15571_));
  INV_X1     g15379(.I(new_n15571_), .ZN(new_n15572_));
  OAI21_X1   g15380(.A1(new_n15567_), .A2(new_n9212_), .B(new_n15572_), .ZN(new_n15573_));
  NAND2_X1   g15381(.A1(new_n15573_), .A2(new_n15566_), .ZN(new_n15574_));
  OAI22_X1   g15382(.A1(new_n15567_), .A2(new_n9212_), .B1(new_n15565_), .B2(new_n15559_), .ZN(new_n15575_));
  NOR4_X1    g15383(.A1(new_n15447_), .A2(\asqrt[27] ), .A3(new_n14959_), .A4(new_n14964_), .ZN(new_n15576_));
  AOI21_X1   g15384(.A1(new_n15568_), .A2(new_n15254_), .B(new_n8763_), .ZN(new_n15577_));
  NOR2_X1    g15385(.A1(new_n15576_), .A2(new_n15577_), .ZN(new_n15578_));
  NAND2_X1   g15386(.A1(new_n15578_), .A2(new_n8319_), .ZN(new_n15579_));
  AOI21_X1   g15387(.A1(new_n15575_), .A2(\asqrt[27] ), .B(new_n15579_), .ZN(new_n15580_));
  NOR2_X1    g15388(.A1(new_n15580_), .A2(new_n15574_), .ZN(new_n15581_));
  AOI22_X1   g15389(.A1(new_n15575_), .A2(\asqrt[27] ), .B1(new_n15573_), .B2(new_n15566_), .ZN(new_n15582_));
  NAND2_X1   g15390(.A1(new_n15262_), .A2(\asqrt[28] ), .ZN(new_n15583_));
  NOR4_X1    g15391(.A1(new_n15447_), .A2(\asqrt[28] ), .A3(new_n14967_), .A4(new_n15262_), .ZN(new_n15584_));
  XOR2_X1    g15392(.A1(new_n15584_), .A2(new_n15583_), .Z(new_n15585_));
  NAND2_X1   g15393(.A1(new_n15585_), .A2(new_n7931_), .ZN(new_n15586_));
  INV_X1     g15394(.I(new_n15586_), .ZN(new_n15587_));
  OAI21_X1   g15395(.A1(new_n15582_), .A2(new_n8319_), .B(new_n15587_), .ZN(new_n15588_));
  NAND2_X1   g15396(.A1(new_n15588_), .A2(new_n15581_), .ZN(new_n15589_));
  OAI22_X1   g15397(.A1(new_n15582_), .A2(new_n8319_), .B1(new_n15580_), .B2(new_n15574_), .ZN(new_n15590_));
  NOR4_X1    g15398(.A1(new_n15447_), .A2(\asqrt[29] ), .A3(new_n14974_), .A4(new_n14979_), .ZN(new_n15591_));
  AOI21_X1   g15399(.A1(new_n15583_), .A2(new_n15261_), .B(new_n7931_), .ZN(new_n15592_));
  NOR2_X1    g15400(.A1(new_n15591_), .A2(new_n15592_), .ZN(new_n15593_));
  NAND2_X1   g15401(.A1(new_n15593_), .A2(new_n7517_), .ZN(new_n15594_));
  AOI21_X1   g15402(.A1(new_n15590_), .A2(\asqrt[29] ), .B(new_n15594_), .ZN(new_n15595_));
  NOR2_X1    g15403(.A1(new_n15595_), .A2(new_n15589_), .ZN(new_n15596_));
  AOI22_X1   g15404(.A1(new_n15590_), .A2(\asqrt[29] ), .B1(new_n15588_), .B2(new_n15581_), .ZN(new_n15597_));
  NAND2_X1   g15405(.A1(new_n15269_), .A2(\asqrt[30] ), .ZN(new_n15598_));
  NOR4_X1    g15406(.A1(new_n15447_), .A2(\asqrt[30] ), .A3(new_n14982_), .A4(new_n15269_), .ZN(new_n15599_));
  XOR2_X1    g15407(.A1(new_n15599_), .A2(new_n15598_), .Z(new_n15600_));
  NAND2_X1   g15408(.A1(new_n15600_), .A2(new_n7110_), .ZN(new_n15601_));
  INV_X1     g15409(.I(new_n15601_), .ZN(new_n15602_));
  OAI21_X1   g15410(.A1(new_n15597_), .A2(new_n7517_), .B(new_n15602_), .ZN(new_n15603_));
  NAND2_X1   g15411(.A1(new_n15603_), .A2(new_n15596_), .ZN(new_n15604_));
  OAI22_X1   g15412(.A1(new_n15597_), .A2(new_n7517_), .B1(new_n15595_), .B2(new_n15589_), .ZN(new_n15605_));
  NOR4_X1    g15413(.A1(new_n15447_), .A2(\asqrt[31] ), .A3(new_n14989_), .A4(new_n14994_), .ZN(new_n15606_));
  AOI21_X1   g15414(.A1(new_n15598_), .A2(new_n15268_), .B(new_n7110_), .ZN(new_n15607_));
  NOR2_X1    g15415(.A1(new_n15606_), .A2(new_n15607_), .ZN(new_n15608_));
  NAND2_X1   g15416(.A1(new_n15608_), .A2(new_n6708_), .ZN(new_n15609_));
  AOI21_X1   g15417(.A1(new_n15605_), .A2(\asqrt[31] ), .B(new_n15609_), .ZN(new_n15610_));
  NOR2_X1    g15418(.A1(new_n15610_), .A2(new_n15604_), .ZN(new_n15611_));
  AOI22_X1   g15419(.A1(new_n15605_), .A2(\asqrt[31] ), .B1(new_n15603_), .B2(new_n15596_), .ZN(new_n15612_));
  NAND2_X1   g15420(.A1(new_n15276_), .A2(\asqrt[32] ), .ZN(new_n15613_));
  NOR4_X1    g15421(.A1(new_n15447_), .A2(\asqrt[32] ), .A3(new_n14997_), .A4(new_n15276_), .ZN(new_n15614_));
  XOR2_X1    g15422(.A1(new_n15614_), .A2(new_n15613_), .Z(new_n15615_));
  NAND2_X1   g15423(.A1(new_n15615_), .A2(new_n6365_), .ZN(new_n15616_));
  INV_X1     g15424(.I(new_n15616_), .ZN(new_n15617_));
  OAI21_X1   g15425(.A1(new_n15612_), .A2(new_n6708_), .B(new_n15617_), .ZN(new_n15618_));
  NAND2_X1   g15426(.A1(new_n15618_), .A2(new_n15611_), .ZN(new_n15619_));
  OAI22_X1   g15427(.A1(new_n15612_), .A2(new_n6708_), .B1(new_n15610_), .B2(new_n15604_), .ZN(new_n15620_));
  NOR4_X1    g15428(.A1(new_n15447_), .A2(\asqrt[33] ), .A3(new_n15004_), .A4(new_n15009_), .ZN(new_n15621_));
  AOI21_X1   g15429(.A1(new_n15613_), .A2(new_n15275_), .B(new_n6365_), .ZN(new_n15622_));
  NOR2_X1    g15430(.A1(new_n15621_), .A2(new_n15622_), .ZN(new_n15623_));
  NAND2_X1   g15431(.A1(new_n15623_), .A2(new_n5991_), .ZN(new_n15624_));
  AOI21_X1   g15432(.A1(new_n15620_), .A2(\asqrt[33] ), .B(new_n15624_), .ZN(new_n15625_));
  NOR2_X1    g15433(.A1(new_n15625_), .A2(new_n15619_), .ZN(new_n15626_));
  AOI22_X1   g15434(.A1(new_n15620_), .A2(\asqrt[33] ), .B1(new_n15618_), .B2(new_n15611_), .ZN(new_n15627_));
  NAND2_X1   g15435(.A1(new_n15283_), .A2(\asqrt[34] ), .ZN(new_n15628_));
  NOR4_X1    g15436(.A1(new_n15447_), .A2(\asqrt[34] ), .A3(new_n15012_), .A4(new_n15283_), .ZN(new_n15629_));
  XOR2_X1    g15437(.A1(new_n15629_), .A2(new_n15628_), .Z(new_n15630_));
  NAND2_X1   g15438(.A1(new_n15630_), .A2(new_n5626_), .ZN(new_n15631_));
  INV_X1     g15439(.I(new_n15631_), .ZN(new_n15632_));
  OAI21_X1   g15440(.A1(new_n15627_), .A2(new_n5991_), .B(new_n15632_), .ZN(new_n15633_));
  NAND2_X1   g15441(.A1(new_n15633_), .A2(new_n15626_), .ZN(new_n15634_));
  OAI22_X1   g15442(.A1(new_n15627_), .A2(new_n5991_), .B1(new_n15625_), .B2(new_n15619_), .ZN(new_n15635_));
  NAND2_X1   g15443(.A1(new_n15024_), .A2(\asqrt[35] ), .ZN(new_n15636_));
  NOR4_X1    g15444(.A1(new_n15447_), .A2(\asqrt[35] ), .A3(new_n15019_), .A4(new_n15024_), .ZN(new_n15637_));
  XOR2_X1    g15445(.A1(new_n15637_), .A2(new_n15636_), .Z(new_n15638_));
  NAND2_X1   g15446(.A1(new_n15638_), .A2(new_n5273_), .ZN(new_n15639_));
  AOI21_X1   g15447(.A1(new_n15635_), .A2(\asqrt[35] ), .B(new_n15639_), .ZN(new_n15640_));
  NOR2_X1    g15448(.A1(new_n15640_), .A2(new_n15634_), .ZN(new_n15641_));
  AOI22_X1   g15449(.A1(new_n15635_), .A2(\asqrt[35] ), .B1(new_n15633_), .B2(new_n15626_), .ZN(new_n15642_));
  NOR4_X1    g15450(.A1(new_n15447_), .A2(\asqrt[36] ), .A3(new_n15027_), .A4(new_n15290_), .ZN(new_n15643_));
  AOI21_X1   g15451(.A1(new_n15636_), .A2(new_n15023_), .B(new_n5273_), .ZN(new_n15644_));
  NOR2_X1    g15452(.A1(new_n15643_), .A2(new_n15644_), .ZN(new_n15645_));
  NAND2_X1   g15453(.A1(new_n15645_), .A2(new_n4973_), .ZN(new_n15646_));
  INV_X1     g15454(.I(new_n15646_), .ZN(new_n15647_));
  OAI21_X1   g15455(.A1(new_n15642_), .A2(new_n5273_), .B(new_n15647_), .ZN(new_n15648_));
  NAND2_X1   g15456(.A1(new_n15648_), .A2(new_n15641_), .ZN(new_n15649_));
  OAI22_X1   g15457(.A1(new_n15642_), .A2(new_n5273_), .B1(new_n15640_), .B2(new_n15634_), .ZN(new_n15650_));
  NAND2_X1   g15458(.A1(new_n15039_), .A2(\asqrt[37] ), .ZN(new_n15651_));
  NOR4_X1    g15459(.A1(new_n15447_), .A2(\asqrt[37] ), .A3(new_n15034_), .A4(new_n15039_), .ZN(new_n15652_));
  XOR2_X1    g15460(.A1(new_n15652_), .A2(new_n15651_), .Z(new_n15653_));
  NAND2_X1   g15461(.A1(new_n15653_), .A2(new_n4645_), .ZN(new_n15654_));
  AOI21_X1   g15462(.A1(new_n15650_), .A2(\asqrt[37] ), .B(new_n15654_), .ZN(new_n15655_));
  NOR2_X1    g15463(.A1(new_n15655_), .A2(new_n15649_), .ZN(new_n15656_));
  AOI22_X1   g15464(.A1(new_n15650_), .A2(\asqrt[37] ), .B1(new_n15648_), .B2(new_n15641_), .ZN(new_n15657_));
  NOR4_X1    g15465(.A1(new_n15447_), .A2(\asqrt[38] ), .A3(new_n15042_), .A4(new_n15297_), .ZN(new_n15658_));
  AOI21_X1   g15466(.A1(new_n15651_), .A2(new_n15038_), .B(new_n4645_), .ZN(new_n15659_));
  NOR2_X1    g15467(.A1(new_n15658_), .A2(new_n15659_), .ZN(new_n15660_));
  NAND2_X1   g15468(.A1(new_n15660_), .A2(new_n4330_), .ZN(new_n15661_));
  INV_X1     g15469(.I(new_n15661_), .ZN(new_n15662_));
  OAI21_X1   g15470(.A1(new_n15657_), .A2(new_n4645_), .B(new_n15662_), .ZN(new_n15663_));
  NAND2_X1   g15471(.A1(new_n15663_), .A2(new_n15656_), .ZN(new_n15664_));
  OAI22_X1   g15472(.A1(new_n15657_), .A2(new_n4645_), .B1(new_n15655_), .B2(new_n15649_), .ZN(new_n15665_));
  NAND2_X1   g15473(.A1(new_n15054_), .A2(\asqrt[39] ), .ZN(new_n15666_));
  NOR4_X1    g15474(.A1(new_n15447_), .A2(\asqrt[39] ), .A3(new_n15049_), .A4(new_n15054_), .ZN(new_n15667_));
  XOR2_X1    g15475(.A1(new_n15667_), .A2(new_n15666_), .Z(new_n15668_));
  NAND2_X1   g15476(.A1(new_n15668_), .A2(new_n4018_), .ZN(new_n15669_));
  AOI21_X1   g15477(.A1(new_n15665_), .A2(\asqrt[39] ), .B(new_n15669_), .ZN(new_n15670_));
  NOR2_X1    g15478(.A1(new_n15670_), .A2(new_n15664_), .ZN(new_n15671_));
  AOI22_X1   g15479(.A1(new_n15665_), .A2(\asqrt[39] ), .B1(new_n15663_), .B2(new_n15656_), .ZN(new_n15672_));
  NAND2_X1   g15480(.A1(new_n15304_), .A2(\asqrt[40] ), .ZN(new_n15673_));
  NOR4_X1    g15481(.A1(new_n15447_), .A2(\asqrt[40] ), .A3(new_n15057_), .A4(new_n15304_), .ZN(new_n15674_));
  XOR2_X1    g15482(.A1(new_n15674_), .A2(new_n15673_), .Z(new_n15675_));
  NAND2_X1   g15483(.A1(new_n15675_), .A2(new_n3760_), .ZN(new_n15676_));
  INV_X1     g15484(.I(new_n15676_), .ZN(new_n15677_));
  OAI21_X1   g15485(.A1(new_n15672_), .A2(new_n4018_), .B(new_n15677_), .ZN(new_n15678_));
  NAND2_X1   g15486(.A1(new_n15678_), .A2(new_n15671_), .ZN(new_n15679_));
  OAI22_X1   g15487(.A1(new_n15672_), .A2(new_n4018_), .B1(new_n15670_), .B2(new_n15664_), .ZN(new_n15680_));
  NOR4_X1    g15488(.A1(new_n15447_), .A2(\asqrt[41] ), .A3(new_n15064_), .A4(new_n15069_), .ZN(new_n15681_));
  AOI21_X1   g15489(.A1(new_n15673_), .A2(new_n15303_), .B(new_n3760_), .ZN(new_n15682_));
  NOR2_X1    g15490(.A1(new_n15681_), .A2(new_n15682_), .ZN(new_n15683_));
  NAND2_X1   g15491(.A1(new_n15683_), .A2(new_n3481_), .ZN(new_n15684_));
  AOI21_X1   g15492(.A1(new_n15680_), .A2(\asqrt[41] ), .B(new_n15684_), .ZN(new_n15685_));
  NOR2_X1    g15493(.A1(new_n15685_), .A2(new_n15679_), .ZN(new_n15686_));
  AOI22_X1   g15494(.A1(new_n15680_), .A2(\asqrt[41] ), .B1(new_n15678_), .B2(new_n15671_), .ZN(new_n15687_));
  NAND2_X1   g15495(.A1(new_n15311_), .A2(\asqrt[42] ), .ZN(new_n15688_));
  NOR4_X1    g15496(.A1(new_n15447_), .A2(\asqrt[42] ), .A3(new_n15072_), .A4(new_n15311_), .ZN(new_n15689_));
  XOR2_X1    g15497(.A1(new_n15689_), .A2(new_n15688_), .Z(new_n15690_));
  NAND2_X1   g15498(.A1(new_n15690_), .A2(new_n3208_), .ZN(new_n15691_));
  INV_X1     g15499(.I(new_n15691_), .ZN(new_n15692_));
  OAI21_X1   g15500(.A1(new_n15687_), .A2(new_n3481_), .B(new_n15692_), .ZN(new_n15693_));
  NAND2_X1   g15501(.A1(new_n15693_), .A2(new_n15686_), .ZN(new_n15694_));
  OAI22_X1   g15502(.A1(new_n15687_), .A2(new_n3481_), .B1(new_n15685_), .B2(new_n15679_), .ZN(new_n15695_));
  NOR4_X1    g15503(.A1(new_n15447_), .A2(\asqrt[43] ), .A3(new_n15079_), .A4(new_n15084_), .ZN(new_n15696_));
  AOI21_X1   g15504(.A1(new_n15688_), .A2(new_n15310_), .B(new_n3208_), .ZN(new_n15697_));
  NOR2_X1    g15505(.A1(new_n15696_), .A2(new_n15697_), .ZN(new_n15698_));
  NAND2_X1   g15506(.A1(new_n15698_), .A2(new_n2941_), .ZN(new_n15699_));
  AOI21_X1   g15507(.A1(new_n15695_), .A2(\asqrt[43] ), .B(new_n15699_), .ZN(new_n15700_));
  NOR2_X1    g15508(.A1(new_n15700_), .A2(new_n15694_), .ZN(new_n15701_));
  AOI22_X1   g15509(.A1(new_n15695_), .A2(\asqrt[43] ), .B1(new_n15693_), .B2(new_n15686_), .ZN(new_n15702_));
  NAND2_X1   g15510(.A1(new_n15318_), .A2(\asqrt[44] ), .ZN(new_n15703_));
  NOR4_X1    g15511(.A1(new_n15447_), .A2(\asqrt[44] ), .A3(new_n15087_), .A4(new_n15318_), .ZN(new_n15704_));
  XOR2_X1    g15512(.A1(new_n15704_), .A2(new_n15703_), .Z(new_n15705_));
  NAND2_X1   g15513(.A1(new_n15705_), .A2(new_n2728_), .ZN(new_n15706_));
  INV_X1     g15514(.I(new_n15706_), .ZN(new_n15707_));
  OAI21_X1   g15515(.A1(new_n15702_), .A2(new_n2941_), .B(new_n15707_), .ZN(new_n15708_));
  NAND2_X1   g15516(.A1(new_n15708_), .A2(new_n15701_), .ZN(new_n15709_));
  OAI22_X1   g15517(.A1(new_n15702_), .A2(new_n2941_), .B1(new_n15700_), .B2(new_n15694_), .ZN(new_n15710_));
  NOR4_X1    g15518(.A1(new_n15447_), .A2(\asqrt[45] ), .A3(new_n15094_), .A4(new_n15099_), .ZN(new_n15711_));
  AOI21_X1   g15519(.A1(new_n15703_), .A2(new_n15317_), .B(new_n2728_), .ZN(new_n15712_));
  NOR2_X1    g15520(.A1(new_n15711_), .A2(new_n15712_), .ZN(new_n15713_));
  NAND2_X1   g15521(.A1(new_n15713_), .A2(new_n2488_), .ZN(new_n15714_));
  AOI21_X1   g15522(.A1(new_n15710_), .A2(\asqrt[45] ), .B(new_n15714_), .ZN(new_n15715_));
  NOR2_X1    g15523(.A1(new_n15715_), .A2(new_n15709_), .ZN(new_n15716_));
  AOI22_X1   g15524(.A1(new_n15710_), .A2(\asqrt[45] ), .B1(new_n15708_), .B2(new_n15701_), .ZN(new_n15717_));
  NAND2_X1   g15525(.A1(new_n15325_), .A2(\asqrt[46] ), .ZN(new_n15718_));
  NOR4_X1    g15526(.A1(new_n15447_), .A2(\asqrt[46] ), .A3(new_n15102_), .A4(new_n15325_), .ZN(new_n15719_));
  XOR2_X1    g15527(.A1(new_n15719_), .A2(new_n15718_), .Z(new_n15720_));
  NAND2_X1   g15528(.A1(new_n15720_), .A2(new_n2253_), .ZN(new_n15721_));
  INV_X1     g15529(.I(new_n15721_), .ZN(new_n15722_));
  OAI21_X1   g15530(.A1(new_n15717_), .A2(new_n2488_), .B(new_n15722_), .ZN(new_n15723_));
  NAND2_X1   g15531(.A1(new_n15723_), .A2(new_n15716_), .ZN(new_n15724_));
  OAI22_X1   g15532(.A1(new_n15717_), .A2(new_n2488_), .B1(new_n15715_), .B2(new_n15709_), .ZN(new_n15725_));
  NAND2_X1   g15533(.A1(new_n15114_), .A2(\asqrt[47] ), .ZN(new_n15726_));
  NOR4_X1    g15534(.A1(new_n15447_), .A2(\asqrt[47] ), .A3(new_n15109_), .A4(new_n15114_), .ZN(new_n15727_));
  XOR2_X1    g15535(.A1(new_n15727_), .A2(new_n15726_), .Z(new_n15728_));
  NAND2_X1   g15536(.A1(new_n15728_), .A2(new_n2046_), .ZN(new_n15729_));
  AOI21_X1   g15537(.A1(new_n15725_), .A2(\asqrt[47] ), .B(new_n15729_), .ZN(new_n15730_));
  NOR2_X1    g15538(.A1(new_n15730_), .A2(new_n15724_), .ZN(new_n15731_));
  AOI22_X1   g15539(.A1(new_n15725_), .A2(\asqrt[47] ), .B1(new_n15723_), .B2(new_n15716_), .ZN(new_n15732_));
  NOR4_X1    g15540(.A1(new_n15447_), .A2(\asqrt[48] ), .A3(new_n15117_), .A4(new_n15332_), .ZN(new_n15733_));
  AOI21_X1   g15541(.A1(new_n15726_), .A2(new_n15113_), .B(new_n2046_), .ZN(new_n15734_));
  NOR2_X1    g15542(.A1(new_n15733_), .A2(new_n15734_), .ZN(new_n15735_));
  NAND2_X1   g15543(.A1(new_n15735_), .A2(new_n1854_), .ZN(new_n15736_));
  INV_X1     g15544(.I(new_n15736_), .ZN(new_n15737_));
  OAI21_X1   g15545(.A1(new_n15732_), .A2(new_n2046_), .B(new_n15737_), .ZN(new_n15738_));
  NAND2_X1   g15546(.A1(new_n15738_), .A2(new_n15731_), .ZN(new_n15739_));
  OAI22_X1   g15547(.A1(new_n15732_), .A2(new_n2046_), .B1(new_n15730_), .B2(new_n15724_), .ZN(new_n15740_));
  NAND2_X1   g15548(.A1(new_n15129_), .A2(\asqrt[49] ), .ZN(new_n15741_));
  NOR4_X1    g15549(.A1(new_n15447_), .A2(\asqrt[49] ), .A3(new_n15124_), .A4(new_n15129_), .ZN(new_n15742_));
  XOR2_X1    g15550(.A1(new_n15742_), .A2(new_n15741_), .Z(new_n15743_));
  NAND2_X1   g15551(.A1(new_n15743_), .A2(new_n1595_), .ZN(new_n15744_));
  AOI21_X1   g15552(.A1(new_n15740_), .A2(\asqrt[49] ), .B(new_n15744_), .ZN(new_n15745_));
  NOR2_X1    g15553(.A1(new_n15745_), .A2(new_n15739_), .ZN(new_n15746_));
  AOI22_X1   g15554(.A1(new_n15740_), .A2(\asqrt[49] ), .B1(new_n15738_), .B2(new_n15731_), .ZN(new_n15747_));
  NOR4_X1    g15555(.A1(new_n15447_), .A2(\asqrt[50] ), .A3(new_n15132_), .A4(new_n15339_), .ZN(new_n15748_));
  AOI21_X1   g15556(.A1(new_n15741_), .A2(new_n15128_), .B(new_n1595_), .ZN(new_n15749_));
  NOR2_X1    g15557(.A1(new_n15748_), .A2(new_n15749_), .ZN(new_n15750_));
  NAND2_X1   g15558(.A1(new_n15750_), .A2(new_n1436_), .ZN(new_n15751_));
  INV_X1     g15559(.I(new_n15751_), .ZN(new_n15752_));
  OAI21_X1   g15560(.A1(new_n15747_), .A2(new_n1595_), .B(new_n15752_), .ZN(new_n15753_));
  NAND2_X1   g15561(.A1(new_n15753_), .A2(new_n15746_), .ZN(new_n15754_));
  OAI22_X1   g15562(.A1(new_n15747_), .A2(new_n1595_), .B1(new_n15745_), .B2(new_n15739_), .ZN(new_n15755_));
  NAND2_X1   g15563(.A1(new_n15144_), .A2(\asqrt[51] ), .ZN(new_n15756_));
  NOR4_X1    g15564(.A1(new_n15447_), .A2(\asqrt[51] ), .A3(new_n15139_), .A4(new_n15144_), .ZN(new_n15757_));
  XOR2_X1    g15565(.A1(new_n15757_), .A2(new_n15756_), .Z(new_n15758_));
  NAND2_X1   g15566(.A1(new_n15758_), .A2(new_n1260_), .ZN(new_n15759_));
  AOI21_X1   g15567(.A1(new_n15755_), .A2(\asqrt[51] ), .B(new_n15759_), .ZN(new_n15760_));
  NOR2_X1    g15568(.A1(new_n15760_), .A2(new_n15754_), .ZN(new_n15761_));
  AOI22_X1   g15569(.A1(new_n15755_), .A2(\asqrt[51] ), .B1(new_n15753_), .B2(new_n15746_), .ZN(new_n15762_));
  NAND2_X1   g15570(.A1(new_n15346_), .A2(\asqrt[52] ), .ZN(new_n15763_));
  NOR4_X1    g15571(.A1(new_n15447_), .A2(\asqrt[52] ), .A3(new_n15147_), .A4(new_n15346_), .ZN(new_n15764_));
  XOR2_X1    g15572(.A1(new_n15764_), .A2(new_n15763_), .Z(new_n15765_));
  NAND2_X1   g15573(.A1(new_n15765_), .A2(new_n1096_), .ZN(new_n15766_));
  INV_X1     g15574(.I(new_n15766_), .ZN(new_n15767_));
  OAI21_X1   g15575(.A1(new_n15762_), .A2(new_n1260_), .B(new_n15767_), .ZN(new_n15768_));
  NAND2_X1   g15576(.A1(new_n15768_), .A2(new_n15761_), .ZN(new_n15769_));
  OAI22_X1   g15577(.A1(new_n15762_), .A2(new_n1260_), .B1(new_n15760_), .B2(new_n15754_), .ZN(new_n15770_));
  NOR4_X1    g15578(.A1(new_n15447_), .A2(\asqrt[53] ), .A3(new_n15153_), .A4(new_n15158_), .ZN(new_n15771_));
  AOI21_X1   g15579(.A1(new_n15763_), .A2(new_n15345_), .B(new_n1096_), .ZN(new_n15772_));
  NOR2_X1    g15580(.A1(new_n15771_), .A2(new_n15772_), .ZN(new_n15773_));
  NAND2_X1   g15581(.A1(new_n15773_), .A2(new_n970_), .ZN(new_n15774_));
  AOI21_X1   g15582(.A1(new_n15770_), .A2(\asqrt[53] ), .B(new_n15774_), .ZN(new_n15775_));
  NOR2_X1    g15583(.A1(new_n15775_), .A2(new_n15769_), .ZN(new_n15776_));
  AOI22_X1   g15584(.A1(new_n15770_), .A2(\asqrt[53] ), .B1(new_n15768_), .B2(new_n15761_), .ZN(new_n15777_));
  NAND2_X1   g15585(.A1(new_n15353_), .A2(\asqrt[54] ), .ZN(new_n15778_));
  NOR4_X1    g15586(.A1(new_n15447_), .A2(\asqrt[54] ), .A3(new_n15160_), .A4(new_n15353_), .ZN(new_n15779_));
  XOR2_X1    g15587(.A1(new_n15779_), .A2(new_n15778_), .Z(new_n15780_));
  NAND2_X1   g15588(.A1(new_n15780_), .A2(new_n825_), .ZN(new_n15781_));
  INV_X1     g15589(.I(new_n15781_), .ZN(new_n15782_));
  OAI21_X1   g15590(.A1(new_n15777_), .A2(new_n970_), .B(new_n15782_), .ZN(new_n15783_));
  NAND2_X1   g15591(.A1(new_n15783_), .A2(new_n15776_), .ZN(new_n15784_));
  OAI22_X1   g15592(.A1(new_n15777_), .A2(new_n970_), .B1(new_n15775_), .B2(new_n15769_), .ZN(new_n15785_));
  NOR4_X1    g15593(.A1(new_n15447_), .A2(\asqrt[55] ), .A3(new_n15166_), .A4(new_n15171_), .ZN(new_n15786_));
  AOI21_X1   g15594(.A1(new_n15778_), .A2(new_n15352_), .B(new_n825_), .ZN(new_n15787_));
  NOR2_X1    g15595(.A1(new_n15786_), .A2(new_n15787_), .ZN(new_n15788_));
  NAND2_X1   g15596(.A1(new_n15788_), .A2(new_n724_), .ZN(new_n15789_));
  AOI21_X1   g15597(.A1(new_n15785_), .A2(\asqrt[55] ), .B(new_n15789_), .ZN(new_n15790_));
  NOR2_X1    g15598(.A1(new_n15790_), .A2(new_n15784_), .ZN(new_n15791_));
  AOI22_X1   g15599(.A1(new_n15785_), .A2(\asqrt[55] ), .B1(new_n15783_), .B2(new_n15776_), .ZN(new_n15792_));
  NAND2_X1   g15600(.A1(new_n15360_), .A2(\asqrt[56] ), .ZN(new_n15793_));
  NOR4_X1    g15601(.A1(new_n15447_), .A2(\asqrt[56] ), .A3(new_n15173_), .A4(new_n15360_), .ZN(new_n15794_));
  XOR2_X1    g15602(.A1(new_n15794_), .A2(new_n15793_), .Z(new_n15795_));
  NAND2_X1   g15603(.A1(new_n15795_), .A2(new_n587_), .ZN(new_n15796_));
  INV_X1     g15604(.I(new_n15796_), .ZN(new_n15797_));
  OAI21_X1   g15605(.A1(new_n15792_), .A2(new_n724_), .B(new_n15797_), .ZN(new_n15798_));
  NAND2_X1   g15606(.A1(new_n15798_), .A2(new_n15791_), .ZN(new_n15799_));
  NAND2_X1   g15607(.A1(new_n15785_), .A2(\asqrt[55] ), .ZN(new_n15800_));
  AOI21_X1   g15608(.A1(new_n15800_), .A2(new_n15784_), .B(new_n724_), .ZN(new_n15801_));
  OAI21_X1   g15609(.A1(new_n15791_), .A2(new_n15801_), .B(\asqrt[57] ), .ZN(new_n15802_));
  NOR2_X1    g15610(.A1(new_n15363_), .A2(new_n587_), .ZN(new_n15803_));
  NOR4_X1    g15611(.A1(new_n15447_), .A2(\asqrt[57] ), .A3(new_n15179_), .A4(new_n15184_), .ZN(new_n15804_));
  XNOR2_X1   g15612(.A1(new_n15804_), .A2(new_n15803_), .ZN(new_n15805_));
  NAND2_X1   g15613(.A1(new_n15805_), .A2(new_n504_), .ZN(new_n15806_));
  INV_X1     g15614(.I(new_n15806_), .ZN(new_n15807_));
  AOI21_X1   g15615(.A1(new_n15802_), .A2(new_n15807_), .B(new_n15799_), .ZN(new_n15808_));
  OAI22_X1   g15616(.A1(new_n15792_), .A2(new_n724_), .B1(new_n15790_), .B2(new_n15784_), .ZN(new_n15809_));
  AOI22_X1   g15617(.A1(new_n15809_), .A2(\asqrt[57] ), .B1(new_n15798_), .B2(new_n15791_), .ZN(new_n15810_));
  NOR4_X1    g15618(.A1(new_n15447_), .A2(\asqrt[58] ), .A3(new_n15186_), .A4(new_n15367_), .ZN(new_n15811_));
  XOR2_X1    g15619(.A1(new_n15811_), .A2(new_n15411_), .Z(new_n15812_));
  NAND2_X1   g15620(.A1(new_n15812_), .A2(new_n376_), .ZN(new_n15813_));
  INV_X1     g15621(.I(new_n15813_), .ZN(new_n15814_));
  OAI21_X1   g15622(.A1(new_n15810_), .A2(new_n504_), .B(new_n15814_), .ZN(new_n15815_));
  NAND2_X1   g15623(.A1(new_n15815_), .A2(new_n15808_), .ZN(new_n15816_));
  AOI21_X1   g15624(.A1(new_n15799_), .A2(new_n15802_), .B(new_n504_), .ZN(new_n15817_));
  OAI21_X1   g15625(.A1(new_n15808_), .A2(new_n15817_), .B(\asqrt[59] ), .ZN(new_n15818_));
  NOR4_X1    g15626(.A1(new_n15447_), .A2(\asqrt[59] ), .A3(new_n15192_), .A4(new_n15197_), .ZN(new_n15819_));
  XOR2_X1    g15627(.A1(new_n15819_), .A2(new_n15389_), .Z(new_n15820_));
  AND2_X2    g15628(.A1(new_n15820_), .A2(new_n275_), .Z(new_n15821_));
  AOI21_X1   g15629(.A1(new_n15818_), .A2(new_n15821_), .B(new_n15816_), .ZN(new_n15822_));
  OAI22_X1   g15630(.A1(new_n15470_), .A2(new_n13760_), .B1(new_n15458_), .B2(new_n15468_), .ZN(new_n15823_));
  AOI22_X1   g15631(.A1(new_n15823_), .A2(\asqrt[18] ), .B1(new_n15477_), .B2(new_n15469_), .ZN(new_n15824_));
  INV_X1     g15632(.I(new_n15511_), .ZN(new_n15825_));
  OAI21_X1   g15633(.A1(new_n15824_), .A2(new_n12657_), .B(new_n15825_), .ZN(new_n15826_));
  AOI21_X1   g15634(.A1(new_n15823_), .A2(\asqrt[18] ), .B(new_n15485_), .ZN(new_n15827_));
  OAI22_X1   g15635(.A1(new_n15824_), .A2(new_n12657_), .B1(new_n15827_), .B2(new_n15514_), .ZN(new_n15828_));
  AOI22_X1   g15636(.A1(new_n15828_), .A2(\asqrt[20] ), .B1(new_n15826_), .B2(new_n15515_), .ZN(new_n15829_));
  INV_X1     g15637(.I(new_n15530_), .ZN(new_n15830_));
  OAI21_X1   g15638(.A1(new_n15829_), .A2(new_n11631_), .B(new_n15830_), .ZN(new_n15831_));
  NAND2_X1   g15639(.A1(new_n15831_), .A2(new_n15534_), .ZN(new_n15832_));
  AOI21_X1   g15640(.A1(new_n15828_), .A2(\asqrt[20] ), .B(new_n15521_), .ZN(new_n15833_));
  OAI22_X1   g15641(.A1(new_n15829_), .A2(new_n11631_), .B1(new_n15833_), .B2(new_n15533_), .ZN(new_n15834_));
  AOI21_X1   g15642(.A1(new_n15834_), .A2(\asqrt[22] ), .B(new_n15540_), .ZN(new_n15835_));
  NOR2_X1    g15643(.A1(new_n15835_), .A2(new_n15832_), .ZN(new_n15836_));
  AOI22_X1   g15644(.A1(new_n15834_), .A2(\asqrt[22] ), .B1(new_n15831_), .B2(new_n15534_), .ZN(new_n15837_));
  INV_X1     g15645(.I(new_n15549_), .ZN(new_n15838_));
  OAI21_X1   g15646(.A1(new_n15837_), .A2(new_n10614_), .B(new_n15838_), .ZN(new_n15839_));
  NAND2_X1   g15647(.A1(new_n15839_), .A2(new_n15836_), .ZN(new_n15840_));
  OAI22_X1   g15648(.A1(new_n15837_), .A2(new_n10614_), .B1(new_n15835_), .B2(new_n15832_), .ZN(new_n15841_));
  AOI21_X1   g15649(.A1(new_n15841_), .A2(\asqrt[24] ), .B(new_n15556_), .ZN(new_n15842_));
  NOR2_X1    g15650(.A1(new_n15842_), .A2(new_n15840_), .ZN(new_n15843_));
  AOI22_X1   g15651(.A1(new_n15841_), .A2(\asqrt[24] ), .B1(new_n15839_), .B2(new_n15836_), .ZN(new_n15844_));
  INV_X1     g15652(.I(new_n15564_), .ZN(new_n15845_));
  OAI21_X1   g15653(.A1(new_n15844_), .A2(new_n9672_), .B(new_n15845_), .ZN(new_n15846_));
  NAND2_X1   g15654(.A1(new_n15846_), .A2(new_n15843_), .ZN(new_n15847_));
  OAI22_X1   g15655(.A1(new_n15844_), .A2(new_n9672_), .B1(new_n15842_), .B2(new_n15840_), .ZN(new_n15848_));
  AOI21_X1   g15656(.A1(new_n15848_), .A2(\asqrt[26] ), .B(new_n15571_), .ZN(new_n15849_));
  NOR2_X1    g15657(.A1(new_n15849_), .A2(new_n15847_), .ZN(new_n15850_));
  AOI22_X1   g15658(.A1(new_n15848_), .A2(\asqrt[26] ), .B1(new_n15846_), .B2(new_n15843_), .ZN(new_n15851_));
  INV_X1     g15659(.I(new_n15579_), .ZN(new_n15852_));
  OAI21_X1   g15660(.A1(new_n15851_), .A2(new_n8763_), .B(new_n15852_), .ZN(new_n15853_));
  NAND2_X1   g15661(.A1(new_n15853_), .A2(new_n15850_), .ZN(new_n15854_));
  OAI22_X1   g15662(.A1(new_n15851_), .A2(new_n8763_), .B1(new_n15849_), .B2(new_n15847_), .ZN(new_n15855_));
  AOI21_X1   g15663(.A1(new_n15855_), .A2(\asqrt[28] ), .B(new_n15586_), .ZN(new_n15856_));
  NOR2_X1    g15664(.A1(new_n15856_), .A2(new_n15854_), .ZN(new_n15857_));
  AOI22_X1   g15665(.A1(new_n15855_), .A2(\asqrt[28] ), .B1(new_n15853_), .B2(new_n15850_), .ZN(new_n15858_));
  INV_X1     g15666(.I(new_n15594_), .ZN(new_n15859_));
  OAI21_X1   g15667(.A1(new_n15858_), .A2(new_n7931_), .B(new_n15859_), .ZN(new_n15860_));
  NAND2_X1   g15668(.A1(new_n15860_), .A2(new_n15857_), .ZN(new_n15861_));
  OAI22_X1   g15669(.A1(new_n15858_), .A2(new_n7931_), .B1(new_n15856_), .B2(new_n15854_), .ZN(new_n15862_));
  AOI21_X1   g15670(.A1(new_n15862_), .A2(\asqrt[30] ), .B(new_n15601_), .ZN(new_n15863_));
  NOR2_X1    g15671(.A1(new_n15863_), .A2(new_n15861_), .ZN(new_n15864_));
  AOI22_X1   g15672(.A1(new_n15862_), .A2(\asqrt[30] ), .B1(new_n15860_), .B2(new_n15857_), .ZN(new_n15865_));
  INV_X1     g15673(.I(new_n15609_), .ZN(new_n15866_));
  OAI21_X1   g15674(.A1(new_n15865_), .A2(new_n7110_), .B(new_n15866_), .ZN(new_n15867_));
  NAND2_X1   g15675(.A1(new_n15867_), .A2(new_n15864_), .ZN(new_n15868_));
  OAI22_X1   g15676(.A1(new_n15865_), .A2(new_n7110_), .B1(new_n15863_), .B2(new_n15861_), .ZN(new_n15869_));
  AOI21_X1   g15677(.A1(new_n15869_), .A2(\asqrt[32] ), .B(new_n15616_), .ZN(new_n15870_));
  NOR2_X1    g15678(.A1(new_n15870_), .A2(new_n15868_), .ZN(new_n15871_));
  AOI22_X1   g15679(.A1(new_n15869_), .A2(\asqrt[32] ), .B1(new_n15867_), .B2(new_n15864_), .ZN(new_n15872_));
  INV_X1     g15680(.I(new_n15624_), .ZN(new_n15873_));
  OAI21_X1   g15681(.A1(new_n15872_), .A2(new_n6365_), .B(new_n15873_), .ZN(new_n15874_));
  NAND2_X1   g15682(.A1(new_n15874_), .A2(new_n15871_), .ZN(new_n15875_));
  OAI22_X1   g15683(.A1(new_n15872_), .A2(new_n6365_), .B1(new_n15870_), .B2(new_n15868_), .ZN(new_n15876_));
  AOI21_X1   g15684(.A1(new_n15876_), .A2(\asqrt[34] ), .B(new_n15631_), .ZN(new_n15877_));
  NOR2_X1    g15685(.A1(new_n15877_), .A2(new_n15875_), .ZN(new_n15878_));
  AOI22_X1   g15686(.A1(new_n15876_), .A2(\asqrt[34] ), .B1(new_n15874_), .B2(new_n15871_), .ZN(new_n15879_));
  INV_X1     g15687(.I(new_n15639_), .ZN(new_n15880_));
  OAI21_X1   g15688(.A1(new_n15879_), .A2(new_n5626_), .B(new_n15880_), .ZN(new_n15881_));
  NAND2_X1   g15689(.A1(new_n15881_), .A2(new_n15878_), .ZN(new_n15882_));
  OAI22_X1   g15690(.A1(new_n15879_), .A2(new_n5626_), .B1(new_n15877_), .B2(new_n15875_), .ZN(new_n15883_));
  AOI21_X1   g15691(.A1(new_n15883_), .A2(\asqrt[36] ), .B(new_n15646_), .ZN(new_n15884_));
  NOR2_X1    g15692(.A1(new_n15884_), .A2(new_n15882_), .ZN(new_n15885_));
  AOI22_X1   g15693(.A1(new_n15883_), .A2(\asqrt[36] ), .B1(new_n15881_), .B2(new_n15878_), .ZN(new_n15886_));
  INV_X1     g15694(.I(new_n15654_), .ZN(new_n15887_));
  OAI21_X1   g15695(.A1(new_n15886_), .A2(new_n4973_), .B(new_n15887_), .ZN(new_n15888_));
  NAND2_X1   g15696(.A1(new_n15888_), .A2(new_n15885_), .ZN(new_n15889_));
  OAI22_X1   g15697(.A1(new_n15886_), .A2(new_n4973_), .B1(new_n15884_), .B2(new_n15882_), .ZN(new_n15890_));
  AOI21_X1   g15698(.A1(new_n15890_), .A2(\asqrt[38] ), .B(new_n15661_), .ZN(new_n15891_));
  NOR2_X1    g15699(.A1(new_n15891_), .A2(new_n15889_), .ZN(new_n15892_));
  AOI22_X1   g15700(.A1(new_n15890_), .A2(\asqrt[38] ), .B1(new_n15888_), .B2(new_n15885_), .ZN(new_n15893_));
  INV_X1     g15701(.I(new_n15669_), .ZN(new_n15894_));
  OAI21_X1   g15702(.A1(new_n15893_), .A2(new_n4330_), .B(new_n15894_), .ZN(new_n15895_));
  NAND2_X1   g15703(.A1(new_n15895_), .A2(new_n15892_), .ZN(new_n15896_));
  OAI22_X1   g15704(.A1(new_n15893_), .A2(new_n4330_), .B1(new_n15891_), .B2(new_n15889_), .ZN(new_n15897_));
  AOI21_X1   g15705(.A1(new_n15897_), .A2(\asqrt[40] ), .B(new_n15676_), .ZN(new_n15898_));
  NOR2_X1    g15706(.A1(new_n15898_), .A2(new_n15896_), .ZN(new_n15899_));
  AOI22_X1   g15707(.A1(new_n15897_), .A2(\asqrt[40] ), .B1(new_n15895_), .B2(new_n15892_), .ZN(new_n15900_));
  INV_X1     g15708(.I(new_n15684_), .ZN(new_n15901_));
  OAI21_X1   g15709(.A1(new_n15900_), .A2(new_n3760_), .B(new_n15901_), .ZN(new_n15902_));
  NAND2_X1   g15710(.A1(new_n15902_), .A2(new_n15899_), .ZN(new_n15903_));
  OAI22_X1   g15711(.A1(new_n15900_), .A2(new_n3760_), .B1(new_n15898_), .B2(new_n15896_), .ZN(new_n15904_));
  AOI21_X1   g15712(.A1(new_n15904_), .A2(\asqrt[42] ), .B(new_n15691_), .ZN(new_n15905_));
  NOR2_X1    g15713(.A1(new_n15905_), .A2(new_n15903_), .ZN(new_n15906_));
  AOI22_X1   g15714(.A1(new_n15904_), .A2(\asqrt[42] ), .B1(new_n15902_), .B2(new_n15899_), .ZN(new_n15907_));
  INV_X1     g15715(.I(new_n15699_), .ZN(new_n15908_));
  OAI21_X1   g15716(.A1(new_n15907_), .A2(new_n3208_), .B(new_n15908_), .ZN(new_n15909_));
  NAND2_X1   g15717(.A1(new_n15909_), .A2(new_n15906_), .ZN(new_n15910_));
  OAI22_X1   g15718(.A1(new_n15907_), .A2(new_n3208_), .B1(new_n15905_), .B2(new_n15903_), .ZN(new_n15911_));
  AOI21_X1   g15719(.A1(new_n15911_), .A2(\asqrt[44] ), .B(new_n15706_), .ZN(new_n15912_));
  NOR2_X1    g15720(.A1(new_n15912_), .A2(new_n15910_), .ZN(new_n15913_));
  AOI22_X1   g15721(.A1(new_n15911_), .A2(\asqrt[44] ), .B1(new_n15909_), .B2(new_n15906_), .ZN(new_n15914_));
  INV_X1     g15722(.I(new_n15714_), .ZN(new_n15915_));
  OAI21_X1   g15723(.A1(new_n15914_), .A2(new_n2728_), .B(new_n15915_), .ZN(new_n15916_));
  NAND2_X1   g15724(.A1(new_n15916_), .A2(new_n15913_), .ZN(new_n15917_));
  OAI22_X1   g15725(.A1(new_n15914_), .A2(new_n2728_), .B1(new_n15912_), .B2(new_n15910_), .ZN(new_n15918_));
  AOI21_X1   g15726(.A1(new_n15918_), .A2(\asqrt[46] ), .B(new_n15721_), .ZN(new_n15919_));
  NOR2_X1    g15727(.A1(new_n15919_), .A2(new_n15917_), .ZN(new_n15920_));
  AOI22_X1   g15728(.A1(new_n15918_), .A2(\asqrt[46] ), .B1(new_n15916_), .B2(new_n15913_), .ZN(new_n15921_));
  INV_X1     g15729(.I(new_n15729_), .ZN(new_n15922_));
  OAI21_X1   g15730(.A1(new_n15921_), .A2(new_n2253_), .B(new_n15922_), .ZN(new_n15923_));
  NAND2_X1   g15731(.A1(new_n15923_), .A2(new_n15920_), .ZN(new_n15924_));
  OAI22_X1   g15732(.A1(new_n15921_), .A2(new_n2253_), .B1(new_n15919_), .B2(new_n15917_), .ZN(new_n15925_));
  AOI21_X1   g15733(.A1(new_n15925_), .A2(\asqrt[48] ), .B(new_n15736_), .ZN(new_n15926_));
  NOR2_X1    g15734(.A1(new_n15926_), .A2(new_n15924_), .ZN(new_n15927_));
  AOI22_X1   g15735(.A1(new_n15925_), .A2(\asqrt[48] ), .B1(new_n15923_), .B2(new_n15920_), .ZN(new_n15928_));
  INV_X1     g15736(.I(new_n15744_), .ZN(new_n15929_));
  OAI21_X1   g15737(.A1(new_n15928_), .A2(new_n1854_), .B(new_n15929_), .ZN(new_n15930_));
  NAND2_X1   g15738(.A1(new_n15930_), .A2(new_n15927_), .ZN(new_n15931_));
  OAI22_X1   g15739(.A1(new_n15928_), .A2(new_n1854_), .B1(new_n15926_), .B2(new_n15924_), .ZN(new_n15932_));
  AOI21_X1   g15740(.A1(new_n15932_), .A2(\asqrt[50] ), .B(new_n15751_), .ZN(new_n15933_));
  NOR2_X1    g15741(.A1(new_n15933_), .A2(new_n15931_), .ZN(new_n15934_));
  AOI22_X1   g15742(.A1(new_n15932_), .A2(\asqrt[50] ), .B1(new_n15930_), .B2(new_n15927_), .ZN(new_n15935_));
  INV_X1     g15743(.I(new_n15759_), .ZN(new_n15936_));
  OAI21_X1   g15744(.A1(new_n15935_), .A2(new_n1436_), .B(new_n15936_), .ZN(new_n15937_));
  NAND2_X1   g15745(.A1(new_n15937_), .A2(new_n15934_), .ZN(new_n15938_));
  OAI22_X1   g15746(.A1(new_n15935_), .A2(new_n1436_), .B1(new_n15933_), .B2(new_n15931_), .ZN(new_n15939_));
  AOI21_X1   g15747(.A1(new_n15939_), .A2(\asqrt[52] ), .B(new_n15766_), .ZN(new_n15940_));
  NOR2_X1    g15748(.A1(new_n15940_), .A2(new_n15938_), .ZN(new_n15941_));
  AOI22_X1   g15749(.A1(new_n15939_), .A2(\asqrt[52] ), .B1(new_n15937_), .B2(new_n15934_), .ZN(new_n15942_));
  INV_X1     g15750(.I(new_n15774_), .ZN(new_n15943_));
  OAI21_X1   g15751(.A1(new_n15942_), .A2(new_n1096_), .B(new_n15943_), .ZN(new_n15944_));
  NAND2_X1   g15752(.A1(new_n15944_), .A2(new_n15941_), .ZN(new_n15945_));
  OAI22_X1   g15753(.A1(new_n15942_), .A2(new_n1096_), .B1(new_n15940_), .B2(new_n15938_), .ZN(new_n15946_));
  AOI21_X1   g15754(.A1(new_n15946_), .A2(\asqrt[54] ), .B(new_n15781_), .ZN(new_n15947_));
  NOR2_X1    g15755(.A1(new_n15947_), .A2(new_n15945_), .ZN(new_n15948_));
  AOI22_X1   g15756(.A1(new_n15946_), .A2(\asqrt[54] ), .B1(new_n15944_), .B2(new_n15941_), .ZN(new_n15949_));
  INV_X1     g15757(.I(new_n15789_), .ZN(new_n15950_));
  OAI21_X1   g15758(.A1(new_n15949_), .A2(new_n825_), .B(new_n15950_), .ZN(new_n15951_));
  NAND2_X1   g15759(.A1(new_n15951_), .A2(new_n15948_), .ZN(new_n15952_));
  OAI22_X1   g15760(.A1(new_n15949_), .A2(new_n825_), .B1(new_n15947_), .B2(new_n15945_), .ZN(new_n15953_));
  AOI21_X1   g15761(.A1(new_n15953_), .A2(\asqrt[56] ), .B(new_n15796_), .ZN(new_n15954_));
  NOR2_X1    g15762(.A1(new_n15954_), .A2(new_n15952_), .ZN(new_n15955_));
  AOI22_X1   g15763(.A1(new_n15953_), .A2(\asqrt[56] ), .B1(new_n15951_), .B2(new_n15948_), .ZN(new_n15956_));
  OAI21_X1   g15764(.A1(new_n15956_), .A2(new_n587_), .B(new_n15807_), .ZN(new_n15957_));
  NAND2_X1   g15765(.A1(new_n15957_), .A2(new_n15955_), .ZN(new_n15958_));
  NAND2_X1   g15766(.A1(new_n15946_), .A2(\asqrt[54] ), .ZN(new_n15959_));
  AOI21_X1   g15767(.A1(new_n15959_), .A2(new_n15945_), .B(new_n825_), .ZN(new_n15960_));
  OAI21_X1   g15768(.A1(new_n15948_), .A2(new_n15960_), .B(\asqrt[56] ), .ZN(new_n15961_));
  AOI21_X1   g15769(.A1(new_n15952_), .A2(new_n15961_), .B(new_n587_), .ZN(new_n15962_));
  OAI21_X1   g15770(.A1(new_n15955_), .A2(new_n15962_), .B(\asqrt[58] ), .ZN(new_n15963_));
  NAND2_X1   g15771(.A1(new_n15958_), .A2(new_n15963_), .ZN(new_n15964_));
  AOI22_X1   g15772(.A1(new_n15964_), .A2(\asqrt[59] ), .B1(new_n15815_), .B2(new_n15808_), .ZN(new_n15965_));
  NOR4_X1    g15773(.A1(new_n15447_), .A2(\asqrt[60] ), .A3(new_n15199_), .A4(new_n15374_), .ZN(new_n15966_));
  XOR2_X1    g15774(.A1(new_n15966_), .A2(new_n15413_), .Z(new_n15967_));
  NAND2_X1   g15775(.A1(new_n15967_), .A2(new_n229_), .ZN(new_n15968_));
  INV_X1     g15776(.I(new_n15968_), .ZN(new_n15969_));
  OAI21_X1   g15777(.A1(new_n15965_), .A2(new_n275_), .B(new_n15969_), .ZN(new_n15970_));
  OAI22_X1   g15778(.A1(new_n15956_), .A2(new_n587_), .B1(new_n15954_), .B2(new_n15952_), .ZN(new_n15971_));
  AOI21_X1   g15779(.A1(new_n15971_), .A2(\asqrt[58] ), .B(new_n15813_), .ZN(new_n15972_));
  NOR2_X1    g15780(.A1(new_n15972_), .A2(new_n15958_), .ZN(new_n15973_));
  AOI22_X1   g15781(.A1(new_n15971_), .A2(\asqrt[58] ), .B1(new_n15957_), .B2(new_n15955_), .ZN(new_n15974_));
  OAI21_X1   g15782(.A1(new_n15974_), .A2(new_n376_), .B(new_n15821_), .ZN(new_n15975_));
  NAND2_X1   g15783(.A1(new_n15975_), .A2(new_n15973_), .ZN(new_n15976_));
  AOI21_X1   g15784(.A1(new_n15958_), .A2(new_n15963_), .B(new_n376_), .ZN(new_n15977_));
  OAI21_X1   g15785(.A1(new_n15973_), .A2(new_n15977_), .B(\asqrt[60] ), .ZN(new_n15978_));
  AOI21_X1   g15786(.A1(new_n15976_), .A2(new_n15978_), .B(new_n229_), .ZN(new_n15979_));
  INV_X1     g15787(.I(new_n15417_), .ZN(new_n15980_));
  NOR2_X1    g15788(.A1(new_n15980_), .A2(\asqrt[62] ), .ZN(new_n15981_));
  INV_X1     g15789(.I(new_n15981_), .ZN(new_n15982_));
  NAND4_X1   g15790(.A1(new_n15979_), .A2(new_n15822_), .A3(new_n15970_), .A4(new_n15982_), .ZN(new_n15983_));
  NAND2_X1   g15791(.A1(new_n15435_), .A2(new_n15385_), .ZN(new_n15984_));
  OAI21_X1   g15792(.A1(\asqrt[14] ), .A2(new_n15984_), .B(new_n15395_), .ZN(new_n15985_));
  NAND2_X1   g15793(.A1(new_n15985_), .A2(new_n231_), .ZN(new_n15986_));
  INV_X1     g15794(.I(new_n15986_), .ZN(new_n15987_));
  NAND3_X1   g15795(.A1(new_n15983_), .A2(new_n15419_), .A3(new_n15987_), .ZN(new_n15988_));
  OAI22_X1   g15796(.A1(new_n15974_), .A2(new_n376_), .B1(new_n15972_), .B2(new_n15958_), .ZN(new_n15989_));
  AOI21_X1   g15797(.A1(new_n15989_), .A2(\asqrt[60] ), .B(new_n15968_), .ZN(new_n15990_));
  AOI22_X1   g15798(.A1(new_n15989_), .A2(\asqrt[60] ), .B1(new_n15975_), .B2(new_n15973_), .ZN(new_n15991_));
  OAI22_X1   g15799(.A1(new_n15991_), .A2(new_n229_), .B1(new_n15990_), .B2(new_n15976_), .ZN(new_n15992_));
  NOR4_X1    g15800(.A1(new_n15992_), .A2(\asqrt[62] ), .A3(new_n15409_), .A4(new_n15417_), .ZN(new_n15993_));
  AOI21_X1   g15801(.A1(new_n15410_), .A2(new_n15988_), .B(new_n15993_), .ZN(new_n15994_));
  INV_X1     g15802(.I(\a[24] ), .ZN(new_n15995_));
  OAI21_X1   g15803(.A1(new_n15386_), .A2(new_n15395_), .B(\asqrt[14] ), .ZN(new_n15996_));
  XOR2_X1    g15804(.A1(new_n15395_), .A2(\asqrt[63] ), .Z(new_n15997_));
  NAND2_X1   g15805(.A1(new_n15996_), .A2(new_n15997_), .ZN(new_n15998_));
  INV_X1     g15806(.I(new_n15998_), .ZN(new_n15999_));
  NAND3_X1   g15807(.A1(new_n15441_), .A2(new_n15379_), .A3(new_n15386_), .ZN(new_n16000_));
  INV_X1     g15808(.I(new_n16000_), .ZN(new_n16001_));
  NOR2_X1    g15809(.A1(new_n15999_), .A2(new_n16001_), .ZN(new_n16002_));
  NOR2_X1    g15810(.A1(\a[22] ), .A2(\a[23] ), .ZN(new_n16003_));
  INV_X1     g15811(.I(new_n16003_), .ZN(new_n16004_));
  NOR3_X1    g15812(.A1(new_n16002_), .A2(new_n15995_), .A3(new_n16004_), .ZN(new_n16005_));
  NAND2_X1   g15813(.A1(new_n15994_), .A2(new_n16005_), .ZN(new_n16006_));
  XOR2_X1    g15814(.A1(new_n16006_), .A2(\a[25] ), .Z(new_n16007_));
  INV_X1     g15815(.I(\a[25] ), .ZN(new_n16008_));
  NAND2_X1   g15816(.A1(new_n15970_), .A2(new_n15822_), .ZN(new_n16009_));
  NAND2_X1   g15817(.A1(new_n15979_), .A2(new_n15982_), .ZN(new_n16010_));
  OAI21_X1   g15818(.A1(new_n16010_), .A2(new_n16009_), .B(new_n15419_), .ZN(new_n16011_));
  OAI21_X1   g15819(.A1(new_n16011_), .A2(new_n15986_), .B(new_n15410_), .ZN(new_n16012_));
  NAND2_X1   g15820(.A1(new_n15993_), .A2(new_n15999_), .ZN(new_n16013_));
  NOR2_X1    g15821(.A1(new_n16013_), .A2(new_n16012_), .ZN(new_n16014_));
  NAND3_X1   g15822(.A1(new_n16014_), .A2(new_n15410_), .A3(new_n16000_), .ZN(new_n16015_));
  NAND2_X1   g15823(.A1(new_n15976_), .A2(new_n15978_), .ZN(new_n16016_));
  AOI22_X1   g15824(.A1(new_n16016_), .A2(\asqrt[61] ), .B1(new_n15970_), .B2(new_n15822_), .ZN(new_n16017_));
  NOR2_X1    g15825(.A1(new_n16017_), .A2(new_n196_), .ZN(new_n16018_));
  AOI21_X1   g15826(.A1(new_n15816_), .A2(new_n15818_), .B(new_n275_), .ZN(new_n16019_));
  OAI21_X1   g15827(.A1(new_n15822_), .A2(new_n16019_), .B(\asqrt[61] ), .ZN(new_n16020_));
  NAND4_X1   g15828(.A1(new_n16009_), .A2(new_n196_), .A3(new_n16020_), .A4(new_n15980_), .ZN(new_n16021_));
  INV_X1     g15829(.I(new_n16021_), .ZN(new_n16022_));
  NOR3_X1    g15830(.A1(new_n16013_), .A2(new_n16012_), .A3(new_n16000_), .ZN(\asqrt[13] ));
  NAND3_X1   g15831(.A1(\asqrt[13] ), .A2(new_n16018_), .A3(new_n16022_), .ZN(new_n16024_));
  OAI21_X1   g15832(.A1(new_n15992_), .A2(\asqrt[62] ), .B(new_n15417_), .ZN(new_n16025_));
  OAI21_X1   g15833(.A1(\asqrt[13] ), .A2(new_n16025_), .B(new_n16018_), .ZN(new_n16026_));
  NAND2_X1   g15834(.A1(new_n16026_), .A2(new_n16024_), .ZN(new_n16027_));
  INV_X1     g15835(.I(new_n16027_), .ZN(new_n16028_));
  NOR3_X1    g15836(.A1(new_n16016_), .A2(\asqrt[61] ), .A3(new_n15967_), .ZN(new_n16029_));
  NAND2_X1   g15837(.A1(\asqrt[13] ), .A2(new_n16029_), .ZN(new_n16030_));
  XOR2_X1    g15838(.A1(new_n16030_), .A2(new_n15979_), .Z(new_n16031_));
  NOR2_X1    g15839(.A1(new_n16031_), .A2(new_n196_), .ZN(new_n16032_));
  INV_X1     g15840(.I(new_n16032_), .ZN(new_n16033_));
  INV_X1     g15841(.I(\a[26] ), .ZN(new_n16034_));
  NOR2_X1    g15842(.A1(\a[24] ), .A2(\a[25] ), .ZN(new_n16035_));
  INV_X1     g15843(.I(new_n16035_), .ZN(new_n16036_));
  NOR3_X1    g15844(.A1(new_n15448_), .A2(new_n16034_), .A3(new_n16036_), .ZN(new_n16037_));
  NAND3_X1   g15845(.A1(new_n15399_), .A2(new_n15435_), .A3(new_n16037_), .ZN(new_n16038_));
  XOR2_X1    g15846(.A1(new_n16038_), .A2(\a[27] ), .Z(new_n16039_));
  INV_X1     g15847(.I(\a[27] ), .ZN(new_n16040_));
  NOR4_X1    g15848(.A1(new_n16013_), .A2(new_n16012_), .A3(new_n16040_), .A4(new_n16000_), .ZN(new_n16041_));
  NOR2_X1    g15849(.A1(new_n16039_), .A2(\a[26] ), .ZN(new_n16042_));
  OAI21_X1   g15850(.A1(new_n16041_), .A2(new_n16042_), .B(new_n16039_), .ZN(new_n16043_));
  INV_X1     g15851(.I(new_n16039_), .ZN(new_n16044_));
  NOR2_X1    g15852(.A1(new_n15990_), .A2(new_n15976_), .ZN(new_n16045_));
  NOR3_X1    g15853(.A1(new_n15991_), .A2(new_n229_), .A3(new_n15981_), .ZN(new_n16046_));
  AOI21_X1   g15854(.A1(new_n16046_), .A2(new_n16045_), .B(new_n15418_), .ZN(new_n16047_));
  AOI21_X1   g15855(.A1(new_n16047_), .A2(new_n15987_), .B(new_n15409_), .ZN(new_n16048_));
  AOI21_X1   g15856(.A1(new_n15992_), .A2(\asqrt[62] ), .B(new_n15410_), .ZN(new_n16049_));
  NOR3_X1    g15857(.A1(new_n16049_), .A2(new_n16021_), .A3(new_n15998_), .ZN(new_n16050_));
  NAND4_X1   g15858(.A1(new_n16050_), .A2(\a[27] ), .A3(new_n16048_), .A4(new_n16001_), .ZN(new_n16051_));
  NAND3_X1   g15859(.A1(new_n16051_), .A2(\a[26] ), .A3(new_n16044_), .ZN(new_n16052_));
  NAND2_X1   g15860(.A1(new_n16043_), .A2(new_n16052_), .ZN(new_n16053_));
  NAND2_X1   g15861(.A1(new_n15433_), .A2(new_n15397_), .ZN(new_n16054_));
  NAND4_X1   g15862(.A1(new_n15437_), .A2(new_n15431_), .A3(new_n15386_), .A4(new_n16054_), .ZN(new_n16055_));
  NOR2_X1    g15863(.A1(new_n15447_), .A2(new_n16034_), .ZN(new_n16056_));
  XOR2_X1    g15864(.A1(new_n16056_), .A2(new_n16055_), .Z(new_n16057_));
  NOR2_X1    g15865(.A1(new_n16057_), .A2(new_n16036_), .ZN(new_n16058_));
  INV_X1     g15866(.I(new_n16058_), .ZN(new_n16059_));
  NAND3_X1   g15867(.A1(new_n16050_), .A2(new_n16048_), .A3(new_n16001_), .ZN(new_n16060_));
  NOR4_X1    g15868(.A1(new_n16020_), .A2(new_n15976_), .A3(new_n15990_), .A4(new_n15981_), .ZN(new_n16061_));
  NOR3_X1    g15869(.A1(new_n16061_), .A2(new_n15418_), .A3(new_n15986_), .ZN(new_n16062_));
  NAND4_X1   g15870(.A1(new_n16017_), .A2(new_n196_), .A3(new_n15410_), .A4(new_n15980_), .ZN(new_n16063_));
  OAI21_X1   g15871(.A1(new_n16062_), .A2(new_n15409_), .B(new_n16063_), .ZN(new_n16064_));
  NAND2_X1   g15872(.A1(new_n16002_), .A2(\asqrt[14] ), .ZN(new_n16065_));
  OAI21_X1   g15873(.A1(new_n16064_), .A2(new_n16065_), .B(new_n15420_), .ZN(new_n16066_));
  NAND3_X1   g15874(.A1(new_n16066_), .A2(new_n15421_), .A3(new_n16060_), .ZN(new_n16067_));
  INV_X1     g15875(.I(new_n16065_), .ZN(new_n16068_));
  AOI21_X1   g15876(.A1(new_n15994_), .A2(new_n16068_), .B(\a[28] ), .ZN(new_n16069_));
  OAI21_X1   g15877(.A1(new_n16069_), .A2(new_n15422_), .B(\asqrt[13] ), .ZN(new_n16070_));
  NAND4_X1   g15878(.A1(new_n16067_), .A2(new_n16070_), .A3(new_n14871_), .A4(new_n16059_), .ZN(new_n16071_));
  NAND2_X1   g15879(.A1(new_n16071_), .A2(new_n16053_), .ZN(new_n16072_));
  NAND3_X1   g15880(.A1(new_n16043_), .A2(new_n16052_), .A3(new_n16059_), .ZN(new_n16073_));
  AOI21_X1   g15881(.A1(\asqrt[14] ), .A2(new_n15420_), .B(\a[29] ), .ZN(new_n16074_));
  NOR2_X1    g15882(.A1(new_n15438_), .A2(\a[28] ), .ZN(new_n16075_));
  AOI21_X1   g15883(.A1(\asqrt[14] ), .A2(\a[28] ), .B(new_n15424_), .ZN(new_n16076_));
  OAI21_X1   g15884(.A1(new_n16075_), .A2(new_n16074_), .B(new_n16076_), .ZN(new_n16077_));
  INV_X1     g15885(.I(new_n16077_), .ZN(new_n16078_));
  NAND3_X1   g15886(.A1(\asqrt[13] ), .A2(new_n15446_), .A3(new_n16078_), .ZN(new_n16079_));
  OAI21_X1   g15887(.A1(new_n16060_), .A2(new_n16077_), .B(new_n15445_), .ZN(new_n16080_));
  NAND3_X1   g15888(.A1(new_n16079_), .A2(new_n16080_), .A3(new_n14273_), .ZN(new_n16081_));
  AOI21_X1   g15889(.A1(new_n16073_), .A2(\asqrt[15] ), .B(new_n16081_), .ZN(new_n16082_));
  NOR2_X1    g15890(.A1(new_n16072_), .A2(new_n16082_), .ZN(new_n16083_));
  AOI22_X1   g15891(.A1(new_n16071_), .A2(new_n16053_), .B1(\asqrt[15] ), .B2(new_n16073_), .ZN(new_n16084_));
  AOI21_X1   g15892(.A1(new_n15456_), .A2(new_n15453_), .B(\asqrt[16] ), .ZN(new_n16085_));
  AND4_X2    g15893(.A1(new_n15497_), .A2(\asqrt[13] ), .A3(new_n15478_), .A4(new_n16085_), .Z(new_n16086_));
  NOR2_X1    g15894(.A1(new_n15497_), .A2(new_n14273_), .ZN(new_n16087_));
  NOR3_X1    g15895(.A1(new_n16086_), .A2(\asqrt[17] ), .A3(new_n16087_), .ZN(new_n16088_));
  OAI21_X1   g15896(.A1(new_n16084_), .A2(new_n14273_), .B(new_n16088_), .ZN(new_n16089_));
  NAND2_X1   g15897(.A1(new_n16089_), .A2(new_n16083_), .ZN(new_n16090_));
  OAI22_X1   g15898(.A1(new_n16084_), .A2(new_n14273_), .B1(new_n16072_), .B2(new_n16082_), .ZN(new_n16091_));
  NAND2_X1   g15899(.A1(new_n15465_), .A2(new_n15466_), .ZN(new_n16092_));
  NAND4_X1   g15900(.A1(\asqrt[13] ), .A2(new_n13760_), .A3(new_n16092_), .A4(new_n15470_), .ZN(new_n16093_));
  XOR2_X1    g15901(.A1(new_n16093_), .A2(new_n15479_), .Z(new_n16094_));
  NAND2_X1   g15902(.A1(new_n16094_), .A2(new_n13192_), .ZN(new_n16095_));
  AOI21_X1   g15903(.A1(new_n16091_), .A2(\asqrt[17] ), .B(new_n16095_), .ZN(new_n16096_));
  NOR2_X1    g15904(.A1(new_n16096_), .A2(new_n16090_), .ZN(new_n16097_));
  AOI22_X1   g15905(.A1(new_n16091_), .A2(\asqrt[17] ), .B1(new_n16089_), .B2(new_n16083_), .ZN(new_n16098_));
  NOR4_X1    g15906(.A1(new_n16060_), .A2(\asqrt[18] ), .A3(new_n15474_), .A4(new_n15823_), .ZN(new_n16099_));
  XOR2_X1    g15907(.A1(new_n16099_), .A2(new_n15480_), .Z(new_n16100_));
  NAND2_X1   g15908(.A1(new_n16100_), .A2(new_n12657_), .ZN(new_n16101_));
  INV_X1     g15909(.I(new_n16101_), .ZN(new_n16102_));
  OAI21_X1   g15910(.A1(new_n16098_), .A2(new_n13192_), .B(new_n16102_), .ZN(new_n16103_));
  NAND2_X1   g15911(.A1(new_n16103_), .A2(new_n16097_), .ZN(new_n16104_));
  OAI22_X1   g15912(.A1(new_n16098_), .A2(new_n13192_), .B1(new_n16096_), .B2(new_n16090_), .ZN(new_n16105_));
  NOR4_X1    g15913(.A1(new_n16060_), .A2(\asqrt[19] ), .A3(new_n15484_), .A4(new_n15506_), .ZN(new_n16106_));
  XNOR2_X1   g15914(.A1(new_n16106_), .A2(new_n15516_), .ZN(new_n16107_));
  NAND2_X1   g15915(.A1(new_n16107_), .A2(new_n12101_), .ZN(new_n16108_));
  AOI21_X1   g15916(.A1(new_n16105_), .A2(\asqrt[19] ), .B(new_n16108_), .ZN(new_n16109_));
  NOR2_X1    g15917(.A1(new_n16109_), .A2(new_n16104_), .ZN(new_n16110_));
  AOI22_X1   g15918(.A1(new_n16105_), .A2(\asqrt[19] ), .B1(new_n16103_), .B2(new_n16097_), .ZN(new_n16111_));
  NOR4_X1    g15919(.A1(new_n16060_), .A2(\asqrt[20] ), .A3(new_n15510_), .A4(new_n15828_), .ZN(new_n16112_));
  XOR2_X1    g15920(.A1(new_n16112_), .A2(new_n15517_), .Z(new_n16113_));
  NAND2_X1   g15921(.A1(new_n16113_), .A2(new_n11631_), .ZN(new_n16114_));
  INV_X1     g15922(.I(new_n16114_), .ZN(new_n16115_));
  OAI21_X1   g15923(.A1(new_n16111_), .A2(new_n12101_), .B(new_n16115_), .ZN(new_n16116_));
  NAND2_X1   g15924(.A1(new_n16116_), .A2(new_n16110_), .ZN(new_n16117_));
  OAI22_X1   g15925(.A1(new_n16111_), .A2(new_n12101_), .B1(new_n16109_), .B2(new_n16104_), .ZN(new_n16118_));
  NOR4_X1    g15926(.A1(new_n16060_), .A2(\asqrt[21] ), .A3(new_n15520_), .A4(new_n15526_), .ZN(new_n16119_));
  XNOR2_X1   g15927(.A1(new_n16119_), .A2(new_n15535_), .ZN(new_n16120_));
  NAND2_X1   g15928(.A1(new_n16120_), .A2(new_n11105_), .ZN(new_n16121_));
  AOI21_X1   g15929(.A1(new_n16118_), .A2(\asqrt[21] ), .B(new_n16121_), .ZN(new_n16122_));
  NOR2_X1    g15930(.A1(new_n16122_), .A2(new_n16117_), .ZN(new_n16123_));
  AOI22_X1   g15931(.A1(new_n16118_), .A2(\asqrt[21] ), .B1(new_n16116_), .B2(new_n16110_), .ZN(new_n16124_));
  NOR4_X1    g15932(.A1(new_n16060_), .A2(\asqrt[22] ), .A3(new_n15529_), .A4(new_n15834_), .ZN(new_n16125_));
  XOR2_X1    g15933(.A1(new_n16125_), .A2(new_n15536_), .Z(new_n16126_));
  NAND2_X1   g15934(.A1(new_n16126_), .A2(new_n10614_), .ZN(new_n16127_));
  INV_X1     g15935(.I(new_n16127_), .ZN(new_n16128_));
  OAI21_X1   g15936(.A1(new_n16124_), .A2(new_n11105_), .B(new_n16128_), .ZN(new_n16129_));
  NAND2_X1   g15937(.A1(new_n16129_), .A2(new_n16123_), .ZN(new_n16130_));
  OAI22_X1   g15938(.A1(new_n16124_), .A2(new_n11105_), .B1(new_n16122_), .B2(new_n16117_), .ZN(new_n16131_));
  NAND2_X1   g15939(.A1(new_n15545_), .A2(\asqrt[23] ), .ZN(new_n16132_));
  NOR4_X1    g15940(.A1(new_n16060_), .A2(\asqrt[23] ), .A3(new_n15539_), .A4(new_n15545_), .ZN(new_n16133_));
  XOR2_X1    g15941(.A1(new_n16133_), .A2(new_n16132_), .Z(new_n16134_));
  NAND2_X1   g15942(.A1(new_n16134_), .A2(new_n10104_), .ZN(new_n16135_));
  AOI21_X1   g15943(.A1(new_n16131_), .A2(\asqrt[23] ), .B(new_n16135_), .ZN(new_n16136_));
  NOR2_X1    g15944(.A1(new_n16136_), .A2(new_n16130_), .ZN(new_n16137_));
  AOI22_X1   g15945(.A1(new_n16131_), .A2(\asqrt[23] ), .B1(new_n16129_), .B2(new_n16123_), .ZN(new_n16138_));
  NOR4_X1    g15946(.A1(new_n16060_), .A2(\asqrt[24] ), .A3(new_n15548_), .A4(new_n15841_), .ZN(new_n16139_));
  AOI21_X1   g15947(.A1(new_n16132_), .A2(new_n15543_), .B(new_n10104_), .ZN(new_n16140_));
  NOR2_X1    g15948(.A1(new_n16139_), .A2(new_n16140_), .ZN(new_n16141_));
  NAND2_X1   g15949(.A1(new_n16141_), .A2(new_n9672_), .ZN(new_n16142_));
  INV_X1     g15950(.I(new_n16142_), .ZN(new_n16143_));
  OAI21_X1   g15951(.A1(new_n16138_), .A2(new_n10104_), .B(new_n16143_), .ZN(new_n16144_));
  NAND2_X1   g15952(.A1(new_n16144_), .A2(new_n16137_), .ZN(new_n16145_));
  OAI22_X1   g15953(.A1(new_n16138_), .A2(new_n10104_), .B1(new_n16136_), .B2(new_n16130_), .ZN(new_n16146_));
  NAND2_X1   g15954(.A1(new_n15560_), .A2(\asqrt[25] ), .ZN(new_n16147_));
  NOR4_X1    g15955(.A1(new_n16060_), .A2(\asqrt[25] ), .A3(new_n15555_), .A4(new_n15560_), .ZN(new_n16148_));
  XOR2_X1    g15956(.A1(new_n16148_), .A2(new_n16147_), .Z(new_n16149_));
  NAND2_X1   g15957(.A1(new_n16149_), .A2(new_n9212_), .ZN(new_n16150_));
  AOI21_X1   g15958(.A1(new_n16146_), .A2(\asqrt[25] ), .B(new_n16150_), .ZN(new_n16151_));
  NOR2_X1    g15959(.A1(new_n16151_), .A2(new_n16145_), .ZN(new_n16152_));
  AOI22_X1   g15960(.A1(new_n16146_), .A2(\asqrt[25] ), .B1(new_n16144_), .B2(new_n16137_), .ZN(new_n16153_));
  NOR4_X1    g15961(.A1(new_n16060_), .A2(\asqrt[26] ), .A3(new_n15563_), .A4(new_n15848_), .ZN(new_n16154_));
  AOI21_X1   g15962(.A1(new_n16147_), .A2(new_n15559_), .B(new_n9212_), .ZN(new_n16155_));
  NOR2_X1    g15963(.A1(new_n16154_), .A2(new_n16155_), .ZN(new_n16156_));
  NAND2_X1   g15964(.A1(new_n16156_), .A2(new_n8763_), .ZN(new_n16157_));
  INV_X1     g15965(.I(new_n16157_), .ZN(new_n16158_));
  OAI21_X1   g15966(.A1(new_n16153_), .A2(new_n9212_), .B(new_n16158_), .ZN(new_n16159_));
  NAND2_X1   g15967(.A1(new_n16159_), .A2(new_n16152_), .ZN(new_n16160_));
  OAI22_X1   g15968(.A1(new_n16153_), .A2(new_n9212_), .B1(new_n16151_), .B2(new_n16145_), .ZN(new_n16161_));
  NAND2_X1   g15969(.A1(new_n15575_), .A2(\asqrt[27] ), .ZN(new_n16162_));
  NOR4_X1    g15970(.A1(new_n16060_), .A2(\asqrt[27] ), .A3(new_n15570_), .A4(new_n15575_), .ZN(new_n16163_));
  XOR2_X1    g15971(.A1(new_n16163_), .A2(new_n16162_), .Z(new_n16164_));
  NAND2_X1   g15972(.A1(new_n16164_), .A2(new_n8319_), .ZN(new_n16165_));
  AOI21_X1   g15973(.A1(new_n16161_), .A2(\asqrt[27] ), .B(new_n16165_), .ZN(new_n16166_));
  NOR2_X1    g15974(.A1(new_n16166_), .A2(new_n16160_), .ZN(new_n16167_));
  AOI22_X1   g15975(.A1(new_n16161_), .A2(\asqrt[27] ), .B1(new_n16159_), .B2(new_n16152_), .ZN(new_n16168_));
  NOR4_X1    g15976(.A1(new_n16060_), .A2(\asqrt[28] ), .A3(new_n15578_), .A4(new_n15855_), .ZN(new_n16169_));
  AOI21_X1   g15977(.A1(new_n16162_), .A2(new_n15574_), .B(new_n8319_), .ZN(new_n16170_));
  NOR2_X1    g15978(.A1(new_n16169_), .A2(new_n16170_), .ZN(new_n16171_));
  NAND2_X1   g15979(.A1(new_n16171_), .A2(new_n7931_), .ZN(new_n16172_));
  INV_X1     g15980(.I(new_n16172_), .ZN(new_n16173_));
  OAI21_X1   g15981(.A1(new_n16168_), .A2(new_n8319_), .B(new_n16173_), .ZN(new_n16174_));
  NAND2_X1   g15982(.A1(new_n16174_), .A2(new_n16167_), .ZN(new_n16175_));
  OAI22_X1   g15983(.A1(new_n16168_), .A2(new_n8319_), .B1(new_n16166_), .B2(new_n16160_), .ZN(new_n16176_));
  NAND2_X1   g15984(.A1(new_n15590_), .A2(\asqrt[29] ), .ZN(new_n16177_));
  NOR4_X1    g15985(.A1(new_n16060_), .A2(\asqrt[29] ), .A3(new_n15585_), .A4(new_n15590_), .ZN(new_n16178_));
  XOR2_X1    g15986(.A1(new_n16178_), .A2(new_n16177_), .Z(new_n16179_));
  NAND2_X1   g15987(.A1(new_n16179_), .A2(new_n7517_), .ZN(new_n16180_));
  AOI21_X1   g15988(.A1(new_n16176_), .A2(\asqrt[29] ), .B(new_n16180_), .ZN(new_n16181_));
  NOR2_X1    g15989(.A1(new_n16181_), .A2(new_n16175_), .ZN(new_n16182_));
  AOI22_X1   g15990(.A1(new_n16176_), .A2(\asqrt[29] ), .B1(new_n16174_), .B2(new_n16167_), .ZN(new_n16183_));
  NOR4_X1    g15991(.A1(new_n16060_), .A2(\asqrt[30] ), .A3(new_n15593_), .A4(new_n15862_), .ZN(new_n16184_));
  AOI21_X1   g15992(.A1(new_n16177_), .A2(new_n15589_), .B(new_n7517_), .ZN(new_n16185_));
  NOR2_X1    g15993(.A1(new_n16184_), .A2(new_n16185_), .ZN(new_n16186_));
  NAND2_X1   g15994(.A1(new_n16186_), .A2(new_n7110_), .ZN(new_n16187_));
  INV_X1     g15995(.I(new_n16187_), .ZN(new_n16188_));
  OAI21_X1   g15996(.A1(new_n16183_), .A2(new_n7517_), .B(new_n16188_), .ZN(new_n16189_));
  NAND2_X1   g15997(.A1(new_n16189_), .A2(new_n16182_), .ZN(new_n16190_));
  OAI22_X1   g15998(.A1(new_n16183_), .A2(new_n7517_), .B1(new_n16181_), .B2(new_n16175_), .ZN(new_n16191_));
  NAND2_X1   g15999(.A1(new_n15605_), .A2(\asqrt[31] ), .ZN(new_n16192_));
  NOR4_X1    g16000(.A1(new_n16060_), .A2(\asqrt[31] ), .A3(new_n15600_), .A4(new_n15605_), .ZN(new_n16193_));
  XOR2_X1    g16001(.A1(new_n16193_), .A2(new_n16192_), .Z(new_n16194_));
  NAND2_X1   g16002(.A1(new_n16194_), .A2(new_n6708_), .ZN(new_n16195_));
  AOI21_X1   g16003(.A1(new_n16191_), .A2(\asqrt[31] ), .B(new_n16195_), .ZN(new_n16196_));
  NOR2_X1    g16004(.A1(new_n16196_), .A2(new_n16190_), .ZN(new_n16197_));
  AOI22_X1   g16005(.A1(new_n16191_), .A2(\asqrt[31] ), .B1(new_n16189_), .B2(new_n16182_), .ZN(new_n16198_));
  NOR4_X1    g16006(.A1(new_n16060_), .A2(\asqrt[32] ), .A3(new_n15608_), .A4(new_n15869_), .ZN(new_n16199_));
  AOI21_X1   g16007(.A1(new_n16192_), .A2(new_n15604_), .B(new_n6708_), .ZN(new_n16200_));
  NOR2_X1    g16008(.A1(new_n16199_), .A2(new_n16200_), .ZN(new_n16201_));
  NAND2_X1   g16009(.A1(new_n16201_), .A2(new_n6365_), .ZN(new_n16202_));
  INV_X1     g16010(.I(new_n16202_), .ZN(new_n16203_));
  OAI21_X1   g16011(.A1(new_n16198_), .A2(new_n6708_), .B(new_n16203_), .ZN(new_n16204_));
  NAND2_X1   g16012(.A1(new_n16204_), .A2(new_n16197_), .ZN(new_n16205_));
  OAI22_X1   g16013(.A1(new_n16198_), .A2(new_n6708_), .B1(new_n16196_), .B2(new_n16190_), .ZN(new_n16206_));
  NAND2_X1   g16014(.A1(new_n15620_), .A2(\asqrt[33] ), .ZN(new_n16207_));
  NOR4_X1    g16015(.A1(new_n16060_), .A2(\asqrt[33] ), .A3(new_n15615_), .A4(new_n15620_), .ZN(new_n16208_));
  XOR2_X1    g16016(.A1(new_n16208_), .A2(new_n16207_), .Z(new_n16209_));
  NAND2_X1   g16017(.A1(new_n16209_), .A2(new_n5991_), .ZN(new_n16210_));
  AOI21_X1   g16018(.A1(new_n16206_), .A2(\asqrt[33] ), .B(new_n16210_), .ZN(new_n16211_));
  NOR2_X1    g16019(.A1(new_n16211_), .A2(new_n16205_), .ZN(new_n16212_));
  AOI22_X1   g16020(.A1(new_n16206_), .A2(\asqrt[33] ), .B1(new_n16204_), .B2(new_n16197_), .ZN(new_n16213_));
  NAND2_X1   g16021(.A1(new_n15876_), .A2(\asqrt[34] ), .ZN(new_n16214_));
  NOR4_X1    g16022(.A1(new_n16060_), .A2(\asqrt[34] ), .A3(new_n15623_), .A4(new_n15876_), .ZN(new_n16215_));
  XOR2_X1    g16023(.A1(new_n16215_), .A2(new_n16214_), .Z(new_n16216_));
  NAND2_X1   g16024(.A1(new_n16216_), .A2(new_n5626_), .ZN(new_n16217_));
  INV_X1     g16025(.I(new_n16217_), .ZN(new_n16218_));
  OAI21_X1   g16026(.A1(new_n16213_), .A2(new_n5991_), .B(new_n16218_), .ZN(new_n16219_));
  NAND2_X1   g16027(.A1(new_n16219_), .A2(new_n16212_), .ZN(new_n16220_));
  OAI22_X1   g16028(.A1(new_n16213_), .A2(new_n5991_), .B1(new_n16211_), .B2(new_n16205_), .ZN(new_n16221_));
  NOR4_X1    g16029(.A1(new_n16060_), .A2(\asqrt[35] ), .A3(new_n15630_), .A4(new_n15635_), .ZN(new_n16222_));
  AOI21_X1   g16030(.A1(new_n16214_), .A2(new_n15875_), .B(new_n5626_), .ZN(new_n16223_));
  NOR2_X1    g16031(.A1(new_n16222_), .A2(new_n16223_), .ZN(new_n16224_));
  NAND2_X1   g16032(.A1(new_n16224_), .A2(new_n5273_), .ZN(new_n16225_));
  AOI21_X1   g16033(.A1(new_n16221_), .A2(\asqrt[35] ), .B(new_n16225_), .ZN(new_n16226_));
  NOR2_X1    g16034(.A1(new_n16226_), .A2(new_n16220_), .ZN(new_n16227_));
  AOI22_X1   g16035(.A1(new_n16221_), .A2(\asqrt[35] ), .B1(new_n16219_), .B2(new_n16212_), .ZN(new_n16228_));
  NAND2_X1   g16036(.A1(new_n15883_), .A2(\asqrt[36] ), .ZN(new_n16229_));
  NOR4_X1    g16037(.A1(new_n16060_), .A2(\asqrt[36] ), .A3(new_n15638_), .A4(new_n15883_), .ZN(new_n16230_));
  XOR2_X1    g16038(.A1(new_n16230_), .A2(new_n16229_), .Z(new_n16231_));
  NAND2_X1   g16039(.A1(new_n16231_), .A2(new_n4973_), .ZN(new_n16232_));
  INV_X1     g16040(.I(new_n16232_), .ZN(new_n16233_));
  OAI21_X1   g16041(.A1(new_n16228_), .A2(new_n5273_), .B(new_n16233_), .ZN(new_n16234_));
  NAND2_X1   g16042(.A1(new_n16234_), .A2(new_n16227_), .ZN(new_n16235_));
  OAI22_X1   g16043(.A1(new_n16228_), .A2(new_n5273_), .B1(new_n16226_), .B2(new_n16220_), .ZN(new_n16236_));
  NOR4_X1    g16044(.A1(new_n16060_), .A2(\asqrt[37] ), .A3(new_n15645_), .A4(new_n15650_), .ZN(new_n16237_));
  AOI21_X1   g16045(.A1(new_n16229_), .A2(new_n15882_), .B(new_n4973_), .ZN(new_n16238_));
  NOR2_X1    g16046(.A1(new_n16237_), .A2(new_n16238_), .ZN(new_n16239_));
  NAND2_X1   g16047(.A1(new_n16239_), .A2(new_n4645_), .ZN(new_n16240_));
  AOI21_X1   g16048(.A1(new_n16236_), .A2(\asqrt[37] ), .B(new_n16240_), .ZN(new_n16241_));
  NOR2_X1    g16049(.A1(new_n16241_), .A2(new_n16235_), .ZN(new_n16242_));
  AOI22_X1   g16050(.A1(new_n16236_), .A2(\asqrt[37] ), .B1(new_n16234_), .B2(new_n16227_), .ZN(new_n16243_));
  NAND2_X1   g16051(.A1(new_n15890_), .A2(\asqrt[38] ), .ZN(new_n16244_));
  NOR4_X1    g16052(.A1(new_n16060_), .A2(\asqrt[38] ), .A3(new_n15653_), .A4(new_n15890_), .ZN(new_n16245_));
  XOR2_X1    g16053(.A1(new_n16245_), .A2(new_n16244_), .Z(new_n16246_));
  NAND2_X1   g16054(.A1(new_n16246_), .A2(new_n4330_), .ZN(new_n16247_));
  INV_X1     g16055(.I(new_n16247_), .ZN(new_n16248_));
  OAI21_X1   g16056(.A1(new_n16243_), .A2(new_n4645_), .B(new_n16248_), .ZN(new_n16249_));
  NAND2_X1   g16057(.A1(new_n16249_), .A2(new_n16242_), .ZN(new_n16250_));
  OAI22_X1   g16058(.A1(new_n16243_), .A2(new_n4645_), .B1(new_n16241_), .B2(new_n16235_), .ZN(new_n16251_));
  NAND2_X1   g16059(.A1(new_n15665_), .A2(\asqrt[39] ), .ZN(new_n16252_));
  NOR4_X1    g16060(.A1(new_n16060_), .A2(\asqrt[39] ), .A3(new_n15660_), .A4(new_n15665_), .ZN(new_n16253_));
  XOR2_X1    g16061(.A1(new_n16253_), .A2(new_n16252_), .Z(new_n16254_));
  NAND2_X1   g16062(.A1(new_n16254_), .A2(new_n4018_), .ZN(new_n16255_));
  AOI21_X1   g16063(.A1(new_n16251_), .A2(\asqrt[39] ), .B(new_n16255_), .ZN(new_n16256_));
  NOR2_X1    g16064(.A1(new_n16256_), .A2(new_n16250_), .ZN(new_n16257_));
  AOI22_X1   g16065(.A1(new_n16251_), .A2(\asqrt[39] ), .B1(new_n16249_), .B2(new_n16242_), .ZN(new_n16258_));
  NOR4_X1    g16066(.A1(new_n16060_), .A2(\asqrt[40] ), .A3(new_n15668_), .A4(new_n15897_), .ZN(new_n16259_));
  AOI21_X1   g16067(.A1(new_n16252_), .A2(new_n15664_), .B(new_n4018_), .ZN(new_n16260_));
  NOR2_X1    g16068(.A1(new_n16259_), .A2(new_n16260_), .ZN(new_n16261_));
  NAND2_X1   g16069(.A1(new_n16261_), .A2(new_n3760_), .ZN(new_n16262_));
  INV_X1     g16070(.I(new_n16262_), .ZN(new_n16263_));
  OAI21_X1   g16071(.A1(new_n16258_), .A2(new_n4018_), .B(new_n16263_), .ZN(new_n16264_));
  NAND2_X1   g16072(.A1(new_n16264_), .A2(new_n16257_), .ZN(new_n16265_));
  OAI22_X1   g16073(.A1(new_n16258_), .A2(new_n4018_), .B1(new_n16256_), .B2(new_n16250_), .ZN(new_n16266_));
  NAND2_X1   g16074(.A1(new_n15680_), .A2(\asqrt[41] ), .ZN(new_n16267_));
  NOR4_X1    g16075(.A1(new_n16060_), .A2(\asqrt[41] ), .A3(new_n15675_), .A4(new_n15680_), .ZN(new_n16268_));
  XOR2_X1    g16076(.A1(new_n16268_), .A2(new_n16267_), .Z(new_n16269_));
  NAND2_X1   g16077(.A1(new_n16269_), .A2(new_n3481_), .ZN(new_n16270_));
  AOI21_X1   g16078(.A1(new_n16266_), .A2(\asqrt[41] ), .B(new_n16270_), .ZN(new_n16271_));
  NOR2_X1    g16079(.A1(new_n16271_), .A2(new_n16265_), .ZN(new_n16272_));
  AOI22_X1   g16080(.A1(new_n16266_), .A2(\asqrt[41] ), .B1(new_n16264_), .B2(new_n16257_), .ZN(new_n16273_));
  NOR4_X1    g16081(.A1(new_n16060_), .A2(\asqrt[42] ), .A3(new_n15683_), .A4(new_n15904_), .ZN(new_n16274_));
  AOI21_X1   g16082(.A1(new_n16267_), .A2(new_n15679_), .B(new_n3481_), .ZN(new_n16275_));
  NOR2_X1    g16083(.A1(new_n16274_), .A2(new_n16275_), .ZN(new_n16276_));
  NAND2_X1   g16084(.A1(new_n16276_), .A2(new_n3208_), .ZN(new_n16277_));
  INV_X1     g16085(.I(new_n16277_), .ZN(new_n16278_));
  OAI21_X1   g16086(.A1(new_n16273_), .A2(new_n3481_), .B(new_n16278_), .ZN(new_n16279_));
  NAND2_X1   g16087(.A1(new_n16279_), .A2(new_n16272_), .ZN(new_n16280_));
  OAI22_X1   g16088(.A1(new_n16273_), .A2(new_n3481_), .B1(new_n16271_), .B2(new_n16265_), .ZN(new_n16281_));
  NAND2_X1   g16089(.A1(new_n15695_), .A2(\asqrt[43] ), .ZN(new_n16282_));
  NOR4_X1    g16090(.A1(new_n16060_), .A2(\asqrt[43] ), .A3(new_n15690_), .A4(new_n15695_), .ZN(new_n16283_));
  XOR2_X1    g16091(.A1(new_n16283_), .A2(new_n16282_), .Z(new_n16284_));
  NAND2_X1   g16092(.A1(new_n16284_), .A2(new_n2941_), .ZN(new_n16285_));
  AOI21_X1   g16093(.A1(new_n16281_), .A2(\asqrt[43] ), .B(new_n16285_), .ZN(new_n16286_));
  NOR2_X1    g16094(.A1(new_n16286_), .A2(new_n16280_), .ZN(new_n16287_));
  AOI22_X1   g16095(.A1(new_n16281_), .A2(\asqrt[43] ), .B1(new_n16279_), .B2(new_n16272_), .ZN(new_n16288_));
  NOR4_X1    g16096(.A1(new_n16060_), .A2(\asqrt[44] ), .A3(new_n15698_), .A4(new_n15911_), .ZN(new_n16289_));
  AOI21_X1   g16097(.A1(new_n16282_), .A2(new_n15694_), .B(new_n2941_), .ZN(new_n16290_));
  NOR2_X1    g16098(.A1(new_n16289_), .A2(new_n16290_), .ZN(new_n16291_));
  NAND2_X1   g16099(.A1(new_n16291_), .A2(new_n2728_), .ZN(new_n16292_));
  INV_X1     g16100(.I(new_n16292_), .ZN(new_n16293_));
  OAI21_X1   g16101(.A1(new_n16288_), .A2(new_n2941_), .B(new_n16293_), .ZN(new_n16294_));
  NAND2_X1   g16102(.A1(new_n16294_), .A2(new_n16287_), .ZN(new_n16295_));
  OAI22_X1   g16103(.A1(new_n16288_), .A2(new_n2941_), .B1(new_n16286_), .B2(new_n16280_), .ZN(new_n16296_));
  NAND2_X1   g16104(.A1(new_n15710_), .A2(\asqrt[45] ), .ZN(new_n16297_));
  NOR4_X1    g16105(.A1(new_n16060_), .A2(\asqrt[45] ), .A3(new_n15705_), .A4(new_n15710_), .ZN(new_n16298_));
  XOR2_X1    g16106(.A1(new_n16298_), .A2(new_n16297_), .Z(new_n16299_));
  NAND2_X1   g16107(.A1(new_n16299_), .A2(new_n2488_), .ZN(new_n16300_));
  AOI21_X1   g16108(.A1(new_n16296_), .A2(\asqrt[45] ), .B(new_n16300_), .ZN(new_n16301_));
  NOR2_X1    g16109(.A1(new_n16301_), .A2(new_n16295_), .ZN(new_n16302_));
  AOI22_X1   g16110(.A1(new_n16296_), .A2(\asqrt[45] ), .B1(new_n16294_), .B2(new_n16287_), .ZN(new_n16303_));
  NAND2_X1   g16111(.A1(new_n15918_), .A2(\asqrt[46] ), .ZN(new_n16304_));
  NOR4_X1    g16112(.A1(new_n16060_), .A2(\asqrt[46] ), .A3(new_n15713_), .A4(new_n15918_), .ZN(new_n16305_));
  XOR2_X1    g16113(.A1(new_n16305_), .A2(new_n16304_), .Z(new_n16306_));
  NAND2_X1   g16114(.A1(new_n16306_), .A2(new_n2253_), .ZN(new_n16307_));
  INV_X1     g16115(.I(new_n16307_), .ZN(new_n16308_));
  OAI21_X1   g16116(.A1(new_n16303_), .A2(new_n2488_), .B(new_n16308_), .ZN(new_n16309_));
  NAND2_X1   g16117(.A1(new_n16309_), .A2(new_n16302_), .ZN(new_n16310_));
  OAI22_X1   g16118(.A1(new_n16303_), .A2(new_n2488_), .B1(new_n16301_), .B2(new_n16295_), .ZN(new_n16311_));
  NOR4_X1    g16119(.A1(new_n16060_), .A2(\asqrt[47] ), .A3(new_n15720_), .A4(new_n15725_), .ZN(new_n16312_));
  AOI21_X1   g16120(.A1(new_n16304_), .A2(new_n15917_), .B(new_n2253_), .ZN(new_n16313_));
  NOR2_X1    g16121(.A1(new_n16312_), .A2(new_n16313_), .ZN(new_n16314_));
  NAND2_X1   g16122(.A1(new_n16314_), .A2(new_n2046_), .ZN(new_n16315_));
  AOI21_X1   g16123(.A1(new_n16311_), .A2(\asqrt[47] ), .B(new_n16315_), .ZN(new_n16316_));
  NOR2_X1    g16124(.A1(new_n16316_), .A2(new_n16310_), .ZN(new_n16317_));
  AOI22_X1   g16125(.A1(new_n16311_), .A2(\asqrt[47] ), .B1(new_n16309_), .B2(new_n16302_), .ZN(new_n16318_));
  NAND2_X1   g16126(.A1(new_n15925_), .A2(\asqrt[48] ), .ZN(new_n16319_));
  NOR4_X1    g16127(.A1(new_n16060_), .A2(\asqrt[48] ), .A3(new_n15728_), .A4(new_n15925_), .ZN(new_n16320_));
  XOR2_X1    g16128(.A1(new_n16320_), .A2(new_n16319_), .Z(new_n16321_));
  NAND2_X1   g16129(.A1(new_n16321_), .A2(new_n1854_), .ZN(new_n16322_));
  INV_X1     g16130(.I(new_n16322_), .ZN(new_n16323_));
  OAI21_X1   g16131(.A1(new_n16318_), .A2(new_n2046_), .B(new_n16323_), .ZN(new_n16324_));
  NAND2_X1   g16132(.A1(new_n16324_), .A2(new_n16317_), .ZN(new_n16325_));
  OAI22_X1   g16133(.A1(new_n16318_), .A2(new_n2046_), .B1(new_n16316_), .B2(new_n16310_), .ZN(new_n16326_));
  NOR4_X1    g16134(.A1(new_n16060_), .A2(\asqrt[49] ), .A3(new_n15735_), .A4(new_n15740_), .ZN(new_n16327_));
  AOI21_X1   g16135(.A1(new_n16319_), .A2(new_n15924_), .B(new_n1854_), .ZN(new_n16328_));
  NOR2_X1    g16136(.A1(new_n16327_), .A2(new_n16328_), .ZN(new_n16329_));
  NAND2_X1   g16137(.A1(new_n16329_), .A2(new_n1595_), .ZN(new_n16330_));
  AOI21_X1   g16138(.A1(new_n16326_), .A2(\asqrt[49] ), .B(new_n16330_), .ZN(new_n16331_));
  NOR2_X1    g16139(.A1(new_n16331_), .A2(new_n16325_), .ZN(new_n16332_));
  AOI22_X1   g16140(.A1(new_n16326_), .A2(\asqrt[49] ), .B1(new_n16324_), .B2(new_n16317_), .ZN(new_n16333_));
  NAND2_X1   g16141(.A1(new_n15932_), .A2(\asqrt[50] ), .ZN(new_n16334_));
  NOR4_X1    g16142(.A1(new_n16060_), .A2(\asqrt[50] ), .A3(new_n15743_), .A4(new_n15932_), .ZN(new_n16335_));
  XOR2_X1    g16143(.A1(new_n16335_), .A2(new_n16334_), .Z(new_n16336_));
  NAND2_X1   g16144(.A1(new_n16336_), .A2(new_n1436_), .ZN(new_n16337_));
  INV_X1     g16145(.I(new_n16337_), .ZN(new_n16338_));
  OAI21_X1   g16146(.A1(new_n16333_), .A2(new_n1595_), .B(new_n16338_), .ZN(new_n16339_));
  NAND2_X1   g16147(.A1(new_n16339_), .A2(new_n16332_), .ZN(new_n16340_));
  OAI22_X1   g16148(.A1(new_n16333_), .A2(new_n1595_), .B1(new_n16331_), .B2(new_n16325_), .ZN(new_n16341_));
  NAND2_X1   g16149(.A1(new_n15755_), .A2(\asqrt[51] ), .ZN(new_n16342_));
  NOR4_X1    g16150(.A1(new_n16060_), .A2(\asqrt[51] ), .A3(new_n15750_), .A4(new_n15755_), .ZN(new_n16343_));
  XOR2_X1    g16151(.A1(new_n16343_), .A2(new_n16342_), .Z(new_n16344_));
  NAND2_X1   g16152(.A1(new_n16344_), .A2(new_n1260_), .ZN(new_n16345_));
  AOI21_X1   g16153(.A1(new_n16341_), .A2(\asqrt[51] ), .B(new_n16345_), .ZN(new_n16346_));
  NOR2_X1    g16154(.A1(new_n16346_), .A2(new_n16340_), .ZN(new_n16347_));
  AOI22_X1   g16155(.A1(new_n16341_), .A2(\asqrt[51] ), .B1(new_n16339_), .B2(new_n16332_), .ZN(new_n16348_));
  NOR4_X1    g16156(.A1(new_n16060_), .A2(\asqrt[52] ), .A3(new_n15758_), .A4(new_n15939_), .ZN(new_n16349_));
  AOI21_X1   g16157(.A1(new_n16342_), .A2(new_n15754_), .B(new_n1260_), .ZN(new_n16350_));
  NOR2_X1    g16158(.A1(new_n16349_), .A2(new_n16350_), .ZN(new_n16351_));
  NAND2_X1   g16159(.A1(new_n16351_), .A2(new_n1096_), .ZN(new_n16352_));
  INV_X1     g16160(.I(new_n16352_), .ZN(new_n16353_));
  OAI21_X1   g16161(.A1(new_n16348_), .A2(new_n1260_), .B(new_n16353_), .ZN(new_n16354_));
  NAND2_X1   g16162(.A1(new_n16354_), .A2(new_n16347_), .ZN(new_n16355_));
  OAI22_X1   g16163(.A1(new_n16348_), .A2(new_n1260_), .B1(new_n16346_), .B2(new_n16340_), .ZN(new_n16356_));
  NOR2_X1    g16164(.A1(new_n15942_), .A2(new_n1096_), .ZN(new_n16357_));
  NOR4_X1    g16165(.A1(new_n16060_), .A2(\asqrt[53] ), .A3(new_n15765_), .A4(new_n15770_), .ZN(new_n16358_));
  XNOR2_X1   g16166(.A1(new_n16358_), .A2(new_n16357_), .ZN(new_n16359_));
  NAND2_X1   g16167(.A1(new_n16359_), .A2(new_n970_), .ZN(new_n16360_));
  AOI21_X1   g16168(.A1(new_n16356_), .A2(\asqrt[53] ), .B(new_n16360_), .ZN(new_n16361_));
  NOR2_X1    g16169(.A1(new_n16361_), .A2(new_n16355_), .ZN(new_n16362_));
  AOI22_X1   g16170(.A1(new_n16356_), .A2(\asqrt[53] ), .B1(new_n16354_), .B2(new_n16347_), .ZN(new_n16363_));
  NOR4_X1    g16171(.A1(new_n16060_), .A2(\asqrt[54] ), .A3(new_n15773_), .A4(new_n15946_), .ZN(new_n16364_));
  XOR2_X1    g16172(.A1(new_n16364_), .A2(new_n15959_), .Z(new_n16365_));
  NAND2_X1   g16173(.A1(new_n16365_), .A2(new_n825_), .ZN(new_n16366_));
  INV_X1     g16174(.I(new_n16366_), .ZN(new_n16367_));
  OAI21_X1   g16175(.A1(new_n16363_), .A2(new_n970_), .B(new_n16367_), .ZN(new_n16368_));
  NAND2_X1   g16176(.A1(new_n16368_), .A2(new_n16362_), .ZN(new_n16369_));
  OAI22_X1   g16177(.A1(new_n16363_), .A2(new_n970_), .B1(new_n16361_), .B2(new_n16355_), .ZN(new_n16370_));
  NOR4_X1    g16178(.A1(new_n16060_), .A2(\asqrt[55] ), .A3(new_n15780_), .A4(new_n15785_), .ZN(new_n16371_));
  XOR2_X1    g16179(.A1(new_n16371_), .A2(new_n15800_), .Z(new_n16372_));
  NAND2_X1   g16180(.A1(new_n16372_), .A2(new_n724_), .ZN(new_n16373_));
  AOI21_X1   g16181(.A1(new_n16370_), .A2(\asqrt[55] ), .B(new_n16373_), .ZN(new_n16374_));
  NOR2_X1    g16182(.A1(new_n16374_), .A2(new_n16369_), .ZN(new_n16375_));
  AOI22_X1   g16183(.A1(new_n16370_), .A2(\asqrt[55] ), .B1(new_n16368_), .B2(new_n16362_), .ZN(new_n16376_));
  NOR4_X1    g16184(.A1(new_n16060_), .A2(\asqrt[56] ), .A3(new_n15788_), .A4(new_n15953_), .ZN(new_n16377_));
  XOR2_X1    g16185(.A1(new_n16377_), .A2(new_n15961_), .Z(new_n16378_));
  NAND2_X1   g16186(.A1(new_n16378_), .A2(new_n587_), .ZN(new_n16379_));
  INV_X1     g16187(.I(new_n16379_), .ZN(new_n16380_));
  OAI21_X1   g16188(.A1(new_n16376_), .A2(new_n724_), .B(new_n16380_), .ZN(new_n16381_));
  NAND2_X1   g16189(.A1(new_n16381_), .A2(new_n16375_), .ZN(new_n16382_));
  OAI22_X1   g16190(.A1(new_n16376_), .A2(new_n724_), .B1(new_n16374_), .B2(new_n16369_), .ZN(new_n16383_));
  NOR4_X1    g16191(.A1(new_n16060_), .A2(\asqrt[57] ), .A3(new_n15795_), .A4(new_n15809_), .ZN(new_n16384_));
  XOR2_X1    g16192(.A1(new_n16384_), .A2(new_n15802_), .Z(new_n16385_));
  NAND2_X1   g16193(.A1(new_n16385_), .A2(new_n504_), .ZN(new_n16386_));
  AOI21_X1   g16194(.A1(new_n16383_), .A2(\asqrt[57] ), .B(new_n16386_), .ZN(new_n16387_));
  NOR2_X1    g16195(.A1(new_n16387_), .A2(new_n16382_), .ZN(new_n16388_));
  AOI22_X1   g16196(.A1(new_n16383_), .A2(\asqrt[57] ), .B1(new_n16381_), .B2(new_n16375_), .ZN(new_n16389_));
  NOR4_X1    g16197(.A1(new_n16060_), .A2(\asqrt[58] ), .A3(new_n15805_), .A4(new_n15971_), .ZN(new_n16390_));
  XOR2_X1    g16198(.A1(new_n16390_), .A2(new_n15963_), .Z(new_n16391_));
  NAND2_X1   g16199(.A1(new_n16391_), .A2(new_n376_), .ZN(new_n16392_));
  INV_X1     g16200(.I(new_n16392_), .ZN(new_n16393_));
  OAI21_X1   g16201(.A1(new_n16389_), .A2(new_n504_), .B(new_n16393_), .ZN(new_n16394_));
  NAND2_X1   g16202(.A1(new_n16394_), .A2(new_n16388_), .ZN(new_n16395_));
  OAI22_X1   g16203(.A1(new_n16389_), .A2(new_n504_), .B1(new_n16387_), .B2(new_n16382_), .ZN(new_n16396_));
  NOR4_X1    g16204(.A1(new_n16060_), .A2(\asqrt[59] ), .A3(new_n15812_), .A4(new_n15964_), .ZN(new_n16397_));
  XOR2_X1    g16205(.A1(new_n16397_), .A2(new_n15818_), .Z(new_n16398_));
  NAND2_X1   g16206(.A1(new_n16398_), .A2(new_n275_), .ZN(new_n16399_));
  AOI21_X1   g16207(.A1(new_n16396_), .A2(\asqrt[59] ), .B(new_n16399_), .ZN(new_n16400_));
  NOR2_X1    g16208(.A1(new_n16400_), .A2(new_n16395_), .ZN(new_n16401_));
  AOI22_X1   g16209(.A1(new_n16396_), .A2(\asqrt[59] ), .B1(new_n16394_), .B2(new_n16388_), .ZN(new_n16402_));
  NOR4_X1    g16210(.A1(new_n16060_), .A2(\asqrt[60] ), .A3(new_n15820_), .A4(new_n15989_), .ZN(new_n16403_));
  XOR2_X1    g16211(.A1(new_n16403_), .A2(new_n15978_), .Z(new_n16404_));
  NAND2_X1   g16212(.A1(new_n16404_), .A2(new_n229_), .ZN(new_n16405_));
  INV_X1     g16213(.I(new_n16405_), .ZN(new_n16406_));
  OAI21_X1   g16214(.A1(new_n16402_), .A2(new_n275_), .B(new_n16406_), .ZN(new_n16407_));
  NAND2_X1   g16215(.A1(new_n16407_), .A2(new_n16401_), .ZN(new_n16408_));
  OAI22_X1   g16216(.A1(new_n16402_), .A2(new_n275_), .B1(new_n16400_), .B2(new_n16395_), .ZN(new_n16409_));
  INV_X1     g16217(.I(new_n16031_), .ZN(new_n16410_));
  NOR2_X1    g16218(.A1(new_n16410_), .A2(\asqrt[62] ), .ZN(new_n16411_));
  INV_X1     g16219(.I(new_n16411_), .ZN(new_n16412_));
  NAND3_X1   g16220(.A1(new_n16409_), .A2(\asqrt[61] ), .A3(new_n16412_), .ZN(new_n16413_));
  OAI21_X1   g16221(.A1(new_n16413_), .A2(new_n16408_), .B(new_n16033_), .ZN(new_n16414_));
  NAND3_X1   g16222(.A1(new_n16060_), .A2(new_n15409_), .A3(new_n16063_), .ZN(new_n16415_));
  AOI21_X1   g16223(.A1(new_n16415_), .A2(new_n16011_), .B(\asqrt[63] ), .ZN(new_n16416_));
  INV_X1     g16224(.I(new_n16416_), .ZN(new_n16417_));
  OAI21_X1   g16225(.A1(new_n16414_), .A2(new_n16417_), .B(new_n16028_), .ZN(new_n16418_));
  INV_X1     g16226(.I(new_n16042_), .ZN(new_n16419_));
  AOI21_X1   g16227(.A1(new_n16051_), .A2(new_n16419_), .B(new_n16044_), .ZN(new_n16420_));
  NOR3_X1    g16228(.A1(new_n16041_), .A2(new_n16034_), .A3(new_n16039_), .ZN(new_n16421_));
  NOR2_X1    g16229(.A1(new_n16421_), .A2(new_n16420_), .ZN(new_n16422_));
  NOR3_X1    g16230(.A1(new_n16069_), .A2(new_n15422_), .A3(\asqrt[13] ), .ZN(new_n16423_));
  AOI21_X1   g16231(.A1(new_n16066_), .A2(new_n15421_), .B(new_n16060_), .ZN(new_n16424_));
  NOR4_X1    g16232(.A1(new_n16424_), .A2(new_n16423_), .A3(\asqrt[15] ), .A4(new_n16058_), .ZN(new_n16425_));
  NOR2_X1    g16233(.A1(new_n16425_), .A2(new_n16422_), .ZN(new_n16426_));
  NOR3_X1    g16234(.A1(new_n16421_), .A2(new_n16420_), .A3(new_n16058_), .ZN(new_n16427_));
  NOR3_X1    g16235(.A1(new_n16060_), .A2(new_n15445_), .A3(new_n16077_), .ZN(new_n16428_));
  AOI21_X1   g16236(.A1(\asqrt[13] ), .A2(new_n16078_), .B(new_n15446_), .ZN(new_n16429_));
  NOR3_X1    g16237(.A1(new_n16429_), .A2(new_n16428_), .A3(\asqrt[16] ), .ZN(new_n16430_));
  OAI21_X1   g16238(.A1(new_n16427_), .A2(new_n14871_), .B(new_n16430_), .ZN(new_n16431_));
  NAND2_X1   g16239(.A1(new_n16426_), .A2(new_n16431_), .ZN(new_n16432_));
  OAI22_X1   g16240(.A1(new_n16425_), .A2(new_n16422_), .B1(new_n14871_), .B2(new_n16427_), .ZN(new_n16433_));
  INV_X1     g16241(.I(new_n16088_), .ZN(new_n16434_));
  AOI21_X1   g16242(.A1(new_n16433_), .A2(\asqrt[16] ), .B(new_n16434_), .ZN(new_n16435_));
  NOR2_X1    g16243(.A1(new_n16435_), .A2(new_n16432_), .ZN(new_n16436_));
  AOI22_X1   g16244(.A1(new_n16433_), .A2(\asqrt[16] ), .B1(new_n16426_), .B2(new_n16431_), .ZN(new_n16437_));
  INV_X1     g16245(.I(new_n16095_), .ZN(new_n16438_));
  OAI21_X1   g16246(.A1(new_n16437_), .A2(new_n13760_), .B(new_n16438_), .ZN(new_n16439_));
  NAND2_X1   g16247(.A1(new_n16439_), .A2(new_n16436_), .ZN(new_n16440_));
  OAI22_X1   g16248(.A1(new_n16437_), .A2(new_n13760_), .B1(new_n16435_), .B2(new_n16432_), .ZN(new_n16441_));
  AOI21_X1   g16249(.A1(new_n16441_), .A2(\asqrt[18] ), .B(new_n16101_), .ZN(new_n16442_));
  NOR2_X1    g16250(.A1(new_n16442_), .A2(new_n16440_), .ZN(new_n16443_));
  AOI22_X1   g16251(.A1(new_n16441_), .A2(\asqrt[18] ), .B1(new_n16439_), .B2(new_n16436_), .ZN(new_n16444_));
  INV_X1     g16252(.I(new_n16108_), .ZN(new_n16445_));
  OAI21_X1   g16253(.A1(new_n16444_), .A2(new_n12657_), .B(new_n16445_), .ZN(new_n16446_));
  NAND2_X1   g16254(.A1(new_n16446_), .A2(new_n16443_), .ZN(new_n16447_));
  OAI22_X1   g16255(.A1(new_n16444_), .A2(new_n12657_), .B1(new_n16442_), .B2(new_n16440_), .ZN(new_n16448_));
  AOI21_X1   g16256(.A1(new_n16448_), .A2(\asqrt[20] ), .B(new_n16114_), .ZN(new_n16449_));
  NOR2_X1    g16257(.A1(new_n16449_), .A2(new_n16447_), .ZN(new_n16450_));
  AOI22_X1   g16258(.A1(new_n16448_), .A2(\asqrt[20] ), .B1(new_n16446_), .B2(new_n16443_), .ZN(new_n16451_));
  INV_X1     g16259(.I(new_n16121_), .ZN(new_n16452_));
  OAI21_X1   g16260(.A1(new_n16451_), .A2(new_n11631_), .B(new_n16452_), .ZN(new_n16453_));
  NAND2_X1   g16261(.A1(new_n16453_), .A2(new_n16450_), .ZN(new_n16454_));
  OAI22_X1   g16262(.A1(new_n16451_), .A2(new_n11631_), .B1(new_n16449_), .B2(new_n16447_), .ZN(new_n16455_));
  AOI21_X1   g16263(.A1(new_n16455_), .A2(\asqrt[22] ), .B(new_n16127_), .ZN(new_n16456_));
  NOR2_X1    g16264(.A1(new_n16456_), .A2(new_n16454_), .ZN(new_n16457_));
  AOI22_X1   g16265(.A1(new_n16455_), .A2(\asqrt[22] ), .B1(new_n16453_), .B2(new_n16450_), .ZN(new_n16458_));
  INV_X1     g16266(.I(new_n16135_), .ZN(new_n16459_));
  OAI21_X1   g16267(.A1(new_n16458_), .A2(new_n10614_), .B(new_n16459_), .ZN(new_n16460_));
  NAND2_X1   g16268(.A1(new_n16460_), .A2(new_n16457_), .ZN(new_n16461_));
  OAI22_X1   g16269(.A1(new_n16458_), .A2(new_n10614_), .B1(new_n16456_), .B2(new_n16454_), .ZN(new_n16462_));
  AOI21_X1   g16270(.A1(new_n16462_), .A2(\asqrt[24] ), .B(new_n16142_), .ZN(new_n16463_));
  NOR2_X1    g16271(.A1(new_n16463_), .A2(new_n16461_), .ZN(new_n16464_));
  AOI22_X1   g16272(.A1(new_n16462_), .A2(\asqrt[24] ), .B1(new_n16460_), .B2(new_n16457_), .ZN(new_n16465_));
  INV_X1     g16273(.I(new_n16150_), .ZN(new_n16466_));
  OAI21_X1   g16274(.A1(new_n16465_), .A2(new_n9672_), .B(new_n16466_), .ZN(new_n16467_));
  NAND2_X1   g16275(.A1(new_n16467_), .A2(new_n16464_), .ZN(new_n16468_));
  OAI22_X1   g16276(.A1(new_n16465_), .A2(new_n9672_), .B1(new_n16463_), .B2(new_n16461_), .ZN(new_n16469_));
  AOI21_X1   g16277(.A1(new_n16469_), .A2(\asqrt[26] ), .B(new_n16157_), .ZN(new_n16470_));
  NOR2_X1    g16278(.A1(new_n16470_), .A2(new_n16468_), .ZN(new_n16471_));
  AOI22_X1   g16279(.A1(new_n16469_), .A2(\asqrt[26] ), .B1(new_n16467_), .B2(new_n16464_), .ZN(new_n16472_));
  INV_X1     g16280(.I(new_n16165_), .ZN(new_n16473_));
  OAI21_X1   g16281(.A1(new_n16472_), .A2(new_n8763_), .B(new_n16473_), .ZN(new_n16474_));
  NAND2_X1   g16282(.A1(new_n16474_), .A2(new_n16471_), .ZN(new_n16475_));
  OAI22_X1   g16283(.A1(new_n16472_), .A2(new_n8763_), .B1(new_n16470_), .B2(new_n16468_), .ZN(new_n16476_));
  AOI21_X1   g16284(.A1(new_n16476_), .A2(\asqrt[28] ), .B(new_n16172_), .ZN(new_n16477_));
  NOR2_X1    g16285(.A1(new_n16477_), .A2(new_n16475_), .ZN(new_n16478_));
  AOI22_X1   g16286(.A1(new_n16476_), .A2(\asqrt[28] ), .B1(new_n16474_), .B2(new_n16471_), .ZN(new_n16479_));
  INV_X1     g16287(.I(new_n16180_), .ZN(new_n16480_));
  OAI21_X1   g16288(.A1(new_n16479_), .A2(new_n7931_), .B(new_n16480_), .ZN(new_n16481_));
  NAND2_X1   g16289(.A1(new_n16481_), .A2(new_n16478_), .ZN(new_n16482_));
  OAI22_X1   g16290(.A1(new_n16479_), .A2(new_n7931_), .B1(new_n16477_), .B2(new_n16475_), .ZN(new_n16483_));
  AOI21_X1   g16291(.A1(new_n16483_), .A2(\asqrt[30] ), .B(new_n16187_), .ZN(new_n16484_));
  NOR2_X1    g16292(.A1(new_n16484_), .A2(new_n16482_), .ZN(new_n16485_));
  AOI22_X1   g16293(.A1(new_n16483_), .A2(\asqrt[30] ), .B1(new_n16481_), .B2(new_n16478_), .ZN(new_n16486_));
  INV_X1     g16294(.I(new_n16195_), .ZN(new_n16487_));
  OAI21_X1   g16295(.A1(new_n16486_), .A2(new_n7110_), .B(new_n16487_), .ZN(new_n16488_));
  NAND2_X1   g16296(.A1(new_n16488_), .A2(new_n16485_), .ZN(new_n16489_));
  OAI22_X1   g16297(.A1(new_n16486_), .A2(new_n7110_), .B1(new_n16484_), .B2(new_n16482_), .ZN(new_n16490_));
  AOI21_X1   g16298(.A1(new_n16490_), .A2(\asqrt[32] ), .B(new_n16202_), .ZN(new_n16491_));
  NOR2_X1    g16299(.A1(new_n16491_), .A2(new_n16489_), .ZN(new_n16492_));
  AOI22_X1   g16300(.A1(new_n16490_), .A2(\asqrt[32] ), .B1(new_n16488_), .B2(new_n16485_), .ZN(new_n16493_));
  INV_X1     g16301(.I(new_n16210_), .ZN(new_n16494_));
  OAI21_X1   g16302(.A1(new_n16493_), .A2(new_n6365_), .B(new_n16494_), .ZN(new_n16495_));
  NAND2_X1   g16303(.A1(new_n16495_), .A2(new_n16492_), .ZN(new_n16496_));
  OAI22_X1   g16304(.A1(new_n16493_), .A2(new_n6365_), .B1(new_n16491_), .B2(new_n16489_), .ZN(new_n16497_));
  AOI21_X1   g16305(.A1(new_n16497_), .A2(\asqrt[34] ), .B(new_n16217_), .ZN(new_n16498_));
  NOR2_X1    g16306(.A1(new_n16498_), .A2(new_n16496_), .ZN(new_n16499_));
  AOI22_X1   g16307(.A1(new_n16497_), .A2(\asqrt[34] ), .B1(new_n16495_), .B2(new_n16492_), .ZN(new_n16500_));
  INV_X1     g16308(.I(new_n16225_), .ZN(new_n16501_));
  OAI21_X1   g16309(.A1(new_n16500_), .A2(new_n5626_), .B(new_n16501_), .ZN(new_n16502_));
  NAND2_X1   g16310(.A1(new_n16502_), .A2(new_n16499_), .ZN(new_n16503_));
  OAI22_X1   g16311(.A1(new_n16500_), .A2(new_n5626_), .B1(new_n16498_), .B2(new_n16496_), .ZN(new_n16504_));
  AOI21_X1   g16312(.A1(new_n16504_), .A2(\asqrt[36] ), .B(new_n16232_), .ZN(new_n16505_));
  NOR2_X1    g16313(.A1(new_n16505_), .A2(new_n16503_), .ZN(new_n16506_));
  AOI22_X1   g16314(.A1(new_n16504_), .A2(\asqrt[36] ), .B1(new_n16502_), .B2(new_n16499_), .ZN(new_n16507_));
  INV_X1     g16315(.I(new_n16240_), .ZN(new_n16508_));
  OAI21_X1   g16316(.A1(new_n16507_), .A2(new_n4973_), .B(new_n16508_), .ZN(new_n16509_));
  NAND2_X1   g16317(.A1(new_n16509_), .A2(new_n16506_), .ZN(new_n16510_));
  OAI22_X1   g16318(.A1(new_n16507_), .A2(new_n4973_), .B1(new_n16505_), .B2(new_n16503_), .ZN(new_n16511_));
  AOI21_X1   g16319(.A1(new_n16511_), .A2(\asqrt[38] ), .B(new_n16247_), .ZN(new_n16512_));
  NOR2_X1    g16320(.A1(new_n16512_), .A2(new_n16510_), .ZN(new_n16513_));
  AOI22_X1   g16321(.A1(new_n16511_), .A2(\asqrt[38] ), .B1(new_n16509_), .B2(new_n16506_), .ZN(new_n16514_));
  INV_X1     g16322(.I(new_n16255_), .ZN(new_n16515_));
  OAI21_X1   g16323(.A1(new_n16514_), .A2(new_n4330_), .B(new_n16515_), .ZN(new_n16516_));
  NAND2_X1   g16324(.A1(new_n16516_), .A2(new_n16513_), .ZN(new_n16517_));
  OAI22_X1   g16325(.A1(new_n16514_), .A2(new_n4330_), .B1(new_n16512_), .B2(new_n16510_), .ZN(new_n16518_));
  AOI21_X1   g16326(.A1(new_n16518_), .A2(\asqrt[40] ), .B(new_n16262_), .ZN(new_n16519_));
  NOR2_X1    g16327(.A1(new_n16519_), .A2(new_n16517_), .ZN(new_n16520_));
  AOI22_X1   g16328(.A1(new_n16518_), .A2(\asqrt[40] ), .B1(new_n16516_), .B2(new_n16513_), .ZN(new_n16521_));
  INV_X1     g16329(.I(new_n16270_), .ZN(new_n16522_));
  OAI21_X1   g16330(.A1(new_n16521_), .A2(new_n3760_), .B(new_n16522_), .ZN(new_n16523_));
  NAND2_X1   g16331(.A1(new_n16523_), .A2(new_n16520_), .ZN(new_n16524_));
  OAI22_X1   g16332(.A1(new_n16521_), .A2(new_n3760_), .B1(new_n16519_), .B2(new_n16517_), .ZN(new_n16525_));
  AOI21_X1   g16333(.A1(new_n16525_), .A2(\asqrt[42] ), .B(new_n16277_), .ZN(new_n16526_));
  NOR2_X1    g16334(.A1(new_n16526_), .A2(new_n16524_), .ZN(new_n16527_));
  AOI22_X1   g16335(.A1(new_n16525_), .A2(\asqrt[42] ), .B1(new_n16523_), .B2(new_n16520_), .ZN(new_n16528_));
  INV_X1     g16336(.I(new_n16285_), .ZN(new_n16529_));
  OAI21_X1   g16337(.A1(new_n16528_), .A2(new_n3208_), .B(new_n16529_), .ZN(new_n16530_));
  NAND2_X1   g16338(.A1(new_n16530_), .A2(new_n16527_), .ZN(new_n16531_));
  OAI22_X1   g16339(.A1(new_n16528_), .A2(new_n3208_), .B1(new_n16526_), .B2(new_n16524_), .ZN(new_n16532_));
  AOI21_X1   g16340(.A1(new_n16532_), .A2(\asqrt[44] ), .B(new_n16292_), .ZN(new_n16533_));
  NOR2_X1    g16341(.A1(new_n16533_), .A2(new_n16531_), .ZN(new_n16534_));
  AOI22_X1   g16342(.A1(new_n16532_), .A2(\asqrt[44] ), .B1(new_n16530_), .B2(new_n16527_), .ZN(new_n16535_));
  INV_X1     g16343(.I(new_n16300_), .ZN(new_n16536_));
  OAI21_X1   g16344(.A1(new_n16535_), .A2(new_n2728_), .B(new_n16536_), .ZN(new_n16537_));
  NAND2_X1   g16345(.A1(new_n16537_), .A2(new_n16534_), .ZN(new_n16538_));
  OAI22_X1   g16346(.A1(new_n16535_), .A2(new_n2728_), .B1(new_n16533_), .B2(new_n16531_), .ZN(new_n16539_));
  AOI21_X1   g16347(.A1(new_n16539_), .A2(\asqrt[46] ), .B(new_n16307_), .ZN(new_n16540_));
  NOR2_X1    g16348(.A1(new_n16540_), .A2(new_n16538_), .ZN(new_n16541_));
  AOI22_X1   g16349(.A1(new_n16539_), .A2(\asqrt[46] ), .B1(new_n16537_), .B2(new_n16534_), .ZN(new_n16542_));
  INV_X1     g16350(.I(new_n16315_), .ZN(new_n16543_));
  OAI21_X1   g16351(.A1(new_n16542_), .A2(new_n2253_), .B(new_n16543_), .ZN(new_n16544_));
  NAND2_X1   g16352(.A1(new_n16544_), .A2(new_n16541_), .ZN(new_n16545_));
  OAI22_X1   g16353(.A1(new_n16542_), .A2(new_n2253_), .B1(new_n16540_), .B2(new_n16538_), .ZN(new_n16546_));
  AOI21_X1   g16354(.A1(new_n16546_), .A2(\asqrt[48] ), .B(new_n16322_), .ZN(new_n16547_));
  NOR2_X1    g16355(.A1(new_n16547_), .A2(new_n16545_), .ZN(new_n16548_));
  AOI22_X1   g16356(.A1(new_n16546_), .A2(\asqrt[48] ), .B1(new_n16544_), .B2(new_n16541_), .ZN(new_n16549_));
  INV_X1     g16357(.I(new_n16330_), .ZN(new_n16550_));
  OAI21_X1   g16358(.A1(new_n16549_), .A2(new_n1854_), .B(new_n16550_), .ZN(new_n16551_));
  NAND2_X1   g16359(.A1(new_n16551_), .A2(new_n16548_), .ZN(new_n16552_));
  OAI22_X1   g16360(.A1(new_n16549_), .A2(new_n1854_), .B1(new_n16547_), .B2(new_n16545_), .ZN(new_n16553_));
  AOI21_X1   g16361(.A1(new_n16553_), .A2(\asqrt[50] ), .B(new_n16337_), .ZN(new_n16554_));
  NOR2_X1    g16362(.A1(new_n16554_), .A2(new_n16552_), .ZN(new_n16555_));
  AOI22_X1   g16363(.A1(new_n16553_), .A2(\asqrt[50] ), .B1(new_n16551_), .B2(new_n16548_), .ZN(new_n16556_));
  INV_X1     g16364(.I(new_n16345_), .ZN(new_n16557_));
  OAI21_X1   g16365(.A1(new_n16556_), .A2(new_n1436_), .B(new_n16557_), .ZN(new_n16558_));
  NAND2_X1   g16366(.A1(new_n16558_), .A2(new_n16555_), .ZN(new_n16559_));
  OAI22_X1   g16367(.A1(new_n16556_), .A2(new_n1436_), .B1(new_n16554_), .B2(new_n16552_), .ZN(new_n16560_));
  AOI21_X1   g16368(.A1(new_n16560_), .A2(\asqrt[52] ), .B(new_n16352_), .ZN(new_n16561_));
  NOR2_X1    g16369(.A1(new_n16561_), .A2(new_n16559_), .ZN(new_n16562_));
  AOI22_X1   g16370(.A1(new_n16560_), .A2(\asqrt[52] ), .B1(new_n16558_), .B2(new_n16555_), .ZN(new_n16563_));
  INV_X1     g16371(.I(new_n16360_), .ZN(new_n16564_));
  OAI21_X1   g16372(.A1(new_n16563_), .A2(new_n1096_), .B(new_n16564_), .ZN(new_n16565_));
  NAND2_X1   g16373(.A1(new_n16565_), .A2(new_n16562_), .ZN(new_n16566_));
  OAI22_X1   g16374(.A1(new_n16563_), .A2(new_n1096_), .B1(new_n16561_), .B2(new_n16559_), .ZN(new_n16567_));
  AOI21_X1   g16375(.A1(new_n16567_), .A2(\asqrt[54] ), .B(new_n16366_), .ZN(new_n16568_));
  NOR2_X1    g16376(.A1(new_n16568_), .A2(new_n16566_), .ZN(new_n16569_));
  AOI22_X1   g16377(.A1(new_n16567_), .A2(\asqrt[54] ), .B1(new_n16565_), .B2(new_n16562_), .ZN(new_n16570_));
  INV_X1     g16378(.I(new_n16373_), .ZN(new_n16571_));
  OAI21_X1   g16379(.A1(new_n16570_), .A2(new_n825_), .B(new_n16571_), .ZN(new_n16572_));
  NAND2_X1   g16380(.A1(new_n16572_), .A2(new_n16569_), .ZN(new_n16573_));
  OAI22_X1   g16381(.A1(new_n16570_), .A2(new_n825_), .B1(new_n16568_), .B2(new_n16566_), .ZN(new_n16574_));
  AOI21_X1   g16382(.A1(new_n16574_), .A2(\asqrt[56] ), .B(new_n16379_), .ZN(new_n16575_));
  NOR2_X1    g16383(.A1(new_n16575_), .A2(new_n16573_), .ZN(new_n16576_));
  AOI22_X1   g16384(.A1(new_n16574_), .A2(\asqrt[56] ), .B1(new_n16572_), .B2(new_n16569_), .ZN(new_n16577_));
  INV_X1     g16385(.I(new_n16386_), .ZN(new_n16578_));
  OAI21_X1   g16386(.A1(new_n16577_), .A2(new_n587_), .B(new_n16578_), .ZN(new_n16579_));
  NAND2_X1   g16387(.A1(new_n16579_), .A2(new_n16576_), .ZN(new_n16580_));
  OAI22_X1   g16388(.A1(new_n16577_), .A2(new_n587_), .B1(new_n16575_), .B2(new_n16573_), .ZN(new_n16581_));
  AOI21_X1   g16389(.A1(new_n16581_), .A2(\asqrt[58] ), .B(new_n16392_), .ZN(new_n16582_));
  NOR2_X1    g16390(.A1(new_n16582_), .A2(new_n16580_), .ZN(new_n16583_));
  AOI22_X1   g16391(.A1(new_n16581_), .A2(\asqrt[58] ), .B1(new_n16579_), .B2(new_n16576_), .ZN(new_n16584_));
  INV_X1     g16392(.I(new_n16399_), .ZN(new_n16585_));
  OAI21_X1   g16393(.A1(new_n16584_), .A2(new_n376_), .B(new_n16585_), .ZN(new_n16586_));
  NAND2_X1   g16394(.A1(new_n16586_), .A2(new_n16583_), .ZN(new_n16587_));
  OAI22_X1   g16395(.A1(new_n16584_), .A2(new_n376_), .B1(new_n16582_), .B2(new_n16580_), .ZN(new_n16588_));
  AOI21_X1   g16396(.A1(new_n16588_), .A2(\asqrt[60] ), .B(new_n16405_), .ZN(new_n16589_));
  AOI22_X1   g16397(.A1(new_n16588_), .A2(\asqrt[60] ), .B1(new_n16586_), .B2(new_n16583_), .ZN(new_n16590_));
  OAI22_X1   g16398(.A1(new_n16590_), .A2(new_n229_), .B1(new_n16589_), .B2(new_n16587_), .ZN(new_n16591_));
  NOR4_X1    g16399(.A1(new_n16591_), .A2(\asqrt[62] ), .A3(new_n16027_), .A4(new_n16031_), .ZN(new_n16592_));
  NAND2_X1   g16400(.A1(new_n16047_), .A2(new_n15409_), .ZN(new_n16593_));
  XOR2_X1    g16401(.A1(new_n16047_), .A2(\asqrt[63] ), .Z(new_n16594_));
  AOI21_X1   g16402(.A1(\asqrt[13] ), .A2(new_n16593_), .B(new_n16594_), .ZN(new_n16595_));
  NAND2_X1   g16403(.A1(new_n16592_), .A2(new_n16595_), .ZN(new_n16596_));
  NOR4_X1    g16404(.A1(new_n16596_), .A2(new_n16008_), .A3(new_n16418_), .A4(new_n16015_), .ZN(new_n16597_));
  NOR2_X1    g16405(.A1(new_n16008_), .A2(\a[24] ), .ZN(new_n16598_));
  OAI21_X1   g16406(.A1(new_n16597_), .A2(new_n16598_), .B(new_n16007_), .ZN(new_n16599_));
  INV_X1     g16407(.I(new_n16007_), .ZN(new_n16600_));
  INV_X1     g16408(.I(new_n16015_), .ZN(new_n16601_));
  NOR2_X1    g16409(.A1(new_n16589_), .A2(new_n16587_), .ZN(new_n16602_));
  NOR3_X1    g16410(.A1(new_n16590_), .A2(new_n229_), .A3(new_n16411_), .ZN(new_n16603_));
  AOI21_X1   g16411(.A1(new_n16603_), .A2(new_n16602_), .B(new_n16032_), .ZN(new_n16604_));
  AOI21_X1   g16412(.A1(new_n16604_), .A2(new_n16416_), .B(new_n16027_), .ZN(new_n16605_));
  AOI22_X1   g16413(.A1(new_n16409_), .A2(\asqrt[61] ), .B1(new_n16407_), .B2(new_n16401_), .ZN(new_n16606_));
  NAND4_X1   g16414(.A1(new_n16606_), .A2(new_n196_), .A3(new_n16028_), .A4(new_n16410_), .ZN(new_n16607_));
  INV_X1     g16415(.I(new_n16595_), .ZN(new_n16608_));
  NOR2_X1    g16416(.A1(new_n16607_), .A2(new_n16608_), .ZN(new_n16609_));
  NAND4_X1   g16417(.A1(new_n16609_), .A2(new_n16605_), .A3(\a[25] ), .A4(new_n16601_), .ZN(new_n16610_));
  NAND3_X1   g16418(.A1(new_n16610_), .A2(\a[24] ), .A3(new_n16600_), .ZN(new_n16611_));
  NAND2_X1   g16419(.A1(new_n16599_), .A2(new_n16611_), .ZN(new_n16612_));
  NOR2_X1    g16420(.A1(new_n16596_), .A2(new_n16418_), .ZN(new_n16613_));
  NOR4_X1    g16421(.A1(new_n16013_), .A2(new_n15409_), .A3(new_n16062_), .A4(new_n16000_), .ZN(new_n16614_));
  NAND2_X1   g16422(.A1(\asqrt[13] ), .A2(\a[24] ), .ZN(new_n16615_));
  XOR2_X1    g16423(.A1(new_n16615_), .A2(new_n16614_), .Z(new_n16616_));
  NOR2_X1    g16424(.A1(new_n16616_), .A2(new_n16004_), .ZN(new_n16617_));
  INV_X1     g16425(.I(new_n16617_), .ZN(new_n16618_));
  NAND3_X1   g16426(.A1(new_n16609_), .A2(new_n16605_), .A3(new_n16601_), .ZN(new_n16619_));
  NAND2_X1   g16427(.A1(new_n16370_), .A2(\asqrt[55] ), .ZN(new_n16620_));
  AOI21_X1   g16428(.A1(new_n16620_), .A2(new_n16369_), .B(new_n724_), .ZN(new_n16621_));
  OAI21_X1   g16429(.A1(new_n16375_), .A2(new_n16621_), .B(\asqrt[57] ), .ZN(new_n16622_));
  AOI21_X1   g16430(.A1(new_n16382_), .A2(new_n16622_), .B(new_n504_), .ZN(new_n16623_));
  OAI21_X1   g16431(.A1(new_n16388_), .A2(new_n16623_), .B(\asqrt[59] ), .ZN(new_n16624_));
  AOI21_X1   g16432(.A1(new_n16395_), .A2(new_n16624_), .B(new_n275_), .ZN(new_n16625_));
  OAI21_X1   g16433(.A1(new_n16401_), .A2(new_n16625_), .B(\asqrt[61] ), .ZN(new_n16626_));
  NOR3_X1    g16434(.A1(new_n16408_), .A2(new_n16626_), .A3(new_n16411_), .ZN(new_n16627_));
  NOR3_X1    g16435(.A1(new_n16627_), .A2(new_n16032_), .A3(new_n16417_), .ZN(new_n16628_));
  OAI21_X1   g16436(.A1(new_n16628_), .A2(new_n16027_), .B(new_n16607_), .ZN(new_n16629_));
  NOR2_X1    g16437(.A1(new_n16601_), .A2(new_n16595_), .ZN(new_n16630_));
  NAND2_X1   g16438(.A1(new_n16630_), .A2(\asqrt[13] ), .ZN(new_n16631_));
  OAI21_X1   g16439(.A1(new_n16629_), .A2(new_n16631_), .B(new_n16034_), .ZN(new_n16632_));
  NAND3_X1   g16440(.A1(new_n16632_), .A2(new_n16035_), .A3(new_n16619_), .ZN(new_n16633_));
  NOR3_X1    g16441(.A1(new_n16596_), .A2(new_n16015_), .A3(new_n16418_), .ZN(\asqrt[12] ));
  NAND2_X1   g16442(.A1(new_n16567_), .A2(\asqrt[54] ), .ZN(new_n16635_));
  AOI21_X1   g16443(.A1(new_n16635_), .A2(new_n16566_), .B(new_n825_), .ZN(new_n16636_));
  OAI21_X1   g16444(.A1(new_n16569_), .A2(new_n16636_), .B(\asqrt[56] ), .ZN(new_n16637_));
  AOI21_X1   g16445(.A1(new_n16573_), .A2(new_n16637_), .B(new_n587_), .ZN(new_n16638_));
  OAI21_X1   g16446(.A1(new_n16576_), .A2(new_n16638_), .B(\asqrt[58] ), .ZN(new_n16639_));
  AOI21_X1   g16447(.A1(new_n16580_), .A2(new_n16639_), .B(new_n376_), .ZN(new_n16640_));
  OAI21_X1   g16448(.A1(new_n16583_), .A2(new_n16640_), .B(\asqrt[60] ), .ZN(new_n16641_));
  AOI21_X1   g16449(.A1(new_n16587_), .A2(new_n16641_), .B(new_n229_), .ZN(new_n16642_));
  NAND4_X1   g16450(.A1(new_n16642_), .A2(new_n16401_), .A3(new_n16407_), .A4(new_n16412_), .ZN(new_n16643_));
  NAND3_X1   g16451(.A1(new_n16643_), .A2(new_n16033_), .A3(new_n16416_), .ZN(new_n16644_));
  AOI21_X1   g16452(.A1(new_n16028_), .A2(new_n16644_), .B(new_n16592_), .ZN(new_n16645_));
  INV_X1     g16453(.I(new_n16631_), .ZN(new_n16646_));
  AOI21_X1   g16454(.A1(new_n16645_), .A2(new_n16646_), .B(\a[26] ), .ZN(new_n16647_));
  OAI21_X1   g16455(.A1(new_n16647_), .A2(new_n16036_), .B(\asqrt[12] ), .ZN(new_n16648_));
  NAND4_X1   g16456(.A1(new_n16648_), .A2(new_n16633_), .A3(new_n15447_), .A4(new_n16618_), .ZN(new_n16649_));
  NAND2_X1   g16457(.A1(new_n16649_), .A2(new_n16612_), .ZN(new_n16650_));
  NAND3_X1   g16458(.A1(new_n16599_), .A2(new_n16611_), .A3(new_n16618_), .ZN(new_n16651_));
  AOI21_X1   g16459(.A1(\asqrt[13] ), .A2(new_n16034_), .B(\a[27] ), .ZN(new_n16652_));
  NOR2_X1    g16460(.A1(new_n16051_), .A2(\a[26] ), .ZN(new_n16653_));
  AOI21_X1   g16461(.A1(\asqrt[13] ), .A2(\a[26] ), .B(new_n16038_), .ZN(new_n16654_));
  OAI21_X1   g16462(.A1(new_n16653_), .A2(new_n16652_), .B(new_n16654_), .ZN(new_n16655_));
  INV_X1     g16463(.I(new_n16655_), .ZN(new_n16656_));
  NAND3_X1   g16464(.A1(\asqrt[12] ), .A2(new_n16059_), .A3(new_n16656_), .ZN(new_n16657_));
  OAI21_X1   g16465(.A1(new_n16619_), .A2(new_n16655_), .B(new_n16058_), .ZN(new_n16658_));
  NAND3_X1   g16466(.A1(new_n16657_), .A2(new_n16658_), .A3(new_n14871_), .ZN(new_n16659_));
  AOI21_X1   g16467(.A1(new_n16651_), .A2(\asqrt[14] ), .B(new_n16659_), .ZN(new_n16660_));
  NOR2_X1    g16468(.A1(new_n16650_), .A2(new_n16660_), .ZN(new_n16661_));
  AOI22_X1   g16469(.A1(new_n16649_), .A2(new_n16612_), .B1(\asqrt[14] ), .B2(new_n16651_), .ZN(new_n16662_));
  NAND2_X1   g16470(.A1(new_n16073_), .A2(\asqrt[15] ), .ZN(new_n16663_));
  INV_X1     g16471(.I(new_n16663_), .ZN(new_n16664_));
  NAND2_X1   g16472(.A1(new_n16067_), .A2(new_n16070_), .ZN(new_n16665_));
  NAND3_X1   g16473(.A1(new_n16665_), .A2(new_n16427_), .A3(new_n14871_), .ZN(new_n16666_));
  NOR3_X1    g16474(.A1(new_n16619_), .A2(new_n16664_), .A3(new_n16666_), .ZN(new_n16667_));
  NOR2_X1    g16475(.A1(new_n16619_), .A2(new_n16666_), .ZN(new_n16668_));
  NOR2_X1    g16476(.A1(new_n16668_), .A2(new_n16663_), .ZN(new_n16669_));
  NOR3_X1    g16477(.A1(new_n16669_), .A2(\asqrt[16] ), .A3(new_n16667_), .ZN(new_n16670_));
  OAI21_X1   g16478(.A1(new_n16662_), .A2(new_n14871_), .B(new_n16670_), .ZN(new_n16671_));
  NAND2_X1   g16479(.A1(new_n16651_), .A2(\asqrt[14] ), .ZN(new_n16672_));
  AOI21_X1   g16480(.A1(new_n16650_), .A2(new_n16672_), .B(new_n14871_), .ZN(new_n16673_));
  OAI21_X1   g16481(.A1(new_n16673_), .A2(new_n16661_), .B(\asqrt[16] ), .ZN(new_n16674_));
  NAND2_X1   g16482(.A1(new_n16433_), .A2(\asqrt[16] ), .ZN(new_n16675_));
  NOR2_X1    g16483(.A1(new_n16429_), .A2(new_n16428_), .ZN(new_n16676_));
  NOR4_X1    g16484(.A1(new_n16619_), .A2(\asqrt[16] ), .A3(new_n16676_), .A4(new_n16433_), .ZN(new_n16677_));
  XOR2_X1    g16485(.A1(new_n16677_), .A2(new_n16675_), .Z(new_n16678_));
  NAND2_X1   g16486(.A1(new_n16678_), .A2(new_n13760_), .ZN(new_n16679_));
  INV_X1     g16487(.I(new_n16679_), .ZN(new_n16680_));
  NAND2_X1   g16488(.A1(new_n16674_), .A2(new_n16680_), .ZN(new_n16681_));
  NAND3_X1   g16489(.A1(new_n16681_), .A2(new_n16661_), .A3(new_n16671_), .ZN(new_n16682_));
  INV_X1     g16490(.I(new_n16598_), .ZN(new_n16683_));
  AOI21_X1   g16491(.A1(new_n16610_), .A2(new_n16683_), .B(new_n16600_), .ZN(new_n16684_));
  NOR3_X1    g16492(.A1(new_n16597_), .A2(new_n15995_), .A3(new_n16007_), .ZN(new_n16685_));
  NOR2_X1    g16493(.A1(new_n16685_), .A2(new_n16684_), .ZN(new_n16686_));
  NOR3_X1    g16494(.A1(new_n16647_), .A2(new_n16036_), .A3(\asqrt[12] ), .ZN(new_n16687_));
  AOI21_X1   g16495(.A1(new_n16632_), .A2(new_n16035_), .B(new_n16619_), .ZN(new_n16688_));
  NOR4_X1    g16496(.A1(new_n16687_), .A2(new_n16688_), .A3(\asqrt[14] ), .A4(new_n16617_), .ZN(new_n16689_));
  NOR2_X1    g16497(.A1(new_n16689_), .A2(new_n16686_), .ZN(new_n16690_));
  NOR3_X1    g16498(.A1(new_n16685_), .A2(new_n16684_), .A3(new_n16617_), .ZN(new_n16691_));
  NOR3_X1    g16499(.A1(new_n16619_), .A2(new_n16058_), .A3(new_n16655_), .ZN(new_n16692_));
  AOI21_X1   g16500(.A1(\asqrt[12] ), .A2(new_n16656_), .B(new_n16059_), .ZN(new_n16693_));
  NOR3_X1    g16501(.A1(new_n16693_), .A2(new_n16692_), .A3(\asqrt[15] ), .ZN(new_n16694_));
  OAI21_X1   g16502(.A1(new_n16691_), .A2(new_n15447_), .B(new_n16694_), .ZN(new_n16695_));
  NAND2_X1   g16503(.A1(new_n16690_), .A2(new_n16695_), .ZN(new_n16696_));
  OAI22_X1   g16504(.A1(new_n16689_), .A2(new_n16686_), .B1(new_n15447_), .B2(new_n16691_), .ZN(new_n16697_));
  INV_X1     g16505(.I(new_n16670_), .ZN(new_n16698_));
  AOI21_X1   g16506(.A1(new_n16697_), .A2(\asqrt[15] ), .B(new_n16698_), .ZN(new_n16699_));
  AOI22_X1   g16507(.A1(new_n16697_), .A2(\asqrt[15] ), .B1(new_n16690_), .B2(new_n16695_), .ZN(new_n16700_));
  OAI22_X1   g16508(.A1(new_n16700_), .A2(new_n14273_), .B1(new_n16699_), .B2(new_n16696_), .ZN(new_n16701_));
  NAND2_X1   g16509(.A1(new_n16091_), .A2(\asqrt[17] ), .ZN(new_n16702_));
  NOR2_X1    g16510(.A1(new_n16086_), .A2(new_n16087_), .ZN(new_n16703_));
  NOR4_X1    g16511(.A1(new_n16619_), .A2(\asqrt[17] ), .A3(new_n16703_), .A4(new_n16091_), .ZN(new_n16704_));
  XOR2_X1    g16512(.A1(new_n16704_), .A2(new_n16702_), .Z(new_n16705_));
  NAND2_X1   g16513(.A1(new_n16705_), .A2(new_n13192_), .ZN(new_n16706_));
  AOI21_X1   g16514(.A1(new_n16701_), .A2(\asqrt[17] ), .B(new_n16706_), .ZN(new_n16707_));
  NOR2_X1    g16515(.A1(new_n16707_), .A2(new_n16682_), .ZN(new_n16708_));
  OAI21_X1   g16516(.A1(new_n16673_), .A2(new_n16698_), .B(new_n16661_), .ZN(new_n16709_));
  AOI21_X1   g16517(.A1(new_n16674_), .A2(new_n16680_), .B(new_n16709_), .ZN(new_n16710_));
  AOI21_X1   g16518(.A1(new_n16709_), .A2(new_n16674_), .B(new_n13760_), .ZN(new_n16711_));
  OAI21_X1   g16519(.A1(new_n16710_), .A2(new_n16711_), .B(\asqrt[18] ), .ZN(new_n16712_));
  NOR4_X1    g16520(.A1(new_n16619_), .A2(\asqrt[18] ), .A3(new_n16094_), .A4(new_n16441_), .ZN(new_n16713_));
  AOI21_X1   g16521(.A1(new_n16702_), .A2(new_n16090_), .B(new_n13192_), .ZN(new_n16714_));
  NOR2_X1    g16522(.A1(new_n16713_), .A2(new_n16714_), .ZN(new_n16715_));
  NAND2_X1   g16523(.A1(new_n16715_), .A2(new_n12657_), .ZN(new_n16716_));
  INV_X1     g16524(.I(new_n16716_), .ZN(new_n16717_));
  NAND2_X1   g16525(.A1(new_n16712_), .A2(new_n16717_), .ZN(new_n16718_));
  NAND2_X1   g16526(.A1(new_n16718_), .A2(new_n16708_), .ZN(new_n16719_));
  NOR2_X1    g16527(.A1(new_n16710_), .A2(new_n16711_), .ZN(new_n16720_));
  OAI22_X1   g16528(.A1(new_n16720_), .A2(new_n13192_), .B1(new_n16707_), .B2(new_n16682_), .ZN(new_n16721_));
  NAND2_X1   g16529(.A1(new_n16105_), .A2(\asqrt[19] ), .ZN(new_n16722_));
  NOR4_X1    g16530(.A1(new_n16619_), .A2(\asqrt[19] ), .A3(new_n16100_), .A4(new_n16105_), .ZN(new_n16723_));
  XOR2_X1    g16531(.A1(new_n16723_), .A2(new_n16722_), .Z(new_n16724_));
  NAND2_X1   g16532(.A1(new_n16724_), .A2(new_n12101_), .ZN(new_n16725_));
  AOI21_X1   g16533(.A1(new_n16721_), .A2(\asqrt[19] ), .B(new_n16725_), .ZN(new_n16726_));
  NOR2_X1    g16534(.A1(new_n16726_), .A2(new_n16719_), .ZN(new_n16727_));
  OAI21_X1   g16535(.A1(new_n16711_), .A2(new_n16706_), .B(new_n16710_), .ZN(new_n16728_));
  AOI21_X1   g16536(.A1(new_n16712_), .A2(new_n16717_), .B(new_n16728_), .ZN(new_n16729_));
  AOI21_X1   g16537(.A1(new_n16728_), .A2(new_n16712_), .B(new_n12657_), .ZN(new_n16730_));
  OAI21_X1   g16538(.A1(new_n16729_), .A2(new_n16730_), .B(\asqrt[20] ), .ZN(new_n16731_));
  NOR4_X1    g16539(.A1(new_n16619_), .A2(\asqrt[20] ), .A3(new_n16107_), .A4(new_n16448_), .ZN(new_n16732_));
  AOI21_X1   g16540(.A1(new_n16722_), .A2(new_n16104_), .B(new_n12101_), .ZN(new_n16733_));
  NOR2_X1    g16541(.A1(new_n16732_), .A2(new_n16733_), .ZN(new_n16734_));
  NAND2_X1   g16542(.A1(new_n16734_), .A2(new_n11631_), .ZN(new_n16735_));
  INV_X1     g16543(.I(new_n16735_), .ZN(new_n16736_));
  NAND2_X1   g16544(.A1(new_n16731_), .A2(new_n16736_), .ZN(new_n16737_));
  NAND2_X1   g16545(.A1(new_n16737_), .A2(new_n16727_), .ZN(new_n16738_));
  AOI22_X1   g16546(.A1(new_n16721_), .A2(\asqrt[19] ), .B1(new_n16718_), .B2(new_n16708_), .ZN(new_n16739_));
  OAI22_X1   g16547(.A1(new_n16739_), .A2(new_n12101_), .B1(new_n16726_), .B2(new_n16719_), .ZN(new_n16740_));
  NAND2_X1   g16548(.A1(new_n16118_), .A2(\asqrt[21] ), .ZN(new_n16741_));
  NOR4_X1    g16549(.A1(new_n16619_), .A2(\asqrt[21] ), .A3(new_n16113_), .A4(new_n16118_), .ZN(new_n16742_));
  XOR2_X1    g16550(.A1(new_n16742_), .A2(new_n16741_), .Z(new_n16743_));
  NAND2_X1   g16551(.A1(new_n16743_), .A2(new_n11105_), .ZN(new_n16744_));
  AOI21_X1   g16552(.A1(new_n16740_), .A2(\asqrt[21] ), .B(new_n16744_), .ZN(new_n16745_));
  NOR2_X1    g16553(.A1(new_n16745_), .A2(new_n16738_), .ZN(new_n16746_));
  AOI22_X1   g16554(.A1(new_n16740_), .A2(\asqrt[21] ), .B1(new_n16737_), .B2(new_n16727_), .ZN(new_n16747_));
  NOR4_X1    g16555(.A1(new_n16619_), .A2(\asqrt[22] ), .A3(new_n16120_), .A4(new_n16455_), .ZN(new_n16748_));
  AOI21_X1   g16556(.A1(new_n16741_), .A2(new_n16117_), .B(new_n11105_), .ZN(new_n16749_));
  NOR2_X1    g16557(.A1(new_n16748_), .A2(new_n16749_), .ZN(new_n16750_));
  NAND2_X1   g16558(.A1(new_n16750_), .A2(new_n10614_), .ZN(new_n16751_));
  INV_X1     g16559(.I(new_n16751_), .ZN(new_n16752_));
  OAI21_X1   g16560(.A1(new_n16747_), .A2(new_n11105_), .B(new_n16752_), .ZN(new_n16753_));
  NAND2_X1   g16561(.A1(new_n16753_), .A2(new_n16746_), .ZN(new_n16754_));
  OAI22_X1   g16562(.A1(new_n16747_), .A2(new_n11105_), .B1(new_n16745_), .B2(new_n16738_), .ZN(new_n16755_));
  NAND2_X1   g16563(.A1(new_n16131_), .A2(\asqrt[23] ), .ZN(new_n16756_));
  NOR4_X1    g16564(.A1(new_n16619_), .A2(\asqrt[23] ), .A3(new_n16126_), .A4(new_n16131_), .ZN(new_n16757_));
  XOR2_X1    g16565(.A1(new_n16757_), .A2(new_n16756_), .Z(new_n16758_));
  NAND2_X1   g16566(.A1(new_n16758_), .A2(new_n10104_), .ZN(new_n16759_));
  AOI21_X1   g16567(.A1(new_n16755_), .A2(\asqrt[23] ), .B(new_n16759_), .ZN(new_n16760_));
  NOR2_X1    g16568(.A1(new_n16760_), .A2(new_n16754_), .ZN(new_n16761_));
  AOI22_X1   g16569(.A1(new_n16755_), .A2(\asqrt[23] ), .B1(new_n16753_), .B2(new_n16746_), .ZN(new_n16762_));
  NAND2_X1   g16570(.A1(new_n16462_), .A2(\asqrt[24] ), .ZN(new_n16763_));
  NOR4_X1    g16571(.A1(new_n16619_), .A2(\asqrt[24] ), .A3(new_n16134_), .A4(new_n16462_), .ZN(new_n16764_));
  XOR2_X1    g16572(.A1(new_n16764_), .A2(new_n16763_), .Z(new_n16765_));
  NAND2_X1   g16573(.A1(new_n16765_), .A2(new_n9672_), .ZN(new_n16766_));
  INV_X1     g16574(.I(new_n16766_), .ZN(new_n16767_));
  OAI21_X1   g16575(.A1(new_n16762_), .A2(new_n10104_), .B(new_n16767_), .ZN(new_n16768_));
  NAND2_X1   g16576(.A1(new_n16768_), .A2(new_n16761_), .ZN(new_n16769_));
  OAI22_X1   g16577(.A1(new_n16762_), .A2(new_n10104_), .B1(new_n16760_), .B2(new_n16754_), .ZN(new_n16770_));
  NOR4_X1    g16578(.A1(new_n16619_), .A2(\asqrt[25] ), .A3(new_n16141_), .A4(new_n16146_), .ZN(new_n16771_));
  AOI21_X1   g16579(.A1(new_n16763_), .A2(new_n16461_), .B(new_n9672_), .ZN(new_n16772_));
  NOR2_X1    g16580(.A1(new_n16771_), .A2(new_n16772_), .ZN(new_n16773_));
  NAND2_X1   g16581(.A1(new_n16773_), .A2(new_n9212_), .ZN(new_n16774_));
  AOI21_X1   g16582(.A1(new_n16770_), .A2(\asqrt[25] ), .B(new_n16774_), .ZN(new_n16775_));
  NOR2_X1    g16583(.A1(new_n16775_), .A2(new_n16769_), .ZN(new_n16776_));
  AOI22_X1   g16584(.A1(new_n16770_), .A2(\asqrt[25] ), .B1(new_n16768_), .B2(new_n16761_), .ZN(new_n16777_));
  NAND2_X1   g16585(.A1(new_n16469_), .A2(\asqrt[26] ), .ZN(new_n16778_));
  NOR4_X1    g16586(.A1(new_n16619_), .A2(\asqrt[26] ), .A3(new_n16149_), .A4(new_n16469_), .ZN(new_n16779_));
  XOR2_X1    g16587(.A1(new_n16779_), .A2(new_n16778_), .Z(new_n16780_));
  NAND2_X1   g16588(.A1(new_n16780_), .A2(new_n8763_), .ZN(new_n16781_));
  INV_X1     g16589(.I(new_n16781_), .ZN(new_n16782_));
  OAI21_X1   g16590(.A1(new_n16777_), .A2(new_n9212_), .B(new_n16782_), .ZN(new_n16783_));
  NAND2_X1   g16591(.A1(new_n16783_), .A2(new_n16776_), .ZN(new_n16784_));
  OAI22_X1   g16592(.A1(new_n16777_), .A2(new_n9212_), .B1(new_n16775_), .B2(new_n16769_), .ZN(new_n16785_));
  NOR4_X1    g16593(.A1(new_n16619_), .A2(\asqrt[27] ), .A3(new_n16156_), .A4(new_n16161_), .ZN(new_n16786_));
  AOI21_X1   g16594(.A1(new_n16778_), .A2(new_n16468_), .B(new_n8763_), .ZN(new_n16787_));
  NOR2_X1    g16595(.A1(new_n16786_), .A2(new_n16787_), .ZN(new_n16788_));
  NAND2_X1   g16596(.A1(new_n16788_), .A2(new_n8319_), .ZN(new_n16789_));
  AOI21_X1   g16597(.A1(new_n16785_), .A2(\asqrt[27] ), .B(new_n16789_), .ZN(new_n16790_));
  NOR2_X1    g16598(.A1(new_n16790_), .A2(new_n16784_), .ZN(new_n16791_));
  AOI22_X1   g16599(.A1(new_n16785_), .A2(\asqrt[27] ), .B1(new_n16783_), .B2(new_n16776_), .ZN(new_n16792_));
  NAND2_X1   g16600(.A1(new_n16476_), .A2(\asqrt[28] ), .ZN(new_n16793_));
  NOR4_X1    g16601(.A1(new_n16619_), .A2(\asqrt[28] ), .A3(new_n16164_), .A4(new_n16476_), .ZN(new_n16794_));
  XOR2_X1    g16602(.A1(new_n16794_), .A2(new_n16793_), .Z(new_n16795_));
  NAND2_X1   g16603(.A1(new_n16795_), .A2(new_n7931_), .ZN(new_n16796_));
  INV_X1     g16604(.I(new_n16796_), .ZN(new_n16797_));
  OAI21_X1   g16605(.A1(new_n16792_), .A2(new_n8319_), .B(new_n16797_), .ZN(new_n16798_));
  NAND2_X1   g16606(.A1(new_n16798_), .A2(new_n16791_), .ZN(new_n16799_));
  OAI22_X1   g16607(.A1(new_n16792_), .A2(new_n8319_), .B1(new_n16790_), .B2(new_n16784_), .ZN(new_n16800_));
  NOR4_X1    g16608(.A1(new_n16619_), .A2(\asqrt[29] ), .A3(new_n16171_), .A4(new_n16176_), .ZN(new_n16801_));
  AOI21_X1   g16609(.A1(new_n16793_), .A2(new_n16475_), .B(new_n7931_), .ZN(new_n16802_));
  NOR2_X1    g16610(.A1(new_n16801_), .A2(new_n16802_), .ZN(new_n16803_));
  NAND2_X1   g16611(.A1(new_n16803_), .A2(new_n7517_), .ZN(new_n16804_));
  AOI21_X1   g16612(.A1(new_n16800_), .A2(\asqrt[29] ), .B(new_n16804_), .ZN(new_n16805_));
  NOR2_X1    g16613(.A1(new_n16805_), .A2(new_n16799_), .ZN(new_n16806_));
  AOI22_X1   g16614(.A1(new_n16800_), .A2(\asqrt[29] ), .B1(new_n16798_), .B2(new_n16791_), .ZN(new_n16807_));
  NAND2_X1   g16615(.A1(new_n16483_), .A2(\asqrt[30] ), .ZN(new_n16808_));
  NOR4_X1    g16616(.A1(new_n16619_), .A2(\asqrt[30] ), .A3(new_n16179_), .A4(new_n16483_), .ZN(new_n16809_));
  XOR2_X1    g16617(.A1(new_n16809_), .A2(new_n16808_), .Z(new_n16810_));
  NAND2_X1   g16618(.A1(new_n16810_), .A2(new_n7110_), .ZN(new_n16811_));
  INV_X1     g16619(.I(new_n16811_), .ZN(new_n16812_));
  OAI21_X1   g16620(.A1(new_n16807_), .A2(new_n7517_), .B(new_n16812_), .ZN(new_n16813_));
  NAND2_X1   g16621(.A1(new_n16813_), .A2(new_n16806_), .ZN(new_n16814_));
  OAI22_X1   g16622(.A1(new_n16807_), .A2(new_n7517_), .B1(new_n16805_), .B2(new_n16799_), .ZN(new_n16815_));
  NOR4_X1    g16623(.A1(new_n16619_), .A2(\asqrt[31] ), .A3(new_n16186_), .A4(new_n16191_), .ZN(new_n16816_));
  AOI21_X1   g16624(.A1(new_n16808_), .A2(new_n16482_), .B(new_n7110_), .ZN(new_n16817_));
  NOR2_X1    g16625(.A1(new_n16816_), .A2(new_n16817_), .ZN(new_n16818_));
  NAND2_X1   g16626(.A1(new_n16818_), .A2(new_n6708_), .ZN(new_n16819_));
  AOI21_X1   g16627(.A1(new_n16815_), .A2(\asqrt[31] ), .B(new_n16819_), .ZN(new_n16820_));
  NOR2_X1    g16628(.A1(new_n16820_), .A2(new_n16814_), .ZN(new_n16821_));
  AOI22_X1   g16629(.A1(new_n16815_), .A2(\asqrt[31] ), .B1(new_n16813_), .B2(new_n16806_), .ZN(new_n16822_));
  NAND2_X1   g16630(.A1(new_n16490_), .A2(\asqrt[32] ), .ZN(new_n16823_));
  NOR4_X1    g16631(.A1(new_n16619_), .A2(\asqrt[32] ), .A3(new_n16194_), .A4(new_n16490_), .ZN(new_n16824_));
  XOR2_X1    g16632(.A1(new_n16824_), .A2(new_n16823_), .Z(new_n16825_));
  NAND2_X1   g16633(.A1(new_n16825_), .A2(new_n6365_), .ZN(new_n16826_));
  INV_X1     g16634(.I(new_n16826_), .ZN(new_n16827_));
  OAI21_X1   g16635(.A1(new_n16822_), .A2(new_n6708_), .B(new_n16827_), .ZN(new_n16828_));
  NAND2_X1   g16636(.A1(new_n16828_), .A2(new_n16821_), .ZN(new_n16829_));
  OAI22_X1   g16637(.A1(new_n16822_), .A2(new_n6708_), .B1(new_n16820_), .B2(new_n16814_), .ZN(new_n16830_));
  NAND2_X1   g16638(.A1(new_n16206_), .A2(\asqrt[33] ), .ZN(new_n16831_));
  NOR4_X1    g16639(.A1(new_n16619_), .A2(\asqrt[33] ), .A3(new_n16201_), .A4(new_n16206_), .ZN(new_n16832_));
  XOR2_X1    g16640(.A1(new_n16832_), .A2(new_n16831_), .Z(new_n16833_));
  NAND2_X1   g16641(.A1(new_n16833_), .A2(new_n5991_), .ZN(new_n16834_));
  AOI21_X1   g16642(.A1(new_n16830_), .A2(\asqrt[33] ), .B(new_n16834_), .ZN(new_n16835_));
  NOR2_X1    g16643(.A1(new_n16835_), .A2(new_n16829_), .ZN(new_n16836_));
  AOI22_X1   g16644(.A1(new_n16830_), .A2(\asqrt[33] ), .B1(new_n16828_), .B2(new_n16821_), .ZN(new_n16837_));
  NOR4_X1    g16645(.A1(new_n16619_), .A2(\asqrt[34] ), .A3(new_n16209_), .A4(new_n16497_), .ZN(new_n16838_));
  AOI21_X1   g16646(.A1(new_n16831_), .A2(new_n16205_), .B(new_n5991_), .ZN(new_n16839_));
  NOR2_X1    g16647(.A1(new_n16838_), .A2(new_n16839_), .ZN(new_n16840_));
  NAND2_X1   g16648(.A1(new_n16840_), .A2(new_n5626_), .ZN(new_n16841_));
  INV_X1     g16649(.I(new_n16841_), .ZN(new_n16842_));
  OAI21_X1   g16650(.A1(new_n16837_), .A2(new_n5991_), .B(new_n16842_), .ZN(new_n16843_));
  NAND2_X1   g16651(.A1(new_n16843_), .A2(new_n16836_), .ZN(new_n16844_));
  OAI22_X1   g16652(.A1(new_n16837_), .A2(new_n5991_), .B1(new_n16835_), .B2(new_n16829_), .ZN(new_n16845_));
  NAND2_X1   g16653(.A1(new_n16221_), .A2(\asqrt[35] ), .ZN(new_n16846_));
  NOR4_X1    g16654(.A1(new_n16619_), .A2(\asqrt[35] ), .A3(new_n16216_), .A4(new_n16221_), .ZN(new_n16847_));
  XOR2_X1    g16655(.A1(new_n16847_), .A2(new_n16846_), .Z(new_n16848_));
  NAND2_X1   g16656(.A1(new_n16848_), .A2(new_n5273_), .ZN(new_n16849_));
  AOI21_X1   g16657(.A1(new_n16845_), .A2(\asqrt[35] ), .B(new_n16849_), .ZN(new_n16850_));
  NOR2_X1    g16658(.A1(new_n16850_), .A2(new_n16844_), .ZN(new_n16851_));
  AOI22_X1   g16659(.A1(new_n16845_), .A2(\asqrt[35] ), .B1(new_n16843_), .B2(new_n16836_), .ZN(new_n16852_));
  NOR4_X1    g16660(.A1(new_n16619_), .A2(\asqrt[36] ), .A3(new_n16224_), .A4(new_n16504_), .ZN(new_n16853_));
  AOI21_X1   g16661(.A1(new_n16846_), .A2(new_n16220_), .B(new_n5273_), .ZN(new_n16854_));
  NOR2_X1    g16662(.A1(new_n16853_), .A2(new_n16854_), .ZN(new_n16855_));
  NAND2_X1   g16663(.A1(new_n16855_), .A2(new_n4973_), .ZN(new_n16856_));
  INV_X1     g16664(.I(new_n16856_), .ZN(new_n16857_));
  OAI21_X1   g16665(.A1(new_n16852_), .A2(new_n5273_), .B(new_n16857_), .ZN(new_n16858_));
  NAND2_X1   g16666(.A1(new_n16858_), .A2(new_n16851_), .ZN(new_n16859_));
  OAI22_X1   g16667(.A1(new_n16852_), .A2(new_n5273_), .B1(new_n16850_), .B2(new_n16844_), .ZN(new_n16860_));
  NAND2_X1   g16668(.A1(new_n16236_), .A2(\asqrt[37] ), .ZN(new_n16861_));
  NOR4_X1    g16669(.A1(new_n16619_), .A2(\asqrt[37] ), .A3(new_n16231_), .A4(new_n16236_), .ZN(new_n16862_));
  XOR2_X1    g16670(.A1(new_n16862_), .A2(new_n16861_), .Z(new_n16863_));
  NAND2_X1   g16671(.A1(new_n16863_), .A2(new_n4645_), .ZN(new_n16864_));
  AOI21_X1   g16672(.A1(new_n16860_), .A2(\asqrt[37] ), .B(new_n16864_), .ZN(new_n16865_));
  NOR2_X1    g16673(.A1(new_n16865_), .A2(new_n16859_), .ZN(new_n16866_));
  AOI22_X1   g16674(.A1(new_n16860_), .A2(\asqrt[37] ), .B1(new_n16858_), .B2(new_n16851_), .ZN(new_n16867_));
  NOR4_X1    g16675(.A1(new_n16619_), .A2(\asqrt[38] ), .A3(new_n16239_), .A4(new_n16511_), .ZN(new_n16868_));
  AOI21_X1   g16676(.A1(new_n16861_), .A2(new_n16235_), .B(new_n4645_), .ZN(new_n16869_));
  NOR2_X1    g16677(.A1(new_n16868_), .A2(new_n16869_), .ZN(new_n16870_));
  NAND2_X1   g16678(.A1(new_n16870_), .A2(new_n4330_), .ZN(new_n16871_));
  INV_X1     g16679(.I(new_n16871_), .ZN(new_n16872_));
  OAI21_X1   g16680(.A1(new_n16867_), .A2(new_n4645_), .B(new_n16872_), .ZN(new_n16873_));
  NAND2_X1   g16681(.A1(new_n16873_), .A2(new_n16866_), .ZN(new_n16874_));
  OAI22_X1   g16682(.A1(new_n16867_), .A2(new_n4645_), .B1(new_n16865_), .B2(new_n16859_), .ZN(new_n16875_));
  NAND2_X1   g16683(.A1(new_n16251_), .A2(\asqrt[39] ), .ZN(new_n16876_));
  NOR4_X1    g16684(.A1(new_n16619_), .A2(\asqrt[39] ), .A3(new_n16246_), .A4(new_n16251_), .ZN(new_n16877_));
  XOR2_X1    g16685(.A1(new_n16877_), .A2(new_n16876_), .Z(new_n16878_));
  NAND2_X1   g16686(.A1(new_n16878_), .A2(new_n4018_), .ZN(new_n16879_));
  AOI21_X1   g16687(.A1(new_n16875_), .A2(\asqrt[39] ), .B(new_n16879_), .ZN(new_n16880_));
  NOR2_X1    g16688(.A1(new_n16880_), .A2(new_n16874_), .ZN(new_n16881_));
  AOI22_X1   g16689(.A1(new_n16875_), .A2(\asqrt[39] ), .B1(new_n16873_), .B2(new_n16866_), .ZN(new_n16882_));
  NAND2_X1   g16690(.A1(new_n16518_), .A2(\asqrt[40] ), .ZN(new_n16883_));
  NOR4_X1    g16691(.A1(new_n16619_), .A2(\asqrt[40] ), .A3(new_n16254_), .A4(new_n16518_), .ZN(new_n16884_));
  XOR2_X1    g16692(.A1(new_n16884_), .A2(new_n16883_), .Z(new_n16885_));
  NAND2_X1   g16693(.A1(new_n16885_), .A2(new_n3760_), .ZN(new_n16886_));
  INV_X1     g16694(.I(new_n16886_), .ZN(new_n16887_));
  OAI21_X1   g16695(.A1(new_n16882_), .A2(new_n4018_), .B(new_n16887_), .ZN(new_n16888_));
  NAND2_X1   g16696(.A1(new_n16888_), .A2(new_n16881_), .ZN(new_n16889_));
  OAI22_X1   g16697(.A1(new_n16882_), .A2(new_n4018_), .B1(new_n16880_), .B2(new_n16874_), .ZN(new_n16890_));
  NOR4_X1    g16698(.A1(new_n16619_), .A2(\asqrt[41] ), .A3(new_n16261_), .A4(new_n16266_), .ZN(new_n16891_));
  AOI21_X1   g16699(.A1(new_n16883_), .A2(new_n16517_), .B(new_n3760_), .ZN(new_n16892_));
  NOR2_X1    g16700(.A1(new_n16891_), .A2(new_n16892_), .ZN(new_n16893_));
  NAND2_X1   g16701(.A1(new_n16893_), .A2(new_n3481_), .ZN(new_n16894_));
  AOI21_X1   g16702(.A1(new_n16890_), .A2(\asqrt[41] ), .B(new_n16894_), .ZN(new_n16895_));
  NOR2_X1    g16703(.A1(new_n16895_), .A2(new_n16889_), .ZN(new_n16896_));
  AOI22_X1   g16704(.A1(new_n16890_), .A2(\asqrt[41] ), .B1(new_n16888_), .B2(new_n16881_), .ZN(new_n16897_));
  NAND2_X1   g16705(.A1(new_n16525_), .A2(\asqrt[42] ), .ZN(new_n16898_));
  NOR4_X1    g16706(.A1(new_n16619_), .A2(\asqrt[42] ), .A3(new_n16269_), .A4(new_n16525_), .ZN(new_n16899_));
  XOR2_X1    g16707(.A1(new_n16899_), .A2(new_n16898_), .Z(new_n16900_));
  NAND2_X1   g16708(.A1(new_n16900_), .A2(new_n3208_), .ZN(new_n16901_));
  INV_X1     g16709(.I(new_n16901_), .ZN(new_n16902_));
  OAI21_X1   g16710(.A1(new_n16897_), .A2(new_n3481_), .B(new_n16902_), .ZN(new_n16903_));
  NAND2_X1   g16711(.A1(new_n16903_), .A2(new_n16896_), .ZN(new_n16904_));
  OAI22_X1   g16712(.A1(new_n16897_), .A2(new_n3481_), .B1(new_n16895_), .B2(new_n16889_), .ZN(new_n16905_));
  NOR4_X1    g16713(.A1(new_n16619_), .A2(\asqrt[43] ), .A3(new_n16276_), .A4(new_n16281_), .ZN(new_n16906_));
  AOI21_X1   g16714(.A1(new_n16898_), .A2(new_n16524_), .B(new_n3208_), .ZN(new_n16907_));
  NOR2_X1    g16715(.A1(new_n16906_), .A2(new_n16907_), .ZN(new_n16908_));
  NAND2_X1   g16716(.A1(new_n16908_), .A2(new_n2941_), .ZN(new_n16909_));
  AOI21_X1   g16717(.A1(new_n16905_), .A2(\asqrt[43] ), .B(new_n16909_), .ZN(new_n16910_));
  NOR2_X1    g16718(.A1(new_n16910_), .A2(new_n16904_), .ZN(new_n16911_));
  AOI22_X1   g16719(.A1(new_n16905_), .A2(\asqrt[43] ), .B1(new_n16903_), .B2(new_n16896_), .ZN(new_n16912_));
  NAND2_X1   g16720(.A1(new_n16532_), .A2(\asqrt[44] ), .ZN(new_n16913_));
  NOR4_X1    g16721(.A1(new_n16619_), .A2(\asqrt[44] ), .A3(new_n16284_), .A4(new_n16532_), .ZN(new_n16914_));
  XOR2_X1    g16722(.A1(new_n16914_), .A2(new_n16913_), .Z(new_n16915_));
  NAND2_X1   g16723(.A1(new_n16915_), .A2(new_n2728_), .ZN(new_n16916_));
  INV_X1     g16724(.I(new_n16916_), .ZN(new_n16917_));
  OAI21_X1   g16725(.A1(new_n16912_), .A2(new_n2941_), .B(new_n16917_), .ZN(new_n16918_));
  NAND2_X1   g16726(.A1(new_n16918_), .A2(new_n16911_), .ZN(new_n16919_));
  OAI22_X1   g16727(.A1(new_n16912_), .A2(new_n2941_), .B1(new_n16910_), .B2(new_n16904_), .ZN(new_n16920_));
  NAND2_X1   g16728(.A1(new_n16296_), .A2(\asqrt[45] ), .ZN(new_n16921_));
  NOR4_X1    g16729(.A1(new_n16619_), .A2(\asqrt[45] ), .A3(new_n16291_), .A4(new_n16296_), .ZN(new_n16922_));
  XOR2_X1    g16730(.A1(new_n16922_), .A2(new_n16921_), .Z(new_n16923_));
  NAND2_X1   g16731(.A1(new_n16923_), .A2(new_n2488_), .ZN(new_n16924_));
  AOI21_X1   g16732(.A1(new_n16920_), .A2(\asqrt[45] ), .B(new_n16924_), .ZN(new_n16925_));
  NOR2_X1    g16733(.A1(new_n16925_), .A2(new_n16919_), .ZN(new_n16926_));
  AOI22_X1   g16734(.A1(new_n16920_), .A2(\asqrt[45] ), .B1(new_n16918_), .B2(new_n16911_), .ZN(new_n16927_));
  NOR4_X1    g16735(.A1(new_n16619_), .A2(\asqrt[46] ), .A3(new_n16299_), .A4(new_n16539_), .ZN(new_n16928_));
  AOI21_X1   g16736(.A1(new_n16921_), .A2(new_n16295_), .B(new_n2488_), .ZN(new_n16929_));
  NOR2_X1    g16737(.A1(new_n16928_), .A2(new_n16929_), .ZN(new_n16930_));
  NAND2_X1   g16738(.A1(new_n16930_), .A2(new_n2253_), .ZN(new_n16931_));
  INV_X1     g16739(.I(new_n16931_), .ZN(new_n16932_));
  OAI21_X1   g16740(.A1(new_n16927_), .A2(new_n2488_), .B(new_n16932_), .ZN(new_n16933_));
  NAND2_X1   g16741(.A1(new_n16933_), .A2(new_n16926_), .ZN(new_n16934_));
  OAI22_X1   g16742(.A1(new_n16927_), .A2(new_n2488_), .B1(new_n16925_), .B2(new_n16919_), .ZN(new_n16935_));
  NAND2_X1   g16743(.A1(new_n16311_), .A2(\asqrt[47] ), .ZN(new_n16936_));
  NOR4_X1    g16744(.A1(new_n16619_), .A2(\asqrt[47] ), .A3(new_n16306_), .A4(new_n16311_), .ZN(new_n16937_));
  XOR2_X1    g16745(.A1(new_n16937_), .A2(new_n16936_), .Z(new_n16938_));
  NAND2_X1   g16746(.A1(new_n16938_), .A2(new_n2046_), .ZN(new_n16939_));
  AOI21_X1   g16747(.A1(new_n16935_), .A2(\asqrt[47] ), .B(new_n16939_), .ZN(new_n16940_));
  NOR2_X1    g16748(.A1(new_n16940_), .A2(new_n16934_), .ZN(new_n16941_));
  AOI22_X1   g16749(.A1(new_n16935_), .A2(\asqrt[47] ), .B1(new_n16933_), .B2(new_n16926_), .ZN(new_n16942_));
  NOR4_X1    g16750(.A1(new_n16619_), .A2(\asqrt[48] ), .A3(new_n16314_), .A4(new_n16546_), .ZN(new_n16943_));
  AOI21_X1   g16751(.A1(new_n16936_), .A2(new_n16310_), .B(new_n2046_), .ZN(new_n16944_));
  NOR2_X1    g16752(.A1(new_n16943_), .A2(new_n16944_), .ZN(new_n16945_));
  NAND2_X1   g16753(.A1(new_n16945_), .A2(new_n1854_), .ZN(new_n16946_));
  INV_X1     g16754(.I(new_n16946_), .ZN(new_n16947_));
  OAI21_X1   g16755(.A1(new_n16942_), .A2(new_n2046_), .B(new_n16947_), .ZN(new_n16948_));
  NAND2_X1   g16756(.A1(new_n16948_), .A2(new_n16941_), .ZN(new_n16949_));
  OAI22_X1   g16757(.A1(new_n16942_), .A2(new_n2046_), .B1(new_n16940_), .B2(new_n16934_), .ZN(new_n16950_));
  NAND2_X1   g16758(.A1(new_n16326_), .A2(\asqrt[49] ), .ZN(new_n16951_));
  NOR4_X1    g16759(.A1(new_n16619_), .A2(\asqrt[49] ), .A3(new_n16321_), .A4(new_n16326_), .ZN(new_n16952_));
  XOR2_X1    g16760(.A1(new_n16952_), .A2(new_n16951_), .Z(new_n16953_));
  NAND2_X1   g16761(.A1(new_n16953_), .A2(new_n1595_), .ZN(new_n16954_));
  AOI21_X1   g16762(.A1(new_n16950_), .A2(\asqrt[49] ), .B(new_n16954_), .ZN(new_n16955_));
  NOR2_X1    g16763(.A1(new_n16955_), .A2(new_n16949_), .ZN(new_n16956_));
  AOI22_X1   g16764(.A1(new_n16950_), .A2(\asqrt[49] ), .B1(new_n16948_), .B2(new_n16941_), .ZN(new_n16957_));
  NOR4_X1    g16765(.A1(new_n16619_), .A2(\asqrt[50] ), .A3(new_n16329_), .A4(new_n16553_), .ZN(new_n16958_));
  AOI21_X1   g16766(.A1(new_n16951_), .A2(new_n16325_), .B(new_n1595_), .ZN(new_n16959_));
  NOR2_X1    g16767(.A1(new_n16958_), .A2(new_n16959_), .ZN(new_n16960_));
  NAND2_X1   g16768(.A1(new_n16960_), .A2(new_n1436_), .ZN(new_n16961_));
  INV_X1     g16769(.I(new_n16961_), .ZN(new_n16962_));
  OAI21_X1   g16770(.A1(new_n16957_), .A2(new_n1595_), .B(new_n16962_), .ZN(new_n16963_));
  NAND2_X1   g16771(.A1(new_n16963_), .A2(new_n16956_), .ZN(new_n16964_));
  OAI22_X1   g16772(.A1(new_n16957_), .A2(new_n1595_), .B1(new_n16955_), .B2(new_n16949_), .ZN(new_n16965_));
  NAND2_X1   g16773(.A1(new_n16341_), .A2(\asqrt[51] ), .ZN(new_n16966_));
  NOR4_X1    g16774(.A1(new_n16619_), .A2(\asqrt[51] ), .A3(new_n16336_), .A4(new_n16341_), .ZN(new_n16967_));
  XOR2_X1    g16775(.A1(new_n16967_), .A2(new_n16966_), .Z(new_n16968_));
  NAND2_X1   g16776(.A1(new_n16968_), .A2(new_n1260_), .ZN(new_n16969_));
  AOI21_X1   g16777(.A1(new_n16965_), .A2(\asqrt[51] ), .B(new_n16969_), .ZN(new_n16970_));
  NOR2_X1    g16778(.A1(new_n16970_), .A2(new_n16964_), .ZN(new_n16971_));
  AOI22_X1   g16779(.A1(new_n16965_), .A2(\asqrt[51] ), .B1(new_n16963_), .B2(new_n16956_), .ZN(new_n16972_));
  NAND2_X1   g16780(.A1(new_n16560_), .A2(\asqrt[52] ), .ZN(new_n16973_));
  NOR4_X1    g16781(.A1(new_n16619_), .A2(\asqrt[52] ), .A3(new_n16344_), .A4(new_n16560_), .ZN(new_n16974_));
  XOR2_X1    g16782(.A1(new_n16974_), .A2(new_n16973_), .Z(new_n16975_));
  NAND2_X1   g16783(.A1(new_n16975_), .A2(new_n1096_), .ZN(new_n16976_));
  INV_X1     g16784(.I(new_n16976_), .ZN(new_n16977_));
  OAI21_X1   g16785(.A1(new_n16972_), .A2(new_n1260_), .B(new_n16977_), .ZN(new_n16978_));
  NAND2_X1   g16786(.A1(new_n16978_), .A2(new_n16971_), .ZN(new_n16979_));
  OAI22_X1   g16787(.A1(new_n16972_), .A2(new_n1260_), .B1(new_n16970_), .B2(new_n16964_), .ZN(new_n16980_));
  NOR4_X1    g16788(.A1(new_n16619_), .A2(\asqrt[53] ), .A3(new_n16351_), .A4(new_n16356_), .ZN(new_n16981_));
  AOI21_X1   g16789(.A1(new_n16973_), .A2(new_n16559_), .B(new_n1096_), .ZN(new_n16982_));
  NOR2_X1    g16790(.A1(new_n16981_), .A2(new_n16982_), .ZN(new_n16983_));
  NAND2_X1   g16791(.A1(new_n16983_), .A2(new_n970_), .ZN(new_n16984_));
  AOI21_X1   g16792(.A1(new_n16980_), .A2(\asqrt[53] ), .B(new_n16984_), .ZN(new_n16985_));
  NOR2_X1    g16793(.A1(new_n16985_), .A2(new_n16979_), .ZN(new_n16986_));
  AOI22_X1   g16794(.A1(new_n16980_), .A2(\asqrt[53] ), .B1(new_n16978_), .B2(new_n16971_), .ZN(new_n16987_));
  NOR4_X1    g16795(.A1(new_n16619_), .A2(\asqrt[54] ), .A3(new_n16359_), .A4(new_n16567_), .ZN(new_n16988_));
  XOR2_X1    g16796(.A1(new_n16988_), .A2(new_n16635_), .Z(new_n16989_));
  NAND2_X1   g16797(.A1(new_n16989_), .A2(new_n825_), .ZN(new_n16990_));
  INV_X1     g16798(.I(new_n16990_), .ZN(new_n16991_));
  OAI21_X1   g16799(.A1(new_n16987_), .A2(new_n970_), .B(new_n16991_), .ZN(new_n16992_));
  NAND2_X1   g16800(.A1(new_n16992_), .A2(new_n16986_), .ZN(new_n16993_));
  OAI22_X1   g16801(.A1(new_n16987_), .A2(new_n970_), .B1(new_n16985_), .B2(new_n16979_), .ZN(new_n16994_));
  NOR4_X1    g16802(.A1(new_n16619_), .A2(\asqrt[55] ), .A3(new_n16365_), .A4(new_n16370_), .ZN(new_n16995_));
  XOR2_X1    g16803(.A1(new_n16995_), .A2(new_n16620_), .Z(new_n16996_));
  NAND2_X1   g16804(.A1(new_n16996_), .A2(new_n724_), .ZN(new_n16997_));
  AOI21_X1   g16805(.A1(new_n16994_), .A2(\asqrt[55] ), .B(new_n16997_), .ZN(new_n16998_));
  NOR2_X1    g16806(.A1(new_n16998_), .A2(new_n16993_), .ZN(new_n16999_));
  AOI22_X1   g16807(.A1(new_n16994_), .A2(\asqrt[55] ), .B1(new_n16992_), .B2(new_n16986_), .ZN(new_n17000_));
  NOR4_X1    g16808(.A1(new_n16619_), .A2(\asqrt[56] ), .A3(new_n16372_), .A4(new_n16574_), .ZN(new_n17001_));
  XOR2_X1    g16809(.A1(new_n17001_), .A2(new_n16637_), .Z(new_n17002_));
  NAND2_X1   g16810(.A1(new_n17002_), .A2(new_n587_), .ZN(new_n17003_));
  INV_X1     g16811(.I(new_n17003_), .ZN(new_n17004_));
  OAI21_X1   g16812(.A1(new_n17000_), .A2(new_n724_), .B(new_n17004_), .ZN(new_n17005_));
  NAND2_X1   g16813(.A1(new_n17005_), .A2(new_n16999_), .ZN(new_n17006_));
  OAI22_X1   g16814(.A1(new_n17000_), .A2(new_n724_), .B1(new_n16998_), .B2(new_n16993_), .ZN(new_n17007_));
  NOR4_X1    g16815(.A1(new_n16619_), .A2(\asqrt[57] ), .A3(new_n16378_), .A4(new_n16383_), .ZN(new_n17008_));
  XOR2_X1    g16816(.A1(new_n17008_), .A2(new_n16622_), .Z(new_n17009_));
  NAND2_X1   g16817(.A1(new_n17009_), .A2(new_n504_), .ZN(new_n17010_));
  AOI21_X1   g16818(.A1(new_n17007_), .A2(\asqrt[57] ), .B(new_n17010_), .ZN(new_n17011_));
  NOR2_X1    g16819(.A1(new_n17011_), .A2(new_n17006_), .ZN(new_n17012_));
  AOI22_X1   g16820(.A1(new_n17007_), .A2(\asqrt[57] ), .B1(new_n17005_), .B2(new_n16999_), .ZN(new_n17013_));
  NOR4_X1    g16821(.A1(new_n16619_), .A2(\asqrt[58] ), .A3(new_n16385_), .A4(new_n16581_), .ZN(new_n17014_));
  XOR2_X1    g16822(.A1(new_n17014_), .A2(new_n16639_), .Z(new_n17015_));
  NAND2_X1   g16823(.A1(new_n17015_), .A2(new_n376_), .ZN(new_n17016_));
  INV_X1     g16824(.I(new_n17016_), .ZN(new_n17017_));
  OAI21_X1   g16825(.A1(new_n17013_), .A2(new_n504_), .B(new_n17017_), .ZN(new_n17018_));
  NAND2_X1   g16826(.A1(new_n17018_), .A2(new_n17012_), .ZN(new_n17019_));
  NAND2_X1   g16827(.A1(new_n16980_), .A2(\asqrt[53] ), .ZN(new_n17020_));
  AOI21_X1   g16828(.A1(new_n17020_), .A2(new_n16979_), .B(new_n970_), .ZN(new_n17021_));
  OAI21_X1   g16829(.A1(new_n16986_), .A2(new_n17021_), .B(\asqrt[55] ), .ZN(new_n17022_));
  AOI21_X1   g16830(.A1(new_n16993_), .A2(new_n17022_), .B(new_n724_), .ZN(new_n17023_));
  OAI21_X1   g16831(.A1(new_n16999_), .A2(new_n17023_), .B(\asqrt[57] ), .ZN(new_n17024_));
  AOI21_X1   g16832(.A1(new_n17006_), .A2(new_n17024_), .B(new_n504_), .ZN(new_n17025_));
  OAI21_X1   g16833(.A1(new_n17012_), .A2(new_n17025_), .B(\asqrt[59] ), .ZN(new_n17026_));
  NOR4_X1    g16834(.A1(new_n16619_), .A2(\asqrt[59] ), .A3(new_n16391_), .A4(new_n16396_), .ZN(new_n17027_));
  XOR2_X1    g16835(.A1(new_n17027_), .A2(new_n16624_), .Z(new_n17028_));
  AND2_X2    g16836(.A1(new_n17028_), .A2(new_n275_), .Z(new_n17029_));
  AOI21_X1   g16837(.A1(new_n17026_), .A2(new_n17029_), .B(new_n17019_), .ZN(new_n17030_));
  OAI22_X1   g16838(.A1(new_n17013_), .A2(new_n504_), .B1(new_n17011_), .B2(new_n17006_), .ZN(new_n17031_));
  AOI22_X1   g16839(.A1(new_n17031_), .A2(\asqrt[59] ), .B1(new_n17018_), .B2(new_n17012_), .ZN(new_n17032_));
  NOR4_X1    g16840(.A1(new_n16619_), .A2(\asqrt[60] ), .A3(new_n16398_), .A4(new_n16588_), .ZN(new_n17033_));
  XOR2_X1    g16841(.A1(new_n17033_), .A2(new_n16641_), .Z(new_n17034_));
  NAND2_X1   g16842(.A1(new_n17034_), .A2(new_n229_), .ZN(new_n17035_));
  INV_X1     g16843(.I(new_n17035_), .ZN(new_n17036_));
  OAI21_X1   g16844(.A1(new_n17032_), .A2(new_n275_), .B(new_n17036_), .ZN(new_n17037_));
  OAI22_X1   g16845(.A1(new_n16662_), .A2(new_n14871_), .B1(new_n16650_), .B2(new_n16660_), .ZN(new_n17038_));
  AOI22_X1   g16846(.A1(new_n17038_), .A2(\asqrt[16] ), .B1(new_n16671_), .B2(new_n16661_), .ZN(new_n17039_));
  INV_X1     g16847(.I(new_n16706_), .ZN(new_n17040_));
  OAI21_X1   g16848(.A1(new_n17039_), .A2(new_n13760_), .B(new_n17040_), .ZN(new_n17041_));
  AOI21_X1   g16849(.A1(new_n17038_), .A2(\asqrt[16] ), .B(new_n16679_), .ZN(new_n17042_));
  OAI22_X1   g16850(.A1(new_n17039_), .A2(new_n13760_), .B1(new_n17042_), .B2(new_n16709_), .ZN(new_n17043_));
  AOI22_X1   g16851(.A1(new_n17043_), .A2(\asqrt[18] ), .B1(new_n17041_), .B2(new_n16710_), .ZN(new_n17044_));
  INV_X1     g16852(.I(new_n16725_), .ZN(new_n17045_));
  OAI21_X1   g16853(.A1(new_n17044_), .A2(new_n12657_), .B(new_n17045_), .ZN(new_n17046_));
  NAND2_X1   g16854(.A1(new_n17046_), .A2(new_n16729_), .ZN(new_n17047_));
  AOI21_X1   g16855(.A1(new_n17043_), .A2(\asqrt[18] ), .B(new_n16716_), .ZN(new_n17048_));
  OAI22_X1   g16856(.A1(new_n17044_), .A2(new_n12657_), .B1(new_n17048_), .B2(new_n16728_), .ZN(new_n17049_));
  AOI21_X1   g16857(.A1(new_n17049_), .A2(\asqrt[20] ), .B(new_n16735_), .ZN(new_n17050_));
  NOR2_X1    g16858(.A1(new_n17050_), .A2(new_n17047_), .ZN(new_n17051_));
  AOI22_X1   g16859(.A1(new_n17049_), .A2(\asqrt[20] ), .B1(new_n17046_), .B2(new_n16729_), .ZN(new_n17052_));
  INV_X1     g16860(.I(new_n16744_), .ZN(new_n17053_));
  OAI21_X1   g16861(.A1(new_n17052_), .A2(new_n11631_), .B(new_n17053_), .ZN(new_n17054_));
  NAND2_X1   g16862(.A1(new_n17054_), .A2(new_n17051_), .ZN(new_n17055_));
  OAI22_X1   g16863(.A1(new_n17052_), .A2(new_n11631_), .B1(new_n17050_), .B2(new_n17047_), .ZN(new_n17056_));
  AOI21_X1   g16864(.A1(new_n17056_), .A2(\asqrt[22] ), .B(new_n16751_), .ZN(new_n17057_));
  NOR2_X1    g16865(.A1(new_n17057_), .A2(new_n17055_), .ZN(new_n17058_));
  AOI22_X1   g16866(.A1(new_n17056_), .A2(\asqrt[22] ), .B1(new_n17054_), .B2(new_n17051_), .ZN(new_n17059_));
  INV_X1     g16867(.I(new_n16759_), .ZN(new_n17060_));
  OAI21_X1   g16868(.A1(new_n17059_), .A2(new_n10614_), .B(new_n17060_), .ZN(new_n17061_));
  NAND2_X1   g16869(.A1(new_n17061_), .A2(new_n17058_), .ZN(new_n17062_));
  OAI22_X1   g16870(.A1(new_n17059_), .A2(new_n10614_), .B1(new_n17057_), .B2(new_n17055_), .ZN(new_n17063_));
  AOI21_X1   g16871(.A1(new_n17063_), .A2(\asqrt[24] ), .B(new_n16766_), .ZN(new_n17064_));
  NOR2_X1    g16872(.A1(new_n17064_), .A2(new_n17062_), .ZN(new_n17065_));
  AOI22_X1   g16873(.A1(new_n17063_), .A2(\asqrt[24] ), .B1(new_n17061_), .B2(new_n17058_), .ZN(new_n17066_));
  INV_X1     g16874(.I(new_n16774_), .ZN(new_n17067_));
  OAI21_X1   g16875(.A1(new_n17066_), .A2(new_n9672_), .B(new_n17067_), .ZN(new_n17068_));
  NAND2_X1   g16876(.A1(new_n17068_), .A2(new_n17065_), .ZN(new_n17069_));
  OAI22_X1   g16877(.A1(new_n17066_), .A2(new_n9672_), .B1(new_n17064_), .B2(new_n17062_), .ZN(new_n17070_));
  AOI21_X1   g16878(.A1(new_n17070_), .A2(\asqrt[26] ), .B(new_n16781_), .ZN(new_n17071_));
  NOR2_X1    g16879(.A1(new_n17071_), .A2(new_n17069_), .ZN(new_n17072_));
  AOI22_X1   g16880(.A1(new_n17070_), .A2(\asqrt[26] ), .B1(new_n17068_), .B2(new_n17065_), .ZN(new_n17073_));
  INV_X1     g16881(.I(new_n16789_), .ZN(new_n17074_));
  OAI21_X1   g16882(.A1(new_n17073_), .A2(new_n8763_), .B(new_n17074_), .ZN(new_n17075_));
  NAND2_X1   g16883(.A1(new_n17075_), .A2(new_n17072_), .ZN(new_n17076_));
  OAI22_X1   g16884(.A1(new_n17073_), .A2(new_n8763_), .B1(new_n17071_), .B2(new_n17069_), .ZN(new_n17077_));
  AOI21_X1   g16885(.A1(new_n17077_), .A2(\asqrt[28] ), .B(new_n16796_), .ZN(new_n17078_));
  NOR2_X1    g16886(.A1(new_n17078_), .A2(new_n17076_), .ZN(new_n17079_));
  AOI22_X1   g16887(.A1(new_n17077_), .A2(\asqrt[28] ), .B1(new_n17075_), .B2(new_n17072_), .ZN(new_n17080_));
  INV_X1     g16888(.I(new_n16804_), .ZN(new_n17081_));
  OAI21_X1   g16889(.A1(new_n17080_), .A2(new_n7931_), .B(new_n17081_), .ZN(new_n17082_));
  NAND2_X1   g16890(.A1(new_n17082_), .A2(new_n17079_), .ZN(new_n17083_));
  OAI22_X1   g16891(.A1(new_n17080_), .A2(new_n7931_), .B1(new_n17078_), .B2(new_n17076_), .ZN(new_n17084_));
  AOI21_X1   g16892(.A1(new_n17084_), .A2(\asqrt[30] ), .B(new_n16811_), .ZN(new_n17085_));
  NOR2_X1    g16893(.A1(new_n17085_), .A2(new_n17083_), .ZN(new_n17086_));
  AOI22_X1   g16894(.A1(new_n17084_), .A2(\asqrt[30] ), .B1(new_n17082_), .B2(new_n17079_), .ZN(new_n17087_));
  INV_X1     g16895(.I(new_n16819_), .ZN(new_n17088_));
  OAI21_X1   g16896(.A1(new_n17087_), .A2(new_n7110_), .B(new_n17088_), .ZN(new_n17089_));
  NAND2_X1   g16897(.A1(new_n17089_), .A2(new_n17086_), .ZN(new_n17090_));
  OAI22_X1   g16898(.A1(new_n17087_), .A2(new_n7110_), .B1(new_n17085_), .B2(new_n17083_), .ZN(new_n17091_));
  AOI21_X1   g16899(.A1(new_n17091_), .A2(\asqrt[32] ), .B(new_n16826_), .ZN(new_n17092_));
  NOR2_X1    g16900(.A1(new_n17092_), .A2(new_n17090_), .ZN(new_n17093_));
  AOI22_X1   g16901(.A1(new_n17091_), .A2(\asqrt[32] ), .B1(new_n17089_), .B2(new_n17086_), .ZN(new_n17094_));
  INV_X1     g16902(.I(new_n16834_), .ZN(new_n17095_));
  OAI21_X1   g16903(.A1(new_n17094_), .A2(new_n6365_), .B(new_n17095_), .ZN(new_n17096_));
  NAND2_X1   g16904(.A1(new_n17096_), .A2(new_n17093_), .ZN(new_n17097_));
  OAI22_X1   g16905(.A1(new_n17094_), .A2(new_n6365_), .B1(new_n17092_), .B2(new_n17090_), .ZN(new_n17098_));
  AOI21_X1   g16906(.A1(new_n17098_), .A2(\asqrt[34] ), .B(new_n16841_), .ZN(new_n17099_));
  NOR2_X1    g16907(.A1(new_n17099_), .A2(new_n17097_), .ZN(new_n17100_));
  AOI22_X1   g16908(.A1(new_n17098_), .A2(\asqrt[34] ), .B1(new_n17096_), .B2(new_n17093_), .ZN(new_n17101_));
  INV_X1     g16909(.I(new_n16849_), .ZN(new_n17102_));
  OAI21_X1   g16910(.A1(new_n17101_), .A2(new_n5626_), .B(new_n17102_), .ZN(new_n17103_));
  NAND2_X1   g16911(.A1(new_n17103_), .A2(new_n17100_), .ZN(new_n17104_));
  OAI22_X1   g16912(.A1(new_n17101_), .A2(new_n5626_), .B1(new_n17099_), .B2(new_n17097_), .ZN(new_n17105_));
  AOI21_X1   g16913(.A1(new_n17105_), .A2(\asqrt[36] ), .B(new_n16856_), .ZN(new_n17106_));
  NOR2_X1    g16914(.A1(new_n17106_), .A2(new_n17104_), .ZN(new_n17107_));
  AOI22_X1   g16915(.A1(new_n17105_), .A2(\asqrt[36] ), .B1(new_n17103_), .B2(new_n17100_), .ZN(new_n17108_));
  INV_X1     g16916(.I(new_n16864_), .ZN(new_n17109_));
  OAI21_X1   g16917(.A1(new_n17108_), .A2(new_n4973_), .B(new_n17109_), .ZN(new_n17110_));
  NAND2_X1   g16918(.A1(new_n17110_), .A2(new_n17107_), .ZN(new_n17111_));
  OAI22_X1   g16919(.A1(new_n17108_), .A2(new_n4973_), .B1(new_n17106_), .B2(new_n17104_), .ZN(new_n17112_));
  AOI21_X1   g16920(.A1(new_n17112_), .A2(\asqrt[38] ), .B(new_n16871_), .ZN(new_n17113_));
  NOR2_X1    g16921(.A1(new_n17113_), .A2(new_n17111_), .ZN(new_n17114_));
  AOI22_X1   g16922(.A1(new_n17112_), .A2(\asqrt[38] ), .B1(new_n17110_), .B2(new_n17107_), .ZN(new_n17115_));
  INV_X1     g16923(.I(new_n16879_), .ZN(new_n17116_));
  OAI21_X1   g16924(.A1(new_n17115_), .A2(new_n4330_), .B(new_n17116_), .ZN(new_n17117_));
  NAND2_X1   g16925(.A1(new_n17117_), .A2(new_n17114_), .ZN(new_n17118_));
  OAI22_X1   g16926(.A1(new_n17115_), .A2(new_n4330_), .B1(new_n17113_), .B2(new_n17111_), .ZN(new_n17119_));
  AOI21_X1   g16927(.A1(new_n17119_), .A2(\asqrt[40] ), .B(new_n16886_), .ZN(new_n17120_));
  NOR2_X1    g16928(.A1(new_n17120_), .A2(new_n17118_), .ZN(new_n17121_));
  AOI22_X1   g16929(.A1(new_n17119_), .A2(\asqrt[40] ), .B1(new_n17117_), .B2(new_n17114_), .ZN(new_n17122_));
  INV_X1     g16930(.I(new_n16894_), .ZN(new_n17123_));
  OAI21_X1   g16931(.A1(new_n17122_), .A2(new_n3760_), .B(new_n17123_), .ZN(new_n17124_));
  NAND2_X1   g16932(.A1(new_n17124_), .A2(new_n17121_), .ZN(new_n17125_));
  OAI22_X1   g16933(.A1(new_n17122_), .A2(new_n3760_), .B1(new_n17120_), .B2(new_n17118_), .ZN(new_n17126_));
  AOI21_X1   g16934(.A1(new_n17126_), .A2(\asqrt[42] ), .B(new_n16901_), .ZN(new_n17127_));
  NOR2_X1    g16935(.A1(new_n17127_), .A2(new_n17125_), .ZN(new_n17128_));
  AOI22_X1   g16936(.A1(new_n17126_), .A2(\asqrt[42] ), .B1(new_n17124_), .B2(new_n17121_), .ZN(new_n17129_));
  INV_X1     g16937(.I(new_n16909_), .ZN(new_n17130_));
  OAI21_X1   g16938(.A1(new_n17129_), .A2(new_n3208_), .B(new_n17130_), .ZN(new_n17131_));
  NAND2_X1   g16939(.A1(new_n17131_), .A2(new_n17128_), .ZN(new_n17132_));
  OAI22_X1   g16940(.A1(new_n17129_), .A2(new_n3208_), .B1(new_n17127_), .B2(new_n17125_), .ZN(new_n17133_));
  AOI21_X1   g16941(.A1(new_n17133_), .A2(\asqrt[44] ), .B(new_n16916_), .ZN(new_n17134_));
  NOR2_X1    g16942(.A1(new_n17134_), .A2(new_n17132_), .ZN(new_n17135_));
  AOI22_X1   g16943(.A1(new_n17133_), .A2(\asqrt[44] ), .B1(new_n17131_), .B2(new_n17128_), .ZN(new_n17136_));
  INV_X1     g16944(.I(new_n16924_), .ZN(new_n17137_));
  OAI21_X1   g16945(.A1(new_n17136_), .A2(new_n2728_), .B(new_n17137_), .ZN(new_n17138_));
  NAND2_X1   g16946(.A1(new_n17138_), .A2(new_n17135_), .ZN(new_n17139_));
  OAI22_X1   g16947(.A1(new_n17136_), .A2(new_n2728_), .B1(new_n17134_), .B2(new_n17132_), .ZN(new_n17140_));
  AOI21_X1   g16948(.A1(new_n17140_), .A2(\asqrt[46] ), .B(new_n16931_), .ZN(new_n17141_));
  NOR2_X1    g16949(.A1(new_n17141_), .A2(new_n17139_), .ZN(new_n17142_));
  AOI22_X1   g16950(.A1(new_n17140_), .A2(\asqrt[46] ), .B1(new_n17138_), .B2(new_n17135_), .ZN(new_n17143_));
  INV_X1     g16951(.I(new_n16939_), .ZN(new_n17144_));
  OAI21_X1   g16952(.A1(new_n17143_), .A2(new_n2253_), .B(new_n17144_), .ZN(new_n17145_));
  NAND2_X1   g16953(.A1(new_n17145_), .A2(new_n17142_), .ZN(new_n17146_));
  OAI22_X1   g16954(.A1(new_n17143_), .A2(new_n2253_), .B1(new_n17141_), .B2(new_n17139_), .ZN(new_n17147_));
  AOI21_X1   g16955(.A1(new_n17147_), .A2(\asqrt[48] ), .B(new_n16946_), .ZN(new_n17148_));
  NOR2_X1    g16956(.A1(new_n17148_), .A2(new_n17146_), .ZN(new_n17149_));
  AOI22_X1   g16957(.A1(new_n17147_), .A2(\asqrt[48] ), .B1(new_n17145_), .B2(new_n17142_), .ZN(new_n17150_));
  INV_X1     g16958(.I(new_n16954_), .ZN(new_n17151_));
  OAI21_X1   g16959(.A1(new_n17150_), .A2(new_n1854_), .B(new_n17151_), .ZN(new_n17152_));
  NAND2_X1   g16960(.A1(new_n17152_), .A2(new_n17149_), .ZN(new_n17153_));
  OAI22_X1   g16961(.A1(new_n17150_), .A2(new_n1854_), .B1(new_n17148_), .B2(new_n17146_), .ZN(new_n17154_));
  AOI21_X1   g16962(.A1(new_n17154_), .A2(\asqrt[50] ), .B(new_n16961_), .ZN(new_n17155_));
  NOR2_X1    g16963(.A1(new_n17155_), .A2(new_n17153_), .ZN(new_n17156_));
  AOI22_X1   g16964(.A1(new_n17154_), .A2(\asqrt[50] ), .B1(new_n17152_), .B2(new_n17149_), .ZN(new_n17157_));
  INV_X1     g16965(.I(new_n16969_), .ZN(new_n17158_));
  OAI21_X1   g16966(.A1(new_n17157_), .A2(new_n1436_), .B(new_n17158_), .ZN(new_n17159_));
  NAND2_X1   g16967(.A1(new_n17159_), .A2(new_n17156_), .ZN(new_n17160_));
  OAI22_X1   g16968(.A1(new_n17157_), .A2(new_n1436_), .B1(new_n17155_), .B2(new_n17153_), .ZN(new_n17161_));
  AOI21_X1   g16969(.A1(new_n17161_), .A2(\asqrt[52] ), .B(new_n16976_), .ZN(new_n17162_));
  NOR2_X1    g16970(.A1(new_n17162_), .A2(new_n17160_), .ZN(new_n17163_));
  AOI22_X1   g16971(.A1(new_n17161_), .A2(\asqrt[52] ), .B1(new_n17159_), .B2(new_n17156_), .ZN(new_n17164_));
  INV_X1     g16972(.I(new_n16984_), .ZN(new_n17165_));
  OAI21_X1   g16973(.A1(new_n17164_), .A2(new_n1096_), .B(new_n17165_), .ZN(new_n17166_));
  NAND2_X1   g16974(.A1(new_n17166_), .A2(new_n17163_), .ZN(new_n17167_));
  OAI22_X1   g16975(.A1(new_n17164_), .A2(new_n1096_), .B1(new_n17162_), .B2(new_n17160_), .ZN(new_n17168_));
  AOI21_X1   g16976(.A1(new_n17168_), .A2(\asqrt[54] ), .B(new_n16990_), .ZN(new_n17169_));
  NOR2_X1    g16977(.A1(new_n17169_), .A2(new_n17167_), .ZN(new_n17170_));
  AOI22_X1   g16978(.A1(new_n17168_), .A2(\asqrt[54] ), .B1(new_n17166_), .B2(new_n17163_), .ZN(new_n17171_));
  INV_X1     g16979(.I(new_n16997_), .ZN(new_n17172_));
  OAI21_X1   g16980(.A1(new_n17171_), .A2(new_n825_), .B(new_n17172_), .ZN(new_n17173_));
  NAND2_X1   g16981(.A1(new_n17173_), .A2(new_n17170_), .ZN(new_n17174_));
  OAI22_X1   g16982(.A1(new_n17171_), .A2(new_n825_), .B1(new_n17169_), .B2(new_n17167_), .ZN(new_n17175_));
  AOI21_X1   g16983(.A1(new_n17175_), .A2(\asqrt[56] ), .B(new_n17003_), .ZN(new_n17176_));
  NOR2_X1    g16984(.A1(new_n17176_), .A2(new_n17174_), .ZN(new_n17177_));
  AOI22_X1   g16985(.A1(new_n17175_), .A2(\asqrt[56] ), .B1(new_n17173_), .B2(new_n17170_), .ZN(new_n17178_));
  INV_X1     g16986(.I(new_n17010_), .ZN(new_n17179_));
  OAI21_X1   g16987(.A1(new_n17178_), .A2(new_n587_), .B(new_n17179_), .ZN(new_n17180_));
  NAND2_X1   g16988(.A1(new_n17180_), .A2(new_n17177_), .ZN(new_n17181_));
  OAI22_X1   g16989(.A1(new_n17178_), .A2(new_n587_), .B1(new_n17176_), .B2(new_n17174_), .ZN(new_n17182_));
  AOI21_X1   g16990(.A1(new_n17182_), .A2(\asqrt[58] ), .B(new_n17016_), .ZN(new_n17183_));
  NOR2_X1    g16991(.A1(new_n17183_), .A2(new_n17181_), .ZN(new_n17184_));
  AOI22_X1   g16992(.A1(new_n17182_), .A2(\asqrt[58] ), .B1(new_n17180_), .B2(new_n17177_), .ZN(new_n17185_));
  OAI21_X1   g16993(.A1(new_n17185_), .A2(new_n376_), .B(new_n17029_), .ZN(new_n17186_));
  NAND2_X1   g16994(.A1(new_n17186_), .A2(new_n17184_), .ZN(new_n17187_));
  NAND2_X1   g16995(.A1(new_n17175_), .A2(\asqrt[56] ), .ZN(new_n17188_));
  AOI21_X1   g16996(.A1(new_n17188_), .A2(new_n17174_), .B(new_n587_), .ZN(new_n17189_));
  OAI21_X1   g16997(.A1(new_n17177_), .A2(new_n17189_), .B(\asqrt[58] ), .ZN(new_n17190_));
  AOI21_X1   g16998(.A1(new_n17181_), .A2(new_n17190_), .B(new_n376_), .ZN(new_n17191_));
  OAI21_X1   g16999(.A1(new_n17184_), .A2(new_n17191_), .B(\asqrt[60] ), .ZN(new_n17192_));
  NAND2_X1   g17000(.A1(new_n17187_), .A2(new_n17192_), .ZN(new_n17193_));
  AOI22_X1   g17001(.A1(new_n17193_), .A2(\asqrt[61] ), .B1(new_n17037_), .B2(new_n17030_), .ZN(new_n17194_));
  NOR2_X1    g17002(.A1(new_n17194_), .A2(new_n196_), .ZN(new_n17195_));
  NOR4_X1    g17003(.A1(new_n16619_), .A2(\asqrt[61] ), .A3(new_n16404_), .A4(new_n16409_), .ZN(new_n17196_));
  XOR2_X1    g17004(.A1(new_n17196_), .A2(new_n16626_), .Z(new_n17197_));
  INV_X1     g17005(.I(new_n17197_), .ZN(new_n17198_));
  NAND2_X1   g17006(.A1(new_n17037_), .A2(new_n17030_), .ZN(new_n17199_));
  AOI21_X1   g17007(.A1(new_n17019_), .A2(new_n17026_), .B(new_n275_), .ZN(new_n17200_));
  OAI21_X1   g17008(.A1(new_n17030_), .A2(new_n17200_), .B(\asqrt[61] ), .ZN(new_n17201_));
  NAND4_X1   g17009(.A1(new_n17199_), .A2(new_n17201_), .A3(new_n196_), .A4(new_n17198_), .ZN(new_n17202_));
  INV_X1     g17010(.I(new_n17202_), .ZN(new_n17203_));
  NOR2_X1    g17011(.A1(new_n16606_), .A2(new_n196_), .ZN(new_n17204_));
  NOR2_X1    g17012(.A1(new_n16591_), .A2(\asqrt[62] ), .ZN(new_n17205_));
  NAND3_X1   g17013(.A1(new_n17205_), .A2(new_n17204_), .A3(new_n16410_), .ZN(new_n17206_));
  NOR2_X1    g17014(.A1(new_n16619_), .A2(new_n17206_), .ZN(new_n17207_));
  OR3_X2     g17015(.A1(\asqrt[12] ), .A2(new_n16410_), .A3(new_n17205_), .Z(new_n17208_));
  AOI21_X1   g17016(.A1(new_n17208_), .A2(new_n17204_), .B(new_n17207_), .ZN(new_n17209_));
  NOR2_X1    g17017(.A1(new_n17197_), .A2(new_n196_), .ZN(new_n17210_));
  INV_X1     g17018(.I(new_n17210_), .ZN(new_n17211_));
  AOI21_X1   g17019(.A1(new_n17187_), .A2(new_n17192_), .B(new_n229_), .ZN(new_n17212_));
  NOR2_X1    g17020(.A1(new_n17198_), .A2(\asqrt[62] ), .ZN(new_n17213_));
  INV_X1     g17021(.I(new_n17213_), .ZN(new_n17214_));
  NAND2_X1   g17022(.A1(new_n17212_), .A2(new_n17214_), .ZN(new_n17215_));
  OAI21_X1   g17023(.A1(new_n17215_), .A2(new_n17199_), .B(new_n17211_), .ZN(new_n17216_));
  NOR3_X1    g17024(.A1(\asqrt[12] ), .A2(new_n16028_), .A3(new_n16592_), .ZN(new_n17217_));
  OAI21_X1   g17025(.A1(new_n17217_), .A2(new_n16604_), .B(new_n231_), .ZN(new_n17218_));
  OAI21_X1   g17026(.A1(new_n17216_), .A2(new_n17218_), .B(new_n17209_), .ZN(new_n17219_));
  OAI21_X1   g17027(.A1(new_n16028_), .A2(new_n16414_), .B(\asqrt[12] ), .ZN(new_n17220_));
  XOR2_X1    g17028(.A1(new_n16414_), .A2(\asqrt[63] ), .Z(new_n17221_));
  NAND2_X1   g17029(.A1(new_n17220_), .A2(new_n17221_), .ZN(new_n17222_));
  INV_X1     g17030(.I(new_n17222_), .ZN(new_n17223_));
  INV_X1     g17031(.I(new_n17209_), .ZN(new_n17224_));
  OAI22_X1   g17032(.A1(new_n17185_), .A2(new_n376_), .B1(new_n17183_), .B2(new_n17181_), .ZN(new_n17225_));
  AOI21_X1   g17033(.A1(new_n17225_), .A2(\asqrt[60] ), .B(new_n17035_), .ZN(new_n17226_));
  AOI22_X1   g17034(.A1(new_n17225_), .A2(\asqrt[60] ), .B1(new_n17186_), .B2(new_n17184_), .ZN(new_n17227_));
  OAI22_X1   g17035(.A1(new_n17227_), .A2(new_n229_), .B1(new_n17226_), .B2(new_n17187_), .ZN(new_n17228_));
  NOR4_X1    g17036(.A1(new_n17228_), .A2(\asqrt[62] ), .A3(new_n17224_), .A4(new_n17197_), .ZN(new_n17229_));
  NAND2_X1   g17037(.A1(new_n17229_), .A2(new_n17223_), .ZN(new_n17230_));
  NAND3_X1   g17038(.A1(new_n16613_), .A2(new_n16015_), .A3(new_n16028_), .ZN(new_n17231_));
  NOR3_X1    g17039(.A1(new_n17230_), .A2(new_n17219_), .A3(new_n17231_), .ZN(\asqrt[11] ));
  NAND3_X1   g17040(.A1(\asqrt[11] ), .A2(new_n17195_), .A3(new_n17203_), .ZN(new_n17233_));
  OAI21_X1   g17041(.A1(new_n17228_), .A2(\asqrt[62] ), .B(new_n17197_), .ZN(new_n17234_));
  OAI21_X1   g17042(.A1(\asqrt[11] ), .A2(new_n17234_), .B(new_n17195_), .ZN(new_n17235_));
  NAND2_X1   g17043(.A1(new_n17235_), .A2(new_n17233_), .ZN(new_n17236_));
  INV_X1     g17044(.I(new_n17236_), .ZN(new_n17237_));
  NOR3_X1    g17045(.A1(new_n17193_), .A2(\asqrt[61] ), .A3(new_n17034_), .ZN(new_n17238_));
  NAND2_X1   g17046(.A1(\asqrt[11] ), .A2(new_n17238_), .ZN(new_n17239_));
  XOR2_X1    g17047(.A1(new_n17239_), .A2(new_n17212_), .Z(new_n17240_));
  NOR2_X1    g17048(.A1(new_n17240_), .A2(new_n196_), .ZN(new_n17241_));
  INV_X1     g17049(.I(new_n17241_), .ZN(new_n17242_));
  INV_X1     g17050(.I(\a[22] ), .ZN(new_n17243_));
  NOR2_X1    g17051(.A1(\a[20] ), .A2(\a[21] ), .ZN(new_n17244_));
  INV_X1     g17052(.I(new_n17244_), .ZN(new_n17245_));
  NOR3_X1    g17053(.A1(new_n16630_), .A2(new_n17243_), .A3(new_n17245_), .ZN(new_n17246_));
  NAND2_X1   g17054(.A1(new_n16645_), .A2(new_n17246_), .ZN(new_n17247_));
  XOR2_X1    g17055(.A1(new_n17247_), .A2(\a[23] ), .Z(new_n17248_));
  INV_X1     g17056(.I(\a[23] ), .ZN(new_n17249_));
  NOR4_X1    g17057(.A1(new_n17230_), .A2(new_n17219_), .A3(new_n17249_), .A4(new_n17231_), .ZN(new_n17250_));
  NOR2_X1    g17058(.A1(new_n17249_), .A2(\a[22] ), .ZN(new_n17251_));
  OAI21_X1   g17059(.A1(new_n17250_), .A2(new_n17251_), .B(new_n17248_), .ZN(new_n17252_));
  INV_X1     g17060(.I(new_n17248_), .ZN(new_n17253_));
  NOR2_X1    g17061(.A1(new_n17226_), .A2(new_n17187_), .ZN(new_n17254_));
  NOR3_X1    g17062(.A1(new_n17227_), .A2(new_n229_), .A3(new_n17213_), .ZN(new_n17255_));
  AOI21_X1   g17063(.A1(new_n17255_), .A2(new_n17254_), .B(new_n17210_), .ZN(new_n17256_));
  INV_X1     g17064(.I(new_n17218_), .ZN(new_n17257_));
  AOI21_X1   g17065(.A1(new_n17256_), .A2(new_n17257_), .B(new_n17224_), .ZN(new_n17258_));
  AOI21_X1   g17066(.A1(new_n17228_), .A2(\asqrt[62] ), .B(new_n17209_), .ZN(new_n17259_));
  NOR3_X1    g17067(.A1(new_n17259_), .A2(new_n17222_), .A3(new_n17202_), .ZN(new_n17260_));
  INV_X1     g17068(.I(new_n17231_), .ZN(new_n17261_));
  NAND4_X1   g17069(.A1(new_n17260_), .A2(\a[23] ), .A3(new_n17258_), .A4(new_n17261_), .ZN(new_n17262_));
  NAND3_X1   g17070(.A1(new_n17262_), .A2(\a[22] ), .A3(new_n17253_), .ZN(new_n17263_));
  NAND2_X1   g17071(.A1(new_n17252_), .A2(new_n17263_), .ZN(new_n17264_));
  NOR2_X1    g17072(.A1(new_n17230_), .A2(new_n17219_), .ZN(new_n17265_));
  NAND4_X1   g17073(.A1(new_n16609_), .A2(new_n16601_), .A3(new_n16028_), .A4(new_n16644_), .ZN(new_n17266_));
  NOR2_X1    g17074(.A1(new_n16619_), .A2(new_n17243_), .ZN(new_n17267_));
  XOR2_X1    g17075(.A1(new_n17267_), .A2(new_n17266_), .Z(new_n17268_));
  NOR2_X1    g17076(.A1(new_n17268_), .A2(new_n17245_), .ZN(new_n17269_));
  INV_X1     g17077(.I(new_n17269_), .ZN(new_n17270_));
  NAND3_X1   g17078(.A1(new_n17260_), .A2(new_n17258_), .A3(new_n17261_), .ZN(new_n17271_));
  NOR4_X1    g17079(.A1(new_n17201_), .A2(new_n17187_), .A3(new_n17226_), .A4(new_n17213_), .ZN(new_n17272_));
  NOR3_X1    g17080(.A1(new_n17272_), .A2(new_n17210_), .A3(new_n17218_), .ZN(new_n17273_));
  NAND4_X1   g17081(.A1(new_n17194_), .A2(new_n196_), .A3(new_n17209_), .A4(new_n17198_), .ZN(new_n17274_));
  OAI21_X1   g17082(.A1(new_n17273_), .A2(new_n17224_), .B(new_n17274_), .ZN(new_n17275_));
  NOR2_X1    g17083(.A1(new_n17223_), .A2(new_n17261_), .ZN(new_n17276_));
  NAND2_X1   g17084(.A1(new_n17276_), .A2(\asqrt[12] ), .ZN(new_n17277_));
  OAI21_X1   g17085(.A1(new_n17275_), .A2(new_n17277_), .B(new_n15995_), .ZN(new_n17278_));
  NAND3_X1   g17086(.A1(new_n17278_), .A2(new_n16003_), .A3(new_n17271_), .ZN(new_n17279_));
  NAND4_X1   g17087(.A1(new_n17212_), .A2(new_n17030_), .A3(new_n17037_), .A4(new_n17214_), .ZN(new_n17280_));
  NAND3_X1   g17088(.A1(new_n17280_), .A2(new_n17211_), .A3(new_n17257_), .ZN(new_n17281_));
  AOI21_X1   g17089(.A1(new_n17209_), .A2(new_n17281_), .B(new_n17229_), .ZN(new_n17282_));
  INV_X1     g17090(.I(new_n17277_), .ZN(new_n17283_));
  AOI21_X1   g17091(.A1(new_n17282_), .A2(new_n17283_), .B(\a[24] ), .ZN(new_n17284_));
  OAI21_X1   g17092(.A1(new_n17284_), .A2(new_n16004_), .B(\asqrt[11] ), .ZN(new_n17285_));
  NAND4_X1   g17093(.A1(new_n17279_), .A2(new_n17285_), .A3(new_n16060_), .A4(new_n17270_), .ZN(new_n17286_));
  NAND2_X1   g17094(.A1(new_n17286_), .A2(new_n17264_), .ZN(new_n17287_));
  NAND3_X1   g17095(.A1(new_n17252_), .A2(new_n17263_), .A3(new_n17270_), .ZN(new_n17288_));
  INV_X1     g17096(.I(new_n16006_), .ZN(new_n17289_));
  NOR2_X1    g17097(.A1(new_n16619_), .A2(\a[24] ), .ZN(new_n17290_));
  OAI22_X1   g17098(.A1(new_n17290_), .A2(\a[25] ), .B1(\a[24] ), .B2(new_n16610_), .ZN(new_n17291_));
  NAND2_X1   g17099(.A1(\asqrt[12] ), .A2(\a[24] ), .ZN(new_n17292_));
  AND3_X2    g17100(.A1(new_n17291_), .A2(new_n17289_), .A3(new_n17292_), .Z(new_n17293_));
  NAND3_X1   g17101(.A1(\asqrt[11] ), .A2(new_n16618_), .A3(new_n17293_), .ZN(new_n17294_));
  INV_X1     g17102(.I(new_n17293_), .ZN(new_n17295_));
  OAI21_X1   g17103(.A1(new_n17271_), .A2(new_n17295_), .B(new_n16617_), .ZN(new_n17296_));
  NAND3_X1   g17104(.A1(new_n17294_), .A2(new_n17296_), .A3(new_n15447_), .ZN(new_n17297_));
  AOI21_X1   g17105(.A1(new_n17288_), .A2(\asqrt[13] ), .B(new_n17297_), .ZN(new_n17298_));
  NOR2_X1    g17106(.A1(new_n17287_), .A2(new_n17298_), .ZN(new_n17299_));
  AOI22_X1   g17107(.A1(new_n17286_), .A2(new_n17264_), .B1(\asqrt[13] ), .B2(new_n17288_), .ZN(new_n17300_));
  AOI21_X1   g17108(.A1(new_n16648_), .A2(new_n16633_), .B(\asqrt[14] ), .ZN(new_n17301_));
  AND4_X2    g17109(.A1(new_n16691_), .A2(\asqrt[11] ), .A3(new_n16672_), .A4(new_n17301_), .Z(new_n17302_));
  NOR2_X1    g17110(.A1(new_n16691_), .A2(new_n15447_), .ZN(new_n17303_));
  NOR3_X1    g17111(.A1(new_n17302_), .A2(\asqrt[15] ), .A3(new_n17303_), .ZN(new_n17304_));
  OAI21_X1   g17112(.A1(new_n17300_), .A2(new_n15447_), .B(new_n17304_), .ZN(new_n17305_));
  NAND2_X1   g17113(.A1(new_n17305_), .A2(new_n17299_), .ZN(new_n17306_));
  OAI22_X1   g17114(.A1(new_n17300_), .A2(new_n15447_), .B1(new_n17287_), .B2(new_n17298_), .ZN(new_n17307_));
  NAND2_X1   g17115(.A1(new_n16657_), .A2(new_n16658_), .ZN(new_n17308_));
  NAND4_X1   g17116(.A1(\asqrt[11] ), .A2(new_n14871_), .A3(new_n17308_), .A4(new_n16662_), .ZN(new_n17309_));
  XOR2_X1    g17117(.A1(new_n17309_), .A2(new_n16673_), .Z(new_n17310_));
  NAND2_X1   g17118(.A1(new_n17310_), .A2(new_n14273_), .ZN(new_n17311_));
  AOI21_X1   g17119(.A1(new_n17307_), .A2(\asqrt[15] ), .B(new_n17311_), .ZN(new_n17312_));
  NOR2_X1    g17120(.A1(new_n17312_), .A2(new_n17306_), .ZN(new_n17313_));
  AOI22_X1   g17121(.A1(new_n17307_), .A2(\asqrt[15] ), .B1(new_n17305_), .B2(new_n17299_), .ZN(new_n17314_));
  NOR2_X1    g17122(.A1(new_n16669_), .A2(new_n16667_), .ZN(new_n17315_));
  NOR4_X1    g17123(.A1(new_n17271_), .A2(\asqrt[16] ), .A3(new_n17315_), .A4(new_n17038_), .ZN(new_n17316_));
  XOR2_X1    g17124(.A1(new_n17316_), .A2(new_n16674_), .Z(new_n17317_));
  NAND2_X1   g17125(.A1(new_n17317_), .A2(new_n13760_), .ZN(new_n17318_));
  INV_X1     g17126(.I(new_n17318_), .ZN(new_n17319_));
  OAI21_X1   g17127(.A1(new_n17314_), .A2(new_n14273_), .B(new_n17319_), .ZN(new_n17320_));
  NAND2_X1   g17128(.A1(new_n17320_), .A2(new_n17313_), .ZN(new_n17321_));
  OAI22_X1   g17129(.A1(new_n17314_), .A2(new_n14273_), .B1(new_n17312_), .B2(new_n17306_), .ZN(new_n17322_));
  NOR4_X1    g17130(.A1(new_n17271_), .A2(\asqrt[17] ), .A3(new_n16678_), .A4(new_n16701_), .ZN(new_n17323_));
  XNOR2_X1   g17131(.A1(new_n17323_), .A2(new_n16711_), .ZN(new_n17324_));
  NAND2_X1   g17132(.A1(new_n17324_), .A2(new_n13192_), .ZN(new_n17325_));
  AOI21_X1   g17133(.A1(new_n17322_), .A2(\asqrt[17] ), .B(new_n17325_), .ZN(new_n17326_));
  NOR2_X1    g17134(.A1(new_n17326_), .A2(new_n17321_), .ZN(new_n17327_));
  AOI22_X1   g17135(.A1(new_n17322_), .A2(\asqrt[17] ), .B1(new_n17320_), .B2(new_n17313_), .ZN(new_n17328_));
  NOR4_X1    g17136(.A1(new_n17271_), .A2(\asqrt[18] ), .A3(new_n16705_), .A4(new_n17043_), .ZN(new_n17329_));
  XOR2_X1    g17137(.A1(new_n17329_), .A2(new_n16712_), .Z(new_n17330_));
  NAND2_X1   g17138(.A1(new_n17330_), .A2(new_n12657_), .ZN(new_n17331_));
  INV_X1     g17139(.I(new_n17331_), .ZN(new_n17332_));
  OAI21_X1   g17140(.A1(new_n17328_), .A2(new_n13192_), .B(new_n17332_), .ZN(new_n17333_));
  NAND2_X1   g17141(.A1(new_n17333_), .A2(new_n17327_), .ZN(new_n17334_));
  OAI22_X1   g17142(.A1(new_n17328_), .A2(new_n13192_), .B1(new_n17326_), .B2(new_n17321_), .ZN(new_n17335_));
  NOR4_X1    g17143(.A1(new_n17271_), .A2(\asqrt[19] ), .A3(new_n16715_), .A4(new_n16721_), .ZN(new_n17336_));
  XNOR2_X1   g17144(.A1(new_n17336_), .A2(new_n16730_), .ZN(new_n17337_));
  NAND2_X1   g17145(.A1(new_n17337_), .A2(new_n12101_), .ZN(new_n17338_));
  AOI21_X1   g17146(.A1(new_n17335_), .A2(\asqrt[19] ), .B(new_n17338_), .ZN(new_n17339_));
  NOR2_X1    g17147(.A1(new_n17339_), .A2(new_n17334_), .ZN(new_n17340_));
  AOI22_X1   g17148(.A1(new_n17335_), .A2(\asqrt[19] ), .B1(new_n17333_), .B2(new_n17327_), .ZN(new_n17341_));
  NOR4_X1    g17149(.A1(new_n17271_), .A2(\asqrt[20] ), .A3(new_n16724_), .A4(new_n17049_), .ZN(new_n17342_));
  XOR2_X1    g17150(.A1(new_n17342_), .A2(new_n16731_), .Z(new_n17343_));
  NAND2_X1   g17151(.A1(new_n17343_), .A2(new_n11631_), .ZN(new_n17344_));
  INV_X1     g17152(.I(new_n17344_), .ZN(new_n17345_));
  OAI21_X1   g17153(.A1(new_n17341_), .A2(new_n12101_), .B(new_n17345_), .ZN(new_n17346_));
  NAND2_X1   g17154(.A1(new_n17346_), .A2(new_n17340_), .ZN(new_n17347_));
  OAI22_X1   g17155(.A1(new_n17341_), .A2(new_n12101_), .B1(new_n17339_), .B2(new_n17334_), .ZN(new_n17348_));
  NAND2_X1   g17156(.A1(new_n16740_), .A2(\asqrt[21] ), .ZN(new_n17349_));
  NOR4_X1    g17157(.A1(new_n17271_), .A2(\asqrt[21] ), .A3(new_n16734_), .A4(new_n16740_), .ZN(new_n17350_));
  XOR2_X1    g17158(.A1(new_n17350_), .A2(new_n17349_), .Z(new_n17351_));
  NAND2_X1   g17159(.A1(new_n17351_), .A2(new_n11105_), .ZN(new_n17352_));
  AOI21_X1   g17160(.A1(new_n17348_), .A2(\asqrt[21] ), .B(new_n17352_), .ZN(new_n17353_));
  NOR2_X1    g17161(.A1(new_n17353_), .A2(new_n17347_), .ZN(new_n17354_));
  AOI22_X1   g17162(.A1(new_n17348_), .A2(\asqrt[21] ), .B1(new_n17346_), .B2(new_n17340_), .ZN(new_n17355_));
  NOR4_X1    g17163(.A1(new_n17271_), .A2(\asqrt[22] ), .A3(new_n16743_), .A4(new_n17056_), .ZN(new_n17356_));
  AOI21_X1   g17164(.A1(new_n17349_), .A2(new_n16738_), .B(new_n11105_), .ZN(new_n17357_));
  NOR2_X1    g17165(.A1(new_n17356_), .A2(new_n17357_), .ZN(new_n17358_));
  NAND2_X1   g17166(.A1(new_n17358_), .A2(new_n10614_), .ZN(new_n17359_));
  INV_X1     g17167(.I(new_n17359_), .ZN(new_n17360_));
  OAI21_X1   g17168(.A1(new_n17355_), .A2(new_n11105_), .B(new_n17360_), .ZN(new_n17361_));
  NAND2_X1   g17169(.A1(new_n17361_), .A2(new_n17354_), .ZN(new_n17362_));
  OAI22_X1   g17170(.A1(new_n17355_), .A2(new_n11105_), .B1(new_n17353_), .B2(new_n17347_), .ZN(new_n17363_));
  NAND2_X1   g17171(.A1(new_n16755_), .A2(\asqrt[23] ), .ZN(new_n17364_));
  NOR4_X1    g17172(.A1(new_n17271_), .A2(\asqrt[23] ), .A3(new_n16750_), .A4(new_n16755_), .ZN(new_n17365_));
  XOR2_X1    g17173(.A1(new_n17365_), .A2(new_n17364_), .Z(new_n17366_));
  NAND2_X1   g17174(.A1(new_n17366_), .A2(new_n10104_), .ZN(new_n17367_));
  AOI21_X1   g17175(.A1(new_n17363_), .A2(\asqrt[23] ), .B(new_n17367_), .ZN(new_n17368_));
  NOR2_X1    g17176(.A1(new_n17368_), .A2(new_n17362_), .ZN(new_n17369_));
  AOI22_X1   g17177(.A1(new_n17363_), .A2(\asqrt[23] ), .B1(new_n17361_), .B2(new_n17354_), .ZN(new_n17370_));
  NOR4_X1    g17178(.A1(new_n17271_), .A2(\asqrt[24] ), .A3(new_n16758_), .A4(new_n17063_), .ZN(new_n17371_));
  AOI21_X1   g17179(.A1(new_n17364_), .A2(new_n16754_), .B(new_n10104_), .ZN(new_n17372_));
  NOR2_X1    g17180(.A1(new_n17371_), .A2(new_n17372_), .ZN(new_n17373_));
  NAND2_X1   g17181(.A1(new_n17373_), .A2(new_n9672_), .ZN(new_n17374_));
  INV_X1     g17182(.I(new_n17374_), .ZN(new_n17375_));
  OAI21_X1   g17183(.A1(new_n17370_), .A2(new_n10104_), .B(new_n17375_), .ZN(new_n17376_));
  NAND2_X1   g17184(.A1(new_n17376_), .A2(new_n17369_), .ZN(new_n17377_));
  OAI22_X1   g17185(.A1(new_n17370_), .A2(new_n10104_), .B1(new_n17368_), .B2(new_n17362_), .ZN(new_n17378_));
  NAND2_X1   g17186(.A1(new_n16770_), .A2(\asqrt[25] ), .ZN(new_n17379_));
  NOR4_X1    g17187(.A1(new_n17271_), .A2(\asqrt[25] ), .A3(new_n16765_), .A4(new_n16770_), .ZN(new_n17380_));
  XOR2_X1    g17188(.A1(new_n17380_), .A2(new_n17379_), .Z(new_n17381_));
  NAND2_X1   g17189(.A1(new_n17381_), .A2(new_n9212_), .ZN(new_n17382_));
  AOI21_X1   g17190(.A1(new_n17378_), .A2(\asqrt[25] ), .B(new_n17382_), .ZN(new_n17383_));
  NOR2_X1    g17191(.A1(new_n17383_), .A2(new_n17377_), .ZN(new_n17384_));
  AOI22_X1   g17192(.A1(new_n17378_), .A2(\asqrt[25] ), .B1(new_n17376_), .B2(new_n17369_), .ZN(new_n17385_));
  NOR4_X1    g17193(.A1(new_n17271_), .A2(\asqrt[26] ), .A3(new_n16773_), .A4(new_n17070_), .ZN(new_n17386_));
  AOI21_X1   g17194(.A1(new_n17379_), .A2(new_n16769_), .B(new_n9212_), .ZN(new_n17387_));
  NOR2_X1    g17195(.A1(new_n17386_), .A2(new_n17387_), .ZN(new_n17388_));
  NAND2_X1   g17196(.A1(new_n17388_), .A2(new_n8763_), .ZN(new_n17389_));
  INV_X1     g17197(.I(new_n17389_), .ZN(new_n17390_));
  OAI21_X1   g17198(.A1(new_n17385_), .A2(new_n9212_), .B(new_n17390_), .ZN(new_n17391_));
  NAND2_X1   g17199(.A1(new_n17391_), .A2(new_n17384_), .ZN(new_n17392_));
  OAI22_X1   g17200(.A1(new_n17385_), .A2(new_n9212_), .B1(new_n17383_), .B2(new_n17377_), .ZN(new_n17393_));
  NAND2_X1   g17201(.A1(new_n16785_), .A2(\asqrt[27] ), .ZN(new_n17394_));
  NOR4_X1    g17202(.A1(new_n17271_), .A2(\asqrt[27] ), .A3(new_n16780_), .A4(new_n16785_), .ZN(new_n17395_));
  XOR2_X1    g17203(.A1(new_n17395_), .A2(new_n17394_), .Z(new_n17396_));
  NAND2_X1   g17204(.A1(new_n17396_), .A2(new_n8319_), .ZN(new_n17397_));
  AOI21_X1   g17205(.A1(new_n17393_), .A2(\asqrt[27] ), .B(new_n17397_), .ZN(new_n17398_));
  NOR2_X1    g17206(.A1(new_n17398_), .A2(new_n17392_), .ZN(new_n17399_));
  AOI22_X1   g17207(.A1(new_n17393_), .A2(\asqrt[27] ), .B1(new_n17391_), .B2(new_n17384_), .ZN(new_n17400_));
  NOR4_X1    g17208(.A1(new_n17271_), .A2(\asqrt[28] ), .A3(new_n16788_), .A4(new_n17077_), .ZN(new_n17401_));
  AOI21_X1   g17209(.A1(new_n17394_), .A2(new_n16784_), .B(new_n8319_), .ZN(new_n17402_));
  NOR2_X1    g17210(.A1(new_n17401_), .A2(new_n17402_), .ZN(new_n17403_));
  NAND2_X1   g17211(.A1(new_n17403_), .A2(new_n7931_), .ZN(new_n17404_));
  INV_X1     g17212(.I(new_n17404_), .ZN(new_n17405_));
  OAI21_X1   g17213(.A1(new_n17400_), .A2(new_n8319_), .B(new_n17405_), .ZN(new_n17406_));
  NAND2_X1   g17214(.A1(new_n17406_), .A2(new_n17399_), .ZN(new_n17407_));
  OAI22_X1   g17215(.A1(new_n17400_), .A2(new_n8319_), .B1(new_n17398_), .B2(new_n17392_), .ZN(new_n17408_));
  NAND2_X1   g17216(.A1(new_n16800_), .A2(\asqrt[29] ), .ZN(new_n17409_));
  NOR4_X1    g17217(.A1(new_n17271_), .A2(\asqrt[29] ), .A3(new_n16795_), .A4(new_n16800_), .ZN(new_n17410_));
  XOR2_X1    g17218(.A1(new_n17410_), .A2(new_n17409_), .Z(new_n17411_));
  NAND2_X1   g17219(.A1(new_n17411_), .A2(new_n7517_), .ZN(new_n17412_));
  AOI21_X1   g17220(.A1(new_n17408_), .A2(\asqrt[29] ), .B(new_n17412_), .ZN(new_n17413_));
  NOR2_X1    g17221(.A1(new_n17413_), .A2(new_n17407_), .ZN(new_n17414_));
  AOI22_X1   g17222(.A1(new_n17408_), .A2(\asqrt[29] ), .B1(new_n17406_), .B2(new_n17399_), .ZN(new_n17415_));
  NOR4_X1    g17223(.A1(new_n17271_), .A2(\asqrt[30] ), .A3(new_n16803_), .A4(new_n17084_), .ZN(new_n17416_));
  AOI21_X1   g17224(.A1(new_n17409_), .A2(new_n16799_), .B(new_n7517_), .ZN(new_n17417_));
  NOR2_X1    g17225(.A1(new_n17416_), .A2(new_n17417_), .ZN(new_n17418_));
  NAND2_X1   g17226(.A1(new_n17418_), .A2(new_n7110_), .ZN(new_n17419_));
  INV_X1     g17227(.I(new_n17419_), .ZN(new_n17420_));
  OAI21_X1   g17228(.A1(new_n17415_), .A2(new_n7517_), .B(new_n17420_), .ZN(new_n17421_));
  NAND2_X1   g17229(.A1(new_n17421_), .A2(new_n17414_), .ZN(new_n17422_));
  OAI22_X1   g17230(.A1(new_n17415_), .A2(new_n7517_), .B1(new_n17413_), .B2(new_n17407_), .ZN(new_n17423_));
  NAND2_X1   g17231(.A1(new_n16815_), .A2(\asqrt[31] ), .ZN(new_n17424_));
  NOR4_X1    g17232(.A1(new_n17271_), .A2(\asqrt[31] ), .A3(new_n16810_), .A4(new_n16815_), .ZN(new_n17425_));
  XOR2_X1    g17233(.A1(new_n17425_), .A2(new_n17424_), .Z(new_n17426_));
  NAND2_X1   g17234(.A1(new_n17426_), .A2(new_n6708_), .ZN(new_n17427_));
  AOI21_X1   g17235(.A1(new_n17423_), .A2(\asqrt[31] ), .B(new_n17427_), .ZN(new_n17428_));
  NOR2_X1    g17236(.A1(new_n17428_), .A2(new_n17422_), .ZN(new_n17429_));
  AOI22_X1   g17237(.A1(new_n17423_), .A2(\asqrt[31] ), .B1(new_n17421_), .B2(new_n17414_), .ZN(new_n17430_));
  NAND2_X1   g17238(.A1(new_n17091_), .A2(\asqrt[32] ), .ZN(new_n17431_));
  NOR4_X1    g17239(.A1(new_n17271_), .A2(\asqrt[32] ), .A3(new_n16818_), .A4(new_n17091_), .ZN(new_n17432_));
  XOR2_X1    g17240(.A1(new_n17432_), .A2(new_n17431_), .Z(new_n17433_));
  NAND2_X1   g17241(.A1(new_n17433_), .A2(new_n6365_), .ZN(new_n17434_));
  INV_X1     g17242(.I(new_n17434_), .ZN(new_n17435_));
  OAI21_X1   g17243(.A1(new_n17430_), .A2(new_n6708_), .B(new_n17435_), .ZN(new_n17436_));
  NAND2_X1   g17244(.A1(new_n17436_), .A2(new_n17429_), .ZN(new_n17437_));
  OAI22_X1   g17245(.A1(new_n17430_), .A2(new_n6708_), .B1(new_n17428_), .B2(new_n17422_), .ZN(new_n17438_));
  NOR4_X1    g17246(.A1(new_n17271_), .A2(\asqrt[33] ), .A3(new_n16825_), .A4(new_n16830_), .ZN(new_n17439_));
  AOI21_X1   g17247(.A1(new_n17431_), .A2(new_n17090_), .B(new_n6365_), .ZN(new_n17440_));
  NOR2_X1    g17248(.A1(new_n17439_), .A2(new_n17440_), .ZN(new_n17441_));
  NAND2_X1   g17249(.A1(new_n17441_), .A2(new_n5991_), .ZN(new_n17442_));
  AOI21_X1   g17250(.A1(new_n17438_), .A2(\asqrt[33] ), .B(new_n17442_), .ZN(new_n17443_));
  NOR2_X1    g17251(.A1(new_n17443_), .A2(new_n17437_), .ZN(new_n17444_));
  AOI22_X1   g17252(.A1(new_n17438_), .A2(\asqrt[33] ), .B1(new_n17436_), .B2(new_n17429_), .ZN(new_n17445_));
  NAND2_X1   g17253(.A1(new_n17098_), .A2(\asqrt[34] ), .ZN(new_n17446_));
  NOR4_X1    g17254(.A1(new_n17271_), .A2(\asqrt[34] ), .A3(new_n16833_), .A4(new_n17098_), .ZN(new_n17447_));
  XOR2_X1    g17255(.A1(new_n17447_), .A2(new_n17446_), .Z(new_n17448_));
  NAND2_X1   g17256(.A1(new_n17448_), .A2(new_n5626_), .ZN(new_n17449_));
  INV_X1     g17257(.I(new_n17449_), .ZN(new_n17450_));
  OAI21_X1   g17258(.A1(new_n17445_), .A2(new_n5991_), .B(new_n17450_), .ZN(new_n17451_));
  NAND2_X1   g17259(.A1(new_n17451_), .A2(new_n17444_), .ZN(new_n17452_));
  OAI22_X1   g17260(.A1(new_n17445_), .A2(new_n5991_), .B1(new_n17443_), .B2(new_n17437_), .ZN(new_n17453_));
  NOR4_X1    g17261(.A1(new_n17271_), .A2(\asqrt[35] ), .A3(new_n16840_), .A4(new_n16845_), .ZN(new_n17454_));
  AOI21_X1   g17262(.A1(new_n17446_), .A2(new_n17097_), .B(new_n5626_), .ZN(new_n17455_));
  NOR2_X1    g17263(.A1(new_n17454_), .A2(new_n17455_), .ZN(new_n17456_));
  NAND2_X1   g17264(.A1(new_n17456_), .A2(new_n5273_), .ZN(new_n17457_));
  AOI21_X1   g17265(.A1(new_n17453_), .A2(\asqrt[35] ), .B(new_n17457_), .ZN(new_n17458_));
  NOR2_X1    g17266(.A1(new_n17458_), .A2(new_n17452_), .ZN(new_n17459_));
  AOI22_X1   g17267(.A1(new_n17453_), .A2(\asqrt[35] ), .B1(new_n17451_), .B2(new_n17444_), .ZN(new_n17460_));
  NAND2_X1   g17268(.A1(new_n17105_), .A2(\asqrt[36] ), .ZN(new_n17461_));
  NOR4_X1    g17269(.A1(new_n17271_), .A2(\asqrt[36] ), .A3(new_n16848_), .A4(new_n17105_), .ZN(new_n17462_));
  XOR2_X1    g17270(.A1(new_n17462_), .A2(new_n17461_), .Z(new_n17463_));
  NAND2_X1   g17271(.A1(new_n17463_), .A2(new_n4973_), .ZN(new_n17464_));
  INV_X1     g17272(.I(new_n17464_), .ZN(new_n17465_));
  OAI21_X1   g17273(.A1(new_n17460_), .A2(new_n5273_), .B(new_n17465_), .ZN(new_n17466_));
  NAND2_X1   g17274(.A1(new_n17466_), .A2(new_n17459_), .ZN(new_n17467_));
  OAI22_X1   g17275(.A1(new_n17460_), .A2(new_n5273_), .B1(new_n17458_), .B2(new_n17452_), .ZN(new_n17468_));
  NAND2_X1   g17276(.A1(new_n16860_), .A2(\asqrt[37] ), .ZN(new_n17469_));
  NOR4_X1    g17277(.A1(new_n17271_), .A2(\asqrt[37] ), .A3(new_n16855_), .A4(new_n16860_), .ZN(new_n17470_));
  XOR2_X1    g17278(.A1(new_n17470_), .A2(new_n17469_), .Z(new_n17471_));
  NAND2_X1   g17279(.A1(new_n17471_), .A2(new_n4645_), .ZN(new_n17472_));
  AOI21_X1   g17280(.A1(new_n17468_), .A2(\asqrt[37] ), .B(new_n17472_), .ZN(new_n17473_));
  NOR2_X1    g17281(.A1(new_n17473_), .A2(new_n17467_), .ZN(new_n17474_));
  AOI22_X1   g17282(.A1(new_n17468_), .A2(\asqrt[37] ), .B1(new_n17466_), .B2(new_n17459_), .ZN(new_n17475_));
  NOR4_X1    g17283(.A1(new_n17271_), .A2(\asqrt[38] ), .A3(new_n16863_), .A4(new_n17112_), .ZN(new_n17476_));
  AOI21_X1   g17284(.A1(new_n17469_), .A2(new_n16859_), .B(new_n4645_), .ZN(new_n17477_));
  NOR2_X1    g17285(.A1(new_n17476_), .A2(new_n17477_), .ZN(new_n17478_));
  NAND2_X1   g17286(.A1(new_n17478_), .A2(new_n4330_), .ZN(new_n17479_));
  INV_X1     g17287(.I(new_n17479_), .ZN(new_n17480_));
  OAI21_X1   g17288(.A1(new_n17475_), .A2(new_n4645_), .B(new_n17480_), .ZN(new_n17481_));
  NAND2_X1   g17289(.A1(new_n17481_), .A2(new_n17474_), .ZN(new_n17482_));
  OAI22_X1   g17290(.A1(new_n17475_), .A2(new_n4645_), .B1(new_n17473_), .B2(new_n17467_), .ZN(new_n17483_));
  NAND2_X1   g17291(.A1(new_n16875_), .A2(\asqrt[39] ), .ZN(new_n17484_));
  NOR4_X1    g17292(.A1(new_n17271_), .A2(\asqrt[39] ), .A3(new_n16870_), .A4(new_n16875_), .ZN(new_n17485_));
  XOR2_X1    g17293(.A1(new_n17485_), .A2(new_n17484_), .Z(new_n17486_));
  NAND2_X1   g17294(.A1(new_n17486_), .A2(new_n4018_), .ZN(new_n17487_));
  AOI21_X1   g17295(.A1(new_n17483_), .A2(\asqrt[39] ), .B(new_n17487_), .ZN(new_n17488_));
  NOR2_X1    g17296(.A1(new_n17488_), .A2(new_n17482_), .ZN(new_n17489_));
  AOI22_X1   g17297(.A1(new_n17483_), .A2(\asqrt[39] ), .B1(new_n17481_), .B2(new_n17474_), .ZN(new_n17490_));
  NOR4_X1    g17298(.A1(new_n17271_), .A2(\asqrt[40] ), .A3(new_n16878_), .A4(new_n17119_), .ZN(new_n17491_));
  AOI21_X1   g17299(.A1(new_n17484_), .A2(new_n16874_), .B(new_n4018_), .ZN(new_n17492_));
  NOR2_X1    g17300(.A1(new_n17491_), .A2(new_n17492_), .ZN(new_n17493_));
  NAND2_X1   g17301(.A1(new_n17493_), .A2(new_n3760_), .ZN(new_n17494_));
  INV_X1     g17302(.I(new_n17494_), .ZN(new_n17495_));
  OAI21_X1   g17303(.A1(new_n17490_), .A2(new_n4018_), .B(new_n17495_), .ZN(new_n17496_));
  NAND2_X1   g17304(.A1(new_n17496_), .A2(new_n17489_), .ZN(new_n17497_));
  OAI22_X1   g17305(.A1(new_n17490_), .A2(new_n4018_), .B1(new_n17488_), .B2(new_n17482_), .ZN(new_n17498_));
  NAND2_X1   g17306(.A1(new_n16890_), .A2(\asqrt[41] ), .ZN(new_n17499_));
  NOR4_X1    g17307(.A1(new_n17271_), .A2(\asqrt[41] ), .A3(new_n16885_), .A4(new_n16890_), .ZN(new_n17500_));
  XOR2_X1    g17308(.A1(new_n17500_), .A2(new_n17499_), .Z(new_n17501_));
  NAND2_X1   g17309(.A1(new_n17501_), .A2(new_n3481_), .ZN(new_n17502_));
  AOI21_X1   g17310(.A1(new_n17498_), .A2(\asqrt[41] ), .B(new_n17502_), .ZN(new_n17503_));
  NOR2_X1    g17311(.A1(new_n17503_), .A2(new_n17497_), .ZN(new_n17504_));
  AOI22_X1   g17312(.A1(new_n17498_), .A2(\asqrt[41] ), .B1(new_n17496_), .B2(new_n17489_), .ZN(new_n17505_));
  NOR4_X1    g17313(.A1(new_n17271_), .A2(\asqrt[42] ), .A3(new_n16893_), .A4(new_n17126_), .ZN(new_n17506_));
  AOI21_X1   g17314(.A1(new_n17499_), .A2(new_n16889_), .B(new_n3481_), .ZN(new_n17507_));
  NOR2_X1    g17315(.A1(new_n17506_), .A2(new_n17507_), .ZN(new_n17508_));
  NAND2_X1   g17316(.A1(new_n17508_), .A2(new_n3208_), .ZN(new_n17509_));
  INV_X1     g17317(.I(new_n17509_), .ZN(new_n17510_));
  OAI21_X1   g17318(.A1(new_n17505_), .A2(new_n3481_), .B(new_n17510_), .ZN(new_n17511_));
  NAND2_X1   g17319(.A1(new_n17511_), .A2(new_n17504_), .ZN(new_n17512_));
  OAI22_X1   g17320(.A1(new_n17505_), .A2(new_n3481_), .B1(new_n17503_), .B2(new_n17497_), .ZN(new_n17513_));
  NAND2_X1   g17321(.A1(new_n16905_), .A2(\asqrt[43] ), .ZN(new_n17514_));
  NOR4_X1    g17322(.A1(new_n17271_), .A2(\asqrt[43] ), .A3(new_n16900_), .A4(new_n16905_), .ZN(new_n17515_));
  XOR2_X1    g17323(.A1(new_n17515_), .A2(new_n17514_), .Z(new_n17516_));
  NAND2_X1   g17324(.A1(new_n17516_), .A2(new_n2941_), .ZN(new_n17517_));
  AOI21_X1   g17325(.A1(new_n17513_), .A2(\asqrt[43] ), .B(new_n17517_), .ZN(new_n17518_));
  NOR2_X1    g17326(.A1(new_n17518_), .A2(new_n17512_), .ZN(new_n17519_));
  AOI22_X1   g17327(.A1(new_n17513_), .A2(\asqrt[43] ), .B1(new_n17511_), .B2(new_n17504_), .ZN(new_n17520_));
  NAND2_X1   g17328(.A1(new_n17133_), .A2(\asqrt[44] ), .ZN(new_n17521_));
  NOR4_X1    g17329(.A1(new_n17271_), .A2(\asqrt[44] ), .A3(new_n16908_), .A4(new_n17133_), .ZN(new_n17522_));
  XOR2_X1    g17330(.A1(new_n17522_), .A2(new_n17521_), .Z(new_n17523_));
  NAND2_X1   g17331(.A1(new_n17523_), .A2(new_n2728_), .ZN(new_n17524_));
  INV_X1     g17332(.I(new_n17524_), .ZN(new_n17525_));
  OAI21_X1   g17333(.A1(new_n17520_), .A2(new_n2941_), .B(new_n17525_), .ZN(new_n17526_));
  NAND2_X1   g17334(.A1(new_n17526_), .A2(new_n17519_), .ZN(new_n17527_));
  OAI22_X1   g17335(.A1(new_n17520_), .A2(new_n2941_), .B1(new_n17518_), .B2(new_n17512_), .ZN(new_n17528_));
  NOR4_X1    g17336(.A1(new_n17271_), .A2(\asqrt[45] ), .A3(new_n16915_), .A4(new_n16920_), .ZN(new_n17529_));
  AOI21_X1   g17337(.A1(new_n17521_), .A2(new_n17132_), .B(new_n2728_), .ZN(new_n17530_));
  NOR2_X1    g17338(.A1(new_n17529_), .A2(new_n17530_), .ZN(new_n17531_));
  NAND2_X1   g17339(.A1(new_n17531_), .A2(new_n2488_), .ZN(new_n17532_));
  AOI21_X1   g17340(.A1(new_n17528_), .A2(\asqrt[45] ), .B(new_n17532_), .ZN(new_n17533_));
  NOR2_X1    g17341(.A1(new_n17533_), .A2(new_n17527_), .ZN(new_n17534_));
  AOI22_X1   g17342(.A1(new_n17528_), .A2(\asqrt[45] ), .B1(new_n17526_), .B2(new_n17519_), .ZN(new_n17535_));
  NAND2_X1   g17343(.A1(new_n17140_), .A2(\asqrt[46] ), .ZN(new_n17536_));
  NOR4_X1    g17344(.A1(new_n17271_), .A2(\asqrt[46] ), .A3(new_n16923_), .A4(new_n17140_), .ZN(new_n17537_));
  XOR2_X1    g17345(.A1(new_n17537_), .A2(new_n17536_), .Z(new_n17538_));
  NAND2_X1   g17346(.A1(new_n17538_), .A2(new_n2253_), .ZN(new_n17539_));
  INV_X1     g17347(.I(new_n17539_), .ZN(new_n17540_));
  OAI21_X1   g17348(.A1(new_n17535_), .A2(new_n2488_), .B(new_n17540_), .ZN(new_n17541_));
  NAND2_X1   g17349(.A1(new_n17541_), .A2(new_n17534_), .ZN(new_n17542_));
  OAI22_X1   g17350(.A1(new_n17535_), .A2(new_n2488_), .B1(new_n17533_), .B2(new_n17527_), .ZN(new_n17543_));
  NOR4_X1    g17351(.A1(new_n17271_), .A2(\asqrt[47] ), .A3(new_n16930_), .A4(new_n16935_), .ZN(new_n17544_));
  AOI21_X1   g17352(.A1(new_n17536_), .A2(new_n17139_), .B(new_n2253_), .ZN(new_n17545_));
  NOR2_X1    g17353(.A1(new_n17544_), .A2(new_n17545_), .ZN(new_n17546_));
  NAND2_X1   g17354(.A1(new_n17546_), .A2(new_n2046_), .ZN(new_n17547_));
  AOI21_X1   g17355(.A1(new_n17543_), .A2(\asqrt[47] ), .B(new_n17547_), .ZN(new_n17548_));
  NOR2_X1    g17356(.A1(new_n17548_), .A2(new_n17542_), .ZN(new_n17549_));
  AOI22_X1   g17357(.A1(new_n17543_), .A2(\asqrt[47] ), .B1(new_n17541_), .B2(new_n17534_), .ZN(new_n17550_));
  NAND2_X1   g17358(.A1(new_n17147_), .A2(\asqrt[48] ), .ZN(new_n17551_));
  NOR4_X1    g17359(.A1(new_n17271_), .A2(\asqrt[48] ), .A3(new_n16938_), .A4(new_n17147_), .ZN(new_n17552_));
  XOR2_X1    g17360(.A1(new_n17552_), .A2(new_n17551_), .Z(new_n17553_));
  NAND2_X1   g17361(.A1(new_n17553_), .A2(new_n1854_), .ZN(new_n17554_));
  INV_X1     g17362(.I(new_n17554_), .ZN(new_n17555_));
  OAI21_X1   g17363(.A1(new_n17550_), .A2(new_n2046_), .B(new_n17555_), .ZN(new_n17556_));
  NAND2_X1   g17364(.A1(new_n17556_), .A2(new_n17549_), .ZN(new_n17557_));
  OAI22_X1   g17365(.A1(new_n17550_), .A2(new_n2046_), .B1(new_n17548_), .B2(new_n17542_), .ZN(new_n17558_));
  NAND2_X1   g17366(.A1(new_n16950_), .A2(\asqrt[49] ), .ZN(new_n17559_));
  NOR4_X1    g17367(.A1(new_n17271_), .A2(\asqrt[49] ), .A3(new_n16945_), .A4(new_n16950_), .ZN(new_n17560_));
  XOR2_X1    g17368(.A1(new_n17560_), .A2(new_n17559_), .Z(new_n17561_));
  NAND2_X1   g17369(.A1(new_n17561_), .A2(new_n1595_), .ZN(new_n17562_));
  AOI21_X1   g17370(.A1(new_n17558_), .A2(\asqrt[49] ), .B(new_n17562_), .ZN(new_n17563_));
  NOR2_X1    g17371(.A1(new_n17563_), .A2(new_n17557_), .ZN(new_n17564_));
  AOI22_X1   g17372(.A1(new_n17558_), .A2(\asqrt[49] ), .B1(new_n17556_), .B2(new_n17549_), .ZN(new_n17565_));
  NOR4_X1    g17373(.A1(new_n17271_), .A2(\asqrt[50] ), .A3(new_n16953_), .A4(new_n17154_), .ZN(new_n17566_));
  AOI21_X1   g17374(.A1(new_n17559_), .A2(new_n16949_), .B(new_n1595_), .ZN(new_n17567_));
  NOR2_X1    g17375(.A1(new_n17566_), .A2(new_n17567_), .ZN(new_n17568_));
  NAND2_X1   g17376(.A1(new_n17568_), .A2(new_n1436_), .ZN(new_n17569_));
  INV_X1     g17377(.I(new_n17569_), .ZN(new_n17570_));
  OAI21_X1   g17378(.A1(new_n17565_), .A2(new_n1595_), .B(new_n17570_), .ZN(new_n17571_));
  NAND2_X1   g17379(.A1(new_n17571_), .A2(new_n17564_), .ZN(new_n17572_));
  OAI22_X1   g17380(.A1(new_n17565_), .A2(new_n1595_), .B1(new_n17563_), .B2(new_n17557_), .ZN(new_n17573_));
  NAND2_X1   g17381(.A1(new_n16965_), .A2(\asqrt[51] ), .ZN(new_n17574_));
  NOR4_X1    g17382(.A1(new_n17271_), .A2(\asqrt[51] ), .A3(new_n16960_), .A4(new_n16965_), .ZN(new_n17575_));
  XOR2_X1    g17383(.A1(new_n17575_), .A2(new_n17574_), .Z(new_n17576_));
  NAND2_X1   g17384(.A1(new_n17576_), .A2(new_n1260_), .ZN(new_n17577_));
  AOI21_X1   g17385(.A1(new_n17573_), .A2(\asqrt[51] ), .B(new_n17577_), .ZN(new_n17578_));
  NOR2_X1    g17386(.A1(new_n17578_), .A2(new_n17572_), .ZN(new_n17579_));
  AOI22_X1   g17387(.A1(new_n17573_), .A2(\asqrt[51] ), .B1(new_n17571_), .B2(new_n17564_), .ZN(new_n17580_));
  NOR4_X1    g17388(.A1(new_n17271_), .A2(\asqrt[52] ), .A3(new_n16968_), .A4(new_n17161_), .ZN(new_n17581_));
  AOI21_X1   g17389(.A1(new_n17574_), .A2(new_n16964_), .B(new_n1260_), .ZN(new_n17582_));
  NOR2_X1    g17390(.A1(new_n17581_), .A2(new_n17582_), .ZN(new_n17583_));
  NAND2_X1   g17391(.A1(new_n17583_), .A2(new_n1096_), .ZN(new_n17584_));
  INV_X1     g17392(.I(new_n17584_), .ZN(new_n17585_));
  OAI21_X1   g17393(.A1(new_n17580_), .A2(new_n1260_), .B(new_n17585_), .ZN(new_n17586_));
  NAND2_X1   g17394(.A1(new_n17586_), .A2(new_n17579_), .ZN(new_n17587_));
  OAI22_X1   g17395(.A1(new_n17580_), .A2(new_n1260_), .B1(new_n17578_), .B2(new_n17572_), .ZN(new_n17588_));
  NOR4_X1    g17396(.A1(new_n17271_), .A2(\asqrt[53] ), .A3(new_n16975_), .A4(new_n16980_), .ZN(new_n17589_));
  XOR2_X1    g17397(.A1(new_n17589_), .A2(new_n17020_), .Z(new_n17590_));
  NAND2_X1   g17398(.A1(new_n17590_), .A2(new_n970_), .ZN(new_n17591_));
  AOI21_X1   g17399(.A1(new_n17588_), .A2(\asqrt[53] ), .B(new_n17591_), .ZN(new_n17592_));
  NOR2_X1    g17400(.A1(new_n17592_), .A2(new_n17587_), .ZN(new_n17593_));
  AOI22_X1   g17401(.A1(new_n17588_), .A2(\asqrt[53] ), .B1(new_n17586_), .B2(new_n17579_), .ZN(new_n17594_));
  NOR4_X1    g17402(.A1(new_n17271_), .A2(\asqrt[54] ), .A3(new_n16983_), .A4(new_n17168_), .ZN(new_n17595_));
  XNOR2_X1   g17403(.A1(new_n17595_), .A2(new_n17021_), .ZN(new_n17596_));
  NAND2_X1   g17404(.A1(new_n17596_), .A2(new_n825_), .ZN(new_n17597_));
  INV_X1     g17405(.I(new_n17597_), .ZN(new_n17598_));
  OAI21_X1   g17406(.A1(new_n17594_), .A2(new_n970_), .B(new_n17598_), .ZN(new_n17599_));
  NAND2_X1   g17407(.A1(new_n17599_), .A2(new_n17593_), .ZN(new_n17600_));
  OAI22_X1   g17408(.A1(new_n17594_), .A2(new_n970_), .B1(new_n17592_), .B2(new_n17587_), .ZN(new_n17601_));
  NOR4_X1    g17409(.A1(new_n17271_), .A2(\asqrt[55] ), .A3(new_n16989_), .A4(new_n16994_), .ZN(new_n17602_));
  XOR2_X1    g17410(.A1(new_n17602_), .A2(new_n17022_), .Z(new_n17603_));
  NAND2_X1   g17411(.A1(new_n17603_), .A2(new_n724_), .ZN(new_n17604_));
  AOI21_X1   g17412(.A1(new_n17601_), .A2(\asqrt[55] ), .B(new_n17604_), .ZN(new_n17605_));
  NOR2_X1    g17413(.A1(new_n17605_), .A2(new_n17600_), .ZN(new_n17606_));
  AOI22_X1   g17414(.A1(new_n17601_), .A2(\asqrt[55] ), .B1(new_n17599_), .B2(new_n17593_), .ZN(new_n17607_));
  NOR4_X1    g17415(.A1(new_n17271_), .A2(\asqrt[56] ), .A3(new_n16996_), .A4(new_n17175_), .ZN(new_n17608_));
  XOR2_X1    g17416(.A1(new_n17608_), .A2(new_n17188_), .Z(new_n17609_));
  NAND2_X1   g17417(.A1(new_n17609_), .A2(new_n587_), .ZN(new_n17610_));
  INV_X1     g17418(.I(new_n17610_), .ZN(new_n17611_));
  OAI21_X1   g17419(.A1(new_n17607_), .A2(new_n724_), .B(new_n17611_), .ZN(new_n17612_));
  NAND2_X1   g17420(.A1(new_n17612_), .A2(new_n17606_), .ZN(new_n17613_));
  OAI22_X1   g17421(.A1(new_n17607_), .A2(new_n724_), .B1(new_n17605_), .B2(new_n17600_), .ZN(new_n17614_));
  NOR4_X1    g17422(.A1(new_n17271_), .A2(\asqrt[57] ), .A3(new_n17002_), .A4(new_n17007_), .ZN(new_n17615_));
  XOR2_X1    g17423(.A1(new_n17615_), .A2(new_n17024_), .Z(new_n17616_));
  NAND2_X1   g17424(.A1(new_n17616_), .A2(new_n504_), .ZN(new_n17617_));
  AOI21_X1   g17425(.A1(new_n17614_), .A2(\asqrt[57] ), .B(new_n17617_), .ZN(new_n17618_));
  NOR2_X1    g17426(.A1(new_n17618_), .A2(new_n17613_), .ZN(new_n17619_));
  AOI22_X1   g17427(.A1(new_n17614_), .A2(\asqrt[57] ), .B1(new_n17612_), .B2(new_n17606_), .ZN(new_n17620_));
  NOR4_X1    g17428(.A1(new_n17271_), .A2(\asqrt[58] ), .A3(new_n17009_), .A4(new_n17182_), .ZN(new_n17621_));
  XOR2_X1    g17429(.A1(new_n17621_), .A2(new_n17190_), .Z(new_n17622_));
  NAND2_X1   g17430(.A1(new_n17622_), .A2(new_n376_), .ZN(new_n17623_));
  INV_X1     g17431(.I(new_n17623_), .ZN(new_n17624_));
  OAI21_X1   g17432(.A1(new_n17620_), .A2(new_n504_), .B(new_n17624_), .ZN(new_n17625_));
  NAND2_X1   g17433(.A1(new_n17625_), .A2(new_n17619_), .ZN(new_n17626_));
  OAI22_X1   g17434(.A1(new_n17620_), .A2(new_n504_), .B1(new_n17618_), .B2(new_n17613_), .ZN(new_n17627_));
  NOR4_X1    g17435(.A1(new_n17271_), .A2(\asqrt[59] ), .A3(new_n17015_), .A4(new_n17031_), .ZN(new_n17628_));
  XOR2_X1    g17436(.A1(new_n17628_), .A2(new_n17026_), .Z(new_n17629_));
  NAND2_X1   g17437(.A1(new_n17629_), .A2(new_n275_), .ZN(new_n17630_));
  AOI21_X1   g17438(.A1(new_n17627_), .A2(\asqrt[59] ), .B(new_n17630_), .ZN(new_n17631_));
  NOR2_X1    g17439(.A1(new_n17631_), .A2(new_n17626_), .ZN(new_n17632_));
  NAND2_X1   g17440(.A1(new_n17614_), .A2(\asqrt[57] ), .ZN(new_n17633_));
  AOI21_X1   g17441(.A1(new_n17633_), .A2(new_n17613_), .B(new_n504_), .ZN(new_n17634_));
  OAI21_X1   g17442(.A1(new_n17619_), .A2(new_n17634_), .B(\asqrt[59] ), .ZN(new_n17635_));
  AOI21_X1   g17443(.A1(new_n17626_), .A2(new_n17635_), .B(new_n275_), .ZN(new_n17636_));
  OAI21_X1   g17444(.A1(new_n17632_), .A2(new_n17636_), .B(\asqrt[61] ), .ZN(new_n17637_));
  AOI22_X1   g17445(.A1(new_n17627_), .A2(\asqrt[59] ), .B1(new_n17625_), .B2(new_n17619_), .ZN(new_n17638_));
  NOR4_X1    g17446(.A1(new_n17271_), .A2(\asqrt[60] ), .A3(new_n17028_), .A4(new_n17225_), .ZN(new_n17639_));
  XOR2_X1    g17447(.A1(new_n17639_), .A2(new_n17192_), .Z(new_n17640_));
  NAND2_X1   g17448(.A1(new_n17640_), .A2(new_n229_), .ZN(new_n17641_));
  INV_X1     g17449(.I(new_n17641_), .ZN(new_n17642_));
  OAI21_X1   g17450(.A1(new_n17638_), .A2(new_n275_), .B(new_n17642_), .ZN(new_n17643_));
  INV_X1     g17451(.I(new_n17240_), .ZN(new_n17644_));
  NOR2_X1    g17452(.A1(new_n17644_), .A2(\asqrt[62] ), .ZN(new_n17645_));
  INV_X1     g17453(.I(new_n17645_), .ZN(new_n17646_));
  NAND3_X1   g17454(.A1(new_n17643_), .A2(new_n17632_), .A3(new_n17646_), .ZN(new_n17647_));
  OAI21_X1   g17455(.A1(new_n17647_), .A2(new_n17637_), .B(new_n17242_), .ZN(new_n17648_));
  NAND3_X1   g17456(.A1(new_n17271_), .A2(new_n17224_), .A3(new_n17274_), .ZN(new_n17649_));
  AOI21_X1   g17457(.A1(new_n17649_), .A2(new_n17216_), .B(\asqrt[63] ), .ZN(new_n17650_));
  INV_X1     g17458(.I(new_n17650_), .ZN(new_n17651_));
  OAI21_X1   g17459(.A1(new_n17648_), .A2(new_n17651_), .B(new_n17237_), .ZN(new_n17652_));
  OAI22_X1   g17460(.A1(new_n17638_), .A2(new_n275_), .B1(new_n17631_), .B2(new_n17626_), .ZN(new_n17653_));
  AOI22_X1   g17461(.A1(new_n17653_), .A2(\asqrt[61] ), .B1(new_n17643_), .B2(new_n17632_), .ZN(new_n17654_));
  NAND4_X1   g17462(.A1(new_n17654_), .A2(new_n196_), .A3(new_n17237_), .A4(new_n17644_), .ZN(new_n17655_));
  INV_X1     g17463(.I(\a[18] ), .ZN(new_n17656_));
  NAND3_X1   g17464(.A1(new_n17265_), .A2(new_n17209_), .A3(new_n17231_), .ZN(new_n17657_));
  INV_X1     g17465(.I(new_n17657_), .ZN(new_n17658_));
  NAND2_X1   g17466(.A1(new_n17256_), .A2(new_n17224_), .ZN(new_n17659_));
  XOR2_X1    g17467(.A1(new_n17256_), .A2(\asqrt[63] ), .Z(new_n17660_));
  AOI21_X1   g17468(.A1(\asqrt[11] ), .A2(new_n17659_), .B(new_n17660_), .ZN(new_n17661_));
  NOR2_X1    g17469(.A1(new_n17658_), .A2(new_n17661_), .ZN(new_n17662_));
  NOR2_X1    g17470(.A1(\a[16] ), .A2(\a[17] ), .ZN(new_n17663_));
  INV_X1     g17471(.I(new_n17663_), .ZN(new_n17664_));
  NOR3_X1    g17472(.A1(new_n17662_), .A2(new_n17656_), .A3(new_n17664_), .ZN(new_n17665_));
  NAND3_X1   g17473(.A1(new_n17652_), .A2(new_n17655_), .A3(new_n17665_), .ZN(new_n17666_));
  XOR2_X1    g17474(.A1(new_n17666_), .A2(\a[19] ), .Z(new_n17667_));
  INV_X1     g17475(.I(\a[19] ), .ZN(new_n17668_));
  NOR2_X1    g17476(.A1(new_n17654_), .A2(new_n196_), .ZN(new_n17669_));
  INV_X1     g17477(.I(new_n17251_), .ZN(new_n17670_));
  AOI21_X1   g17478(.A1(new_n17262_), .A2(new_n17670_), .B(new_n17253_), .ZN(new_n17671_));
  NOR3_X1    g17479(.A1(new_n17250_), .A2(new_n17243_), .A3(new_n17248_), .ZN(new_n17672_));
  NOR2_X1    g17480(.A1(new_n17672_), .A2(new_n17671_), .ZN(new_n17673_));
  NOR3_X1    g17481(.A1(new_n17284_), .A2(new_n16004_), .A3(\asqrt[11] ), .ZN(new_n17674_));
  AOI21_X1   g17482(.A1(new_n17278_), .A2(new_n16003_), .B(new_n17271_), .ZN(new_n17675_));
  NOR4_X1    g17483(.A1(new_n17675_), .A2(new_n17674_), .A3(\asqrt[13] ), .A4(new_n17269_), .ZN(new_n17676_));
  NOR2_X1    g17484(.A1(new_n17676_), .A2(new_n17673_), .ZN(new_n17677_));
  NOR3_X1    g17485(.A1(new_n17672_), .A2(new_n17671_), .A3(new_n17269_), .ZN(new_n17678_));
  NOR3_X1    g17486(.A1(new_n17271_), .A2(new_n16617_), .A3(new_n17295_), .ZN(new_n17679_));
  AOI21_X1   g17487(.A1(\asqrt[11] ), .A2(new_n17293_), .B(new_n16618_), .ZN(new_n17680_));
  NOR3_X1    g17488(.A1(new_n17680_), .A2(new_n17679_), .A3(\asqrt[14] ), .ZN(new_n17681_));
  OAI21_X1   g17489(.A1(new_n17678_), .A2(new_n16060_), .B(new_n17681_), .ZN(new_n17682_));
  NAND2_X1   g17490(.A1(new_n17677_), .A2(new_n17682_), .ZN(new_n17683_));
  OAI22_X1   g17491(.A1(new_n17676_), .A2(new_n17673_), .B1(new_n16060_), .B2(new_n17678_), .ZN(new_n17684_));
  INV_X1     g17492(.I(new_n17304_), .ZN(new_n17685_));
  AOI21_X1   g17493(.A1(new_n17684_), .A2(\asqrt[14] ), .B(new_n17685_), .ZN(new_n17686_));
  NOR2_X1    g17494(.A1(new_n17686_), .A2(new_n17683_), .ZN(new_n17687_));
  AOI22_X1   g17495(.A1(new_n17684_), .A2(\asqrt[14] ), .B1(new_n17677_), .B2(new_n17682_), .ZN(new_n17688_));
  INV_X1     g17496(.I(new_n17311_), .ZN(new_n17689_));
  OAI21_X1   g17497(.A1(new_n17688_), .A2(new_n14871_), .B(new_n17689_), .ZN(new_n17690_));
  NAND2_X1   g17498(.A1(new_n17690_), .A2(new_n17687_), .ZN(new_n17691_));
  OAI22_X1   g17499(.A1(new_n17688_), .A2(new_n14871_), .B1(new_n17686_), .B2(new_n17683_), .ZN(new_n17692_));
  AOI21_X1   g17500(.A1(new_n17692_), .A2(\asqrt[16] ), .B(new_n17318_), .ZN(new_n17693_));
  NOR2_X1    g17501(.A1(new_n17693_), .A2(new_n17691_), .ZN(new_n17694_));
  AOI22_X1   g17502(.A1(new_n17692_), .A2(\asqrt[16] ), .B1(new_n17690_), .B2(new_n17687_), .ZN(new_n17695_));
  INV_X1     g17503(.I(new_n17325_), .ZN(new_n17696_));
  OAI21_X1   g17504(.A1(new_n17695_), .A2(new_n13760_), .B(new_n17696_), .ZN(new_n17697_));
  NAND2_X1   g17505(.A1(new_n17697_), .A2(new_n17694_), .ZN(new_n17698_));
  OAI22_X1   g17506(.A1(new_n17695_), .A2(new_n13760_), .B1(new_n17693_), .B2(new_n17691_), .ZN(new_n17699_));
  AOI21_X1   g17507(.A1(new_n17699_), .A2(\asqrt[18] ), .B(new_n17331_), .ZN(new_n17700_));
  NOR2_X1    g17508(.A1(new_n17700_), .A2(new_n17698_), .ZN(new_n17701_));
  AOI22_X1   g17509(.A1(new_n17699_), .A2(\asqrt[18] ), .B1(new_n17697_), .B2(new_n17694_), .ZN(new_n17702_));
  INV_X1     g17510(.I(new_n17338_), .ZN(new_n17703_));
  OAI21_X1   g17511(.A1(new_n17702_), .A2(new_n12657_), .B(new_n17703_), .ZN(new_n17704_));
  NAND2_X1   g17512(.A1(new_n17704_), .A2(new_n17701_), .ZN(new_n17705_));
  OAI22_X1   g17513(.A1(new_n17702_), .A2(new_n12657_), .B1(new_n17700_), .B2(new_n17698_), .ZN(new_n17706_));
  AOI21_X1   g17514(.A1(new_n17706_), .A2(\asqrt[20] ), .B(new_n17344_), .ZN(new_n17707_));
  NOR2_X1    g17515(.A1(new_n17707_), .A2(new_n17705_), .ZN(new_n17708_));
  AOI22_X1   g17516(.A1(new_n17706_), .A2(\asqrt[20] ), .B1(new_n17704_), .B2(new_n17701_), .ZN(new_n17709_));
  INV_X1     g17517(.I(new_n17352_), .ZN(new_n17710_));
  OAI21_X1   g17518(.A1(new_n17709_), .A2(new_n11631_), .B(new_n17710_), .ZN(new_n17711_));
  NAND2_X1   g17519(.A1(new_n17711_), .A2(new_n17708_), .ZN(new_n17712_));
  OAI22_X1   g17520(.A1(new_n17709_), .A2(new_n11631_), .B1(new_n17707_), .B2(new_n17705_), .ZN(new_n17713_));
  AOI21_X1   g17521(.A1(new_n17713_), .A2(\asqrt[22] ), .B(new_n17359_), .ZN(new_n17714_));
  NOR2_X1    g17522(.A1(new_n17714_), .A2(new_n17712_), .ZN(new_n17715_));
  AOI22_X1   g17523(.A1(new_n17713_), .A2(\asqrt[22] ), .B1(new_n17711_), .B2(new_n17708_), .ZN(new_n17716_));
  INV_X1     g17524(.I(new_n17367_), .ZN(new_n17717_));
  OAI21_X1   g17525(.A1(new_n17716_), .A2(new_n10614_), .B(new_n17717_), .ZN(new_n17718_));
  NAND2_X1   g17526(.A1(new_n17718_), .A2(new_n17715_), .ZN(new_n17719_));
  OAI22_X1   g17527(.A1(new_n17716_), .A2(new_n10614_), .B1(new_n17714_), .B2(new_n17712_), .ZN(new_n17720_));
  AOI21_X1   g17528(.A1(new_n17720_), .A2(\asqrt[24] ), .B(new_n17374_), .ZN(new_n17721_));
  NOR2_X1    g17529(.A1(new_n17721_), .A2(new_n17719_), .ZN(new_n17722_));
  AOI22_X1   g17530(.A1(new_n17720_), .A2(\asqrt[24] ), .B1(new_n17718_), .B2(new_n17715_), .ZN(new_n17723_));
  INV_X1     g17531(.I(new_n17382_), .ZN(new_n17724_));
  OAI21_X1   g17532(.A1(new_n17723_), .A2(new_n9672_), .B(new_n17724_), .ZN(new_n17725_));
  NAND2_X1   g17533(.A1(new_n17725_), .A2(new_n17722_), .ZN(new_n17726_));
  OAI22_X1   g17534(.A1(new_n17723_), .A2(new_n9672_), .B1(new_n17721_), .B2(new_n17719_), .ZN(new_n17727_));
  AOI21_X1   g17535(.A1(new_n17727_), .A2(\asqrt[26] ), .B(new_n17389_), .ZN(new_n17728_));
  NOR2_X1    g17536(.A1(new_n17728_), .A2(new_n17726_), .ZN(new_n17729_));
  AOI22_X1   g17537(.A1(new_n17727_), .A2(\asqrt[26] ), .B1(new_n17725_), .B2(new_n17722_), .ZN(new_n17730_));
  INV_X1     g17538(.I(new_n17397_), .ZN(new_n17731_));
  OAI21_X1   g17539(.A1(new_n17730_), .A2(new_n8763_), .B(new_n17731_), .ZN(new_n17732_));
  NAND2_X1   g17540(.A1(new_n17732_), .A2(new_n17729_), .ZN(new_n17733_));
  OAI22_X1   g17541(.A1(new_n17730_), .A2(new_n8763_), .B1(new_n17728_), .B2(new_n17726_), .ZN(new_n17734_));
  AOI21_X1   g17542(.A1(new_n17734_), .A2(\asqrt[28] ), .B(new_n17404_), .ZN(new_n17735_));
  NOR2_X1    g17543(.A1(new_n17735_), .A2(new_n17733_), .ZN(new_n17736_));
  AOI22_X1   g17544(.A1(new_n17734_), .A2(\asqrt[28] ), .B1(new_n17732_), .B2(new_n17729_), .ZN(new_n17737_));
  INV_X1     g17545(.I(new_n17412_), .ZN(new_n17738_));
  OAI21_X1   g17546(.A1(new_n17737_), .A2(new_n7931_), .B(new_n17738_), .ZN(new_n17739_));
  NAND2_X1   g17547(.A1(new_n17739_), .A2(new_n17736_), .ZN(new_n17740_));
  OAI22_X1   g17548(.A1(new_n17737_), .A2(new_n7931_), .B1(new_n17735_), .B2(new_n17733_), .ZN(new_n17741_));
  AOI21_X1   g17549(.A1(new_n17741_), .A2(\asqrt[30] ), .B(new_n17419_), .ZN(new_n17742_));
  NOR2_X1    g17550(.A1(new_n17742_), .A2(new_n17740_), .ZN(new_n17743_));
  AOI22_X1   g17551(.A1(new_n17741_), .A2(\asqrt[30] ), .B1(new_n17739_), .B2(new_n17736_), .ZN(new_n17744_));
  INV_X1     g17552(.I(new_n17427_), .ZN(new_n17745_));
  OAI21_X1   g17553(.A1(new_n17744_), .A2(new_n7110_), .B(new_n17745_), .ZN(new_n17746_));
  NAND2_X1   g17554(.A1(new_n17746_), .A2(new_n17743_), .ZN(new_n17747_));
  OAI22_X1   g17555(.A1(new_n17744_), .A2(new_n7110_), .B1(new_n17742_), .B2(new_n17740_), .ZN(new_n17748_));
  AOI21_X1   g17556(.A1(new_n17748_), .A2(\asqrt[32] ), .B(new_n17434_), .ZN(new_n17749_));
  NOR2_X1    g17557(.A1(new_n17749_), .A2(new_n17747_), .ZN(new_n17750_));
  AOI22_X1   g17558(.A1(new_n17748_), .A2(\asqrt[32] ), .B1(new_n17746_), .B2(new_n17743_), .ZN(new_n17751_));
  INV_X1     g17559(.I(new_n17442_), .ZN(new_n17752_));
  OAI21_X1   g17560(.A1(new_n17751_), .A2(new_n6365_), .B(new_n17752_), .ZN(new_n17753_));
  NAND2_X1   g17561(.A1(new_n17753_), .A2(new_n17750_), .ZN(new_n17754_));
  OAI22_X1   g17562(.A1(new_n17751_), .A2(new_n6365_), .B1(new_n17749_), .B2(new_n17747_), .ZN(new_n17755_));
  AOI21_X1   g17563(.A1(new_n17755_), .A2(\asqrt[34] ), .B(new_n17449_), .ZN(new_n17756_));
  NOR2_X1    g17564(.A1(new_n17756_), .A2(new_n17754_), .ZN(new_n17757_));
  AOI22_X1   g17565(.A1(new_n17755_), .A2(\asqrt[34] ), .B1(new_n17753_), .B2(new_n17750_), .ZN(new_n17758_));
  INV_X1     g17566(.I(new_n17457_), .ZN(new_n17759_));
  OAI21_X1   g17567(.A1(new_n17758_), .A2(new_n5626_), .B(new_n17759_), .ZN(new_n17760_));
  NAND2_X1   g17568(.A1(new_n17760_), .A2(new_n17757_), .ZN(new_n17761_));
  OAI22_X1   g17569(.A1(new_n17758_), .A2(new_n5626_), .B1(new_n17756_), .B2(new_n17754_), .ZN(new_n17762_));
  AOI21_X1   g17570(.A1(new_n17762_), .A2(\asqrt[36] ), .B(new_n17464_), .ZN(new_n17763_));
  NOR2_X1    g17571(.A1(new_n17763_), .A2(new_n17761_), .ZN(new_n17764_));
  AOI22_X1   g17572(.A1(new_n17762_), .A2(\asqrt[36] ), .B1(new_n17760_), .B2(new_n17757_), .ZN(new_n17765_));
  INV_X1     g17573(.I(new_n17472_), .ZN(new_n17766_));
  OAI21_X1   g17574(.A1(new_n17765_), .A2(new_n4973_), .B(new_n17766_), .ZN(new_n17767_));
  NAND2_X1   g17575(.A1(new_n17767_), .A2(new_n17764_), .ZN(new_n17768_));
  OAI22_X1   g17576(.A1(new_n17765_), .A2(new_n4973_), .B1(new_n17763_), .B2(new_n17761_), .ZN(new_n17769_));
  AOI21_X1   g17577(.A1(new_n17769_), .A2(\asqrt[38] ), .B(new_n17479_), .ZN(new_n17770_));
  NOR2_X1    g17578(.A1(new_n17770_), .A2(new_n17768_), .ZN(new_n17771_));
  AOI22_X1   g17579(.A1(new_n17769_), .A2(\asqrt[38] ), .B1(new_n17767_), .B2(new_n17764_), .ZN(new_n17772_));
  INV_X1     g17580(.I(new_n17487_), .ZN(new_n17773_));
  OAI21_X1   g17581(.A1(new_n17772_), .A2(new_n4330_), .B(new_n17773_), .ZN(new_n17774_));
  NAND2_X1   g17582(.A1(new_n17774_), .A2(new_n17771_), .ZN(new_n17775_));
  OAI22_X1   g17583(.A1(new_n17772_), .A2(new_n4330_), .B1(new_n17770_), .B2(new_n17768_), .ZN(new_n17776_));
  AOI21_X1   g17584(.A1(new_n17776_), .A2(\asqrt[40] ), .B(new_n17494_), .ZN(new_n17777_));
  NOR2_X1    g17585(.A1(new_n17777_), .A2(new_n17775_), .ZN(new_n17778_));
  AOI22_X1   g17586(.A1(new_n17776_), .A2(\asqrt[40] ), .B1(new_n17774_), .B2(new_n17771_), .ZN(new_n17779_));
  INV_X1     g17587(.I(new_n17502_), .ZN(new_n17780_));
  OAI21_X1   g17588(.A1(new_n17779_), .A2(new_n3760_), .B(new_n17780_), .ZN(new_n17781_));
  NAND2_X1   g17589(.A1(new_n17781_), .A2(new_n17778_), .ZN(new_n17782_));
  OAI22_X1   g17590(.A1(new_n17779_), .A2(new_n3760_), .B1(new_n17777_), .B2(new_n17775_), .ZN(new_n17783_));
  AOI21_X1   g17591(.A1(new_n17783_), .A2(\asqrt[42] ), .B(new_n17509_), .ZN(new_n17784_));
  NOR2_X1    g17592(.A1(new_n17784_), .A2(new_n17782_), .ZN(new_n17785_));
  AOI22_X1   g17593(.A1(new_n17783_), .A2(\asqrt[42] ), .B1(new_n17781_), .B2(new_n17778_), .ZN(new_n17786_));
  INV_X1     g17594(.I(new_n17517_), .ZN(new_n17787_));
  OAI21_X1   g17595(.A1(new_n17786_), .A2(new_n3208_), .B(new_n17787_), .ZN(new_n17788_));
  NAND2_X1   g17596(.A1(new_n17788_), .A2(new_n17785_), .ZN(new_n17789_));
  OAI22_X1   g17597(.A1(new_n17786_), .A2(new_n3208_), .B1(new_n17784_), .B2(new_n17782_), .ZN(new_n17790_));
  AOI21_X1   g17598(.A1(new_n17790_), .A2(\asqrt[44] ), .B(new_n17524_), .ZN(new_n17791_));
  NOR2_X1    g17599(.A1(new_n17791_), .A2(new_n17789_), .ZN(new_n17792_));
  AOI22_X1   g17600(.A1(new_n17790_), .A2(\asqrt[44] ), .B1(new_n17788_), .B2(new_n17785_), .ZN(new_n17793_));
  INV_X1     g17601(.I(new_n17532_), .ZN(new_n17794_));
  OAI21_X1   g17602(.A1(new_n17793_), .A2(new_n2728_), .B(new_n17794_), .ZN(new_n17795_));
  NAND2_X1   g17603(.A1(new_n17795_), .A2(new_n17792_), .ZN(new_n17796_));
  OAI22_X1   g17604(.A1(new_n17793_), .A2(new_n2728_), .B1(new_n17791_), .B2(new_n17789_), .ZN(new_n17797_));
  AOI21_X1   g17605(.A1(new_n17797_), .A2(\asqrt[46] ), .B(new_n17539_), .ZN(new_n17798_));
  NOR2_X1    g17606(.A1(new_n17798_), .A2(new_n17796_), .ZN(new_n17799_));
  AOI22_X1   g17607(.A1(new_n17797_), .A2(\asqrt[46] ), .B1(new_n17795_), .B2(new_n17792_), .ZN(new_n17800_));
  INV_X1     g17608(.I(new_n17547_), .ZN(new_n17801_));
  OAI21_X1   g17609(.A1(new_n17800_), .A2(new_n2253_), .B(new_n17801_), .ZN(new_n17802_));
  NAND2_X1   g17610(.A1(new_n17802_), .A2(new_n17799_), .ZN(new_n17803_));
  OAI22_X1   g17611(.A1(new_n17800_), .A2(new_n2253_), .B1(new_n17798_), .B2(new_n17796_), .ZN(new_n17804_));
  AOI21_X1   g17612(.A1(new_n17804_), .A2(\asqrt[48] ), .B(new_n17554_), .ZN(new_n17805_));
  NOR2_X1    g17613(.A1(new_n17805_), .A2(new_n17803_), .ZN(new_n17806_));
  AOI22_X1   g17614(.A1(new_n17804_), .A2(\asqrt[48] ), .B1(new_n17802_), .B2(new_n17799_), .ZN(new_n17807_));
  INV_X1     g17615(.I(new_n17562_), .ZN(new_n17808_));
  OAI21_X1   g17616(.A1(new_n17807_), .A2(new_n1854_), .B(new_n17808_), .ZN(new_n17809_));
  NAND2_X1   g17617(.A1(new_n17809_), .A2(new_n17806_), .ZN(new_n17810_));
  OAI22_X1   g17618(.A1(new_n17807_), .A2(new_n1854_), .B1(new_n17805_), .B2(new_n17803_), .ZN(new_n17811_));
  AOI21_X1   g17619(.A1(new_n17811_), .A2(\asqrt[50] ), .B(new_n17569_), .ZN(new_n17812_));
  NOR2_X1    g17620(.A1(new_n17812_), .A2(new_n17810_), .ZN(new_n17813_));
  AOI22_X1   g17621(.A1(new_n17811_), .A2(\asqrt[50] ), .B1(new_n17809_), .B2(new_n17806_), .ZN(new_n17814_));
  INV_X1     g17622(.I(new_n17577_), .ZN(new_n17815_));
  OAI21_X1   g17623(.A1(new_n17814_), .A2(new_n1436_), .B(new_n17815_), .ZN(new_n17816_));
  NAND2_X1   g17624(.A1(new_n17816_), .A2(new_n17813_), .ZN(new_n17817_));
  OAI22_X1   g17625(.A1(new_n17814_), .A2(new_n1436_), .B1(new_n17812_), .B2(new_n17810_), .ZN(new_n17818_));
  AOI21_X1   g17626(.A1(new_n17818_), .A2(\asqrt[52] ), .B(new_n17584_), .ZN(new_n17819_));
  NOR2_X1    g17627(.A1(new_n17819_), .A2(new_n17817_), .ZN(new_n17820_));
  AOI22_X1   g17628(.A1(new_n17818_), .A2(\asqrt[52] ), .B1(new_n17816_), .B2(new_n17813_), .ZN(new_n17821_));
  INV_X1     g17629(.I(new_n17591_), .ZN(new_n17822_));
  OAI21_X1   g17630(.A1(new_n17821_), .A2(new_n1096_), .B(new_n17822_), .ZN(new_n17823_));
  NAND2_X1   g17631(.A1(new_n17823_), .A2(new_n17820_), .ZN(new_n17824_));
  OAI22_X1   g17632(.A1(new_n17821_), .A2(new_n1096_), .B1(new_n17819_), .B2(new_n17817_), .ZN(new_n17825_));
  AOI21_X1   g17633(.A1(new_n17825_), .A2(\asqrt[54] ), .B(new_n17597_), .ZN(new_n17826_));
  NOR2_X1    g17634(.A1(new_n17826_), .A2(new_n17824_), .ZN(new_n17827_));
  AOI22_X1   g17635(.A1(new_n17825_), .A2(\asqrt[54] ), .B1(new_n17823_), .B2(new_n17820_), .ZN(new_n17828_));
  INV_X1     g17636(.I(new_n17604_), .ZN(new_n17829_));
  OAI21_X1   g17637(.A1(new_n17828_), .A2(new_n825_), .B(new_n17829_), .ZN(new_n17830_));
  NAND2_X1   g17638(.A1(new_n17830_), .A2(new_n17827_), .ZN(new_n17831_));
  OAI22_X1   g17639(.A1(new_n17828_), .A2(new_n825_), .B1(new_n17826_), .B2(new_n17824_), .ZN(new_n17832_));
  AOI21_X1   g17640(.A1(new_n17832_), .A2(\asqrt[56] ), .B(new_n17610_), .ZN(new_n17833_));
  NOR2_X1    g17641(.A1(new_n17833_), .A2(new_n17831_), .ZN(new_n17834_));
  AOI22_X1   g17642(.A1(new_n17832_), .A2(\asqrt[56] ), .B1(new_n17830_), .B2(new_n17827_), .ZN(new_n17835_));
  INV_X1     g17643(.I(new_n17617_), .ZN(new_n17836_));
  OAI21_X1   g17644(.A1(new_n17835_), .A2(new_n587_), .B(new_n17836_), .ZN(new_n17837_));
  NAND2_X1   g17645(.A1(new_n17837_), .A2(new_n17834_), .ZN(new_n17838_));
  OAI22_X1   g17646(.A1(new_n17835_), .A2(new_n587_), .B1(new_n17833_), .B2(new_n17831_), .ZN(new_n17839_));
  AOI21_X1   g17647(.A1(new_n17839_), .A2(\asqrt[58] ), .B(new_n17623_), .ZN(new_n17840_));
  NOR2_X1    g17648(.A1(new_n17840_), .A2(new_n17838_), .ZN(new_n17841_));
  AOI22_X1   g17649(.A1(new_n17839_), .A2(\asqrt[58] ), .B1(new_n17837_), .B2(new_n17834_), .ZN(new_n17842_));
  INV_X1     g17650(.I(new_n17630_), .ZN(new_n17843_));
  OAI21_X1   g17651(.A1(new_n17842_), .A2(new_n376_), .B(new_n17843_), .ZN(new_n17844_));
  NAND2_X1   g17652(.A1(new_n17844_), .A2(new_n17841_), .ZN(new_n17845_));
  OAI22_X1   g17653(.A1(new_n17842_), .A2(new_n376_), .B1(new_n17840_), .B2(new_n17838_), .ZN(new_n17846_));
  AOI22_X1   g17654(.A1(new_n17846_), .A2(\asqrt[60] ), .B1(new_n17844_), .B2(new_n17841_), .ZN(new_n17847_));
  AOI21_X1   g17655(.A1(new_n17846_), .A2(\asqrt[60] ), .B(new_n17641_), .ZN(new_n17848_));
  OAI22_X1   g17656(.A1(new_n17847_), .A2(new_n229_), .B1(new_n17848_), .B2(new_n17845_), .ZN(new_n17849_));
  NOR2_X1    g17657(.A1(new_n17849_), .A2(\asqrt[62] ), .ZN(new_n17850_));
  NOR4_X1    g17658(.A1(new_n17849_), .A2(\asqrt[62] ), .A3(new_n17236_), .A4(new_n17240_), .ZN(new_n17851_));
  NAND2_X1   g17659(.A1(new_n17851_), .A2(new_n17661_), .ZN(new_n17852_));
  NOR3_X1    g17660(.A1(new_n17852_), .A2(new_n17657_), .A3(new_n17652_), .ZN(\asqrt[10] ));
  NAND4_X1   g17661(.A1(\asqrt[10] ), .A2(new_n17644_), .A3(new_n17669_), .A4(new_n17850_), .ZN(new_n17854_));
  OAI21_X1   g17662(.A1(new_n17849_), .A2(\asqrt[62] ), .B(new_n17240_), .ZN(new_n17855_));
  OAI21_X1   g17663(.A1(\asqrt[10] ), .A2(new_n17855_), .B(new_n17669_), .ZN(new_n17856_));
  NAND2_X1   g17664(.A1(new_n17854_), .A2(new_n17856_), .ZN(new_n17857_));
  INV_X1     g17665(.I(new_n17857_), .ZN(new_n17858_));
  NAND2_X1   g17666(.A1(new_n17839_), .A2(\asqrt[58] ), .ZN(new_n17859_));
  AOI21_X1   g17667(.A1(new_n17859_), .A2(new_n17838_), .B(new_n376_), .ZN(new_n17860_));
  OAI21_X1   g17668(.A1(new_n17841_), .A2(new_n17860_), .B(\asqrt[60] ), .ZN(new_n17861_));
  AOI21_X1   g17669(.A1(new_n17845_), .A2(new_n17861_), .B(new_n229_), .ZN(new_n17862_));
  NOR3_X1    g17670(.A1(new_n17653_), .A2(\asqrt[61] ), .A3(new_n17640_), .ZN(new_n17863_));
  NAND2_X1   g17671(.A1(\asqrt[10] ), .A2(new_n17863_), .ZN(new_n17864_));
  XOR2_X1    g17672(.A1(new_n17864_), .A2(new_n17862_), .Z(new_n17865_));
  NOR2_X1    g17673(.A1(new_n17865_), .A2(new_n196_), .ZN(new_n17866_));
  INV_X1     g17674(.I(new_n17866_), .ZN(new_n17867_));
  INV_X1     g17675(.I(\a[20] ), .ZN(new_n17868_));
  NOR2_X1    g17676(.A1(\a[18] ), .A2(\a[19] ), .ZN(new_n17869_));
  INV_X1     g17677(.I(new_n17869_), .ZN(new_n17870_));
  NOR3_X1    g17678(.A1(new_n17276_), .A2(new_n17868_), .A3(new_n17870_), .ZN(new_n17871_));
  NAND2_X1   g17679(.A1(new_n17282_), .A2(new_n17871_), .ZN(new_n17872_));
  XOR2_X1    g17680(.A1(new_n17872_), .A2(\a[21] ), .Z(new_n17873_));
  INV_X1     g17681(.I(\a[21] ), .ZN(new_n17874_));
  NOR4_X1    g17682(.A1(new_n17852_), .A2(new_n17874_), .A3(new_n17657_), .A4(new_n17652_), .ZN(new_n17875_));
  NOR2_X1    g17683(.A1(new_n17874_), .A2(\a[20] ), .ZN(new_n17876_));
  OAI21_X1   g17684(.A1(new_n17875_), .A2(new_n17876_), .B(new_n17873_), .ZN(new_n17877_));
  INV_X1     g17685(.I(new_n17873_), .ZN(new_n17878_));
  NOR3_X1    g17686(.A1(new_n17848_), .A2(new_n17845_), .A3(new_n17645_), .ZN(new_n17879_));
  AOI21_X1   g17687(.A1(new_n17879_), .A2(new_n17862_), .B(new_n17241_), .ZN(new_n17880_));
  AOI21_X1   g17688(.A1(new_n17880_), .A2(new_n17650_), .B(new_n17236_), .ZN(new_n17881_));
  INV_X1     g17689(.I(new_n17661_), .ZN(new_n17882_));
  NOR2_X1    g17690(.A1(new_n17655_), .A2(new_n17882_), .ZN(new_n17883_));
  NAND4_X1   g17691(.A1(new_n17883_), .A2(\a[21] ), .A3(new_n17881_), .A4(new_n17658_), .ZN(new_n17884_));
  NAND3_X1   g17692(.A1(new_n17884_), .A2(\a[20] ), .A3(new_n17878_), .ZN(new_n17885_));
  NAND2_X1   g17693(.A1(new_n17877_), .A2(new_n17885_), .ZN(new_n17886_));
  NOR2_X1    g17694(.A1(new_n17852_), .A2(new_n17652_), .ZN(new_n17887_));
  NOR4_X1    g17695(.A1(new_n17230_), .A2(new_n17224_), .A3(new_n17273_), .A4(new_n17231_), .ZN(new_n17888_));
  NAND2_X1   g17696(.A1(\asqrt[11] ), .A2(\a[20] ), .ZN(new_n17889_));
  XOR2_X1    g17697(.A1(new_n17889_), .A2(new_n17888_), .Z(new_n17890_));
  NOR2_X1    g17698(.A1(new_n17890_), .A2(new_n17870_), .ZN(new_n17891_));
  INV_X1     g17699(.I(new_n17891_), .ZN(new_n17892_));
  NAND3_X1   g17700(.A1(new_n17883_), .A2(new_n17658_), .A3(new_n17881_), .ZN(new_n17893_));
  NAND2_X1   g17701(.A1(new_n17662_), .A2(\asqrt[11] ), .ZN(new_n17894_));
  INV_X1     g17702(.I(new_n17894_), .ZN(new_n17895_));
  NAND3_X1   g17703(.A1(new_n17652_), .A2(new_n17655_), .A3(new_n17895_), .ZN(new_n17896_));
  NAND2_X1   g17704(.A1(new_n17896_), .A2(new_n17243_), .ZN(new_n17897_));
  NAND3_X1   g17705(.A1(new_n17897_), .A2(new_n17244_), .A3(new_n17893_), .ZN(new_n17898_));
  NOR3_X1    g17706(.A1(new_n17881_), .A2(new_n17851_), .A3(new_n17894_), .ZN(new_n17899_));
  OAI21_X1   g17707(.A1(new_n17899_), .A2(\a[22] ), .B(new_n17244_), .ZN(new_n17900_));
  NAND2_X1   g17708(.A1(new_n17900_), .A2(\asqrt[10] ), .ZN(new_n17901_));
  NAND4_X1   g17709(.A1(new_n17901_), .A2(new_n16619_), .A3(new_n17898_), .A4(new_n17892_), .ZN(new_n17902_));
  NAND2_X1   g17710(.A1(new_n17902_), .A2(new_n17886_), .ZN(new_n17903_));
  NAND3_X1   g17711(.A1(new_n17877_), .A2(new_n17885_), .A3(new_n17892_), .ZN(new_n17904_));
  AOI21_X1   g17712(.A1(\asqrt[11] ), .A2(new_n17243_), .B(\a[23] ), .ZN(new_n17905_));
  NOR2_X1    g17713(.A1(new_n17262_), .A2(\a[22] ), .ZN(new_n17906_));
  AOI21_X1   g17714(.A1(\asqrt[11] ), .A2(\a[22] ), .B(new_n17247_), .ZN(new_n17907_));
  OAI21_X1   g17715(.A1(new_n17906_), .A2(new_n17905_), .B(new_n17907_), .ZN(new_n17908_));
  INV_X1     g17716(.I(new_n17908_), .ZN(new_n17909_));
  NAND3_X1   g17717(.A1(\asqrt[10] ), .A2(new_n17270_), .A3(new_n17909_), .ZN(new_n17910_));
  OAI21_X1   g17718(.A1(new_n17893_), .A2(new_n17908_), .B(new_n17269_), .ZN(new_n17911_));
  NAND3_X1   g17719(.A1(new_n17910_), .A2(new_n17911_), .A3(new_n16060_), .ZN(new_n17912_));
  AOI21_X1   g17720(.A1(new_n17904_), .A2(\asqrt[12] ), .B(new_n17912_), .ZN(new_n17913_));
  NOR2_X1    g17721(.A1(new_n17903_), .A2(new_n17913_), .ZN(new_n17914_));
  NAND2_X1   g17722(.A1(new_n17904_), .A2(\asqrt[12] ), .ZN(new_n17915_));
  AOI21_X1   g17723(.A1(new_n17903_), .A2(new_n17915_), .B(new_n16060_), .ZN(new_n17916_));
  NOR2_X1    g17724(.A1(new_n17675_), .A2(new_n17674_), .ZN(new_n17917_));
  NOR4_X1    g17725(.A1(new_n17893_), .A2(\asqrt[13] ), .A3(new_n17917_), .A4(new_n17288_), .ZN(new_n17918_));
  AOI21_X1   g17726(.A1(new_n17673_), .A2(new_n17270_), .B(new_n16060_), .ZN(new_n17919_));
  NOR2_X1    g17727(.A1(new_n17918_), .A2(new_n17919_), .ZN(new_n17920_));
  NAND2_X1   g17728(.A1(new_n17920_), .A2(new_n15447_), .ZN(new_n17921_));
  OAI21_X1   g17729(.A1(new_n17916_), .A2(new_n17921_), .B(new_n17914_), .ZN(new_n17922_));
  AOI22_X1   g17730(.A1(new_n17902_), .A2(new_n17886_), .B1(\asqrt[12] ), .B2(new_n17904_), .ZN(new_n17923_));
  OAI22_X1   g17731(.A1(new_n17923_), .A2(new_n16060_), .B1(new_n17903_), .B2(new_n17913_), .ZN(new_n17924_));
  NOR2_X1    g17732(.A1(new_n17300_), .A2(new_n15447_), .ZN(new_n17925_));
  NAND2_X1   g17733(.A1(new_n17294_), .A2(new_n17296_), .ZN(new_n17926_));
  NAND4_X1   g17734(.A1(\asqrt[10] ), .A2(new_n15447_), .A3(new_n17926_), .A4(new_n17300_), .ZN(new_n17927_));
  XOR2_X1    g17735(.A1(new_n17927_), .A2(new_n17925_), .Z(new_n17928_));
  NAND2_X1   g17736(.A1(new_n17928_), .A2(new_n14871_), .ZN(new_n17929_));
  AOI21_X1   g17737(.A1(new_n17924_), .A2(\asqrt[14] ), .B(new_n17929_), .ZN(new_n17930_));
  OAI21_X1   g17738(.A1(new_n17916_), .A2(new_n17914_), .B(\asqrt[14] ), .ZN(new_n17931_));
  AOI21_X1   g17739(.A1(new_n17922_), .A2(new_n17931_), .B(new_n14871_), .ZN(new_n17932_));
  NAND2_X1   g17740(.A1(new_n17307_), .A2(\asqrt[15] ), .ZN(new_n17933_));
  NOR2_X1    g17741(.A1(new_n17302_), .A2(new_n17303_), .ZN(new_n17934_));
  NOR4_X1    g17742(.A1(new_n17893_), .A2(\asqrt[15] ), .A3(new_n17934_), .A4(new_n17307_), .ZN(new_n17935_));
  XOR2_X1    g17743(.A1(new_n17935_), .A2(new_n17933_), .Z(new_n17936_));
  NAND2_X1   g17744(.A1(new_n17936_), .A2(new_n14273_), .ZN(new_n17937_));
  NOR2_X1    g17745(.A1(new_n17932_), .A2(new_n17937_), .ZN(new_n17938_));
  NOR3_X1    g17746(.A1(new_n17938_), .A2(new_n17922_), .A3(new_n17930_), .ZN(new_n17939_));
  INV_X1     g17747(.I(new_n17929_), .ZN(new_n17940_));
  AOI21_X1   g17748(.A1(new_n17931_), .A2(new_n17940_), .B(new_n17922_), .ZN(new_n17941_));
  OAI21_X1   g17749(.A1(new_n17941_), .A2(new_n17932_), .B(\asqrt[16] ), .ZN(new_n17942_));
  NOR4_X1    g17750(.A1(new_n17893_), .A2(\asqrt[16] ), .A3(new_n17310_), .A4(new_n17692_), .ZN(new_n17943_));
  AOI21_X1   g17751(.A1(new_n17933_), .A2(new_n17306_), .B(new_n14273_), .ZN(new_n17944_));
  NOR2_X1    g17752(.A1(new_n17943_), .A2(new_n17944_), .ZN(new_n17945_));
  NAND2_X1   g17753(.A1(new_n17945_), .A2(new_n13760_), .ZN(new_n17946_));
  INV_X1     g17754(.I(new_n17946_), .ZN(new_n17947_));
  NAND2_X1   g17755(.A1(new_n17942_), .A2(new_n17947_), .ZN(new_n17948_));
  NAND2_X1   g17756(.A1(new_n17948_), .A2(new_n17939_), .ZN(new_n17949_));
  OAI21_X1   g17757(.A1(new_n17932_), .A2(new_n17937_), .B(new_n17941_), .ZN(new_n17950_));
  NAND2_X1   g17758(.A1(new_n17950_), .A2(new_n17942_), .ZN(new_n17951_));
  NAND2_X1   g17759(.A1(new_n17322_), .A2(\asqrt[17] ), .ZN(new_n17952_));
  NOR4_X1    g17760(.A1(new_n17893_), .A2(\asqrt[17] ), .A3(new_n17317_), .A4(new_n17322_), .ZN(new_n17953_));
  XOR2_X1    g17761(.A1(new_n17953_), .A2(new_n17952_), .Z(new_n17954_));
  NAND2_X1   g17762(.A1(new_n17954_), .A2(new_n13192_), .ZN(new_n17955_));
  AOI21_X1   g17763(.A1(new_n17951_), .A2(\asqrt[17] ), .B(new_n17955_), .ZN(new_n17956_));
  NOR2_X1    g17764(.A1(new_n17956_), .A2(new_n17949_), .ZN(new_n17957_));
  AOI21_X1   g17765(.A1(new_n17942_), .A2(new_n17947_), .B(new_n17950_), .ZN(new_n17958_));
  AOI21_X1   g17766(.A1(new_n17950_), .A2(new_n17942_), .B(new_n13760_), .ZN(new_n17959_));
  OAI21_X1   g17767(.A1(new_n17958_), .A2(new_n17959_), .B(\asqrt[18] ), .ZN(new_n17960_));
  NOR4_X1    g17768(.A1(new_n17893_), .A2(\asqrt[18] ), .A3(new_n17324_), .A4(new_n17699_), .ZN(new_n17961_));
  AOI21_X1   g17769(.A1(new_n17952_), .A2(new_n17321_), .B(new_n13192_), .ZN(new_n17962_));
  NOR2_X1    g17770(.A1(new_n17961_), .A2(new_n17962_), .ZN(new_n17963_));
  NAND2_X1   g17771(.A1(new_n17963_), .A2(new_n12657_), .ZN(new_n17964_));
  INV_X1     g17772(.I(new_n17964_), .ZN(new_n17965_));
  NAND2_X1   g17773(.A1(new_n17960_), .A2(new_n17965_), .ZN(new_n17966_));
  NAND2_X1   g17774(.A1(new_n17966_), .A2(new_n17957_), .ZN(new_n17967_));
  AOI22_X1   g17775(.A1(new_n17951_), .A2(\asqrt[17] ), .B1(new_n17948_), .B2(new_n17939_), .ZN(new_n17968_));
  OAI22_X1   g17776(.A1(new_n17968_), .A2(new_n13192_), .B1(new_n17956_), .B2(new_n17949_), .ZN(new_n17969_));
  NAND2_X1   g17777(.A1(new_n17335_), .A2(\asqrt[19] ), .ZN(new_n17970_));
  NOR4_X1    g17778(.A1(new_n17893_), .A2(\asqrt[19] ), .A3(new_n17330_), .A4(new_n17335_), .ZN(new_n17971_));
  XOR2_X1    g17779(.A1(new_n17971_), .A2(new_n17970_), .Z(new_n17972_));
  NAND2_X1   g17780(.A1(new_n17972_), .A2(new_n12101_), .ZN(new_n17973_));
  AOI21_X1   g17781(.A1(new_n17969_), .A2(\asqrt[19] ), .B(new_n17973_), .ZN(new_n17974_));
  NOR2_X1    g17782(.A1(new_n17974_), .A2(new_n17967_), .ZN(new_n17975_));
  AOI22_X1   g17783(.A1(new_n17969_), .A2(\asqrt[19] ), .B1(new_n17966_), .B2(new_n17957_), .ZN(new_n17976_));
  NOR4_X1    g17784(.A1(new_n17893_), .A2(\asqrt[20] ), .A3(new_n17337_), .A4(new_n17706_), .ZN(new_n17977_));
  AOI21_X1   g17785(.A1(new_n17970_), .A2(new_n17334_), .B(new_n12101_), .ZN(new_n17978_));
  NOR2_X1    g17786(.A1(new_n17977_), .A2(new_n17978_), .ZN(new_n17979_));
  NAND2_X1   g17787(.A1(new_n17979_), .A2(new_n11631_), .ZN(new_n17980_));
  INV_X1     g17788(.I(new_n17980_), .ZN(new_n17981_));
  OAI21_X1   g17789(.A1(new_n17976_), .A2(new_n12101_), .B(new_n17981_), .ZN(new_n17982_));
  NAND2_X1   g17790(.A1(new_n17982_), .A2(new_n17975_), .ZN(new_n17983_));
  OAI22_X1   g17791(.A1(new_n17976_), .A2(new_n12101_), .B1(new_n17974_), .B2(new_n17967_), .ZN(new_n17984_));
  NAND2_X1   g17792(.A1(new_n17348_), .A2(\asqrt[21] ), .ZN(new_n17985_));
  NOR4_X1    g17793(.A1(new_n17893_), .A2(\asqrt[21] ), .A3(new_n17343_), .A4(new_n17348_), .ZN(new_n17986_));
  XOR2_X1    g17794(.A1(new_n17986_), .A2(new_n17985_), .Z(new_n17987_));
  NAND2_X1   g17795(.A1(new_n17987_), .A2(new_n11105_), .ZN(new_n17988_));
  AOI21_X1   g17796(.A1(new_n17984_), .A2(\asqrt[21] ), .B(new_n17988_), .ZN(new_n17989_));
  NOR2_X1    g17797(.A1(new_n17989_), .A2(new_n17983_), .ZN(new_n17990_));
  AOI22_X1   g17798(.A1(new_n17984_), .A2(\asqrt[21] ), .B1(new_n17982_), .B2(new_n17975_), .ZN(new_n17991_));
  NAND2_X1   g17799(.A1(new_n17713_), .A2(\asqrt[22] ), .ZN(new_n17992_));
  NOR4_X1    g17800(.A1(new_n17893_), .A2(\asqrt[22] ), .A3(new_n17351_), .A4(new_n17713_), .ZN(new_n17993_));
  XOR2_X1    g17801(.A1(new_n17993_), .A2(new_n17992_), .Z(new_n17994_));
  NAND2_X1   g17802(.A1(new_n17994_), .A2(new_n10614_), .ZN(new_n17995_));
  INV_X1     g17803(.I(new_n17995_), .ZN(new_n17996_));
  OAI21_X1   g17804(.A1(new_n17991_), .A2(new_n11105_), .B(new_n17996_), .ZN(new_n17997_));
  NAND2_X1   g17805(.A1(new_n17997_), .A2(new_n17990_), .ZN(new_n17998_));
  OAI22_X1   g17806(.A1(new_n17991_), .A2(new_n11105_), .B1(new_n17989_), .B2(new_n17983_), .ZN(new_n17999_));
  NOR4_X1    g17807(.A1(new_n17893_), .A2(\asqrt[23] ), .A3(new_n17358_), .A4(new_n17363_), .ZN(new_n18000_));
  AOI21_X1   g17808(.A1(new_n17992_), .A2(new_n17712_), .B(new_n10614_), .ZN(new_n18001_));
  NOR2_X1    g17809(.A1(new_n18000_), .A2(new_n18001_), .ZN(new_n18002_));
  NAND2_X1   g17810(.A1(new_n18002_), .A2(new_n10104_), .ZN(new_n18003_));
  AOI21_X1   g17811(.A1(new_n17999_), .A2(\asqrt[23] ), .B(new_n18003_), .ZN(new_n18004_));
  NOR2_X1    g17812(.A1(new_n18004_), .A2(new_n17998_), .ZN(new_n18005_));
  AOI22_X1   g17813(.A1(new_n17999_), .A2(\asqrt[23] ), .B1(new_n17997_), .B2(new_n17990_), .ZN(new_n18006_));
  NAND2_X1   g17814(.A1(new_n17720_), .A2(\asqrt[24] ), .ZN(new_n18007_));
  NOR4_X1    g17815(.A1(new_n17893_), .A2(\asqrt[24] ), .A3(new_n17366_), .A4(new_n17720_), .ZN(new_n18008_));
  XOR2_X1    g17816(.A1(new_n18008_), .A2(new_n18007_), .Z(new_n18009_));
  NAND2_X1   g17817(.A1(new_n18009_), .A2(new_n9672_), .ZN(new_n18010_));
  INV_X1     g17818(.I(new_n18010_), .ZN(new_n18011_));
  OAI21_X1   g17819(.A1(new_n18006_), .A2(new_n10104_), .B(new_n18011_), .ZN(new_n18012_));
  NAND2_X1   g17820(.A1(new_n18012_), .A2(new_n18005_), .ZN(new_n18013_));
  OAI22_X1   g17821(.A1(new_n18006_), .A2(new_n10104_), .B1(new_n18004_), .B2(new_n17998_), .ZN(new_n18014_));
  NOR4_X1    g17822(.A1(new_n17893_), .A2(\asqrt[25] ), .A3(new_n17373_), .A4(new_n17378_), .ZN(new_n18015_));
  AOI21_X1   g17823(.A1(new_n18007_), .A2(new_n17719_), .B(new_n9672_), .ZN(new_n18016_));
  NOR2_X1    g17824(.A1(new_n18015_), .A2(new_n18016_), .ZN(new_n18017_));
  NAND2_X1   g17825(.A1(new_n18017_), .A2(new_n9212_), .ZN(new_n18018_));
  AOI21_X1   g17826(.A1(new_n18014_), .A2(\asqrt[25] ), .B(new_n18018_), .ZN(new_n18019_));
  NOR2_X1    g17827(.A1(new_n18019_), .A2(new_n18013_), .ZN(new_n18020_));
  AOI22_X1   g17828(.A1(new_n18014_), .A2(\asqrt[25] ), .B1(new_n18012_), .B2(new_n18005_), .ZN(new_n18021_));
  NAND2_X1   g17829(.A1(new_n17727_), .A2(\asqrt[26] ), .ZN(new_n18022_));
  NOR4_X1    g17830(.A1(new_n17893_), .A2(\asqrt[26] ), .A3(new_n17381_), .A4(new_n17727_), .ZN(new_n18023_));
  XOR2_X1    g17831(.A1(new_n18023_), .A2(new_n18022_), .Z(new_n18024_));
  NAND2_X1   g17832(.A1(new_n18024_), .A2(new_n8763_), .ZN(new_n18025_));
  INV_X1     g17833(.I(new_n18025_), .ZN(new_n18026_));
  OAI21_X1   g17834(.A1(new_n18021_), .A2(new_n9212_), .B(new_n18026_), .ZN(new_n18027_));
  NAND2_X1   g17835(.A1(new_n18027_), .A2(new_n18020_), .ZN(new_n18028_));
  OAI22_X1   g17836(.A1(new_n18021_), .A2(new_n9212_), .B1(new_n18019_), .B2(new_n18013_), .ZN(new_n18029_));
  NOR4_X1    g17837(.A1(new_n17893_), .A2(\asqrt[27] ), .A3(new_n17388_), .A4(new_n17393_), .ZN(new_n18030_));
  AOI21_X1   g17838(.A1(new_n18022_), .A2(new_n17726_), .B(new_n8763_), .ZN(new_n18031_));
  NOR2_X1    g17839(.A1(new_n18030_), .A2(new_n18031_), .ZN(new_n18032_));
  NAND2_X1   g17840(.A1(new_n18032_), .A2(new_n8319_), .ZN(new_n18033_));
  AOI21_X1   g17841(.A1(new_n18029_), .A2(\asqrt[27] ), .B(new_n18033_), .ZN(new_n18034_));
  NOR2_X1    g17842(.A1(new_n18034_), .A2(new_n18028_), .ZN(new_n18035_));
  AOI22_X1   g17843(.A1(new_n18029_), .A2(\asqrt[27] ), .B1(new_n18027_), .B2(new_n18020_), .ZN(new_n18036_));
  NAND2_X1   g17844(.A1(new_n17734_), .A2(\asqrt[28] ), .ZN(new_n18037_));
  NOR4_X1    g17845(.A1(new_n17893_), .A2(\asqrt[28] ), .A3(new_n17396_), .A4(new_n17734_), .ZN(new_n18038_));
  XOR2_X1    g17846(.A1(new_n18038_), .A2(new_n18037_), .Z(new_n18039_));
  NAND2_X1   g17847(.A1(new_n18039_), .A2(new_n7931_), .ZN(new_n18040_));
  INV_X1     g17848(.I(new_n18040_), .ZN(new_n18041_));
  OAI21_X1   g17849(.A1(new_n18036_), .A2(new_n8319_), .B(new_n18041_), .ZN(new_n18042_));
  NAND2_X1   g17850(.A1(new_n18042_), .A2(new_n18035_), .ZN(new_n18043_));
  OAI22_X1   g17851(.A1(new_n18036_), .A2(new_n8319_), .B1(new_n18034_), .B2(new_n18028_), .ZN(new_n18044_));
  NOR4_X1    g17852(.A1(new_n17893_), .A2(\asqrt[29] ), .A3(new_n17403_), .A4(new_n17408_), .ZN(new_n18045_));
  AOI21_X1   g17853(.A1(new_n18037_), .A2(new_n17733_), .B(new_n7931_), .ZN(new_n18046_));
  NOR2_X1    g17854(.A1(new_n18045_), .A2(new_n18046_), .ZN(new_n18047_));
  NAND2_X1   g17855(.A1(new_n18047_), .A2(new_n7517_), .ZN(new_n18048_));
  AOI21_X1   g17856(.A1(new_n18044_), .A2(\asqrt[29] ), .B(new_n18048_), .ZN(new_n18049_));
  NOR2_X1    g17857(.A1(new_n18049_), .A2(new_n18043_), .ZN(new_n18050_));
  AOI22_X1   g17858(.A1(new_n18044_), .A2(\asqrt[29] ), .B1(new_n18042_), .B2(new_n18035_), .ZN(new_n18051_));
  NAND2_X1   g17859(.A1(new_n17741_), .A2(\asqrt[30] ), .ZN(new_n18052_));
  NOR4_X1    g17860(.A1(new_n17893_), .A2(\asqrt[30] ), .A3(new_n17411_), .A4(new_n17741_), .ZN(new_n18053_));
  XOR2_X1    g17861(.A1(new_n18053_), .A2(new_n18052_), .Z(new_n18054_));
  NAND2_X1   g17862(.A1(new_n18054_), .A2(new_n7110_), .ZN(new_n18055_));
  INV_X1     g17863(.I(new_n18055_), .ZN(new_n18056_));
  OAI21_X1   g17864(.A1(new_n18051_), .A2(new_n7517_), .B(new_n18056_), .ZN(new_n18057_));
  NAND2_X1   g17865(.A1(new_n18057_), .A2(new_n18050_), .ZN(new_n18058_));
  OAI22_X1   g17866(.A1(new_n18051_), .A2(new_n7517_), .B1(new_n18049_), .B2(new_n18043_), .ZN(new_n18059_));
  NAND2_X1   g17867(.A1(new_n17423_), .A2(\asqrt[31] ), .ZN(new_n18060_));
  NOR4_X1    g17868(.A1(new_n17893_), .A2(\asqrt[31] ), .A3(new_n17418_), .A4(new_n17423_), .ZN(new_n18061_));
  XOR2_X1    g17869(.A1(new_n18061_), .A2(new_n18060_), .Z(new_n18062_));
  NAND2_X1   g17870(.A1(new_n18062_), .A2(new_n6708_), .ZN(new_n18063_));
  AOI21_X1   g17871(.A1(new_n18059_), .A2(\asqrt[31] ), .B(new_n18063_), .ZN(new_n18064_));
  NOR2_X1    g17872(.A1(new_n18064_), .A2(new_n18058_), .ZN(new_n18065_));
  AOI22_X1   g17873(.A1(new_n18059_), .A2(\asqrt[31] ), .B1(new_n18057_), .B2(new_n18050_), .ZN(new_n18066_));
  NOR4_X1    g17874(.A1(new_n17893_), .A2(\asqrt[32] ), .A3(new_n17426_), .A4(new_n17748_), .ZN(new_n18067_));
  AOI21_X1   g17875(.A1(new_n18060_), .A2(new_n17422_), .B(new_n6708_), .ZN(new_n18068_));
  NOR2_X1    g17876(.A1(new_n18067_), .A2(new_n18068_), .ZN(new_n18069_));
  NAND2_X1   g17877(.A1(new_n18069_), .A2(new_n6365_), .ZN(new_n18070_));
  INV_X1     g17878(.I(new_n18070_), .ZN(new_n18071_));
  OAI21_X1   g17879(.A1(new_n18066_), .A2(new_n6708_), .B(new_n18071_), .ZN(new_n18072_));
  NAND2_X1   g17880(.A1(new_n18072_), .A2(new_n18065_), .ZN(new_n18073_));
  OAI22_X1   g17881(.A1(new_n18066_), .A2(new_n6708_), .B1(new_n18064_), .B2(new_n18058_), .ZN(new_n18074_));
  NAND2_X1   g17882(.A1(new_n17438_), .A2(\asqrt[33] ), .ZN(new_n18075_));
  NOR4_X1    g17883(.A1(new_n17893_), .A2(\asqrt[33] ), .A3(new_n17433_), .A4(new_n17438_), .ZN(new_n18076_));
  XOR2_X1    g17884(.A1(new_n18076_), .A2(new_n18075_), .Z(new_n18077_));
  NAND2_X1   g17885(.A1(new_n18077_), .A2(new_n5991_), .ZN(new_n18078_));
  AOI21_X1   g17886(.A1(new_n18074_), .A2(\asqrt[33] ), .B(new_n18078_), .ZN(new_n18079_));
  NOR2_X1    g17887(.A1(new_n18079_), .A2(new_n18073_), .ZN(new_n18080_));
  AOI22_X1   g17888(.A1(new_n18074_), .A2(\asqrt[33] ), .B1(new_n18072_), .B2(new_n18065_), .ZN(new_n18081_));
  NOR4_X1    g17889(.A1(new_n17893_), .A2(\asqrt[34] ), .A3(new_n17441_), .A4(new_n17755_), .ZN(new_n18082_));
  AOI21_X1   g17890(.A1(new_n18075_), .A2(new_n17437_), .B(new_n5991_), .ZN(new_n18083_));
  NOR2_X1    g17891(.A1(new_n18082_), .A2(new_n18083_), .ZN(new_n18084_));
  NAND2_X1   g17892(.A1(new_n18084_), .A2(new_n5626_), .ZN(new_n18085_));
  INV_X1     g17893(.I(new_n18085_), .ZN(new_n18086_));
  OAI21_X1   g17894(.A1(new_n18081_), .A2(new_n5991_), .B(new_n18086_), .ZN(new_n18087_));
  NAND2_X1   g17895(.A1(new_n18087_), .A2(new_n18080_), .ZN(new_n18088_));
  OAI22_X1   g17896(.A1(new_n18081_), .A2(new_n5991_), .B1(new_n18079_), .B2(new_n18073_), .ZN(new_n18089_));
  NAND2_X1   g17897(.A1(new_n17453_), .A2(\asqrt[35] ), .ZN(new_n18090_));
  NOR4_X1    g17898(.A1(new_n17893_), .A2(\asqrt[35] ), .A3(new_n17448_), .A4(new_n17453_), .ZN(new_n18091_));
  XOR2_X1    g17899(.A1(new_n18091_), .A2(new_n18090_), .Z(new_n18092_));
  NAND2_X1   g17900(.A1(new_n18092_), .A2(new_n5273_), .ZN(new_n18093_));
  AOI21_X1   g17901(.A1(new_n18089_), .A2(\asqrt[35] ), .B(new_n18093_), .ZN(new_n18094_));
  NOR2_X1    g17902(.A1(new_n18094_), .A2(new_n18088_), .ZN(new_n18095_));
  AOI22_X1   g17903(.A1(new_n18089_), .A2(\asqrt[35] ), .B1(new_n18087_), .B2(new_n18080_), .ZN(new_n18096_));
  NAND2_X1   g17904(.A1(new_n17762_), .A2(\asqrt[36] ), .ZN(new_n18097_));
  NOR4_X1    g17905(.A1(new_n17893_), .A2(\asqrt[36] ), .A3(new_n17456_), .A4(new_n17762_), .ZN(new_n18098_));
  XOR2_X1    g17906(.A1(new_n18098_), .A2(new_n18097_), .Z(new_n18099_));
  NAND2_X1   g17907(.A1(new_n18099_), .A2(new_n4973_), .ZN(new_n18100_));
  INV_X1     g17908(.I(new_n18100_), .ZN(new_n18101_));
  OAI21_X1   g17909(.A1(new_n18096_), .A2(new_n5273_), .B(new_n18101_), .ZN(new_n18102_));
  NAND2_X1   g17910(.A1(new_n18102_), .A2(new_n18095_), .ZN(new_n18103_));
  OAI22_X1   g17911(.A1(new_n18096_), .A2(new_n5273_), .B1(new_n18094_), .B2(new_n18088_), .ZN(new_n18104_));
  NOR4_X1    g17912(.A1(new_n17893_), .A2(\asqrt[37] ), .A3(new_n17463_), .A4(new_n17468_), .ZN(new_n18105_));
  AOI21_X1   g17913(.A1(new_n18097_), .A2(new_n17761_), .B(new_n4973_), .ZN(new_n18106_));
  NOR2_X1    g17914(.A1(new_n18105_), .A2(new_n18106_), .ZN(new_n18107_));
  NAND2_X1   g17915(.A1(new_n18107_), .A2(new_n4645_), .ZN(new_n18108_));
  AOI21_X1   g17916(.A1(new_n18104_), .A2(\asqrt[37] ), .B(new_n18108_), .ZN(new_n18109_));
  NOR2_X1    g17917(.A1(new_n18109_), .A2(new_n18103_), .ZN(new_n18110_));
  AOI22_X1   g17918(.A1(new_n18104_), .A2(\asqrt[37] ), .B1(new_n18102_), .B2(new_n18095_), .ZN(new_n18111_));
  NAND2_X1   g17919(.A1(new_n17769_), .A2(\asqrt[38] ), .ZN(new_n18112_));
  NOR4_X1    g17920(.A1(new_n17893_), .A2(\asqrt[38] ), .A3(new_n17471_), .A4(new_n17769_), .ZN(new_n18113_));
  XOR2_X1    g17921(.A1(new_n18113_), .A2(new_n18112_), .Z(new_n18114_));
  NAND2_X1   g17922(.A1(new_n18114_), .A2(new_n4330_), .ZN(new_n18115_));
  INV_X1     g17923(.I(new_n18115_), .ZN(new_n18116_));
  OAI21_X1   g17924(.A1(new_n18111_), .A2(new_n4645_), .B(new_n18116_), .ZN(new_n18117_));
  NAND2_X1   g17925(.A1(new_n18117_), .A2(new_n18110_), .ZN(new_n18118_));
  OAI22_X1   g17926(.A1(new_n18111_), .A2(new_n4645_), .B1(new_n18109_), .B2(new_n18103_), .ZN(new_n18119_));
  NOR4_X1    g17927(.A1(new_n17893_), .A2(\asqrt[39] ), .A3(new_n17478_), .A4(new_n17483_), .ZN(new_n18120_));
  AOI21_X1   g17928(.A1(new_n18112_), .A2(new_n17768_), .B(new_n4330_), .ZN(new_n18121_));
  NOR2_X1    g17929(.A1(new_n18120_), .A2(new_n18121_), .ZN(new_n18122_));
  NAND2_X1   g17930(.A1(new_n18122_), .A2(new_n4018_), .ZN(new_n18123_));
  AOI21_X1   g17931(.A1(new_n18119_), .A2(\asqrt[39] ), .B(new_n18123_), .ZN(new_n18124_));
  NOR2_X1    g17932(.A1(new_n18124_), .A2(new_n18118_), .ZN(new_n18125_));
  AOI22_X1   g17933(.A1(new_n18119_), .A2(\asqrt[39] ), .B1(new_n18117_), .B2(new_n18110_), .ZN(new_n18126_));
  NAND2_X1   g17934(.A1(new_n17776_), .A2(\asqrt[40] ), .ZN(new_n18127_));
  NOR4_X1    g17935(.A1(new_n17893_), .A2(\asqrt[40] ), .A3(new_n17486_), .A4(new_n17776_), .ZN(new_n18128_));
  XOR2_X1    g17936(.A1(new_n18128_), .A2(new_n18127_), .Z(new_n18129_));
  NAND2_X1   g17937(.A1(new_n18129_), .A2(new_n3760_), .ZN(new_n18130_));
  INV_X1     g17938(.I(new_n18130_), .ZN(new_n18131_));
  OAI21_X1   g17939(.A1(new_n18126_), .A2(new_n4018_), .B(new_n18131_), .ZN(new_n18132_));
  NAND2_X1   g17940(.A1(new_n18132_), .A2(new_n18125_), .ZN(new_n18133_));
  OAI22_X1   g17941(.A1(new_n18126_), .A2(new_n4018_), .B1(new_n18124_), .B2(new_n18118_), .ZN(new_n18134_));
  NOR4_X1    g17942(.A1(new_n17893_), .A2(\asqrt[41] ), .A3(new_n17493_), .A4(new_n17498_), .ZN(new_n18135_));
  AOI21_X1   g17943(.A1(new_n18127_), .A2(new_n17775_), .B(new_n3760_), .ZN(new_n18136_));
  NOR2_X1    g17944(.A1(new_n18135_), .A2(new_n18136_), .ZN(new_n18137_));
  NAND2_X1   g17945(.A1(new_n18137_), .A2(new_n3481_), .ZN(new_n18138_));
  AOI21_X1   g17946(.A1(new_n18134_), .A2(\asqrt[41] ), .B(new_n18138_), .ZN(new_n18139_));
  NOR2_X1    g17947(.A1(new_n18139_), .A2(new_n18133_), .ZN(new_n18140_));
  AOI22_X1   g17948(.A1(new_n18134_), .A2(\asqrt[41] ), .B1(new_n18132_), .B2(new_n18125_), .ZN(new_n18141_));
  NAND2_X1   g17949(.A1(new_n17783_), .A2(\asqrt[42] ), .ZN(new_n18142_));
  NOR4_X1    g17950(.A1(new_n17893_), .A2(\asqrt[42] ), .A3(new_n17501_), .A4(new_n17783_), .ZN(new_n18143_));
  XOR2_X1    g17951(.A1(new_n18143_), .A2(new_n18142_), .Z(new_n18144_));
  NAND2_X1   g17952(.A1(new_n18144_), .A2(new_n3208_), .ZN(new_n18145_));
  INV_X1     g17953(.I(new_n18145_), .ZN(new_n18146_));
  OAI21_X1   g17954(.A1(new_n18141_), .A2(new_n3481_), .B(new_n18146_), .ZN(new_n18147_));
  NAND2_X1   g17955(.A1(new_n18147_), .A2(new_n18140_), .ZN(new_n18148_));
  OAI22_X1   g17956(.A1(new_n18141_), .A2(new_n3481_), .B1(new_n18139_), .B2(new_n18133_), .ZN(new_n18149_));
  NAND2_X1   g17957(.A1(new_n17513_), .A2(\asqrt[43] ), .ZN(new_n18150_));
  NOR4_X1    g17958(.A1(new_n17893_), .A2(\asqrt[43] ), .A3(new_n17508_), .A4(new_n17513_), .ZN(new_n18151_));
  XOR2_X1    g17959(.A1(new_n18151_), .A2(new_n18150_), .Z(new_n18152_));
  NAND2_X1   g17960(.A1(new_n18152_), .A2(new_n2941_), .ZN(new_n18153_));
  AOI21_X1   g17961(.A1(new_n18149_), .A2(\asqrt[43] ), .B(new_n18153_), .ZN(new_n18154_));
  NOR2_X1    g17962(.A1(new_n18154_), .A2(new_n18148_), .ZN(new_n18155_));
  AOI22_X1   g17963(.A1(new_n18149_), .A2(\asqrt[43] ), .B1(new_n18147_), .B2(new_n18140_), .ZN(new_n18156_));
  NOR4_X1    g17964(.A1(new_n17893_), .A2(\asqrt[44] ), .A3(new_n17516_), .A4(new_n17790_), .ZN(new_n18157_));
  AOI21_X1   g17965(.A1(new_n18150_), .A2(new_n17512_), .B(new_n2941_), .ZN(new_n18158_));
  NOR2_X1    g17966(.A1(new_n18157_), .A2(new_n18158_), .ZN(new_n18159_));
  NAND2_X1   g17967(.A1(new_n18159_), .A2(new_n2728_), .ZN(new_n18160_));
  INV_X1     g17968(.I(new_n18160_), .ZN(new_n18161_));
  OAI21_X1   g17969(.A1(new_n18156_), .A2(new_n2941_), .B(new_n18161_), .ZN(new_n18162_));
  NAND2_X1   g17970(.A1(new_n18162_), .A2(new_n18155_), .ZN(new_n18163_));
  OAI22_X1   g17971(.A1(new_n18156_), .A2(new_n2941_), .B1(new_n18154_), .B2(new_n18148_), .ZN(new_n18164_));
  NAND2_X1   g17972(.A1(new_n17528_), .A2(\asqrt[45] ), .ZN(new_n18165_));
  NOR4_X1    g17973(.A1(new_n17893_), .A2(\asqrt[45] ), .A3(new_n17523_), .A4(new_n17528_), .ZN(new_n18166_));
  XOR2_X1    g17974(.A1(new_n18166_), .A2(new_n18165_), .Z(new_n18167_));
  NAND2_X1   g17975(.A1(new_n18167_), .A2(new_n2488_), .ZN(new_n18168_));
  AOI21_X1   g17976(.A1(new_n18164_), .A2(\asqrt[45] ), .B(new_n18168_), .ZN(new_n18169_));
  NOR2_X1    g17977(.A1(new_n18169_), .A2(new_n18163_), .ZN(new_n18170_));
  AOI22_X1   g17978(.A1(new_n18164_), .A2(\asqrt[45] ), .B1(new_n18162_), .B2(new_n18155_), .ZN(new_n18171_));
  NOR4_X1    g17979(.A1(new_n17893_), .A2(\asqrt[46] ), .A3(new_n17531_), .A4(new_n17797_), .ZN(new_n18172_));
  AOI21_X1   g17980(.A1(new_n18165_), .A2(new_n17527_), .B(new_n2488_), .ZN(new_n18173_));
  NOR2_X1    g17981(.A1(new_n18172_), .A2(new_n18173_), .ZN(new_n18174_));
  NAND2_X1   g17982(.A1(new_n18174_), .A2(new_n2253_), .ZN(new_n18175_));
  INV_X1     g17983(.I(new_n18175_), .ZN(new_n18176_));
  OAI21_X1   g17984(.A1(new_n18171_), .A2(new_n2488_), .B(new_n18176_), .ZN(new_n18177_));
  NAND2_X1   g17985(.A1(new_n18177_), .A2(new_n18170_), .ZN(new_n18178_));
  OAI22_X1   g17986(.A1(new_n18171_), .A2(new_n2488_), .B1(new_n18169_), .B2(new_n18163_), .ZN(new_n18179_));
  NAND2_X1   g17987(.A1(new_n17543_), .A2(\asqrt[47] ), .ZN(new_n18180_));
  NOR4_X1    g17988(.A1(new_n17893_), .A2(\asqrt[47] ), .A3(new_n17538_), .A4(new_n17543_), .ZN(new_n18181_));
  XOR2_X1    g17989(.A1(new_n18181_), .A2(new_n18180_), .Z(new_n18182_));
  NAND2_X1   g17990(.A1(new_n18182_), .A2(new_n2046_), .ZN(new_n18183_));
  AOI21_X1   g17991(.A1(new_n18179_), .A2(\asqrt[47] ), .B(new_n18183_), .ZN(new_n18184_));
  NOR2_X1    g17992(.A1(new_n18184_), .A2(new_n18178_), .ZN(new_n18185_));
  AOI22_X1   g17993(.A1(new_n18179_), .A2(\asqrt[47] ), .B1(new_n18177_), .B2(new_n18170_), .ZN(new_n18186_));
  NAND2_X1   g17994(.A1(new_n17804_), .A2(\asqrt[48] ), .ZN(new_n18187_));
  NOR4_X1    g17995(.A1(new_n17893_), .A2(\asqrt[48] ), .A3(new_n17546_), .A4(new_n17804_), .ZN(new_n18188_));
  XOR2_X1    g17996(.A1(new_n18188_), .A2(new_n18187_), .Z(new_n18189_));
  NAND2_X1   g17997(.A1(new_n18189_), .A2(new_n1854_), .ZN(new_n18190_));
  INV_X1     g17998(.I(new_n18190_), .ZN(new_n18191_));
  OAI21_X1   g17999(.A1(new_n18186_), .A2(new_n2046_), .B(new_n18191_), .ZN(new_n18192_));
  NAND2_X1   g18000(.A1(new_n18192_), .A2(new_n18185_), .ZN(new_n18193_));
  OAI22_X1   g18001(.A1(new_n18186_), .A2(new_n2046_), .B1(new_n18184_), .B2(new_n18178_), .ZN(new_n18194_));
  NOR4_X1    g18002(.A1(new_n17893_), .A2(\asqrt[49] ), .A3(new_n17553_), .A4(new_n17558_), .ZN(new_n18195_));
  AOI21_X1   g18003(.A1(new_n18187_), .A2(new_n17803_), .B(new_n1854_), .ZN(new_n18196_));
  NOR2_X1    g18004(.A1(new_n18195_), .A2(new_n18196_), .ZN(new_n18197_));
  NAND2_X1   g18005(.A1(new_n18197_), .A2(new_n1595_), .ZN(new_n18198_));
  AOI21_X1   g18006(.A1(new_n18194_), .A2(\asqrt[49] ), .B(new_n18198_), .ZN(new_n18199_));
  NOR2_X1    g18007(.A1(new_n18199_), .A2(new_n18193_), .ZN(new_n18200_));
  AOI22_X1   g18008(.A1(new_n18194_), .A2(\asqrt[49] ), .B1(new_n18192_), .B2(new_n18185_), .ZN(new_n18201_));
  NAND2_X1   g18009(.A1(new_n17811_), .A2(\asqrt[50] ), .ZN(new_n18202_));
  NOR4_X1    g18010(.A1(new_n17893_), .A2(\asqrt[50] ), .A3(new_n17561_), .A4(new_n17811_), .ZN(new_n18203_));
  XOR2_X1    g18011(.A1(new_n18203_), .A2(new_n18202_), .Z(new_n18204_));
  NAND2_X1   g18012(.A1(new_n18204_), .A2(new_n1436_), .ZN(new_n18205_));
  INV_X1     g18013(.I(new_n18205_), .ZN(new_n18206_));
  OAI21_X1   g18014(.A1(new_n18201_), .A2(new_n1595_), .B(new_n18206_), .ZN(new_n18207_));
  NAND2_X1   g18015(.A1(new_n18207_), .A2(new_n18200_), .ZN(new_n18208_));
  OAI22_X1   g18016(.A1(new_n18201_), .A2(new_n1595_), .B1(new_n18199_), .B2(new_n18193_), .ZN(new_n18209_));
  NOR4_X1    g18017(.A1(new_n17893_), .A2(\asqrt[51] ), .A3(new_n17568_), .A4(new_n17573_), .ZN(new_n18210_));
  AOI21_X1   g18018(.A1(new_n18202_), .A2(new_n17810_), .B(new_n1436_), .ZN(new_n18211_));
  NOR2_X1    g18019(.A1(new_n18210_), .A2(new_n18211_), .ZN(new_n18212_));
  NAND2_X1   g18020(.A1(new_n18212_), .A2(new_n1260_), .ZN(new_n18213_));
  AOI21_X1   g18021(.A1(new_n18209_), .A2(\asqrt[51] ), .B(new_n18213_), .ZN(new_n18214_));
  NOR2_X1    g18022(.A1(new_n18214_), .A2(new_n18208_), .ZN(new_n18215_));
  AOI22_X1   g18023(.A1(new_n18209_), .A2(\asqrt[51] ), .B1(new_n18207_), .B2(new_n18200_), .ZN(new_n18216_));
  NAND2_X1   g18024(.A1(new_n17818_), .A2(\asqrt[52] ), .ZN(new_n18217_));
  NOR4_X1    g18025(.A1(new_n17893_), .A2(\asqrt[52] ), .A3(new_n17576_), .A4(new_n17818_), .ZN(new_n18218_));
  XOR2_X1    g18026(.A1(new_n18218_), .A2(new_n18217_), .Z(new_n18219_));
  NAND2_X1   g18027(.A1(new_n18219_), .A2(new_n1096_), .ZN(new_n18220_));
  INV_X1     g18028(.I(new_n18220_), .ZN(new_n18221_));
  OAI21_X1   g18029(.A1(new_n18216_), .A2(new_n1260_), .B(new_n18221_), .ZN(new_n18222_));
  NAND2_X1   g18030(.A1(new_n18222_), .A2(new_n18215_), .ZN(new_n18223_));
  OAI22_X1   g18031(.A1(new_n18216_), .A2(new_n1260_), .B1(new_n18214_), .B2(new_n18208_), .ZN(new_n18224_));
  NOR4_X1    g18032(.A1(new_n17893_), .A2(\asqrt[53] ), .A3(new_n17583_), .A4(new_n17588_), .ZN(new_n18225_));
  AOI21_X1   g18033(.A1(new_n18217_), .A2(new_n17817_), .B(new_n1096_), .ZN(new_n18226_));
  NOR2_X1    g18034(.A1(new_n18225_), .A2(new_n18226_), .ZN(new_n18227_));
  NAND2_X1   g18035(.A1(new_n18227_), .A2(new_n970_), .ZN(new_n18228_));
  AOI21_X1   g18036(.A1(new_n18224_), .A2(\asqrt[53] ), .B(new_n18228_), .ZN(new_n18229_));
  NOR2_X1    g18037(.A1(new_n18229_), .A2(new_n18223_), .ZN(new_n18230_));
  AOI22_X1   g18038(.A1(new_n18224_), .A2(\asqrt[53] ), .B1(new_n18222_), .B2(new_n18215_), .ZN(new_n18231_));
  NAND2_X1   g18039(.A1(new_n17825_), .A2(\asqrt[54] ), .ZN(new_n18232_));
  NOR4_X1    g18040(.A1(new_n17893_), .A2(\asqrt[54] ), .A3(new_n17590_), .A4(new_n17825_), .ZN(new_n18233_));
  XOR2_X1    g18041(.A1(new_n18233_), .A2(new_n18232_), .Z(new_n18234_));
  NAND2_X1   g18042(.A1(new_n18234_), .A2(new_n825_), .ZN(new_n18235_));
  INV_X1     g18043(.I(new_n18235_), .ZN(new_n18236_));
  OAI21_X1   g18044(.A1(new_n18231_), .A2(new_n970_), .B(new_n18236_), .ZN(new_n18237_));
  NAND2_X1   g18045(.A1(new_n18237_), .A2(new_n18230_), .ZN(new_n18238_));
  OAI22_X1   g18046(.A1(new_n18231_), .A2(new_n970_), .B1(new_n18229_), .B2(new_n18223_), .ZN(new_n18239_));
  NAND2_X1   g18047(.A1(new_n17601_), .A2(\asqrt[55] ), .ZN(new_n18240_));
  NOR4_X1    g18048(.A1(new_n17893_), .A2(\asqrt[55] ), .A3(new_n17596_), .A4(new_n17601_), .ZN(new_n18241_));
  XOR2_X1    g18049(.A1(new_n18241_), .A2(new_n18240_), .Z(new_n18242_));
  NAND2_X1   g18050(.A1(new_n18242_), .A2(new_n724_), .ZN(new_n18243_));
  AOI21_X1   g18051(.A1(new_n18239_), .A2(\asqrt[55] ), .B(new_n18243_), .ZN(new_n18244_));
  NOR2_X1    g18052(.A1(new_n18244_), .A2(new_n18238_), .ZN(new_n18245_));
  AOI22_X1   g18053(.A1(new_n18239_), .A2(\asqrt[55] ), .B1(new_n18237_), .B2(new_n18230_), .ZN(new_n18246_));
  NOR4_X1    g18054(.A1(new_n17893_), .A2(\asqrt[56] ), .A3(new_n17603_), .A4(new_n17832_), .ZN(new_n18247_));
  AOI21_X1   g18055(.A1(new_n18240_), .A2(new_n17600_), .B(new_n724_), .ZN(new_n18248_));
  NOR2_X1    g18056(.A1(new_n18247_), .A2(new_n18248_), .ZN(new_n18249_));
  NAND2_X1   g18057(.A1(new_n18249_), .A2(new_n587_), .ZN(new_n18250_));
  INV_X1     g18058(.I(new_n18250_), .ZN(new_n18251_));
  OAI21_X1   g18059(.A1(new_n18246_), .A2(new_n724_), .B(new_n18251_), .ZN(new_n18252_));
  NAND2_X1   g18060(.A1(new_n18252_), .A2(new_n18245_), .ZN(new_n18253_));
  NAND2_X1   g18061(.A1(new_n18224_), .A2(\asqrt[53] ), .ZN(new_n18254_));
  AOI21_X1   g18062(.A1(new_n18254_), .A2(new_n18223_), .B(new_n970_), .ZN(new_n18255_));
  OAI21_X1   g18063(.A1(new_n18230_), .A2(new_n18255_), .B(\asqrt[55] ), .ZN(new_n18256_));
  AOI21_X1   g18064(.A1(new_n18238_), .A2(new_n18256_), .B(new_n724_), .ZN(new_n18257_));
  OAI21_X1   g18065(.A1(new_n18245_), .A2(new_n18257_), .B(\asqrt[57] ), .ZN(new_n18258_));
  NOR4_X1    g18066(.A1(new_n17893_), .A2(\asqrt[57] ), .A3(new_n17609_), .A4(new_n17614_), .ZN(new_n18259_));
  XOR2_X1    g18067(.A1(new_n18259_), .A2(new_n17633_), .Z(new_n18260_));
  NAND2_X1   g18068(.A1(new_n18260_), .A2(new_n504_), .ZN(new_n18261_));
  INV_X1     g18069(.I(new_n18261_), .ZN(new_n18262_));
  AOI21_X1   g18070(.A1(new_n18258_), .A2(new_n18262_), .B(new_n18253_), .ZN(new_n18263_));
  OAI22_X1   g18071(.A1(new_n18246_), .A2(new_n724_), .B1(new_n18244_), .B2(new_n18238_), .ZN(new_n18264_));
  AOI22_X1   g18072(.A1(new_n18264_), .A2(\asqrt[57] ), .B1(new_n18252_), .B2(new_n18245_), .ZN(new_n18265_));
  NOR4_X1    g18073(.A1(new_n17893_), .A2(\asqrt[58] ), .A3(new_n17616_), .A4(new_n17839_), .ZN(new_n18266_));
  XOR2_X1    g18074(.A1(new_n18266_), .A2(new_n17859_), .Z(new_n18267_));
  NAND2_X1   g18075(.A1(new_n18267_), .A2(new_n376_), .ZN(new_n18268_));
  INV_X1     g18076(.I(new_n18268_), .ZN(new_n18269_));
  OAI21_X1   g18077(.A1(new_n18265_), .A2(new_n504_), .B(new_n18269_), .ZN(new_n18270_));
  NAND2_X1   g18078(.A1(new_n18270_), .A2(new_n18263_), .ZN(new_n18271_));
  AOI21_X1   g18079(.A1(new_n18253_), .A2(new_n18258_), .B(new_n504_), .ZN(new_n18272_));
  OAI21_X1   g18080(.A1(new_n18263_), .A2(new_n18272_), .B(\asqrt[59] ), .ZN(new_n18273_));
  NOR4_X1    g18081(.A1(new_n17893_), .A2(\asqrt[59] ), .A3(new_n17622_), .A4(new_n17627_), .ZN(new_n18274_));
  XOR2_X1    g18082(.A1(new_n18274_), .A2(new_n17635_), .Z(new_n18275_));
  AND2_X2    g18083(.A1(new_n18275_), .A2(new_n275_), .Z(new_n18276_));
  AOI21_X1   g18084(.A1(new_n18273_), .A2(new_n18276_), .B(new_n18271_), .ZN(new_n18277_));
  INV_X1     g18085(.I(new_n17921_), .ZN(new_n18278_));
  OAI21_X1   g18086(.A1(new_n17923_), .A2(new_n16060_), .B(new_n18278_), .ZN(new_n18279_));
  AOI22_X1   g18087(.A1(new_n17924_), .A2(\asqrt[14] ), .B1(new_n18279_), .B2(new_n17914_), .ZN(new_n18280_));
  INV_X1     g18088(.I(new_n17937_), .ZN(new_n18281_));
  OAI21_X1   g18089(.A1(new_n18280_), .A2(new_n14871_), .B(new_n18281_), .ZN(new_n18282_));
  OAI22_X1   g18090(.A1(new_n18280_), .A2(new_n14871_), .B1(new_n17930_), .B2(new_n17922_), .ZN(new_n18283_));
  AOI22_X1   g18091(.A1(new_n18283_), .A2(\asqrt[16] ), .B1(new_n18282_), .B2(new_n17941_), .ZN(new_n18284_));
  INV_X1     g18092(.I(new_n17955_), .ZN(new_n18285_));
  OAI21_X1   g18093(.A1(new_n18284_), .A2(new_n13760_), .B(new_n18285_), .ZN(new_n18286_));
  NAND2_X1   g18094(.A1(new_n18286_), .A2(new_n17958_), .ZN(new_n18287_));
  AOI21_X1   g18095(.A1(new_n18283_), .A2(\asqrt[16] ), .B(new_n17946_), .ZN(new_n18288_));
  OAI22_X1   g18096(.A1(new_n18284_), .A2(new_n13760_), .B1(new_n18288_), .B2(new_n17950_), .ZN(new_n18289_));
  AOI21_X1   g18097(.A1(new_n18289_), .A2(\asqrt[18] ), .B(new_n17964_), .ZN(new_n18290_));
  NOR2_X1    g18098(.A1(new_n18290_), .A2(new_n18287_), .ZN(new_n18291_));
  AOI22_X1   g18099(.A1(new_n18289_), .A2(\asqrt[18] ), .B1(new_n18286_), .B2(new_n17958_), .ZN(new_n18292_));
  INV_X1     g18100(.I(new_n17973_), .ZN(new_n18293_));
  OAI21_X1   g18101(.A1(new_n18292_), .A2(new_n12657_), .B(new_n18293_), .ZN(new_n18294_));
  NAND2_X1   g18102(.A1(new_n18294_), .A2(new_n18291_), .ZN(new_n18295_));
  OAI22_X1   g18103(.A1(new_n18292_), .A2(new_n12657_), .B1(new_n18290_), .B2(new_n18287_), .ZN(new_n18296_));
  AOI21_X1   g18104(.A1(new_n18296_), .A2(\asqrt[20] ), .B(new_n17980_), .ZN(new_n18297_));
  NOR2_X1    g18105(.A1(new_n18297_), .A2(new_n18295_), .ZN(new_n18298_));
  AOI22_X1   g18106(.A1(new_n18296_), .A2(\asqrt[20] ), .B1(new_n18294_), .B2(new_n18291_), .ZN(new_n18299_));
  INV_X1     g18107(.I(new_n17988_), .ZN(new_n18300_));
  OAI21_X1   g18108(.A1(new_n18299_), .A2(new_n11631_), .B(new_n18300_), .ZN(new_n18301_));
  NAND2_X1   g18109(.A1(new_n18301_), .A2(new_n18298_), .ZN(new_n18302_));
  OAI22_X1   g18110(.A1(new_n18299_), .A2(new_n11631_), .B1(new_n18297_), .B2(new_n18295_), .ZN(new_n18303_));
  AOI21_X1   g18111(.A1(new_n18303_), .A2(\asqrt[22] ), .B(new_n17995_), .ZN(new_n18304_));
  NOR2_X1    g18112(.A1(new_n18304_), .A2(new_n18302_), .ZN(new_n18305_));
  AOI22_X1   g18113(.A1(new_n18303_), .A2(\asqrt[22] ), .B1(new_n18301_), .B2(new_n18298_), .ZN(new_n18306_));
  INV_X1     g18114(.I(new_n18003_), .ZN(new_n18307_));
  OAI21_X1   g18115(.A1(new_n18306_), .A2(new_n10614_), .B(new_n18307_), .ZN(new_n18308_));
  NAND2_X1   g18116(.A1(new_n18308_), .A2(new_n18305_), .ZN(new_n18309_));
  OAI22_X1   g18117(.A1(new_n18306_), .A2(new_n10614_), .B1(new_n18304_), .B2(new_n18302_), .ZN(new_n18310_));
  AOI21_X1   g18118(.A1(new_n18310_), .A2(\asqrt[24] ), .B(new_n18010_), .ZN(new_n18311_));
  NOR2_X1    g18119(.A1(new_n18311_), .A2(new_n18309_), .ZN(new_n18312_));
  AOI22_X1   g18120(.A1(new_n18310_), .A2(\asqrt[24] ), .B1(new_n18308_), .B2(new_n18305_), .ZN(new_n18313_));
  INV_X1     g18121(.I(new_n18018_), .ZN(new_n18314_));
  OAI21_X1   g18122(.A1(new_n18313_), .A2(new_n9672_), .B(new_n18314_), .ZN(new_n18315_));
  NAND2_X1   g18123(.A1(new_n18315_), .A2(new_n18312_), .ZN(new_n18316_));
  OAI22_X1   g18124(.A1(new_n18313_), .A2(new_n9672_), .B1(new_n18311_), .B2(new_n18309_), .ZN(new_n18317_));
  AOI21_X1   g18125(.A1(new_n18317_), .A2(\asqrt[26] ), .B(new_n18025_), .ZN(new_n18318_));
  NOR2_X1    g18126(.A1(new_n18318_), .A2(new_n18316_), .ZN(new_n18319_));
  AOI22_X1   g18127(.A1(new_n18317_), .A2(\asqrt[26] ), .B1(new_n18315_), .B2(new_n18312_), .ZN(new_n18320_));
  INV_X1     g18128(.I(new_n18033_), .ZN(new_n18321_));
  OAI21_X1   g18129(.A1(new_n18320_), .A2(new_n8763_), .B(new_n18321_), .ZN(new_n18322_));
  NAND2_X1   g18130(.A1(new_n18322_), .A2(new_n18319_), .ZN(new_n18323_));
  OAI22_X1   g18131(.A1(new_n18320_), .A2(new_n8763_), .B1(new_n18318_), .B2(new_n18316_), .ZN(new_n18324_));
  AOI21_X1   g18132(.A1(new_n18324_), .A2(\asqrt[28] ), .B(new_n18040_), .ZN(new_n18325_));
  NOR2_X1    g18133(.A1(new_n18325_), .A2(new_n18323_), .ZN(new_n18326_));
  AOI22_X1   g18134(.A1(new_n18324_), .A2(\asqrt[28] ), .B1(new_n18322_), .B2(new_n18319_), .ZN(new_n18327_));
  INV_X1     g18135(.I(new_n18048_), .ZN(new_n18328_));
  OAI21_X1   g18136(.A1(new_n18327_), .A2(new_n7931_), .B(new_n18328_), .ZN(new_n18329_));
  NAND2_X1   g18137(.A1(new_n18329_), .A2(new_n18326_), .ZN(new_n18330_));
  OAI22_X1   g18138(.A1(new_n18327_), .A2(new_n7931_), .B1(new_n18325_), .B2(new_n18323_), .ZN(new_n18331_));
  AOI21_X1   g18139(.A1(new_n18331_), .A2(\asqrt[30] ), .B(new_n18055_), .ZN(new_n18332_));
  NOR2_X1    g18140(.A1(new_n18332_), .A2(new_n18330_), .ZN(new_n18333_));
  AOI22_X1   g18141(.A1(new_n18331_), .A2(\asqrt[30] ), .B1(new_n18329_), .B2(new_n18326_), .ZN(new_n18334_));
  INV_X1     g18142(.I(new_n18063_), .ZN(new_n18335_));
  OAI21_X1   g18143(.A1(new_n18334_), .A2(new_n7110_), .B(new_n18335_), .ZN(new_n18336_));
  NAND2_X1   g18144(.A1(new_n18336_), .A2(new_n18333_), .ZN(new_n18337_));
  OAI22_X1   g18145(.A1(new_n18334_), .A2(new_n7110_), .B1(new_n18332_), .B2(new_n18330_), .ZN(new_n18338_));
  AOI21_X1   g18146(.A1(new_n18338_), .A2(\asqrt[32] ), .B(new_n18070_), .ZN(new_n18339_));
  NOR2_X1    g18147(.A1(new_n18339_), .A2(new_n18337_), .ZN(new_n18340_));
  AOI22_X1   g18148(.A1(new_n18338_), .A2(\asqrt[32] ), .B1(new_n18336_), .B2(new_n18333_), .ZN(new_n18341_));
  INV_X1     g18149(.I(new_n18078_), .ZN(new_n18342_));
  OAI21_X1   g18150(.A1(new_n18341_), .A2(new_n6365_), .B(new_n18342_), .ZN(new_n18343_));
  NAND2_X1   g18151(.A1(new_n18343_), .A2(new_n18340_), .ZN(new_n18344_));
  OAI22_X1   g18152(.A1(new_n18341_), .A2(new_n6365_), .B1(new_n18339_), .B2(new_n18337_), .ZN(new_n18345_));
  AOI21_X1   g18153(.A1(new_n18345_), .A2(\asqrt[34] ), .B(new_n18085_), .ZN(new_n18346_));
  NOR2_X1    g18154(.A1(new_n18346_), .A2(new_n18344_), .ZN(new_n18347_));
  AOI22_X1   g18155(.A1(new_n18345_), .A2(\asqrt[34] ), .B1(new_n18343_), .B2(new_n18340_), .ZN(new_n18348_));
  INV_X1     g18156(.I(new_n18093_), .ZN(new_n18349_));
  OAI21_X1   g18157(.A1(new_n18348_), .A2(new_n5626_), .B(new_n18349_), .ZN(new_n18350_));
  NAND2_X1   g18158(.A1(new_n18350_), .A2(new_n18347_), .ZN(new_n18351_));
  OAI22_X1   g18159(.A1(new_n18348_), .A2(new_n5626_), .B1(new_n18346_), .B2(new_n18344_), .ZN(new_n18352_));
  AOI21_X1   g18160(.A1(new_n18352_), .A2(\asqrt[36] ), .B(new_n18100_), .ZN(new_n18353_));
  NOR2_X1    g18161(.A1(new_n18353_), .A2(new_n18351_), .ZN(new_n18354_));
  AOI22_X1   g18162(.A1(new_n18352_), .A2(\asqrt[36] ), .B1(new_n18350_), .B2(new_n18347_), .ZN(new_n18355_));
  INV_X1     g18163(.I(new_n18108_), .ZN(new_n18356_));
  OAI21_X1   g18164(.A1(new_n18355_), .A2(new_n4973_), .B(new_n18356_), .ZN(new_n18357_));
  NAND2_X1   g18165(.A1(new_n18357_), .A2(new_n18354_), .ZN(new_n18358_));
  OAI22_X1   g18166(.A1(new_n18355_), .A2(new_n4973_), .B1(new_n18353_), .B2(new_n18351_), .ZN(new_n18359_));
  AOI21_X1   g18167(.A1(new_n18359_), .A2(\asqrt[38] ), .B(new_n18115_), .ZN(new_n18360_));
  NOR2_X1    g18168(.A1(new_n18360_), .A2(new_n18358_), .ZN(new_n18361_));
  AOI22_X1   g18169(.A1(new_n18359_), .A2(\asqrt[38] ), .B1(new_n18357_), .B2(new_n18354_), .ZN(new_n18362_));
  INV_X1     g18170(.I(new_n18123_), .ZN(new_n18363_));
  OAI21_X1   g18171(.A1(new_n18362_), .A2(new_n4330_), .B(new_n18363_), .ZN(new_n18364_));
  NAND2_X1   g18172(.A1(new_n18364_), .A2(new_n18361_), .ZN(new_n18365_));
  OAI22_X1   g18173(.A1(new_n18362_), .A2(new_n4330_), .B1(new_n18360_), .B2(new_n18358_), .ZN(new_n18366_));
  AOI21_X1   g18174(.A1(new_n18366_), .A2(\asqrt[40] ), .B(new_n18130_), .ZN(new_n18367_));
  NOR2_X1    g18175(.A1(new_n18367_), .A2(new_n18365_), .ZN(new_n18368_));
  AOI22_X1   g18176(.A1(new_n18366_), .A2(\asqrt[40] ), .B1(new_n18364_), .B2(new_n18361_), .ZN(new_n18369_));
  INV_X1     g18177(.I(new_n18138_), .ZN(new_n18370_));
  OAI21_X1   g18178(.A1(new_n18369_), .A2(new_n3760_), .B(new_n18370_), .ZN(new_n18371_));
  NAND2_X1   g18179(.A1(new_n18371_), .A2(new_n18368_), .ZN(new_n18372_));
  OAI22_X1   g18180(.A1(new_n18369_), .A2(new_n3760_), .B1(new_n18367_), .B2(new_n18365_), .ZN(new_n18373_));
  AOI21_X1   g18181(.A1(new_n18373_), .A2(\asqrt[42] ), .B(new_n18145_), .ZN(new_n18374_));
  NOR2_X1    g18182(.A1(new_n18374_), .A2(new_n18372_), .ZN(new_n18375_));
  AOI22_X1   g18183(.A1(new_n18373_), .A2(\asqrt[42] ), .B1(new_n18371_), .B2(new_n18368_), .ZN(new_n18376_));
  INV_X1     g18184(.I(new_n18153_), .ZN(new_n18377_));
  OAI21_X1   g18185(.A1(new_n18376_), .A2(new_n3208_), .B(new_n18377_), .ZN(new_n18378_));
  NAND2_X1   g18186(.A1(new_n18378_), .A2(new_n18375_), .ZN(new_n18379_));
  OAI22_X1   g18187(.A1(new_n18376_), .A2(new_n3208_), .B1(new_n18374_), .B2(new_n18372_), .ZN(new_n18380_));
  AOI21_X1   g18188(.A1(new_n18380_), .A2(\asqrt[44] ), .B(new_n18160_), .ZN(new_n18381_));
  NOR2_X1    g18189(.A1(new_n18381_), .A2(new_n18379_), .ZN(new_n18382_));
  AOI22_X1   g18190(.A1(new_n18380_), .A2(\asqrt[44] ), .B1(new_n18378_), .B2(new_n18375_), .ZN(new_n18383_));
  INV_X1     g18191(.I(new_n18168_), .ZN(new_n18384_));
  OAI21_X1   g18192(.A1(new_n18383_), .A2(new_n2728_), .B(new_n18384_), .ZN(new_n18385_));
  NAND2_X1   g18193(.A1(new_n18385_), .A2(new_n18382_), .ZN(new_n18386_));
  OAI22_X1   g18194(.A1(new_n18383_), .A2(new_n2728_), .B1(new_n18381_), .B2(new_n18379_), .ZN(new_n18387_));
  AOI21_X1   g18195(.A1(new_n18387_), .A2(\asqrt[46] ), .B(new_n18175_), .ZN(new_n18388_));
  NOR2_X1    g18196(.A1(new_n18388_), .A2(new_n18386_), .ZN(new_n18389_));
  AOI22_X1   g18197(.A1(new_n18387_), .A2(\asqrt[46] ), .B1(new_n18385_), .B2(new_n18382_), .ZN(new_n18390_));
  INV_X1     g18198(.I(new_n18183_), .ZN(new_n18391_));
  OAI21_X1   g18199(.A1(new_n18390_), .A2(new_n2253_), .B(new_n18391_), .ZN(new_n18392_));
  NAND2_X1   g18200(.A1(new_n18392_), .A2(new_n18389_), .ZN(new_n18393_));
  OAI22_X1   g18201(.A1(new_n18390_), .A2(new_n2253_), .B1(new_n18388_), .B2(new_n18386_), .ZN(new_n18394_));
  AOI21_X1   g18202(.A1(new_n18394_), .A2(\asqrt[48] ), .B(new_n18190_), .ZN(new_n18395_));
  NOR2_X1    g18203(.A1(new_n18395_), .A2(new_n18393_), .ZN(new_n18396_));
  AOI22_X1   g18204(.A1(new_n18394_), .A2(\asqrt[48] ), .B1(new_n18392_), .B2(new_n18389_), .ZN(new_n18397_));
  INV_X1     g18205(.I(new_n18198_), .ZN(new_n18398_));
  OAI21_X1   g18206(.A1(new_n18397_), .A2(new_n1854_), .B(new_n18398_), .ZN(new_n18399_));
  NAND2_X1   g18207(.A1(new_n18399_), .A2(new_n18396_), .ZN(new_n18400_));
  OAI22_X1   g18208(.A1(new_n18397_), .A2(new_n1854_), .B1(new_n18395_), .B2(new_n18393_), .ZN(new_n18401_));
  AOI21_X1   g18209(.A1(new_n18401_), .A2(\asqrt[50] ), .B(new_n18205_), .ZN(new_n18402_));
  NOR2_X1    g18210(.A1(new_n18402_), .A2(new_n18400_), .ZN(new_n18403_));
  AOI22_X1   g18211(.A1(new_n18401_), .A2(\asqrt[50] ), .B1(new_n18399_), .B2(new_n18396_), .ZN(new_n18404_));
  INV_X1     g18212(.I(new_n18213_), .ZN(new_n18405_));
  OAI21_X1   g18213(.A1(new_n18404_), .A2(new_n1436_), .B(new_n18405_), .ZN(new_n18406_));
  NAND2_X1   g18214(.A1(new_n18406_), .A2(new_n18403_), .ZN(new_n18407_));
  OAI22_X1   g18215(.A1(new_n18404_), .A2(new_n1436_), .B1(new_n18402_), .B2(new_n18400_), .ZN(new_n18408_));
  AOI21_X1   g18216(.A1(new_n18408_), .A2(\asqrt[52] ), .B(new_n18220_), .ZN(new_n18409_));
  NOR2_X1    g18217(.A1(new_n18409_), .A2(new_n18407_), .ZN(new_n18410_));
  AOI22_X1   g18218(.A1(new_n18408_), .A2(\asqrt[52] ), .B1(new_n18406_), .B2(new_n18403_), .ZN(new_n18411_));
  INV_X1     g18219(.I(new_n18228_), .ZN(new_n18412_));
  OAI21_X1   g18220(.A1(new_n18411_), .A2(new_n1096_), .B(new_n18412_), .ZN(new_n18413_));
  NAND2_X1   g18221(.A1(new_n18413_), .A2(new_n18410_), .ZN(new_n18414_));
  OAI22_X1   g18222(.A1(new_n18411_), .A2(new_n1096_), .B1(new_n18409_), .B2(new_n18407_), .ZN(new_n18415_));
  AOI21_X1   g18223(.A1(new_n18415_), .A2(\asqrt[54] ), .B(new_n18235_), .ZN(new_n18416_));
  NOR2_X1    g18224(.A1(new_n18416_), .A2(new_n18414_), .ZN(new_n18417_));
  AOI22_X1   g18225(.A1(new_n18415_), .A2(\asqrt[54] ), .B1(new_n18413_), .B2(new_n18410_), .ZN(new_n18418_));
  INV_X1     g18226(.I(new_n18243_), .ZN(new_n18419_));
  OAI21_X1   g18227(.A1(new_n18418_), .A2(new_n825_), .B(new_n18419_), .ZN(new_n18420_));
  NAND2_X1   g18228(.A1(new_n18420_), .A2(new_n18417_), .ZN(new_n18421_));
  OAI22_X1   g18229(.A1(new_n18418_), .A2(new_n825_), .B1(new_n18416_), .B2(new_n18414_), .ZN(new_n18422_));
  AOI21_X1   g18230(.A1(new_n18422_), .A2(\asqrt[56] ), .B(new_n18250_), .ZN(new_n18423_));
  NOR2_X1    g18231(.A1(new_n18423_), .A2(new_n18421_), .ZN(new_n18424_));
  AOI22_X1   g18232(.A1(new_n18422_), .A2(\asqrt[56] ), .B1(new_n18420_), .B2(new_n18417_), .ZN(new_n18425_));
  OAI21_X1   g18233(.A1(new_n18425_), .A2(new_n587_), .B(new_n18262_), .ZN(new_n18426_));
  NAND2_X1   g18234(.A1(new_n18426_), .A2(new_n18424_), .ZN(new_n18427_));
  NAND2_X1   g18235(.A1(new_n18415_), .A2(\asqrt[54] ), .ZN(new_n18428_));
  AOI21_X1   g18236(.A1(new_n18428_), .A2(new_n18414_), .B(new_n825_), .ZN(new_n18429_));
  OAI21_X1   g18237(.A1(new_n18417_), .A2(new_n18429_), .B(\asqrt[56] ), .ZN(new_n18430_));
  AOI21_X1   g18238(.A1(new_n18421_), .A2(new_n18430_), .B(new_n587_), .ZN(new_n18431_));
  OAI21_X1   g18239(.A1(new_n18424_), .A2(new_n18431_), .B(\asqrt[58] ), .ZN(new_n18432_));
  NAND2_X1   g18240(.A1(new_n18427_), .A2(new_n18432_), .ZN(new_n18433_));
  AOI22_X1   g18241(.A1(new_n18433_), .A2(\asqrt[59] ), .B1(new_n18270_), .B2(new_n18263_), .ZN(new_n18434_));
  NOR4_X1    g18242(.A1(new_n17893_), .A2(\asqrt[60] ), .A3(new_n17629_), .A4(new_n17846_), .ZN(new_n18435_));
  XOR2_X1    g18243(.A1(new_n18435_), .A2(new_n17861_), .Z(new_n18436_));
  NAND2_X1   g18244(.A1(new_n18436_), .A2(new_n229_), .ZN(new_n18437_));
  INV_X1     g18245(.I(new_n18437_), .ZN(new_n18438_));
  OAI21_X1   g18246(.A1(new_n18434_), .A2(new_n275_), .B(new_n18438_), .ZN(new_n18439_));
  NAND2_X1   g18247(.A1(new_n18439_), .A2(new_n18277_), .ZN(new_n18440_));
  OAI22_X1   g18248(.A1(new_n18425_), .A2(new_n587_), .B1(new_n18423_), .B2(new_n18421_), .ZN(new_n18441_));
  AOI21_X1   g18249(.A1(new_n18441_), .A2(\asqrt[58] ), .B(new_n18268_), .ZN(new_n18442_));
  NOR2_X1    g18250(.A1(new_n18442_), .A2(new_n18427_), .ZN(new_n18443_));
  AOI22_X1   g18251(.A1(new_n18441_), .A2(\asqrt[58] ), .B1(new_n18426_), .B2(new_n18424_), .ZN(new_n18444_));
  OAI21_X1   g18252(.A1(new_n18444_), .A2(new_n376_), .B(new_n18276_), .ZN(new_n18445_));
  NAND2_X1   g18253(.A1(new_n18445_), .A2(new_n18443_), .ZN(new_n18446_));
  AOI21_X1   g18254(.A1(new_n18427_), .A2(new_n18432_), .B(new_n376_), .ZN(new_n18447_));
  OAI21_X1   g18255(.A1(new_n18443_), .A2(new_n18447_), .B(\asqrt[60] ), .ZN(new_n18448_));
  AOI21_X1   g18256(.A1(new_n18446_), .A2(new_n18448_), .B(new_n229_), .ZN(new_n18449_));
  INV_X1     g18257(.I(new_n17865_), .ZN(new_n18450_));
  NOR2_X1    g18258(.A1(new_n18450_), .A2(\asqrt[62] ), .ZN(new_n18451_));
  INV_X1     g18259(.I(new_n18451_), .ZN(new_n18452_));
  NAND2_X1   g18260(.A1(new_n18449_), .A2(new_n18452_), .ZN(new_n18453_));
  OAI21_X1   g18261(.A1(new_n18453_), .A2(new_n18440_), .B(new_n17867_), .ZN(new_n18454_));
  NAND2_X1   g18262(.A1(new_n17655_), .A2(new_n17236_), .ZN(new_n18455_));
  OAI21_X1   g18263(.A1(\asqrt[10] ), .A2(new_n18455_), .B(new_n17648_), .ZN(new_n18456_));
  NAND2_X1   g18264(.A1(new_n18456_), .A2(new_n231_), .ZN(new_n18457_));
  OAI21_X1   g18265(.A1(new_n18454_), .A2(new_n18457_), .B(new_n17858_), .ZN(new_n18458_));
  OAI22_X1   g18266(.A1(new_n18444_), .A2(new_n376_), .B1(new_n18442_), .B2(new_n18427_), .ZN(new_n18459_));
  AOI21_X1   g18267(.A1(new_n18459_), .A2(\asqrt[60] ), .B(new_n18437_), .ZN(new_n18460_));
  AOI22_X1   g18268(.A1(new_n18459_), .A2(\asqrt[60] ), .B1(new_n18445_), .B2(new_n18443_), .ZN(new_n18461_));
  OAI22_X1   g18269(.A1(new_n18461_), .A2(new_n229_), .B1(new_n18460_), .B2(new_n18446_), .ZN(new_n18462_));
  NOR4_X1    g18270(.A1(new_n18462_), .A2(\asqrt[62] ), .A3(new_n17857_), .A4(new_n17865_), .ZN(new_n18463_));
  OAI21_X1   g18271(.A1(new_n17237_), .A2(new_n17648_), .B(\asqrt[10] ), .ZN(new_n18464_));
  XOR2_X1    g18272(.A1(new_n17648_), .A2(\asqrt[63] ), .Z(new_n18465_));
  NAND2_X1   g18273(.A1(new_n18464_), .A2(new_n18465_), .ZN(new_n18466_));
  INV_X1     g18274(.I(new_n18466_), .ZN(new_n18467_));
  NAND2_X1   g18275(.A1(new_n18463_), .A2(new_n18467_), .ZN(new_n18468_));
  NAND3_X1   g18276(.A1(new_n17887_), .A2(new_n17657_), .A3(new_n17237_), .ZN(new_n18469_));
  NOR4_X1    g18277(.A1(new_n18468_), .A2(new_n18458_), .A3(new_n17668_), .A4(new_n18469_), .ZN(new_n18470_));
  NOR2_X1    g18278(.A1(new_n17667_), .A2(\a[18] ), .ZN(new_n18471_));
  OAI21_X1   g18279(.A1(new_n18470_), .A2(new_n18471_), .B(new_n17667_), .ZN(new_n18472_));
  INV_X1     g18280(.I(new_n17667_), .ZN(new_n18473_));
  NOR2_X1    g18281(.A1(new_n18460_), .A2(new_n18446_), .ZN(new_n18474_));
  NOR3_X1    g18282(.A1(new_n18461_), .A2(new_n229_), .A3(new_n18451_), .ZN(new_n18475_));
  AOI21_X1   g18283(.A1(new_n18475_), .A2(new_n18474_), .B(new_n17866_), .ZN(new_n18476_));
  INV_X1     g18284(.I(new_n18457_), .ZN(new_n18477_));
  AOI21_X1   g18285(.A1(new_n18476_), .A2(new_n18477_), .B(new_n17857_), .ZN(new_n18478_));
  AOI21_X1   g18286(.A1(new_n18462_), .A2(\asqrt[62] ), .B(new_n17858_), .ZN(new_n18479_));
  AOI21_X1   g18287(.A1(new_n18271_), .A2(new_n18273_), .B(new_n275_), .ZN(new_n18480_));
  OAI21_X1   g18288(.A1(new_n18277_), .A2(new_n18480_), .B(\asqrt[61] ), .ZN(new_n18481_));
  NAND4_X1   g18289(.A1(new_n18440_), .A2(new_n196_), .A3(new_n18481_), .A4(new_n18450_), .ZN(new_n18482_));
  NOR3_X1    g18290(.A1(new_n18479_), .A2(new_n18482_), .A3(new_n18466_), .ZN(new_n18483_));
  INV_X1     g18291(.I(new_n18469_), .ZN(new_n18484_));
  NAND4_X1   g18292(.A1(new_n18483_), .A2(\a[19] ), .A3(new_n18478_), .A4(new_n18484_), .ZN(new_n18485_));
  NAND3_X1   g18293(.A1(new_n18485_), .A2(\a[18] ), .A3(new_n18473_), .ZN(new_n18486_));
  NAND2_X1   g18294(.A1(new_n18472_), .A2(new_n18486_), .ZN(new_n18487_));
  NAND2_X1   g18295(.A1(new_n17880_), .A2(new_n17650_), .ZN(new_n18488_));
  NOR2_X1    g18296(.A1(new_n18468_), .A2(new_n18458_), .ZN(new_n18489_));
  NAND4_X1   g18297(.A1(new_n17883_), .A2(new_n17658_), .A3(new_n17237_), .A4(new_n18488_), .ZN(new_n18490_));
  NOR2_X1    g18298(.A1(new_n17893_), .A2(new_n17656_), .ZN(new_n18491_));
  XOR2_X1    g18299(.A1(new_n18491_), .A2(new_n18490_), .Z(new_n18492_));
  NOR2_X1    g18300(.A1(new_n18492_), .A2(new_n17664_), .ZN(new_n18493_));
  INV_X1     g18301(.I(new_n18493_), .ZN(new_n18494_));
  NAND3_X1   g18302(.A1(new_n18483_), .A2(new_n18478_), .A3(new_n18484_), .ZN(new_n18495_));
  NOR4_X1    g18303(.A1(new_n18481_), .A2(new_n18446_), .A3(new_n18460_), .A4(new_n18451_), .ZN(new_n18496_));
  NOR3_X1    g18304(.A1(new_n18496_), .A2(new_n17866_), .A3(new_n18457_), .ZN(new_n18497_));
  NAND2_X1   g18305(.A1(new_n18446_), .A2(new_n18448_), .ZN(new_n18498_));
  AOI22_X1   g18306(.A1(new_n18498_), .A2(\asqrt[61] ), .B1(new_n18439_), .B2(new_n18277_), .ZN(new_n18499_));
  NAND4_X1   g18307(.A1(new_n18499_), .A2(new_n196_), .A3(new_n17858_), .A4(new_n18450_), .ZN(new_n18500_));
  OAI21_X1   g18308(.A1(new_n18497_), .A2(new_n17857_), .B(new_n18500_), .ZN(new_n18501_));
  NOR2_X1    g18309(.A1(new_n18467_), .A2(new_n18484_), .ZN(new_n18502_));
  NAND2_X1   g18310(.A1(new_n18502_), .A2(\asqrt[10] ), .ZN(new_n18503_));
  OAI21_X1   g18311(.A1(new_n18501_), .A2(new_n18503_), .B(new_n17868_), .ZN(new_n18504_));
  NAND3_X1   g18312(.A1(new_n18504_), .A2(new_n17869_), .A3(new_n18495_), .ZN(new_n18505_));
  NOR3_X1    g18313(.A1(new_n18468_), .A2(new_n18458_), .A3(new_n18469_), .ZN(\asqrt[9] ));
  NAND3_X1   g18314(.A1(new_n18474_), .A2(new_n18449_), .A3(new_n18452_), .ZN(new_n18507_));
  NAND3_X1   g18315(.A1(new_n18507_), .A2(new_n17867_), .A3(new_n18477_), .ZN(new_n18508_));
  AOI21_X1   g18316(.A1(new_n18508_), .A2(new_n17858_), .B(new_n18463_), .ZN(new_n18509_));
  INV_X1     g18317(.I(new_n18503_), .ZN(new_n18510_));
  AOI21_X1   g18318(.A1(new_n18509_), .A2(new_n18510_), .B(\a[20] ), .ZN(new_n18511_));
  OAI21_X1   g18319(.A1(new_n18511_), .A2(new_n17870_), .B(\asqrt[9] ), .ZN(new_n18512_));
  NAND4_X1   g18320(.A1(new_n18505_), .A2(new_n18512_), .A3(new_n17271_), .A4(new_n18494_), .ZN(new_n18513_));
  NAND2_X1   g18321(.A1(new_n18513_), .A2(new_n18487_), .ZN(new_n18514_));
  NAND3_X1   g18322(.A1(new_n18472_), .A2(new_n18486_), .A3(new_n18494_), .ZN(new_n18515_));
  AOI21_X1   g18323(.A1(\asqrt[10] ), .A2(new_n17868_), .B(\a[21] ), .ZN(new_n18516_));
  NOR2_X1    g18324(.A1(new_n17884_), .A2(\a[20] ), .ZN(new_n18517_));
  AOI21_X1   g18325(.A1(\asqrt[10] ), .A2(\a[20] ), .B(new_n17872_), .ZN(new_n18518_));
  OAI21_X1   g18326(.A1(new_n18517_), .A2(new_n18516_), .B(new_n18518_), .ZN(new_n18519_));
  INV_X1     g18327(.I(new_n18519_), .ZN(new_n18520_));
  NAND3_X1   g18328(.A1(\asqrt[9] ), .A2(new_n17892_), .A3(new_n18520_), .ZN(new_n18521_));
  OAI21_X1   g18329(.A1(new_n18495_), .A2(new_n18519_), .B(new_n17891_), .ZN(new_n18522_));
  NAND3_X1   g18330(.A1(new_n18521_), .A2(new_n18522_), .A3(new_n16619_), .ZN(new_n18523_));
  AOI21_X1   g18331(.A1(new_n18515_), .A2(\asqrt[11] ), .B(new_n18523_), .ZN(new_n18524_));
  NOR2_X1    g18332(.A1(new_n18514_), .A2(new_n18524_), .ZN(new_n18525_));
  AOI22_X1   g18333(.A1(new_n18513_), .A2(new_n18487_), .B1(\asqrt[11] ), .B2(new_n18515_), .ZN(new_n18526_));
  INV_X1     g18334(.I(new_n17876_), .ZN(new_n18527_));
  AOI21_X1   g18335(.A1(new_n17884_), .A2(new_n18527_), .B(new_n17878_), .ZN(new_n18528_));
  INV_X1     g18336(.I(new_n17885_), .ZN(new_n18529_));
  NOR3_X1    g18337(.A1(new_n18529_), .A2(new_n18528_), .A3(new_n17891_), .ZN(new_n18530_));
  AOI21_X1   g18338(.A1(new_n17901_), .A2(new_n17898_), .B(\asqrt[12] ), .ZN(new_n18531_));
  AND4_X2    g18339(.A1(new_n18530_), .A2(\asqrt[9] ), .A3(new_n17915_), .A4(new_n18531_), .Z(new_n18532_));
  NOR2_X1    g18340(.A1(new_n18530_), .A2(new_n16619_), .ZN(new_n18533_));
  NOR3_X1    g18341(.A1(new_n18532_), .A2(\asqrt[13] ), .A3(new_n18533_), .ZN(new_n18534_));
  OAI21_X1   g18342(.A1(new_n18526_), .A2(new_n16619_), .B(new_n18534_), .ZN(new_n18535_));
  NAND2_X1   g18343(.A1(new_n18535_), .A2(new_n18525_), .ZN(new_n18536_));
  OAI22_X1   g18344(.A1(new_n18526_), .A2(new_n16619_), .B1(new_n18514_), .B2(new_n18524_), .ZN(new_n18537_));
  NAND2_X1   g18345(.A1(new_n17910_), .A2(new_n17911_), .ZN(new_n18538_));
  NAND4_X1   g18346(.A1(\asqrt[9] ), .A2(new_n16060_), .A3(new_n18538_), .A4(new_n17923_), .ZN(new_n18539_));
  XOR2_X1    g18347(.A1(new_n18539_), .A2(new_n17916_), .Z(new_n18540_));
  NAND2_X1   g18348(.A1(new_n18540_), .A2(new_n15447_), .ZN(new_n18541_));
  AOI21_X1   g18349(.A1(new_n18537_), .A2(\asqrt[13] ), .B(new_n18541_), .ZN(new_n18542_));
  NOR2_X1    g18350(.A1(new_n18542_), .A2(new_n18536_), .ZN(new_n18543_));
  AOI22_X1   g18351(.A1(new_n18537_), .A2(\asqrt[13] ), .B1(new_n18535_), .B2(new_n18525_), .ZN(new_n18544_));
  NOR4_X1    g18352(.A1(new_n18495_), .A2(\asqrt[14] ), .A3(new_n17920_), .A4(new_n17924_), .ZN(new_n18545_));
  XOR2_X1    g18353(.A1(new_n18545_), .A2(new_n17931_), .Z(new_n18546_));
  NAND2_X1   g18354(.A1(new_n18546_), .A2(new_n14871_), .ZN(new_n18547_));
  INV_X1     g18355(.I(new_n18547_), .ZN(new_n18548_));
  OAI21_X1   g18356(.A1(new_n18544_), .A2(new_n15447_), .B(new_n18548_), .ZN(new_n18549_));
  NAND2_X1   g18357(.A1(new_n18549_), .A2(new_n18543_), .ZN(new_n18550_));
  OAI22_X1   g18358(.A1(new_n18544_), .A2(new_n15447_), .B1(new_n18542_), .B2(new_n18536_), .ZN(new_n18551_));
  NOR2_X1    g18359(.A1(new_n17928_), .A2(\asqrt[15] ), .ZN(new_n18552_));
  NAND3_X1   g18360(.A1(\asqrt[9] ), .A2(new_n18280_), .A3(new_n18552_), .ZN(new_n18553_));
  XOR2_X1    g18361(.A1(new_n18553_), .A2(new_n17932_), .Z(new_n18554_));
  NAND2_X1   g18362(.A1(new_n18554_), .A2(new_n14273_), .ZN(new_n18555_));
  AOI21_X1   g18363(.A1(new_n18551_), .A2(\asqrt[15] ), .B(new_n18555_), .ZN(new_n18556_));
  NOR2_X1    g18364(.A1(new_n18556_), .A2(new_n18550_), .ZN(new_n18557_));
  AOI22_X1   g18365(.A1(new_n18551_), .A2(\asqrt[15] ), .B1(new_n18549_), .B2(new_n18543_), .ZN(new_n18558_));
  NOR4_X1    g18366(.A1(new_n18495_), .A2(\asqrt[16] ), .A3(new_n17936_), .A4(new_n18283_), .ZN(new_n18559_));
  XOR2_X1    g18367(.A1(new_n18559_), .A2(new_n17942_), .Z(new_n18560_));
  NAND2_X1   g18368(.A1(new_n18560_), .A2(new_n13760_), .ZN(new_n18561_));
  INV_X1     g18369(.I(new_n18561_), .ZN(new_n18562_));
  OAI21_X1   g18370(.A1(new_n18558_), .A2(new_n14273_), .B(new_n18562_), .ZN(new_n18563_));
  NAND2_X1   g18371(.A1(new_n18563_), .A2(new_n18557_), .ZN(new_n18564_));
  OAI22_X1   g18372(.A1(new_n18558_), .A2(new_n14273_), .B1(new_n18556_), .B2(new_n18550_), .ZN(new_n18565_));
  NOR4_X1    g18373(.A1(new_n18495_), .A2(\asqrt[17] ), .A3(new_n17945_), .A4(new_n17951_), .ZN(new_n18566_));
  XNOR2_X1   g18374(.A1(new_n18566_), .A2(new_n17959_), .ZN(new_n18567_));
  NAND2_X1   g18375(.A1(new_n18567_), .A2(new_n13192_), .ZN(new_n18568_));
  AOI21_X1   g18376(.A1(new_n18565_), .A2(\asqrt[17] ), .B(new_n18568_), .ZN(new_n18569_));
  NOR2_X1    g18377(.A1(new_n18569_), .A2(new_n18564_), .ZN(new_n18570_));
  AOI22_X1   g18378(.A1(new_n18565_), .A2(\asqrt[17] ), .B1(new_n18563_), .B2(new_n18557_), .ZN(new_n18571_));
  NOR4_X1    g18379(.A1(new_n18495_), .A2(\asqrt[18] ), .A3(new_n17954_), .A4(new_n18289_), .ZN(new_n18572_));
  XOR2_X1    g18380(.A1(new_n18572_), .A2(new_n17960_), .Z(new_n18573_));
  NAND2_X1   g18381(.A1(new_n18573_), .A2(new_n12657_), .ZN(new_n18574_));
  INV_X1     g18382(.I(new_n18574_), .ZN(new_n18575_));
  OAI21_X1   g18383(.A1(new_n18571_), .A2(new_n13192_), .B(new_n18575_), .ZN(new_n18576_));
  NAND2_X1   g18384(.A1(new_n18576_), .A2(new_n18570_), .ZN(new_n18577_));
  OAI22_X1   g18385(.A1(new_n18571_), .A2(new_n13192_), .B1(new_n18569_), .B2(new_n18564_), .ZN(new_n18578_));
  NAND2_X1   g18386(.A1(new_n17969_), .A2(\asqrt[19] ), .ZN(new_n18579_));
  NOR4_X1    g18387(.A1(new_n18495_), .A2(\asqrt[19] ), .A3(new_n17963_), .A4(new_n17969_), .ZN(new_n18580_));
  XOR2_X1    g18388(.A1(new_n18580_), .A2(new_n18579_), .Z(new_n18581_));
  NAND2_X1   g18389(.A1(new_n18581_), .A2(new_n12101_), .ZN(new_n18582_));
  AOI21_X1   g18390(.A1(new_n18578_), .A2(\asqrt[19] ), .B(new_n18582_), .ZN(new_n18583_));
  NOR2_X1    g18391(.A1(new_n18583_), .A2(new_n18577_), .ZN(new_n18584_));
  AOI22_X1   g18392(.A1(new_n18578_), .A2(\asqrt[19] ), .B1(new_n18576_), .B2(new_n18570_), .ZN(new_n18585_));
  NOR4_X1    g18393(.A1(new_n18495_), .A2(\asqrt[20] ), .A3(new_n17972_), .A4(new_n18296_), .ZN(new_n18586_));
  AOI21_X1   g18394(.A1(new_n18579_), .A2(new_n17967_), .B(new_n12101_), .ZN(new_n18587_));
  NOR2_X1    g18395(.A1(new_n18586_), .A2(new_n18587_), .ZN(new_n18588_));
  NAND2_X1   g18396(.A1(new_n18588_), .A2(new_n11631_), .ZN(new_n18589_));
  INV_X1     g18397(.I(new_n18589_), .ZN(new_n18590_));
  OAI21_X1   g18398(.A1(new_n18585_), .A2(new_n12101_), .B(new_n18590_), .ZN(new_n18591_));
  NAND2_X1   g18399(.A1(new_n18591_), .A2(new_n18584_), .ZN(new_n18592_));
  OAI22_X1   g18400(.A1(new_n18585_), .A2(new_n12101_), .B1(new_n18583_), .B2(new_n18577_), .ZN(new_n18593_));
  NAND2_X1   g18401(.A1(new_n17984_), .A2(\asqrt[21] ), .ZN(new_n18594_));
  NOR4_X1    g18402(.A1(new_n18495_), .A2(\asqrt[21] ), .A3(new_n17979_), .A4(new_n17984_), .ZN(new_n18595_));
  XOR2_X1    g18403(.A1(new_n18595_), .A2(new_n18594_), .Z(new_n18596_));
  NAND2_X1   g18404(.A1(new_n18596_), .A2(new_n11105_), .ZN(new_n18597_));
  AOI21_X1   g18405(.A1(new_n18593_), .A2(\asqrt[21] ), .B(new_n18597_), .ZN(new_n18598_));
  NOR2_X1    g18406(.A1(new_n18598_), .A2(new_n18592_), .ZN(new_n18599_));
  AOI22_X1   g18407(.A1(new_n18593_), .A2(\asqrt[21] ), .B1(new_n18591_), .B2(new_n18584_), .ZN(new_n18600_));
  NOR4_X1    g18408(.A1(new_n18495_), .A2(\asqrt[22] ), .A3(new_n17987_), .A4(new_n18303_), .ZN(new_n18601_));
  AOI21_X1   g18409(.A1(new_n18594_), .A2(new_n17983_), .B(new_n11105_), .ZN(new_n18602_));
  NOR2_X1    g18410(.A1(new_n18601_), .A2(new_n18602_), .ZN(new_n18603_));
  NAND2_X1   g18411(.A1(new_n18603_), .A2(new_n10614_), .ZN(new_n18604_));
  INV_X1     g18412(.I(new_n18604_), .ZN(new_n18605_));
  OAI21_X1   g18413(.A1(new_n18600_), .A2(new_n11105_), .B(new_n18605_), .ZN(new_n18606_));
  NAND2_X1   g18414(.A1(new_n18606_), .A2(new_n18599_), .ZN(new_n18607_));
  OAI22_X1   g18415(.A1(new_n18600_), .A2(new_n11105_), .B1(new_n18598_), .B2(new_n18592_), .ZN(new_n18608_));
  NAND2_X1   g18416(.A1(new_n17999_), .A2(\asqrt[23] ), .ZN(new_n18609_));
  NOR4_X1    g18417(.A1(new_n18495_), .A2(\asqrt[23] ), .A3(new_n17994_), .A4(new_n17999_), .ZN(new_n18610_));
  XOR2_X1    g18418(.A1(new_n18610_), .A2(new_n18609_), .Z(new_n18611_));
  NAND2_X1   g18419(.A1(new_n18611_), .A2(new_n10104_), .ZN(new_n18612_));
  AOI21_X1   g18420(.A1(new_n18608_), .A2(\asqrt[23] ), .B(new_n18612_), .ZN(new_n18613_));
  NOR2_X1    g18421(.A1(new_n18613_), .A2(new_n18607_), .ZN(new_n18614_));
  AOI22_X1   g18422(.A1(new_n18608_), .A2(\asqrt[23] ), .B1(new_n18606_), .B2(new_n18599_), .ZN(new_n18615_));
  NOR4_X1    g18423(.A1(new_n18495_), .A2(\asqrt[24] ), .A3(new_n18002_), .A4(new_n18310_), .ZN(new_n18616_));
  AOI21_X1   g18424(.A1(new_n18609_), .A2(new_n17998_), .B(new_n10104_), .ZN(new_n18617_));
  NOR2_X1    g18425(.A1(new_n18616_), .A2(new_n18617_), .ZN(new_n18618_));
  NAND2_X1   g18426(.A1(new_n18618_), .A2(new_n9672_), .ZN(new_n18619_));
  INV_X1     g18427(.I(new_n18619_), .ZN(new_n18620_));
  OAI21_X1   g18428(.A1(new_n18615_), .A2(new_n10104_), .B(new_n18620_), .ZN(new_n18621_));
  NAND2_X1   g18429(.A1(new_n18621_), .A2(new_n18614_), .ZN(new_n18622_));
  OAI22_X1   g18430(.A1(new_n18615_), .A2(new_n10104_), .B1(new_n18613_), .B2(new_n18607_), .ZN(new_n18623_));
  NAND2_X1   g18431(.A1(new_n18014_), .A2(\asqrt[25] ), .ZN(new_n18624_));
  NOR4_X1    g18432(.A1(new_n18495_), .A2(\asqrt[25] ), .A3(new_n18009_), .A4(new_n18014_), .ZN(new_n18625_));
  XOR2_X1    g18433(.A1(new_n18625_), .A2(new_n18624_), .Z(new_n18626_));
  NAND2_X1   g18434(.A1(new_n18626_), .A2(new_n9212_), .ZN(new_n18627_));
  AOI21_X1   g18435(.A1(new_n18623_), .A2(\asqrt[25] ), .B(new_n18627_), .ZN(new_n18628_));
  NOR2_X1    g18436(.A1(new_n18628_), .A2(new_n18622_), .ZN(new_n18629_));
  AOI22_X1   g18437(.A1(new_n18623_), .A2(\asqrt[25] ), .B1(new_n18621_), .B2(new_n18614_), .ZN(new_n18630_));
  NOR4_X1    g18438(.A1(new_n18495_), .A2(\asqrt[26] ), .A3(new_n18017_), .A4(new_n18317_), .ZN(new_n18631_));
  AOI21_X1   g18439(.A1(new_n18624_), .A2(new_n18013_), .B(new_n9212_), .ZN(new_n18632_));
  NOR2_X1    g18440(.A1(new_n18631_), .A2(new_n18632_), .ZN(new_n18633_));
  NAND2_X1   g18441(.A1(new_n18633_), .A2(new_n8763_), .ZN(new_n18634_));
  INV_X1     g18442(.I(new_n18634_), .ZN(new_n18635_));
  OAI21_X1   g18443(.A1(new_n18630_), .A2(new_n9212_), .B(new_n18635_), .ZN(new_n18636_));
  NAND2_X1   g18444(.A1(new_n18636_), .A2(new_n18629_), .ZN(new_n18637_));
  OAI22_X1   g18445(.A1(new_n18630_), .A2(new_n9212_), .B1(new_n18628_), .B2(new_n18622_), .ZN(new_n18638_));
  NAND2_X1   g18446(.A1(new_n18029_), .A2(\asqrt[27] ), .ZN(new_n18639_));
  NOR4_X1    g18447(.A1(new_n18495_), .A2(\asqrt[27] ), .A3(new_n18024_), .A4(new_n18029_), .ZN(new_n18640_));
  XOR2_X1    g18448(.A1(new_n18640_), .A2(new_n18639_), .Z(new_n18641_));
  NAND2_X1   g18449(.A1(new_n18641_), .A2(new_n8319_), .ZN(new_n18642_));
  AOI21_X1   g18450(.A1(new_n18638_), .A2(\asqrt[27] ), .B(new_n18642_), .ZN(new_n18643_));
  NOR2_X1    g18451(.A1(new_n18643_), .A2(new_n18637_), .ZN(new_n18644_));
  AOI22_X1   g18452(.A1(new_n18638_), .A2(\asqrt[27] ), .B1(new_n18636_), .B2(new_n18629_), .ZN(new_n18645_));
  NOR4_X1    g18453(.A1(new_n18495_), .A2(\asqrt[28] ), .A3(new_n18032_), .A4(new_n18324_), .ZN(new_n18646_));
  AOI21_X1   g18454(.A1(new_n18639_), .A2(new_n18028_), .B(new_n8319_), .ZN(new_n18647_));
  NOR2_X1    g18455(.A1(new_n18646_), .A2(new_n18647_), .ZN(new_n18648_));
  NAND2_X1   g18456(.A1(new_n18648_), .A2(new_n7931_), .ZN(new_n18649_));
  INV_X1     g18457(.I(new_n18649_), .ZN(new_n18650_));
  OAI21_X1   g18458(.A1(new_n18645_), .A2(new_n8319_), .B(new_n18650_), .ZN(new_n18651_));
  NAND2_X1   g18459(.A1(new_n18651_), .A2(new_n18644_), .ZN(new_n18652_));
  OAI22_X1   g18460(.A1(new_n18645_), .A2(new_n8319_), .B1(new_n18643_), .B2(new_n18637_), .ZN(new_n18653_));
  NAND2_X1   g18461(.A1(new_n18044_), .A2(\asqrt[29] ), .ZN(new_n18654_));
  NOR4_X1    g18462(.A1(new_n18495_), .A2(\asqrt[29] ), .A3(new_n18039_), .A4(new_n18044_), .ZN(new_n18655_));
  XOR2_X1    g18463(.A1(new_n18655_), .A2(new_n18654_), .Z(new_n18656_));
  NAND2_X1   g18464(.A1(new_n18656_), .A2(new_n7517_), .ZN(new_n18657_));
  AOI21_X1   g18465(.A1(new_n18653_), .A2(\asqrt[29] ), .B(new_n18657_), .ZN(new_n18658_));
  NOR2_X1    g18466(.A1(new_n18658_), .A2(new_n18652_), .ZN(new_n18659_));
  AOI22_X1   g18467(.A1(new_n18653_), .A2(\asqrt[29] ), .B1(new_n18651_), .B2(new_n18644_), .ZN(new_n18660_));
  NAND2_X1   g18468(.A1(new_n18331_), .A2(\asqrt[30] ), .ZN(new_n18661_));
  NOR4_X1    g18469(.A1(new_n18495_), .A2(\asqrt[30] ), .A3(new_n18047_), .A4(new_n18331_), .ZN(new_n18662_));
  XOR2_X1    g18470(.A1(new_n18662_), .A2(new_n18661_), .Z(new_n18663_));
  NAND2_X1   g18471(.A1(new_n18663_), .A2(new_n7110_), .ZN(new_n18664_));
  INV_X1     g18472(.I(new_n18664_), .ZN(new_n18665_));
  OAI21_X1   g18473(.A1(new_n18660_), .A2(new_n7517_), .B(new_n18665_), .ZN(new_n18666_));
  NAND2_X1   g18474(.A1(new_n18666_), .A2(new_n18659_), .ZN(new_n18667_));
  OAI22_X1   g18475(.A1(new_n18660_), .A2(new_n7517_), .B1(new_n18658_), .B2(new_n18652_), .ZN(new_n18668_));
  NOR4_X1    g18476(.A1(new_n18495_), .A2(\asqrt[31] ), .A3(new_n18054_), .A4(new_n18059_), .ZN(new_n18669_));
  AOI21_X1   g18477(.A1(new_n18661_), .A2(new_n18330_), .B(new_n7110_), .ZN(new_n18670_));
  NOR2_X1    g18478(.A1(new_n18669_), .A2(new_n18670_), .ZN(new_n18671_));
  NAND2_X1   g18479(.A1(new_n18671_), .A2(new_n6708_), .ZN(new_n18672_));
  AOI21_X1   g18480(.A1(new_n18668_), .A2(\asqrt[31] ), .B(new_n18672_), .ZN(new_n18673_));
  NOR2_X1    g18481(.A1(new_n18673_), .A2(new_n18667_), .ZN(new_n18674_));
  AOI22_X1   g18482(.A1(new_n18668_), .A2(\asqrt[31] ), .B1(new_n18666_), .B2(new_n18659_), .ZN(new_n18675_));
  NAND2_X1   g18483(.A1(new_n18338_), .A2(\asqrt[32] ), .ZN(new_n18676_));
  NOR4_X1    g18484(.A1(new_n18495_), .A2(\asqrt[32] ), .A3(new_n18062_), .A4(new_n18338_), .ZN(new_n18677_));
  XOR2_X1    g18485(.A1(new_n18677_), .A2(new_n18676_), .Z(new_n18678_));
  NAND2_X1   g18486(.A1(new_n18678_), .A2(new_n6365_), .ZN(new_n18679_));
  INV_X1     g18487(.I(new_n18679_), .ZN(new_n18680_));
  OAI21_X1   g18488(.A1(new_n18675_), .A2(new_n6708_), .B(new_n18680_), .ZN(new_n18681_));
  NAND2_X1   g18489(.A1(new_n18681_), .A2(new_n18674_), .ZN(new_n18682_));
  OAI22_X1   g18490(.A1(new_n18675_), .A2(new_n6708_), .B1(new_n18673_), .B2(new_n18667_), .ZN(new_n18683_));
  NOR4_X1    g18491(.A1(new_n18495_), .A2(\asqrt[33] ), .A3(new_n18069_), .A4(new_n18074_), .ZN(new_n18684_));
  AOI21_X1   g18492(.A1(new_n18676_), .A2(new_n18337_), .B(new_n6365_), .ZN(new_n18685_));
  NOR2_X1    g18493(.A1(new_n18684_), .A2(new_n18685_), .ZN(new_n18686_));
  NAND2_X1   g18494(.A1(new_n18686_), .A2(new_n5991_), .ZN(new_n18687_));
  AOI21_X1   g18495(.A1(new_n18683_), .A2(\asqrt[33] ), .B(new_n18687_), .ZN(new_n18688_));
  NOR2_X1    g18496(.A1(new_n18688_), .A2(new_n18682_), .ZN(new_n18689_));
  AOI22_X1   g18497(.A1(new_n18683_), .A2(\asqrt[33] ), .B1(new_n18681_), .B2(new_n18674_), .ZN(new_n18690_));
  NAND2_X1   g18498(.A1(new_n18345_), .A2(\asqrt[34] ), .ZN(new_n18691_));
  NOR4_X1    g18499(.A1(new_n18495_), .A2(\asqrt[34] ), .A3(new_n18077_), .A4(new_n18345_), .ZN(new_n18692_));
  XOR2_X1    g18500(.A1(new_n18692_), .A2(new_n18691_), .Z(new_n18693_));
  NAND2_X1   g18501(.A1(new_n18693_), .A2(new_n5626_), .ZN(new_n18694_));
  INV_X1     g18502(.I(new_n18694_), .ZN(new_n18695_));
  OAI21_X1   g18503(.A1(new_n18690_), .A2(new_n5991_), .B(new_n18695_), .ZN(new_n18696_));
  NAND2_X1   g18504(.A1(new_n18696_), .A2(new_n18689_), .ZN(new_n18697_));
  OAI22_X1   g18505(.A1(new_n18690_), .A2(new_n5991_), .B1(new_n18688_), .B2(new_n18682_), .ZN(new_n18698_));
  NAND2_X1   g18506(.A1(new_n18089_), .A2(\asqrt[35] ), .ZN(new_n18699_));
  NOR4_X1    g18507(.A1(new_n18495_), .A2(\asqrt[35] ), .A3(new_n18084_), .A4(new_n18089_), .ZN(new_n18700_));
  XOR2_X1    g18508(.A1(new_n18700_), .A2(new_n18699_), .Z(new_n18701_));
  NAND2_X1   g18509(.A1(new_n18701_), .A2(new_n5273_), .ZN(new_n18702_));
  AOI21_X1   g18510(.A1(new_n18698_), .A2(\asqrt[35] ), .B(new_n18702_), .ZN(new_n18703_));
  NOR2_X1    g18511(.A1(new_n18703_), .A2(new_n18697_), .ZN(new_n18704_));
  AOI22_X1   g18512(.A1(new_n18698_), .A2(\asqrt[35] ), .B1(new_n18696_), .B2(new_n18689_), .ZN(new_n18705_));
  NOR4_X1    g18513(.A1(new_n18495_), .A2(\asqrt[36] ), .A3(new_n18092_), .A4(new_n18352_), .ZN(new_n18706_));
  AOI21_X1   g18514(.A1(new_n18699_), .A2(new_n18088_), .B(new_n5273_), .ZN(new_n18707_));
  NOR2_X1    g18515(.A1(new_n18706_), .A2(new_n18707_), .ZN(new_n18708_));
  NAND2_X1   g18516(.A1(new_n18708_), .A2(new_n4973_), .ZN(new_n18709_));
  INV_X1     g18517(.I(new_n18709_), .ZN(new_n18710_));
  OAI21_X1   g18518(.A1(new_n18705_), .A2(new_n5273_), .B(new_n18710_), .ZN(new_n18711_));
  NAND2_X1   g18519(.A1(new_n18711_), .A2(new_n18704_), .ZN(new_n18712_));
  OAI22_X1   g18520(.A1(new_n18705_), .A2(new_n5273_), .B1(new_n18703_), .B2(new_n18697_), .ZN(new_n18713_));
  NAND2_X1   g18521(.A1(new_n18104_), .A2(\asqrt[37] ), .ZN(new_n18714_));
  NOR4_X1    g18522(.A1(new_n18495_), .A2(\asqrt[37] ), .A3(new_n18099_), .A4(new_n18104_), .ZN(new_n18715_));
  XOR2_X1    g18523(.A1(new_n18715_), .A2(new_n18714_), .Z(new_n18716_));
  NAND2_X1   g18524(.A1(new_n18716_), .A2(new_n4645_), .ZN(new_n18717_));
  AOI21_X1   g18525(.A1(new_n18713_), .A2(\asqrt[37] ), .B(new_n18717_), .ZN(new_n18718_));
  NOR2_X1    g18526(.A1(new_n18718_), .A2(new_n18712_), .ZN(new_n18719_));
  AOI22_X1   g18527(.A1(new_n18713_), .A2(\asqrt[37] ), .B1(new_n18711_), .B2(new_n18704_), .ZN(new_n18720_));
  NOR4_X1    g18528(.A1(new_n18495_), .A2(\asqrt[38] ), .A3(new_n18107_), .A4(new_n18359_), .ZN(new_n18721_));
  AOI21_X1   g18529(.A1(new_n18714_), .A2(new_n18103_), .B(new_n4645_), .ZN(new_n18722_));
  NOR2_X1    g18530(.A1(new_n18721_), .A2(new_n18722_), .ZN(new_n18723_));
  NAND2_X1   g18531(.A1(new_n18723_), .A2(new_n4330_), .ZN(new_n18724_));
  INV_X1     g18532(.I(new_n18724_), .ZN(new_n18725_));
  OAI21_X1   g18533(.A1(new_n18720_), .A2(new_n4645_), .B(new_n18725_), .ZN(new_n18726_));
  NAND2_X1   g18534(.A1(new_n18726_), .A2(new_n18719_), .ZN(new_n18727_));
  OAI22_X1   g18535(.A1(new_n18720_), .A2(new_n4645_), .B1(new_n18718_), .B2(new_n18712_), .ZN(new_n18728_));
  NAND2_X1   g18536(.A1(new_n18119_), .A2(\asqrt[39] ), .ZN(new_n18729_));
  NOR4_X1    g18537(.A1(new_n18495_), .A2(\asqrt[39] ), .A3(new_n18114_), .A4(new_n18119_), .ZN(new_n18730_));
  XOR2_X1    g18538(.A1(new_n18730_), .A2(new_n18729_), .Z(new_n18731_));
  NAND2_X1   g18539(.A1(new_n18731_), .A2(new_n4018_), .ZN(new_n18732_));
  AOI21_X1   g18540(.A1(new_n18728_), .A2(\asqrt[39] ), .B(new_n18732_), .ZN(new_n18733_));
  NOR2_X1    g18541(.A1(new_n18733_), .A2(new_n18727_), .ZN(new_n18734_));
  AOI22_X1   g18542(.A1(new_n18728_), .A2(\asqrt[39] ), .B1(new_n18726_), .B2(new_n18719_), .ZN(new_n18735_));
  NOR4_X1    g18543(.A1(new_n18495_), .A2(\asqrt[40] ), .A3(new_n18122_), .A4(new_n18366_), .ZN(new_n18736_));
  AOI21_X1   g18544(.A1(new_n18729_), .A2(new_n18118_), .B(new_n4018_), .ZN(new_n18737_));
  NOR2_X1    g18545(.A1(new_n18736_), .A2(new_n18737_), .ZN(new_n18738_));
  NAND2_X1   g18546(.A1(new_n18738_), .A2(new_n3760_), .ZN(new_n18739_));
  INV_X1     g18547(.I(new_n18739_), .ZN(new_n18740_));
  OAI21_X1   g18548(.A1(new_n18735_), .A2(new_n4018_), .B(new_n18740_), .ZN(new_n18741_));
  NAND2_X1   g18549(.A1(new_n18741_), .A2(new_n18734_), .ZN(new_n18742_));
  OAI22_X1   g18550(.A1(new_n18735_), .A2(new_n4018_), .B1(new_n18733_), .B2(new_n18727_), .ZN(new_n18743_));
  NAND2_X1   g18551(.A1(new_n18134_), .A2(\asqrt[41] ), .ZN(new_n18744_));
  NOR4_X1    g18552(.A1(new_n18495_), .A2(\asqrt[41] ), .A3(new_n18129_), .A4(new_n18134_), .ZN(new_n18745_));
  XOR2_X1    g18553(.A1(new_n18745_), .A2(new_n18744_), .Z(new_n18746_));
  NAND2_X1   g18554(.A1(new_n18746_), .A2(new_n3481_), .ZN(new_n18747_));
  AOI21_X1   g18555(.A1(new_n18743_), .A2(\asqrt[41] ), .B(new_n18747_), .ZN(new_n18748_));
  NOR2_X1    g18556(.A1(new_n18748_), .A2(new_n18742_), .ZN(new_n18749_));
  AOI22_X1   g18557(.A1(new_n18743_), .A2(\asqrt[41] ), .B1(new_n18741_), .B2(new_n18734_), .ZN(new_n18750_));
  NAND2_X1   g18558(.A1(new_n18373_), .A2(\asqrt[42] ), .ZN(new_n18751_));
  NOR4_X1    g18559(.A1(new_n18495_), .A2(\asqrt[42] ), .A3(new_n18137_), .A4(new_n18373_), .ZN(new_n18752_));
  XOR2_X1    g18560(.A1(new_n18752_), .A2(new_n18751_), .Z(new_n18753_));
  NAND2_X1   g18561(.A1(new_n18753_), .A2(new_n3208_), .ZN(new_n18754_));
  INV_X1     g18562(.I(new_n18754_), .ZN(new_n18755_));
  OAI21_X1   g18563(.A1(new_n18750_), .A2(new_n3481_), .B(new_n18755_), .ZN(new_n18756_));
  NAND2_X1   g18564(.A1(new_n18756_), .A2(new_n18749_), .ZN(new_n18757_));
  OAI22_X1   g18565(.A1(new_n18750_), .A2(new_n3481_), .B1(new_n18748_), .B2(new_n18742_), .ZN(new_n18758_));
  NOR4_X1    g18566(.A1(new_n18495_), .A2(\asqrt[43] ), .A3(new_n18144_), .A4(new_n18149_), .ZN(new_n18759_));
  AOI21_X1   g18567(.A1(new_n18751_), .A2(new_n18372_), .B(new_n3208_), .ZN(new_n18760_));
  NOR2_X1    g18568(.A1(new_n18759_), .A2(new_n18760_), .ZN(new_n18761_));
  NAND2_X1   g18569(.A1(new_n18761_), .A2(new_n2941_), .ZN(new_n18762_));
  AOI21_X1   g18570(.A1(new_n18758_), .A2(\asqrt[43] ), .B(new_n18762_), .ZN(new_n18763_));
  NOR2_X1    g18571(.A1(new_n18763_), .A2(new_n18757_), .ZN(new_n18764_));
  AOI22_X1   g18572(.A1(new_n18758_), .A2(\asqrt[43] ), .B1(new_n18756_), .B2(new_n18749_), .ZN(new_n18765_));
  NAND2_X1   g18573(.A1(new_n18380_), .A2(\asqrt[44] ), .ZN(new_n18766_));
  NOR4_X1    g18574(.A1(new_n18495_), .A2(\asqrt[44] ), .A3(new_n18152_), .A4(new_n18380_), .ZN(new_n18767_));
  XOR2_X1    g18575(.A1(new_n18767_), .A2(new_n18766_), .Z(new_n18768_));
  NAND2_X1   g18576(.A1(new_n18768_), .A2(new_n2728_), .ZN(new_n18769_));
  INV_X1     g18577(.I(new_n18769_), .ZN(new_n18770_));
  OAI21_X1   g18578(.A1(new_n18765_), .A2(new_n2941_), .B(new_n18770_), .ZN(new_n18771_));
  NAND2_X1   g18579(.A1(new_n18771_), .A2(new_n18764_), .ZN(new_n18772_));
  OAI22_X1   g18580(.A1(new_n18765_), .A2(new_n2941_), .B1(new_n18763_), .B2(new_n18757_), .ZN(new_n18773_));
  NOR4_X1    g18581(.A1(new_n18495_), .A2(\asqrt[45] ), .A3(new_n18159_), .A4(new_n18164_), .ZN(new_n18774_));
  AOI21_X1   g18582(.A1(new_n18766_), .A2(new_n18379_), .B(new_n2728_), .ZN(new_n18775_));
  NOR2_X1    g18583(.A1(new_n18774_), .A2(new_n18775_), .ZN(new_n18776_));
  NAND2_X1   g18584(.A1(new_n18776_), .A2(new_n2488_), .ZN(new_n18777_));
  AOI21_X1   g18585(.A1(new_n18773_), .A2(\asqrt[45] ), .B(new_n18777_), .ZN(new_n18778_));
  NOR2_X1    g18586(.A1(new_n18778_), .A2(new_n18772_), .ZN(new_n18779_));
  AOI22_X1   g18587(.A1(new_n18773_), .A2(\asqrt[45] ), .B1(new_n18771_), .B2(new_n18764_), .ZN(new_n18780_));
  NAND2_X1   g18588(.A1(new_n18387_), .A2(\asqrt[46] ), .ZN(new_n18781_));
  NOR4_X1    g18589(.A1(new_n18495_), .A2(\asqrt[46] ), .A3(new_n18167_), .A4(new_n18387_), .ZN(new_n18782_));
  XOR2_X1    g18590(.A1(new_n18782_), .A2(new_n18781_), .Z(new_n18783_));
  NAND2_X1   g18591(.A1(new_n18783_), .A2(new_n2253_), .ZN(new_n18784_));
  INV_X1     g18592(.I(new_n18784_), .ZN(new_n18785_));
  OAI21_X1   g18593(.A1(new_n18780_), .A2(new_n2488_), .B(new_n18785_), .ZN(new_n18786_));
  NAND2_X1   g18594(.A1(new_n18786_), .A2(new_n18779_), .ZN(new_n18787_));
  OAI22_X1   g18595(.A1(new_n18780_), .A2(new_n2488_), .B1(new_n18778_), .B2(new_n18772_), .ZN(new_n18788_));
  NAND2_X1   g18596(.A1(new_n18179_), .A2(\asqrt[47] ), .ZN(new_n18789_));
  NOR4_X1    g18597(.A1(new_n18495_), .A2(\asqrt[47] ), .A3(new_n18174_), .A4(new_n18179_), .ZN(new_n18790_));
  XOR2_X1    g18598(.A1(new_n18790_), .A2(new_n18789_), .Z(new_n18791_));
  NAND2_X1   g18599(.A1(new_n18791_), .A2(new_n2046_), .ZN(new_n18792_));
  AOI21_X1   g18600(.A1(new_n18788_), .A2(\asqrt[47] ), .B(new_n18792_), .ZN(new_n18793_));
  NOR2_X1    g18601(.A1(new_n18793_), .A2(new_n18787_), .ZN(new_n18794_));
  AOI22_X1   g18602(.A1(new_n18788_), .A2(\asqrt[47] ), .B1(new_n18786_), .B2(new_n18779_), .ZN(new_n18795_));
  NOR4_X1    g18603(.A1(new_n18495_), .A2(\asqrt[48] ), .A3(new_n18182_), .A4(new_n18394_), .ZN(new_n18796_));
  AOI21_X1   g18604(.A1(new_n18789_), .A2(new_n18178_), .B(new_n2046_), .ZN(new_n18797_));
  NOR2_X1    g18605(.A1(new_n18796_), .A2(new_n18797_), .ZN(new_n18798_));
  NAND2_X1   g18606(.A1(new_n18798_), .A2(new_n1854_), .ZN(new_n18799_));
  INV_X1     g18607(.I(new_n18799_), .ZN(new_n18800_));
  OAI21_X1   g18608(.A1(new_n18795_), .A2(new_n2046_), .B(new_n18800_), .ZN(new_n18801_));
  NAND2_X1   g18609(.A1(new_n18801_), .A2(new_n18794_), .ZN(new_n18802_));
  OAI22_X1   g18610(.A1(new_n18795_), .A2(new_n2046_), .B1(new_n18793_), .B2(new_n18787_), .ZN(new_n18803_));
  NAND2_X1   g18611(.A1(new_n18194_), .A2(\asqrt[49] ), .ZN(new_n18804_));
  NOR4_X1    g18612(.A1(new_n18495_), .A2(\asqrt[49] ), .A3(new_n18189_), .A4(new_n18194_), .ZN(new_n18805_));
  XOR2_X1    g18613(.A1(new_n18805_), .A2(new_n18804_), .Z(new_n18806_));
  NAND2_X1   g18614(.A1(new_n18806_), .A2(new_n1595_), .ZN(new_n18807_));
  AOI21_X1   g18615(.A1(new_n18803_), .A2(\asqrt[49] ), .B(new_n18807_), .ZN(new_n18808_));
  NOR2_X1    g18616(.A1(new_n18808_), .A2(new_n18802_), .ZN(new_n18809_));
  AOI22_X1   g18617(.A1(new_n18803_), .A2(\asqrt[49] ), .B1(new_n18801_), .B2(new_n18794_), .ZN(new_n18810_));
  NOR4_X1    g18618(.A1(new_n18495_), .A2(\asqrt[50] ), .A3(new_n18197_), .A4(new_n18401_), .ZN(new_n18811_));
  AOI21_X1   g18619(.A1(new_n18804_), .A2(new_n18193_), .B(new_n1595_), .ZN(new_n18812_));
  NOR2_X1    g18620(.A1(new_n18811_), .A2(new_n18812_), .ZN(new_n18813_));
  NAND2_X1   g18621(.A1(new_n18813_), .A2(new_n1436_), .ZN(new_n18814_));
  INV_X1     g18622(.I(new_n18814_), .ZN(new_n18815_));
  OAI21_X1   g18623(.A1(new_n18810_), .A2(new_n1595_), .B(new_n18815_), .ZN(new_n18816_));
  NAND2_X1   g18624(.A1(new_n18816_), .A2(new_n18809_), .ZN(new_n18817_));
  OAI22_X1   g18625(.A1(new_n18810_), .A2(new_n1595_), .B1(new_n18808_), .B2(new_n18802_), .ZN(new_n18818_));
  NAND2_X1   g18626(.A1(new_n18209_), .A2(\asqrt[51] ), .ZN(new_n18819_));
  NOR4_X1    g18627(.A1(new_n18495_), .A2(\asqrt[51] ), .A3(new_n18204_), .A4(new_n18209_), .ZN(new_n18820_));
  XOR2_X1    g18628(.A1(new_n18820_), .A2(new_n18819_), .Z(new_n18821_));
  NAND2_X1   g18629(.A1(new_n18821_), .A2(new_n1260_), .ZN(new_n18822_));
  AOI21_X1   g18630(.A1(new_n18818_), .A2(\asqrt[51] ), .B(new_n18822_), .ZN(new_n18823_));
  NOR2_X1    g18631(.A1(new_n18823_), .A2(new_n18817_), .ZN(new_n18824_));
  AOI22_X1   g18632(.A1(new_n18818_), .A2(\asqrt[51] ), .B1(new_n18816_), .B2(new_n18809_), .ZN(new_n18825_));
  NAND2_X1   g18633(.A1(new_n18408_), .A2(\asqrt[52] ), .ZN(new_n18826_));
  NOR4_X1    g18634(.A1(new_n18495_), .A2(\asqrt[52] ), .A3(new_n18212_), .A4(new_n18408_), .ZN(new_n18827_));
  XOR2_X1    g18635(.A1(new_n18827_), .A2(new_n18826_), .Z(new_n18828_));
  NAND2_X1   g18636(.A1(new_n18828_), .A2(new_n1096_), .ZN(new_n18829_));
  INV_X1     g18637(.I(new_n18829_), .ZN(new_n18830_));
  OAI21_X1   g18638(.A1(new_n18825_), .A2(new_n1260_), .B(new_n18830_), .ZN(new_n18831_));
  NAND2_X1   g18639(.A1(new_n18831_), .A2(new_n18824_), .ZN(new_n18832_));
  OAI22_X1   g18640(.A1(new_n18825_), .A2(new_n1260_), .B1(new_n18823_), .B2(new_n18817_), .ZN(new_n18833_));
  NOR4_X1    g18641(.A1(new_n18495_), .A2(\asqrt[53] ), .A3(new_n18219_), .A4(new_n18224_), .ZN(new_n18834_));
  XOR2_X1    g18642(.A1(new_n18834_), .A2(new_n18254_), .Z(new_n18835_));
  NAND2_X1   g18643(.A1(new_n18835_), .A2(new_n970_), .ZN(new_n18836_));
  AOI21_X1   g18644(.A1(new_n18833_), .A2(\asqrt[53] ), .B(new_n18836_), .ZN(new_n18837_));
  NOR2_X1    g18645(.A1(new_n18837_), .A2(new_n18832_), .ZN(new_n18838_));
  AOI22_X1   g18646(.A1(new_n18833_), .A2(\asqrt[53] ), .B1(new_n18831_), .B2(new_n18824_), .ZN(new_n18839_));
  NOR4_X1    g18647(.A1(new_n18495_), .A2(\asqrt[54] ), .A3(new_n18227_), .A4(new_n18415_), .ZN(new_n18840_));
  XOR2_X1    g18648(.A1(new_n18840_), .A2(new_n18428_), .Z(new_n18841_));
  NAND2_X1   g18649(.A1(new_n18841_), .A2(new_n825_), .ZN(new_n18842_));
  INV_X1     g18650(.I(new_n18842_), .ZN(new_n18843_));
  OAI21_X1   g18651(.A1(new_n18839_), .A2(new_n970_), .B(new_n18843_), .ZN(new_n18844_));
  NAND2_X1   g18652(.A1(new_n18844_), .A2(new_n18838_), .ZN(new_n18845_));
  OAI22_X1   g18653(.A1(new_n18839_), .A2(new_n970_), .B1(new_n18837_), .B2(new_n18832_), .ZN(new_n18846_));
  NOR4_X1    g18654(.A1(new_n18495_), .A2(\asqrt[55] ), .A3(new_n18234_), .A4(new_n18239_), .ZN(new_n18847_));
  XOR2_X1    g18655(.A1(new_n18847_), .A2(new_n18256_), .Z(new_n18848_));
  NAND2_X1   g18656(.A1(new_n18848_), .A2(new_n724_), .ZN(new_n18849_));
  AOI21_X1   g18657(.A1(new_n18846_), .A2(\asqrt[55] ), .B(new_n18849_), .ZN(new_n18850_));
  NOR2_X1    g18658(.A1(new_n18850_), .A2(new_n18845_), .ZN(new_n18851_));
  AOI22_X1   g18659(.A1(new_n18846_), .A2(\asqrt[55] ), .B1(new_n18844_), .B2(new_n18838_), .ZN(new_n18852_));
  NOR4_X1    g18660(.A1(new_n18495_), .A2(\asqrt[56] ), .A3(new_n18242_), .A4(new_n18422_), .ZN(new_n18853_));
  XOR2_X1    g18661(.A1(new_n18853_), .A2(new_n18430_), .Z(new_n18854_));
  NAND2_X1   g18662(.A1(new_n18854_), .A2(new_n587_), .ZN(new_n18855_));
  INV_X1     g18663(.I(new_n18855_), .ZN(new_n18856_));
  OAI21_X1   g18664(.A1(new_n18852_), .A2(new_n724_), .B(new_n18856_), .ZN(new_n18857_));
  NAND2_X1   g18665(.A1(new_n18857_), .A2(new_n18851_), .ZN(new_n18858_));
  OAI22_X1   g18666(.A1(new_n18852_), .A2(new_n724_), .B1(new_n18850_), .B2(new_n18845_), .ZN(new_n18859_));
  NOR4_X1    g18667(.A1(new_n18495_), .A2(\asqrt[57] ), .A3(new_n18249_), .A4(new_n18264_), .ZN(new_n18860_));
  XOR2_X1    g18668(.A1(new_n18860_), .A2(new_n18258_), .Z(new_n18861_));
  NAND2_X1   g18669(.A1(new_n18861_), .A2(new_n504_), .ZN(new_n18862_));
  AOI21_X1   g18670(.A1(new_n18859_), .A2(\asqrt[57] ), .B(new_n18862_), .ZN(new_n18863_));
  NOR2_X1    g18671(.A1(new_n18863_), .A2(new_n18858_), .ZN(new_n18864_));
  AOI22_X1   g18672(.A1(new_n18859_), .A2(\asqrt[57] ), .B1(new_n18857_), .B2(new_n18851_), .ZN(new_n18865_));
  NOR4_X1    g18673(.A1(new_n18495_), .A2(\asqrt[58] ), .A3(new_n18260_), .A4(new_n18441_), .ZN(new_n18866_));
  XOR2_X1    g18674(.A1(new_n18866_), .A2(new_n18432_), .Z(new_n18867_));
  NAND2_X1   g18675(.A1(new_n18867_), .A2(new_n376_), .ZN(new_n18868_));
  INV_X1     g18676(.I(new_n18868_), .ZN(new_n18869_));
  OAI21_X1   g18677(.A1(new_n18865_), .A2(new_n504_), .B(new_n18869_), .ZN(new_n18870_));
  NAND2_X1   g18678(.A1(new_n18870_), .A2(new_n18864_), .ZN(new_n18871_));
  OAI22_X1   g18679(.A1(new_n18865_), .A2(new_n504_), .B1(new_n18863_), .B2(new_n18858_), .ZN(new_n18872_));
  NOR4_X1    g18680(.A1(new_n18495_), .A2(\asqrt[59] ), .A3(new_n18267_), .A4(new_n18433_), .ZN(new_n18873_));
  XOR2_X1    g18681(.A1(new_n18873_), .A2(new_n18273_), .Z(new_n18874_));
  NAND2_X1   g18682(.A1(new_n18874_), .A2(new_n275_), .ZN(new_n18875_));
  AOI21_X1   g18683(.A1(new_n18872_), .A2(\asqrt[59] ), .B(new_n18875_), .ZN(new_n18876_));
  NOR2_X1    g18684(.A1(new_n18876_), .A2(new_n18871_), .ZN(new_n18877_));
  AOI22_X1   g18685(.A1(new_n18872_), .A2(\asqrt[59] ), .B1(new_n18870_), .B2(new_n18864_), .ZN(new_n18878_));
  NOR4_X1    g18686(.A1(new_n18495_), .A2(\asqrt[60] ), .A3(new_n18275_), .A4(new_n18459_), .ZN(new_n18879_));
  XOR2_X1    g18687(.A1(new_n18879_), .A2(new_n18448_), .Z(new_n18880_));
  NAND2_X1   g18688(.A1(new_n18880_), .A2(new_n229_), .ZN(new_n18881_));
  INV_X1     g18689(.I(new_n18881_), .ZN(new_n18882_));
  OAI21_X1   g18690(.A1(new_n18878_), .A2(new_n275_), .B(new_n18882_), .ZN(new_n18883_));
  OAI22_X1   g18691(.A1(new_n18878_), .A2(new_n275_), .B1(new_n18876_), .B2(new_n18871_), .ZN(new_n18884_));
  AOI22_X1   g18692(.A1(new_n18884_), .A2(\asqrt[61] ), .B1(new_n18883_), .B2(new_n18877_), .ZN(new_n18885_));
  NOR2_X1    g18693(.A1(new_n18885_), .A2(new_n196_), .ZN(new_n18886_));
  NAND3_X1   g18694(.A1(new_n18489_), .A2(new_n17858_), .A3(new_n18469_), .ZN(new_n18887_));
  INV_X1     g18695(.I(new_n18887_), .ZN(new_n18888_));
  NOR2_X1    g18696(.A1(new_n18499_), .A2(new_n196_), .ZN(new_n18889_));
  INV_X1     g18697(.I(new_n18482_), .ZN(new_n18890_));
  NAND3_X1   g18698(.A1(\asqrt[9] ), .A2(new_n18889_), .A3(new_n18890_), .ZN(new_n18891_));
  OAI21_X1   g18699(.A1(new_n18462_), .A2(\asqrt[62] ), .B(new_n17865_), .ZN(new_n18892_));
  OAI21_X1   g18700(.A1(\asqrt[9] ), .A2(new_n18892_), .B(new_n18889_), .ZN(new_n18893_));
  NAND2_X1   g18701(.A1(new_n18893_), .A2(new_n18891_), .ZN(new_n18894_));
  NOR3_X1    g18702(.A1(new_n18498_), .A2(\asqrt[61] ), .A3(new_n18436_), .ZN(new_n18895_));
  NAND2_X1   g18703(.A1(\asqrt[9] ), .A2(new_n18895_), .ZN(new_n18896_));
  XOR2_X1    g18704(.A1(new_n18896_), .A2(new_n18449_), .Z(new_n18897_));
  NOR2_X1    g18705(.A1(new_n18897_), .A2(new_n196_), .ZN(new_n18898_));
  INV_X1     g18706(.I(new_n18471_), .ZN(new_n18899_));
  AOI21_X1   g18707(.A1(new_n18485_), .A2(new_n18899_), .B(new_n18473_), .ZN(new_n18900_));
  NOR3_X1    g18708(.A1(new_n18470_), .A2(new_n17656_), .A3(new_n17667_), .ZN(new_n18901_));
  NOR2_X1    g18709(.A1(new_n18901_), .A2(new_n18900_), .ZN(new_n18902_));
  NOR3_X1    g18710(.A1(new_n18511_), .A2(new_n17870_), .A3(\asqrt[9] ), .ZN(new_n18903_));
  AOI21_X1   g18711(.A1(new_n18504_), .A2(new_n17869_), .B(new_n18495_), .ZN(new_n18904_));
  NOR4_X1    g18712(.A1(new_n18904_), .A2(new_n18903_), .A3(\asqrt[11] ), .A4(new_n18493_), .ZN(new_n18905_));
  NOR2_X1    g18713(.A1(new_n18905_), .A2(new_n18902_), .ZN(new_n18906_));
  NOR3_X1    g18714(.A1(new_n18901_), .A2(new_n18900_), .A3(new_n18493_), .ZN(new_n18907_));
  NOR3_X1    g18715(.A1(new_n18495_), .A2(new_n17891_), .A3(new_n18519_), .ZN(new_n18908_));
  AOI21_X1   g18716(.A1(\asqrt[9] ), .A2(new_n18520_), .B(new_n17892_), .ZN(new_n18909_));
  NOR3_X1    g18717(.A1(new_n18909_), .A2(new_n18908_), .A3(\asqrt[12] ), .ZN(new_n18910_));
  OAI21_X1   g18718(.A1(new_n18907_), .A2(new_n17271_), .B(new_n18910_), .ZN(new_n18911_));
  NAND2_X1   g18719(.A1(new_n18906_), .A2(new_n18911_), .ZN(new_n18912_));
  OAI22_X1   g18720(.A1(new_n18905_), .A2(new_n18902_), .B1(new_n17271_), .B2(new_n18907_), .ZN(new_n18913_));
  INV_X1     g18721(.I(new_n18534_), .ZN(new_n18914_));
  AOI21_X1   g18722(.A1(new_n18913_), .A2(\asqrt[12] ), .B(new_n18914_), .ZN(new_n18915_));
  NOR2_X1    g18723(.A1(new_n18915_), .A2(new_n18912_), .ZN(new_n18916_));
  AOI22_X1   g18724(.A1(new_n18913_), .A2(\asqrt[12] ), .B1(new_n18906_), .B2(new_n18911_), .ZN(new_n18917_));
  INV_X1     g18725(.I(new_n18541_), .ZN(new_n18918_));
  OAI21_X1   g18726(.A1(new_n18917_), .A2(new_n16060_), .B(new_n18918_), .ZN(new_n18919_));
  NAND2_X1   g18727(.A1(new_n18919_), .A2(new_n18916_), .ZN(new_n18920_));
  OAI22_X1   g18728(.A1(new_n18917_), .A2(new_n16060_), .B1(new_n18915_), .B2(new_n18912_), .ZN(new_n18921_));
  AOI21_X1   g18729(.A1(new_n18921_), .A2(\asqrt[14] ), .B(new_n18547_), .ZN(new_n18922_));
  NOR2_X1    g18730(.A1(new_n18922_), .A2(new_n18920_), .ZN(new_n18923_));
  AOI22_X1   g18731(.A1(new_n18921_), .A2(\asqrt[14] ), .B1(new_n18919_), .B2(new_n18916_), .ZN(new_n18924_));
  INV_X1     g18732(.I(new_n18555_), .ZN(new_n18925_));
  OAI21_X1   g18733(.A1(new_n18924_), .A2(new_n14871_), .B(new_n18925_), .ZN(new_n18926_));
  NAND2_X1   g18734(.A1(new_n18926_), .A2(new_n18923_), .ZN(new_n18927_));
  OAI22_X1   g18735(.A1(new_n18924_), .A2(new_n14871_), .B1(new_n18922_), .B2(new_n18920_), .ZN(new_n18928_));
  AOI21_X1   g18736(.A1(new_n18928_), .A2(\asqrt[16] ), .B(new_n18561_), .ZN(new_n18929_));
  NOR2_X1    g18737(.A1(new_n18929_), .A2(new_n18927_), .ZN(new_n18930_));
  AOI22_X1   g18738(.A1(new_n18928_), .A2(\asqrt[16] ), .B1(new_n18926_), .B2(new_n18923_), .ZN(new_n18931_));
  INV_X1     g18739(.I(new_n18568_), .ZN(new_n18932_));
  OAI21_X1   g18740(.A1(new_n18931_), .A2(new_n13760_), .B(new_n18932_), .ZN(new_n18933_));
  NAND2_X1   g18741(.A1(new_n18933_), .A2(new_n18930_), .ZN(new_n18934_));
  OAI22_X1   g18742(.A1(new_n18931_), .A2(new_n13760_), .B1(new_n18929_), .B2(new_n18927_), .ZN(new_n18935_));
  AOI21_X1   g18743(.A1(new_n18935_), .A2(\asqrt[18] ), .B(new_n18574_), .ZN(new_n18936_));
  NOR2_X1    g18744(.A1(new_n18936_), .A2(new_n18934_), .ZN(new_n18937_));
  AOI22_X1   g18745(.A1(new_n18935_), .A2(\asqrt[18] ), .B1(new_n18933_), .B2(new_n18930_), .ZN(new_n18938_));
  INV_X1     g18746(.I(new_n18582_), .ZN(new_n18939_));
  OAI21_X1   g18747(.A1(new_n18938_), .A2(new_n12657_), .B(new_n18939_), .ZN(new_n18940_));
  NAND2_X1   g18748(.A1(new_n18940_), .A2(new_n18937_), .ZN(new_n18941_));
  OAI22_X1   g18749(.A1(new_n18938_), .A2(new_n12657_), .B1(new_n18936_), .B2(new_n18934_), .ZN(new_n18942_));
  AOI21_X1   g18750(.A1(new_n18942_), .A2(\asqrt[20] ), .B(new_n18589_), .ZN(new_n18943_));
  NOR2_X1    g18751(.A1(new_n18943_), .A2(new_n18941_), .ZN(new_n18944_));
  AOI22_X1   g18752(.A1(new_n18942_), .A2(\asqrt[20] ), .B1(new_n18940_), .B2(new_n18937_), .ZN(new_n18945_));
  INV_X1     g18753(.I(new_n18597_), .ZN(new_n18946_));
  OAI21_X1   g18754(.A1(new_n18945_), .A2(new_n11631_), .B(new_n18946_), .ZN(new_n18947_));
  NAND2_X1   g18755(.A1(new_n18947_), .A2(new_n18944_), .ZN(new_n18948_));
  OAI22_X1   g18756(.A1(new_n18945_), .A2(new_n11631_), .B1(new_n18943_), .B2(new_n18941_), .ZN(new_n18949_));
  AOI21_X1   g18757(.A1(new_n18949_), .A2(\asqrt[22] ), .B(new_n18604_), .ZN(new_n18950_));
  NOR2_X1    g18758(.A1(new_n18950_), .A2(new_n18948_), .ZN(new_n18951_));
  AOI22_X1   g18759(.A1(new_n18949_), .A2(\asqrt[22] ), .B1(new_n18947_), .B2(new_n18944_), .ZN(new_n18952_));
  INV_X1     g18760(.I(new_n18612_), .ZN(new_n18953_));
  OAI21_X1   g18761(.A1(new_n18952_), .A2(new_n10614_), .B(new_n18953_), .ZN(new_n18954_));
  NAND2_X1   g18762(.A1(new_n18954_), .A2(new_n18951_), .ZN(new_n18955_));
  OAI22_X1   g18763(.A1(new_n18952_), .A2(new_n10614_), .B1(new_n18950_), .B2(new_n18948_), .ZN(new_n18956_));
  AOI21_X1   g18764(.A1(new_n18956_), .A2(\asqrt[24] ), .B(new_n18619_), .ZN(new_n18957_));
  NOR2_X1    g18765(.A1(new_n18957_), .A2(new_n18955_), .ZN(new_n18958_));
  AOI22_X1   g18766(.A1(new_n18956_), .A2(\asqrt[24] ), .B1(new_n18954_), .B2(new_n18951_), .ZN(new_n18959_));
  INV_X1     g18767(.I(new_n18627_), .ZN(new_n18960_));
  OAI21_X1   g18768(.A1(new_n18959_), .A2(new_n9672_), .B(new_n18960_), .ZN(new_n18961_));
  NAND2_X1   g18769(.A1(new_n18961_), .A2(new_n18958_), .ZN(new_n18962_));
  OAI22_X1   g18770(.A1(new_n18959_), .A2(new_n9672_), .B1(new_n18957_), .B2(new_n18955_), .ZN(new_n18963_));
  AOI21_X1   g18771(.A1(new_n18963_), .A2(\asqrt[26] ), .B(new_n18634_), .ZN(new_n18964_));
  NOR2_X1    g18772(.A1(new_n18964_), .A2(new_n18962_), .ZN(new_n18965_));
  AOI22_X1   g18773(.A1(new_n18963_), .A2(\asqrt[26] ), .B1(new_n18961_), .B2(new_n18958_), .ZN(new_n18966_));
  INV_X1     g18774(.I(new_n18642_), .ZN(new_n18967_));
  OAI21_X1   g18775(.A1(new_n18966_), .A2(new_n8763_), .B(new_n18967_), .ZN(new_n18968_));
  NAND2_X1   g18776(.A1(new_n18968_), .A2(new_n18965_), .ZN(new_n18969_));
  OAI22_X1   g18777(.A1(new_n18966_), .A2(new_n8763_), .B1(new_n18964_), .B2(new_n18962_), .ZN(new_n18970_));
  AOI21_X1   g18778(.A1(new_n18970_), .A2(\asqrt[28] ), .B(new_n18649_), .ZN(new_n18971_));
  NOR2_X1    g18779(.A1(new_n18971_), .A2(new_n18969_), .ZN(new_n18972_));
  AOI22_X1   g18780(.A1(new_n18970_), .A2(\asqrt[28] ), .B1(new_n18968_), .B2(new_n18965_), .ZN(new_n18973_));
  INV_X1     g18781(.I(new_n18657_), .ZN(new_n18974_));
  OAI21_X1   g18782(.A1(new_n18973_), .A2(new_n7931_), .B(new_n18974_), .ZN(new_n18975_));
  NAND2_X1   g18783(.A1(new_n18975_), .A2(new_n18972_), .ZN(new_n18976_));
  OAI22_X1   g18784(.A1(new_n18973_), .A2(new_n7931_), .B1(new_n18971_), .B2(new_n18969_), .ZN(new_n18977_));
  AOI21_X1   g18785(.A1(new_n18977_), .A2(\asqrt[30] ), .B(new_n18664_), .ZN(new_n18978_));
  NOR2_X1    g18786(.A1(new_n18978_), .A2(new_n18976_), .ZN(new_n18979_));
  AOI22_X1   g18787(.A1(new_n18977_), .A2(\asqrt[30] ), .B1(new_n18975_), .B2(new_n18972_), .ZN(new_n18980_));
  INV_X1     g18788(.I(new_n18672_), .ZN(new_n18981_));
  OAI21_X1   g18789(.A1(new_n18980_), .A2(new_n7110_), .B(new_n18981_), .ZN(new_n18982_));
  NAND2_X1   g18790(.A1(new_n18982_), .A2(new_n18979_), .ZN(new_n18983_));
  OAI22_X1   g18791(.A1(new_n18980_), .A2(new_n7110_), .B1(new_n18978_), .B2(new_n18976_), .ZN(new_n18984_));
  AOI21_X1   g18792(.A1(new_n18984_), .A2(\asqrt[32] ), .B(new_n18679_), .ZN(new_n18985_));
  NOR2_X1    g18793(.A1(new_n18985_), .A2(new_n18983_), .ZN(new_n18986_));
  AOI22_X1   g18794(.A1(new_n18984_), .A2(\asqrt[32] ), .B1(new_n18982_), .B2(new_n18979_), .ZN(new_n18987_));
  INV_X1     g18795(.I(new_n18687_), .ZN(new_n18988_));
  OAI21_X1   g18796(.A1(new_n18987_), .A2(new_n6365_), .B(new_n18988_), .ZN(new_n18989_));
  NAND2_X1   g18797(.A1(new_n18989_), .A2(new_n18986_), .ZN(new_n18990_));
  OAI22_X1   g18798(.A1(new_n18987_), .A2(new_n6365_), .B1(new_n18985_), .B2(new_n18983_), .ZN(new_n18991_));
  AOI21_X1   g18799(.A1(new_n18991_), .A2(\asqrt[34] ), .B(new_n18694_), .ZN(new_n18992_));
  NOR2_X1    g18800(.A1(new_n18992_), .A2(new_n18990_), .ZN(new_n18993_));
  AOI22_X1   g18801(.A1(new_n18991_), .A2(\asqrt[34] ), .B1(new_n18989_), .B2(new_n18986_), .ZN(new_n18994_));
  INV_X1     g18802(.I(new_n18702_), .ZN(new_n18995_));
  OAI21_X1   g18803(.A1(new_n18994_), .A2(new_n5626_), .B(new_n18995_), .ZN(new_n18996_));
  NAND2_X1   g18804(.A1(new_n18996_), .A2(new_n18993_), .ZN(new_n18997_));
  OAI22_X1   g18805(.A1(new_n18994_), .A2(new_n5626_), .B1(new_n18992_), .B2(new_n18990_), .ZN(new_n18998_));
  AOI21_X1   g18806(.A1(new_n18998_), .A2(\asqrt[36] ), .B(new_n18709_), .ZN(new_n18999_));
  NOR2_X1    g18807(.A1(new_n18999_), .A2(new_n18997_), .ZN(new_n19000_));
  AOI22_X1   g18808(.A1(new_n18998_), .A2(\asqrt[36] ), .B1(new_n18996_), .B2(new_n18993_), .ZN(new_n19001_));
  INV_X1     g18809(.I(new_n18717_), .ZN(new_n19002_));
  OAI21_X1   g18810(.A1(new_n19001_), .A2(new_n4973_), .B(new_n19002_), .ZN(new_n19003_));
  NAND2_X1   g18811(.A1(new_n19003_), .A2(new_n19000_), .ZN(new_n19004_));
  OAI22_X1   g18812(.A1(new_n19001_), .A2(new_n4973_), .B1(new_n18999_), .B2(new_n18997_), .ZN(new_n19005_));
  AOI21_X1   g18813(.A1(new_n19005_), .A2(\asqrt[38] ), .B(new_n18724_), .ZN(new_n19006_));
  NOR2_X1    g18814(.A1(new_n19006_), .A2(new_n19004_), .ZN(new_n19007_));
  AOI22_X1   g18815(.A1(new_n19005_), .A2(\asqrt[38] ), .B1(new_n19003_), .B2(new_n19000_), .ZN(new_n19008_));
  INV_X1     g18816(.I(new_n18732_), .ZN(new_n19009_));
  OAI21_X1   g18817(.A1(new_n19008_), .A2(new_n4330_), .B(new_n19009_), .ZN(new_n19010_));
  NAND2_X1   g18818(.A1(new_n19010_), .A2(new_n19007_), .ZN(new_n19011_));
  OAI22_X1   g18819(.A1(new_n19008_), .A2(new_n4330_), .B1(new_n19006_), .B2(new_n19004_), .ZN(new_n19012_));
  AOI21_X1   g18820(.A1(new_n19012_), .A2(\asqrt[40] ), .B(new_n18739_), .ZN(new_n19013_));
  NOR2_X1    g18821(.A1(new_n19013_), .A2(new_n19011_), .ZN(new_n19014_));
  AOI22_X1   g18822(.A1(new_n19012_), .A2(\asqrt[40] ), .B1(new_n19010_), .B2(new_n19007_), .ZN(new_n19015_));
  INV_X1     g18823(.I(new_n18747_), .ZN(new_n19016_));
  OAI21_X1   g18824(.A1(new_n19015_), .A2(new_n3760_), .B(new_n19016_), .ZN(new_n19017_));
  NAND2_X1   g18825(.A1(new_n19017_), .A2(new_n19014_), .ZN(new_n19018_));
  OAI22_X1   g18826(.A1(new_n19015_), .A2(new_n3760_), .B1(new_n19013_), .B2(new_n19011_), .ZN(new_n19019_));
  AOI21_X1   g18827(.A1(new_n19019_), .A2(\asqrt[42] ), .B(new_n18754_), .ZN(new_n19020_));
  NOR2_X1    g18828(.A1(new_n19020_), .A2(new_n19018_), .ZN(new_n19021_));
  AOI22_X1   g18829(.A1(new_n19019_), .A2(\asqrt[42] ), .B1(new_n19017_), .B2(new_n19014_), .ZN(new_n19022_));
  INV_X1     g18830(.I(new_n18762_), .ZN(new_n19023_));
  OAI21_X1   g18831(.A1(new_n19022_), .A2(new_n3208_), .B(new_n19023_), .ZN(new_n19024_));
  NAND2_X1   g18832(.A1(new_n19024_), .A2(new_n19021_), .ZN(new_n19025_));
  OAI22_X1   g18833(.A1(new_n19022_), .A2(new_n3208_), .B1(new_n19020_), .B2(new_n19018_), .ZN(new_n19026_));
  AOI21_X1   g18834(.A1(new_n19026_), .A2(\asqrt[44] ), .B(new_n18769_), .ZN(new_n19027_));
  NOR2_X1    g18835(.A1(new_n19027_), .A2(new_n19025_), .ZN(new_n19028_));
  AOI22_X1   g18836(.A1(new_n19026_), .A2(\asqrt[44] ), .B1(new_n19024_), .B2(new_n19021_), .ZN(new_n19029_));
  INV_X1     g18837(.I(new_n18777_), .ZN(new_n19030_));
  OAI21_X1   g18838(.A1(new_n19029_), .A2(new_n2728_), .B(new_n19030_), .ZN(new_n19031_));
  NAND2_X1   g18839(.A1(new_n19031_), .A2(new_n19028_), .ZN(new_n19032_));
  OAI22_X1   g18840(.A1(new_n19029_), .A2(new_n2728_), .B1(new_n19027_), .B2(new_n19025_), .ZN(new_n19033_));
  AOI21_X1   g18841(.A1(new_n19033_), .A2(\asqrt[46] ), .B(new_n18784_), .ZN(new_n19034_));
  NOR2_X1    g18842(.A1(new_n19034_), .A2(new_n19032_), .ZN(new_n19035_));
  AOI22_X1   g18843(.A1(new_n19033_), .A2(\asqrt[46] ), .B1(new_n19031_), .B2(new_n19028_), .ZN(new_n19036_));
  INV_X1     g18844(.I(new_n18792_), .ZN(new_n19037_));
  OAI21_X1   g18845(.A1(new_n19036_), .A2(new_n2253_), .B(new_n19037_), .ZN(new_n19038_));
  NAND2_X1   g18846(.A1(new_n19038_), .A2(new_n19035_), .ZN(new_n19039_));
  OAI22_X1   g18847(.A1(new_n19036_), .A2(new_n2253_), .B1(new_n19034_), .B2(new_n19032_), .ZN(new_n19040_));
  AOI21_X1   g18848(.A1(new_n19040_), .A2(\asqrt[48] ), .B(new_n18799_), .ZN(new_n19041_));
  NOR2_X1    g18849(.A1(new_n19041_), .A2(new_n19039_), .ZN(new_n19042_));
  AOI22_X1   g18850(.A1(new_n19040_), .A2(\asqrt[48] ), .B1(new_n19038_), .B2(new_n19035_), .ZN(new_n19043_));
  INV_X1     g18851(.I(new_n18807_), .ZN(new_n19044_));
  OAI21_X1   g18852(.A1(new_n19043_), .A2(new_n1854_), .B(new_n19044_), .ZN(new_n19045_));
  NAND2_X1   g18853(.A1(new_n19045_), .A2(new_n19042_), .ZN(new_n19046_));
  OAI22_X1   g18854(.A1(new_n19043_), .A2(new_n1854_), .B1(new_n19041_), .B2(new_n19039_), .ZN(new_n19047_));
  AOI21_X1   g18855(.A1(new_n19047_), .A2(\asqrt[50] ), .B(new_n18814_), .ZN(new_n19048_));
  NOR2_X1    g18856(.A1(new_n19048_), .A2(new_n19046_), .ZN(new_n19049_));
  AOI22_X1   g18857(.A1(new_n19047_), .A2(\asqrt[50] ), .B1(new_n19045_), .B2(new_n19042_), .ZN(new_n19050_));
  INV_X1     g18858(.I(new_n18822_), .ZN(new_n19051_));
  OAI21_X1   g18859(.A1(new_n19050_), .A2(new_n1436_), .B(new_n19051_), .ZN(new_n19052_));
  NAND2_X1   g18860(.A1(new_n19052_), .A2(new_n19049_), .ZN(new_n19053_));
  OAI22_X1   g18861(.A1(new_n19050_), .A2(new_n1436_), .B1(new_n19048_), .B2(new_n19046_), .ZN(new_n19054_));
  AOI21_X1   g18862(.A1(new_n19054_), .A2(\asqrt[52] ), .B(new_n18829_), .ZN(new_n19055_));
  NOR2_X1    g18863(.A1(new_n19055_), .A2(new_n19053_), .ZN(new_n19056_));
  AOI22_X1   g18864(.A1(new_n19054_), .A2(\asqrt[52] ), .B1(new_n19052_), .B2(new_n19049_), .ZN(new_n19057_));
  INV_X1     g18865(.I(new_n18836_), .ZN(new_n19058_));
  OAI21_X1   g18866(.A1(new_n19057_), .A2(new_n1096_), .B(new_n19058_), .ZN(new_n19059_));
  NAND2_X1   g18867(.A1(new_n19059_), .A2(new_n19056_), .ZN(new_n19060_));
  OAI22_X1   g18868(.A1(new_n19057_), .A2(new_n1096_), .B1(new_n19055_), .B2(new_n19053_), .ZN(new_n19061_));
  AOI21_X1   g18869(.A1(new_n19061_), .A2(\asqrt[54] ), .B(new_n18842_), .ZN(new_n19062_));
  NOR2_X1    g18870(.A1(new_n19062_), .A2(new_n19060_), .ZN(new_n19063_));
  AOI22_X1   g18871(.A1(new_n19061_), .A2(\asqrt[54] ), .B1(new_n19059_), .B2(new_n19056_), .ZN(new_n19064_));
  INV_X1     g18872(.I(new_n18849_), .ZN(new_n19065_));
  OAI21_X1   g18873(.A1(new_n19064_), .A2(new_n825_), .B(new_n19065_), .ZN(new_n19066_));
  NAND2_X1   g18874(.A1(new_n19066_), .A2(new_n19063_), .ZN(new_n19067_));
  OAI22_X1   g18875(.A1(new_n19064_), .A2(new_n825_), .B1(new_n19062_), .B2(new_n19060_), .ZN(new_n19068_));
  AOI21_X1   g18876(.A1(new_n19068_), .A2(\asqrt[56] ), .B(new_n18855_), .ZN(new_n19069_));
  NOR2_X1    g18877(.A1(new_n19069_), .A2(new_n19067_), .ZN(new_n19070_));
  AOI22_X1   g18878(.A1(new_n19068_), .A2(\asqrt[56] ), .B1(new_n19066_), .B2(new_n19063_), .ZN(new_n19071_));
  INV_X1     g18879(.I(new_n18862_), .ZN(new_n19072_));
  OAI21_X1   g18880(.A1(new_n19071_), .A2(new_n587_), .B(new_n19072_), .ZN(new_n19073_));
  NAND2_X1   g18881(.A1(new_n19073_), .A2(new_n19070_), .ZN(new_n19074_));
  OAI22_X1   g18882(.A1(new_n19071_), .A2(new_n587_), .B1(new_n19069_), .B2(new_n19067_), .ZN(new_n19075_));
  AOI21_X1   g18883(.A1(new_n19075_), .A2(\asqrt[58] ), .B(new_n18868_), .ZN(new_n19076_));
  NOR2_X1    g18884(.A1(new_n19076_), .A2(new_n19074_), .ZN(new_n19077_));
  AOI22_X1   g18885(.A1(new_n19075_), .A2(\asqrt[58] ), .B1(new_n19073_), .B2(new_n19070_), .ZN(new_n19078_));
  INV_X1     g18886(.I(new_n18875_), .ZN(new_n19079_));
  OAI21_X1   g18887(.A1(new_n19078_), .A2(new_n376_), .B(new_n19079_), .ZN(new_n19080_));
  NAND2_X1   g18888(.A1(new_n19080_), .A2(new_n19077_), .ZN(new_n19081_));
  OAI22_X1   g18889(.A1(new_n19078_), .A2(new_n376_), .B1(new_n19076_), .B2(new_n19074_), .ZN(new_n19082_));
  AOI21_X1   g18890(.A1(new_n19082_), .A2(\asqrt[60] ), .B(new_n18881_), .ZN(new_n19083_));
  NOR2_X1    g18891(.A1(new_n19083_), .A2(new_n19081_), .ZN(new_n19084_));
  AOI22_X1   g18892(.A1(new_n19082_), .A2(\asqrt[60] ), .B1(new_n19080_), .B2(new_n19077_), .ZN(new_n19085_));
  INV_X1     g18893(.I(new_n18897_), .ZN(new_n19086_));
  NOR2_X1    g18894(.A1(new_n19086_), .A2(\asqrt[62] ), .ZN(new_n19087_));
  NOR3_X1    g18895(.A1(new_n19085_), .A2(new_n229_), .A3(new_n19087_), .ZN(new_n19088_));
  AOI21_X1   g18896(.A1(new_n19088_), .A2(new_n19084_), .B(new_n18898_), .ZN(new_n19089_));
  NAND3_X1   g18897(.A1(new_n18495_), .A2(new_n17857_), .A3(new_n18500_), .ZN(new_n19090_));
  AOI21_X1   g18898(.A1(new_n19090_), .A2(new_n18454_), .B(\asqrt[63] ), .ZN(new_n19091_));
  AOI21_X1   g18899(.A1(new_n19089_), .A2(new_n19091_), .B(new_n18894_), .ZN(new_n19092_));
  INV_X1     g18900(.I(new_n18894_), .ZN(new_n19093_));
  NAND4_X1   g18901(.A1(new_n18885_), .A2(new_n196_), .A3(new_n19093_), .A4(new_n19086_), .ZN(new_n19094_));
  NAND2_X1   g18902(.A1(new_n18476_), .A2(new_n17857_), .ZN(new_n19095_));
  XOR2_X1    g18903(.A1(new_n18476_), .A2(\asqrt[63] ), .Z(new_n19096_));
  AOI21_X1   g18904(.A1(\asqrt[9] ), .A2(new_n19095_), .B(new_n19096_), .ZN(new_n19097_));
  INV_X1     g18905(.I(new_n19097_), .ZN(new_n19098_));
  NOR2_X1    g18906(.A1(new_n19094_), .A2(new_n19098_), .ZN(new_n19099_));
  NAND3_X1   g18907(.A1(new_n19099_), .A2(new_n19092_), .A3(new_n18888_), .ZN(new_n19100_));
  OAI22_X1   g18908(.A1(new_n19085_), .A2(new_n229_), .B1(new_n19083_), .B2(new_n19081_), .ZN(new_n19101_));
  NOR2_X1    g18909(.A1(new_n19101_), .A2(\asqrt[62] ), .ZN(new_n19102_));
  NAND3_X1   g18910(.A1(new_n19102_), .A2(new_n18886_), .A3(new_n19086_), .ZN(new_n19103_));
  NOR2_X1    g18911(.A1(new_n19100_), .A2(new_n19103_), .ZN(new_n19104_));
  INV_X1     g18912(.I(new_n18898_), .ZN(new_n19105_));
  NAND2_X1   g18913(.A1(new_n18883_), .A2(new_n18877_), .ZN(new_n19106_));
  INV_X1     g18914(.I(new_n19087_), .ZN(new_n19107_));
  NAND3_X1   g18915(.A1(new_n18884_), .A2(\asqrt[61] ), .A3(new_n19107_), .ZN(new_n19108_));
  OAI21_X1   g18916(.A1(new_n19108_), .A2(new_n19106_), .B(new_n19105_), .ZN(new_n19109_));
  INV_X1     g18917(.I(new_n19091_), .ZN(new_n19110_));
  OAI21_X1   g18918(.A1(new_n19109_), .A2(new_n19110_), .B(new_n19093_), .ZN(new_n19111_));
  NOR4_X1    g18919(.A1(new_n19111_), .A2(new_n18887_), .A3(new_n19094_), .A4(new_n19098_), .ZN(\asqrt[8] ));
  OR3_X2     g18920(.A1(\asqrt[8] ), .A2(new_n19086_), .A3(new_n19102_), .Z(new_n19113_));
  AOI21_X1   g18921(.A1(new_n19113_), .A2(new_n18886_), .B(new_n19104_), .ZN(new_n19114_));
  INV_X1     g18922(.I(new_n19114_), .ZN(new_n19115_));
  INV_X1     g18923(.I(\a[16] ), .ZN(new_n19116_));
  NOR2_X1    g18924(.A1(\a[14] ), .A2(\a[15] ), .ZN(new_n19117_));
  INV_X1     g18925(.I(new_n19117_), .ZN(new_n19118_));
  NOR3_X1    g18926(.A1(new_n18502_), .A2(new_n19116_), .A3(new_n19118_), .ZN(new_n19119_));
  NAND2_X1   g18927(.A1(new_n18509_), .A2(new_n19119_), .ZN(new_n19120_));
  XOR2_X1    g18928(.A1(new_n19120_), .A2(\a[17] ), .Z(new_n19121_));
  INV_X1     g18929(.I(\a[17] ), .ZN(new_n19122_));
  NOR4_X1    g18930(.A1(new_n19101_), .A2(\asqrt[62] ), .A3(new_n18894_), .A4(new_n18897_), .ZN(new_n19123_));
  NAND2_X1   g18931(.A1(new_n19123_), .A2(new_n19097_), .ZN(new_n19124_));
  NOR4_X1    g18932(.A1(new_n19124_), .A2(new_n19122_), .A3(new_n19111_), .A4(new_n18887_), .ZN(new_n19125_));
  NOR2_X1    g18933(.A1(new_n19122_), .A2(\a[16] ), .ZN(new_n19126_));
  OAI21_X1   g18934(.A1(new_n19125_), .A2(new_n19126_), .B(new_n19121_), .ZN(new_n19127_));
  INV_X1     g18935(.I(new_n19121_), .ZN(new_n19128_));
  NAND4_X1   g18936(.A1(new_n19099_), .A2(new_n19092_), .A3(\a[17] ), .A4(new_n18888_), .ZN(new_n19129_));
  NAND3_X1   g18937(.A1(new_n19129_), .A2(\a[16] ), .A3(new_n19128_), .ZN(new_n19130_));
  NAND2_X1   g18938(.A1(new_n19127_), .A2(new_n19130_), .ZN(new_n19131_));
  NOR2_X1    g18939(.A1(new_n19124_), .A2(new_n19111_), .ZN(new_n19132_));
  NOR4_X1    g18940(.A1(new_n18468_), .A2(new_n17857_), .A3(new_n18497_), .A4(new_n18469_), .ZN(new_n19133_));
  NAND2_X1   g18941(.A1(\asqrt[9] ), .A2(\a[16] ), .ZN(new_n19134_));
  XOR2_X1    g18942(.A1(new_n19134_), .A2(new_n19133_), .Z(new_n19135_));
  NOR2_X1    g18943(.A1(new_n19135_), .A2(new_n19118_), .ZN(new_n19136_));
  INV_X1     g18944(.I(new_n19136_), .ZN(new_n19137_));
  NAND2_X1   g18945(.A1(new_n18846_), .A2(\asqrt[55] ), .ZN(new_n19138_));
  AOI21_X1   g18946(.A1(new_n19138_), .A2(new_n18845_), .B(new_n724_), .ZN(new_n19139_));
  OAI21_X1   g18947(.A1(new_n18851_), .A2(new_n19139_), .B(\asqrt[57] ), .ZN(new_n19140_));
  AOI21_X1   g18948(.A1(new_n18858_), .A2(new_n19140_), .B(new_n504_), .ZN(new_n19141_));
  OAI21_X1   g18949(.A1(new_n18864_), .A2(new_n19141_), .B(\asqrt[59] ), .ZN(new_n19142_));
  AOI21_X1   g18950(.A1(new_n18871_), .A2(new_n19142_), .B(new_n275_), .ZN(new_n19143_));
  OAI21_X1   g18951(.A1(new_n18877_), .A2(new_n19143_), .B(\asqrt[61] ), .ZN(new_n19144_));
  NOR3_X1    g18952(.A1(new_n19106_), .A2(new_n19144_), .A3(new_n19087_), .ZN(new_n19145_));
  NOR3_X1    g18953(.A1(new_n19145_), .A2(new_n18898_), .A3(new_n19110_), .ZN(new_n19146_));
  OAI21_X1   g18954(.A1(new_n19146_), .A2(new_n18894_), .B(new_n19094_), .ZN(new_n19147_));
  NOR2_X1    g18955(.A1(new_n18888_), .A2(new_n19097_), .ZN(new_n19148_));
  NAND2_X1   g18956(.A1(new_n19148_), .A2(\asqrt[9] ), .ZN(new_n19149_));
  OAI21_X1   g18957(.A1(new_n19147_), .A2(new_n19149_), .B(new_n17656_), .ZN(new_n19150_));
  NAND3_X1   g18958(.A1(new_n19150_), .A2(new_n17663_), .A3(new_n19100_), .ZN(new_n19151_));
  NAND2_X1   g18959(.A1(new_n19061_), .A2(\asqrt[54] ), .ZN(new_n19152_));
  AOI21_X1   g18960(.A1(new_n19152_), .A2(new_n19060_), .B(new_n825_), .ZN(new_n19153_));
  OAI21_X1   g18961(.A1(new_n19063_), .A2(new_n19153_), .B(\asqrt[56] ), .ZN(new_n19154_));
  AOI21_X1   g18962(.A1(new_n19067_), .A2(new_n19154_), .B(new_n587_), .ZN(new_n19155_));
  OAI21_X1   g18963(.A1(new_n19070_), .A2(new_n19155_), .B(\asqrt[58] ), .ZN(new_n19156_));
  AOI21_X1   g18964(.A1(new_n19074_), .A2(new_n19156_), .B(new_n376_), .ZN(new_n19157_));
  OAI21_X1   g18965(.A1(new_n19077_), .A2(new_n19157_), .B(\asqrt[60] ), .ZN(new_n19158_));
  AOI21_X1   g18966(.A1(new_n19081_), .A2(new_n19158_), .B(new_n229_), .ZN(new_n19159_));
  NAND4_X1   g18967(.A1(new_n19159_), .A2(new_n18877_), .A3(new_n18883_), .A4(new_n19107_), .ZN(new_n19160_));
  NAND3_X1   g18968(.A1(new_n19160_), .A2(new_n19105_), .A3(new_n19091_), .ZN(new_n19161_));
  AOI21_X1   g18969(.A1(new_n19093_), .A2(new_n19161_), .B(new_n19123_), .ZN(new_n19162_));
  INV_X1     g18970(.I(new_n19149_), .ZN(new_n19163_));
  AOI21_X1   g18971(.A1(new_n19162_), .A2(new_n19163_), .B(\a[18] ), .ZN(new_n19164_));
  OAI21_X1   g18972(.A1(new_n19164_), .A2(new_n17664_), .B(\asqrt[8] ), .ZN(new_n19165_));
  NAND4_X1   g18973(.A1(new_n19165_), .A2(new_n19151_), .A3(new_n17893_), .A4(new_n19137_), .ZN(new_n19166_));
  NAND2_X1   g18974(.A1(new_n19166_), .A2(new_n19131_), .ZN(new_n19167_));
  NAND3_X1   g18975(.A1(new_n19127_), .A2(new_n19130_), .A3(new_n19137_), .ZN(new_n19168_));
  AOI21_X1   g18976(.A1(\asqrt[9] ), .A2(new_n17656_), .B(\a[19] ), .ZN(new_n19169_));
  NOR2_X1    g18977(.A1(new_n18485_), .A2(\a[18] ), .ZN(new_n19170_));
  AOI21_X1   g18978(.A1(\asqrt[9] ), .A2(\a[18] ), .B(new_n17666_), .ZN(new_n19171_));
  OAI21_X1   g18979(.A1(new_n19170_), .A2(new_n19169_), .B(new_n19171_), .ZN(new_n19172_));
  INV_X1     g18980(.I(new_n19172_), .ZN(new_n19173_));
  NAND3_X1   g18981(.A1(\asqrt[8] ), .A2(new_n18494_), .A3(new_n19173_), .ZN(new_n19174_));
  OAI21_X1   g18982(.A1(new_n19100_), .A2(new_n19172_), .B(new_n18493_), .ZN(new_n19175_));
  NAND3_X1   g18983(.A1(new_n19175_), .A2(new_n19174_), .A3(new_n17271_), .ZN(new_n19176_));
  AOI21_X1   g18984(.A1(new_n19168_), .A2(\asqrt[10] ), .B(new_n19176_), .ZN(new_n19177_));
  NOR2_X1    g18985(.A1(new_n19167_), .A2(new_n19177_), .ZN(new_n19178_));
  NAND2_X1   g18986(.A1(new_n19168_), .A2(\asqrt[10] ), .ZN(new_n19179_));
  AOI21_X1   g18987(.A1(new_n19167_), .A2(new_n19179_), .B(new_n17271_), .ZN(new_n19180_));
  NAND2_X1   g18988(.A1(new_n18515_), .A2(\asqrt[11] ), .ZN(new_n19181_));
  NAND2_X1   g18989(.A1(new_n18505_), .A2(new_n18512_), .ZN(new_n19182_));
  NAND3_X1   g18990(.A1(new_n19182_), .A2(new_n18907_), .A3(new_n17271_), .ZN(new_n19183_));
  NOR2_X1    g18991(.A1(new_n19100_), .A2(new_n19183_), .ZN(new_n19184_));
  AND2_X2    g18992(.A1(new_n19184_), .A2(new_n19181_), .Z(new_n19185_));
  NOR2_X1    g18993(.A1(new_n19184_), .A2(new_n19181_), .ZN(new_n19186_));
  NOR3_X1    g18994(.A1(new_n19185_), .A2(\asqrt[12] ), .A3(new_n19186_), .ZN(new_n19187_));
  INV_X1     g18995(.I(new_n19187_), .ZN(new_n19188_));
  OAI21_X1   g18996(.A1(new_n19180_), .A2(new_n19188_), .B(new_n19178_), .ZN(new_n19189_));
  OAI21_X1   g18997(.A1(new_n19180_), .A2(new_n19178_), .B(\asqrt[12] ), .ZN(new_n19190_));
  NAND2_X1   g18998(.A1(new_n18913_), .A2(\asqrt[12] ), .ZN(new_n19191_));
  NOR2_X1    g18999(.A1(new_n18909_), .A2(new_n18908_), .ZN(new_n19192_));
  NOR4_X1    g19000(.A1(new_n19100_), .A2(\asqrt[12] ), .A3(new_n19192_), .A4(new_n18913_), .ZN(new_n19193_));
  XOR2_X1    g19001(.A1(new_n19193_), .A2(new_n19191_), .Z(new_n19194_));
  NAND2_X1   g19002(.A1(new_n19194_), .A2(new_n16060_), .ZN(new_n19195_));
  INV_X1     g19003(.I(new_n19195_), .ZN(new_n19196_));
  AOI21_X1   g19004(.A1(new_n19190_), .A2(new_n19196_), .B(new_n19189_), .ZN(new_n19197_));
  AOI21_X1   g19005(.A1(new_n19189_), .A2(new_n19190_), .B(new_n16060_), .ZN(new_n19198_));
  NAND2_X1   g19006(.A1(new_n18537_), .A2(\asqrt[13] ), .ZN(new_n19199_));
  NOR2_X1    g19007(.A1(new_n18532_), .A2(new_n18533_), .ZN(new_n19200_));
  NOR4_X1    g19008(.A1(new_n19100_), .A2(\asqrt[13] ), .A3(new_n19200_), .A4(new_n18537_), .ZN(new_n19201_));
  XOR2_X1    g19009(.A1(new_n19201_), .A2(new_n19199_), .Z(new_n19202_));
  NAND2_X1   g19010(.A1(new_n19202_), .A2(new_n15447_), .ZN(new_n19203_));
  OAI21_X1   g19011(.A1(new_n19198_), .A2(new_n19203_), .B(new_n19197_), .ZN(new_n19204_));
  OAI21_X1   g19012(.A1(new_n19197_), .A2(new_n19198_), .B(\asqrt[14] ), .ZN(new_n19205_));
  NOR4_X1    g19013(.A1(new_n19100_), .A2(\asqrt[14] ), .A3(new_n18540_), .A4(new_n18921_), .ZN(new_n19206_));
  AOI21_X1   g19014(.A1(new_n19199_), .A2(new_n18536_), .B(new_n15447_), .ZN(new_n19207_));
  NOR2_X1    g19015(.A1(new_n19206_), .A2(new_n19207_), .ZN(new_n19208_));
  NAND2_X1   g19016(.A1(new_n19208_), .A2(new_n14871_), .ZN(new_n19209_));
  INV_X1     g19017(.I(new_n19209_), .ZN(new_n19210_));
  AOI21_X1   g19018(.A1(new_n19205_), .A2(new_n19210_), .B(new_n19204_), .ZN(new_n19211_));
  AOI22_X1   g19019(.A1(new_n19166_), .A2(new_n19131_), .B1(\asqrt[10] ), .B2(new_n19168_), .ZN(new_n19212_));
  OAI21_X1   g19020(.A1(new_n19212_), .A2(new_n17271_), .B(new_n19187_), .ZN(new_n19213_));
  OAI22_X1   g19021(.A1(new_n19212_), .A2(new_n17271_), .B1(new_n19167_), .B2(new_n19177_), .ZN(new_n19214_));
  AOI22_X1   g19022(.A1(new_n19214_), .A2(\asqrt[12] ), .B1(new_n19213_), .B2(new_n19178_), .ZN(new_n19215_));
  INV_X1     g19023(.I(new_n19203_), .ZN(new_n19216_));
  OAI21_X1   g19024(.A1(new_n19215_), .A2(new_n16060_), .B(new_n19216_), .ZN(new_n19217_));
  AOI21_X1   g19025(.A1(new_n19214_), .A2(\asqrt[12] ), .B(new_n19195_), .ZN(new_n19218_));
  OAI22_X1   g19026(.A1(new_n19215_), .A2(new_n16060_), .B1(new_n19218_), .B2(new_n19189_), .ZN(new_n19219_));
  AOI22_X1   g19027(.A1(new_n19219_), .A2(\asqrt[14] ), .B1(new_n19217_), .B2(new_n19197_), .ZN(new_n19220_));
  NAND2_X1   g19028(.A1(new_n18551_), .A2(\asqrt[15] ), .ZN(new_n19221_));
  NOR4_X1    g19029(.A1(new_n19100_), .A2(\asqrt[15] ), .A3(new_n18546_), .A4(new_n18551_), .ZN(new_n19222_));
  XOR2_X1    g19030(.A1(new_n19222_), .A2(new_n19221_), .Z(new_n19223_));
  NAND2_X1   g19031(.A1(new_n19223_), .A2(new_n14273_), .ZN(new_n19224_));
  INV_X1     g19032(.I(new_n19224_), .ZN(new_n19225_));
  OAI21_X1   g19033(.A1(new_n19220_), .A2(new_n14871_), .B(new_n19225_), .ZN(new_n19226_));
  NAND2_X1   g19034(.A1(new_n19226_), .A2(new_n19211_), .ZN(new_n19227_));
  AOI21_X1   g19035(.A1(new_n19219_), .A2(\asqrt[14] ), .B(new_n19209_), .ZN(new_n19228_));
  OAI22_X1   g19036(.A1(new_n19220_), .A2(new_n14871_), .B1(new_n19228_), .B2(new_n19204_), .ZN(new_n19229_));
  NOR4_X1    g19037(.A1(new_n19100_), .A2(\asqrt[16] ), .A3(new_n18554_), .A4(new_n18928_), .ZN(new_n19230_));
  AOI21_X1   g19038(.A1(new_n19221_), .A2(new_n18550_), .B(new_n14273_), .ZN(new_n19231_));
  NOR2_X1    g19039(.A1(new_n19230_), .A2(new_n19231_), .ZN(new_n19232_));
  NAND2_X1   g19040(.A1(new_n19232_), .A2(new_n13760_), .ZN(new_n19233_));
  AOI21_X1   g19041(.A1(new_n19229_), .A2(\asqrt[16] ), .B(new_n19233_), .ZN(new_n19234_));
  NOR2_X1    g19042(.A1(new_n19234_), .A2(new_n19227_), .ZN(new_n19235_));
  AOI22_X1   g19043(.A1(new_n19229_), .A2(\asqrt[16] ), .B1(new_n19226_), .B2(new_n19211_), .ZN(new_n19236_));
  NAND2_X1   g19044(.A1(new_n18565_), .A2(\asqrt[17] ), .ZN(new_n19237_));
  NOR4_X1    g19045(.A1(new_n19100_), .A2(\asqrt[17] ), .A3(new_n18560_), .A4(new_n18565_), .ZN(new_n19238_));
  XOR2_X1    g19046(.A1(new_n19238_), .A2(new_n19237_), .Z(new_n19239_));
  NAND2_X1   g19047(.A1(new_n19239_), .A2(new_n13192_), .ZN(new_n19240_));
  INV_X1     g19048(.I(new_n19240_), .ZN(new_n19241_));
  OAI21_X1   g19049(.A1(new_n19236_), .A2(new_n13760_), .B(new_n19241_), .ZN(new_n19242_));
  NAND2_X1   g19050(.A1(new_n19242_), .A2(new_n19235_), .ZN(new_n19243_));
  OAI22_X1   g19051(.A1(new_n19236_), .A2(new_n13760_), .B1(new_n19234_), .B2(new_n19227_), .ZN(new_n19244_));
  NOR4_X1    g19052(.A1(new_n19100_), .A2(\asqrt[18] ), .A3(new_n18567_), .A4(new_n18935_), .ZN(new_n19245_));
  AOI21_X1   g19053(.A1(new_n19237_), .A2(new_n18564_), .B(new_n13192_), .ZN(new_n19246_));
  NOR2_X1    g19054(.A1(new_n19245_), .A2(new_n19246_), .ZN(new_n19247_));
  NAND2_X1   g19055(.A1(new_n19247_), .A2(new_n12657_), .ZN(new_n19248_));
  AOI21_X1   g19056(.A1(new_n19244_), .A2(\asqrt[18] ), .B(new_n19248_), .ZN(new_n19249_));
  NOR2_X1    g19057(.A1(new_n19249_), .A2(new_n19243_), .ZN(new_n19250_));
  AOI22_X1   g19058(.A1(new_n19244_), .A2(\asqrt[18] ), .B1(new_n19242_), .B2(new_n19235_), .ZN(new_n19251_));
  NAND2_X1   g19059(.A1(new_n18578_), .A2(\asqrt[19] ), .ZN(new_n19252_));
  NOR4_X1    g19060(.A1(new_n19100_), .A2(\asqrt[19] ), .A3(new_n18573_), .A4(new_n18578_), .ZN(new_n19253_));
  XOR2_X1    g19061(.A1(new_n19253_), .A2(new_n19252_), .Z(new_n19254_));
  NAND2_X1   g19062(.A1(new_n19254_), .A2(new_n12101_), .ZN(new_n19255_));
  INV_X1     g19063(.I(new_n19255_), .ZN(new_n19256_));
  OAI21_X1   g19064(.A1(new_n19251_), .A2(new_n12657_), .B(new_n19256_), .ZN(new_n19257_));
  NAND2_X1   g19065(.A1(new_n19257_), .A2(new_n19250_), .ZN(new_n19258_));
  OAI22_X1   g19066(.A1(new_n19251_), .A2(new_n12657_), .B1(new_n19249_), .B2(new_n19243_), .ZN(new_n19259_));
  NAND2_X1   g19067(.A1(new_n18942_), .A2(\asqrt[20] ), .ZN(new_n19260_));
  NOR4_X1    g19068(.A1(new_n19100_), .A2(\asqrt[20] ), .A3(new_n18581_), .A4(new_n18942_), .ZN(new_n19261_));
  XOR2_X1    g19069(.A1(new_n19261_), .A2(new_n19260_), .Z(new_n19262_));
  NAND2_X1   g19070(.A1(new_n19262_), .A2(new_n11631_), .ZN(new_n19263_));
  AOI21_X1   g19071(.A1(new_n19259_), .A2(\asqrt[20] ), .B(new_n19263_), .ZN(new_n19264_));
  NOR2_X1    g19072(.A1(new_n19264_), .A2(new_n19258_), .ZN(new_n19265_));
  AOI22_X1   g19073(.A1(new_n19259_), .A2(\asqrt[20] ), .B1(new_n19257_), .B2(new_n19250_), .ZN(new_n19266_));
  NOR4_X1    g19074(.A1(new_n19100_), .A2(\asqrt[21] ), .A3(new_n18588_), .A4(new_n18593_), .ZN(new_n19267_));
  AOI21_X1   g19075(.A1(new_n19260_), .A2(new_n18941_), .B(new_n11631_), .ZN(new_n19268_));
  NOR2_X1    g19076(.A1(new_n19267_), .A2(new_n19268_), .ZN(new_n19269_));
  NAND2_X1   g19077(.A1(new_n19269_), .A2(new_n11105_), .ZN(new_n19270_));
  INV_X1     g19078(.I(new_n19270_), .ZN(new_n19271_));
  OAI21_X1   g19079(.A1(new_n19266_), .A2(new_n11631_), .B(new_n19271_), .ZN(new_n19272_));
  NAND2_X1   g19080(.A1(new_n19272_), .A2(new_n19265_), .ZN(new_n19273_));
  OAI22_X1   g19081(.A1(new_n19266_), .A2(new_n11631_), .B1(new_n19264_), .B2(new_n19258_), .ZN(new_n19274_));
  NAND2_X1   g19082(.A1(new_n18949_), .A2(\asqrt[22] ), .ZN(new_n19275_));
  NOR4_X1    g19083(.A1(new_n19100_), .A2(\asqrt[22] ), .A3(new_n18596_), .A4(new_n18949_), .ZN(new_n19276_));
  XOR2_X1    g19084(.A1(new_n19276_), .A2(new_n19275_), .Z(new_n19277_));
  NAND2_X1   g19085(.A1(new_n19277_), .A2(new_n10614_), .ZN(new_n19278_));
  AOI21_X1   g19086(.A1(new_n19274_), .A2(\asqrt[22] ), .B(new_n19278_), .ZN(new_n19279_));
  NOR2_X1    g19087(.A1(new_n19279_), .A2(new_n19273_), .ZN(new_n19280_));
  AOI22_X1   g19088(.A1(new_n19274_), .A2(\asqrt[22] ), .B1(new_n19272_), .B2(new_n19265_), .ZN(new_n19281_));
  NOR4_X1    g19089(.A1(new_n19100_), .A2(\asqrt[23] ), .A3(new_n18603_), .A4(new_n18608_), .ZN(new_n19282_));
  AOI21_X1   g19090(.A1(new_n19275_), .A2(new_n18948_), .B(new_n10614_), .ZN(new_n19283_));
  NOR2_X1    g19091(.A1(new_n19282_), .A2(new_n19283_), .ZN(new_n19284_));
  NAND2_X1   g19092(.A1(new_n19284_), .A2(new_n10104_), .ZN(new_n19285_));
  INV_X1     g19093(.I(new_n19285_), .ZN(new_n19286_));
  OAI21_X1   g19094(.A1(new_n19281_), .A2(new_n10614_), .B(new_n19286_), .ZN(new_n19287_));
  NAND2_X1   g19095(.A1(new_n19287_), .A2(new_n19280_), .ZN(new_n19288_));
  OAI22_X1   g19096(.A1(new_n19281_), .A2(new_n10614_), .B1(new_n19279_), .B2(new_n19273_), .ZN(new_n19289_));
  NAND2_X1   g19097(.A1(new_n18956_), .A2(\asqrt[24] ), .ZN(new_n19290_));
  NOR4_X1    g19098(.A1(new_n19100_), .A2(\asqrt[24] ), .A3(new_n18611_), .A4(new_n18956_), .ZN(new_n19291_));
  XOR2_X1    g19099(.A1(new_n19291_), .A2(new_n19290_), .Z(new_n19292_));
  NAND2_X1   g19100(.A1(new_n19292_), .A2(new_n9672_), .ZN(new_n19293_));
  AOI21_X1   g19101(.A1(new_n19289_), .A2(\asqrt[24] ), .B(new_n19293_), .ZN(new_n19294_));
  NOR2_X1    g19102(.A1(new_n19294_), .A2(new_n19288_), .ZN(new_n19295_));
  AOI22_X1   g19103(.A1(new_n19289_), .A2(\asqrt[24] ), .B1(new_n19287_), .B2(new_n19280_), .ZN(new_n19296_));
  NOR4_X1    g19104(.A1(new_n19100_), .A2(\asqrt[25] ), .A3(new_n18618_), .A4(new_n18623_), .ZN(new_n19297_));
  AOI21_X1   g19105(.A1(new_n19290_), .A2(new_n18955_), .B(new_n9672_), .ZN(new_n19298_));
  NOR2_X1    g19106(.A1(new_n19297_), .A2(new_n19298_), .ZN(new_n19299_));
  NAND2_X1   g19107(.A1(new_n19299_), .A2(new_n9212_), .ZN(new_n19300_));
  INV_X1     g19108(.I(new_n19300_), .ZN(new_n19301_));
  OAI21_X1   g19109(.A1(new_n19296_), .A2(new_n9672_), .B(new_n19301_), .ZN(new_n19302_));
  NAND2_X1   g19110(.A1(new_n19302_), .A2(new_n19295_), .ZN(new_n19303_));
  OAI22_X1   g19111(.A1(new_n19296_), .A2(new_n9672_), .B1(new_n19294_), .B2(new_n19288_), .ZN(new_n19304_));
  NAND2_X1   g19112(.A1(new_n18963_), .A2(\asqrt[26] ), .ZN(new_n19305_));
  NOR4_X1    g19113(.A1(new_n19100_), .A2(\asqrt[26] ), .A3(new_n18626_), .A4(new_n18963_), .ZN(new_n19306_));
  XOR2_X1    g19114(.A1(new_n19306_), .A2(new_n19305_), .Z(new_n19307_));
  NAND2_X1   g19115(.A1(new_n19307_), .A2(new_n8763_), .ZN(new_n19308_));
  AOI21_X1   g19116(.A1(new_n19304_), .A2(\asqrt[26] ), .B(new_n19308_), .ZN(new_n19309_));
  NOR2_X1    g19117(.A1(new_n19309_), .A2(new_n19303_), .ZN(new_n19310_));
  AOI22_X1   g19118(.A1(new_n19304_), .A2(\asqrt[26] ), .B1(new_n19302_), .B2(new_n19295_), .ZN(new_n19311_));
  NOR4_X1    g19119(.A1(new_n19100_), .A2(\asqrt[27] ), .A3(new_n18633_), .A4(new_n18638_), .ZN(new_n19312_));
  AOI21_X1   g19120(.A1(new_n19305_), .A2(new_n18962_), .B(new_n8763_), .ZN(new_n19313_));
  NOR2_X1    g19121(.A1(new_n19312_), .A2(new_n19313_), .ZN(new_n19314_));
  NAND2_X1   g19122(.A1(new_n19314_), .A2(new_n8319_), .ZN(new_n19315_));
  INV_X1     g19123(.I(new_n19315_), .ZN(new_n19316_));
  OAI21_X1   g19124(.A1(new_n19311_), .A2(new_n8763_), .B(new_n19316_), .ZN(new_n19317_));
  NAND2_X1   g19125(.A1(new_n19317_), .A2(new_n19310_), .ZN(new_n19318_));
  OAI22_X1   g19126(.A1(new_n19311_), .A2(new_n8763_), .B1(new_n19309_), .B2(new_n19303_), .ZN(new_n19319_));
  NAND2_X1   g19127(.A1(new_n18970_), .A2(\asqrt[28] ), .ZN(new_n19320_));
  NOR4_X1    g19128(.A1(new_n19100_), .A2(\asqrt[28] ), .A3(new_n18641_), .A4(new_n18970_), .ZN(new_n19321_));
  XOR2_X1    g19129(.A1(new_n19321_), .A2(new_n19320_), .Z(new_n19322_));
  NAND2_X1   g19130(.A1(new_n19322_), .A2(new_n7931_), .ZN(new_n19323_));
  AOI21_X1   g19131(.A1(new_n19319_), .A2(\asqrt[28] ), .B(new_n19323_), .ZN(new_n19324_));
  NOR2_X1    g19132(.A1(new_n19324_), .A2(new_n19318_), .ZN(new_n19325_));
  AOI22_X1   g19133(.A1(new_n19319_), .A2(\asqrt[28] ), .B1(new_n19317_), .B2(new_n19310_), .ZN(new_n19326_));
  NAND2_X1   g19134(.A1(new_n18653_), .A2(\asqrt[29] ), .ZN(new_n19327_));
  NOR4_X1    g19135(.A1(new_n19100_), .A2(\asqrt[29] ), .A3(new_n18648_), .A4(new_n18653_), .ZN(new_n19328_));
  XOR2_X1    g19136(.A1(new_n19328_), .A2(new_n19327_), .Z(new_n19329_));
  NAND2_X1   g19137(.A1(new_n19329_), .A2(new_n7517_), .ZN(new_n19330_));
  INV_X1     g19138(.I(new_n19330_), .ZN(new_n19331_));
  OAI21_X1   g19139(.A1(new_n19326_), .A2(new_n7931_), .B(new_n19331_), .ZN(new_n19332_));
  NAND2_X1   g19140(.A1(new_n19332_), .A2(new_n19325_), .ZN(new_n19333_));
  OAI22_X1   g19141(.A1(new_n19326_), .A2(new_n7931_), .B1(new_n19324_), .B2(new_n19318_), .ZN(new_n19334_));
  NOR4_X1    g19142(.A1(new_n19100_), .A2(\asqrt[30] ), .A3(new_n18656_), .A4(new_n18977_), .ZN(new_n19335_));
  AOI21_X1   g19143(.A1(new_n19327_), .A2(new_n18652_), .B(new_n7517_), .ZN(new_n19336_));
  NOR2_X1    g19144(.A1(new_n19335_), .A2(new_n19336_), .ZN(new_n19337_));
  NAND2_X1   g19145(.A1(new_n19337_), .A2(new_n7110_), .ZN(new_n19338_));
  AOI21_X1   g19146(.A1(new_n19334_), .A2(\asqrt[30] ), .B(new_n19338_), .ZN(new_n19339_));
  NOR2_X1    g19147(.A1(new_n19339_), .A2(new_n19333_), .ZN(new_n19340_));
  AOI22_X1   g19148(.A1(new_n19334_), .A2(\asqrt[30] ), .B1(new_n19332_), .B2(new_n19325_), .ZN(new_n19341_));
  NAND2_X1   g19149(.A1(new_n18668_), .A2(\asqrt[31] ), .ZN(new_n19342_));
  NOR4_X1    g19150(.A1(new_n19100_), .A2(\asqrt[31] ), .A3(new_n18663_), .A4(new_n18668_), .ZN(new_n19343_));
  XOR2_X1    g19151(.A1(new_n19343_), .A2(new_n19342_), .Z(new_n19344_));
  NAND2_X1   g19152(.A1(new_n19344_), .A2(new_n6708_), .ZN(new_n19345_));
  INV_X1     g19153(.I(new_n19345_), .ZN(new_n19346_));
  OAI21_X1   g19154(.A1(new_n19341_), .A2(new_n7110_), .B(new_n19346_), .ZN(new_n19347_));
  NAND2_X1   g19155(.A1(new_n19347_), .A2(new_n19340_), .ZN(new_n19348_));
  OAI22_X1   g19156(.A1(new_n19341_), .A2(new_n7110_), .B1(new_n19339_), .B2(new_n19333_), .ZN(new_n19349_));
  NOR4_X1    g19157(.A1(new_n19100_), .A2(\asqrt[32] ), .A3(new_n18671_), .A4(new_n18984_), .ZN(new_n19350_));
  AOI21_X1   g19158(.A1(new_n19342_), .A2(new_n18667_), .B(new_n6708_), .ZN(new_n19351_));
  NOR2_X1    g19159(.A1(new_n19350_), .A2(new_n19351_), .ZN(new_n19352_));
  NAND2_X1   g19160(.A1(new_n19352_), .A2(new_n6365_), .ZN(new_n19353_));
  AOI21_X1   g19161(.A1(new_n19349_), .A2(\asqrt[32] ), .B(new_n19353_), .ZN(new_n19354_));
  NOR2_X1    g19162(.A1(new_n19354_), .A2(new_n19348_), .ZN(new_n19355_));
  AOI22_X1   g19163(.A1(new_n19349_), .A2(\asqrt[32] ), .B1(new_n19347_), .B2(new_n19340_), .ZN(new_n19356_));
  NAND2_X1   g19164(.A1(new_n18683_), .A2(\asqrt[33] ), .ZN(new_n19357_));
  NOR4_X1    g19165(.A1(new_n19100_), .A2(\asqrt[33] ), .A3(new_n18678_), .A4(new_n18683_), .ZN(new_n19358_));
  XOR2_X1    g19166(.A1(new_n19358_), .A2(new_n19357_), .Z(new_n19359_));
  NAND2_X1   g19167(.A1(new_n19359_), .A2(new_n5991_), .ZN(new_n19360_));
  INV_X1     g19168(.I(new_n19360_), .ZN(new_n19361_));
  OAI21_X1   g19169(.A1(new_n19356_), .A2(new_n6365_), .B(new_n19361_), .ZN(new_n19362_));
  NAND2_X1   g19170(.A1(new_n19362_), .A2(new_n19355_), .ZN(new_n19363_));
  OAI22_X1   g19171(.A1(new_n19356_), .A2(new_n6365_), .B1(new_n19354_), .B2(new_n19348_), .ZN(new_n19364_));
  NOR4_X1    g19172(.A1(new_n19100_), .A2(\asqrt[34] ), .A3(new_n18686_), .A4(new_n18991_), .ZN(new_n19365_));
  AOI21_X1   g19173(.A1(new_n19357_), .A2(new_n18682_), .B(new_n5991_), .ZN(new_n19366_));
  NOR2_X1    g19174(.A1(new_n19365_), .A2(new_n19366_), .ZN(new_n19367_));
  NAND2_X1   g19175(.A1(new_n19367_), .A2(new_n5626_), .ZN(new_n19368_));
  AOI21_X1   g19176(.A1(new_n19364_), .A2(\asqrt[34] ), .B(new_n19368_), .ZN(new_n19369_));
  NOR2_X1    g19177(.A1(new_n19369_), .A2(new_n19363_), .ZN(new_n19370_));
  AOI22_X1   g19178(.A1(new_n19364_), .A2(\asqrt[34] ), .B1(new_n19362_), .B2(new_n19355_), .ZN(new_n19371_));
  NAND2_X1   g19179(.A1(new_n18698_), .A2(\asqrt[35] ), .ZN(new_n19372_));
  NOR4_X1    g19180(.A1(new_n19100_), .A2(\asqrt[35] ), .A3(new_n18693_), .A4(new_n18698_), .ZN(new_n19373_));
  XOR2_X1    g19181(.A1(new_n19373_), .A2(new_n19372_), .Z(new_n19374_));
  NAND2_X1   g19182(.A1(new_n19374_), .A2(new_n5273_), .ZN(new_n19375_));
  INV_X1     g19183(.I(new_n19375_), .ZN(new_n19376_));
  OAI21_X1   g19184(.A1(new_n19371_), .A2(new_n5626_), .B(new_n19376_), .ZN(new_n19377_));
  NAND2_X1   g19185(.A1(new_n19377_), .A2(new_n19370_), .ZN(new_n19378_));
  OAI22_X1   g19186(.A1(new_n19371_), .A2(new_n5626_), .B1(new_n19369_), .B2(new_n19363_), .ZN(new_n19379_));
  NAND2_X1   g19187(.A1(new_n18998_), .A2(\asqrt[36] ), .ZN(new_n19380_));
  NOR4_X1    g19188(.A1(new_n19100_), .A2(\asqrt[36] ), .A3(new_n18701_), .A4(new_n18998_), .ZN(new_n19381_));
  XOR2_X1    g19189(.A1(new_n19381_), .A2(new_n19380_), .Z(new_n19382_));
  NAND2_X1   g19190(.A1(new_n19382_), .A2(new_n4973_), .ZN(new_n19383_));
  AOI21_X1   g19191(.A1(new_n19379_), .A2(\asqrt[36] ), .B(new_n19383_), .ZN(new_n19384_));
  NOR2_X1    g19192(.A1(new_n19384_), .A2(new_n19378_), .ZN(new_n19385_));
  AOI22_X1   g19193(.A1(new_n19379_), .A2(\asqrt[36] ), .B1(new_n19377_), .B2(new_n19370_), .ZN(new_n19386_));
  NOR4_X1    g19194(.A1(new_n19100_), .A2(\asqrt[37] ), .A3(new_n18708_), .A4(new_n18713_), .ZN(new_n19387_));
  AOI21_X1   g19195(.A1(new_n19380_), .A2(new_n18997_), .B(new_n4973_), .ZN(new_n19388_));
  NOR2_X1    g19196(.A1(new_n19387_), .A2(new_n19388_), .ZN(new_n19389_));
  NAND2_X1   g19197(.A1(new_n19389_), .A2(new_n4645_), .ZN(new_n19390_));
  INV_X1     g19198(.I(new_n19390_), .ZN(new_n19391_));
  OAI21_X1   g19199(.A1(new_n19386_), .A2(new_n4973_), .B(new_n19391_), .ZN(new_n19392_));
  NAND2_X1   g19200(.A1(new_n19392_), .A2(new_n19385_), .ZN(new_n19393_));
  OAI22_X1   g19201(.A1(new_n19386_), .A2(new_n4973_), .B1(new_n19384_), .B2(new_n19378_), .ZN(new_n19394_));
  NAND2_X1   g19202(.A1(new_n19005_), .A2(\asqrt[38] ), .ZN(new_n19395_));
  NOR4_X1    g19203(.A1(new_n19100_), .A2(\asqrt[38] ), .A3(new_n18716_), .A4(new_n19005_), .ZN(new_n19396_));
  XOR2_X1    g19204(.A1(new_n19396_), .A2(new_n19395_), .Z(new_n19397_));
  NAND2_X1   g19205(.A1(new_n19397_), .A2(new_n4330_), .ZN(new_n19398_));
  AOI21_X1   g19206(.A1(new_n19394_), .A2(\asqrt[38] ), .B(new_n19398_), .ZN(new_n19399_));
  NOR2_X1    g19207(.A1(new_n19399_), .A2(new_n19393_), .ZN(new_n19400_));
  AOI22_X1   g19208(.A1(new_n19394_), .A2(\asqrt[38] ), .B1(new_n19392_), .B2(new_n19385_), .ZN(new_n19401_));
  NOR4_X1    g19209(.A1(new_n19100_), .A2(\asqrt[39] ), .A3(new_n18723_), .A4(new_n18728_), .ZN(new_n19402_));
  AOI21_X1   g19210(.A1(new_n19395_), .A2(new_n19004_), .B(new_n4330_), .ZN(new_n19403_));
  NOR2_X1    g19211(.A1(new_n19402_), .A2(new_n19403_), .ZN(new_n19404_));
  NAND2_X1   g19212(.A1(new_n19404_), .A2(new_n4018_), .ZN(new_n19405_));
  INV_X1     g19213(.I(new_n19405_), .ZN(new_n19406_));
  OAI21_X1   g19214(.A1(new_n19401_), .A2(new_n4330_), .B(new_n19406_), .ZN(new_n19407_));
  NAND2_X1   g19215(.A1(new_n19407_), .A2(new_n19400_), .ZN(new_n19408_));
  OAI22_X1   g19216(.A1(new_n19401_), .A2(new_n4330_), .B1(new_n19399_), .B2(new_n19393_), .ZN(new_n19409_));
  NAND2_X1   g19217(.A1(new_n19012_), .A2(\asqrt[40] ), .ZN(new_n19410_));
  NOR4_X1    g19218(.A1(new_n19100_), .A2(\asqrt[40] ), .A3(new_n18731_), .A4(new_n19012_), .ZN(new_n19411_));
  XOR2_X1    g19219(.A1(new_n19411_), .A2(new_n19410_), .Z(new_n19412_));
  NAND2_X1   g19220(.A1(new_n19412_), .A2(new_n3760_), .ZN(new_n19413_));
  AOI21_X1   g19221(.A1(new_n19409_), .A2(\asqrt[40] ), .B(new_n19413_), .ZN(new_n19414_));
  NOR2_X1    g19222(.A1(new_n19414_), .A2(new_n19408_), .ZN(new_n19415_));
  AOI22_X1   g19223(.A1(new_n19409_), .A2(\asqrt[40] ), .B1(new_n19407_), .B2(new_n19400_), .ZN(new_n19416_));
  NAND2_X1   g19224(.A1(new_n18743_), .A2(\asqrt[41] ), .ZN(new_n19417_));
  NOR4_X1    g19225(.A1(new_n19100_), .A2(\asqrt[41] ), .A3(new_n18738_), .A4(new_n18743_), .ZN(new_n19418_));
  XOR2_X1    g19226(.A1(new_n19418_), .A2(new_n19417_), .Z(new_n19419_));
  NAND2_X1   g19227(.A1(new_n19419_), .A2(new_n3481_), .ZN(new_n19420_));
  INV_X1     g19228(.I(new_n19420_), .ZN(new_n19421_));
  OAI21_X1   g19229(.A1(new_n19416_), .A2(new_n3760_), .B(new_n19421_), .ZN(new_n19422_));
  NAND2_X1   g19230(.A1(new_n19422_), .A2(new_n19415_), .ZN(new_n19423_));
  OAI22_X1   g19231(.A1(new_n19416_), .A2(new_n3760_), .B1(new_n19414_), .B2(new_n19408_), .ZN(new_n19424_));
  NOR4_X1    g19232(.A1(new_n19100_), .A2(\asqrt[42] ), .A3(new_n18746_), .A4(new_n19019_), .ZN(new_n19425_));
  AOI21_X1   g19233(.A1(new_n19417_), .A2(new_n18742_), .B(new_n3481_), .ZN(new_n19426_));
  NOR2_X1    g19234(.A1(new_n19425_), .A2(new_n19426_), .ZN(new_n19427_));
  NAND2_X1   g19235(.A1(new_n19427_), .A2(new_n3208_), .ZN(new_n19428_));
  AOI21_X1   g19236(.A1(new_n19424_), .A2(\asqrt[42] ), .B(new_n19428_), .ZN(new_n19429_));
  NOR2_X1    g19237(.A1(new_n19429_), .A2(new_n19423_), .ZN(new_n19430_));
  AOI22_X1   g19238(.A1(new_n19424_), .A2(\asqrt[42] ), .B1(new_n19422_), .B2(new_n19415_), .ZN(new_n19431_));
  NAND2_X1   g19239(.A1(new_n18758_), .A2(\asqrt[43] ), .ZN(new_n19432_));
  NOR4_X1    g19240(.A1(new_n19100_), .A2(\asqrt[43] ), .A3(new_n18753_), .A4(new_n18758_), .ZN(new_n19433_));
  XOR2_X1    g19241(.A1(new_n19433_), .A2(new_n19432_), .Z(new_n19434_));
  NAND2_X1   g19242(.A1(new_n19434_), .A2(new_n2941_), .ZN(new_n19435_));
  INV_X1     g19243(.I(new_n19435_), .ZN(new_n19436_));
  OAI21_X1   g19244(.A1(new_n19431_), .A2(new_n3208_), .B(new_n19436_), .ZN(new_n19437_));
  NAND2_X1   g19245(.A1(new_n19437_), .A2(new_n19430_), .ZN(new_n19438_));
  OAI22_X1   g19246(.A1(new_n19431_), .A2(new_n3208_), .B1(new_n19429_), .B2(new_n19423_), .ZN(new_n19439_));
  NOR4_X1    g19247(.A1(new_n19100_), .A2(\asqrt[44] ), .A3(new_n18761_), .A4(new_n19026_), .ZN(new_n19440_));
  AOI21_X1   g19248(.A1(new_n19432_), .A2(new_n18757_), .B(new_n2941_), .ZN(new_n19441_));
  NOR2_X1    g19249(.A1(new_n19440_), .A2(new_n19441_), .ZN(new_n19442_));
  NAND2_X1   g19250(.A1(new_n19442_), .A2(new_n2728_), .ZN(new_n19443_));
  AOI21_X1   g19251(.A1(new_n19439_), .A2(\asqrt[44] ), .B(new_n19443_), .ZN(new_n19444_));
  NOR2_X1    g19252(.A1(new_n19444_), .A2(new_n19438_), .ZN(new_n19445_));
  AOI22_X1   g19253(.A1(new_n19439_), .A2(\asqrt[44] ), .B1(new_n19437_), .B2(new_n19430_), .ZN(new_n19446_));
  NAND2_X1   g19254(.A1(new_n18773_), .A2(\asqrt[45] ), .ZN(new_n19447_));
  NOR4_X1    g19255(.A1(new_n19100_), .A2(\asqrt[45] ), .A3(new_n18768_), .A4(new_n18773_), .ZN(new_n19448_));
  XOR2_X1    g19256(.A1(new_n19448_), .A2(new_n19447_), .Z(new_n19449_));
  NAND2_X1   g19257(.A1(new_n19449_), .A2(new_n2488_), .ZN(new_n19450_));
  INV_X1     g19258(.I(new_n19450_), .ZN(new_n19451_));
  OAI21_X1   g19259(.A1(new_n19446_), .A2(new_n2728_), .B(new_n19451_), .ZN(new_n19452_));
  NAND2_X1   g19260(.A1(new_n19452_), .A2(new_n19445_), .ZN(new_n19453_));
  OAI22_X1   g19261(.A1(new_n19446_), .A2(new_n2728_), .B1(new_n19444_), .B2(new_n19438_), .ZN(new_n19454_));
  NOR4_X1    g19262(.A1(new_n19100_), .A2(\asqrt[46] ), .A3(new_n18776_), .A4(new_n19033_), .ZN(new_n19455_));
  AOI21_X1   g19263(.A1(new_n19447_), .A2(new_n18772_), .B(new_n2488_), .ZN(new_n19456_));
  NOR2_X1    g19264(.A1(new_n19455_), .A2(new_n19456_), .ZN(new_n19457_));
  NAND2_X1   g19265(.A1(new_n19457_), .A2(new_n2253_), .ZN(new_n19458_));
  AOI21_X1   g19266(.A1(new_n19454_), .A2(\asqrt[46] ), .B(new_n19458_), .ZN(new_n19459_));
  NOR2_X1    g19267(.A1(new_n19459_), .A2(new_n19453_), .ZN(new_n19460_));
  AOI22_X1   g19268(.A1(new_n19454_), .A2(\asqrt[46] ), .B1(new_n19452_), .B2(new_n19445_), .ZN(new_n19461_));
  NAND2_X1   g19269(.A1(new_n18788_), .A2(\asqrt[47] ), .ZN(new_n19462_));
  NOR4_X1    g19270(.A1(new_n19100_), .A2(\asqrt[47] ), .A3(new_n18783_), .A4(new_n18788_), .ZN(new_n19463_));
  XOR2_X1    g19271(.A1(new_n19463_), .A2(new_n19462_), .Z(new_n19464_));
  NAND2_X1   g19272(.A1(new_n19464_), .A2(new_n2046_), .ZN(new_n19465_));
  INV_X1     g19273(.I(new_n19465_), .ZN(new_n19466_));
  OAI21_X1   g19274(.A1(new_n19461_), .A2(new_n2253_), .B(new_n19466_), .ZN(new_n19467_));
  NAND2_X1   g19275(.A1(new_n19467_), .A2(new_n19460_), .ZN(new_n19468_));
  OAI22_X1   g19276(.A1(new_n19461_), .A2(new_n2253_), .B1(new_n19459_), .B2(new_n19453_), .ZN(new_n19469_));
  NAND2_X1   g19277(.A1(new_n19040_), .A2(\asqrt[48] ), .ZN(new_n19470_));
  NOR4_X1    g19278(.A1(new_n19100_), .A2(\asqrt[48] ), .A3(new_n18791_), .A4(new_n19040_), .ZN(new_n19471_));
  XOR2_X1    g19279(.A1(new_n19471_), .A2(new_n19470_), .Z(new_n19472_));
  NAND2_X1   g19280(.A1(new_n19472_), .A2(new_n1854_), .ZN(new_n19473_));
  AOI21_X1   g19281(.A1(new_n19469_), .A2(\asqrt[48] ), .B(new_n19473_), .ZN(new_n19474_));
  NOR2_X1    g19282(.A1(new_n19474_), .A2(new_n19468_), .ZN(new_n19475_));
  AOI22_X1   g19283(.A1(new_n19469_), .A2(\asqrt[48] ), .B1(new_n19467_), .B2(new_n19460_), .ZN(new_n19476_));
  NOR4_X1    g19284(.A1(new_n19100_), .A2(\asqrt[49] ), .A3(new_n18798_), .A4(new_n18803_), .ZN(new_n19477_));
  AOI21_X1   g19285(.A1(new_n19470_), .A2(new_n19039_), .B(new_n1854_), .ZN(new_n19478_));
  NOR2_X1    g19286(.A1(new_n19477_), .A2(new_n19478_), .ZN(new_n19479_));
  NAND2_X1   g19287(.A1(new_n19479_), .A2(new_n1595_), .ZN(new_n19480_));
  INV_X1     g19288(.I(new_n19480_), .ZN(new_n19481_));
  OAI21_X1   g19289(.A1(new_n19476_), .A2(new_n1854_), .B(new_n19481_), .ZN(new_n19482_));
  NAND2_X1   g19290(.A1(new_n19482_), .A2(new_n19475_), .ZN(new_n19483_));
  OAI22_X1   g19291(.A1(new_n19476_), .A2(new_n1854_), .B1(new_n19474_), .B2(new_n19468_), .ZN(new_n19484_));
  NAND2_X1   g19292(.A1(new_n19047_), .A2(\asqrt[50] ), .ZN(new_n19485_));
  NOR4_X1    g19293(.A1(new_n19100_), .A2(\asqrt[50] ), .A3(new_n18806_), .A4(new_n19047_), .ZN(new_n19486_));
  XOR2_X1    g19294(.A1(new_n19486_), .A2(new_n19485_), .Z(new_n19487_));
  NAND2_X1   g19295(.A1(new_n19487_), .A2(new_n1436_), .ZN(new_n19488_));
  AOI21_X1   g19296(.A1(new_n19484_), .A2(\asqrt[50] ), .B(new_n19488_), .ZN(new_n19489_));
  NOR2_X1    g19297(.A1(new_n19489_), .A2(new_n19483_), .ZN(new_n19490_));
  AOI22_X1   g19298(.A1(new_n19484_), .A2(\asqrt[50] ), .B1(new_n19482_), .B2(new_n19475_), .ZN(new_n19491_));
  NOR4_X1    g19299(.A1(new_n19100_), .A2(\asqrt[51] ), .A3(new_n18813_), .A4(new_n18818_), .ZN(new_n19492_));
  AOI21_X1   g19300(.A1(new_n19485_), .A2(new_n19046_), .B(new_n1436_), .ZN(new_n19493_));
  NOR2_X1    g19301(.A1(new_n19492_), .A2(new_n19493_), .ZN(new_n19494_));
  NAND2_X1   g19302(.A1(new_n19494_), .A2(new_n1260_), .ZN(new_n19495_));
  INV_X1     g19303(.I(new_n19495_), .ZN(new_n19496_));
  OAI21_X1   g19304(.A1(new_n19491_), .A2(new_n1436_), .B(new_n19496_), .ZN(new_n19497_));
  NAND2_X1   g19305(.A1(new_n19497_), .A2(new_n19490_), .ZN(new_n19498_));
  OAI22_X1   g19306(.A1(new_n19491_), .A2(new_n1436_), .B1(new_n19489_), .B2(new_n19483_), .ZN(new_n19499_));
  NAND2_X1   g19307(.A1(new_n19054_), .A2(\asqrt[52] ), .ZN(new_n19500_));
  NOR4_X1    g19308(.A1(new_n19100_), .A2(\asqrt[52] ), .A3(new_n18821_), .A4(new_n19054_), .ZN(new_n19501_));
  XOR2_X1    g19309(.A1(new_n19501_), .A2(new_n19500_), .Z(new_n19502_));
  NAND2_X1   g19310(.A1(new_n19502_), .A2(new_n1096_), .ZN(new_n19503_));
  AOI21_X1   g19311(.A1(new_n19499_), .A2(\asqrt[52] ), .B(new_n19503_), .ZN(new_n19504_));
  NOR2_X1    g19312(.A1(new_n19504_), .A2(new_n19498_), .ZN(new_n19505_));
  AOI22_X1   g19313(.A1(new_n19499_), .A2(\asqrt[52] ), .B1(new_n19497_), .B2(new_n19490_), .ZN(new_n19506_));
  NOR2_X1    g19314(.A1(new_n19057_), .A2(new_n1096_), .ZN(new_n19507_));
  NOR4_X1    g19315(.A1(new_n19100_), .A2(\asqrt[53] ), .A3(new_n18828_), .A4(new_n18833_), .ZN(new_n19508_));
  XNOR2_X1   g19316(.A1(new_n19508_), .A2(new_n19507_), .ZN(new_n19509_));
  NAND2_X1   g19317(.A1(new_n19509_), .A2(new_n970_), .ZN(new_n19510_));
  INV_X1     g19318(.I(new_n19510_), .ZN(new_n19511_));
  OAI21_X1   g19319(.A1(new_n19506_), .A2(new_n1096_), .B(new_n19511_), .ZN(new_n19512_));
  NAND2_X1   g19320(.A1(new_n19512_), .A2(new_n19505_), .ZN(new_n19513_));
  OAI22_X1   g19321(.A1(new_n19506_), .A2(new_n1096_), .B1(new_n19504_), .B2(new_n19498_), .ZN(new_n19514_));
  NOR4_X1    g19322(.A1(new_n19100_), .A2(\asqrt[54] ), .A3(new_n18835_), .A4(new_n19061_), .ZN(new_n19515_));
  XOR2_X1    g19323(.A1(new_n19515_), .A2(new_n19152_), .Z(new_n19516_));
  NAND2_X1   g19324(.A1(new_n19516_), .A2(new_n825_), .ZN(new_n19517_));
  AOI21_X1   g19325(.A1(new_n19514_), .A2(\asqrt[54] ), .B(new_n19517_), .ZN(new_n19518_));
  NOR2_X1    g19326(.A1(new_n19518_), .A2(new_n19513_), .ZN(new_n19519_));
  AOI22_X1   g19327(.A1(new_n19514_), .A2(\asqrt[54] ), .B1(new_n19512_), .B2(new_n19505_), .ZN(new_n19520_));
  NOR4_X1    g19328(.A1(new_n19100_), .A2(\asqrt[55] ), .A3(new_n18841_), .A4(new_n18846_), .ZN(new_n19521_));
  XOR2_X1    g19329(.A1(new_n19521_), .A2(new_n19138_), .Z(new_n19522_));
  NAND2_X1   g19330(.A1(new_n19522_), .A2(new_n724_), .ZN(new_n19523_));
  INV_X1     g19331(.I(new_n19523_), .ZN(new_n19524_));
  OAI21_X1   g19332(.A1(new_n19520_), .A2(new_n825_), .B(new_n19524_), .ZN(new_n19525_));
  NAND2_X1   g19333(.A1(new_n19525_), .A2(new_n19519_), .ZN(new_n19526_));
  OAI22_X1   g19334(.A1(new_n19520_), .A2(new_n825_), .B1(new_n19518_), .B2(new_n19513_), .ZN(new_n19527_));
  NOR4_X1    g19335(.A1(new_n19100_), .A2(\asqrt[56] ), .A3(new_n18848_), .A4(new_n19068_), .ZN(new_n19528_));
  XOR2_X1    g19336(.A1(new_n19528_), .A2(new_n19154_), .Z(new_n19529_));
  NAND2_X1   g19337(.A1(new_n19529_), .A2(new_n587_), .ZN(new_n19530_));
  AOI21_X1   g19338(.A1(new_n19527_), .A2(\asqrt[56] ), .B(new_n19530_), .ZN(new_n19531_));
  NOR2_X1    g19339(.A1(new_n19531_), .A2(new_n19526_), .ZN(new_n19532_));
  AOI22_X1   g19340(.A1(new_n19527_), .A2(\asqrt[56] ), .B1(new_n19525_), .B2(new_n19519_), .ZN(new_n19533_));
  NOR4_X1    g19341(.A1(new_n19100_), .A2(\asqrt[57] ), .A3(new_n18854_), .A4(new_n18859_), .ZN(new_n19534_));
  XOR2_X1    g19342(.A1(new_n19534_), .A2(new_n19140_), .Z(new_n19535_));
  NAND2_X1   g19343(.A1(new_n19535_), .A2(new_n504_), .ZN(new_n19536_));
  INV_X1     g19344(.I(new_n19536_), .ZN(new_n19537_));
  OAI21_X1   g19345(.A1(new_n19533_), .A2(new_n587_), .B(new_n19537_), .ZN(new_n19538_));
  NAND2_X1   g19346(.A1(new_n19538_), .A2(new_n19532_), .ZN(new_n19539_));
  OAI22_X1   g19347(.A1(new_n19533_), .A2(new_n587_), .B1(new_n19531_), .B2(new_n19526_), .ZN(new_n19540_));
  NOR4_X1    g19348(.A1(new_n19100_), .A2(\asqrt[58] ), .A3(new_n18861_), .A4(new_n19075_), .ZN(new_n19541_));
  XOR2_X1    g19349(.A1(new_n19541_), .A2(new_n19156_), .Z(new_n19542_));
  NAND2_X1   g19350(.A1(new_n19542_), .A2(new_n376_), .ZN(new_n19543_));
  AOI21_X1   g19351(.A1(new_n19540_), .A2(\asqrt[58] ), .B(new_n19543_), .ZN(new_n19544_));
  NOR2_X1    g19352(.A1(new_n19544_), .A2(new_n19539_), .ZN(new_n19545_));
  AOI22_X1   g19353(.A1(new_n19540_), .A2(\asqrt[58] ), .B1(new_n19538_), .B2(new_n19532_), .ZN(new_n19546_));
  NOR4_X1    g19354(.A1(new_n19100_), .A2(\asqrt[59] ), .A3(new_n18867_), .A4(new_n18872_), .ZN(new_n19547_));
  XOR2_X1    g19355(.A1(new_n19547_), .A2(new_n19142_), .Z(new_n19548_));
  AND2_X2    g19356(.A1(new_n19548_), .A2(new_n275_), .Z(new_n19549_));
  OAI21_X1   g19357(.A1(new_n19546_), .A2(new_n376_), .B(new_n19549_), .ZN(new_n19550_));
  NAND2_X1   g19358(.A1(new_n19550_), .A2(new_n19545_), .ZN(new_n19551_));
  OAI22_X1   g19359(.A1(new_n19546_), .A2(new_n376_), .B1(new_n19544_), .B2(new_n19539_), .ZN(new_n19552_));
  AOI22_X1   g19360(.A1(new_n19552_), .A2(\asqrt[60] ), .B1(new_n19550_), .B2(new_n19545_), .ZN(new_n19553_));
  NOR4_X1    g19361(.A1(new_n19100_), .A2(\asqrt[60] ), .A3(new_n18874_), .A4(new_n19082_), .ZN(new_n19554_));
  XOR2_X1    g19362(.A1(new_n19554_), .A2(new_n19158_), .Z(new_n19555_));
  NAND2_X1   g19363(.A1(new_n19555_), .A2(new_n229_), .ZN(new_n19556_));
  AOI21_X1   g19364(.A1(new_n19552_), .A2(\asqrt[60] ), .B(new_n19556_), .ZN(new_n19557_));
  OAI22_X1   g19365(.A1(new_n19553_), .A2(new_n229_), .B1(new_n19557_), .B2(new_n19551_), .ZN(new_n19558_));
  NOR4_X1    g19366(.A1(new_n19100_), .A2(\asqrt[61] ), .A3(new_n18880_), .A4(new_n18884_), .ZN(new_n19559_));
  XOR2_X1    g19367(.A1(new_n19559_), .A2(new_n19144_), .Z(new_n19560_));
  NOR4_X1    g19368(.A1(new_n19558_), .A2(\asqrt[62] ), .A3(new_n19115_), .A4(new_n19560_), .ZN(new_n19561_));
  NOR2_X1    g19369(.A1(new_n19560_), .A2(new_n196_), .ZN(new_n19562_));
  INV_X1     g19370(.I(new_n19562_), .ZN(new_n19563_));
  NOR2_X1    g19371(.A1(new_n19198_), .A2(new_n19203_), .ZN(new_n19564_));
  NOR3_X1    g19372(.A1(new_n19564_), .A2(new_n19189_), .A3(new_n19218_), .ZN(new_n19565_));
  NAND2_X1   g19373(.A1(new_n19205_), .A2(new_n19210_), .ZN(new_n19566_));
  NAND2_X1   g19374(.A1(new_n19566_), .A2(new_n19565_), .ZN(new_n19567_));
  NAND2_X1   g19375(.A1(new_n19204_), .A2(new_n19205_), .ZN(new_n19568_));
  AOI21_X1   g19376(.A1(new_n19568_), .A2(\asqrt[15] ), .B(new_n19224_), .ZN(new_n19569_));
  NOR2_X1    g19377(.A1(new_n19569_), .A2(new_n19567_), .ZN(new_n19570_));
  AOI21_X1   g19378(.A1(new_n19204_), .A2(new_n19205_), .B(new_n14871_), .ZN(new_n19571_));
  OAI21_X1   g19379(.A1(new_n19211_), .A2(new_n19571_), .B(\asqrt[16] ), .ZN(new_n19572_));
  INV_X1     g19380(.I(new_n19233_), .ZN(new_n19573_));
  NAND2_X1   g19381(.A1(new_n19572_), .A2(new_n19573_), .ZN(new_n19574_));
  NAND2_X1   g19382(.A1(new_n19574_), .A2(new_n19570_), .ZN(new_n19575_));
  AOI22_X1   g19383(.A1(new_n19568_), .A2(\asqrt[15] ), .B1(new_n19566_), .B2(new_n19565_), .ZN(new_n19576_));
  OAI22_X1   g19384(.A1(new_n19576_), .A2(new_n14273_), .B1(new_n19569_), .B2(new_n19567_), .ZN(new_n19577_));
  AOI21_X1   g19385(.A1(new_n19577_), .A2(\asqrt[17] ), .B(new_n19240_), .ZN(new_n19578_));
  NOR2_X1    g19386(.A1(new_n19578_), .A2(new_n19575_), .ZN(new_n19579_));
  AOI22_X1   g19387(.A1(new_n19577_), .A2(\asqrt[17] ), .B1(new_n19574_), .B2(new_n19570_), .ZN(new_n19580_));
  INV_X1     g19388(.I(new_n19248_), .ZN(new_n19581_));
  OAI21_X1   g19389(.A1(new_n19580_), .A2(new_n13192_), .B(new_n19581_), .ZN(new_n19582_));
  NAND2_X1   g19390(.A1(new_n19582_), .A2(new_n19579_), .ZN(new_n19583_));
  OAI22_X1   g19391(.A1(new_n19580_), .A2(new_n13192_), .B1(new_n19578_), .B2(new_n19575_), .ZN(new_n19584_));
  AOI21_X1   g19392(.A1(new_n19584_), .A2(\asqrt[19] ), .B(new_n19255_), .ZN(new_n19585_));
  NOR2_X1    g19393(.A1(new_n19585_), .A2(new_n19583_), .ZN(new_n19586_));
  AOI22_X1   g19394(.A1(new_n19584_), .A2(\asqrt[19] ), .B1(new_n19582_), .B2(new_n19579_), .ZN(new_n19587_));
  INV_X1     g19395(.I(new_n19263_), .ZN(new_n19588_));
  OAI21_X1   g19396(.A1(new_n19587_), .A2(new_n12101_), .B(new_n19588_), .ZN(new_n19589_));
  NAND2_X1   g19397(.A1(new_n19589_), .A2(new_n19586_), .ZN(new_n19590_));
  OAI22_X1   g19398(.A1(new_n19587_), .A2(new_n12101_), .B1(new_n19585_), .B2(new_n19583_), .ZN(new_n19591_));
  AOI21_X1   g19399(.A1(new_n19591_), .A2(\asqrt[21] ), .B(new_n19270_), .ZN(new_n19592_));
  NOR2_X1    g19400(.A1(new_n19592_), .A2(new_n19590_), .ZN(new_n19593_));
  AOI22_X1   g19401(.A1(new_n19591_), .A2(\asqrt[21] ), .B1(new_n19589_), .B2(new_n19586_), .ZN(new_n19594_));
  INV_X1     g19402(.I(new_n19278_), .ZN(new_n19595_));
  OAI21_X1   g19403(.A1(new_n19594_), .A2(new_n11105_), .B(new_n19595_), .ZN(new_n19596_));
  NAND2_X1   g19404(.A1(new_n19596_), .A2(new_n19593_), .ZN(new_n19597_));
  OAI22_X1   g19405(.A1(new_n19594_), .A2(new_n11105_), .B1(new_n19592_), .B2(new_n19590_), .ZN(new_n19598_));
  AOI21_X1   g19406(.A1(new_n19598_), .A2(\asqrt[23] ), .B(new_n19285_), .ZN(new_n19599_));
  NOR2_X1    g19407(.A1(new_n19599_), .A2(new_n19597_), .ZN(new_n19600_));
  AOI22_X1   g19408(.A1(new_n19598_), .A2(\asqrt[23] ), .B1(new_n19596_), .B2(new_n19593_), .ZN(new_n19601_));
  INV_X1     g19409(.I(new_n19293_), .ZN(new_n19602_));
  OAI21_X1   g19410(.A1(new_n19601_), .A2(new_n10104_), .B(new_n19602_), .ZN(new_n19603_));
  NAND2_X1   g19411(.A1(new_n19603_), .A2(new_n19600_), .ZN(new_n19604_));
  OAI22_X1   g19412(.A1(new_n19601_), .A2(new_n10104_), .B1(new_n19599_), .B2(new_n19597_), .ZN(new_n19605_));
  AOI21_X1   g19413(.A1(new_n19605_), .A2(\asqrt[25] ), .B(new_n19300_), .ZN(new_n19606_));
  NOR2_X1    g19414(.A1(new_n19606_), .A2(new_n19604_), .ZN(new_n19607_));
  AOI22_X1   g19415(.A1(new_n19605_), .A2(\asqrt[25] ), .B1(new_n19603_), .B2(new_n19600_), .ZN(new_n19608_));
  INV_X1     g19416(.I(new_n19308_), .ZN(new_n19609_));
  OAI21_X1   g19417(.A1(new_n19608_), .A2(new_n9212_), .B(new_n19609_), .ZN(new_n19610_));
  NAND2_X1   g19418(.A1(new_n19610_), .A2(new_n19607_), .ZN(new_n19611_));
  OAI22_X1   g19419(.A1(new_n19608_), .A2(new_n9212_), .B1(new_n19606_), .B2(new_n19604_), .ZN(new_n19612_));
  AOI21_X1   g19420(.A1(new_n19612_), .A2(\asqrt[27] ), .B(new_n19315_), .ZN(new_n19613_));
  NOR2_X1    g19421(.A1(new_n19613_), .A2(new_n19611_), .ZN(new_n19614_));
  AOI22_X1   g19422(.A1(new_n19612_), .A2(\asqrt[27] ), .B1(new_n19610_), .B2(new_n19607_), .ZN(new_n19615_));
  INV_X1     g19423(.I(new_n19323_), .ZN(new_n19616_));
  OAI21_X1   g19424(.A1(new_n19615_), .A2(new_n8319_), .B(new_n19616_), .ZN(new_n19617_));
  NAND2_X1   g19425(.A1(new_n19617_), .A2(new_n19614_), .ZN(new_n19618_));
  OAI22_X1   g19426(.A1(new_n19615_), .A2(new_n8319_), .B1(new_n19613_), .B2(new_n19611_), .ZN(new_n19619_));
  AOI21_X1   g19427(.A1(new_n19619_), .A2(\asqrt[29] ), .B(new_n19330_), .ZN(new_n19620_));
  NOR2_X1    g19428(.A1(new_n19620_), .A2(new_n19618_), .ZN(new_n19621_));
  AOI22_X1   g19429(.A1(new_n19619_), .A2(\asqrt[29] ), .B1(new_n19617_), .B2(new_n19614_), .ZN(new_n19622_));
  INV_X1     g19430(.I(new_n19338_), .ZN(new_n19623_));
  OAI21_X1   g19431(.A1(new_n19622_), .A2(new_n7517_), .B(new_n19623_), .ZN(new_n19624_));
  NAND2_X1   g19432(.A1(new_n19624_), .A2(new_n19621_), .ZN(new_n19625_));
  OAI22_X1   g19433(.A1(new_n19622_), .A2(new_n7517_), .B1(new_n19620_), .B2(new_n19618_), .ZN(new_n19626_));
  AOI21_X1   g19434(.A1(new_n19626_), .A2(\asqrt[31] ), .B(new_n19345_), .ZN(new_n19627_));
  NOR2_X1    g19435(.A1(new_n19627_), .A2(new_n19625_), .ZN(new_n19628_));
  AOI22_X1   g19436(.A1(new_n19626_), .A2(\asqrt[31] ), .B1(new_n19624_), .B2(new_n19621_), .ZN(new_n19629_));
  INV_X1     g19437(.I(new_n19353_), .ZN(new_n19630_));
  OAI21_X1   g19438(.A1(new_n19629_), .A2(new_n6708_), .B(new_n19630_), .ZN(new_n19631_));
  NAND2_X1   g19439(.A1(new_n19631_), .A2(new_n19628_), .ZN(new_n19632_));
  OAI22_X1   g19440(.A1(new_n19629_), .A2(new_n6708_), .B1(new_n19627_), .B2(new_n19625_), .ZN(new_n19633_));
  AOI21_X1   g19441(.A1(new_n19633_), .A2(\asqrt[33] ), .B(new_n19360_), .ZN(new_n19634_));
  NOR2_X1    g19442(.A1(new_n19634_), .A2(new_n19632_), .ZN(new_n19635_));
  AOI22_X1   g19443(.A1(new_n19633_), .A2(\asqrt[33] ), .B1(new_n19631_), .B2(new_n19628_), .ZN(new_n19636_));
  INV_X1     g19444(.I(new_n19368_), .ZN(new_n19637_));
  OAI21_X1   g19445(.A1(new_n19636_), .A2(new_n5991_), .B(new_n19637_), .ZN(new_n19638_));
  NAND2_X1   g19446(.A1(new_n19638_), .A2(new_n19635_), .ZN(new_n19639_));
  OAI22_X1   g19447(.A1(new_n19636_), .A2(new_n5991_), .B1(new_n19634_), .B2(new_n19632_), .ZN(new_n19640_));
  AOI21_X1   g19448(.A1(new_n19640_), .A2(\asqrt[35] ), .B(new_n19375_), .ZN(new_n19641_));
  NOR2_X1    g19449(.A1(new_n19641_), .A2(new_n19639_), .ZN(new_n19642_));
  AOI22_X1   g19450(.A1(new_n19640_), .A2(\asqrt[35] ), .B1(new_n19638_), .B2(new_n19635_), .ZN(new_n19643_));
  INV_X1     g19451(.I(new_n19383_), .ZN(new_n19644_));
  OAI21_X1   g19452(.A1(new_n19643_), .A2(new_n5273_), .B(new_n19644_), .ZN(new_n19645_));
  NAND2_X1   g19453(.A1(new_n19645_), .A2(new_n19642_), .ZN(new_n19646_));
  OAI22_X1   g19454(.A1(new_n19643_), .A2(new_n5273_), .B1(new_n19641_), .B2(new_n19639_), .ZN(new_n19647_));
  AOI21_X1   g19455(.A1(new_n19647_), .A2(\asqrt[37] ), .B(new_n19390_), .ZN(new_n19648_));
  NOR2_X1    g19456(.A1(new_n19648_), .A2(new_n19646_), .ZN(new_n19649_));
  AOI22_X1   g19457(.A1(new_n19647_), .A2(\asqrt[37] ), .B1(new_n19645_), .B2(new_n19642_), .ZN(new_n19650_));
  INV_X1     g19458(.I(new_n19398_), .ZN(new_n19651_));
  OAI21_X1   g19459(.A1(new_n19650_), .A2(new_n4645_), .B(new_n19651_), .ZN(new_n19652_));
  NAND2_X1   g19460(.A1(new_n19652_), .A2(new_n19649_), .ZN(new_n19653_));
  OAI22_X1   g19461(.A1(new_n19650_), .A2(new_n4645_), .B1(new_n19648_), .B2(new_n19646_), .ZN(new_n19654_));
  AOI21_X1   g19462(.A1(new_n19654_), .A2(\asqrt[39] ), .B(new_n19405_), .ZN(new_n19655_));
  NOR2_X1    g19463(.A1(new_n19655_), .A2(new_n19653_), .ZN(new_n19656_));
  AOI22_X1   g19464(.A1(new_n19654_), .A2(\asqrt[39] ), .B1(new_n19652_), .B2(new_n19649_), .ZN(new_n19657_));
  INV_X1     g19465(.I(new_n19413_), .ZN(new_n19658_));
  OAI21_X1   g19466(.A1(new_n19657_), .A2(new_n4018_), .B(new_n19658_), .ZN(new_n19659_));
  NAND2_X1   g19467(.A1(new_n19659_), .A2(new_n19656_), .ZN(new_n19660_));
  OAI22_X1   g19468(.A1(new_n19657_), .A2(new_n4018_), .B1(new_n19655_), .B2(new_n19653_), .ZN(new_n19661_));
  AOI21_X1   g19469(.A1(new_n19661_), .A2(\asqrt[41] ), .B(new_n19420_), .ZN(new_n19662_));
  NOR2_X1    g19470(.A1(new_n19662_), .A2(new_n19660_), .ZN(new_n19663_));
  AOI22_X1   g19471(.A1(new_n19661_), .A2(\asqrt[41] ), .B1(new_n19659_), .B2(new_n19656_), .ZN(new_n19664_));
  INV_X1     g19472(.I(new_n19428_), .ZN(new_n19665_));
  OAI21_X1   g19473(.A1(new_n19664_), .A2(new_n3481_), .B(new_n19665_), .ZN(new_n19666_));
  NAND2_X1   g19474(.A1(new_n19666_), .A2(new_n19663_), .ZN(new_n19667_));
  OAI22_X1   g19475(.A1(new_n19664_), .A2(new_n3481_), .B1(new_n19662_), .B2(new_n19660_), .ZN(new_n19668_));
  AOI21_X1   g19476(.A1(new_n19668_), .A2(\asqrt[43] ), .B(new_n19435_), .ZN(new_n19669_));
  NOR2_X1    g19477(.A1(new_n19669_), .A2(new_n19667_), .ZN(new_n19670_));
  AOI22_X1   g19478(.A1(new_n19668_), .A2(\asqrt[43] ), .B1(new_n19666_), .B2(new_n19663_), .ZN(new_n19671_));
  INV_X1     g19479(.I(new_n19443_), .ZN(new_n19672_));
  OAI21_X1   g19480(.A1(new_n19671_), .A2(new_n2941_), .B(new_n19672_), .ZN(new_n19673_));
  NAND2_X1   g19481(.A1(new_n19673_), .A2(new_n19670_), .ZN(new_n19674_));
  OAI22_X1   g19482(.A1(new_n19671_), .A2(new_n2941_), .B1(new_n19669_), .B2(new_n19667_), .ZN(new_n19675_));
  AOI21_X1   g19483(.A1(new_n19675_), .A2(\asqrt[45] ), .B(new_n19450_), .ZN(new_n19676_));
  NOR2_X1    g19484(.A1(new_n19676_), .A2(new_n19674_), .ZN(new_n19677_));
  AOI22_X1   g19485(.A1(new_n19675_), .A2(\asqrt[45] ), .B1(new_n19673_), .B2(new_n19670_), .ZN(new_n19678_));
  INV_X1     g19486(.I(new_n19458_), .ZN(new_n19679_));
  OAI21_X1   g19487(.A1(new_n19678_), .A2(new_n2488_), .B(new_n19679_), .ZN(new_n19680_));
  NAND2_X1   g19488(.A1(new_n19680_), .A2(new_n19677_), .ZN(new_n19681_));
  OAI22_X1   g19489(.A1(new_n19678_), .A2(new_n2488_), .B1(new_n19676_), .B2(new_n19674_), .ZN(new_n19682_));
  AOI21_X1   g19490(.A1(new_n19682_), .A2(\asqrt[47] ), .B(new_n19465_), .ZN(new_n19683_));
  NOR2_X1    g19491(.A1(new_n19683_), .A2(new_n19681_), .ZN(new_n19684_));
  AOI22_X1   g19492(.A1(new_n19682_), .A2(\asqrt[47] ), .B1(new_n19680_), .B2(new_n19677_), .ZN(new_n19685_));
  INV_X1     g19493(.I(new_n19473_), .ZN(new_n19686_));
  OAI21_X1   g19494(.A1(new_n19685_), .A2(new_n2046_), .B(new_n19686_), .ZN(new_n19687_));
  NAND2_X1   g19495(.A1(new_n19687_), .A2(new_n19684_), .ZN(new_n19688_));
  OAI22_X1   g19496(.A1(new_n19685_), .A2(new_n2046_), .B1(new_n19683_), .B2(new_n19681_), .ZN(new_n19689_));
  AOI21_X1   g19497(.A1(new_n19689_), .A2(\asqrt[49] ), .B(new_n19480_), .ZN(new_n19690_));
  NOR2_X1    g19498(.A1(new_n19690_), .A2(new_n19688_), .ZN(new_n19691_));
  AOI22_X1   g19499(.A1(new_n19689_), .A2(\asqrt[49] ), .B1(new_n19687_), .B2(new_n19684_), .ZN(new_n19692_));
  INV_X1     g19500(.I(new_n19488_), .ZN(new_n19693_));
  OAI21_X1   g19501(.A1(new_n19692_), .A2(new_n1595_), .B(new_n19693_), .ZN(new_n19694_));
  NAND2_X1   g19502(.A1(new_n19694_), .A2(new_n19691_), .ZN(new_n19695_));
  OAI22_X1   g19503(.A1(new_n19692_), .A2(new_n1595_), .B1(new_n19690_), .B2(new_n19688_), .ZN(new_n19696_));
  AOI21_X1   g19504(.A1(new_n19696_), .A2(\asqrt[51] ), .B(new_n19495_), .ZN(new_n19697_));
  NOR2_X1    g19505(.A1(new_n19697_), .A2(new_n19695_), .ZN(new_n19698_));
  AOI22_X1   g19506(.A1(new_n19696_), .A2(\asqrt[51] ), .B1(new_n19694_), .B2(new_n19691_), .ZN(new_n19699_));
  INV_X1     g19507(.I(new_n19503_), .ZN(new_n19700_));
  OAI21_X1   g19508(.A1(new_n19699_), .A2(new_n1260_), .B(new_n19700_), .ZN(new_n19701_));
  NAND2_X1   g19509(.A1(new_n19701_), .A2(new_n19698_), .ZN(new_n19702_));
  OAI22_X1   g19510(.A1(new_n19699_), .A2(new_n1260_), .B1(new_n19697_), .B2(new_n19695_), .ZN(new_n19703_));
  AOI21_X1   g19511(.A1(new_n19703_), .A2(\asqrt[53] ), .B(new_n19510_), .ZN(new_n19704_));
  NOR2_X1    g19512(.A1(new_n19704_), .A2(new_n19702_), .ZN(new_n19705_));
  AOI22_X1   g19513(.A1(new_n19703_), .A2(\asqrt[53] ), .B1(new_n19701_), .B2(new_n19698_), .ZN(new_n19706_));
  INV_X1     g19514(.I(new_n19517_), .ZN(new_n19707_));
  OAI21_X1   g19515(.A1(new_n19706_), .A2(new_n970_), .B(new_n19707_), .ZN(new_n19708_));
  NAND2_X1   g19516(.A1(new_n19708_), .A2(new_n19705_), .ZN(new_n19709_));
  OAI22_X1   g19517(.A1(new_n19706_), .A2(new_n970_), .B1(new_n19704_), .B2(new_n19702_), .ZN(new_n19710_));
  AOI21_X1   g19518(.A1(new_n19710_), .A2(\asqrt[55] ), .B(new_n19523_), .ZN(new_n19711_));
  NOR2_X1    g19519(.A1(new_n19711_), .A2(new_n19709_), .ZN(new_n19712_));
  AOI22_X1   g19520(.A1(new_n19710_), .A2(\asqrt[55] ), .B1(new_n19708_), .B2(new_n19705_), .ZN(new_n19713_));
  INV_X1     g19521(.I(new_n19530_), .ZN(new_n19714_));
  OAI21_X1   g19522(.A1(new_n19713_), .A2(new_n724_), .B(new_n19714_), .ZN(new_n19715_));
  NAND2_X1   g19523(.A1(new_n19715_), .A2(new_n19712_), .ZN(new_n19716_));
  NAND2_X1   g19524(.A1(new_n19710_), .A2(\asqrt[55] ), .ZN(new_n19717_));
  AOI21_X1   g19525(.A1(new_n19717_), .A2(new_n19709_), .B(new_n724_), .ZN(new_n19718_));
  OAI21_X1   g19526(.A1(new_n19712_), .A2(new_n19718_), .B(\asqrt[57] ), .ZN(new_n19719_));
  AOI21_X1   g19527(.A1(new_n19719_), .A2(new_n19537_), .B(new_n19716_), .ZN(new_n19720_));
  OAI22_X1   g19528(.A1(new_n19713_), .A2(new_n724_), .B1(new_n19711_), .B2(new_n19709_), .ZN(new_n19721_));
  AOI22_X1   g19529(.A1(new_n19721_), .A2(\asqrt[57] ), .B1(new_n19715_), .B2(new_n19712_), .ZN(new_n19722_));
  INV_X1     g19530(.I(new_n19543_), .ZN(new_n19723_));
  OAI21_X1   g19531(.A1(new_n19722_), .A2(new_n504_), .B(new_n19723_), .ZN(new_n19724_));
  NAND2_X1   g19532(.A1(new_n19724_), .A2(new_n19720_), .ZN(new_n19725_));
  AOI21_X1   g19533(.A1(new_n19716_), .A2(new_n19719_), .B(new_n504_), .ZN(new_n19726_));
  OAI21_X1   g19534(.A1(new_n19720_), .A2(new_n19726_), .B(\asqrt[59] ), .ZN(new_n19727_));
  AOI21_X1   g19535(.A1(new_n19727_), .A2(new_n19549_), .B(new_n19725_), .ZN(new_n19728_));
  NAND2_X1   g19536(.A1(new_n19514_), .A2(\asqrt[54] ), .ZN(new_n19729_));
  AOI21_X1   g19537(.A1(new_n19729_), .A2(new_n19513_), .B(new_n825_), .ZN(new_n19730_));
  OAI21_X1   g19538(.A1(new_n19519_), .A2(new_n19730_), .B(\asqrt[56] ), .ZN(new_n19731_));
  AOI21_X1   g19539(.A1(new_n19526_), .A2(new_n19731_), .B(new_n587_), .ZN(new_n19732_));
  OAI21_X1   g19540(.A1(new_n19532_), .A2(new_n19732_), .B(\asqrt[58] ), .ZN(new_n19733_));
  AOI21_X1   g19541(.A1(new_n19539_), .A2(new_n19733_), .B(new_n376_), .ZN(new_n19734_));
  OAI21_X1   g19542(.A1(new_n19545_), .A2(new_n19734_), .B(\asqrt[60] ), .ZN(new_n19735_));
  AOI21_X1   g19543(.A1(new_n19551_), .A2(new_n19735_), .B(new_n229_), .ZN(new_n19736_));
  NAND2_X1   g19544(.A1(new_n19539_), .A2(new_n19733_), .ZN(new_n19737_));
  AOI22_X1   g19545(.A1(new_n19737_), .A2(\asqrt[59] ), .B1(new_n19724_), .B2(new_n19720_), .ZN(new_n19738_));
  INV_X1     g19546(.I(new_n19556_), .ZN(new_n19739_));
  OAI21_X1   g19547(.A1(new_n19738_), .A2(new_n275_), .B(new_n19739_), .ZN(new_n19740_));
  INV_X1     g19548(.I(new_n19560_), .ZN(new_n19741_));
  NOR2_X1    g19549(.A1(new_n19741_), .A2(\asqrt[62] ), .ZN(new_n19742_));
  INV_X1     g19550(.I(new_n19742_), .ZN(new_n19743_));
  NAND4_X1   g19551(.A1(new_n19736_), .A2(new_n19728_), .A3(new_n19740_), .A4(new_n19743_), .ZN(new_n19744_));
  NOR3_X1    g19552(.A1(\asqrt[8] ), .A2(new_n19093_), .A3(new_n19123_), .ZN(new_n19745_));
  OAI21_X1   g19553(.A1(new_n19745_), .A2(new_n19089_), .B(new_n231_), .ZN(new_n19746_));
  INV_X1     g19554(.I(new_n19746_), .ZN(new_n19747_));
  NAND3_X1   g19555(.A1(new_n19744_), .A2(new_n19563_), .A3(new_n19747_), .ZN(new_n19748_));
  AOI21_X1   g19556(.A1(new_n19114_), .A2(new_n19748_), .B(new_n19561_), .ZN(new_n19749_));
  INV_X1     g19557(.I(\a[12] ), .ZN(new_n19750_));
  NAND3_X1   g19558(.A1(new_n19132_), .A2(new_n18887_), .A3(new_n19093_), .ZN(new_n19751_));
  INV_X1     g19559(.I(new_n19751_), .ZN(new_n19752_));
  OAI21_X1   g19560(.A1(new_n19093_), .A2(new_n19109_), .B(\asqrt[8] ), .ZN(new_n19753_));
  XOR2_X1    g19561(.A1(new_n19109_), .A2(\asqrt[63] ), .Z(new_n19754_));
  NAND2_X1   g19562(.A1(new_n19753_), .A2(new_n19754_), .ZN(new_n19755_));
  INV_X1     g19563(.I(new_n19755_), .ZN(new_n19756_));
  NOR2_X1    g19564(.A1(new_n19756_), .A2(new_n19752_), .ZN(new_n19757_));
  NOR2_X1    g19565(.A1(\a[10] ), .A2(\a[11] ), .ZN(new_n19758_));
  INV_X1     g19566(.I(new_n19758_), .ZN(new_n19759_));
  NOR3_X1    g19567(.A1(new_n19757_), .A2(new_n19750_), .A3(new_n19759_), .ZN(new_n19760_));
  NAND2_X1   g19568(.A1(new_n19749_), .A2(new_n19760_), .ZN(new_n19761_));
  XOR2_X1    g19569(.A1(new_n19761_), .A2(\a[13] ), .Z(new_n19762_));
  INV_X1     g19570(.I(new_n19762_), .ZN(new_n19763_));
  NAND2_X1   g19571(.A1(new_n19740_), .A2(new_n19728_), .ZN(new_n19764_));
  NAND2_X1   g19572(.A1(new_n19736_), .A2(new_n19743_), .ZN(new_n19765_));
  OAI21_X1   g19573(.A1(new_n19765_), .A2(new_n19764_), .B(new_n19563_), .ZN(new_n19766_));
  OAI21_X1   g19574(.A1(new_n19766_), .A2(new_n19746_), .B(new_n19114_), .ZN(new_n19767_));
  NAND2_X1   g19575(.A1(new_n19561_), .A2(new_n19756_), .ZN(new_n19768_));
  NOR2_X1    g19576(.A1(new_n19768_), .A2(new_n19767_), .ZN(new_n19769_));
  NOR2_X1    g19577(.A1(new_n19115_), .A2(new_n19752_), .ZN(new_n19770_));
  NAND2_X1   g19578(.A1(new_n19769_), .A2(new_n19770_), .ZN(new_n19771_));
  INV_X1     g19579(.I(new_n19771_), .ZN(new_n19772_));
  NAND2_X1   g19580(.A1(new_n19551_), .A2(new_n19735_), .ZN(new_n19773_));
  AOI22_X1   g19581(.A1(new_n19773_), .A2(\asqrt[61] ), .B1(new_n19740_), .B2(new_n19728_), .ZN(new_n19774_));
  NOR2_X1    g19582(.A1(new_n19774_), .A2(new_n196_), .ZN(new_n19775_));
  NOR2_X1    g19583(.A1(new_n19557_), .A2(new_n19551_), .ZN(new_n19776_));
  NOR3_X1    g19584(.A1(new_n19553_), .A2(new_n229_), .A3(new_n19742_), .ZN(new_n19777_));
  AOI21_X1   g19585(.A1(new_n19777_), .A2(new_n19776_), .B(new_n19562_), .ZN(new_n19778_));
  AOI21_X1   g19586(.A1(new_n19778_), .A2(new_n19747_), .B(new_n19115_), .ZN(new_n19779_));
  NAND4_X1   g19587(.A1(new_n19774_), .A2(new_n196_), .A3(new_n19114_), .A4(new_n19741_), .ZN(new_n19780_));
  NOR2_X1    g19588(.A1(new_n19780_), .A2(new_n19755_), .ZN(new_n19781_));
  NAND3_X1   g19589(.A1(new_n19781_), .A2(new_n19779_), .A3(new_n19752_), .ZN(new_n19782_));
  NOR4_X1    g19590(.A1(new_n19782_), .A2(\asqrt[62] ), .A3(new_n19558_), .A4(new_n19560_), .ZN(new_n19783_));
  XNOR2_X1   g19591(.A1(new_n19783_), .A2(new_n19775_), .ZN(new_n19784_));
  NOR3_X1    g19592(.A1(new_n19768_), .A2(new_n19767_), .A3(new_n19751_), .ZN(\asqrt[7] ));
  NOR3_X1    g19593(.A1(new_n19773_), .A2(\asqrt[61] ), .A3(new_n19555_), .ZN(new_n19786_));
  NAND2_X1   g19594(.A1(\asqrt[7] ), .A2(new_n19786_), .ZN(new_n19787_));
  XOR2_X1    g19595(.A1(new_n19787_), .A2(new_n19736_), .Z(new_n19788_));
  NOR2_X1    g19596(.A1(new_n19788_), .A2(new_n196_), .ZN(new_n19789_));
  INV_X1     g19597(.I(\a[14] ), .ZN(new_n19790_));
  NOR2_X1    g19598(.A1(\a[12] ), .A2(\a[13] ), .ZN(new_n19791_));
  INV_X1     g19599(.I(new_n19791_), .ZN(new_n19792_));
  NOR3_X1    g19600(.A1(new_n19148_), .A2(new_n19790_), .A3(new_n19792_), .ZN(new_n19793_));
  NAND2_X1   g19601(.A1(new_n19162_), .A2(new_n19793_), .ZN(new_n19794_));
  XOR2_X1    g19602(.A1(new_n19794_), .A2(\a[15] ), .Z(new_n19795_));
  INV_X1     g19603(.I(new_n19795_), .ZN(new_n19796_));
  NAND4_X1   g19604(.A1(new_n19781_), .A2(\a[15] ), .A3(new_n19779_), .A4(new_n19752_), .ZN(new_n19797_));
  INV_X1     g19605(.I(\a[15] ), .ZN(new_n19798_));
  NOR2_X1    g19606(.A1(new_n19798_), .A2(\a[14] ), .ZN(new_n19799_));
  INV_X1     g19607(.I(new_n19799_), .ZN(new_n19800_));
  AOI21_X1   g19608(.A1(new_n19797_), .A2(new_n19800_), .B(new_n19796_), .ZN(new_n19801_));
  NOR4_X1    g19609(.A1(new_n19768_), .A2(new_n19767_), .A3(new_n19798_), .A4(new_n19751_), .ZN(new_n19802_));
  NOR3_X1    g19610(.A1(new_n19802_), .A2(new_n19790_), .A3(new_n19795_), .ZN(new_n19803_));
  NOR2_X1    g19611(.A1(new_n19803_), .A2(new_n19801_), .ZN(new_n19804_));
  NAND4_X1   g19612(.A1(new_n19099_), .A2(new_n18888_), .A3(new_n19093_), .A4(new_n19161_), .ZN(new_n19805_));
  NOR2_X1    g19613(.A1(new_n19100_), .A2(new_n19790_), .ZN(new_n19806_));
  XOR2_X1    g19614(.A1(new_n19806_), .A2(new_n19805_), .Z(new_n19807_));
  NOR2_X1    g19615(.A1(new_n19807_), .A2(new_n19792_), .ZN(new_n19808_));
  NAND2_X1   g19616(.A1(new_n19757_), .A2(\asqrt[8] ), .ZN(new_n19809_));
  INV_X1     g19617(.I(new_n19809_), .ZN(new_n19810_));
  AOI21_X1   g19618(.A1(new_n19749_), .A2(new_n19810_), .B(\a[16] ), .ZN(new_n19811_));
  NOR3_X1    g19619(.A1(new_n19811_), .A2(new_n19118_), .A3(\asqrt[7] ), .ZN(new_n19812_));
  AOI21_X1   g19620(.A1(new_n19725_), .A2(new_n19727_), .B(new_n275_), .ZN(new_n19813_));
  OAI21_X1   g19621(.A1(new_n19728_), .A2(new_n19813_), .B(\asqrt[61] ), .ZN(new_n19814_));
  NOR4_X1    g19622(.A1(new_n19814_), .A2(new_n19551_), .A3(new_n19557_), .A4(new_n19742_), .ZN(new_n19815_));
  NOR3_X1    g19623(.A1(new_n19815_), .A2(new_n19562_), .A3(new_n19746_), .ZN(new_n19816_));
  OAI21_X1   g19624(.A1(new_n19816_), .A2(new_n19115_), .B(new_n19780_), .ZN(new_n19817_));
  OAI21_X1   g19625(.A1(new_n19817_), .A2(new_n19809_), .B(new_n19116_), .ZN(new_n19818_));
  AOI21_X1   g19626(.A1(new_n19818_), .A2(new_n19117_), .B(new_n19782_), .ZN(new_n19819_));
  NOR4_X1    g19627(.A1(new_n19819_), .A2(new_n19812_), .A3(\asqrt[9] ), .A4(new_n19808_), .ZN(new_n19820_));
  NOR2_X1    g19628(.A1(new_n19820_), .A2(new_n19804_), .ZN(new_n19821_));
  NOR3_X1    g19629(.A1(new_n19803_), .A2(new_n19801_), .A3(new_n19808_), .ZN(new_n19822_));
  INV_X1     g19630(.I(new_n19120_), .ZN(new_n19823_));
  NOR2_X1    g19631(.A1(new_n19100_), .A2(\a[16] ), .ZN(new_n19824_));
  OAI22_X1   g19632(.A1(new_n19824_), .A2(\a[17] ), .B1(\a[16] ), .B2(new_n19129_), .ZN(new_n19825_));
  NAND2_X1   g19633(.A1(\asqrt[8] ), .A2(\a[16] ), .ZN(new_n19826_));
  AND3_X2    g19634(.A1(new_n19825_), .A2(new_n19823_), .A3(new_n19826_), .Z(new_n19827_));
  INV_X1     g19635(.I(new_n19827_), .ZN(new_n19828_));
  NOR3_X1    g19636(.A1(new_n19782_), .A2(new_n19136_), .A3(new_n19828_), .ZN(new_n19829_));
  AOI21_X1   g19637(.A1(\asqrt[7] ), .A2(new_n19827_), .B(new_n19137_), .ZN(new_n19830_));
  NOR3_X1    g19638(.A1(new_n19830_), .A2(new_n19829_), .A3(\asqrt[10] ), .ZN(new_n19831_));
  OAI21_X1   g19639(.A1(new_n19822_), .A2(new_n18495_), .B(new_n19831_), .ZN(new_n19832_));
  NAND2_X1   g19640(.A1(new_n19821_), .A2(new_n19832_), .ZN(new_n19833_));
  OAI22_X1   g19641(.A1(new_n19820_), .A2(new_n19804_), .B1(new_n19822_), .B2(new_n18495_), .ZN(new_n19834_));
  INV_X1     g19642(.I(new_n19126_), .ZN(new_n19835_));
  AOI21_X1   g19643(.A1(new_n19129_), .A2(new_n19835_), .B(new_n19128_), .ZN(new_n19836_));
  INV_X1     g19644(.I(new_n19130_), .ZN(new_n19837_));
  NOR3_X1    g19645(.A1(new_n19837_), .A2(new_n19836_), .A3(new_n19136_), .ZN(new_n19838_));
  AOI21_X1   g19646(.A1(new_n19165_), .A2(new_n19151_), .B(\asqrt[10] ), .ZN(new_n19839_));
  AND4_X2    g19647(.A1(new_n19838_), .A2(\asqrt[7] ), .A3(new_n19179_), .A4(new_n19839_), .Z(new_n19840_));
  NOR2_X1    g19648(.A1(new_n19838_), .A2(new_n17893_), .ZN(new_n19841_));
  NOR3_X1    g19649(.A1(new_n19840_), .A2(\asqrt[11] ), .A3(new_n19841_), .ZN(new_n19842_));
  INV_X1     g19650(.I(new_n19842_), .ZN(new_n19843_));
  AOI21_X1   g19651(.A1(new_n19834_), .A2(\asqrt[10] ), .B(new_n19843_), .ZN(new_n19844_));
  NOR2_X1    g19652(.A1(new_n19844_), .A2(new_n19833_), .ZN(new_n19845_));
  AOI22_X1   g19653(.A1(new_n19834_), .A2(\asqrt[10] ), .B1(new_n19821_), .B2(new_n19832_), .ZN(new_n19846_));
  NAND2_X1   g19654(.A1(new_n19175_), .A2(new_n19174_), .ZN(new_n19847_));
  NAND4_X1   g19655(.A1(\asqrt[7] ), .A2(new_n17271_), .A3(new_n19847_), .A4(new_n19212_), .ZN(new_n19848_));
  XOR2_X1    g19656(.A1(new_n19848_), .A2(new_n19180_), .Z(new_n19849_));
  NAND2_X1   g19657(.A1(new_n19849_), .A2(new_n16619_), .ZN(new_n19850_));
  INV_X1     g19658(.I(new_n19850_), .ZN(new_n19851_));
  OAI21_X1   g19659(.A1(new_n19846_), .A2(new_n17271_), .B(new_n19851_), .ZN(new_n19852_));
  NAND2_X1   g19660(.A1(new_n19852_), .A2(new_n19845_), .ZN(new_n19853_));
  OAI22_X1   g19661(.A1(new_n19846_), .A2(new_n17271_), .B1(new_n19844_), .B2(new_n19833_), .ZN(new_n19854_));
  NOR2_X1    g19662(.A1(new_n19185_), .A2(new_n19186_), .ZN(new_n19855_));
  NOR4_X1    g19663(.A1(new_n19782_), .A2(\asqrt[12] ), .A3(new_n19855_), .A4(new_n19214_), .ZN(new_n19856_));
  XOR2_X1    g19664(.A1(new_n19856_), .A2(new_n19190_), .Z(new_n19857_));
  NAND2_X1   g19665(.A1(new_n19857_), .A2(new_n16060_), .ZN(new_n19858_));
  AOI21_X1   g19666(.A1(new_n19854_), .A2(\asqrt[12] ), .B(new_n19858_), .ZN(new_n19859_));
  NOR2_X1    g19667(.A1(new_n19859_), .A2(new_n19853_), .ZN(new_n19860_));
  AOI22_X1   g19668(.A1(new_n19854_), .A2(\asqrt[12] ), .B1(new_n19852_), .B2(new_n19845_), .ZN(new_n19861_));
  NOR2_X1    g19669(.A1(new_n19194_), .A2(\asqrt[13] ), .ZN(new_n19862_));
  NAND3_X1   g19670(.A1(\asqrt[7] ), .A2(new_n19215_), .A3(new_n19862_), .ZN(new_n19863_));
  XOR2_X1    g19671(.A1(new_n19863_), .A2(new_n19198_), .Z(new_n19864_));
  NAND2_X1   g19672(.A1(new_n19864_), .A2(new_n15447_), .ZN(new_n19865_));
  INV_X1     g19673(.I(new_n19865_), .ZN(new_n19866_));
  OAI21_X1   g19674(.A1(new_n19861_), .A2(new_n16060_), .B(new_n19866_), .ZN(new_n19867_));
  NAND2_X1   g19675(.A1(new_n19867_), .A2(new_n19860_), .ZN(new_n19868_));
  OAI22_X1   g19676(.A1(new_n19861_), .A2(new_n16060_), .B1(new_n19859_), .B2(new_n19853_), .ZN(new_n19869_));
  NOR4_X1    g19677(.A1(new_n19782_), .A2(\asqrt[14] ), .A3(new_n19202_), .A4(new_n19219_), .ZN(new_n19870_));
  XOR2_X1    g19678(.A1(new_n19870_), .A2(new_n19205_), .Z(new_n19871_));
  NAND2_X1   g19679(.A1(new_n19871_), .A2(new_n14871_), .ZN(new_n19872_));
  AOI21_X1   g19680(.A1(new_n19869_), .A2(\asqrt[14] ), .B(new_n19872_), .ZN(new_n19873_));
  NOR2_X1    g19681(.A1(new_n19873_), .A2(new_n19868_), .ZN(new_n19874_));
  AOI22_X1   g19682(.A1(new_n19869_), .A2(\asqrt[14] ), .B1(new_n19867_), .B2(new_n19860_), .ZN(new_n19875_));
  NOR4_X1    g19683(.A1(new_n19782_), .A2(\asqrt[15] ), .A3(new_n19208_), .A4(new_n19568_), .ZN(new_n19876_));
  XNOR2_X1   g19684(.A1(new_n19876_), .A2(new_n19571_), .ZN(new_n19877_));
  NAND2_X1   g19685(.A1(new_n19877_), .A2(new_n14273_), .ZN(new_n19878_));
  INV_X1     g19686(.I(new_n19878_), .ZN(new_n19879_));
  OAI21_X1   g19687(.A1(new_n19875_), .A2(new_n14871_), .B(new_n19879_), .ZN(new_n19880_));
  NAND2_X1   g19688(.A1(new_n19880_), .A2(new_n19874_), .ZN(new_n19881_));
  OAI22_X1   g19689(.A1(new_n19875_), .A2(new_n14871_), .B1(new_n19873_), .B2(new_n19868_), .ZN(new_n19882_));
  NOR4_X1    g19690(.A1(new_n19782_), .A2(\asqrt[16] ), .A3(new_n19223_), .A4(new_n19229_), .ZN(new_n19883_));
  XOR2_X1    g19691(.A1(new_n19883_), .A2(new_n19572_), .Z(new_n19884_));
  NAND2_X1   g19692(.A1(new_n19884_), .A2(new_n13760_), .ZN(new_n19885_));
  AOI21_X1   g19693(.A1(new_n19882_), .A2(\asqrt[16] ), .B(new_n19885_), .ZN(new_n19886_));
  NOR2_X1    g19694(.A1(new_n19886_), .A2(new_n19881_), .ZN(new_n19887_));
  AOI22_X1   g19695(.A1(new_n19882_), .A2(\asqrt[16] ), .B1(new_n19880_), .B2(new_n19874_), .ZN(new_n19888_));
  NAND2_X1   g19696(.A1(new_n19577_), .A2(\asqrt[17] ), .ZN(new_n19889_));
  NOR4_X1    g19697(.A1(new_n19782_), .A2(\asqrt[17] ), .A3(new_n19232_), .A4(new_n19577_), .ZN(new_n19890_));
  XOR2_X1    g19698(.A1(new_n19890_), .A2(new_n19889_), .Z(new_n19891_));
  NAND2_X1   g19699(.A1(new_n19891_), .A2(new_n13192_), .ZN(new_n19892_));
  INV_X1     g19700(.I(new_n19892_), .ZN(new_n19893_));
  OAI21_X1   g19701(.A1(new_n19888_), .A2(new_n13760_), .B(new_n19893_), .ZN(new_n19894_));
  NAND2_X1   g19702(.A1(new_n19894_), .A2(new_n19887_), .ZN(new_n19895_));
  OAI22_X1   g19703(.A1(new_n19888_), .A2(new_n13760_), .B1(new_n19886_), .B2(new_n19881_), .ZN(new_n19896_));
  NOR4_X1    g19704(.A1(new_n19782_), .A2(\asqrt[18] ), .A3(new_n19239_), .A4(new_n19244_), .ZN(new_n19897_));
  AOI21_X1   g19705(.A1(new_n19889_), .A2(new_n19575_), .B(new_n13192_), .ZN(new_n19898_));
  NOR2_X1    g19706(.A1(new_n19897_), .A2(new_n19898_), .ZN(new_n19899_));
  NAND2_X1   g19707(.A1(new_n19899_), .A2(new_n12657_), .ZN(new_n19900_));
  AOI21_X1   g19708(.A1(new_n19896_), .A2(\asqrt[18] ), .B(new_n19900_), .ZN(new_n19901_));
  NOR2_X1    g19709(.A1(new_n19901_), .A2(new_n19895_), .ZN(new_n19902_));
  AOI22_X1   g19710(.A1(new_n19896_), .A2(\asqrt[18] ), .B1(new_n19894_), .B2(new_n19887_), .ZN(new_n19903_));
  NAND2_X1   g19711(.A1(new_n19584_), .A2(\asqrt[19] ), .ZN(new_n19904_));
  NOR4_X1    g19712(.A1(new_n19782_), .A2(\asqrt[19] ), .A3(new_n19247_), .A4(new_n19584_), .ZN(new_n19905_));
  XOR2_X1    g19713(.A1(new_n19905_), .A2(new_n19904_), .Z(new_n19906_));
  NAND2_X1   g19714(.A1(new_n19906_), .A2(new_n12101_), .ZN(new_n19907_));
  INV_X1     g19715(.I(new_n19907_), .ZN(new_n19908_));
  OAI21_X1   g19716(.A1(new_n19903_), .A2(new_n12657_), .B(new_n19908_), .ZN(new_n19909_));
  NAND2_X1   g19717(.A1(new_n19909_), .A2(new_n19902_), .ZN(new_n19910_));
  OAI22_X1   g19718(.A1(new_n19903_), .A2(new_n12657_), .B1(new_n19901_), .B2(new_n19895_), .ZN(new_n19911_));
  NOR4_X1    g19719(.A1(new_n19782_), .A2(\asqrt[20] ), .A3(new_n19254_), .A4(new_n19259_), .ZN(new_n19912_));
  AOI21_X1   g19720(.A1(new_n19904_), .A2(new_n19583_), .B(new_n12101_), .ZN(new_n19913_));
  NOR2_X1    g19721(.A1(new_n19912_), .A2(new_n19913_), .ZN(new_n19914_));
  NAND2_X1   g19722(.A1(new_n19914_), .A2(new_n11631_), .ZN(new_n19915_));
  AOI21_X1   g19723(.A1(new_n19911_), .A2(\asqrt[20] ), .B(new_n19915_), .ZN(new_n19916_));
  NOR2_X1    g19724(.A1(new_n19916_), .A2(new_n19910_), .ZN(new_n19917_));
  AOI22_X1   g19725(.A1(new_n19911_), .A2(\asqrt[20] ), .B1(new_n19909_), .B2(new_n19902_), .ZN(new_n19918_));
  NAND2_X1   g19726(.A1(new_n19591_), .A2(\asqrt[21] ), .ZN(new_n19919_));
  NOR4_X1    g19727(.A1(new_n19782_), .A2(\asqrt[21] ), .A3(new_n19262_), .A4(new_n19591_), .ZN(new_n19920_));
  XOR2_X1    g19728(.A1(new_n19920_), .A2(new_n19919_), .Z(new_n19921_));
  NAND2_X1   g19729(.A1(new_n19921_), .A2(new_n11105_), .ZN(new_n19922_));
  INV_X1     g19730(.I(new_n19922_), .ZN(new_n19923_));
  OAI21_X1   g19731(.A1(new_n19918_), .A2(new_n11631_), .B(new_n19923_), .ZN(new_n19924_));
  NAND2_X1   g19732(.A1(new_n19924_), .A2(new_n19917_), .ZN(new_n19925_));
  OAI22_X1   g19733(.A1(new_n19918_), .A2(new_n11631_), .B1(new_n19916_), .B2(new_n19910_), .ZN(new_n19926_));
  NOR4_X1    g19734(.A1(new_n19782_), .A2(\asqrt[22] ), .A3(new_n19269_), .A4(new_n19274_), .ZN(new_n19927_));
  AOI21_X1   g19735(.A1(new_n19919_), .A2(new_n19590_), .B(new_n11105_), .ZN(new_n19928_));
  NOR2_X1    g19736(.A1(new_n19927_), .A2(new_n19928_), .ZN(new_n19929_));
  NAND2_X1   g19737(.A1(new_n19929_), .A2(new_n10614_), .ZN(new_n19930_));
  AOI21_X1   g19738(.A1(new_n19926_), .A2(\asqrt[22] ), .B(new_n19930_), .ZN(new_n19931_));
  NOR2_X1    g19739(.A1(new_n19931_), .A2(new_n19925_), .ZN(new_n19932_));
  AOI22_X1   g19740(.A1(new_n19926_), .A2(\asqrt[22] ), .B1(new_n19924_), .B2(new_n19917_), .ZN(new_n19933_));
  NAND2_X1   g19741(.A1(new_n19598_), .A2(\asqrt[23] ), .ZN(new_n19934_));
  NOR4_X1    g19742(.A1(new_n19782_), .A2(\asqrt[23] ), .A3(new_n19277_), .A4(new_n19598_), .ZN(new_n19935_));
  XOR2_X1    g19743(.A1(new_n19935_), .A2(new_n19934_), .Z(new_n19936_));
  NAND2_X1   g19744(.A1(new_n19936_), .A2(new_n10104_), .ZN(new_n19937_));
  INV_X1     g19745(.I(new_n19937_), .ZN(new_n19938_));
  OAI21_X1   g19746(.A1(new_n19933_), .A2(new_n10614_), .B(new_n19938_), .ZN(new_n19939_));
  NAND2_X1   g19747(.A1(new_n19939_), .A2(new_n19932_), .ZN(new_n19940_));
  OAI22_X1   g19748(.A1(new_n19933_), .A2(new_n10614_), .B1(new_n19931_), .B2(new_n19925_), .ZN(new_n19941_));
  NOR4_X1    g19749(.A1(new_n19782_), .A2(\asqrt[24] ), .A3(new_n19284_), .A4(new_n19289_), .ZN(new_n19942_));
  AOI21_X1   g19750(.A1(new_n19934_), .A2(new_n19597_), .B(new_n10104_), .ZN(new_n19943_));
  NOR2_X1    g19751(.A1(new_n19942_), .A2(new_n19943_), .ZN(new_n19944_));
  NAND2_X1   g19752(.A1(new_n19944_), .A2(new_n9672_), .ZN(new_n19945_));
  AOI21_X1   g19753(.A1(new_n19941_), .A2(\asqrt[24] ), .B(new_n19945_), .ZN(new_n19946_));
  NOR2_X1    g19754(.A1(new_n19946_), .A2(new_n19940_), .ZN(new_n19947_));
  AOI22_X1   g19755(.A1(new_n19941_), .A2(\asqrt[24] ), .B1(new_n19939_), .B2(new_n19932_), .ZN(new_n19948_));
  NAND2_X1   g19756(.A1(new_n19605_), .A2(\asqrt[25] ), .ZN(new_n19949_));
  NOR4_X1    g19757(.A1(new_n19782_), .A2(\asqrt[25] ), .A3(new_n19292_), .A4(new_n19605_), .ZN(new_n19950_));
  XOR2_X1    g19758(.A1(new_n19950_), .A2(new_n19949_), .Z(new_n19951_));
  NAND2_X1   g19759(.A1(new_n19951_), .A2(new_n9212_), .ZN(new_n19952_));
  INV_X1     g19760(.I(new_n19952_), .ZN(new_n19953_));
  OAI21_X1   g19761(.A1(new_n19948_), .A2(new_n9672_), .B(new_n19953_), .ZN(new_n19954_));
  NAND2_X1   g19762(.A1(new_n19954_), .A2(new_n19947_), .ZN(new_n19955_));
  OAI22_X1   g19763(.A1(new_n19948_), .A2(new_n9672_), .B1(new_n19946_), .B2(new_n19940_), .ZN(new_n19956_));
  NOR4_X1    g19764(.A1(new_n19782_), .A2(\asqrt[26] ), .A3(new_n19299_), .A4(new_n19304_), .ZN(new_n19957_));
  AOI21_X1   g19765(.A1(new_n19949_), .A2(new_n19604_), .B(new_n9212_), .ZN(new_n19958_));
  NOR2_X1    g19766(.A1(new_n19957_), .A2(new_n19958_), .ZN(new_n19959_));
  NAND2_X1   g19767(.A1(new_n19959_), .A2(new_n8763_), .ZN(new_n19960_));
  AOI21_X1   g19768(.A1(new_n19956_), .A2(\asqrt[26] ), .B(new_n19960_), .ZN(new_n19961_));
  NOR2_X1    g19769(.A1(new_n19961_), .A2(new_n19955_), .ZN(new_n19962_));
  AOI22_X1   g19770(.A1(new_n19956_), .A2(\asqrt[26] ), .B1(new_n19954_), .B2(new_n19947_), .ZN(new_n19963_));
  NAND2_X1   g19771(.A1(new_n19612_), .A2(\asqrt[27] ), .ZN(new_n19964_));
  NOR4_X1    g19772(.A1(new_n19782_), .A2(\asqrt[27] ), .A3(new_n19307_), .A4(new_n19612_), .ZN(new_n19965_));
  XOR2_X1    g19773(.A1(new_n19965_), .A2(new_n19964_), .Z(new_n19966_));
  NAND2_X1   g19774(.A1(new_n19966_), .A2(new_n8319_), .ZN(new_n19967_));
  INV_X1     g19775(.I(new_n19967_), .ZN(new_n19968_));
  OAI21_X1   g19776(.A1(new_n19963_), .A2(new_n8763_), .B(new_n19968_), .ZN(new_n19969_));
  NAND2_X1   g19777(.A1(new_n19969_), .A2(new_n19962_), .ZN(new_n19970_));
  OAI22_X1   g19778(.A1(new_n19963_), .A2(new_n8763_), .B1(new_n19961_), .B2(new_n19955_), .ZN(new_n19971_));
  NOR4_X1    g19779(.A1(new_n19782_), .A2(\asqrt[28] ), .A3(new_n19314_), .A4(new_n19319_), .ZN(new_n19972_));
  AOI21_X1   g19780(.A1(new_n19964_), .A2(new_n19611_), .B(new_n8319_), .ZN(new_n19973_));
  NOR2_X1    g19781(.A1(new_n19972_), .A2(new_n19973_), .ZN(new_n19974_));
  NAND2_X1   g19782(.A1(new_n19974_), .A2(new_n7931_), .ZN(new_n19975_));
  AOI21_X1   g19783(.A1(new_n19971_), .A2(\asqrt[28] ), .B(new_n19975_), .ZN(new_n19976_));
  NOR2_X1    g19784(.A1(new_n19976_), .A2(new_n19970_), .ZN(new_n19977_));
  AOI22_X1   g19785(.A1(new_n19971_), .A2(\asqrt[28] ), .B1(new_n19969_), .B2(new_n19962_), .ZN(new_n19978_));
  NAND2_X1   g19786(.A1(new_n19619_), .A2(\asqrt[29] ), .ZN(new_n19979_));
  NOR4_X1    g19787(.A1(new_n19782_), .A2(\asqrt[29] ), .A3(new_n19322_), .A4(new_n19619_), .ZN(new_n19980_));
  XOR2_X1    g19788(.A1(new_n19980_), .A2(new_n19979_), .Z(new_n19981_));
  NAND2_X1   g19789(.A1(new_n19981_), .A2(new_n7517_), .ZN(new_n19982_));
  INV_X1     g19790(.I(new_n19982_), .ZN(new_n19983_));
  OAI21_X1   g19791(.A1(new_n19978_), .A2(new_n7931_), .B(new_n19983_), .ZN(new_n19984_));
  NAND2_X1   g19792(.A1(new_n19984_), .A2(new_n19977_), .ZN(new_n19985_));
  OAI22_X1   g19793(.A1(new_n19978_), .A2(new_n7931_), .B1(new_n19976_), .B2(new_n19970_), .ZN(new_n19986_));
  NAND2_X1   g19794(.A1(new_n19334_), .A2(\asqrt[30] ), .ZN(new_n19987_));
  NOR4_X1    g19795(.A1(new_n19782_), .A2(\asqrt[30] ), .A3(new_n19329_), .A4(new_n19334_), .ZN(new_n19988_));
  XOR2_X1    g19796(.A1(new_n19988_), .A2(new_n19987_), .Z(new_n19989_));
  NAND2_X1   g19797(.A1(new_n19989_), .A2(new_n7110_), .ZN(new_n19990_));
  AOI21_X1   g19798(.A1(new_n19986_), .A2(\asqrt[30] ), .B(new_n19990_), .ZN(new_n19991_));
  NOR2_X1    g19799(.A1(new_n19991_), .A2(new_n19985_), .ZN(new_n19992_));
  AOI22_X1   g19800(.A1(new_n19986_), .A2(\asqrt[30] ), .B1(new_n19984_), .B2(new_n19977_), .ZN(new_n19993_));
  NOR4_X1    g19801(.A1(new_n19782_), .A2(\asqrt[31] ), .A3(new_n19337_), .A4(new_n19626_), .ZN(new_n19994_));
  AOI21_X1   g19802(.A1(new_n19987_), .A2(new_n19333_), .B(new_n7110_), .ZN(new_n19995_));
  NOR2_X1    g19803(.A1(new_n19994_), .A2(new_n19995_), .ZN(new_n19996_));
  NAND2_X1   g19804(.A1(new_n19996_), .A2(new_n6708_), .ZN(new_n19997_));
  INV_X1     g19805(.I(new_n19997_), .ZN(new_n19998_));
  OAI21_X1   g19806(.A1(new_n19993_), .A2(new_n7110_), .B(new_n19998_), .ZN(new_n19999_));
  NAND2_X1   g19807(.A1(new_n19999_), .A2(new_n19992_), .ZN(new_n20000_));
  OAI22_X1   g19808(.A1(new_n19993_), .A2(new_n7110_), .B1(new_n19991_), .B2(new_n19985_), .ZN(new_n20001_));
  NAND2_X1   g19809(.A1(new_n19349_), .A2(\asqrt[32] ), .ZN(new_n20002_));
  NOR4_X1    g19810(.A1(new_n19782_), .A2(\asqrt[32] ), .A3(new_n19344_), .A4(new_n19349_), .ZN(new_n20003_));
  XOR2_X1    g19811(.A1(new_n20003_), .A2(new_n20002_), .Z(new_n20004_));
  NAND2_X1   g19812(.A1(new_n20004_), .A2(new_n6365_), .ZN(new_n20005_));
  AOI21_X1   g19813(.A1(new_n20001_), .A2(\asqrt[32] ), .B(new_n20005_), .ZN(new_n20006_));
  NOR2_X1    g19814(.A1(new_n20006_), .A2(new_n20000_), .ZN(new_n20007_));
  AOI22_X1   g19815(.A1(new_n20001_), .A2(\asqrt[32] ), .B1(new_n19999_), .B2(new_n19992_), .ZN(new_n20008_));
  NAND2_X1   g19816(.A1(new_n19633_), .A2(\asqrt[33] ), .ZN(new_n20009_));
  NOR4_X1    g19817(.A1(new_n19782_), .A2(\asqrt[33] ), .A3(new_n19352_), .A4(new_n19633_), .ZN(new_n20010_));
  XOR2_X1    g19818(.A1(new_n20010_), .A2(new_n20009_), .Z(new_n20011_));
  NAND2_X1   g19819(.A1(new_n20011_), .A2(new_n5991_), .ZN(new_n20012_));
  INV_X1     g19820(.I(new_n20012_), .ZN(new_n20013_));
  OAI21_X1   g19821(.A1(new_n20008_), .A2(new_n6365_), .B(new_n20013_), .ZN(new_n20014_));
  NAND2_X1   g19822(.A1(new_n20014_), .A2(new_n20007_), .ZN(new_n20015_));
  OAI22_X1   g19823(.A1(new_n20008_), .A2(new_n6365_), .B1(new_n20006_), .B2(new_n20000_), .ZN(new_n20016_));
  NOR4_X1    g19824(.A1(new_n19782_), .A2(\asqrt[34] ), .A3(new_n19359_), .A4(new_n19364_), .ZN(new_n20017_));
  AOI21_X1   g19825(.A1(new_n20009_), .A2(new_n19632_), .B(new_n5991_), .ZN(new_n20018_));
  NOR2_X1    g19826(.A1(new_n20017_), .A2(new_n20018_), .ZN(new_n20019_));
  NAND2_X1   g19827(.A1(new_n20019_), .A2(new_n5626_), .ZN(new_n20020_));
  AOI21_X1   g19828(.A1(new_n20016_), .A2(\asqrt[34] ), .B(new_n20020_), .ZN(new_n20021_));
  NOR2_X1    g19829(.A1(new_n20021_), .A2(new_n20015_), .ZN(new_n20022_));
  AOI22_X1   g19830(.A1(new_n20016_), .A2(\asqrt[34] ), .B1(new_n20014_), .B2(new_n20007_), .ZN(new_n20023_));
  NAND2_X1   g19831(.A1(new_n19640_), .A2(\asqrt[35] ), .ZN(new_n20024_));
  NOR4_X1    g19832(.A1(new_n19782_), .A2(\asqrt[35] ), .A3(new_n19367_), .A4(new_n19640_), .ZN(new_n20025_));
  XOR2_X1    g19833(.A1(new_n20025_), .A2(new_n20024_), .Z(new_n20026_));
  NAND2_X1   g19834(.A1(new_n20026_), .A2(new_n5273_), .ZN(new_n20027_));
  INV_X1     g19835(.I(new_n20027_), .ZN(new_n20028_));
  OAI21_X1   g19836(.A1(new_n20023_), .A2(new_n5626_), .B(new_n20028_), .ZN(new_n20029_));
  NAND2_X1   g19837(.A1(new_n20029_), .A2(new_n20022_), .ZN(new_n20030_));
  OAI22_X1   g19838(.A1(new_n20023_), .A2(new_n5626_), .B1(new_n20021_), .B2(new_n20015_), .ZN(new_n20031_));
  NOR4_X1    g19839(.A1(new_n19782_), .A2(\asqrt[36] ), .A3(new_n19374_), .A4(new_n19379_), .ZN(new_n20032_));
  AOI21_X1   g19840(.A1(new_n20024_), .A2(new_n19639_), .B(new_n5273_), .ZN(new_n20033_));
  NOR2_X1    g19841(.A1(new_n20032_), .A2(new_n20033_), .ZN(new_n20034_));
  NAND2_X1   g19842(.A1(new_n20034_), .A2(new_n4973_), .ZN(new_n20035_));
  AOI21_X1   g19843(.A1(new_n20031_), .A2(\asqrt[36] ), .B(new_n20035_), .ZN(new_n20036_));
  NOR2_X1    g19844(.A1(new_n20036_), .A2(new_n20030_), .ZN(new_n20037_));
  AOI22_X1   g19845(.A1(new_n20031_), .A2(\asqrt[36] ), .B1(new_n20029_), .B2(new_n20022_), .ZN(new_n20038_));
  NAND2_X1   g19846(.A1(new_n19647_), .A2(\asqrt[37] ), .ZN(new_n20039_));
  NOR4_X1    g19847(.A1(new_n19782_), .A2(\asqrt[37] ), .A3(new_n19382_), .A4(new_n19647_), .ZN(new_n20040_));
  XOR2_X1    g19848(.A1(new_n20040_), .A2(new_n20039_), .Z(new_n20041_));
  NAND2_X1   g19849(.A1(new_n20041_), .A2(new_n4645_), .ZN(new_n20042_));
  INV_X1     g19850(.I(new_n20042_), .ZN(new_n20043_));
  OAI21_X1   g19851(.A1(new_n20038_), .A2(new_n4973_), .B(new_n20043_), .ZN(new_n20044_));
  NAND2_X1   g19852(.A1(new_n20044_), .A2(new_n20037_), .ZN(new_n20045_));
  OAI22_X1   g19853(.A1(new_n20038_), .A2(new_n4973_), .B1(new_n20036_), .B2(new_n20030_), .ZN(new_n20046_));
  NOR4_X1    g19854(.A1(new_n19782_), .A2(\asqrt[38] ), .A3(new_n19389_), .A4(new_n19394_), .ZN(new_n20047_));
  AOI21_X1   g19855(.A1(new_n20039_), .A2(new_n19646_), .B(new_n4645_), .ZN(new_n20048_));
  NOR2_X1    g19856(.A1(new_n20047_), .A2(new_n20048_), .ZN(new_n20049_));
  NAND2_X1   g19857(.A1(new_n20049_), .A2(new_n4330_), .ZN(new_n20050_));
  AOI21_X1   g19858(.A1(new_n20046_), .A2(\asqrt[38] ), .B(new_n20050_), .ZN(new_n20051_));
  NOR2_X1    g19859(.A1(new_n20051_), .A2(new_n20045_), .ZN(new_n20052_));
  AOI22_X1   g19860(.A1(new_n20046_), .A2(\asqrt[38] ), .B1(new_n20044_), .B2(new_n20037_), .ZN(new_n20053_));
  NAND2_X1   g19861(.A1(new_n19654_), .A2(\asqrt[39] ), .ZN(new_n20054_));
  NOR4_X1    g19862(.A1(new_n19782_), .A2(\asqrt[39] ), .A3(new_n19397_), .A4(new_n19654_), .ZN(new_n20055_));
  XOR2_X1    g19863(.A1(new_n20055_), .A2(new_n20054_), .Z(new_n20056_));
  NAND2_X1   g19864(.A1(new_n20056_), .A2(new_n4018_), .ZN(new_n20057_));
  INV_X1     g19865(.I(new_n20057_), .ZN(new_n20058_));
  OAI21_X1   g19866(.A1(new_n20053_), .A2(new_n4330_), .B(new_n20058_), .ZN(new_n20059_));
  NAND2_X1   g19867(.A1(new_n20059_), .A2(new_n20052_), .ZN(new_n20060_));
  OAI22_X1   g19868(.A1(new_n20053_), .A2(new_n4330_), .B1(new_n20051_), .B2(new_n20045_), .ZN(new_n20061_));
  NOR4_X1    g19869(.A1(new_n19782_), .A2(\asqrt[40] ), .A3(new_n19404_), .A4(new_n19409_), .ZN(new_n20062_));
  AOI21_X1   g19870(.A1(new_n20054_), .A2(new_n19653_), .B(new_n4018_), .ZN(new_n20063_));
  NOR2_X1    g19871(.A1(new_n20062_), .A2(new_n20063_), .ZN(new_n20064_));
  NAND2_X1   g19872(.A1(new_n20064_), .A2(new_n3760_), .ZN(new_n20065_));
  AOI21_X1   g19873(.A1(new_n20061_), .A2(\asqrt[40] ), .B(new_n20065_), .ZN(new_n20066_));
  NOR2_X1    g19874(.A1(new_n20066_), .A2(new_n20060_), .ZN(new_n20067_));
  AOI22_X1   g19875(.A1(new_n20061_), .A2(\asqrt[40] ), .B1(new_n20059_), .B2(new_n20052_), .ZN(new_n20068_));
  NAND2_X1   g19876(.A1(new_n19661_), .A2(\asqrt[41] ), .ZN(new_n20069_));
  NOR4_X1    g19877(.A1(new_n19782_), .A2(\asqrt[41] ), .A3(new_n19412_), .A4(new_n19661_), .ZN(new_n20070_));
  XOR2_X1    g19878(.A1(new_n20070_), .A2(new_n20069_), .Z(new_n20071_));
  NAND2_X1   g19879(.A1(new_n20071_), .A2(new_n3481_), .ZN(new_n20072_));
  INV_X1     g19880(.I(new_n20072_), .ZN(new_n20073_));
  OAI21_X1   g19881(.A1(new_n20068_), .A2(new_n3760_), .B(new_n20073_), .ZN(new_n20074_));
  NAND2_X1   g19882(.A1(new_n20074_), .A2(new_n20067_), .ZN(new_n20075_));
  OAI22_X1   g19883(.A1(new_n20068_), .A2(new_n3760_), .B1(new_n20066_), .B2(new_n20060_), .ZN(new_n20076_));
  NAND2_X1   g19884(.A1(new_n19424_), .A2(\asqrt[42] ), .ZN(new_n20077_));
  NOR4_X1    g19885(.A1(new_n19782_), .A2(\asqrt[42] ), .A3(new_n19419_), .A4(new_n19424_), .ZN(new_n20078_));
  XOR2_X1    g19886(.A1(new_n20078_), .A2(new_n20077_), .Z(new_n20079_));
  NAND2_X1   g19887(.A1(new_n20079_), .A2(new_n3208_), .ZN(new_n20080_));
  AOI21_X1   g19888(.A1(new_n20076_), .A2(\asqrt[42] ), .B(new_n20080_), .ZN(new_n20081_));
  NOR2_X1    g19889(.A1(new_n20081_), .A2(new_n20075_), .ZN(new_n20082_));
  AOI22_X1   g19890(.A1(new_n20076_), .A2(\asqrt[42] ), .B1(new_n20074_), .B2(new_n20067_), .ZN(new_n20083_));
  NOR4_X1    g19891(.A1(new_n19782_), .A2(\asqrt[43] ), .A3(new_n19427_), .A4(new_n19668_), .ZN(new_n20084_));
  AOI21_X1   g19892(.A1(new_n20077_), .A2(new_n19423_), .B(new_n3208_), .ZN(new_n20085_));
  NOR2_X1    g19893(.A1(new_n20084_), .A2(new_n20085_), .ZN(new_n20086_));
  NAND2_X1   g19894(.A1(new_n20086_), .A2(new_n2941_), .ZN(new_n20087_));
  INV_X1     g19895(.I(new_n20087_), .ZN(new_n20088_));
  OAI21_X1   g19896(.A1(new_n20083_), .A2(new_n3208_), .B(new_n20088_), .ZN(new_n20089_));
  NAND2_X1   g19897(.A1(new_n20089_), .A2(new_n20082_), .ZN(new_n20090_));
  OAI22_X1   g19898(.A1(new_n20083_), .A2(new_n3208_), .B1(new_n20081_), .B2(new_n20075_), .ZN(new_n20091_));
  NAND2_X1   g19899(.A1(new_n19439_), .A2(\asqrt[44] ), .ZN(new_n20092_));
  NOR4_X1    g19900(.A1(new_n19782_), .A2(\asqrt[44] ), .A3(new_n19434_), .A4(new_n19439_), .ZN(new_n20093_));
  XOR2_X1    g19901(.A1(new_n20093_), .A2(new_n20092_), .Z(new_n20094_));
  NAND2_X1   g19902(.A1(new_n20094_), .A2(new_n2728_), .ZN(new_n20095_));
  AOI21_X1   g19903(.A1(new_n20091_), .A2(\asqrt[44] ), .B(new_n20095_), .ZN(new_n20096_));
  NOR2_X1    g19904(.A1(new_n20096_), .A2(new_n20090_), .ZN(new_n20097_));
  AOI22_X1   g19905(.A1(new_n20091_), .A2(\asqrt[44] ), .B1(new_n20089_), .B2(new_n20082_), .ZN(new_n20098_));
  NAND2_X1   g19906(.A1(new_n19675_), .A2(\asqrt[45] ), .ZN(new_n20099_));
  NOR4_X1    g19907(.A1(new_n19782_), .A2(\asqrt[45] ), .A3(new_n19442_), .A4(new_n19675_), .ZN(new_n20100_));
  XOR2_X1    g19908(.A1(new_n20100_), .A2(new_n20099_), .Z(new_n20101_));
  NAND2_X1   g19909(.A1(new_n20101_), .A2(new_n2488_), .ZN(new_n20102_));
  INV_X1     g19910(.I(new_n20102_), .ZN(new_n20103_));
  OAI21_X1   g19911(.A1(new_n20098_), .A2(new_n2728_), .B(new_n20103_), .ZN(new_n20104_));
  NAND2_X1   g19912(.A1(new_n20104_), .A2(new_n20097_), .ZN(new_n20105_));
  OAI22_X1   g19913(.A1(new_n20098_), .A2(new_n2728_), .B1(new_n20096_), .B2(new_n20090_), .ZN(new_n20106_));
  NOR4_X1    g19914(.A1(new_n19782_), .A2(\asqrt[46] ), .A3(new_n19449_), .A4(new_n19454_), .ZN(new_n20107_));
  AOI21_X1   g19915(.A1(new_n20099_), .A2(new_n19674_), .B(new_n2488_), .ZN(new_n20108_));
  NOR2_X1    g19916(.A1(new_n20107_), .A2(new_n20108_), .ZN(new_n20109_));
  NAND2_X1   g19917(.A1(new_n20109_), .A2(new_n2253_), .ZN(new_n20110_));
  AOI21_X1   g19918(.A1(new_n20106_), .A2(\asqrt[46] ), .B(new_n20110_), .ZN(new_n20111_));
  NOR2_X1    g19919(.A1(new_n20111_), .A2(new_n20105_), .ZN(new_n20112_));
  AOI22_X1   g19920(.A1(new_n20106_), .A2(\asqrt[46] ), .B1(new_n20104_), .B2(new_n20097_), .ZN(new_n20113_));
  NAND2_X1   g19921(.A1(new_n19682_), .A2(\asqrt[47] ), .ZN(new_n20114_));
  NOR4_X1    g19922(.A1(new_n19782_), .A2(\asqrt[47] ), .A3(new_n19457_), .A4(new_n19682_), .ZN(new_n20115_));
  XOR2_X1    g19923(.A1(new_n20115_), .A2(new_n20114_), .Z(new_n20116_));
  NAND2_X1   g19924(.A1(new_n20116_), .A2(new_n2046_), .ZN(new_n20117_));
  INV_X1     g19925(.I(new_n20117_), .ZN(new_n20118_));
  OAI21_X1   g19926(.A1(new_n20113_), .A2(new_n2253_), .B(new_n20118_), .ZN(new_n20119_));
  NAND2_X1   g19927(.A1(new_n20119_), .A2(new_n20112_), .ZN(new_n20120_));
  OAI22_X1   g19928(.A1(new_n20113_), .A2(new_n2253_), .B1(new_n20111_), .B2(new_n20105_), .ZN(new_n20121_));
  NOR4_X1    g19929(.A1(new_n19782_), .A2(\asqrt[48] ), .A3(new_n19464_), .A4(new_n19469_), .ZN(new_n20122_));
  AOI21_X1   g19930(.A1(new_n20114_), .A2(new_n19681_), .B(new_n2046_), .ZN(new_n20123_));
  NOR2_X1    g19931(.A1(new_n20122_), .A2(new_n20123_), .ZN(new_n20124_));
  NAND2_X1   g19932(.A1(new_n20124_), .A2(new_n1854_), .ZN(new_n20125_));
  AOI21_X1   g19933(.A1(new_n20121_), .A2(\asqrt[48] ), .B(new_n20125_), .ZN(new_n20126_));
  NOR2_X1    g19934(.A1(new_n20126_), .A2(new_n20120_), .ZN(new_n20127_));
  AOI22_X1   g19935(.A1(new_n20121_), .A2(\asqrt[48] ), .B1(new_n20119_), .B2(new_n20112_), .ZN(new_n20128_));
  NAND2_X1   g19936(.A1(new_n19689_), .A2(\asqrt[49] ), .ZN(new_n20129_));
  NOR4_X1    g19937(.A1(new_n19782_), .A2(\asqrt[49] ), .A3(new_n19472_), .A4(new_n19689_), .ZN(new_n20130_));
  XOR2_X1    g19938(.A1(new_n20130_), .A2(new_n20129_), .Z(new_n20131_));
  NAND2_X1   g19939(.A1(new_n20131_), .A2(new_n1595_), .ZN(new_n20132_));
  INV_X1     g19940(.I(new_n20132_), .ZN(new_n20133_));
  OAI21_X1   g19941(.A1(new_n20128_), .A2(new_n1854_), .B(new_n20133_), .ZN(new_n20134_));
  NAND2_X1   g19942(.A1(new_n20134_), .A2(new_n20127_), .ZN(new_n20135_));
  OAI22_X1   g19943(.A1(new_n20128_), .A2(new_n1854_), .B1(new_n20126_), .B2(new_n20120_), .ZN(new_n20136_));
  NOR4_X1    g19944(.A1(new_n19782_), .A2(\asqrt[50] ), .A3(new_n19479_), .A4(new_n19484_), .ZN(new_n20137_));
  AOI21_X1   g19945(.A1(new_n20129_), .A2(new_n19688_), .B(new_n1595_), .ZN(new_n20138_));
  NOR2_X1    g19946(.A1(new_n20137_), .A2(new_n20138_), .ZN(new_n20139_));
  NAND2_X1   g19947(.A1(new_n20139_), .A2(new_n1436_), .ZN(new_n20140_));
  AOI21_X1   g19948(.A1(new_n20136_), .A2(\asqrt[50] ), .B(new_n20140_), .ZN(new_n20141_));
  NOR2_X1    g19949(.A1(new_n20141_), .A2(new_n20135_), .ZN(new_n20142_));
  AOI22_X1   g19950(.A1(new_n20136_), .A2(\asqrt[50] ), .B1(new_n20134_), .B2(new_n20127_), .ZN(new_n20143_));
  NAND2_X1   g19951(.A1(new_n19696_), .A2(\asqrt[51] ), .ZN(new_n20144_));
  NOR4_X1    g19952(.A1(new_n19782_), .A2(\asqrt[51] ), .A3(new_n19487_), .A4(new_n19696_), .ZN(new_n20145_));
  XOR2_X1    g19953(.A1(new_n20145_), .A2(new_n20144_), .Z(new_n20146_));
  NAND2_X1   g19954(.A1(new_n20146_), .A2(new_n1260_), .ZN(new_n20147_));
  INV_X1     g19955(.I(new_n20147_), .ZN(new_n20148_));
  OAI21_X1   g19956(.A1(new_n20143_), .A2(new_n1436_), .B(new_n20148_), .ZN(new_n20149_));
  NAND2_X1   g19957(.A1(new_n20149_), .A2(new_n20142_), .ZN(new_n20150_));
  OAI22_X1   g19958(.A1(new_n20143_), .A2(new_n1436_), .B1(new_n20141_), .B2(new_n20135_), .ZN(new_n20151_));
  NAND2_X1   g19959(.A1(new_n19499_), .A2(\asqrt[52] ), .ZN(new_n20152_));
  NOR4_X1    g19960(.A1(new_n19782_), .A2(\asqrt[52] ), .A3(new_n19494_), .A4(new_n19499_), .ZN(new_n20153_));
  XOR2_X1    g19961(.A1(new_n20153_), .A2(new_n20152_), .Z(new_n20154_));
  NAND2_X1   g19962(.A1(new_n20154_), .A2(new_n1096_), .ZN(new_n20155_));
  AOI21_X1   g19963(.A1(new_n20151_), .A2(\asqrt[52] ), .B(new_n20155_), .ZN(new_n20156_));
  NOR2_X1    g19964(.A1(new_n20156_), .A2(new_n20150_), .ZN(new_n20157_));
  AOI22_X1   g19965(.A1(new_n20151_), .A2(\asqrt[52] ), .B1(new_n20149_), .B2(new_n20142_), .ZN(new_n20158_));
  NOR4_X1    g19966(.A1(new_n19782_), .A2(\asqrt[53] ), .A3(new_n19502_), .A4(new_n19703_), .ZN(new_n20159_));
  AOI21_X1   g19967(.A1(new_n20152_), .A2(new_n19498_), .B(new_n1096_), .ZN(new_n20160_));
  NOR2_X1    g19968(.A1(new_n20159_), .A2(new_n20160_), .ZN(new_n20161_));
  NAND2_X1   g19969(.A1(new_n20161_), .A2(new_n970_), .ZN(new_n20162_));
  INV_X1     g19970(.I(new_n20162_), .ZN(new_n20163_));
  OAI21_X1   g19971(.A1(new_n20158_), .A2(new_n1096_), .B(new_n20163_), .ZN(new_n20164_));
  NAND2_X1   g19972(.A1(new_n20164_), .A2(new_n20157_), .ZN(new_n20165_));
  OAI22_X1   g19973(.A1(new_n20158_), .A2(new_n1096_), .B1(new_n20156_), .B2(new_n20150_), .ZN(new_n20166_));
  NOR4_X1    g19974(.A1(new_n19782_), .A2(\asqrt[54] ), .A3(new_n19509_), .A4(new_n19514_), .ZN(new_n20167_));
  XOR2_X1    g19975(.A1(new_n20167_), .A2(new_n19729_), .Z(new_n20168_));
  NAND2_X1   g19976(.A1(new_n20168_), .A2(new_n825_), .ZN(new_n20169_));
  AOI21_X1   g19977(.A1(new_n20166_), .A2(\asqrt[54] ), .B(new_n20169_), .ZN(new_n20170_));
  NOR2_X1    g19978(.A1(new_n20170_), .A2(new_n20165_), .ZN(new_n20171_));
  AOI22_X1   g19979(.A1(new_n20166_), .A2(\asqrt[54] ), .B1(new_n20164_), .B2(new_n20157_), .ZN(new_n20172_));
  NOR4_X1    g19980(.A1(new_n19782_), .A2(\asqrt[55] ), .A3(new_n19516_), .A4(new_n19710_), .ZN(new_n20173_));
  XOR2_X1    g19981(.A1(new_n20173_), .A2(new_n19717_), .Z(new_n20174_));
  NAND2_X1   g19982(.A1(new_n20174_), .A2(new_n724_), .ZN(new_n20175_));
  INV_X1     g19983(.I(new_n20175_), .ZN(new_n20176_));
  OAI21_X1   g19984(.A1(new_n20172_), .A2(new_n825_), .B(new_n20176_), .ZN(new_n20177_));
  NAND2_X1   g19985(.A1(new_n20177_), .A2(new_n20171_), .ZN(new_n20178_));
  OAI22_X1   g19986(.A1(new_n20172_), .A2(new_n825_), .B1(new_n20170_), .B2(new_n20165_), .ZN(new_n20179_));
  NOR4_X1    g19987(.A1(new_n19782_), .A2(\asqrt[56] ), .A3(new_n19522_), .A4(new_n19527_), .ZN(new_n20180_));
  XOR2_X1    g19988(.A1(new_n20180_), .A2(new_n19731_), .Z(new_n20181_));
  NAND2_X1   g19989(.A1(new_n20181_), .A2(new_n587_), .ZN(new_n20182_));
  AOI21_X1   g19990(.A1(new_n20179_), .A2(\asqrt[56] ), .B(new_n20182_), .ZN(new_n20183_));
  NOR2_X1    g19991(.A1(new_n20183_), .A2(new_n20178_), .ZN(new_n20184_));
  AOI22_X1   g19992(.A1(new_n20179_), .A2(\asqrt[56] ), .B1(new_n20177_), .B2(new_n20171_), .ZN(new_n20185_));
  NOR4_X1    g19993(.A1(new_n19782_), .A2(\asqrt[57] ), .A3(new_n19529_), .A4(new_n19721_), .ZN(new_n20186_));
  XOR2_X1    g19994(.A1(new_n20186_), .A2(new_n19719_), .Z(new_n20187_));
  NAND2_X1   g19995(.A1(new_n20187_), .A2(new_n504_), .ZN(new_n20188_));
  INV_X1     g19996(.I(new_n20188_), .ZN(new_n20189_));
  OAI21_X1   g19997(.A1(new_n20185_), .A2(new_n587_), .B(new_n20189_), .ZN(new_n20190_));
  NAND2_X1   g19998(.A1(new_n20190_), .A2(new_n20184_), .ZN(new_n20191_));
  OAI22_X1   g19999(.A1(new_n20185_), .A2(new_n587_), .B1(new_n20183_), .B2(new_n20178_), .ZN(new_n20192_));
  NOR4_X1    g20000(.A1(new_n19782_), .A2(\asqrt[58] ), .A3(new_n19535_), .A4(new_n19540_), .ZN(new_n20193_));
  XOR2_X1    g20001(.A1(new_n20193_), .A2(new_n19733_), .Z(new_n20194_));
  NAND2_X1   g20002(.A1(new_n20194_), .A2(new_n376_), .ZN(new_n20195_));
  AOI21_X1   g20003(.A1(new_n20192_), .A2(\asqrt[58] ), .B(new_n20195_), .ZN(new_n20196_));
  NOR2_X1    g20004(.A1(new_n20196_), .A2(new_n20191_), .ZN(new_n20197_));
  NAND2_X1   g20005(.A1(new_n20192_), .A2(\asqrt[58] ), .ZN(new_n20198_));
  AOI21_X1   g20006(.A1(new_n20198_), .A2(new_n20191_), .B(new_n376_), .ZN(new_n20199_));
  NOR4_X1    g20007(.A1(new_n19782_), .A2(\asqrt[59] ), .A3(new_n19542_), .A4(new_n19737_), .ZN(new_n20200_));
  XOR2_X1    g20008(.A1(new_n20200_), .A2(new_n19727_), .Z(new_n20201_));
  NAND2_X1   g20009(.A1(new_n20201_), .A2(new_n275_), .ZN(new_n20202_));
  OAI21_X1   g20010(.A1(new_n20199_), .A2(new_n20202_), .B(new_n20197_), .ZN(new_n20203_));
  OAI21_X1   g20011(.A1(new_n20197_), .A2(new_n20199_), .B(\asqrt[60] ), .ZN(new_n20204_));
  AOI21_X1   g20012(.A1(new_n20203_), .A2(new_n20204_), .B(new_n229_), .ZN(new_n20205_));
  AOI22_X1   g20013(.A1(new_n20192_), .A2(\asqrt[58] ), .B1(new_n20190_), .B2(new_n20184_), .ZN(new_n20206_));
  OAI22_X1   g20014(.A1(new_n20206_), .A2(new_n376_), .B1(new_n20196_), .B2(new_n20191_), .ZN(new_n20207_));
  NOR4_X1    g20015(.A1(new_n19782_), .A2(\asqrt[60] ), .A3(new_n19548_), .A4(new_n19552_), .ZN(new_n20208_));
  XOR2_X1    g20016(.A1(new_n20208_), .A2(new_n19735_), .Z(new_n20209_));
  NAND2_X1   g20017(.A1(new_n20209_), .A2(new_n229_), .ZN(new_n20210_));
  AOI21_X1   g20018(.A1(new_n20207_), .A2(\asqrt[60] ), .B(new_n20210_), .ZN(new_n20211_));
  INV_X1     g20019(.I(new_n19788_), .ZN(new_n20212_));
  NOR2_X1    g20020(.A1(new_n20212_), .A2(\asqrt[62] ), .ZN(new_n20213_));
  NOR3_X1    g20021(.A1(new_n20211_), .A2(new_n20203_), .A3(new_n20213_), .ZN(new_n20214_));
  AOI21_X1   g20022(.A1(new_n20214_), .A2(new_n20205_), .B(new_n19789_), .ZN(new_n20215_));
  NAND2_X1   g20023(.A1(new_n19780_), .A2(new_n19115_), .ZN(new_n20216_));
  AOI21_X1   g20024(.A1(new_n20216_), .A2(new_n19766_), .B(\asqrt[63] ), .ZN(new_n20217_));
  AOI21_X1   g20025(.A1(new_n20215_), .A2(new_n20217_), .B(new_n19784_), .ZN(new_n20218_));
  INV_X1     g20026(.I(new_n19784_), .ZN(new_n20219_));
  OAI21_X1   g20027(.A1(new_n19802_), .A2(new_n19799_), .B(new_n19795_), .ZN(new_n20220_));
  NAND3_X1   g20028(.A1(new_n19797_), .A2(\a[14] ), .A3(new_n19796_), .ZN(new_n20221_));
  NAND2_X1   g20029(.A1(new_n20220_), .A2(new_n20221_), .ZN(new_n20222_));
  INV_X1     g20030(.I(new_n19808_), .ZN(new_n20223_));
  NAND3_X1   g20031(.A1(new_n19818_), .A2(new_n19117_), .A3(new_n19782_), .ZN(new_n20224_));
  OAI21_X1   g20032(.A1(new_n19811_), .A2(new_n19118_), .B(\asqrt[7] ), .ZN(new_n20225_));
  NAND4_X1   g20033(.A1(new_n20224_), .A2(new_n20225_), .A3(new_n18495_), .A4(new_n20223_), .ZN(new_n20226_));
  NAND2_X1   g20034(.A1(new_n20226_), .A2(new_n20222_), .ZN(new_n20227_));
  NAND3_X1   g20035(.A1(new_n20220_), .A2(new_n20221_), .A3(new_n20223_), .ZN(new_n20228_));
  NAND3_X1   g20036(.A1(\asqrt[7] ), .A2(new_n19137_), .A3(new_n19827_), .ZN(new_n20229_));
  OAI21_X1   g20037(.A1(new_n19782_), .A2(new_n19828_), .B(new_n19136_), .ZN(new_n20230_));
  NAND3_X1   g20038(.A1(new_n20230_), .A2(new_n20229_), .A3(new_n17893_), .ZN(new_n20231_));
  AOI21_X1   g20039(.A1(new_n20228_), .A2(\asqrt[9] ), .B(new_n20231_), .ZN(new_n20232_));
  NOR2_X1    g20040(.A1(new_n20227_), .A2(new_n20232_), .ZN(new_n20233_));
  AOI22_X1   g20041(.A1(new_n20226_), .A2(new_n20222_), .B1(\asqrt[9] ), .B2(new_n20228_), .ZN(new_n20234_));
  OAI21_X1   g20042(.A1(new_n20234_), .A2(new_n17893_), .B(new_n19842_), .ZN(new_n20235_));
  NAND2_X1   g20043(.A1(new_n20235_), .A2(new_n20233_), .ZN(new_n20236_));
  OAI22_X1   g20044(.A1(new_n20234_), .A2(new_n17893_), .B1(new_n20227_), .B2(new_n20232_), .ZN(new_n20237_));
  AOI21_X1   g20045(.A1(new_n20237_), .A2(\asqrt[11] ), .B(new_n19850_), .ZN(new_n20238_));
  NOR2_X1    g20046(.A1(new_n20238_), .A2(new_n20236_), .ZN(new_n20239_));
  AOI22_X1   g20047(.A1(new_n20237_), .A2(\asqrt[11] ), .B1(new_n20235_), .B2(new_n20233_), .ZN(new_n20240_));
  INV_X1     g20048(.I(new_n19858_), .ZN(new_n20241_));
  OAI21_X1   g20049(.A1(new_n20240_), .A2(new_n16619_), .B(new_n20241_), .ZN(new_n20242_));
  NAND2_X1   g20050(.A1(new_n20242_), .A2(new_n20239_), .ZN(new_n20243_));
  OAI22_X1   g20051(.A1(new_n20240_), .A2(new_n16619_), .B1(new_n20238_), .B2(new_n20236_), .ZN(new_n20244_));
  AOI21_X1   g20052(.A1(new_n20244_), .A2(\asqrt[13] ), .B(new_n19865_), .ZN(new_n20245_));
  NOR2_X1    g20053(.A1(new_n20245_), .A2(new_n20243_), .ZN(new_n20246_));
  AOI22_X1   g20054(.A1(new_n20244_), .A2(\asqrt[13] ), .B1(new_n20242_), .B2(new_n20239_), .ZN(new_n20247_));
  INV_X1     g20055(.I(new_n19872_), .ZN(new_n20248_));
  OAI21_X1   g20056(.A1(new_n20247_), .A2(new_n15447_), .B(new_n20248_), .ZN(new_n20249_));
  NAND2_X1   g20057(.A1(new_n20249_), .A2(new_n20246_), .ZN(new_n20250_));
  OAI22_X1   g20058(.A1(new_n20247_), .A2(new_n15447_), .B1(new_n20245_), .B2(new_n20243_), .ZN(new_n20251_));
  AOI21_X1   g20059(.A1(new_n20251_), .A2(\asqrt[15] ), .B(new_n19878_), .ZN(new_n20252_));
  NOR2_X1    g20060(.A1(new_n20252_), .A2(new_n20250_), .ZN(new_n20253_));
  AOI22_X1   g20061(.A1(new_n20251_), .A2(\asqrt[15] ), .B1(new_n20249_), .B2(new_n20246_), .ZN(new_n20254_));
  INV_X1     g20062(.I(new_n19885_), .ZN(new_n20255_));
  OAI21_X1   g20063(.A1(new_n20254_), .A2(new_n14273_), .B(new_n20255_), .ZN(new_n20256_));
  NAND2_X1   g20064(.A1(new_n20256_), .A2(new_n20253_), .ZN(new_n20257_));
  OAI22_X1   g20065(.A1(new_n20254_), .A2(new_n14273_), .B1(new_n20252_), .B2(new_n20250_), .ZN(new_n20258_));
  AOI21_X1   g20066(.A1(new_n20258_), .A2(\asqrt[17] ), .B(new_n19892_), .ZN(new_n20259_));
  NOR2_X1    g20067(.A1(new_n20259_), .A2(new_n20257_), .ZN(new_n20260_));
  AOI22_X1   g20068(.A1(new_n20258_), .A2(\asqrt[17] ), .B1(new_n20256_), .B2(new_n20253_), .ZN(new_n20261_));
  INV_X1     g20069(.I(new_n19900_), .ZN(new_n20262_));
  OAI21_X1   g20070(.A1(new_n20261_), .A2(new_n13192_), .B(new_n20262_), .ZN(new_n20263_));
  NAND2_X1   g20071(.A1(new_n20263_), .A2(new_n20260_), .ZN(new_n20264_));
  OAI22_X1   g20072(.A1(new_n20261_), .A2(new_n13192_), .B1(new_n20259_), .B2(new_n20257_), .ZN(new_n20265_));
  AOI21_X1   g20073(.A1(new_n20265_), .A2(\asqrt[19] ), .B(new_n19907_), .ZN(new_n20266_));
  NOR2_X1    g20074(.A1(new_n20266_), .A2(new_n20264_), .ZN(new_n20267_));
  AOI22_X1   g20075(.A1(new_n20265_), .A2(\asqrt[19] ), .B1(new_n20263_), .B2(new_n20260_), .ZN(new_n20268_));
  INV_X1     g20076(.I(new_n19915_), .ZN(new_n20269_));
  OAI21_X1   g20077(.A1(new_n20268_), .A2(new_n12101_), .B(new_n20269_), .ZN(new_n20270_));
  NAND2_X1   g20078(.A1(new_n20270_), .A2(new_n20267_), .ZN(new_n20271_));
  OAI22_X1   g20079(.A1(new_n20268_), .A2(new_n12101_), .B1(new_n20266_), .B2(new_n20264_), .ZN(new_n20272_));
  AOI21_X1   g20080(.A1(new_n20272_), .A2(\asqrt[21] ), .B(new_n19922_), .ZN(new_n20273_));
  NOR2_X1    g20081(.A1(new_n20273_), .A2(new_n20271_), .ZN(new_n20274_));
  AOI22_X1   g20082(.A1(new_n20272_), .A2(\asqrt[21] ), .B1(new_n20270_), .B2(new_n20267_), .ZN(new_n20275_));
  INV_X1     g20083(.I(new_n19930_), .ZN(new_n20276_));
  OAI21_X1   g20084(.A1(new_n20275_), .A2(new_n11105_), .B(new_n20276_), .ZN(new_n20277_));
  NAND2_X1   g20085(.A1(new_n20277_), .A2(new_n20274_), .ZN(new_n20278_));
  OAI22_X1   g20086(.A1(new_n20275_), .A2(new_n11105_), .B1(new_n20273_), .B2(new_n20271_), .ZN(new_n20279_));
  AOI21_X1   g20087(.A1(new_n20279_), .A2(\asqrt[23] ), .B(new_n19937_), .ZN(new_n20280_));
  NOR2_X1    g20088(.A1(new_n20280_), .A2(new_n20278_), .ZN(new_n20281_));
  AOI22_X1   g20089(.A1(new_n20279_), .A2(\asqrt[23] ), .B1(new_n20277_), .B2(new_n20274_), .ZN(new_n20282_));
  INV_X1     g20090(.I(new_n19945_), .ZN(new_n20283_));
  OAI21_X1   g20091(.A1(new_n20282_), .A2(new_n10104_), .B(new_n20283_), .ZN(new_n20284_));
  NAND2_X1   g20092(.A1(new_n20284_), .A2(new_n20281_), .ZN(new_n20285_));
  OAI22_X1   g20093(.A1(new_n20282_), .A2(new_n10104_), .B1(new_n20280_), .B2(new_n20278_), .ZN(new_n20286_));
  AOI21_X1   g20094(.A1(new_n20286_), .A2(\asqrt[25] ), .B(new_n19952_), .ZN(new_n20287_));
  NOR2_X1    g20095(.A1(new_n20287_), .A2(new_n20285_), .ZN(new_n20288_));
  AOI22_X1   g20096(.A1(new_n20286_), .A2(\asqrt[25] ), .B1(new_n20284_), .B2(new_n20281_), .ZN(new_n20289_));
  INV_X1     g20097(.I(new_n19960_), .ZN(new_n20290_));
  OAI21_X1   g20098(.A1(new_n20289_), .A2(new_n9212_), .B(new_n20290_), .ZN(new_n20291_));
  NAND2_X1   g20099(.A1(new_n20291_), .A2(new_n20288_), .ZN(new_n20292_));
  OAI22_X1   g20100(.A1(new_n20289_), .A2(new_n9212_), .B1(new_n20287_), .B2(new_n20285_), .ZN(new_n20293_));
  AOI21_X1   g20101(.A1(new_n20293_), .A2(\asqrt[27] ), .B(new_n19967_), .ZN(new_n20294_));
  NOR2_X1    g20102(.A1(new_n20294_), .A2(new_n20292_), .ZN(new_n20295_));
  AOI22_X1   g20103(.A1(new_n20293_), .A2(\asqrt[27] ), .B1(new_n20291_), .B2(new_n20288_), .ZN(new_n20296_));
  INV_X1     g20104(.I(new_n19975_), .ZN(new_n20297_));
  OAI21_X1   g20105(.A1(new_n20296_), .A2(new_n8319_), .B(new_n20297_), .ZN(new_n20298_));
  NAND2_X1   g20106(.A1(new_n20298_), .A2(new_n20295_), .ZN(new_n20299_));
  OAI22_X1   g20107(.A1(new_n20296_), .A2(new_n8319_), .B1(new_n20294_), .B2(new_n20292_), .ZN(new_n20300_));
  AOI21_X1   g20108(.A1(new_n20300_), .A2(\asqrt[29] ), .B(new_n19982_), .ZN(new_n20301_));
  NOR2_X1    g20109(.A1(new_n20301_), .A2(new_n20299_), .ZN(new_n20302_));
  AOI22_X1   g20110(.A1(new_n20300_), .A2(\asqrt[29] ), .B1(new_n20298_), .B2(new_n20295_), .ZN(new_n20303_));
  INV_X1     g20111(.I(new_n19990_), .ZN(new_n20304_));
  OAI21_X1   g20112(.A1(new_n20303_), .A2(new_n7517_), .B(new_n20304_), .ZN(new_n20305_));
  NAND2_X1   g20113(.A1(new_n20305_), .A2(new_n20302_), .ZN(new_n20306_));
  OAI22_X1   g20114(.A1(new_n20303_), .A2(new_n7517_), .B1(new_n20301_), .B2(new_n20299_), .ZN(new_n20307_));
  AOI21_X1   g20115(.A1(new_n20307_), .A2(\asqrt[31] ), .B(new_n19997_), .ZN(new_n20308_));
  NOR2_X1    g20116(.A1(new_n20308_), .A2(new_n20306_), .ZN(new_n20309_));
  AOI22_X1   g20117(.A1(new_n20307_), .A2(\asqrt[31] ), .B1(new_n20305_), .B2(new_n20302_), .ZN(new_n20310_));
  INV_X1     g20118(.I(new_n20005_), .ZN(new_n20311_));
  OAI21_X1   g20119(.A1(new_n20310_), .A2(new_n6708_), .B(new_n20311_), .ZN(new_n20312_));
  NAND2_X1   g20120(.A1(new_n20312_), .A2(new_n20309_), .ZN(new_n20313_));
  OAI22_X1   g20121(.A1(new_n20310_), .A2(new_n6708_), .B1(new_n20308_), .B2(new_n20306_), .ZN(new_n20314_));
  AOI21_X1   g20122(.A1(new_n20314_), .A2(\asqrt[33] ), .B(new_n20012_), .ZN(new_n20315_));
  NOR2_X1    g20123(.A1(new_n20315_), .A2(new_n20313_), .ZN(new_n20316_));
  AOI22_X1   g20124(.A1(new_n20314_), .A2(\asqrt[33] ), .B1(new_n20312_), .B2(new_n20309_), .ZN(new_n20317_));
  INV_X1     g20125(.I(new_n20020_), .ZN(new_n20318_));
  OAI21_X1   g20126(.A1(new_n20317_), .A2(new_n5991_), .B(new_n20318_), .ZN(new_n20319_));
  NAND2_X1   g20127(.A1(new_n20319_), .A2(new_n20316_), .ZN(new_n20320_));
  OAI22_X1   g20128(.A1(new_n20317_), .A2(new_n5991_), .B1(new_n20315_), .B2(new_n20313_), .ZN(new_n20321_));
  AOI21_X1   g20129(.A1(new_n20321_), .A2(\asqrt[35] ), .B(new_n20027_), .ZN(new_n20322_));
  NOR2_X1    g20130(.A1(new_n20322_), .A2(new_n20320_), .ZN(new_n20323_));
  AOI22_X1   g20131(.A1(new_n20321_), .A2(\asqrt[35] ), .B1(new_n20319_), .B2(new_n20316_), .ZN(new_n20324_));
  INV_X1     g20132(.I(new_n20035_), .ZN(new_n20325_));
  OAI21_X1   g20133(.A1(new_n20324_), .A2(new_n5273_), .B(new_n20325_), .ZN(new_n20326_));
  NAND2_X1   g20134(.A1(new_n20326_), .A2(new_n20323_), .ZN(new_n20327_));
  OAI22_X1   g20135(.A1(new_n20324_), .A2(new_n5273_), .B1(new_n20322_), .B2(new_n20320_), .ZN(new_n20328_));
  AOI21_X1   g20136(.A1(new_n20328_), .A2(\asqrt[37] ), .B(new_n20042_), .ZN(new_n20329_));
  NOR2_X1    g20137(.A1(new_n20329_), .A2(new_n20327_), .ZN(new_n20330_));
  AOI22_X1   g20138(.A1(new_n20328_), .A2(\asqrt[37] ), .B1(new_n20326_), .B2(new_n20323_), .ZN(new_n20331_));
  INV_X1     g20139(.I(new_n20050_), .ZN(new_n20332_));
  OAI21_X1   g20140(.A1(new_n20331_), .A2(new_n4645_), .B(new_n20332_), .ZN(new_n20333_));
  NAND2_X1   g20141(.A1(new_n20333_), .A2(new_n20330_), .ZN(new_n20334_));
  OAI22_X1   g20142(.A1(new_n20331_), .A2(new_n4645_), .B1(new_n20329_), .B2(new_n20327_), .ZN(new_n20335_));
  AOI21_X1   g20143(.A1(new_n20335_), .A2(\asqrt[39] ), .B(new_n20057_), .ZN(new_n20336_));
  NOR2_X1    g20144(.A1(new_n20336_), .A2(new_n20334_), .ZN(new_n20337_));
  AOI22_X1   g20145(.A1(new_n20335_), .A2(\asqrt[39] ), .B1(new_n20333_), .B2(new_n20330_), .ZN(new_n20338_));
  INV_X1     g20146(.I(new_n20065_), .ZN(new_n20339_));
  OAI21_X1   g20147(.A1(new_n20338_), .A2(new_n4018_), .B(new_n20339_), .ZN(new_n20340_));
  NAND2_X1   g20148(.A1(new_n20340_), .A2(new_n20337_), .ZN(new_n20341_));
  OAI22_X1   g20149(.A1(new_n20338_), .A2(new_n4018_), .B1(new_n20336_), .B2(new_n20334_), .ZN(new_n20342_));
  AOI21_X1   g20150(.A1(new_n20342_), .A2(\asqrt[41] ), .B(new_n20072_), .ZN(new_n20343_));
  NOR2_X1    g20151(.A1(new_n20343_), .A2(new_n20341_), .ZN(new_n20344_));
  AOI22_X1   g20152(.A1(new_n20342_), .A2(\asqrt[41] ), .B1(new_n20340_), .B2(new_n20337_), .ZN(new_n20345_));
  INV_X1     g20153(.I(new_n20080_), .ZN(new_n20346_));
  OAI21_X1   g20154(.A1(new_n20345_), .A2(new_n3481_), .B(new_n20346_), .ZN(new_n20347_));
  NAND2_X1   g20155(.A1(new_n20347_), .A2(new_n20344_), .ZN(new_n20348_));
  OAI22_X1   g20156(.A1(new_n20345_), .A2(new_n3481_), .B1(new_n20343_), .B2(new_n20341_), .ZN(new_n20349_));
  AOI21_X1   g20157(.A1(new_n20349_), .A2(\asqrt[43] ), .B(new_n20087_), .ZN(new_n20350_));
  NOR2_X1    g20158(.A1(new_n20350_), .A2(new_n20348_), .ZN(new_n20351_));
  AOI22_X1   g20159(.A1(new_n20349_), .A2(\asqrt[43] ), .B1(new_n20347_), .B2(new_n20344_), .ZN(new_n20352_));
  INV_X1     g20160(.I(new_n20095_), .ZN(new_n20353_));
  OAI21_X1   g20161(.A1(new_n20352_), .A2(new_n2941_), .B(new_n20353_), .ZN(new_n20354_));
  NAND2_X1   g20162(.A1(new_n20354_), .A2(new_n20351_), .ZN(new_n20355_));
  OAI22_X1   g20163(.A1(new_n20352_), .A2(new_n2941_), .B1(new_n20350_), .B2(new_n20348_), .ZN(new_n20356_));
  AOI21_X1   g20164(.A1(new_n20356_), .A2(\asqrt[45] ), .B(new_n20102_), .ZN(new_n20357_));
  NOR2_X1    g20165(.A1(new_n20357_), .A2(new_n20355_), .ZN(new_n20358_));
  AOI22_X1   g20166(.A1(new_n20356_), .A2(\asqrt[45] ), .B1(new_n20354_), .B2(new_n20351_), .ZN(new_n20359_));
  INV_X1     g20167(.I(new_n20110_), .ZN(new_n20360_));
  OAI21_X1   g20168(.A1(new_n20359_), .A2(new_n2488_), .B(new_n20360_), .ZN(new_n20361_));
  NAND2_X1   g20169(.A1(new_n20361_), .A2(new_n20358_), .ZN(new_n20362_));
  OAI22_X1   g20170(.A1(new_n20359_), .A2(new_n2488_), .B1(new_n20357_), .B2(new_n20355_), .ZN(new_n20363_));
  AOI21_X1   g20171(.A1(new_n20363_), .A2(\asqrt[47] ), .B(new_n20117_), .ZN(new_n20364_));
  NOR2_X1    g20172(.A1(new_n20364_), .A2(new_n20362_), .ZN(new_n20365_));
  AOI22_X1   g20173(.A1(new_n20363_), .A2(\asqrt[47] ), .B1(new_n20361_), .B2(new_n20358_), .ZN(new_n20366_));
  INV_X1     g20174(.I(new_n20125_), .ZN(new_n20367_));
  OAI21_X1   g20175(.A1(new_n20366_), .A2(new_n2046_), .B(new_n20367_), .ZN(new_n20368_));
  NAND2_X1   g20176(.A1(new_n20368_), .A2(new_n20365_), .ZN(new_n20369_));
  OAI22_X1   g20177(.A1(new_n20366_), .A2(new_n2046_), .B1(new_n20364_), .B2(new_n20362_), .ZN(new_n20370_));
  AOI21_X1   g20178(.A1(new_n20370_), .A2(\asqrt[49] ), .B(new_n20132_), .ZN(new_n20371_));
  NOR2_X1    g20179(.A1(new_n20371_), .A2(new_n20369_), .ZN(new_n20372_));
  AOI22_X1   g20180(.A1(new_n20370_), .A2(\asqrt[49] ), .B1(new_n20368_), .B2(new_n20365_), .ZN(new_n20373_));
  INV_X1     g20181(.I(new_n20140_), .ZN(new_n20374_));
  OAI21_X1   g20182(.A1(new_n20373_), .A2(new_n1595_), .B(new_n20374_), .ZN(new_n20375_));
  NAND2_X1   g20183(.A1(new_n20375_), .A2(new_n20372_), .ZN(new_n20376_));
  OAI22_X1   g20184(.A1(new_n20373_), .A2(new_n1595_), .B1(new_n20371_), .B2(new_n20369_), .ZN(new_n20377_));
  AOI21_X1   g20185(.A1(new_n20377_), .A2(\asqrt[51] ), .B(new_n20147_), .ZN(new_n20378_));
  NOR2_X1    g20186(.A1(new_n20378_), .A2(new_n20376_), .ZN(new_n20379_));
  AOI22_X1   g20187(.A1(new_n20377_), .A2(\asqrt[51] ), .B1(new_n20375_), .B2(new_n20372_), .ZN(new_n20380_));
  INV_X1     g20188(.I(new_n20155_), .ZN(new_n20381_));
  OAI21_X1   g20189(.A1(new_n20380_), .A2(new_n1260_), .B(new_n20381_), .ZN(new_n20382_));
  NAND2_X1   g20190(.A1(new_n20382_), .A2(new_n20379_), .ZN(new_n20383_));
  OAI22_X1   g20191(.A1(new_n20380_), .A2(new_n1260_), .B1(new_n20378_), .B2(new_n20376_), .ZN(new_n20384_));
  AOI21_X1   g20192(.A1(new_n20384_), .A2(\asqrt[53] ), .B(new_n20162_), .ZN(new_n20385_));
  NOR2_X1    g20193(.A1(new_n20385_), .A2(new_n20383_), .ZN(new_n20386_));
  AOI22_X1   g20194(.A1(new_n20384_), .A2(\asqrt[53] ), .B1(new_n20382_), .B2(new_n20379_), .ZN(new_n20387_));
  INV_X1     g20195(.I(new_n20169_), .ZN(new_n20388_));
  OAI21_X1   g20196(.A1(new_n20387_), .A2(new_n970_), .B(new_n20388_), .ZN(new_n20389_));
  NAND2_X1   g20197(.A1(new_n20389_), .A2(new_n20386_), .ZN(new_n20390_));
  OAI22_X1   g20198(.A1(new_n20387_), .A2(new_n970_), .B1(new_n20385_), .B2(new_n20383_), .ZN(new_n20391_));
  AOI21_X1   g20199(.A1(new_n20391_), .A2(\asqrt[55] ), .B(new_n20175_), .ZN(new_n20392_));
  NOR2_X1    g20200(.A1(new_n20392_), .A2(new_n20390_), .ZN(new_n20393_));
  AOI22_X1   g20201(.A1(new_n20391_), .A2(\asqrt[55] ), .B1(new_n20389_), .B2(new_n20386_), .ZN(new_n20394_));
  INV_X1     g20202(.I(new_n20182_), .ZN(new_n20395_));
  OAI21_X1   g20203(.A1(new_n20394_), .A2(new_n724_), .B(new_n20395_), .ZN(new_n20396_));
  NAND2_X1   g20204(.A1(new_n20396_), .A2(new_n20393_), .ZN(new_n20397_));
  OAI22_X1   g20205(.A1(new_n20394_), .A2(new_n724_), .B1(new_n20392_), .B2(new_n20390_), .ZN(new_n20398_));
  AOI21_X1   g20206(.A1(new_n20398_), .A2(\asqrt[57] ), .B(new_n20188_), .ZN(new_n20399_));
  NOR2_X1    g20207(.A1(new_n20399_), .A2(new_n20397_), .ZN(new_n20400_));
  AOI22_X1   g20208(.A1(new_n20398_), .A2(\asqrt[57] ), .B1(new_n20396_), .B2(new_n20393_), .ZN(new_n20401_));
  INV_X1     g20209(.I(new_n20195_), .ZN(new_n20402_));
  OAI21_X1   g20210(.A1(new_n20401_), .A2(new_n504_), .B(new_n20402_), .ZN(new_n20403_));
  NAND2_X1   g20211(.A1(new_n20403_), .A2(new_n20400_), .ZN(new_n20404_));
  OAI22_X1   g20212(.A1(new_n20401_), .A2(new_n504_), .B1(new_n20399_), .B2(new_n20397_), .ZN(new_n20405_));
  AOI21_X1   g20213(.A1(new_n20405_), .A2(\asqrt[59] ), .B(new_n20202_), .ZN(new_n20406_));
  NOR2_X1    g20214(.A1(new_n20406_), .A2(new_n20404_), .ZN(new_n20407_));
  AOI22_X1   g20215(.A1(new_n20405_), .A2(\asqrt[59] ), .B1(new_n20403_), .B2(new_n20400_), .ZN(new_n20408_));
  OAI22_X1   g20216(.A1(new_n20408_), .A2(new_n275_), .B1(new_n20406_), .B2(new_n20404_), .ZN(new_n20409_));
  INV_X1     g20217(.I(new_n20210_), .ZN(new_n20410_));
  OAI21_X1   g20218(.A1(new_n20408_), .A2(new_n275_), .B(new_n20410_), .ZN(new_n20411_));
  AOI22_X1   g20219(.A1(new_n20409_), .A2(\asqrt[61] ), .B1(new_n20411_), .B2(new_n20407_), .ZN(new_n20412_));
  NAND4_X1   g20220(.A1(new_n20412_), .A2(new_n196_), .A3(new_n20219_), .A4(new_n20212_), .ZN(new_n20413_));
  NAND2_X1   g20221(.A1(new_n19778_), .A2(new_n19115_), .ZN(new_n20414_));
  XOR2_X1    g20222(.A1(new_n19778_), .A2(\asqrt[63] ), .Z(new_n20415_));
  AOI21_X1   g20223(.A1(\asqrt[7] ), .A2(new_n20414_), .B(new_n20415_), .ZN(new_n20416_));
  INV_X1     g20224(.I(new_n20416_), .ZN(new_n20417_));
  NOR2_X1    g20225(.A1(new_n20413_), .A2(new_n20417_), .ZN(new_n20418_));
  NAND4_X1   g20226(.A1(new_n20418_), .A2(\a[13] ), .A3(new_n20218_), .A4(new_n19772_), .ZN(new_n20419_));
  INV_X1     g20227(.I(\a[13] ), .ZN(new_n20420_));
  NOR2_X1    g20228(.A1(new_n20420_), .A2(\a[12] ), .ZN(new_n20421_));
  INV_X1     g20229(.I(new_n20421_), .ZN(new_n20422_));
  AOI21_X1   g20230(.A1(new_n20419_), .A2(new_n20422_), .B(new_n19763_), .ZN(new_n20423_));
  INV_X1     g20231(.I(new_n19789_), .ZN(new_n20424_));
  NAND2_X1   g20232(.A1(new_n20405_), .A2(\asqrt[59] ), .ZN(new_n20425_));
  AOI21_X1   g20233(.A1(new_n20425_), .A2(new_n20404_), .B(new_n275_), .ZN(new_n20426_));
  OAI21_X1   g20234(.A1(new_n20407_), .A2(new_n20426_), .B(\asqrt[61] ), .ZN(new_n20427_));
  INV_X1     g20235(.I(new_n20213_), .ZN(new_n20428_));
  NAND3_X1   g20236(.A1(new_n20411_), .A2(new_n20407_), .A3(new_n20428_), .ZN(new_n20429_));
  OAI21_X1   g20237(.A1(new_n20429_), .A2(new_n20427_), .B(new_n20424_), .ZN(new_n20430_));
  INV_X1     g20238(.I(new_n20217_), .ZN(new_n20431_));
  OAI21_X1   g20239(.A1(new_n20430_), .A2(new_n20431_), .B(new_n20219_), .ZN(new_n20432_));
  OAI21_X1   g20240(.A1(new_n20412_), .A2(new_n196_), .B(new_n19784_), .ZN(new_n20433_));
  NOR2_X1    g20241(.A1(new_n20211_), .A2(new_n20203_), .ZN(new_n20434_));
  NOR4_X1    g20242(.A1(new_n20434_), .A2(new_n20205_), .A3(\asqrt[62] ), .A4(new_n19788_), .ZN(new_n20435_));
  NAND3_X1   g20243(.A1(new_n20433_), .A2(new_n20435_), .A3(new_n20416_), .ZN(new_n20436_));
  NOR4_X1    g20244(.A1(new_n20436_), .A2(new_n20420_), .A3(new_n19771_), .A4(new_n20432_), .ZN(new_n20437_));
  NOR3_X1    g20245(.A1(new_n20437_), .A2(new_n19750_), .A3(new_n19762_), .ZN(new_n20438_));
  NOR2_X1    g20246(.A1(new_n20438_), .A2(new_n20423_), .ZN(new_n20439_));
  NAND4_X1   g20247(.A1(new_n19781_), .A2(new_n19114_), .A3(new_n19748_), .A4(new_n19752_), .ZN(new_n20441_));
  NOR2_X1    g20248(.A1(new_n19782_), .A2(new_n19750_), .ZN(new_n20442_));
  XOR2_X1    g20249(.A1(new_n20442_), .A2(new_n20441_), .Z(new_n20443_));
  NOR2_X1    g20250(.A1(new_n20443_), .A2(new_n19759_), .ZN(new_n20444_));
  NOR4_X1    g20251(.A1(new_n20432_), .A2(new_n19771_), .A3(new_n20413_), .A4(new_n20417_), .ZN(\asqrt[6] ));
  NAND2_X1   g20252(.A1(new_n19771_), .A2(\asqrt[7] ), .ZN(new_n20446_));
  NOR2_X1    g20253(.A1(new_n20446_), .A2(new_n20416_), .ZN(new_n20447_));
  INV_X1     g20254(.I(new_n20447_), .ZN(new_n20448_));
  AOI21_X1   g20255(.A1(new_n20433_), .A2(new_n20435_), .B(new_n20448_), .ZN(new_n20449_));
  AOI21_X1   g20256(.A1(new_n20449_), .A2(new_n20432_), .B(\a[14] ), .ZN(new_n20450_));
  NOR3_X1    g20257(.A1(new_n20450_), .A2(new_n19792_), .A3(\asqrt[6] ), .ZN(new_n20451_));
  NAND2_X1   g20258(.A1(new_n20411_), .A2(new_n20407_), .ZN(new_n20452_));
  NAND2_X1   g20259(.A1(new_n20452_), .A2(new_n20427_), .ZN(new_n20453_));
  NOR4_X1    g20260(.A1(new_n20453_), .A2(\asqrt[62] ), .A3(new_n19784_), .A4(new_n19788_), .ZN(new_n20454_));
  NAND4_X1   g20261(.A1(new_n20218_), .A2(new_n20454_), .A3(new_n19772_), .A4(new_n20416_), .ZN(new_n20455_));
  NAND2_X1   g20262(.A1(new_n20413_), .A2(new_n20447_), .ZN(new_n20456_));
  OAI21_X1   g20263(.A1(new_n20456_), .A2(new_n20218_), .B(new_n19790_), .ZN(new_n20457_));
  AOI21_X1   g20264(.A1(new_n20457_), .A2(new_n19791_), .B(new_n20455_), .ZN(new_n20458_));
  NOR4_X1    g20265(.A1(new_n20458_), .A2(new_n20451_), .A3(\asqrt[8] ), .A4(new_n20444_), .ZN(new_n20459_));
  NOR2_X1    g20266(.A1(new_n20459_), .A2(new_n20439_), .ZN(new_n20460_));
  NOR3_X1    g20267(.A1(new_n20438_), .A2(new_n20423_), .A3(new_n20444_), .ZN(new_n20461_));
  AOI21_X1   g20268(.A1(\asqrt[7] ), .A2(new_n19790_), .B(\a[15] ), .ZN(new_n20462_));
  NOR2_X1    g20269(.A1(new_n19797_), .A2(\a[14] ), .ZN(new_n20463_));
  AOI21_X1   g20270(.A1(\asqrt[7] ), .A2(\a[14] ), .B(new_n19794_), .ZN(new_n20464_));
  OAI21_X1   g20271(.A1(new_n20463_), .A2(new_n20462_), .B(new_n20464_), .ZN(new_n20465_));
  NOR3_X1    g20272(.A1(new_n20455_), .A2(new_n19808_), .A3(new_n20465_), .ZN(new_n20466_));
  INV_X1     g20273(.I(new_n20465_), .ZN(new_n20467_));
  AOI21_X1   g20274(.A1(\asqrt[6] ), .A2(new_n20467_), .B(new_n20223_), .ZN(new_n20468_));
  NOR3_X1    g20275(.A1(new_n20466_), .A2(new_n20468_), .A3(\asqrt[9] ), .ZN(new_n20469_));
  OAI21_X1   g20276(.A1(new_n20461_), .A2(new_n19100_), .B(new_n20469_), .ZN(new_n20470_));
  NAND2_X1   g20277(.A1(new_n20470_), .A2(new_n20460_), .ZN(new_n20471_));
  OAI22_X1   g20278(.A1(new_n20439_), .A2(new_n20459_), .B1(new_n20461_), .B2(new_n19100_), .ZN(new_n20472_));
  NOR2_X1    g20279(.A1(new_n19819_), .A2(new_n19812_), .ZN(new_n20473_));
  NOR4_X1    g20280(.A1(new_n20455_), .A2(\asqrt[9] ), .A3(new_n20473_), .A4(new_n20228_), .ZN(new_n20474_));
  AOI21_X1   g20281(.A1(new_n19804_), .A2(new_n20223_), .B(new_n18495_), .ZN(new_n20475_));
  NOR2_X1    g20282(.A1(new_n20474_), .A2(new_n20475_), .ZN(new_n20476_));
  NAND2_X1   g20283(.A1(new_n20476_), .A2(new_n17893_), .ZN(new_n20477_));
  AOI21_X1   g20284(.A1(new_n20472_), .A2(\asqrt[9] ), .B(new_n20477_), .ZN(new_n20478_));
  NOR2_X1    g20285(.A1(new_n20478_), .A2(new_n20471_), .ZN(new_n20479_));
  AOI22_X1   g20286(.A1(new_n20472_), .A2(\asqrt[9] ), .B1(new_n20460_), .B2(new_n20470_), .ZN(new_n20480_));
  NOR2_X1    g20287(.A1(new_n20234_), .A2(new_n17893_), .ZN(new_n20481_));
  NAND2_X1   g20288(.A1(new_n20230_), .A2(new_n20229_), .ZN(new_n20482_));
  NAND4_X1   g20289(.A1(\asqrt[6] ), .A2(new_n17893_), .A3(new_n20482_), .A4(new_n20234_), .ZN(new_n20483_));
  XOR2_X1    g20290(.A1(new_n20483_), .A2(new_n20481_), .Z(new_n20484_));
  NAND2_X1   g20291(.A1(new_n20484_), .A2(new_n17271_), .ZN(new_n20485_));
  INV_X1     g20292(.I(new_n20485_), .ZN(new_n20486_));
  OAI21_X1   g20293(.A1(new_n20480_), .A2(new_n17893_), .B(new_n20486_), .ZN(new_n20487_));
  NAND2_X1   g20294(.A1(new_n20487_), .A2(new_n20479_), .ZN(new_n20488_));
  OAI22_X1   g20295(.A1(new_n20480_), .A2(new_n17893_), .B1(new_n20478_), .B2(new_n20471_), .ZN(new_n20489_));
  NAND2_X1   g20296(.A1(new_n20237_), .A2(\asqrt[11] ), .ZN(new_n20490_));
  NOR2_X1    g20297(.A1(new_n19840_), .A2(new_n19841_), .ZN(new_n20491_));
  NOR4_X1    g20298(.A1(new_n20455_), .A2(\asqrt[11] ), .A3(new_n20491_), .A4(new_n20237_), .ZN(new_n20492_));
  XOR2_X1    g20299(.A1(new_n20492_), .A2(new_n20490_), .Z(new_n20493_));
  NAND2_X1   g20300(.A1(new_n20493_), .A2(new_n16619_), .ZN(new_n20494_));
  AOI21_X1   g20301(.A1(new_n20489_), .A2(\asqrt[11] ), .B(new_n20494_), .ZN(new_n20495_));
  NOR2_X1    g20302(.A1(new_n20495_), .A2(new_n20488_), .ZN(new_n20496_));
  AOI22_X1   g20303(.A1(new_n20489_), .A2(\asqrt[11] ), .B1(new_n20487_), .B2(new_n20479_), .ZN(new_n20497_));
  NOR4_X1    g20304(.A1(new_n20455_), .A2(\asqrt[12] ), .A3(new_n19849_), .A4(new_n19854_), .ZN(new_n20498_));
  AOI21_X1   g20305(.A1(new_n20490_), .A2(new_n20236_), .B(new_n16619_), .ZN(new_n20499_));
  NOR2_X1    g20306(.A1(new_n20498_), .A2(new_n20499_), .ZN(new_n20500_));
  NAND2_X1   g20307(.A1(new_n20500_), .A2(new_n16060_), .ZN(new_n20501_));
  INV_X1     g20308(.I(new_n20501_), .ZN(new_n20502_));
  OAI21_X1   g20309(.A1(new_n20497_), .A2(new_n16619_), .B(new_n20502_), .ZN(new_n20503_));
  NAND2_X1   g20310(.A1(new_n20503_), .A2(new_n20496_), .ZN(new_n20504_));
  OAI22_X1   g20311(.A1(new_n20497_), .A2(new_n16619_), .B1(new_n20495_), .B2(new_n20488_), .ZN(new_n20505_));
  NAND2_X1   g20312(.A1(new_n20244_), .A2(\asqrt[13] ), .ZN(new_n20506_));
  NOR4_X1    g20313(.A1(new_n20455_), .A2(\asqrt[13] ), .A3(new_n19857_), .A4(new_n20244_), .ZN(new_n20507_));
  XOR2_X1    g20314(.A1(new_n20507_), .A2(new_n20506_), .Z(new_n20508_));
  NAND2_X1   g20315(.A1(new_n20508_), .A2(new_n15447_), .ZN(new_n20509_));
  AOI21_X1   g20316(.A1(new_n20505_), .A2(\asqrt[13] ), .B(new_n20509_), .ZN(new_n20510_));
  NOR2_X1    g20317(.A1(new_n20510_), .A2(new_n20504_), .ZN(new_n20511_));
  AOI22_X1   g20318(.A1(new_n20505_), .A2(\asqrt[13] ), .B1(new_n20503_), .B2(new_n20496_), .ZN(new_n20512_));
  NOR4_X1    g20319(.A1(new_n20455_), .A2(\asqrt[14] ), .A3(new_n19864_), .A4(new_n19869_), .ZN(new_n20513_));
  AOI21_X1   g20320(.A1(new_n20506_), .A2(new_n20243_), .B(new_n15447_), .ZN(new_n20514_));
  NOR2_X1    g20321(.A1(new_n20513_), .A2(new_n20514_), .ZN(new_n20515_));
  NAND2_X1   g20322(.A1(new_n20515_), .A2(new_n14871_), .ZN(new_n20516_));
  INV_X1     g20323(.I(new_n20516_), .ZN(new_n20517_));
  OAI21_X1   g20324(.A1(new_n20512_), .A2(new_n15447_), .B(new_n20517_), .ZN(new_n20518_));
  NAND2_X1   g20325(.A1(new_n20518_), .A2(new_n20511_), .ZN(new_n20519_));
  OAI22_X1   g20326(.A1(new_n20512_), .A2(new_n15447_), .B1(new_n20510_), .B2(new_n20504_), .ZN(new_n20520_));
  NAND2_X1   g20327(.A1(new_n20251_), .A2(\asqrt[15] ), .ZN(new_n20521_));
  NOR4_X1    g20328(.A1(new_n20455_), .A2(\asqrt[15] ), .A3(new_n19871_), .A4(new_n20251_), .ZN(new_n20522_));
  XOR2_X1    g20329(.A1(new_n20522_), .A2(new_n20521_), .Z(new_n20523_));
  NAND2_X1   g20330(.A1(new_n20523_), .A2(new_n14273_), .ZN(new_n20524_));
  AOI21_X1   g20331(.A1(new_n20520_), .A2(\asqrt[15] ), .B(new_n20524_), .ZN(new_n20525_));
  NOR2_X1    g20332(.A1(new_n20525_), .A2(new_n20519_), .ZN(new_n20526_));
  AOI22_X1   g20333(.A1(new_n20520_), .A2(\asqrt[15] ), .B1(new_n20518_), .B2(new_n20511_), .ZN(new_n20527_));
  NOR4_X1    g20334(.A1(new_n20455_), .A2(\asqrt[16] ), .A3(new_n19877_), .A4(new_n19882_), .ZN(new_n20528_));
  AOI21_X1   g20335(.A1(new_n20521_), .A2(new_n20250_), .B(new_n14273_), .ZN(new_n20529_));
  NOR2_X1    g20336(.A1(new_n20528_), .A2(new_n20529_), .ZN(new_n20530_));
  NAND2_X1   g20337(.A1(new_n20530_), .A2(new_n13760_), .ZN(new_n20531_));
  INV_X1     g20338(.I(new_n20531_), .ZN(new_n20532_));
  OAI21_X1   g20339(.A1(new_n20527_), .A2(new_n14273_), .B(new_n20532_), .ZN(new_n20533_));
  NAND2_X1   g20340(.A1(new_n20533_), .A2(new_n20526_), .ZN(new_n20534_));
  OAI22_X1   g20341(.A1(new_n20527_), .A2(new_n14273_), .B1(new_n20525_), .B2(new_n20519_), .ZN(new_n20535_));
  NAND2_X1   g20342(.A1(new_n20258_), .A2(\asqrt[17] ), .ZN(new_n20536_));
  NOR4_X1    g20343(.A1(new_n20455_), .A2(\asqrt[17] ), .A3(new_n19884_), .A4(new_n20258_), .ZN(new_n20537_));
  XOR2_X1    g20344(.A1(new_n20537_), .A2(new_n20536_), .Z(new_n20538_));
  NAND2_X1   g20345(.A1(new_n20538_), .A2(new_n13192_), .ZN(new_n20539_));
  AOI21_X1   g20346(.A1(new_n20535_), .A2(\asqrt[17] ), .B(new_n20539_), .ZN(new_n20540_));
  NOR2_X1    g20347(.A1(new_n20540_), .A2(new_n20534_), .ZN(new_n20541_));
  AOI22_X1   g20348(.A1(new_n20535_), .A2(\asqrt[17] ), .B1(new_n20533_), .B2(new_n20526_), .ZN(new_n20542_));
  NAND2_X1   g20349(.A1(new_n19896_), .A2(\asqrt[18] ), .ZN(new_n20543_));
  NOR4_X1    g20350(.A1(new_n20455_), .A2(\asqrt[18] ), .A3(new_n19891_), .A4(new_n19896_), .ZN(new_n20544_));
  XOR2_X1    g20351(.A1(new_n20544_), .A2(new_n20543_), .Z(new_n20545_));
  NAND2_X1   g20352(.A1(new_n20545_), .A2(new_n12657_), .ZN(new_n20546_));
  INV_X1     g20353(.I(new_n20546_), .ZN(new_n20547_));
  OAI21_X1   g20354(.A1(new_n20542_), .A2(new_n13192_), .B(new_n20547_), .ZN(new_n20548_));
  NAND2_X1   g20355(.A1(new_n20548_), .A2(new_n20541_), .ZN(new_n20549_));
  OAI22_X1   g20356(.A1(new_n20542_), .A2(new_n13192_), .B1(new_n20540_), .B2(new_n20534_), .ZN(new_n20550_));
  NOR4_X1    g20357(.A1(new_n20455_), .A2(\asqrt[19] ), .A3(new_n19899_), .A4(new_n20265_), .ZN(new_n20551_));
  AOI21_X1   g20358(.A1(new_n20543_), .A2(new_n19895_), .B(new_n12657_), .ZN(new_n20552_));
  NOR2_X1    g20359(.A1(new_n20551_), .A2(new_n20552_), .ZN(new_n20553_));
  NAND2_X1   g20360(.A1(new_n20553_), .A2(new_n12101_), .ZN(new_n20554_));
  AOI21_X1   g20361(.A1(new_n20550_), .A2(\asqrt[19] ), .B(new_n20554_), .ZN(new_n20555_));
  NOR2_X1    g20362(.A1(new_n20555_), .A2(new_n20549_), .ZN(new_n20556_));
  AOI22_X1   g20363(.A1(new_n20550_), .A2(\asqrt[19] ), .B1(new_n20548_), .B2(new_n20541_), .ZN(new_n20557_));
  NAND2_X1   g20364(.A1(new_n19911_), .A2(\asqrt[20] ), .ZN(new_n20558_));
  NOR4_X1    g20365(.A1(new_n20455_), .A2(\asqrt[20] ), .A3(new_n19906_), .A4(new_n19911_), .ZN(new_n20559_));
  XOR2_X1    g20366(.A1(new_n20559_), .A2(new_n20558_), .Z(new_n20560_));
  NAND2_X1   g20367(.A1(new_n20560_), .A2(new_n11631_), .ZN(new_n20561_));
  INV_X1     g20368(.I(new_n20561_), .ZN(new_n20562_));
  OAI21_X1   g20369(.A1(new_n20557_), .A2(new_n12101_), .B(new_n20562_), .ZN(new_n20563_));
  NAND2_X1   g20370(.A1(new_n20563_), .A2(new_n20556_), .ZN(new_n20564_));
  OAI22_X1   g20371(.A1(new_n20557_), .A2(new_n12101_), .B1(new_n20555_), .B2(new_n20549_), .ZN(new_n20565_));
  NOR4_X1    g20372(.A1(new_n20455_), .A2(\asqrt[21] ), .A3(new_n19914_), .A4(new_n20272_), .ZN(new_n20566_));
  AOI21_X1   g20373(.A1(new_n20558_), .A2(new_n19910_), .B(new_n11631_), .ZN(new_n20567_));
  NOR2_X1    g20374(.A1(new_n20566_), .A2(new_n20567_), .ZN(new_n20568_));
  NAND2_X1   g20375(.A1(new_n20568_), .A2(new_n11105_), .ZN(new_n20569_));
  AOI21_X1   g20376(.A1(new_n20565_), .A2(\asqrt[21] ), .B(new_n20569_), .ZN(new_n20570_));
  NOR2_X1    g20377(.A1(new_n20570_), .A2(new_n20564_), .ZN(new_n20571_));
  AOI22_X1   g20378(.A1(new_n20565_), .A2(\asqrt[21] ), .B1(new_n20563_), .B2(new_n20556_), .ZN(new_n20572_));
  NAND2_X1   g20379(.A1(new_n19926_), .A2(\asqrt[22] ), .ZN(new_n20573_));
  NOR4_X1    g20380(.A1(new_n20455_), .A2(\asqrt[22] ), .A3(new_n19921_), .A4(new_n19926_), .ZN(new_n20574_));
  XOR2_X1    g20381(.A1(new_n20574_), .A2(new_n20573_), .Z(new_n20575_));
  NAND2_X1   g20382(.A1(new_n20575_), .A2(new_n10614_), .ZN(new_n20576_));
  INV_X1     g20383(.I(new_n20576_), .ZN(new_n20577_));
  OAI21_X1   g20384(.A1(new_n20572_), .A2(new_n11105_), .B(new_n20577_), .ZN(new_n20578_));
  NAND2_X1   g20385(.A1(new_n20578_), .A2(new_n20571_), .ZN(new_n20579_));
  OAI22_X1   g20386(.A1(new_n20572_), .A2(new_n11105_), .B1(new_n20570_), .B2(new_n20564_), .ZN(new_n20580_));
  NOR4_X1    g20387(.A1(new_n20455_), .A2(\asqrt[23] ), .A3(new_n19929_), .A4(new_n20279_), .ZN(new_n20581_));
  AOI21_X1   g20388(.A1(new_n20573_), .A2(new_n19925_), .B(new_n10614_), .ZN(new_n20582_));
  NOR2_X1    g20389(.A1(new_n20581_), .A2(new_n20582_), .ZN(new_n20583_));
  NAND2_X1   g20390(.A1(new_n20583_), .A2(new_n10104_), .ZN(new_n20584_));
  AOI21_X1   g20391(.A1(new_n20580_), .A2(\asqrt[23] ), .B(new_n20584_), .ZN(new_n20585_));
  NOR2_X1    g20392(.A1(new_n20585_), .A2(new_n20579_), .ZN(new_n20586_));
  AOI22_X1   g20393(.A1(new_n20580_), .A2(\asqrt[23] ), .B1(new_n20578_), .B2(new_n20571_), .ZN(new_n20587_));
  NAND2_X1   g20394(.A1(new_n19941_), .A2(\asqrt[24] ), .ZN(new_n20588_));
  NOR4_X1    g20395(.A1(new_n20455_), .A2(\asqrt[24] ), .A3(new_n19936_), .A4(new_n19941_), .ZN(new_n20589_));
  XOR2_X1    g20396(.A1(new_n20589_), .A2(new_n20588_), .Z(new_n20590_));
  NAND2_X1   g20397(.A1(new_n20590_), .A2(new_n9672_), .ZN(new_n20591_));
  INV_X1     g20398(.I(new_n20591_), .ZN(new_n20592_));
  OAI21_X1   g20399(.A1(new_n20587_), .A2(new_n10104_), .B(new_n20592_), .ZN(new_n20593_));
  NAND2_X1   g20400(.A1(new_n20593_), .A2(new_n20586_), .ZN(new_n20594_));
  OAI22_X1   g20401(.A1(new_n20587_), .A2(new_n10104_), .B1(new_n20585_), .B2(new_n20579_), .ZN(new_n20595_));
  NOR4_X1    g20402(.A1(new_n20455_), .A2(\asqrt[25] ), .A3(new_n19944_), .A4(new_n20286_), .ZN(new_n20596_));
  AOI21_X1   g20403(.A1(new_n20588_), .A2(new_n19940_), .B(new_n9672_), .ZN(new_n20597_));
  NOR2_X1    g20404(.A1(new_n20596_), .A2(new_n20597_), .ZN(new_n20598_));
  NAND2_X1   g20405(.A1(new_n20598_), .A2(new_n9212_), .ZN(new_n20599_));
  AOI21_X1   g20406(.A1(new_n20595_), .A2(\asqrt[25] ), .B(new_n20599_), .ZN(new_n20600_));
  NOR2_X1    g20407(.A1(new_n20600_), .A2(new_n20594_), .ZN(new_n20601_));
  AOI22_X1   g20408(.A1(new_n20595_), .A2(\asqrt[25] ), .B1(new_n20593_), .B2(new_n20586_), .ZN(new_n20602_));
  NAND2_X1   g20409(.A1(new_n19956_), .A2(\asqrt[26] ), .ZN(new_n20603_));
  NOR4_X1    g20410(.A1(new_n20455_), .A2(\asqrt[26] ), .A3(new_n19951_), .A4(new_n19956_), .ZN(new_n20604_));
  XOR2_X1    g20411(.A1(new_n20604_), .A2(new_n20603_), .Z(new_n20605_));
  NAND2_X1   g20412(.A1(new_n20605_), .A2(new_n8763_), .ZN(new_n20606_));
  INV_X1     g20413(.I(new_n20606_), .ZN(new_n20607_));
  OAI21_X1   g20414(.A1(new_n20602_), .A2(new_n9212_), .B(new_n20607_), .ZN(new_n20608_));
  NAND2_X1   g20415(.A1(new_n20608_), .A2(new_n20601_), .ZN(new_n20609_));
  OAI22_X1   g20416(.A1(new_n20602_), .A2(new_n9212_), .B1(new_n20600_), .B2(new_n20594_), .ZN(new_n20610_));
  NAND2_X1   g20417(.A1(new_n20293_), .A2(\asqrt[27] ), .ZN(new_n20611_));
  NOR4_X1    g20418(.A1(new_n20455_), .A2(\asqrt[27] ), .A3(new_n19959_), .A4(new_n20293_), .ZN(new_n20612_));
  XOR2_X1    g20419(.A1(new_n20612_), .A2(new_n20611_), .Z(new_n20613_));
  NAND2_X1   g20420(.A1(new_n20613_), .A2(new_n8319_), .ZN(new_n20614_));
  AOI21_X1   g20421(.A1(new_n20610_), .A2(\asqrt[27] ), .B(new_n20614_), .ZN(new_n20615_));
  NOR2_X1    g20422(.A1(new_n20615_), .A2(new_n20609_), .ZN(new_n20616_));
  AOI22_X1   g20423(.A1(new_n20610_), .A2(\asqrt[27] ), .B1(new_n20608_), .B2(new_n20601_), .ZN(new_n20617_));
  NOR4_X1    g20424(.A1(new_n20455_), .A2(\asqrt[28] ), .A3(new_n19966_), .A4(new_n19971_), .ZN(new_n20618_));
  AOI21_X1   g20425(.A1(new_n20611_), .A2(new_n20292_), .B(new_n8319_), .ZN(new_n20619_));
  NOR2_X1    g20426(.A1(new_n20618_), .A2(new_n20619_), .ZN(new_n20620_));
  NAND2_X1   g20427(.A1(new_n20620_), .A2(new_n7931_), .ZN(new_n20621_));
  INV_X1     g20428(.I(new_n20621_), .ZN(new_n20622_));
  OAI21_X1   g20429(.A1(new_n20617_), .A2(new_n8319_), .B(new_n20622_), .ZN(new_n20623_));
  NAND2_X1   g20430(.A1(new_n20623_), .A2(new_n20616_), .ZN(new_n20624_));
  OAI22_X1   g20431(.A1(new_n20617_), .A2(new_n8319_), .B1(new_n20615_), .B2(new_n20609_), .ZN(new_n20625_));
  NAND2_X1   g20432(.A1(new_n20300_), .A2(\asqrt[29] ), .ZN(new_n20626_));
  NOR4_X1    g20433(.A1(new_n20455_), .A2(\asqrt[29] ), .A3(new_n19974_), .A4(new_n20300_), .ZN(new_n20627_));
  XOR2_X1    g20434(.A1(new_n20627_), .A2(new_n20626_), .Z(new_n20628_));
  NAND2_X1   g20435(.A1(new_n20628_), .A2(new_n7517_), .ZN(new_n20629_));
  AOI21_X1   g20436(.A1(new_n20625_), .A2(\asqrt[29] ), .B(new_n20629_), .ZN(new_n20630_));
  NOR2_X1    g20437(.A1(new_n20630_), .A2(new_n20624_), .ZN(new_n20631_));
  AOI22_X1   g20438(.A1(new_n20625_), .A2(\asqrt[29] ), .B1(new_n20623_), .B2(new_n20616_), .ZN(new_n20632_));
  NOR4_X1    g20439(.A1(new_n20455_), .A2(\asqrt[30] ), .A3(new_n19981_), .A4(new_n19986_), .ZN(new_n20633_));
  AOI21_X1   g20440(.A1(new_n20626_), .A2(new_n20299_), .B(new_n7517_), .ZN(new_n20634_));
  NOR2_X1    g20441(.A1(new_n20633_), .A2(new_n20634_), .ZN(new_n20635_));
  NAND2_X1   g20442(.A1(new_n20635_), .A2(new_n7110_), .ZN(new_n20636_));
  INV_X1     g20443(.I(new_n20636_), .ZN(new_n20637_));
  OAI21_X1   g20444(.A1(new_n20632_), .A2(new_n7517_), .B(new_n20637_), .ZN(new_n20638_));
  NAND2_X1   g20445(.A1(new_n20638_), .A2(new_n20631_), .ZN(new_n20639_));
  OAI22_X1   g20446(.A1(new_n20632_), .A2(new_n7517_), .B1(new_n20630_), .B2(new_n20624_), .ZN(new_n20640_));
  NAND2_X1   g20447(.A1(new_n20307_), .A2(\asqrt[31] ), .ZN(new_n20641_));
  NOR4_X1    g20448(.A1(new_n20455_), .A2(\asqrt[31] ), .A3(new_n19989_), .A4(new_n20307_), .ZN(new_n20642_));
  XOR2_X1    g20449(.A1(new_n20642_), .A2(new_n20641_), .Z(new_n20643_));
  NAND2_X1   g20450(.A1(new_n20643_), .A2(new_n6708_), .ZN(new_n20644_));
  AOI21_X1   g20451(.A1(new_n20640_), .A2(\asqrt[31] ), .B(new_n20644_), .ZN(new_n20645_));
  NOR2_X1    g20452(.A1(new_n20645_), .A2(new_n20639_), .ZN(new_n20646_));
  AOI22_X1   g20453(.A1(new_n20640_), .A2(\asqrt[31] ), .B1(new_n20638_), .B2(new_n20631_), .ZN(new_n20647_));
  NOR4_X1    g20454(.A1(new_n20455_), .A2(\asqrt[32] ), .A3(new_n19996_), .A4(new_n20001_), .ZN(new_n20648_));
  AOI21_X1   g20455(.A1(new_n20641_), .A2(new_n20306_), .B(new_n6708_), .ZN(new_n20649_));
  NOR2_X1    g20456(.A1(new_n20648_), .A2(new_n20649_), .ZN(new_n20650_));
  NAND2_X1   g20457(.A1(new_n20650_), .A2(new_n6365_), .ZN(new_n20651_));
  INV_X1     g20458(.I(new_n20651_), .ZN(new_n20652_));
  OAI21_X1   g20459(.A1(new_n20647_), .A2(new_n6708_), .B(new_n20652_), .ZN(new_n20653_));
  NAND2_X1   g20460(.A1(new_n20653_), .A2(new_n20646_), .ZN(new_n20654_));
  OAI22_X1   g20461(.A1(new_n20647_), .A2(new_n6708_), .B1(new_n20645_), .B2(new_n20639_), .ZN(new_n20655_));
  NAND2_X1   g20462(.A1(new_n20314_), .A2(\asqrt[33] ), .ZN(new_n20656_));
  NOR4_X1    g20463(.A1(new_n20455_), .A2(\asqrt[33] ), .A3(new_n20004_), .A4(new_n20314_), .ZN(new_n20657_));
  XOR2_X1    g20464(.A1(new_n20657_), .A2(new_n20656_), .Z(new_n20658_));
  NAND2_X1   g20465(.A1(new_n20658_), .A2(new_n5991_), .ZN(new_n20659_));
  AOI21_X1   g20466(.A1(new_n20655_), .A2(\asqrt[33] ), .B(new_n20659_), .ZN(new_n20660_));
  NOR2_X1    g20467(.A1(new_n20660_), .A2(new_n20654_), .ZN(new_n20661_));
  AOI22_X1   g20468(.A1(new_n20655_), .A2(\asqrt[33] ), .B1(new_n20653_), .B2(new_n20646_), .ZN(new_n20662_));
  NOR4_X1    g20469(.A1(new_n20455_), .A2(\asqrt[34] ), .A3(new_n20011_), .A4(new_n20016_), .ZN(new_n20663_));
  AOI21_X1   g20470(.A1(new_n20656_), .A2(new_n20313_), .B(new_n5991_), .ZN(new_n20664_));
  NOR2_X1    g20471(.A1(new_n20663_), .A2(new_n20664_), .ZN(new_n20665_));
  NAND2_X1   g20472(.A1(new_n20665_), .A2(new_n5626_), .ZN(new_n20666_));
  INV_X1     g20473(.I(new_n20666_), .ZN(new_n20667_));
  OAI21_X1   g20474(.A1(new_n20662_), .A2(new_n5991_), .B(new_n20667_), .ZN(new_n20668_));
  NAND2_X1   g20475(.A1(new_n20668_), .A2(new_n20661_), .ZN(new_n20669_));
  OAI22_X1   g20476(.A1(new_n20662_), .A2(new_n5991_), .B1(new_n20660_), .B2(new_n20654_), .ZN(new_n20670_));
  NAND2_X1   g20477(.A1(new_n20321_), .A2(\asqrt[35] ), .ZN(new_n20671_));
  NOR4_X1    g20478(.A1(new_n20455_), .A2(\asqrt[35] ), .A3(new_n20019_), .A4(new_n20321_), .ZN(new_n20672_));
  XOR2_X1    g20479(.A1(new_n20672_), .A2(new_n20671_), .Z(new_n20673_));
  NAND2_X1   g20480(.A1(new_n20673_), .A2(new_n5273_), .ZN(new_n20674_));
  AOI21_X1   g20481(.A1(new_n20670_), .A2(\asqrt[35] ), .B(new_n20674_), .ZN(new_n20675_));
  NOR2_X1    g20482(.A1(new_n20675_), .A2(new_n20669_), .ZN(new_n20676_));
  AOI22_X1   g20483(.A1(new_n20670_), .A2(\asqrt[35] ), .B1(new_n20668_), .B2(new_n20661_), .ZN(new_n20677_));
  NOR4_X1    g20484(.A1(new_n20455_), .A2(\asqrt[36] ), .A3(new_n20026_), .A4(new_n20031_), .ZN(new_n20678_));
  AOI21_X1   g20485(.A1(new_n20671_), .A2(new_n20320_), .B(new_n5273_), .ZN(new_n20679_));
  NOR2_X1    g20486(.A1(new_n20678_), .A2(new_n20679_), .ZN(new_n20680_));
  NAND2_X1   g20487(.A1(new_n20680_), .A2(new_n4973_), .ZN(new_n20681_));
  INV_X1     g20488(.I(new_n20681_), .ZN(new_n20682_));
  OAI21_X1   g20489(.A1(new_n20677_), .A2(new_n5273_), .B(new_n20682_), .ZN(new_n20683_));
  NAND2_X1   g20490(.A1(new_n20683_), .A2(new_n20676_), .ZN(new_n20684_));
  OAI22_X1   g20491(.A1(new_n20677_), .A2(new_n5273_), .B1(new_n20675_), .B2(new_n20669_), .ZN(new_n20685_));
  NAND2_X1   g20492(.A1(new_n20328_), .A2(\asqrt[37] ), .ZN(new_n20686_));
  NOR4_X1    g20493(.A1(new_n20455_), .A2(\asqrt[37] ), .A3(new_n20034_), .A4(new_n20328_), .ZN(new_n20687_));
  XOR2_X1    g20494(.A1(new_n20687_), .A2(new_n20686_), .Z(new_n20688_));
  NAND2_X1   g20495(.A1(new_n20688_), .A2(new_n4645_), .ZN(new_n20689_));
  AOI21_X1   g20496(.A1(new_n20685_), .A2(\asqrt[37] ), .B(new_n20689_), .ZN(new_n20690_));
  NOR2_X1    g20497(.A1(new_n20690_), .A2(new_n20684_), .ZN(new_n20691_));
  AOI22_X1   g20498(.A1(new_n20685_), .A2(\asqrt[37] ), .B1(new_n20683_), .B2(new_n20676_), .ZN(new_n20692_));
  NOR4_X1    g20499(.A1(new_n20455_), .A2(\asqrt[38] ), .A3(new_n20041_), .A4(new_n20046_), .ZN(new_n20693_));
  AOI21_X1   g20500(.A1(new_n20686_), .A2(new_n20327_), .B(new_n4645_), .ZN(new_n20694_));
  NOR2_X1    g20501(.A1(new_n20693_), .A2(new_n20694_), .ZN(new_n20695_));
  NAND2_X1   g20502(.A1(new_n20695_), .A2(new_n4330_), .ZN(new_n20696_));
  INV_X1     g20503(.I(new_n20696_), .ZN(new_n20697_));
  OAI21_X1   g20504(.A1(new_n20692_), .A2(new_n4645_), .B(new_n20697_), .ZN(new_n20698_));
  NAND2_X1   g20505(.A1(new_n20698_), .A2(new_n20691_), .ZN(new_n20699_));
  OAI22_X1   g20506(.A1(new_n20692_), .A2(new_n4645_), .B1(new_n20690_), .B2(new_n20684_), .ZN(new_n20700_));
  NAND2_X1   g20507(.A1(new_n20335_), .A2(\asqrt[39] ), .ZN(new_n20701_));
  NOR4_X1    g20508(.A1(new_n20455_), .A2(\asqrt[39] ), .A3(new_n20049_), .A4(new_n20335_), .ZN(new_n20702_));
  XOR2_X1    g20509(.A1(new_n20702_), .A2(new_n20701_), .Z(new_n20703_));
  NAND2_X1   g20510(.A1(new_n20703_), .A2(new_n4018_), .ZN(new_n20704_));
  AOI21_X1   g20511(.A1(new_n20700_), .A2(\asqrt[39] ), .B(new_n20704_), .ZN(new_n20705_));
  NOR2_X1    g20512(.A1(new_n20705_), .A2(new_n20699_), .ZN(new_n20706_));
  AOI22_X1   g20513(.A1(new_n20700_), .A2(\asqrt[39] ), .B1(new_n20698_), .B2(new_n20691_), .ZN(new_n20707_));
  NOR4_X1    g20514(.A1(new_n20455_), .A2(\asqrt[40] ), .A3(new_n20056_), .A4(new_n20061_), .ZN(new_n20708_));
  AOI21_X1   g20515(.A1(new_n20701_), .A2(new_n20334_), .B(new_n4018_), .ZN(new_n20709_));
  NOR2_X1    g20516(.A1(new_n20708_), .A2(new_n20709_), .ZN(new_n20710_));
  NAND2_X1   g20517(.A1(new_n20710_), .A2(new_n3760_), .ZN(new_n20711_));
  INV_X1     g20518(.I(new_n20711_), .ZN(new_n20712_));
  OAI21_X1   g20519(.A1(new_n20707_), .A2(new_n4018_), .B(new_n20712_), .ZN(new_n20713_));
  NAND2_X1   g20520(.A1(new_n20713_), .A2(new_n20706_), .ZN(new_n20714_));
  OAI22_X1   g20521(.A1(new_n20707_), .A2(new_n4018_), .B1(new_n20705_), .B2(new_n20699_), .ZN(new_n20715_));
  NAND2_X1   g20522(.A1(new_n20342_), .A2(\asqrt[41] ), .ZN(new_n20716_));
  NOR4_X1    g20523(.A1(new_n20455_), .A2(\asqrt[41] ), .A3(new_n20064_), .A4(new_n20342_), .ZN(new_n20717_));
  XOR2_X1    g20524(.A1(new_n20717_), .A2(new_n20716_), .Z(new_n20718_));
  NAND2_X1   g20525(.A1(new_n20718_), .A2(new_n3481_), .ZN(new_n20719_));
  AOI21_X1   g20526(.A1(new_n20715_), .A2(\asqrt[41] ), .B(new_n20719_), .ZN(new_n20720_));
  NOR2_X1    g20527(.A1(new_n20720_), .A2(new_n20714_), .ZN(new_n20721_));
  AOI22_X1   g20528(.A1(new_n20715_), .A2(\asqrt[41] ), .B1(new_n20713_), .B2(new_n20706_), .ZN(new_n20722_));
  NOR4_X1    g20529(.A1(new_n20455_), .A2(\asqrt[42] ), .A3(new_n20071_), .A4(new_n20076_), .ZN(new_n20723_));
  AOI21_X1   g20530(.A1(new_n20716_), .A2(new_n20341_), .B(new_n3481_), .ZN(new_n20724_));
  NOR2_X1    g20531(.A1(new_n20723_), .A2(new_n20724_), .ZN(new_n20725_));
  NAND2_X1   g20532(.A1(new_n20725_), .A2(new_n3208_), .ZN(new_n20726_));
  INV_X1     g20533(.I(new_n20726_), .ZN(new_n20727_));
  OAI21_X1   g20534(.A1(new_n20722_), .A2(new_n3481_), .B(new_n20727_), .ZN(new_n20728_));
  NAND2_X1   g20535(.A1(new_n20728_), .A2(new_n20721_), .ZN(new_n20729_));
  OAI22_X1   g20536(.A1(new_n20722_), .A2(new_n3481_), .B1(new_n20720_), .B2(new_n20714_), .ZN(new_n20730_));
  NAND2_X1   g20537(.A1(new_n20349_), .A2(\asqrt[43] ), .ZN(new_n20731_));
  NOR4_X1    g20538(.A1(new_n20455_), .A2(\asqrt[43] ), .A3(new_n20079_), .A4(new_n20349_), .ZN(new_n20732_));
  XOR2_X1    g20539(.A1(new_n20732_), .A2(new_n20731_), .Z(new_n20733_));
  NAND2_X1   g20540(.A1(new_n20733_), .A2(new_n2941_), .ZN(new_n20734_));
  AOI21_X1   g20541(.A1(new_n20730_), .A2(\asqrt[43] ), .B(new_n20734_), .ZN(new_n20735_));
  NOR2_X1    g20542(.A1(new_n20735_), .A2(new_n20729_), .ZN(new_n20736_));
  AOI22_X1   g20543(.A1(new_n20730_), .A2(\asqrt[43] ), .B1(new_n20728_), .B2(new_n20721_), .ZN(new_n20737_));
  NOR4_X1    g20544(.A1(new_n20455_), .A2(\asqrt[44] ), .A3(new_n20086_), .A4(new_n20091_), .ZN(new_n20738_));
  AOI21_X1   g20545(.A1(new_n20731_), .A2(new_n20348_), .B(new_n2941_), .ZN(new_n20739_));
  NOR2_X1    g20546(.A1(new_n20738_), .A2(new_n20739_), .ZN(new_n20740_));
  NAND2_X1   g20547(.A1(new_n20740_), .A2(new_n2728_), .ZN(new_n20741_));
  INV_X1     g20548(.I(new_n20741_), .ZN(new_n20742_));
  OAI21_X1   g20549(.A1(new_n20737_), .A2(new_n2941_), .B(new_n20742_), .ZN(new_n20743_));
  NAND2_X1   g20550(.A1(new_n20743_), .A2(new_n20736_), .ZN(new_n20744_));
  OAI22_X1   g20551(.A1(new_n20737_), .A2(new_n2941_), .B1(new_n20735_), .B2(new_n20729_), .ZN(new_n20745_));
  NAND2_X1   g20552(.A1(new_n20356_), .A2(\asqrt[45] ), .ZN(new_n20746_));
  NOR4_X1    g20553(.A1(new_n20455_), .A2(\asqrt[45] ), .A3(new_n20094_), .A4(new_n20356_), .ZN(new_n20747_));
  XOR2_X1    g20554(.A1(new_n20747_), .A2(new_n20746_), .Z(new_n20748_));
  NAND2_X1   g20555(.A1(new_n20748_), .A2(new_n2488_), .ZN(new_n20749_));
  AOI21_X1   g20556(.A1(new_n20745_), .A2(\asqrt[45] ), .B(new_n20749_), .ZN(new_n20750_));
  NOR2_X1    g20557(.A1(new_n20750_), .A2(new_n20744_), .ZN(new_n20751_));
  AOI22_X1   g20558(.A1(new_n20745_), .A2(\asqrt[45] ), .B1(new_n20743_), .B2(new_n20736_), .ZN(new_n20752_));
  NOR4_X1    g20559(.A1(new_n20455_), .A2(\asqrt[46] ), .A3(new_n20101_), .A4(new_n20106_), .ZN(new_n20753_));
  AOI21_X1   g20560(.A1(new_n20746_), .A2(new_n20355_), .B(new_n2488_), .ZN(new_n20754_));
  NOR2_X1    g20561(.A1(new_n20753_), .A2(new_n20754_), .ZN(new_n20755_));
  NAND2_X1   g20562(.A1(new_n20755_), .A2(new_n2253_), .ZN(new_n20756_));
  INV_X1     g20563(.I(new_n20756_), .ZN(new_n20757_));
  OAI21_X1   g20564(.A1(new_n20752_), .A2(new_n2488_), .B(new_n20757_), .ZN(new_n20758_));
  NAND2_X1   g20565(.A1(new_n20758_), .A2(new_n20751_), .ZN(new_n20759_));
  OAI22_X1   g20566(.A1(new_n20752_), .A2(new_n2488_), .B1(new_n20750_), .B2(new_n20744_), .ZN(new_n20760_));
  NAND2_X1   g20567(.A1(new_n20363_), .A2(\asqrt[47] ), .ZN(new_n20761_));
  NOR4_X1    g20568(.A1(new_n20455_), .A2(\asqrt[47] ), .A3(new_n20109_), .A4(new_n20363_), .ZN(new_n20762_));
  XOR2_X1    g20569(.A1(new_n20762_), .A2(new_n20761_), .Z(new_n20763_));
  NAND2_X1   g20570(.A1(new_n20763_), .A2(new_n2046_), .ZN(new_n20764_));
  AOI21_X1   g20571(.A1(new_n20760_), .A2(\asqrt[47] ), .B(new_n20764_), .ZN(new_n20765_));
  NOR2_X1    g20572(.A1(new_n20765_), .A2(new_n20759_), .ZN(new_n20766_));
  AOI22_X1   g20573(.A1(new_n20760_), .A2(\asqrt[47] ), .B1(new_n20758_), .B2(new_n20751_), .ZN(new_n20767_));
  NOR4_X1    g20574(.A1(new_n20455_), .A2(\asqrt[48] ), .A3(new_n20116_), .A4(new_n20121_), .ZN(new_n20768_));
  AOI21_X1   g20575(.A1(new_n20761_), .A2(new_n20362_), .B(new_n2046_), .ZN(new_n20769_));
  NOR2_X1    g20576(.A1(new_n20768_), .A2(new_n20769_), .ZN(new_n20770_));
  NAND2_X1   g20577(.A1(new_n20770_), .A2(new_n1854_), .ZN(new_n20771_));
  INV_X1     g20578(.I(new_n20771_), .ZN(new_n20772_));
  OAI21_X1   g20579(.A1(new_n20767_), .A2(new_n2046_), .B(new_n20772_), .ZN(new_n20773_));
  NAND2_X1   g20580(.A1(new_n20773_), .A2(new_n20766_), .ZN(new_n20774_));
  OAI22_X1   g20581(.A1(new_n20767_), .A2(new_n2046_), .B1(new_n20765_), .B2(new_n20759_), .ZN(new_n20775_));
  NAND2_X1   g20582(.A1(new_n20370_), .A2(\asqrt[49] ), .ZN(new_n20776_));
  NOR4_X1    g20583(.A1(new_n20455_), .A2(\asqrt[49] ), .A3(new_n20124_), .A4(new_n20370_), .ZN(new_n20777_));
  XOR2_X1    g20584(.A1(new_n20777_), .A2(new_n20776_), .Z(new_n20778_));
  NAND2_X1   g20585(.A1(new_n20778_), .A2(new_n1595_), .ZN(new_n20779_));
  AOI21_X1   g20586(.A1(new_n20775_), .A2(\asqrt[49] ), .B(new_n20779_), .ZN(new_n20780_));
  NOR2_X1    g20587(.A1(new_n20780_), .A2(new_n20774_), .ZN(new_n20781_));
  AOI22_X1   g20588(.A1(new_n20775_), .A2(\asqrt[49] ), .B1(new_n20773_), .B2(new_n20766_), .ZN(new_n20782_));
  NOR4_X1    g20589(.A1(new_n20455_), .A2(\asqrt[50] ), .A3(new_n20131_), .A4(new_n20136_), .ZN(new_n20783_));
  AOI21_X1   g20590(.A1(new_n20776_), .A2(new_n20369_), .B(new_n1595_), .ZN(new_n20784_));
  NOR2_X1    g20591(.A1(new_n20783_), .A2(new_n20784_), .ZN(new_n20785_));
  NAND2_X1   g20592(.A1(new_n20785_), .A2(new_n1436_), .ZN(new_n20786_));
  INV_X1     g20593(.I(new_n20786_), .ZN(new_n20787_));
  OAI21_X1   g20594(.A1(new_n20782_), .A2(new_n1595_), .B(new_n20787_), .ZN(new_n20788_));
  NAND2_X1   g20595(.A1(new_n20788_), .A2(new_n20781_), .ZN(new_n20789_));
  OAI22_X1   g20596(.A1(new_n20782_), .A2(new_n1595_), .B1(new_n20780_), .B2(new_n20774_), .ZN(new_n20790_));
  NAND2_X1   g20597(.A1(new_n20377_), .A2(\asqrt[51] ), .ZN(new_n20791_));
  NOR4_X1    g20598(.A1(new_n20455_), .A2(\asqrt[51] ), .A3(new_n20139_), .A4(new_n20377_), .ZN(new_n20792_));
  XOR2_X1    g20599(.A1(new_n20792_), .A2(new_n20791_), .Z(new_n20793_));
  NAND2_X1   g20600(.A1(new_n20793_), .A2(new_n1260_), .ZN(new_n20794_));
  AOI21_X1   g20601(.A1(new_n20790_), .A2(\asqrt[51] ), .B(new_n20794_), .ZN(new_n20795_));
  NOR2_X1    g20602(.A1(new_n20795_), .A2(new_n20789_), .ZN(new_n20796_));
  AOI22_X1   g20603(.A1(new_n20790_), .A2(\asqrt[51] ), .B1(new_n20788_), .B2(new_n20781_), .ZN(new_n20797_));
  NOR4_X1    g20604(.A1(new_n20455_), .A2(\asqrt[52] ), .A3(new_n20146_), .A4(new_n20151_), .ZN(new_n20798_));
  AOI21_X1   g20605(.A1(new_n20791_), .A2(new_n20376_), .B(new_n1260_), .ZN(new_n20799_));
  NOR2_X1    g20606(.A1(new_n20798_), .A2(new_n20799_), .ZN(new_n20800_));
  NAND2_X1   g20607(.A1(new_n20800_), .A2(new_n1096_), .ZN(new_n20801_));
  INV_X1     g20608(.I(new_n20801_), .ZN(new_n20802_));
  OAI21_X1   g20609(.A1(new_n20797_), .A2(new_n1260_), .B(new_n20802_), .ZN(new_n20803_));
  NAND2_X1   g20610(.A1(new_n20803_), .A2(new_n20796_), .ZN(new_n20804_));
  OAI22_X1   g20611(.A1(new_n20797_), .A2(new_n1260_), .B1(new_n20795_), .B2(new_n20789_), .ZN(new_n20805_));
  NAND2_X1   g20612(.A1(new_n20384_), .A2(\asqrt[53] ), .ZN(new_n20806_));
  NOR4_X1    g20613(.A1(new_n20455_), .A2(\asqrt[53] ), .A3(new_n20154_), .A4(new_n20384_), .ZN(new_n20807_));
  XOR2_X1    g20614(.A1(new_n20807_), .A2(new_n20806_), .Z(new_n20808_));
  NAND2_X1   g20615(.A1(new_n20808_), .A2(new_n970_), .ZN(new_n20809_));
  AOI21_X1   g20616(.A1(new_n20805_), .A2(\asqrt[53] ), .B(new_n20809_), .ZN(new_n20810_));
  NOR2_X1    g20617(.A1(new_n20810_), .A2(new_n20804_), .ZN(new_n20811_));
  AOI22_X1   g20618(.A1(new_n20805_), .A2(\asqrt[53] ), .B1(new_n20803_), .B2(new_n20796_), .ZN(new_n20812_));
  NOR4_X1    g20619(.A1(new_n20455_), .A2(\asqrt[54] ), .A3(new_n20161_), .A4(new_n20166_), .ZN(new_n20813_));
  AOI21_X1   g20620(.A1(new_n20806_), .A2(new_n20383_), .B(new_n970_), .ZN(new_n20814_));
  NOR2_X1    g20621(.A1(new_n20813_), .A2(new_n20814_), .ZN(new_n20815_));
  NAND2_X1   g20622(.A1(new_n20815_), .A2(new_n825_), .ZN(new_n20816_));
  INV_X1     g20623(.I(new_n20816_), .ZN(new_n20817_));
  OAI21_X1   g20624(.A1(new_n20812_), .A2(new_n970_), .B(new_n20817_), .ZN(new_n20818_));
  NAND2_X1   g20625(.A1(new_n20818_), .A2(new_n20811_), .ZN(new_n20819_));
  OAI22_X1   g20626(.A1(new_n20812_), .A2(new_n970_), .B1(new_n20810_), .B2(new_n20804_), .ZN(new_n20820_));
  NAND2_X1   g20627(.A1(new_n20391_), .A2(\asqrt[55] ), .ZN(new_n20821_));
  NOR4_X1    g20628(.A1(new_n20455_), .A2(\asqrt[55] ), .A3(new_n20168_), .A4(new_n20391_), .ZN(new_n20822_));
  XOR2_X1    g20629(.A1(new_n20822_), .A2(new_n20821_), .Z(new_n20823_));
  NAND2_X1   g20630(.A1(new_n20823_), .A2(new_n724_), .ZN(new_n20824_));
  AOI21_X1   g20631(.A1(new_n20820_), .A2(\asqrt[55] ), .B(new_n20824_), .ZN(new_n20825_));
  NOR2_X1    g20632(.A1(new_n20825_), .A2(new_n20819_), .ZN(new_n20826_));
  AOI22_X1   g20633(.A1(new_n20820_), .A2(\asqrt[55] ), .B1(new_n20818_), .B2(new_n20811_), .ZN(new_n20827_));
  NOR4_X1    g20634(.A1(new_n20455_), .A2(\asqrt[56] ), .A3(new_n20174_), .A4(new_n20179_), .ZN(new_n20828_));
  AOI21_X1   g20635(.A1(new_n20821_), .A2(new_n20390_), .B(new_n724_), .ZN(new_n20829_));
  NOR2_X1    g20636(.A1(new_n20828_), .A2(new_n20829_), .ZN(new_n20830_));
  NAND2_X1   g20637(.A1(new_n20830_), .A2(new_n587_), .ZN(new_n20831_));
  INV_X1     g20638(.I(new_n20831_), .ZN(new_n20832_));
  OAI21_X1   g20639(.A1(new_n20827_), .A2(new_n724_), .B(new_n20832_), .ZN(new_n20833_));
  NAND2_X1   g20640(.A1(new_n20833_), .A2(new_n20826_), .ZN(new_n20834_));
  OAI22_X1   g20641(.A1(new_n20827_), .A2(new_n724_), .B1(new_n20825_), .B2(new_n20819_), .ZN(new_n20835_));
  NAND2_X1   g20642(.A1(new_n20398_), .A2(\asqrt[57] ), .ZN(new_n20836_));
  NOR4_X1    g20643(.A1(new_n20455_), .A2(\asqrt[57] ), .A3(new_n20181_), .A4(new_n20398_), .ZN(new_n20837_));
  XOR2_X1    g20644(.A1(new_n20837_), .A2(new_n20836_), .Z(new_n20838_));
  NAND2_X1   g20645(.A1(new_n20838_), .A2(new_n504_), .ZN(new_n20839_));
  AOI21_X1   g20646(.A1(new_n20835_), .A2(\asqrt[57] ), .B(new_n20839_), .ZN(new_n20840_));
  NOR2_X1    g20647(.A1(new_n20840_), .A2(new_n20834_), .ZN(new_n20841_));
  AOI22_X1   g20648(.A1(new_n20835_), .A2(\asqrt[57] ), .B1(new_n20833_), .B2(new_n20826_), .ZN(new_n20842_));
  NOR4_X1    g20649(.A1(new_n20455_), .A2(\asqrt[58] ), .A3(new_n20187_), .A4(new_n20192_), .ZN(new_n20843_));
  XOR2_X1    g20650(.A1(new_n20843_), .A2(new_n20198_), .Z(new_n20844_));
  NAND2_X1   g20651(.A1(new_n20844_), .A2(new_n376_), .ZN(new_n20845_));
  INV_X1     g20652(.I(new_n20845_), .ZN(new_n20846_));
  OAI21_X1   g20653(.A1(new_n20842_), .A2(new_n504_), .B(new_n20846_), .ZN(new_n20847_));
  NAND2_X1   g20654(.A1(new_n20847_), .A2(new_n20841_), .ZN(new_n20848_));
  OAI22_X1   g20655(.A1(new_n20842_), .A2(new_n504_), .B1(new_n20840_), .B2(new_n20834_), .ZN(new_n20849_));
  NOR4_X1    g20656(.A1(new_n20455_), .A2(\asqrt[59] ), .A3(new_n20194_), .A4(new_n20405_), .ZN(new_n20850_));
  XOR2_X1    g20657(.A1(new_n20850_), .A2(new_n20425_), .Z(new_n20851_));
  NAND2_X1   g20658(.A1(new_n20851_), .A2(new_n275_), .ZN(new_n20852_));
  AOI21_X1   g20659(.A1(new_n20849_), .A2(\asqrt[59] ), .B(new_n20852_), .ZN(new_n20853_));
  NOR2_X1    g20660(.A1(new_n20853_), .A2(new_n20848_), .ZN(new_n20854_));
  AOI22_X1   g20661(.A1(new_n20849_), .A2(\asqrt[59] ), .B1(new_n20847_), .B2(new_n20841_), .ZN(new_n20855_));
  OAI22_X1   g20662(.A1(new_n20855_), .A2(new_n275_), .B1(new_n20853_), .B2(new_n20848_), .ZN(new_n20856_));
  NOR4_X1    g20663(.A1(new_n20455_), .A2(\asqrt[60] ), .A3(new_n20201_), .A4(new_n20207_), .ZN(new_n20857_));
  XOR2_X1    g20664(.A1(new_n20857_), .A2(new_n20204_), .Z(new_n20858_));
  NAND2_X1   g20665(.A1(new_n20858_), .A2(new_n229_), .ZN(new_n20859_));
  INV_X1     g20666(.I(new_n20859_), .ZN(new_n20860_));
  OAI21_X1   g20667(.A1(new_n20855_), .A2(new_n275_), .B(new_n20860_), .ZN(new_n20861_));
  AOI22_X1   g20668(.A1(new_n20856_), .A2(\asqrt[61] ), .B1(new_n20861_), .B2(new_n20854_), .ZN(new_n20862_));
  NOR2_X1    g20669(.A1(new_n20862_), .A2(new_n196_), .ZN(new_n20863_));
  OAI21_X1   g20670(.A1(new_n20437_), .A2(new_n20421_), .B(new_n19762_), .ZN(new_n20864_));
  NAND3_X1   g20671(.A1(new_n20419_), .A2(\a[12] ), .A3(new_n19763_), .ZN(new_n20865_));
  NAND2_X1   g20672(.A1(new_n20864_), .A2(new_n20865_), .ZN(new_n20866_));
  INV_X1     g20673(.I(new_n20444_), .ZN(new_n20867_));
  NAND3_X1   g20674(.A1(new_n20457_), .A2(new_n20455_), .A3(new_n19791_), .ZN(new_n20868_));
  OAI21_X1   g20675(.A1(new_n20450_), .A2(new_n19792_), .B(\asqrt[6] ), .ZN(new_n20869_));
  NAND4_X1   g20676(.A1(new_n20869_), .A2(new_n20868_), .A3(new_n19100_), .A4(new_n20867_), .ZN(new_n20870_));
  NAND2_X1   g20677(.A1(new_n20870_), .A2(new_n20866_), .ZN(new_n20871_));
  NAND3_X1   g20678(.A1(new_n20864_), .A2(new_n20865_), .A3(new_n20867_), .ZN(new_n20872_));
  NAND3_X1   g20679(.A1(\asqrt[6] ), .A2(new_n20223_), .A3(new_n20467_), .ZN(new_n20873_));
  OAI21_X1   g20680(.A1(new_n20455_), .A2(new_n20465_), .B(new_n19808_), .ZN(new_n20874_));
  NAND3_X1   g20681(.A1(new_n20874_), .A2(new_n20873_), .A3(new_n18495_), .ZN(new_n20875_));
  AOI21_X1   g20682(.A1(new_n20872_), .A2(\asqrt[8] ), .B(new_n20875_), .ZN(new_n20876_));
  NOR2_X1    g20683(.A1(new_n20876_), .A2(new_n20871_), .ZN(new_n20877_));
  AOI22_X1   g20684(.A1(new_n20866_), .A2(new_n20870_), .B1(new_n20872_), .B2(\asqrt[8] ), .ZN(new_n20878_));
  INV_X1     g20685(.I(new_n20477_), .ZN(new_n20879_));
  OAI21_X1   g20686(.A1(new_n20878_), .A2(new_n18495_), .B(new_n20879_), .ZN(new_n20880_));
  NAND2_X1   g20687(.A1(new_n20880_), .A2(new_n20877_), .ZN(new_n20881_));
  OAI22_X1   g20688(.A1(new_n20878_), .A2(new_n18495_), .B1(new_n20871_), .B2(new_n20876_), .ZN(new_n20882_));
  AOI21_X1   g20689(.A1(new_n20882_), .A2(\asqrt[10] ), .B(new_n20485_), .ZN(new_n20883_));
  NOR2_X1    g20690(.A1(new_n20883_), .A2(new_n20881_), .ZN(new_n20884_));
  AOI22_X1   g20691(.A1(new_n20882_), .A2(\asqrt[10] ), .B1(new_n20880_), .B2(new_n20877_), .ZN(new_n20885_));
  INV_X1     g20692(.I(new_n20494_), .ZN(new_n20886_));
  OAI21_X1   g20693(.A1(new_n20885_), .A2(new_n17271_), .B(new_n20886_), .ZN(new_n20887_));
  NAND2_X1   g20694(.A1(new_n20887_), .A2(new_n20884_), .ZN(new_n20888_));
  OAI22_X1   g20695(.A1(new_n20885_), .A2(new_n17271_), .B1(new_n20883_), .B2(new_n20881_), .ZN(new_n20889_));
  AOI21_X1   g20696(.A1(new_n20889_), .A2(\asqrt[12] ), .B(new_n20501_), .ZN(new_n20890_));
  NOR2_X1    g20697(.A1(new_n20890_), .A2(new_n20888_), .ZN(new_n20891_));
  AOI22_X1   g20698(.A1(new_n20889_), .A2(\asqrt[12] ), .B1(new_n20887_), .B2(new_n20884_), .ZN(new_n20892_));
  INV_X1     g20699(.I(new_n20509_), .ZN(new_n20893_));
  OAI21_X1   g20700(.A1(new_n20892_), .A2(new_n16060_), .B(new_n20893_), .ZN(new_n20894_));
  NAND2_X1   g20701(.A1(new_n20894_), .A2(new_n20891_), .ZN(new_n20895_));
  OAI22_X1   g20702(.A1(new_n20892_), .A2(new_n16060_), .B1(new_n20890_), .B2(new_n20888_), .ZN(new_n20896_));
  AOI21_X1   g20703(.A1(new_n20896_), .A2(\asqrt[14] ), .B(new_n20516_), .ZN(new_n20897_));
  NOR2_X1    g20704(.A1(new_n20897_), .A2(new_n20895_), .ZN(new_n20898_));
  AOI22_X1   g20705(.A1(new_n20896_), .A2(\asqrt[14] ), .B1(new_n20894_), .B2(new_n20891_), .ZN(new_n20899_));
  INV_X1     g20706(.I(new_n20524_), .ZN(new_n20900_));
  OAI21_X1   g20707(.A1(new_n20899_), .A2(new_n14871_), .B(new_n20900_), .ZN(new_n20901_));
  NAND2_X1   g20708(.A1(new_n20901_), .A2(new_n20898_), .ZN(new_n20902_));
  OAI22_X1   g20709(.A1(new_n20899_), .A2(new_n14871_), .B1(new_n20897_), .B2(new_n20895_), .ZN(new_n20903_));
  AOI21_X1   g20710(.A1(new_n20903_), .A2(\asqrt[16] ), .B(new_n20531_), .ZN(new_n20904_));
  NOR2_X1    g20711(.A1(new_n20904_), .A2(new_n20902_), .ZN(new_n20905_));
  AOI22_X1   g20712(.A1(new_n20903_), .A2(\asqrt[16] ), .B1(new_n20901_), .B2(new_n20898_), .ZN(new_n20906_));
  INV_X1     g20713(.I(new_n20539_), .ZN(new_n20907_));
  OAI21_X1   g20714(.A1(new_n20906_), .A2(new_n13760_), .B(new_n20907_), .ZN(new_n20908_));
  NAND2_X1   g20715(.A1(new_n20908_), .A2(new_n20905_), .ZN(new_n20909_));
  OAI22_X1   g20716(.A1(new_n20906_), .A2(new_n13760_), .B1(new_n20904_), .B2(new_n20902_), .ZN(new_n20910_));
  AOI21_X1   g20717(.A1(new_n20910_), .A2(\asqrt[18] ), .B(new_n20546_), .ZN(new_n20911_));
  NOR2_X1    g20718(.A1(new_n20911_), .A2(new_n20909_), .ZN(new_n20912_));
  AOI22_X1   g20719(.A1(new_n20910_), .A2(\asqrt[18] ), .B1(new_n20908_), .B2(new_n20905_), .ZN(new_n20913_));
  INV_X1     g20720(.I(new_n20554_), .ZN(new_n20914_));
  OAI21_X1   g20721(.A1(new_n20913_), .A2(new_n12657_), .B(new_n20914_), .ZN(new_n20915_));
  NAND2_X1   g20722(.A1(new_n20915_), .A2(new_n20912_), .ZN(new_n20916_));
  OAI22_X1   g20723(.A1(new_n20913_), .A2(new_n12657_), .B1(new_n20911_), .B2(new_n20909_), .ZN(new_n20917_));
  AOI21_X1   g20724(.A1(new_n20917_), .A2(\asqrt[20] ), .B(new_n20561_), .ZN(new_n20918_));
  NOR2_X1    g20725(.A1(new_n20918_), .A2(new_n20916_), .ZN(new_n20919_));
  AOI22_X1   g20726(.A1(new_n20917_), .A2(\asqrt[20] ), .B1(new_n20915_), .B2(new_n20912_), .ZN(new_n20920_));
  INV_X1     g20727(.I(new_n20569_), .ZN(new_n20921_));
  OAI21_X1   g20728(.A1(new_n20920_), .A2(new_n11631_), .B(new_n20921_), .ZN(new_n20922_));
  NAND2_X1   g20729(.A1(new_n20922_), .A2(new_n20919_), .ZN(new_n20923_));
  OAI22_X1   g20730(.A1(new_n20920_), .A2(new_n11631_), .B1(new_n20918_), .B2(new_n20916_), .ZN(new_n20924_));
  AOI21_X1   g20731(.A1(new_n20924_), .A2(\asqrt[22] ), .B(new_n20576_), .ZN(new_n20925_));
  NOR2_X1    g20732(.A1(new_n20925_), .A2(new_n20923_), .ZN(new_n20926_));
  AOI22_X1   g20733(.A1(new_n20924_), .A2(\asqrt[22] ), .B1(new_n20922_), .B2(new_n20919_), .ZN(new_n20927_));
  INV_X1     g20734(.I(new_n20584_), .ZN(new_n20928_));
  OAI21_X1   g20735(.A1(new_n20927_), .A2(new_n10614_), .B(new_n20928_), .ZN(new_n20929_));
  NAND2_X1   g20736(.A1(new_n20929_), .A2(new_n20926_), .ZN(new_n20930_));
  OAI22_X1   g20737(.A1(new_n20927_), .A2(new_n10614_), .B1(new_n20925_), .B2(new_n20923_), .ZN(new_n20931_));
  AOI21_X1   g20738(.A1(new_n20931_), .A2(\asqrt[24] ), .B(new_n20591_), .ZN(new_n20932_));
  NOR2_X1    g20739(.A1(new_n20932_), .A2(new_n20930_), .ZN(new_n20933_));
  AOI22_X1   g20740(.A1(new_n20931_), .A2(\asqrt[24] ), .B1(new_n20929_), .B2(new_n20926_), .ZN(new_n20934_));
  INV_X1     g20741(.I(new_n20599_), .ZN(new_n20935_));
  OAI21_X1   g20742(.A1(new_n20934_), .A2(new_n9672_), .B(new_n20935_), .ZN(new_n20936_));
  NAND2_X1   g20743(.A1(new_n20936_), .A2(new_n20933_), .ZN(new_n20937_));
  OAI22_X1   g20744(.A1(new_n20934_), .A2(new_n9672_), .B1(new_n20932_), .B2(new_n20930_), .ZN(new_n20938_));
  AOI21_X1   g20745(.A1(new_n20938_), .A2(\asqrt[26] ), .B(new_n20606_), .ZN(new_n20939_));
  NOR2_X1    g20746(.A1(new_n20939_), .A2(new_n20937_), .ZN(new_n20940_));
  AOI22_X1   g20747(.A1(new_n20938_), .A2(\asqrt[26] ), .B1(new_n20936_), .B2(new_n20933_), .ZN(new_n20941_));
  INV_X1     g20748(.I(new_n20614_), .ZN(new_n20942_));
  OAI21_X1   g20749(.A1(new_n20941_), .A2(new_n8763_), .B(new_n20942_), .ZN(new_n20943_));
  NAND2_X1   g20750(.A1(new_n20943_), .A2(new_n20940_), .ZN(new_n20944_));
  OAI22_X1   g20751(.A1(new_n20941_), .A2(new_n8763_), .B1(new_n20939_), .B2(new_n20937_), .ZN(new_n20945_));
  AOI21_X1   g20752(.A1(new_n20945_), .A2(\asqrt[28] ), .B(new_n20621_), .ZN(new_n20946_));
  NOR2_X1    g20753(.A1(new_n20946_), .A2(new_n20944_), .ZN(new_n20947_));
  AOI22_X1   g20754(.A1(new_n20945_), .A2(\asqrt[28] ), .B1(new_n20943_), .B2(new_n20940_), .ZN(new_n20948_));
  INV_X1     g20755(.I(new_n20629_), .ZN(new_n20949_));
  OAI21_X1   g20756(.A1(new_n20948_), .A2(new_n7931_), .B(new_n20949_), .ZN(new_n20950_));
  NAND2_X1   g20757(.A1(new_n20950_), .A2(new_n20947_), .ZN(new_n20951_));
  OAI22_X1   g20758(.A1(new_n20948_), .A2(new_n7931_), .B1(new_n20946_), .B2(new_n20944_), .ZN(new_n20952_));
  AOI21_X1   g20759(.A1(new_n20952_), .A2(\asqrt[30] ), .B(new_n20636_), .ZN(new_n20953_));
  NOR2_X1    g20760(.A1(new_n20953_), .A2(new_n20951_), .ZN(new_n20954_));
  AOI22_X1   g20761(.A1(new_n20952_), .A2(\asqrt[30] ), .B1(new_n20950_), .B2(new_n20947_), .ZN(new_n20955_));
  INV_X1     g20762(.I(new_n20644_), .ZN(new_n20956_));
  OAI21_X1   g20763(.A1(new_n20955_), .A2(new_n7110_), .B(new_n20956_), .ZN(new_n20957_));
  NAND2_X1   g20764(.A1(new_n20957_), .A2(new_n20954_), .ZN(new_n20958_));
  OAI22_X1   g20765(.A1(new_n20955_), .A2(new_n7110_), .B1(new_n20953_), .B2(new_n20951_), .ZN(new_n20959_));
  AOI21_X1   g20766(.A1(new_n20959_), .A2(\asqrt[32] ), .B(new_n20651_), .ZN(new_n20960_));
  NOR2_X1    g20767(.A1(new_n20960_), .A2(new_n20958_), .ZN(new_n20961_));
  AOI22_X1   g20768(.A1(new_n20959_), .A2(\asqrt[32] ), .B1(new_n20957_), .B2(new_n20954_), .ZN(new_n20962_));
  INV_X1     g20769(.I(new_n20659_), .ZN(new_n20963_));
  OAI21_X1   g20770(.A1(new_n20962_), .A2(new_n6365_), .B(new_n20963_), .ZN(new_n20964_));
  NAND2_X1   g20771(.A1(new_n20964_), .A2(new_n20961_), .ZN(new_n20965_));
  OAI22_X1   g20772(.A1(new_n20962_), .A2(new_n6365_), .B1(new_n20960_), .B2(new_n20958_), .ZN(new_n20966_));
  AOI21_X1   g20773(.A1(new_n20966_), .A2(\asqrt[34] ), .B(new_n20666_), .ZN(new_n20967_));
  NOR2_X1    g20774(.A1(new_n20967_), .A2(new_n20965_), .ZN(new_n20968_));
  AOI22_X1   g20775(.A1(new_n20966_), .A2(\asqrt[34] ), .B1(new_n20964_), .B2(new_n20961_), .ZN(new_n20969_));
  INV_X1     g20776(.I(new_n20674_), .ZN(new_n20970_));
  OAI21_X1   g20777(.A1(new_n20969_), .A2(new_n5626_), .B(new_n20970_), .ZN(new_n20971_));
  NAND2_X1   g20778(.A1(new_n20971_), .A2(new_n20968_), .ZN(new_n20972_));
  OAI22_X1   g20779(.A1(new_n20969_), .A2(new_n5626_), .B1(new_n20967_), .B2(new_n20965_), .ZN(new_n20973_));
  AOI21_X1   g20780(.A1(new_n20973_), .A2(\asqrt[36] ), .B(new_n20681_), .ZN(new_n20974_));
  NOR2_X1    g20781(.A1(new_n20974_), .A2(new_n20972_), .ZN(new_n20975_));
  AOI22_X1   g20782(.A1(new_n20973_), .A2(\asqrt[36] ), .B1(new_n20971_), .B2(new_n20968_), .ZN(new_n20976_));
  INV_X1     g20783(.I(new_n20689_), .ZN(new_n20977_));
  OAI21_X1   g20784(.A1(new_n20976_), .A2(new_n4973_), .B(new_n20977_), .ZN(new_n20978_));
  NAND2_X1   g20785(.A1(new_n20978_), .A2(new_n20975_), .ZN(new_n20979_));
  OAI22_X1   g20786(.A1(new_n20976_), .A2(new_n4973_), .B1(new_n20974_), .B2(new_n20972_), .ZN(new_n20980_));
  AOI21_X1   g20787(.A1(new_n20980_), .A2(\asqrt[38] ), .B(new_n20696_), .ZN(new_n20981_));
  NOR2_X1    g20788(.A1(new_n20981_), .A2(new_n20979_), .ZN(new_n20982_));
  AOI22_X1   g20789(.A1(new_n20980_), .A2(\asqrt[38] ), .B1(new_n20978_), .B2(new_n20975_), .ZN(new_n20983_));
  INV_X1     g20790(.I(new_n20704_), .ZN(new_n20984_));
  OAI21_X1   g20791(.A1(new_n20983_), .A2(new_n4330_), .B(new_n20984_), .ZN(new_n20985_));
  NAND2_X1   g20792(.A1(new_n20985_), .A2(new_n20982_), .ZN(new_n20986_));
  OAI22_X1   g20793(.A1(new_n20983_), .A2(new_n4330_), .B1(new_n20981_), .B2(new_n20979_), .ZN(new_n20987_));
  AOI21_X1   g20794(.A1(new_n20987_), .A2(\asqrt[40] ), .B(new_n20711_), .ZN(new_n20988_));
  NOR2_X1    g20795(.A1(new_n20988_), .A2(new_n20986_), .ZN(new_n20989_));
  AOI22_X1   g20796(.A1(new_n20987_), .A2(\asqrt[40] ), .B1(new_n20985_), .B2(new_n20982_), .ZN(new_n20990_));
  INV_X1     g20797(.I(new_n20719_), .ZN(new_n20991_));
  OAI21_X1   g20798(.A1(new_n20990_), .A2(new_n3760_), .B(new_n20991_), .ZN(new_n20992_));
  NAND2_X1   g20799(.A1(new_n20992_), .A2(new_n20989_), .ZN(new_n20993_));
  OAI22_X1   g20800(.A1(new_n20990_), .A2(new_n3760_), .B1(new_n20988_), .B2(new_n20986_), .ZN(new_n20994_));
  AOI21_X1   g20801(.A1(new_n20994_), .A2(\asqrt[42] ), .B(new_n20726_), .ZN(new_n20995_));
  NOR2_X1    g20802(.A1(new_n20995_), .A2(new_n20993_), .ZN(new_n20996_));
  AOI22_X1   g20803(.A1(new_n20994_), .A2(\asqrt[42] ), .B1(new_n20992_), .B2(new_n20989_), .ZN(new_n20997_));
  INV_X1     g20804(.I(new_n20734_), .ZN(new_n20998_));
  OAI21_X1   g20805(.A1(new_n20997_), .A2(new_n3208_), .B(new_n20998_), .ZN(new_n20999_));
  NAND2_X1   g20806(.A1(new_n20999_), .A2(new_n20996_), .ZN(new_n21000_));
  OAI22_X1   g20807(.A1(new_n20997_), .A2(new_n3208_), .B1(new_n20995_), .B2(new_n20993_), .ZN(new_n21001_));
  AOI21_X1   g20808(.A1(new_n21001_), .A2(\asqrt[44] ), .B(new_n20741_), .ZN(new_n21002_));
  NOR2_X1    g20809(.A1(new_n21002_), .A2(new_n21000_), .ZN(new_n21003_));
  AOI22_X1   g20810(.A1(new_n21001_), .A2(\asqrt[44] ), .B1(new_n20999_), .B2(new_n20996_), .ZN(new_n21004_));
  INV_X1     g20811(.I(new_n20749_), .ZN(new_n21005_));
  OAI21_X1   g20812(.A1(new_n21004_), .A2(new_n2728_), .B(new_n21005_), .ZN(new_n21006_));
  NAND2_X1   g20813(.A1(new_n21006_), .A2(new_n21003_), .ZN(new_n21007_));
  OAI22_X1   g20814(.A1(new_n21004_), .A2(new_n2728_), .B1(new_n21002_), .B2(new_n21000_), .ZN(new_n21008_));
  AOI21_X1   g20815(.A1(new_n21008_), .A2(\asqrt[46] ), .B(new_n20756_), .ZN(new_n21009_));
  NOR2_X1    g20816(.A1(new_n21009_), .A2(new_n21007_), .ZN(new_n21010_));
  AOI22_X1   g20817(.A1(new_n21008_), .A2(\asqrt[46] ), .B1(new_n21006_), .B2(new_n21003_), .ZN(new_n21011_));
  INV_X1     g20818(.I(new_n20764_), .ZN(new_n21012_));
  OAI21_X1   g20819(.A1(new_n21011_), .A2(new_n2253_), .B(new_n21012_), .ZN(new_n21013_));
  NAND2_X1   g20820(.A1(new_n21013_), .A2(new_n21010_), .ZN(new_n21014_));
  OAI22_X1   g20821(.A1(new_n21011_), .A2(new_n2253_), .B1(new_n21009_), .B2(new_n21007_), .ZN(new_n21015_));
  AOI21_X1   g20822(.A1(new_n21015_), .A2(\asqrt[48] ), .B(new_n20771_), .ZN(new_n21016_));
  NOR2_X1    g20823(.A1(new_n21016_), .A2(new_n21014_), .ZN(new_n21017_));
  AOI22_X1   g20824(.A1(new_n21015_), .A2(\asqrt[48] ), .B1(new_n21013_), .B2(new_n21010_), .ZN(new_n21018_));
  INV_X1     g20825(.I(new_n20779_), .ZN(new_n21019_));
  OAI21_X1   g20826(.A1(new_n21018_), .A2(new_n1854_), .B(new_n21019_), .ZN(new_n21020_));
  NAND2_X1   g20827(.A1(new_n21020_), .A2(new_n21017_), .ZN(new_n21021_));
  OAI22_X1   g20828(.A1(new_n21018_), .A2(new_n1854_), .B1(new_n21016_), .B2(new_n21014_), .ZN(new_n21022_));
  AOI21_X1   g20829(.A1(new_n21022_), .A2(\asqrt[50] ), .B(new_n20786_), .ZN(new_n21023_));
  NOR2_X1    g20830(.A1(new_n21023_), .A2(new_n21021_), .ZN(new_n21024_));
  AOI22_X1   g20831(.A1(new_n21022_), .A2(\asqrt[50] ), .B1(new_n21020_), .B2(new_n21017_), .ZN(new_n21025_));
  INV_X1     g20832(.I(new_n20794_), .ZN(new_n21026_));
  OAI21_X1   g20833(.A1(new_n21025_), .A2(new_n1436_), .B(new_n21026_), .ZN(new_n21027_));
  NAND2_X1   g20834(.A1(new_n21027_), .A2(new_n21024_), .ZN(new_n21028_));
  OAI22_X1   g20835(.A1(new_n21025_), .A2(new_n1436_), .B1(new_n21023_), .B2(new_n21021_), .ZN(new_n21029_));
  AOI21_X1   g20836(.A1(new_n21029_), .A2(\asqrt[52] ), .B(new_n20801_), .ZN(new_n21030_));
  NOR2_X1    g20837(.A1(new_n21030_), .A2(new_n21028_), .ZN(new_n21031_));
  AOI22_X1   g20838(.A1(new_n21029_), .A2(\asqrt[52] ), .B1(new_n21027_), .B2(new_n21024_), .ZN(new_n21032_));
  INV_X1     g20839(.I(new_n20809_), .ZN(new_n21033_));
  OAI21_X1   g20840(.A1(new_n21032_), .A2(new_n1096_), .B(new_n21033_), .ZN(new_n21034_));
  NAND2_X1   g20841(.A1(new_n21034_), .A2(new_n21031_), .ZN(new_n21035_));
  OAI22_X1   g20842(.A1(new_n21032_), .A2(new_n1096_), .B1(new_n21030_), .B2(new_n21028_), .ZN(new_n21036_));
  AOI21_X1   g20843(.A1(new_n21036_), .A2(\asqrt[54] ), .B(new_n20816_), .ZN(new_n21037_));
  NOR2_X1    g20844(.A1(new_n21037_), .A2(new_n21035_), .ZN(new_n21038_));
  AOI22_X1   g20845(.A1(new_n21036_), .A2(\asqrt[54] ), .B1(new_n21034_), .B2(new_n21031_), .ZN(new_n21039_));
  INV_X1     g20846(.I(new_n20824_), .ZN(new_n21040_));
  OAI21_X1   g20847(.A1(new_n21039_), .A2(new_n825_), .B(new_n21040_), .ZN(new_n21041_));
  NAND2_X1   g20848(.A1(new_n21041_), .A2(new_n21038_), .ZN(new_n21042_));
  OAI22_X1   g20849(.A1(new_n21039_), .A2(new_n825_), .B1(new_n21037_), .B2(new_n21035_), .ZN(new_n21043_));
  AOI21_X1   g20850(.A1(new_n21043_), .A2(\asqrt[56] ), .B(new_n20831_), .ZN(new_n21044_));
  NOR2_X1    g20851(.A1(new_n21044_), .A2(new_n21042_), .ZN(new_n21045_));
  AOI22_X1   g20852(.A1(new_n21043_), .A2(\asqrt[56] ), .B1(new_n21041_), .B2(new_n21038_), .ZN(new_n21046_));
  INV_X1     g20853(.I(new_n20839_), .ZN(new_n21047_));
  OAI21_X1   g20854(.A1(new_n21046_), .A2(new_n587_), .B(new_n21047_), .ZN(new_n21048_));
  NAND2_X1   g20855(.A1(new_n21048_), .A2(new_n21045_), .ZN(new_n21049_));
  OAI22_X1   g20856(.A1(new_n21046_), .A2(new_n587_), .B1(new_n21044_), .B2(new_n21042_), .ZN(new_n21050_));
  AOI21_X1   g20857(.A1(new_n21050_), .A2(\asqrt[58] ), .B(new_n20845_), .ZN(new_n21051_));
  NOR2_X1    g20858(.A1(new_n21051_), .A2(new_n21049_), .ZN(new_n21052_));
  AOI22_X1   g20859(.A1(new_n21050_), .A2(\asqrt[58] ), .B1(new_n21048_), .B2(new_n21045_), .ZN(new_n21053_));
  INV_X1     g20860(.I(new_n20852_), .ZN(new_n21054_));
  OAI21_X1   g20861(.A1(new_n21053_), .A2(new_n376_), .B(new_n21054_), .ZN(new_n21055_));
  NAND2_X1   g20862(.A1(new_n21055_), .A2(new_n21052_), .ZN(new_n21056_));
  OAI22_X1   g20863(.A1(new_n21053_), .A2(new_n376_), .B1(new_n21051_), .B2(new_n21049_), .ZN(new_n21057_));
  AOI22_X1   g20864(.A1(new_n21057_), .A2(\asqrt[60] ), .B1(new_n21055_), .B2(new_n21052_), .ZN(new_n21058_));
  AOI21_X1   g20865(.A1(new_n21057_), .A2(\asqrt[60] ), .B(new_n20859_), .ZN(new_n21059_));
  OAI22_X1   g20866(.A1(new_n21058_), .A2(new_n229_), .B1(new_n21059_), .B2(new_n21056_), .ZN(new_n21060_));
  NOR4_X1    g20867(.A1(new_n20455_), .A2(\asqrt[61] ), .A3(new_n20409_), .A4(new_n20209_), .ZN(new_n21061_));
  XOR2_X1    g20868(.A1(new_n21061_), .A2(new_n20427_), .Z(new_n21062_));
  AOI21_X1   g20869(.A1(new_n19784_), .A2(new_n20215_), .B(new_n20455_), .ZN(new_n21063_));
  XOR2_X1    g20870(.A1(new_n20430_), .A2(new_n231_), .Z(new_n21064_));
  NOR2_X1    g20871(.A1(new_n21063_), .A2(new_n21064_), .ZN(new_n21065_));
  NAND2_X1   g20872(.A1(new_n20453_), .A2(\asqrt[62] ), .ZN(new_n21066_));
  NAND2_X1   g20873(.A1(\asqrt[6] ), .A2(new_n20435_), .ZN(new_n21067_));
  XNOR2_X1   g20874(.A1(new_n21067_), .A2(new_n21066_), .ZN(new_n21068_));
  NOR2_X1    g20875(.A1(new_n21059_), .A2(new_n21056_), .ZN(new_n21069_));
  NOR2_X1    g20876(.A1(new_n21062_), .A2(new_n196_), .ZN(new_n21070_));
  INV_X1     g20877(.I(new_n21062_), .ZN(new_n21071_));
  NOR2_X1    g20878(.A1(new_n21071_), .A2(\asqrt[62] ), .ZN(new_n21072_));
  NOR3_X1    g20879(.A1(new_n21058_), .A2(new_n229_), .A3(new_n21072_), .ZN(new_n21073_));
  AOI21_X1   g20880(.A1(new_n21073_), .A2(new_n21069_), .B(new_n21070_), .ZN(new_n21074_));
  NAND3_X1   g20881(.A1(new_n20455_), .A2(new_n19784_), .A3(new_n20413_), .ZN(new_n21075_));
  AOI21_X1   g20882(.A1(new_n21075_), .A2(new_n20430_), .B(\asqrt[63] ), .ZN(new_n21076_));
  AOI21_X1   g20883(.A1(new_n21074_), .A2(new_n21076_), .B(new_n21068_), .ZN(new_n21077_));
  NOR4_X1    g20884(.A1(new_n21060_), .A2(\asqrt[62] ), .A3(new_n21062_), .A4(new_n21068_), .ZN(new_n21078_));
  NOR3_X1    g20885(.A1(new_n21077_), .A2(new_n21065_), .A3(new_n21078_), .ZN(new_n21079_));
  NOR4_X1    g20886(.A1(new_n21079_), .A2(\asqrt[62] ), .A3(new_n21060_), .A4(new_n21062_), .ZN(new_n21080_));
  XNOR2_X1   g20887(.A1(new_n21080_), .A2(new_n20863_), .ZN(new_n21081_));
  NAND2_X1   g20888(.A1(new_n20820_), .A2(\asqrt[55] ), .ZN(new_n21082_));
  AOI21_X1   g20889(.A1(new_n21082_), .A2(new_n20819_), .B(new_n724_), .ZN(new_n21083_));
  OAI21_X1   g20890(.A1(new_n20826_), .A2(new_n21083_), .B(\asqrt[57] ), .ZN(new_n21084_));
  AOI21_X1   g20891(.A1(new_n20834_), .A2(new_n21084_), .B(new_n504_), .ZN(new_n21085_));
  OAI21_X1   g20892(.A1(new_n20841_), .A2(new_n21085_), .B(\asqrt[59] ), .ZN(new_n21086_));
  AOI21_X1   g20893(.A1(new_n20848_), .A2(new_n21086_), .B(new_n275_), .ZN(new_n21087_));
  OAI21_X1   g20894(.A1(new_n20854_), .A2(new_n21087_), .B(\asqrt[61] ), .ZN(new_n21088_));
  NOR4_X1    g20895(.A1(new_n21079_), .A2(\asqrt[61] ), .A3(new_n20856_), .A4(new_n20858_), .ZN(new_n21089_));
  XOR2_X1    g20896(.A1(new_n21089_), .A2(new_n21088_), .Z(new_n21090_));
  NOR2_X1    g20897(.A1(new_n21090_), .A2(new_n196_), .ZN(new_n21091_));
  INV_X1     g20898(.I(\a[11] ), .ZN(new_n21092_));
  NOR2_X1    g20899(.A1(\a[8] ), .A2(\a[9] ), .ZN(new_n21093_));
  INV_X1     g20900(.I(new_n21093_), .ZN(new_n21094_));
  NOR2_X1    g20901(.A1(new_n21094_), .A2(\a[10] ), .ZN(new_n21095_));
  NOR4_X1    g20902(.A1(new_n20436_), .A2(new_n19772_), .A3(new_n20432_), .A4(new_n21095_), .ZN(new_n21096_));
  XOR2_X1    g20903(.A1(new_n21096_), .A2(new_n21092_), .Z(new_n21097_));
  INV_X1     g20904(.I(new_n21097_), .ZN(new_n21098_));
  NAND2_X1   g20905(.A1(new_n20861_), .A2(new_n20854_), .ZN(new_n21099_));
  NOR3_X1    g20906(.A1(new_n21099_), .A2(new_n21088_), .A3(new_n21072_), .ZN(new_n21100_));
  INV_X1     g20907(.I(new_n21076_), .ZN(new_n21101_));
  NOR3_X1    g20908(.A1(new_n21100_), .A2(new_n21070_), .A3(new_n21101_), .ZN(new_n21102_));
  INV_X1     g20909(.I(new_n21068_), .ZN(new_n21103_));
  NAND4_X1   g20910(.A1(new_n20862_), .A2(new_n196_), .A3(new_n21071_), .A4(new_n21103_), .ZN(new_n21104_));
  OAI21_X1   g20911(.A1(new_n21102_), .A2(new_n21068_), .B(new_n21104_), .ZN(new_n21105_));
  OAI21_X1   g20912(.A1(new_n21105_), .A2(new_n21065_), .B(\a[11] ), .ZN(new_n21106_));
  NOR2_X1    g20913(.A1(new_n21097_), .A2(\a[10] ), .ZN(new_n21107_));
  INV_X1     g20914(.I(new_n21107_), .ZN(new_n21108_));
  AOI21_X1   g20915(.A1(new_n21106_), .A2(new_n21108_), .B(new_n21098_), .ZN(new_n21109_));
  INV_X1     g20916(.I(\a[10] ), .ZN(new_n21110_));
  INV_X1     g20917(.I(new_n21065_), .ZN(new_n21111_));
  INV_X1     g20918(.I(new_n21070_), .ZN(new_n21112_));
  NAND2_X1   g20919(.A1(new_n21043_), .A2(\asqrt[56] ), .ZN(new_n21113_));
  AOI21_X1   g20920(.A1(new_n21113_), .A2(new_n21042_), .B(new_n587_), .ZN(new_n21114_));
  OAI21_X1   g20921(.A1(new_n21045_), .A2(new_n21114_), .B(\asqrt[58] ), .ZN(new_n21115_));
  AOI21_X1   g20922(.A1(new_n21049_), .A2(new_n21115_), .B(new_n376_), .ZN(new_n21116_));
  OAI21_X1   g20923(.A1(new_n21052_), .A2(new_n21116_), .B(\asqrt[60] ), .ZN(new_n21117_));
  AOI21_X1   g20924(.A1(new_n21056_), .A2(new_n21117_), .B(new_n229_), .ZN(new_n21118_));
  INV_X1     g20925(.I(new_n21072_), .ZN(new_n21119_));
  NAND3_X1   g20926(.A1(new_n21069_), .A2(new_n21118_), .A3(new_n21119_), .ZN(new_n21120_));
  NAND3_X1   g20927(.A1(new_n21120_), .A2(new_n21112_), .A3(new_n21076_), .ZN(new_n21121_));
  AOI21_X1   g20928(.A1(new_n21121_), .A2(new_n21103_), .B(new_n21078_), .ZN(new_n21122_));
  AOI21_X1   g20929(.A1(new_n21122_), .A2(new_n21111_), .B(new_n21092_), .ZN(new_n21123_));
  NOR3_X1    g20930(.A1(new_n21123_), .A2(new_n21110_), .A3(new_n21097_), .ZN(new_n21124_));
  NAND3_X1   g20931(.A1(new_n20856_), .A2(\asqrt[61] ), .A3(new_n21119_), .ZN(new_n21125_));
  OAI21_X1   g20932(.A1(new_n21125_), .A2(new_n21099_), .B(new_n21112_), .ZN(new_n21126_));
  OAI21_X1   g20933(.A1(new_n21126_), .A2(new_n21101_), .B(new_n21103_), .ZN(new_n21127_));
  NAND3_X1   g20934(.A1(new_n21127_), .A2(new_n21111_), .A3(new_n21104_), .ZN(\asqrt[5] ));
  NAND3_X1   g20935(.A1(\asqrt[5] ), .A2(\a[10] ), .A3(\asqrt[6] ), .ZN(new_n21129_));
  NAND3_X1   g20936(.A1(new_n21079_), .A2(new_n21110_), .A3(\asqrt[6] ), .ZN(new_n21130_));
  AOI21_X1   g20937(.A1(new_n21129_), .A2(new_n21130_), .B(new_n21094_), .ZN(new_n21131_));
  NOR2_X1    g20938(.A1(new_n21111_), .A2(new_n20455_), .ZN(new_n21132_));
  NAND2_X1   g20939(.A1(new_n21078_), .A2(new_n21132_), .ZN(new_n21133_));
  OAI21_X1   g20940(.A1(new_n21133_), .A2(new_n21127_), .B(new_n19750_), .ZN(new_n21134_));
  NAND3_X1   g20941(.A1(new_n21134_), .A2(new_n21079_), .A3(new_n19758_), .ZN(new_n21135_));
  INV_X1     g20942(.I(new_n21132_), .ZN(new_n21136_));
  NOR2_X1    g20943(.A1(new_n21104_), .A2(new_n21136_), .ZN(new_n21137_));
  AOI21_X1   g20944(.A1(new_n21137_), .A2(new_n21077_), .B(\a[12] ), .ZN(new_n21138_));
  OAI21_X1   g20945(.A1(new_n21138_), .A2(new_n19759_), .B(\asqrt[5] ), .ZN(new_n21139_));
  NAND3_X1   g20946(.A1(new_n21139_), .A2(new_n21135_), .A3(new_n19782_), .ZN(new_n21140_));
  OAI22_X1   g20947(.A1(new_n21140_), .A2(new_n21131_), .B1(new_n21109_), .B2(new_n21124_), .ZN(new_n21141_));
  OAI21_X1   g20948(.A1(new_n21123_), .A2(new_n21107_), .B(new_n21097_), .ZN(new_n21142_));
  NAND3_X1   g20949(.A1(new_n21106_), .A2(\a[10] ), .A3(new_n21098_), .ZN(new_n21143_));
  NAND2_X1   g20950(.A1(new_n21143_), .A2(new_n21142_), .ZN(new_n21144_));
  OAI21_X1   g20951(.A1(new_n21144_), .A2(new_n21131_), .B(\asqrt[7] ), .ZN(new_n21145_));
  AOI21_X1   g20952(.A1(\asqrt[6] ), .A2(new_n19750_), .B(\a[13] ), .ZN(new_n21146_));
  NOR2_X1    g20953(.A1(new_n20419_), .A2(\a[12] ), .ZN(new_n21147_));
  AOI21_X1   g20954(.A1(\asqrt[6] ), .A2(\a[12] ), .B(new_n19761_), .ZN(new_n21148_));
  OAI21_X1   g20955(.A1(new_n21147_), .A2(new_n21146_), .B(new_n21148_), .ZN(new_n21149_));
  NOR3_X1    g20956(.A1(new_n21079_), .A2(new_n20444_), .A3(new_n21149_), .ZN(new_n21150_));
  INV_X1     g20957(.I(new_n21150_), .ZN(new_n21151_));
  OAI21_X1   g20958(.A1(new_n21079_), .A2(new_n21149_), .B(new_n20444_), .ZN(new_n21152_));
  NAND3_X1   g20959(.A1(new_n21151_), .A2(new_n19100_), .A3(new_n21152_), .ZN(new_n21153_));
  INV_X1     g20960(.I(new_n21153_), .ZN(new_n21154_));
  AOI21_X1   g20961(.A1(new_n21145_), .A2(new_n21154_), .B(new_n21141_), .ZN(new_n21155_));
  AOI21_X1   g20962(.A1(new_n21145_), .A2(new_n21141_), .B(new_n19100_), .ZN(new_n21156_));
  NOR2_X1    g20963(.A1(new_n20458_), .A2(new_n20451_), .ZN(new_n21157_));
  NOR4_X1    g20964(.A1(new_n21079_), .A2(\asqrt[8] ), .A3(new_n21157_), .A4(new_n20872_), .ZN(new_n21158_));
  NAND2_X1   g20965(.A1(new_n20872_), .A2(\asqrt[8] ), .ZN(new_n21159_));
  NOR4_X1    g20966(.A1(new_n21079_), .A2(\asqrt[8] ), .A3(new_n21157_), .A4(new_n20872_), .ZN(new_n21160_));
  NOR2_X1    g20967(.A1(new_n21160_), .A2(new_n21159_), .ZN(new_n21161_));
  NOR3_X1    g20968(.A1(new_n21161_), .A2(\asqrt[9] ), .A3(new_n21158_), .ZN(new_n21162_));
  INV_X1     g20969(.I(new_n21162_), .ZN(new_n21163_));
  OAI21_X1   g20970(.A1(new_n21156_), .A2(new_n21163_), .B(new_n21155_), .ZN(new_n21164_));
  OAI21_X1   g20971(.A1(new_n21155_), .A2(new_n21156_), .B(\asqrt[9] ), .ZN(new_n21165_));
  NOR2_X1    g20972(.A1(new_n20466_), .A2(new_n20468_), .ZN(new_n21166_));
  NOR4_X1    g20973(.A1(new_n21079_), .A2(\asqrt[9] ), .A3(new_n21166_), .A4(new_n20472_), .ZN(new_n21167_));
  AOI21_X1   g20974(.A1(new_n20871_), .A2(new_n21159_), .B(new_n18495_), .ZN(new_n21168_));
  NOR2_X1    g20975(.A1(new_n21167_), .A2(new_n21168_), .ZN(new_n21169_));
  NAND2_X1   g20976(.A1(new_n21169_), .A2(new_n17893_), .ZN(new_n21170_));
  INV_X1     g20977(.I(new_n21170_), .ZN(new_n21171_));
  AOI21_X1   g20978(.A1(new_n21165_), .A2(new_n21171_), .B(new_n21164_), .ZN(new_n21172_));
  NOR3_X1    g20979(.A1(new_n21079_), .A2(new_n21110_), .A3(new_n20455_), .ZN(new_n21173_));
  NOR4_X1    g20980(.A1(new_n21105_), .A2(\a[10] ), .A3(new_n20455_), .A4(new_n21065_), .ZN(new_n21174_));
  OAI21_X1   g20981(.A1(new_n21173_), .A2(new_n21174_), .B(new_n21093_), .ZN(new_n21175_));
  NOR3_X1    g20982(.A1(new_n21138_), .A2(\asqrt[5] ), .A3(new_n19759_), .ZN(new_n21176_));
  AOI21_X1   g20983(.A1(new_n21134_), .A2(new_n19758_), .B(new_n21079_), .ZN(new_n21177_));
  NOR3_X1    g20984(.A1(new_n21176_), .A2(new_n21177_), .A3(\asqrt[7] ), .ZN(new_n21178_));
  NAND2_X1   g20985(.A1(new_n21178_), .A2(new_n21175_), .ZN(new_n21179_));
  NAND3_X1   g20986(.A1(new_n21175_), .A2(new_n21142_), .A3(new_n21143_), .ZN(new_n21180_));
  AOI22_X1   g20987(.A1(new_n21179_), .A2(new_n21144_), .B1(new_n21180_), .B2(\asqrt[7] ), .ZN(new_n21181_));
  OAI21_X1   g20988(.A1(new_n21181_), .A2(new_n19100_), .B(new_n21162_), .ZN(new_n21182_));
  AOI21_X1   g20989(.A1(new_n21180_), .A2(\asqrt[7] ), .B(new_n21153_), .ZN(new_n21183_));
  OAI22_X1   g20990(.A1(new_n21181_), .A2(new_n19100_), .B1(new_n21141_), .B2(new_n21183_), .ZN(new_n21184_));
  AOI22_X1   g20991(.A1(new_n21184_), .A2(\asqrt[9] ), .B1(new_n21182_), .B2(new_n21155_), .ZN(new_n21185_));
  NAND2_X1   g20992(.A1(new_n20882_), .A2(\asqrt[10] ), .ZN(new_n21186_));
  NOR4_X1    g20993(.A1(new_n21079_), .A2(\asqrt[10] ), .A3(new_n20476_), .A4(new_n20882_), .ZN(new_n21187_));
  XOR2_X1    g20994(.A1(new_n21187_), .A2(new_n21186_), .Z(new_n21188_));
  NAND2_X1   g20995(.A1(new_n21188_), .A2(new_n17271_), .ZN(new_n21189_));
  INV_X1     g20996(.I(new_n21189_), .ZN(new_n21190_));
  OAI21_X1   g20997(.A1(new_n21185_), .A2(new_n17893_), .B(new_n21190_), .ZN(new_n21191_));
  NAND2_X1   g20998(.A1(new_n21191_), .A2(new_n21172_), .ZN(new_n21192_));
  AOI21_X1   g20999(.A1(new_n21184_), .A2(\asqrt[9] ), .B(new_n21170_), .ZN(new_n21193_));
  OAI22_X1   g21000(.A1(new_n21185_), .A2(new_n17893_), .B1(new_n21193_), .B2(new_n21164_), .ZN(new_n21194_));
  NAND2_X1   g21001(.A1(new_n20489_), .A2(\asqrt[11] ), .ZN(new_n21195_));
  NOR4_X1    g21002(.A1(new_n21079_), .A2(\asqrt[11] ), .A3(new_n20484_), .A4(new_n20489_), .ZN(new_n21196_));
  XOR2_X1    g21003(.A1(new_n21196_), .A2(new_n21195_), .Z(new_n21197_));
  NAND2_X1   g21004(.A1(new_n21197_), .A2(new_n16619_), .ZN(new_n21198_));
  AOI21_X1   g21005(.A1(new_n21194_), .A2(\asqrt[11] ), .B(new_n21198_), .ZN(new_n21199_));
  NOR2_X1    g21006(.A1(new_n21199_), .A2(new_n21192_), .ZN(new_n21200_));
  AOI22_X1   g21007(.A1(new_n21194_), .A2(\asqrt[11] ), .B1(new_n21191_), .B2(new_n21172_), .ZN(new_n21201_));
  NOR4_X1    g21008(.A1(new_n21079_), .A2(\asqrt[12] ), .A3(new_n20493_), .A4(new_n20889_), .ZN(new_n21202_));
  AOI21_X1   g21009(.A1(new_n21195_), .A2(new_n20488_), .B(new_n16619_), .ZN(new_n21203_));
  NOR2_X1    g21010(.A1(new_n21202_), .A2(new_n21203_), .ZN(new_n21204_));
  NAND2_X1   g21011(.A1(new_n21204_), .A2(new_n16060_), .ZN(new_n21205_));
  INV_X1     g21012(.I(new_n21205_), .ZN(new_n21206_));
  OAI21_X1   g21013(.A1(new_n21201_), .A2(new_n16619_), .B(new_n21206_), .ZN(new_n21207_));
  NAND2_X1   g21014(.A1(new_n21207_), .A2(new_n21200_), .ZN(new_n21208_));
  OAI22_X1   g21015(.A1(new_n21201_), .A2(new_n16619_), .B1(new_n21199_), .B2(new_n21192_), .ZN(new_n21209_));
  NAND2_X1   g21016(.A1(new_n20505_), .A2(\asqrt[13] ), .ZN(new_n21210_));
  NOR4_X1    g21017(.A1(new_n21079_), .A2(\asqrt[13] ), .A3(new_n20500_), .A4(new_n20505_), .ZN(new_n21211_));
  XOR2_X1    g21018(.A1(new_n21211_), .A2(new_n21210_), .Z(new_n21212_));
  NAND2_X1   g21019(.A1(new_n21212_), .A2(new_n15447_), .ZN(new_n21213_));
  AOI21_X1   g21020(.A1(new_n21209_), .A2(\asqrt[13] ), .B(new_n21213_), .ZN(new_n21214_));
  NOR2_X1    g21021(.A1(new_n21214_), .A2(new_n21208_), .ZN(new_n21215_));
  AOI22_X1   g21022(.A1(new_n21209_), .A2(\asqrt[13] ), .B1(new_n21207_), .B2(new_n21200_), .ZN(new_n21216_));
  NAND2_X1   g21023(.A1(new_n20896_), .A2(\asqrt[14] ), .ZN(new_n21217_));
  NOR4_X1    g21024(.A1(new_n21079_), .A2(\asqrt[14] ), .A3(new_n20508_), .A4(new_n20896_), .ZN(new_n21218_));
  XOR2_X1    g21025(.A1(new_n21218_), .A2(new_n21217_), .Z(new_n21219_));
  NAND2_X1   g21026(.A1(new_n21219_), .A2(new_n14871_), .ZN(new_n21220_));
  INV_X1     g21027(.I(new_n21220_), .ZN(new_n21221_));
  OAI21_X1   g21028(.A1(new_n21216_), .A2(new_n15447_), .B(new_n21221_), .ZN(new_n21222_));
  NAND2_X1   g21029(.A1(new_n21222_), .A2(new_n21215_), .ZN(new_n21223_));
  OAI22_X1   g21030(.A1(new_n21216_), .A2(new_n15447_), .B1(new_n21214_), .B2(new_n21208_), .ZN(new_n21224_));
  NOR4_X1    g21031(.A1(new_n21079_), .A2(\asqrt[15] ), .A3(new_n20515_), .A4(new_n20520_), .ZN(new_n21225_));
  AOI21_X1   g21032(.A1(new_n21217_), .A2(new_n20895_), .B(new_n14871_), .ZN(new_n21226_));
  NOR2_X1    g21033(.A1(new_n21225_), .A2(new_n21226_), .ZN(new_n21227_));
  NAND2_X1   g21034(.A1(new_n21227_), .A2(new_n14273_), .ZN(new_n21228_));
  AOI21_X1   g21035(.A1(new_n21224_), .A2(\asqrt[15] ), .B(new_n21228_), .ZN(new_n21229_));
  NOR2_X1    g21036(.A1(new_n21229_), .A2(new_n21223_), .ZN(new_n21230_));
  AOI22_X1   g21037(.A1(new_n21224_), .A2(\asqrt[15] ), .B1(new_n21222_), .B2(new_n21215_), .ZN(new_n21231_));
  NAND2_X1   g21038(.A1(new_n20903_), .A2(\asqrt[16] ), .ZN(new_n21232_));
  NOR4_X1    g21039(.A1(new_n21079_), .A2(\asqrt[16] ), .A3(new_n20523_), .A4(new_n20903_), .ZN(new_n21233_));
  XOR2_X1    g21040(.A1(new_n21233_), .A2(new_n21232_), .Z(new_n21234_));
  NAND2_X1   g21041(.A1(new_n21234_), .A2(new_n13760_), .ZN(new_n21235_));
  INV_X1     g21042(.I(new_n21235_), .ZN(new_n21236_));
  OAI21_X1   g21043(.A1(new_n21231_), .A2(new_n14273_), .B(new_n21236_), .ZN(new_n21237_));
  NAND2_X1   g21044(.A1(new_n21237_), .A2(new_n21230_), .ZN(new_n21238_));
  OAI22_X1   g21045(.A1(new_n21231_), .A2(new_n14273_), .B1(new_n21229_), .B2(new_n21223_), .ZN(new_n21239_));
  NOR4_X1    g21046(.A1(new_n21079_), .A2(\asqrt[17] ), .A3(new_n20530_), .A4(new_n20535_), .ZN(new_n21240_));
  AOI21_X1   g21047(.A1(new_n21232_), .A2(new_n20902_), .B(new_n13760_), .ZN(new_n21241_));
  NOR2_X1    g21048(.A1(new_n21240_), .A2(new_n21241_), .ZN(new_n21242_));
  NAND2_X1   g21049(.A1(new_n21242_), .A2(new_n13192_), .ZN(new_n21243_));
  AOI21_X1   g21050(.A1(new_n21239_), .A2(\asqrt[17] ), .B(new_n21243_), .ZN(new_n21244_));
  NOR2_X1    g21051(.A1(new_n21244_), .A2(new_n21238_), .ZN(new_n21245_));
  AOI22_X1   g21052(.A1(new_n21239_), .A2(\asqrt[17] ), .B1(new_n21237_), .B2(new_n21230_), .ZN(new_n21246_));
  NAND2_X1   g21053(.A1(new_n20910_), .A2(\asqrt[18] ), .ZN(new_n21247_));
  NOR4_X1    g21054(.A1(new_n21079_), .A2(\asqrt[18] ), .A3(new_n20538_), .A4(new_n20910_), .ZN(new_n21248_));
  XOR2_X1    g21055(.A1(new_n21248_), .A2(new_n21247_), .Z(new_n21249_));
  NAND2_X1   g21056(.A1(new_n21249_), .A2(new_n12657_), .ZN(new_n21250_));
  INV_X1     g21057(.I(new_n21250_), .ZN(new_n21251_));
  OAI21_X1   g21058(.A1(new_n21246_), .A2(new_n13192_), .B(new_n21251_), .ZN(new_n21252_));
  NAND2_X1   g21059(.A1(new_n21252_), .A2(new_n21245_), .ZN(new_n21253_));
  OAI22_X1   g21060(.A1(new_n21246_), .A2(new_n13192_), .B1(new_n21244_), .B2(new_n21238_), .ZN(new_n21254_));
  NOR4_X1    g21061(.A1(new_n21079_), .A2(\asqrt[19] ), .A3(new_n20545_), .A4(new_n20550_), .ZN(new_n21255_));
  AOI21_X1   g21062(.A1(new_n21247_), .A2(new_n20909_), .B(new_n12657_), .ZN(new_n21256_));
  NOR2_X1    g21063(.A1(new_n21255_), .A2(new_n21256_), .ZN(new_n21257_));
  NAND2_X1   g21064(.A1(new_n21257_), .A2(new_n12101_), .ZN(new_n21258_));
  AOI21_X1   g21065(.A1(new_n21254_), .A2(\asqrt[19] ), .B(new_n21258_), .ZN(new_n21259_));
  NOR2_X1    g21066(.A1(new_n21259_), .A2(new_n21253_), .ZN(new_n21260_));
  AOI22_X1   g21067(.A1(new_n21254_), .A2(\asqrt[19] ), .B1(new_n21252_), .B2(new_n21245_), .ZN(new_n21261_));
  NAND2_X1   g21068(.A1(new_n20917_), .A2(\asqrt[20] ), .ZN(new_n21262_));
  NOR4_X1    g21069(.A1(new_n21079_), .A2(\asqrt[20] ), .A3(new_n20553_), .A4(new_n20917_), .ZN(new_n21263_));
  XOR2_X1    g21070(.A1(new_n21263_), .A2(new_n21262_), .Z(new_n21264_));
  NAND2_X1   g21071(.A1(new_n21264_), .A2(new_n11631_), .ZN(new_n21265_));
  INV_X1     g21072(.I(new_n21265_), .ZN(new_n21266_));
  OAI21_X1   g21073(.A1(new_n21261_), .A2(new_n12101_), .B(new_n21266_), .ZN(new_n21267_));
  NAND2_X1   g21074(.A1(new_n21267_), .A2(new_n21260_), .ZN(new_n21268_));
  OAI22_X1   g21075(.A1(new_n21261_), .A2(new_n12101_), .B1(new_n21259_), .B2(new_n21253_), .ZN(new_n21269_));
  NAND2_X1   g21076(.A1(new_n20565_), .A2(\asqrt[21] ), .ZN(new_n21270_));
  NOR4_X1    g21077(.A1(new_n21079_), .A2(\asqrt[21] ), .A3(new_n20560_), .A4(new_n20565_), .ZN(new_n21271_));
  XOR2_X1    g21078(.A1(new_n21271_), .A2(new_n21270_), .Z(new_n21272_));
  NAND2_X1   g21079(.A1(new_n21272_), .A2(new_n11105_), .ZN(new_n21273_));
  AOI21_X1   g21080(.A1(new_n21269_), .A2(\asqrt[21] ), .B(new_n21273_), .ZN(new_n21274_));
  NOR2_X1    g21081(.A1(new_n21274_), .A2(new_n21268_), .ZN(new_n21275_));
  AOI22_X1   g21082(.A1(new_n21269_), .A2(\asqrt[21] ), .B1(new_n21267_), .B2(new_n21260_), .ZN(new_n21276_));
  NOR4_X1    g21083(.A1(new_n21079_), .A2(\asqrt[22] ), .A3(new_n20568_), .A4(new_n20924_), .ZN(new_n21277_));
  AOI21_X1   g21084(.A1(new_n21270_), .A2(new_n20564_), .B(new_n11105_), .ZN(new_n21278_));
  NOR2_X1    g21085(.A1(new_n21277_), .A2(new_n21278_), .ZN(new_n21279_));
  NAND2_X1   g21086(.A1(new_n21279_), .A2(new_n10614_), .ZN(new_n21280_));
  INV_X1     g21087(.I(new_n21280_), .ZN(new_n21281_));
  OAI21_X1   g21088(.A1(new_n21276_), .A2(new_n11105_), .B(new_n21281_), .ZN(new_n21282_));
  NAND2_X1   g21089(.A1(new_n21282_), .A2(new_n21275_), .ZN(new_n21283_));
  OAI22_X1   g21090(.A1(new_n21276_), .A2(new_n11105_), .B1(new_n21274_), .B2(new_n21268_), .ZN(new_n21284_));
  NAND2_X1   g21091(.A1(new_n20580_), .A2(\asqrt[23] ), .ZN(new_n21285_));
  NOR4_X1    g21092(.A1(new_n21079_), .A2(\asqrt[23] ), .A3(new_n20575_), .A4(new_n20580_), .ZN(new_n21286_));
  XOR2_X1    g21093(.A1(new_n21286_), .A2(new_n21285_), .Z(new_n21287_));
  NAND2_X1   g21094(.A1(new_n21287_), .A2(new_n10104_), .ZN(new_n21288_));
  AOI21_X1   g21095(.A1(new_n21284_), .A2(\asqrt[23] ), .B(new_n21288_), .ZN(new_n21289_));
  NOR2_X1    g21096(.A1(new_n21289_), .A2(new_n21283_), .ZN(new_n21290_));
  AOI22_X1   g21097(.A1(new_n21284_), .A2(\asqrt[23] ), .B1(new_n21282_), .B2(new_n21275_), .ZN(new_n21291_));
  NOR4_X1    g21098(.A1(new_n21079_), .A2(\asqrt[24] ), .A3(new_n20583_), .A4(new_n20931_), .ZN(new_n21292_));
  AOI21_X1   g21099(.A1(new_n21285_), .A2(new_n20579_), .B(new_n10104_), .ZN(new_n21293_));
  NOR2_X1    g21100(.A1(new_n21292_), .A2(new_n21293_), .ZN(new_n21294_));
  NAND2_X1   g21101(.A1(new_n21294_), .A2(new_n9672_), .ZN(new_n21295_));
  INV_X1     g21102(.I(new_n21295_), .ZN(new_n21296_));
  OAI21_X1   g21103(.A1(new_n21291_), .A2(new_n10104_), .B(new_n21296_), .ZN(new_n21297_));
  NAND2_X1   g21104(.A1(new_n21297_), .A2(new_n21290_), .ZN(new_n21298_));
  OAI22_X1   g21105(.A1(new_n21291_), .A2(new_n10104_), .B1(new_n21289_), .B2(new_n21283_), .ZN(new_n21299_));
  NAND2_X1   g21106(.A1(new_n20595_), .A2(\asqrt[25] ), .ZN(new_n21300_));
  NOR4_X1    g21107(.A1(new_n21079_), .A2(\asqrt[25] ), .A3(new_n20590_), .A4(new_n20595_), .ZN(new_n21301_));
  XOR2_X1    g21108(.A1(new_n21301_), .A2(new_n21300_), .Z(new_n21302_));
  NAND2_X1   g21109(.A1(new_n21302_), .A2(new_n9212_), .ZN(new_n21303_));
  AOI21_X1   g21110(.A1(new_n21299_), .A2(\asqrt[25] ), .B(new_n21303_), .ZN(new_n21304_));
  NOR2_X1    g21111(.A1(new_n21304_), .A2(new_n21298_), .ZN(new_n21305_));
  AOI22_X1   g21112(.A1(new_n21299_), .A2(\asqrt[25] ), .B1(new_n21297_), .B2(new_n21290_), .ZN(new_n21306_));
  NOR4_X1    g21113(.A1(new_n21079_), .A2(\asqrt[26] ), .A3(new_n20598_), .A4(new_n20938_), .ZN(new_n21307_));
  AOI21_X1   g21114(.A1(new_n21300_), .A2(new_n20594_), .B(new_n9212_), .ZN(new_n21308_));
  NOR2_X1    g21115(.A1(new_n21307_), .A2(new_n21308_), .ZN(new_n21309_));
  NAND2_X1   g21116(.A1(new_n21309_), .A2(new_n8763_), .ZN(new_n21310_));
  INV_X1     g21117(.I(new_n21310_), .ZN(new_n21311_));
  OAI21_X1   g21118(.A1(new_n21306_), .A2(new_n9212_), .B(new_n21311_), .ZN(new_n21312_));
  NAND2_X1   g21119(.A1(new_n21312_), .A2(new_n21305_), .ZN(new_n21313_));
  OAI22_X1   g21120(.A1(new_n21306_), .A2(new_n9212_), .B1(new_n21304_), .B2(new_n21298_), .ZN(new_n21314_));
  NAND2_X1   g21121(.A1(new_n20610_), .A2(\asqrt[27] ), .ZN(new_n21315_));
  NOR4_X1    g21122(.A1(new_n21079_), .A2(\asqrt[27] ), .A3(new_n20605_), .A4(new_n20610_), .ZN(new_n21316_));
  XOR2_X1    g21123(.A1(new_n21316_), .A2(new_n21315_), .Z(new_n21317_));
  NAND2_X1   g21124(.A1(new_n21317_), .A2(new_n8319_), .ZN(new_n21318_));
  AOI21_X1   g21125(.A1(new_n21314_), .A2(\asqrt[27] ), .B(new_n21318_), .ZN(new_n21319_));
  NOR2_X1    g21126(.A1(new_n21319_), .A2(new_n21313_), .ZN(new_n21320_));
  AOI22_X1   g21127(.A1(new_n21314_), .A2(\asqrt[27] ), .B1(new_n21312_), .B2(new_n21305_), .ZN(new_n21321_));
  NOR4_X1    g21128(.A1(new_n21079_), .A2(\asqrt[28] ), .A3(new_n20613_), .A4(new_n20945_), .ZN(new_n21322_));
  AOI21_X1   g21129(.A1(new_n21315_), .A2(new_n20609_), .B(new_n8319_), .ZN(new_n21323_));
  NOR2_X1    g21130(.A1(new_n21322_), .A2(new_n21323_), .ZN(new_n21324_));
  NAND2_X1   g21131(.A1(new_n21324_), .A2(new_n7931_), .ZN(new_n21325_));
  INV_X1     g21132(.I(new_n21325_), .ZN(new_n21326_));
  OAI21_X1   g21133(.A1(new_n21321_), .A2(new_n8319_), .B(new_n21326_), .ZN(new_n21327_));
  NAND2_X1   g21134(.A1(new_n21327_), .A2(new_n21320_), .ZN(new_n21328_));
  OAI22_X1   g21135(.A1(new_n21321_), .A2(new_n8319_), .B1(new_n21319_), .B2(new_n21313_), .ZN(new_n21329_));
  NAND2_X1   g21136(.A1(new_n20625_), .A2(\asqrt[29] ), .ZN(new_n21330_));
  NOR4_X1    g21137(.A1(new_n21079_), .A2(\asqrt[29] ), .A3(new_n20620_), .A4(new_n20625_), .ZN(new_n21331_));
  XOR2_X1    g21138(.A1(new_n21331_), .A2(new_n21330_), .Z(new_n21332_));
  NAND2_X1   g21139(.A1(new_n21332_), .A2(new_n7517_), .ZN(new_n21333_));
  AOI21_X1   g21140(.A1(new_n21329_), .A2(\asqrt[29] ), .B(new_n21333_), .ZN(new_n21334_));
  NOR2_X1    g21141(.A1(new_n21334_), .A2(new_n21328_), .ZN(new_n21335_));
  AOI22_X1   g21142(.A1(new_n21329_), .A2(\asqrt[29] ), .B1(new_n21327_), .B2(new_n21320_), .ZN(new_n21336_));
  NOR4_X1    g21143(.A1(new_n21079_), .A2(\asqrt[30] ), .A3(new_n20628_), .A4(new_n20952_), .ZN(new_n21337_));
  AOI21_X1   g21144(.A1(new_n21330_), .A2(new_n20624_), .B(new_n7517_), .ZN(new_n21338_));
  NOR2_X1    g21145(.A1(new_n21337_), .A2(new_n21338_), .ZN(new_n21339_));
  NAND2_X1   g21146(.A1(new_n21339_), .A2(new_n7110_), .ZN(new_n21340_));
  INV_X1     g21147(.I(new_n21340_), .ZN(new_n21341_));
  OAI21_X1   g21148(.A1(new_n21336_), .A2(new_n7517_), .B(new_n21341_), .ZN(new_n21342_));
  NAND2_X1   g21149(.A1(new_n21342_), .A2(new_n21335_), .ZN(new_n21343_));
  OAI22_X1   g21150(.A1(new_n21336_), .A2(new_n7517_), .B1(new_n21334_), .B2(new_n21328_), .ZN(new_n21344_));
  NAND2_X1   g21151(.A1(new_n20640_), .A2(\asqrt[31] ), .ZN(new_n21345_));
  NOR4_X1    g21152(.A1(new_n21079_), .A2(\asqrt[31] ), .A3(new_n20635_), .A4(new_n20640_), .ZN(new_n21346_));
  XOR2_X1    g21153(.A1(new_n21346_), .A2(new_n21345_), .Z(new_n21347_));
  NAND2_X1   g21154(.A1(new_n21347_), .A2(new_n6708_), .ZN(new_n21348_));
  AOI21_X1   g21155(.A1(new_n21344_), .A2(\asqrt[31] ), .B(new_n21348_), .ZN(new_n21349_));
  NOR2_X1    g21156(.A1(new_n21349_), .A2(new_n21343_), .ZN(new_n21350_));
  AOI22_X1   g21157(.A1(new_n21344_), .A2(\asqrt[31] ), .B1(new_n21342_), .B2(new_n21335_), .ZN(new_n21351_));
  NOR4_X1    g21158(.A1(new_n21079_), .A2(\asqrt[32] ), .A3(new_n20643_), .A4(new_n20959_), .ZN(new_n21352_));
  AOI21_X1   g21159(.A1(new_n21345_), .A2(new_n20639_), .B(new_n6708_), .ZN(new_n21353_));
  NOR2_X1    g21160(.A1(new_n21352_), .A2(new_n21353_), .ZN(new_n21354_));
  NAND2_X1   g21161(.A1(new_n21354_), .A2(new_n6365_), .ZN(new_n21355_));
  INV_X1     g21162(.I(new_n21355_), .ZN(new_n21356_));
  OAI21_X1   g21163(.A1(new_n21351_), .A2(new_n6708_), .B(new_n21356_), .ZN(new_n21357_));
  NAND2_X1   g21164(.A1(new_n21357_), .A2(new_n21350_), .ZN(new_n21358_));
  OAI22_X1   g21165(.A1(new_n21351_), .A2(new_n6708_), .B1(new_n21349_), .B2(new_n21343_), .ZN(new_n21359_));
  NAND2_X1   g21166(.A1(new_n20655_), .A2(\asqrt[33] ), .ZN(new_n21360_));
  NOR4_X1    g21167(.A1(new_n21079_), .A2(\asqrt[33] ), .A3(new_n20650_), .A4(new_n20655_), .ZN(new_n21361_));
  XOR2_X1    g21168(.A1(new_n21361_), .A2(new_n21360_), .Z(new_n21362_));
  NAND2_X1   g21169(.A1(new_n21362_), .A2(new_n5991_), .ZN(new_n21363_));
  AOI21_X1   g21170(.A1(new_n21359_), .A2(\asqrt[33] ), .B(new_n21363_), .ZN(new_n21364_));
  NOR2_X1    g21171(.A1(new_n21364_), .A2(new_n21358_), .ZN(new_n21365_));
  AOI22_X1   g21172(.A1(new_n21359_), .A2(\asqrt[33] ), .B1(new_n21357_), .B2(new_n21350_), .ZN(new_n21366_));
  NOR4_X1    g21173(.A1(new_n21079_), .A2(\asqrt[34] ), .A3(new_n20658_), .A4(new_n20966_), .ZN(new_n21367_));
  AOI21_X1   g21174(.A1(new_n21360_), .A2(new_n20654_), .B(new_n5991_), .ZN(new_n21368_));
  NOR2_X1    g21175(.A1(new_n21367_), .A2(new_n21368_), .ZN(new_n21369_));
  NAND2_X1   g21176(.A1(new_n21369_), .A2(new_n5626_), .ZN(new_n21370_));
  INV_X1     g21177(.I(new_n21370_), .ZN(new_n21371_));
  OAI21_X1   g21178(.A1(new_n21366_), .A2(new_n5991_), .B(new_n21371_), .ZN(new_n21372_));
  NAND2_X1   g21179(.A1(new_n21372_), .A2(new_n21365_), .ZN(new_n21373_));
  OAI22_X1   g21180(.A1(new_n21366_), .A2(new_n5991_), .B1(new_n21364_), .B2(new_n21358_), .ZN(new_n21374_));
  NAND2_X1   g21181(.A1(new_n20670_), .A2(\asqrt[35] ), .ZN(new_n21375_));
  NOR4_X1    g21182(.A1(new_n21079_), .A2(\asqrt[35] ), .A3(new_n20665_), .A4(new_n20670_), .ZN(new_n21376_));
  XOR2_X1    g21183(.A1(new_n21376_), .A2(new_n21375_), .Z(new_n21377_));
  NAND2_X1   g21184(.A1(new_n21377_), .A2(new_n5273_), .ZN(new_n21378_));
  AOI21_X1   g21185(.A1(new_n21374_), .A2(\asqrt[35] ), .B(new_n21378_), .ZN(new_n21379_));
  NOR2_X1    g21186(.A1(new_n21379_), .A2(new_n21373_), .ZN(new_n21380_));
  AOI22_X1   g21187(.A1(new_n21374_), .A2(\asqrt[35] ), .B1(new_n21372_), .B2(new_n21365_), .ZN(new_n21381_));
  NOR4_X1    g21188(.A1(new_n21079_), .A2(\asqrt[36] ), .A3(new_n20673_), .A4(new_n20973_), .ZN(new_n21382_));
  AOI21_X1   g21189(.A1(new_n21375_), .A2(new_n20669_), .B(new_n5273_), .ZN(new_n21383_));
  NOR2_X1    g21190(.A1(new_n21382_), .A2(new_n21383_), .ZN(new_n21384_));
  NAND2_X1   g21191(.A1(new_n21384_), .A2(new_n4973_), .ZN(new_n21385_));
  INV_X1     g21192(.I(new_n21385_), .ZN(new_n21386_));
  OAI21_X1   g21193(.A1(new_n21381_), .A2(new_n5273_), .B(new_n21386_), .ZN(new_n21387_));
  NAND2_X1   g21194(.A1(new_n21387_), .A2(new_n21380_), .ZN(new_n21388_));
  OAI22_X1   g21195(.A1(new_n21381_), .A2(new_n5273_), .B1(new_n21379_), .B2(new_n21373_), .ZN(new_n21389_));
  NAND2_X1   g21196(.A1(new_n20685_), .A2(\asqrt[37] ), .ZN(new_n21390_));
  NOR4_X1    g21197(.A1(new_n21079_), .A2(\asqrt[37] ), .A3(new_n20680_), .A4(new_n20685_), .ZN(new_n21391_));
  XOR2_X1    g21198(.A1(new_n21391_), .A2(new_n21390_), .Z(new_n21392_));
  NAND2_X1   g21199(.A1(new_n21392_), .A2(new_n4645_), .ZN(new_n21393_));
  AOI21_X1   g21200(.A1(new_n21389_), .A2(\asqrt[37] ), .B(new_n21393_), .ZN(new_n21394_));
  NOR2_X1    g21201(.A1(new_n21394_), .A2(new_n21388_), .ZN(new_n21395_));
  AOI22_X1   g21202(.A1(new_n21389_), .A2(\asqrt[37] ), .B1(new_n21387_), .B2(new_n21380_), .ZN(new_n21396_));
  NOR4_X1    g21203(.A1(new_n21079_), .A2(\asqrt[38] ), .A3(new_n20688_), .A4(new_n20980_), .ZN(new_n21397_));
  AOI21_X1   g21204(.A1(new_n21390_), .A2(new_n20684_), .B(new_n4645_), .ZN(new_n21398_));
  NOR2_X1    g21205(.A1(new_n21397_), .A2(new_n21398_), .ZN(new_n21399_));
  NAND2_X1   g21206(.A1(new_n21399_), .A2(new_n4330_), .ZN(new_n21400_));
  INV_X1     g21207(.I(new_n21400_), .ZN(new_n21401_));
  OAI21_X1   g21208(.A1(new_n21396_), .A2(new_n4645_), .B(new_n21401_), .ZN(new_n21402_));
  NAND2_X1   g21209(.A1(new_n21402_), .A2(new_n21395_), .ZN(new_n21403_));
  OAI22_X1   g21210(.A1(new_n21396_), .A2(new_n4645_), .B1(new_n21394_), .B2(new_n21388_), .ZN(new_n21404_));
  NAND2_X1   g21211(.A1(new_n20700_), .A2(\asqrt[39] ), .ZN(new_n21405_));
  NOR4_X1    g21212(.A1(new_n21079_), .A2(\asqrt[39] ), .A3(new_n20695_), .A4(new_n20700_), .ZN(new_n21406_));
  XOR2_X1    g21213(.A1(new_n21406_), .A2(new_n21405_), .Z(new_n21407_));
  NAND2_X1   g21214(.A1(new_n21407_), .A2(new_n4018_), .ZN(new_n21408_));
  AOI21_X1   g21215(.A1(new_n21404_), .A2(\asqrt[39] ), .B(new_n21408_), .ZN(new_n21409_));
  NOR2_X1    g21216(.A1(new_n21409_), .A2(new_n21403_), .ZN(new_n21410_));
  AOI22_X1   g21217(.A1(new_n21404_), .A2(\asqrt[39] ), .B1(new_n21402_), .B2(new_n21395_), .ZN(new_n21411_));
  NOR4_X1    g21218(.A1(new_n21079_), .A2(\asqrt[40] ), .A3(new_n20703_), .A4(new_n20987_), .ZN(new_n21412_));
  AOI21_X1   g21219(.A1(new_n21405_), .A2(new_n20699_), .B(new_n4018_), .ZN(new_n21413_));
  NOR2_X1    g21220(.A1(new_n21412_), .A2(new_n21413_), .ZN(new_n21414_));
  NAND2_X1   g21221(.A1(new_n21414_), .A2(new_n3760_), .ZN(new_n21415_));
  INV_X1     g21222(.I(new_n21415_), .ZN(new_n21416_));
  OAI21_X1   g21223(.A1(new_n21411_), .A2(new_n4018_), .B(new_n21416_), .ZN(new_n21417_));
  NAND2_X1   g21224(.A1(new_n21417_), .A2(new_n21410_), .ZN(new_n21418_));
  OAI22_X1   g21225(.A1(new_n21411_), .A2(new_n4018_), .B1(new_n21409_), .B2(new_n21403_), .ZN(new_n21419_));
  NAND2_X1   g21226(.A1(new_n20715_), .A2(\asqrt[41] ), .ZN(new_n21420_));
  NOR4_X1    g21227(.A1(new_n21079_), .A2(\asqrt[41] ), .A3(new_n20710_), .A4(new_n20715_), .ZN(new_n21421_));
  XOR2_X1    g21228(.A1(new_n21421_), .A2(new_n21420_), .Z(new_n21422_));
  NAND2_X1   g21229(.A1(new_n21422_), .A2(new_n3481_), .ZN(new_n21423_));
  AOI21_X1   g21230(.A1(new_n21419_), .A2(\asqrt[41] ), .B(new_n21423_), .ZN(new_n21424_));
  NOR2_X1    g21231(.A1(new_n21424_), .A2(new_n21418_), .ZN(new_n21425_));
  AOI22_X1   g21232(.A1(new_n21419_), .A2(\asqrt[41] ), .B1(new_n21417_), .B2(new_n21410_), .ZN(new_n21426_));
  NOR4_X1    g21233(.A1(new_n21079_), .A2(\asqrt[42] ), .A3(new_n20718_), .A4(new_n20994_), .ZN(new_n21427_));
  AOI21_X1   g21234(.A1(new_n21420_), .A2(new_n20714_), .B(new_n3481_), .ZN(new_n21428_));
  NOR2_X1    g21235(.A1(new_n21427_), .A2(new_n21428_), .ZN(new_n21429_));
  NAND2_X1   g21236(.A1(new_n21429_), .A2(new_n3208_), .ZN(new_n21430_));
  INV_X1     g21237(.I(new_n21430_), .ZN(new_n21431_));
  OAI21_X1   g21238(.A1(new_n21426_), .A2(new_n3481_), .B(new_n21431_), .ZN(new_n21432_));
  NAND2_X1   g21239(.A1(new_n21432_), .A2(new_n21425_), .ZN(new_n21433_));
  OAI22_X1   g21240(.A1(new_n21426_), .A2(new_n3481_), .B1(new_n21424_), .B2(new_n21418_), .ZN(new_n21434_));
  NAND2_X1   g21241(.A1(new_n20730_), .A2(\asqrt[43] ), .ZN(new_n21435_));
  NOR4_X1    g21242(.A1(new_n21079_), .A2(\asqrt[43] ), .A3(new_n20725_), .A4(new_n20730_), .ZN(new_n21436_));
  XOR2_X1    g21243(.A1(new_n21436_), .A2(new_n21435_), .Z(new_n21437_));
  NAND2_X1   g21244(.A1(new_n21437_), .A2(new_n2941_), .ZN(new_n21438_));
  AOI21_X1   g21245(.A1(new_n21434_), .A2(\asqrt[43] ), .B(new_n21438_), .ZN(new_n21439_));
  NOR2_X1    g21246(.A1(new_n21439_), .A2(new_n21433_), .ZN(new_n21440_));
  AOI22_X1   g21247(.A1(new_n21434_), .A2(\asqrt[43] ), .B1(new_n21432_), .B2(new_n21425_), .ZN(new_n21441_));
  NOR4_X1    g21248(.A1(new_n21079_), .A2(\asqrt[44] ), .A3(new_n20733_), .A4(new_n21001_), .ZN(new_n21442_));
  AOI21_X1   g21249(.A1(new_n21435_), .A2(new_n20729_), .B(new_n2941_), .ZN(new_n21443_));
  NOR2_X1    g21250(.A1(new_n21442_), .A2(new_n21443_), .ZN(new_n21444_));
  NAND2_X1   g21251(.A1(new_n21444_), .A2(new_n2728_), .ZN(new_n21445_));
  INV_X1     g21252(.I(new_n21445_), .ZN(new_n21446_));
  OAI21_X1   g21253(.A1(new_n21441_), .A2(new_n2941_), .B(new_n21446_), .ZN(new_n21447_));
  NAND2_X1   g21254(.A1(new_n21447_), .A2(new_n21440_), .ZN(new_n21448_));
  OAI22_X1   g21255(.A1(new_n21441_), .A2(new_n2941_), .B1(new_n21439_), .B2(new_n21433_), .ZN(new_n21449_));
  NAND2_X1   g21256(.A1(new_n20745_), .A2(\asqrt[45] ), .ZN(new_n21450_));
  NOR4_X1    g21257(.A1(new_n21079_), .A2(\asqrt[45] ), .A3(new_n20740_), .A4(new_n20745_), .ZN(new_n21451_));
  XOR2_X1    g21258(.A1(new_n21451_), .A2(new_n21450_), .Z(new_n21452_));
  NAND2_X1   g21259(.A1(new_n21452_), .A2(new_n2488_), .ZN(new_n21453_));
  AOI21_X1   g21260(.A1(new_n21449_), .A2(\asqrt[45] ), .B(new_n21453_), .ZN(new_n21454_));
  NOR2_X1    g21261(.A1(new_n21454_), .A2(new_n21448_), .ZN(new_n21455_));
  AOI22_X1   g21262(.A1(new_n21449_), .A2(\asqrt[45] ), .B1(new_n21447_), .B2(new_n21440_), .ZN(new_n21456_));
  NOR4_X1    g21263(.A1(new_n21079_), .A2(\asqrt[46] ), .A3(new_n20748_), .A4(new_n21008_), .ZN(new_n21457_));
  AOI21_X1   g21264(.A1(new_n21450_), .A2(new_n20744_), .B(new_n2488_), .ZN(new_n21458_));
  NOR2_X1    g21265(.A1(new_n21457_), .A2(new_n21458_), .ZN(new_n21459_));
  NAND2_X1   g21266(.A1(new_n21459_), .A2(new_n2253_), .ZN(new_n21460_));
  INV_X1     g21267(.I(new_n21460_), .ZN(new_n21461_));
  OAI21_X1   g21268(.A1(new_n21456_), .A2(new_n2488_), .B(new_n21461_), .ZN(new_n21462_));
  NAND2_X1   g21269(.A1(new_n21462_), .A2(new_n21455_), .ZN(new_n21463_));
  OAI22_X1   g21270(.A1(new_n21456_), .A2(new_n2488_), .B1(new_n21454_), .B2(new_n21448_), .ZN(new_n21464_));
  NAND2_X1   g21271(.A1(new_n20760_), .A2(\asqrt[47] ), .ZN(new_n21465_));
  NOR4_X1    g21272(.A1(new_n21079_), .A2(\asqrt[47] ), .A3(new_n20755_), .A4(new_n20760_), .ZN(new_n21466_));
  XOR2_X1    g21273(.A1(new_n21466_), .A2(new_n21465_), .Z(new_n21467_));
  NAND2_X1   g21274(.A1(new_n21467_), .A2(new_n2046_), .ZN(new_n21468_));
  AOI21_X1   g21275(.A1(new_n21464_), .A2(\asqrt[47] ), .B(new_n21468_), .ZN(new_n21469_));
  NOR2_X1    g21276(.A1(new_n21469_), .A2(new_n21463_), .ZN(new_n21470_));
  AOI22_X1   g21277(.A1(new_n21464_), .A2(\asqrt[47] ), .B1(new_n21462_), .B2(new_n21455_), .ZN(new_n21471_));
  NOR4_X1    g21278(.A1(new_n21079_), .A2(\asqrt[48] ), .A3(new_n20763_), .A4(new_n21015_), .ZN(new_n21472_));
  AOI21_X1   g21279(.A1(new_n21465_), .A2(new_n20759_), .B(new_n2046_), .ZN(new_n21473_));
  NOR2_X1    g21280(.A1(new_n21472_), .A2(new_n21473_), .ZN(new_n21474_));
  NAND2_X1   g21281(.A1(new_n21474_), .A2(new_n1854_), .ZN(new_n21475_));
  INV_X1     g21282(.I(new_n21475_), .ZN(new_n21476_));
  OAI21_X1   g21283(.A1(new_n21471_), .A2(new_n2046_), .B(new_n21476_), .ZN(new_n21477_));
  NAND2_X1   g21284(.A1(new_n21477_), .A2(new_n21470_), .ZN(new_n21478_));
  OAI22_X1   g21285(.A1(new_n21471_), .A2(new_n2046_), .B1(new_n21469_), .B2(new_n21463_), .ZN(new_n21479_));
  NAND2_X1   g21286(.A1(new_n20775_), .A2(\asqrt[49] ), .ZN(new_n21480_));
  NOR4_X1    g21287(.A1(new_n21079_), .A2(\asqrt[49] ), .A3(new_n20770_), .A4(new_n20775_), .ZN(new_n21481_));
  XOR2_X1    g21288(.A1(new_n21481_), .A2(new_n21480_), .Z(new_n21482_));
  NAND2_X1   g21289(.A1(new_n21482_), .A2(new_n1595_), .ZN(new_n21483_));
  AOI21_X1   g21290(.A1(new_n21479_), .A2(\asqrt[49] ), .B(new_n21483_), .ZN(new_n21484_));
  NOR2_X1    g21291(.A1(new_n21484_), .A2(new_n21478_), .ZN(new_n21485_));
  AOI22_X1   g21292(.A1(new_n21479_), .A2(\asqrt[49] ), .B1(new_n21477_), .B2(new_n21470_), .ZN(new_n21486_));
  NOR4_X1    g21293(.A1(new_n21079_), .A2(\asqrt[50] ), .A3(new_n20778_), .A4(new_n21022_), .ZN(new_n21487_));
  AOI21_X1   g21294(.A1(new_n21480_), .A2(new_n20774_), .B(new_n1595_), .ZN(new_n21488_));
  NOR2_X1    g21295(.A1(new_n21487_), .A2(new_n21488_), .ZN(new_n21489_));
  NAND2_X1   g21296(.A1(new_n21489_), .A2(new_n1436_), .ZN(new_n21490_));
  INV_X1     g21297(.I(new_n21490_), .ZN(new_n21491_));
  OAI21_X1   g21298(.A1(new_n21486_), .A2(new_n1595_), .B(new_n21491_), .ZN(new_n21492_));
  NAND2_X1   g21299(.A1(new_n21492_), .A2(new_n21485_), .ZN(new_n21493_));
  OAI22_X1   g21300(.A1(new_n21486_), .A2(new_n1595_), .B1(new_n21484_), .B2(new_n21478_), .ZN(new_n21494_));
  NAND2_X1   g21301(.A1(new_n20790_), .A2(\asqrt[51] ), .ZN(new_n21495_));
  NOR4_X1    g21302(.A1(new_n21079_), .A2(\asqrt[51] ), .A3(new_n20785_), .A4(new_n20790_), .ZN(new_n21496_));
  XOR2_X1    g21303(.A1(new_n21496_), .A2(new_n21495_), .Z(new_n21497_));
  NAND2_X1   g21304(.A1(new_n21497_), .A2(new_n1260_), .ZN(new_n21498_));
  AOI21_X1   g21305(.A1(new_n21494_), .A2(\asqrt[51] ), .B(new_n21498_), .ZN(new_n21499_));
  NOR2_X1    g21306(.A1(new_n21499_), .A2(new_n21493_), .ZN(new_n21500_));
  AOI22_X1   g21307(.A1(new_n21494_), .A2(\asqrt[51] ), .B1(new_n21492_), .B2(new_n21485_), .ZN(new_n21501_));
  NOR4_X1    g21308(.A1(new_n21079_), .A2(\asqrt[52] ), .A3(new_n20793_), .A4(new_n21029_), .ZN(new_n21502_));
  AOI21_X1   g21309(.A1(new_n21495_), .A2(new_n20789_), .B(new_n1260_), .ZN(new_n21503_));
  NOR2_X1    g21310(.A1(new_n21502_), .A2(new_n21503_), .ZN(new_n21504_));
  NAND2_X1   g21311(.A1(new_n21504_), .A2(new_n1096_), .ZN(new_n21505_));
  INV_X1     g21312(.I(new_n21505_), .ZN(new_n21506_));
  OAI21_X1   g21313(.A1(new_n21501_), .A2(new_n1260_), .B(new_n21506_), .ZN(new_n21507_));
  NAND2_X1   g21314(.A1(new_n21507_), .A2(new_n21500_), .ZN(new_n21508_));
  OAI22_X1   g21315(.A1(new_n21501_), .A2(new_n1260_), .B1(new_n21499_), .B2(new_n21493_), .ZN(new_n21509_));
  NAND2_X1   g21316(.A1(new_n20805_), .A2(\asqrt[53] ), .ZN(new_n21510_));
  NOR4_X1    g21317(.A1(new_n21079_), .A2(\asqrt[53] ), .A3(new_n20800_), .A4(new_n20805_), .ZN(new_n21511_));
  XOR2_X1    g21318(.A1(new_n21511_), .A2(new_n21510_), .Z(new_n21512_));
  NAND2_X1   g21319(.A1(new_n21512_), .A2(new_n970_), .ZN(new_n21513_));
  AOI21_X1   g21320(.A1(new_n21509_), .A2(\asqrt[53] ), .B(new_n21513_), .ZN(new_n21514_));
  NOR2_X1    g21321(.A1(new_n21514_), .A2(new_n21508_), .ZN(new_n21515_));
  AOI22_X1   g21322(.A1(new_n21509_), .A2(\asqrt[53] ), .B1(new_n21507_), .B2(new_n21500_), .ZN(new_n21516_));
  NOR2_X1    g21323(.A1(new_n20812_), .A2(new_n970_), .ZN(new_n21517_));
  NOR4_X1    g21324(.A1(new_n21079_), .A2(\asqrt[54] ), .A3(new_n20808_), .A4(new_n21036_), .ZN(new_n21518_));
  XNOR2_X1   g21325(.A1(new_n21518_), .A2(new_n21517_), .ZN(new_n21519_));
  NAND2_X1   g21326(.A1(new_n21519_), .A2(new_n825_), .ZN(new_n21520_));
  INV_X1     g21327(.I(new_n21520_), .ZN(new_n21521_));
  OAI21_X1   g21328(.A1(new_n21516_), .A2(new_n970_), .B(new_n21521_), .ZN(new_n21522_));
  NAND2_X1   g21329(.A1(new_n21522_), .A2(new_n21515_), .ZN(new_n21523_));
  OAI22_X1   g21330(.A1(new_n21516_), .A2(new_n970_), .B1(new_n21514_), .B2(new_n21508_), .ZN(new_n21524_));
  NOR4_X1    g21331(.A1(new_n21079_), .A2(\asqrt[55] ), .A3(new_n20815_), .A4(new_n20820_), .ZN(new_n21525_));
  XOR2_X1    g21332(.A1(new_n21525_), .A2(new_n21082_), .Z(new_n21526_));
  NAND2_X1   g21333(.A1(new_n21526_), .A2(new_n724_), .ZN(new_n21527_));
  AOI21_X1   g21334(.A1(new_n21524_), .A2(\asqrt[55] ), .B(new_n21527_), .ZN(new_n21528_));
  NOR2_X1    g21335(.A1(new_n21528_), .A2(new_n21523_), .ZN(new_n21529_));
  AOI22_X1   g21336(.A1(new_n21524_), .A2(\asqrt[55] ), .B1(new_n21522_), .B2(new_n21515_), .ZN(new_n21530_));
  NOR4_X1    g21337(.A1(new_n21079_), .A2(\asqrt[56] ), .A3(new_n20823_), .A4(new_n21043_), .ZN(new_n21531_));
  XOR2_X1    g21338(.A1(new_n21531_), .A2(new_n21113_), .Z(new_n21532_));
  NAND2_X1   g21339(.A1(new_n21532_), .A2(new_n587_), .ZN(new_n21533_));
  INV_X1     g21340(.I(new_n21533_), .ZN(new_n21534_));
  OAI21_X1   g21341(.A1(new_n21530_), .A2(new_n724_), .B(new_n21534_), .ZN(new_n21535_));
  NAND2_X1   g21342(.A1(new_n21535_), .A2(new_n21529_), .ZN(new_n21536_));
  OAI22_X1   g21343(.A1(new_n21530_), .A2(new_n724_), .B1(new_n21528_), .B2(new_n21523_), .ZN(new_n21537_));
  NOR4_X1    g21344(.A1(new_n21079_), .A2(\asqrt[57] ), .A3(new_n20830_), .A4(new_n20835_), .ZN(new_n21538_));
  XOR2_X1    g21345(.A1(new_n21538_), .A2(new_n21084_), .Z(new_n21539_));
  NAND2_X1   g21346(.A1(new_n21539_), .A2(new_n504_), .ZN(new_n21540_));
  AOI21_X1   g21347(.A1(new_n21537_), .A2(\asqrt[57] ), .B(new_n21540_), .ZN(new_n21541_));
  NOR2_X1    g21348(.A1(new_n21541_), .A2(new_n21536_), .ZN(new_n21542_));
  AOI22_X1   g21349(.A1(new_n21537_), .A2(\asqrt[57] ), .B1(new_n21535_), .B2(new_n21529_), .ZN(new_n21543_));
  NOR4_X1    g21350(.A1(new_n21079_), .A2(\asqrt[58] ), .A3(new_n20838_), .A4(new_n21050_), .ZN(new_n21544_));
  XOR2_X1    g21351(.A1(new_n21544_), .A2(new_n21115_), .Z(new_n21545_));
  NAND2_X1   g21352(.A1(new_n21545_), .A2(new_n376_), .ZN(new_n21546_));
  INV_X1     g21353(.I(new_n21546_), .ZN(new_n21547_));
  OAI21_X1   g21354(.A1(new_n21543_), .A2(new_n504_), .B(new_n21547_), .ZN(new_n21548_));
  NAND2_X1   g21355(.A1(new_n21548_), .A2(new_n21542_), .ZN(new_n21549_));
  OAI22_X1   g21356(.A1(new_n21543_), .A2(new_n504_), .B1(new_n21541_), .B2(new_n21536_), .ZN(new_n21550_));
  NOR4_X1    g21357(.A1(new_n21079_), .A2(\asqrt[59] ), .A3(new_n20844_), .A4(new_n20849_), .ZN(new_n21551_));
  XOR2_X1    g21358(.A1(new_n21551_), .A2(new_n21086_), .Z(new_n21552_));
  NAND2_X1   g21359(.A1(new_n21552_), .A2(new_n275_), .ZN(new_n21553_));
  AOI21_X1   g21360(.A1(new_n21550_), .A2(\asqrt[59] ), .B(new_n21553_), .ZN(new_n21554_));
  NOR2_X1    g21361(.A1(new_n21554_), .A2(new_n21549_), .ZN(new_n21555_));
  AOI22_X1   g21362(.A1(new_n21550_), .A2(\asqrt[59] ), .B1(new_n21548_), .B2(new_n21542_), .ZN(new_n21556_));
  NOR4_X1    g21363(.A1(new_n21079_), .A2(\asqrt[60] ), .A3(new_n20851_), .A4(new_n21057_), .ZN(new_n21557_));
  XOR2_X1    g21364(.A1(new_n21557_), .A2(new_n21117_), .Z(new_n21558_));
  NAND2_X1   g21365(.A1(new_n21558_), .A2(new_n229_), .ZN(new_n21559_));
  INV_X1     g21366(.I(new_n21559_), .ZN(new_n21560_));
  OAI21_X1   g21367(.A1(new_n21556_), .A2(new_n275_), .B(new_n21560_), .ZN(new_n21561_));
  NAND2_X1   g21368(.A1(new_n21561_), .A2(new_n21555_), .ZN(new_n21562_));
  NAND2_X1   g21369(.A1(new_n21537_), .A2(\asqrt[57] ), .ZN(new_n21563_));
  AOI21_X1   g21370(.A1(new_n21563_), .A2(new_n21536_), .B(new_n504_), .ZN(new_n21564_));
  OAI21_X1   g21371(.A1(new_n21542_), .A2(new_n21564_), .B(\asqrt[59] ), .ZN(new_n21565_));
  AOI21_X1   g21372(.A1(new_n21549_), .A2(new_n21565_), .B(new_n275_), .ZN(new_n21566_));
  OAI21_X1   g21373(.A1(new_n21555_), .A2(new_n21566_), .B(\asqrt[61] ), .ZN(new_n21567_));
  INV_X1     g21374(.I(new_n21090_), .ZN(new_n21568_));
  NOR2_X1    g21375(.A1(new_n21568_), .A2(\asqrt[62] ), .ZN(new_n21569_));
  NOR3_X1    g21376(.A1(new_n21562_), .A2(new_n21567_), .A3(new_n21569_), .ZN(new_n21570_));
  NAND3_X1   g21377(.A1(new_n21079_), .A2(new_n21068_), .A3(new_n21104_), .ZN(new_n21571_));
  AOI21_X1   g21378(.A1(new_n21571_), .A2(new_n21126_), .B(\asqrt[63] ), .ZN(new_n21572_));
  INV_X1     g21379(.I(new_n21572_), .ZN(new_n21573_));
  NOR3_X1    g21380(.A1(new_n21570_), .A2(new_n21091_), .A3(new_n21573_), .ZN(new_n21574_));
  INV_X1     g21381(.I(new_n21081_), .ZN(new_n21575_));
  OAI22_X1   g21382(.A1(new_n21556_), .A2(new_n275_), .B1(new_n21554_), .B2(new_n21549_), .ZN(new_n21576_));
  AOI22_X1   g21383(.A1(new_n21576_), .A2(\asqrt[61] ), .B1(new_n21561_), .B2(new_n21555_), .ZN(new_n21577_));
  NAND4_X1   g21384(.A1(new_n21577_), .A2(new_n196_), .A3(new_n21575_), .A4(new_n21568_), .ZN(new_n21578_));
  OAI21_X1   g21385(.A1(new_n21574_), .A2(new_n21081_), .B(new_n21578_), .ZN(new_n21579_));
  AOI21_X1   g21386(.A1(new_n21068_), .A2(new_n21074_), .B(new_n21079_), .ZN(new_n21580_));
  XOR2_X1    g21387(.A1(new_n21074_), .A2(\asqrt[63] ), .Z(new_n21581_));
  NOR2_X1    g21388(.A1(new_n21580_), .A2(new_n21581_), .ZN(new_n21582_));
  INV_X1     g21389(.I(new_n21582_), .ZN(new_n21583_));
  NOR2_X1    g21390(.A1(\a[4] ), .A2(\a[5] ), .ZN(new_n21584_));
  INV_X1     g21391(.I(new_n21584_), .ZN(new_n21585_));
  OAI21_X1   g21392(.A1(\a[6] ), .A2(new_n21585_), .B(new_n21583_), .ZN(new_n21586_));
  NOR2_X1    g21393(.A1(new_n21579_), .A2(new_n21586_), .ZN(new_n21587_));
  XOR2_X1    g21394(.A1(new_n21587_), .A2(new_n217_), .Z(new_n21588_));
  INV_X1     g21395(.I(new_n21588_), .ZN(new_n21589_));
  NOR2_X1    g21396(.A1(new_n21156_), .A2(new_n21163_), .ZN(new_n21590_));
  NOR3_X1    g21397(.A1(new_n21590_), .A2(new_n21141_), .A3(new_n21183_), .ZN(new_n21591_));
  NAND2_X1   g21398(.A1(new_n21165_), .A2(new_n21171_), .ZN(new_n21592_));
  NAND2_X1   g21399(.A1(new_n21592_), .A2(new_n21591_), .ZN(new_n21593_));
  NAND2_X1   g21400(.A1(new_n21164_), .A2(new_n21165_), .ZN(new_n21594_));
  AOI21_X1   g21401(.A1(new_n21594_), .A2(\asqrt[10] ), .B(new_n21189_), .ZN(new_n21595_));
  NOR2_X1    g21402(.A1(new_n21595_), .A2(new_n21593_), .ZN(new_n21596_));
  AOI21_X1   g21403(.A1(new_n21164_), .A2(new_n21165_), .B(new_n17893_), .ZN(new_n21597_));
  OAI21_X1   g21404(.A1(new_n21172_), .A2(new_n21597_), .B(\asqrt[11] ), .ZN(new_n21598_));
  INV_X1     g21405(.I(new_n21198_), .ZN(new_n21599_));
  NAND2_X1   g21406(.A1(new_n21598_), .A2(new_n21599_), .ZN(new_n21600_));
  NAND2_X1   g21407(.A1(new_n21600_), .A2(new_n21596_), .ZN(new_n21601_));
  AOI22_X1   g21408(.A1(new_n21594_), .A2(\asqrt[10] ), .B1(new_n21592_), .B2(new_n21591_), .ZN(new_n21602_));
  OAI22_X1   g21409(.A1(new_n21602_), .A2(new_n17271_), .B1(new_n21595_), .B2(new_n21593_), .ZN(new_n21603_));
  AOI21_X1   g21410(.A1(new_n21603_), .A2(\asqrt[12] ), .B(new_n21205_), .ZN(new_n21604_));
  NOR2_X1    g21411(.A1(new_n21604_), .A2(new_n21601_), .ZN(new_n21605_));
  AOI22_X1   g21412(.A1(new_n21603_), .A2(\asqrt[12] ), .B1(new_n21600_), .B2(new_n21596_), .ZN(new_n21606_));
  INV_X1     g21413(.I(new_n21213_), .ZN(new_n21607_));
  OAI21_X1   g21414(.A1(new_n21606_), .A2(new_n16060_), .B(new_n21607_), .ZN(new_n21608_));
  NAND2_X1   g21415(.A1(new_n21608_), .A2(new_n21605_), .ZN(new_n21609_));
  OAI22_X1   g21416(.A1(new_n21606_), .A2(new_n16060_), .B1(new_n21604_), .B2(new_n21601_), .ZN(new_n21610_));
  AOI21_X1   g21417(.A1(new_n21610_), .A2(\asqrt[14] ), .B(new_n21220_), .ZN(new_n21611_));
  NOR2_X1    g21418(.A1(new_n21611_), .A2(new_n21609_), .ZN(new_n21612_));
  AOI22_X1   g21419(.A1(new_n21610_), .A2(\asqrt[14] ), .B1(new_n21608_), .B2(new_n21605_), .ZN(new_n21613_));
  INV_X1     g21420(.I(new_n21228_), .ZN(new_n21614_));
  OAI21_X1   g21421(.A1(new_n21613_), .A2(new_n14871_), .B(new_n21614_), .ZN(new_n21615_));
  NAND2_X1   g21422(.A1(new_n21615_), .A2(new_n21612_), .ZN(new_n21616_));
  OAI22_X1   g21423(.A1(new_n21613_), .A2(new_n14871_), .B1(new_n21611_), .B2(new_n21609_), .ZN(new_n21617_));
  AOI21_X1   g21424(.A1(new_n21617_), .A2(\asqrt[16] ), .B(new_n21235_), .ZN(new_n21618_));
  NOR2_X1    g21425(.A1(new_n21618_), .A2(new_n21616_), .ZN(new_n21619_));
  AOI22_X1   g21426(.A1(new_n21617_), .A2(\asqrt[16] ), .B1(new_n21615_), .B2(new_n21612_), .ZN(new_n21620_));
  INV_X1     g21427(.I(new_n21243_), .ZN(new_n21621_));
  OAI21_X1   g21428(.A1(new_n21620_), .A2(new_n13760_), .B(new_n21621_), .ZN(new_n21622_));
  NAND2_X1   g21429(.A1(new_n21622_), .A2(new_n21619_), .ZN(new_n21623_));
  OAI22_X1   g21430(.A1(new_n21620_), .A2(new_n13760_), .B1(new_n21618_), .B2(new_n21616_), .ZN(new_n21624_));
  AOI21_X1   g21431(.A1(new_n21624_), .A2(\asqrt[18] ), .B(new_n21250_), .ZN(new_n21625_));
  NOR2_X1    g21432(.A1(new_n21625_), .A2(new_n21623_), .ZN(new_n21626_));
  AOI22_X1   g21433(.A1(new_n21624_), .A2(\asqrt[18] ), .B1(new_n21622_), .B2(new_n21619_), .ZN(new_n21627_));
  INV_X1     g21434(.I(new_n21258_), .ZN(new_n21628_));
  OAI21_X1   g21435(.A1(new_n21627_), .A2(new_n12657_), .B(new_n21628_), .ZN(new_n21629_));
  NAND2_X1   g21436(.A1(new_n21629_), .A2(new_n21626_), .ZN(new_n21630_));
  OAI22_X1   g21437(.A1(new_n21627_), .A2(new_n12657_), .B1(new_n21625_), .B2(new_n21623_), .ZN(new_n21631_));
  AOI21_X1   g21438(.A1(new_n21631_), .A2(\asqrt[20] ), .B(new_n21265_), .ZN(new_n21632_));
  NOR2_X1    g21439(.A1(new_n21632_), .A2(new_n21630_), .ZN(new_n21633_));
  AOI22_X1   g21440(.A1(new_n21631_), .A2(\asqrt[20] ), .B1(new_n21629_), .B2(new_n21626_), .ZN(new_n21634_));
  INV_X1     g21441(.I(new_n21273_), .ZN(new_n21635_));
  OAI21_X1   g21442(.A1(new_n21634_), .A2(new_n11631_), .B(new_n21635_), .ZN(new_n21636_));
  NAND2_X1   g21443(.A1(new_n21636_), .A2(new_n21633_), .ZN(new_n21637_));
  OAI22_X1   g21444(.A1(new_n21634_), .A2(new_n11631_), .B1(new_n21632_), .B2(new_n21630_), .ZN(new_n21638_));
  AOI21_X1   g21445(.A1(new_n21638_), .A2(\asqrt[22] ), .B(new_n21280_), .ZN(new_n21639_));
  NOR2_X1    g21446(.A1(new_n21639_), .A2(new_n21637_), .ZN(new_n21640_));
  AOI22_X1   g21447(.A1(new_n21638_), .A2(\asqrt[22] ), .B1(new_n21636_), .B2(new_n21633_), .ZN(new_n21641_));
  INV_X1     g21448(.I(new_n21288_), .ZN(new_n21642_));
  OAI21_X1   g21449(.A1(new_n21641_), .A2(new_n10614_), .B(new_n21642_), .ZN(new_n21643_));
  NAND2_X1   g21450(.A1(new_n21643_), .A2(new_n21640_), .ZN(new_n21644_));
  OAI22_X1   g21451(.A1(new_n21641_), .A2(new_n10614_), .B1(new_n21639_), .B2(new_n21637_), .ZN(new_n21645_));
  AOI21_X1   g21452(.A1(new_n21645_), .A2(\asqrt[24] ), .B(new_n21295_), .ZN(new_n21646_));
  NOR2_X1    g21453(.A1(new_n21646_), .A2(new_n21644_), .ZN(new_n21647_));
  AOI22_X1   g21454(.A1(new_n21645_), .A2(\asqrt[24] ), .B1(new_n21643_), .B2(new_n21640_), .ZN(new_n21648_));
  INV_X1     g21455(.I(new_n21303_), .ZN(new_n21649_));
  OAI21_X1   g21456(.A1(new_n21648_), .A2(new_n9672_), .B(new_n21649_), .ZN(new_n21650_));
  NAND2_X1   g21457(.A1(new_n21650_), .A2(new_n21647_), .ZN(new_n21651_));
  OAI22_X1   g21458(.A1(new_n21648_), .A2(new_n9672_), .B1(new_n21646_), .B2(new_n21644_), .ZN(new_n21652_));
  AOI21_X1   g21459(.A1(new_n21652_), .A2(\asqrt[26] ), .B(new_n21310_), .ZN(new_n21653_));
  NOR2_X1    g21460(.A1(new_n21653_), .A2(new_n21651_), .ZN(new_n21654_));
  AOI22_X1   g21461(.A1(new_n21652_), .A2(\asqrt[26] ), .B1(new_n21650_), .B2(new_n21647_), .ZN(new_n21655_));
  INV_X1     g21462(.I(new_n21318_), .ZN(new_n21656_));
  OAI21_X1   g21463(.A1(new_n21655_), .A2(new_n8763_), .B(new_n21656_), .ZN(new_n21657_));
  NAND2_X1   g21464(.A1(new_n21657_), .A2(new_n21654_), .ZN(new_n21658_));
  OAI22_X1   g21465(.A1(new_n21655_), .A2(new_n8763_), .B1(new_n21653_), .B2(new_n21651_), .ZN(new_n21659_));
  AOI21_X1   g21466(.A1(new_n21659_), .A2(\asqrt[28] ), .B(new_n21325_), .ZN(new_n21660_));
  NOR2_X1    g21467(.A1(new_n21660_), .A2(new_n21658_), .ZN(new_n21661_));
  AOI22_X1   g21468(.A1(new_n21659_), .A2(\asqrt[28] ), .B1(new_n21657_), .B2(new_n21654_), .ZN(new_n21662_));
  INV_X1     g21469(.I(new_n21333_), .ZN(new_n21663_));
  OAI21_X1   g21470(.A1(new_n21662_), .A2(new_n7931_), .B(new_n21663_), .ZN(new_n21664_));
  NAND2_X1   g21471(.A1(new_n21664_), .A2(new_n21661_), .ZN(new_n21665_));
  OAI22_X1   g21472(.A1(new_n21662_), .A2(new_n7931_), .B1(new_n21660_), .B2(new_n21658_), .ZN(new_n21666_));
  AOI21_X1   g21473(.A1(new_n21666_), .A2(\asqrt[30] ), .B(new_n21340_), .ZN(new_n21667_));
  NOR2_X1    g21474(.A1(new_n21667_), .A2(new_n21665_), .ZN(new_n21668_));
  AOI22_X1   g21475(.A1(new_n21666_), .A2(\asqrt[30] ), .B1(new_n21664_), .B2(new_n21661_), .ZN(new_n21669_));
  INV_X1     g21476(.I(new_n21348_), .ZN(new_n21670_));
  OAI21_X1   g21477(.A1(new_n21669_), .A2(new_n7110_), .B(new_n21670_), .ZN(new_n21671_));
  NAND2_X1   g21478(.A1(new_n21671_), .A2(new_n21668_), .ZN(new_n21672_));
  OAI22_X1   g21479(.A1(new_n21669_), .A2(new_n7110_), .B1(new_n21667_), .B2(new_n21665_), .ZN(new_n21673_));
  AOI21_X1   g21480(.A1(new_n21673_), .A2(\asqrt[32] ), .B(new_n21355_), .ZN(new_n21674_));
  NOR2_X1    g21481(.A1(new_n21674_), .A2(new_n21672_), .ZN(new_n21675_));
  AOI22_X1   g21482(.A1(new_n21673_), .A2(\asqrt[32] ), .B1(new_n21671_), .B2(new_n21668_), .ZN(new_n21676_));
  INV_X1     g21483(.I(new_n21363_), .ZN(new_n21677_));
  OAI21_X1   g21484(.A1(new_n21676_), .A2(new_n6365_), .B(new_n21677_), .ZN(new_n21678_));
  NAND2_X1   g21485(.A1(new_n21678_), .A2(new_n21675_), .ZN(new_n21679_));
  OAI22_X1   g21486(.A1(new_n21676_), .A2(new_n6365_), .B1(new_n21674_), .B2(new_n21672_), .ZN(new_n21680_));
  AOI21_X1   g21487(.A1(new_n21680_), .A2(\asqrt[34] ), .B(new_n21370_), .ZN(new_n21681_));
  NOR2_X1    g21488(.A1(new_n21681_), .A2(new_n21679_), .ZN(new_n21682_));
  AOI22_X1   g21489(.A1(new_n21680_), .A2(\asqrt[34] ), .B1(new_n21678_), .B2(new_n21675_), .ZN(new_n21683_));
  INV_X1     g21490(.I(new_n21378_), .ZN(new_n21684_));
  OAI21_X1   g21491(.A1(new_n21683_), .A2(new_n5626_), .B(new_n21684_), .ZN(new_n21685_));
  NAND2_X1   g21492(.A1(new_n21685_), .A2(new_n21682_), .ZN(new_n21686_));
  OAI22_X1   g21493(.A1(new_n21683_), .A2(new_n5626_), .B1(new_n21681_), .B2(new_n21679_), .ZN(new_n21687_));
  AOI21_X1   g21494(.A1(new_n21687_), .A2(\asqrt[36] ), .B(new_n21385_), .ZN(new_n21688_));
  NOR2_X1    g21495(.A1(new_n21688_), .A2(new_n21686_), .ZN(new_n21689_));
  AOI22_X1   g21496(.A1(new_n21687_), .A2(\asqrt[36] ), .B1(new_n21685_), .B2(new_n21682_), .ZN(new_n21690_));
  INV_X1     g21497(.I(new_n21393_), .ZN(new_n21691_));
  OAI21_X1   g21498(.A1(new_n21690_), .A2(new_n4973_), .B(new_n21691_), .ZN(new_n21692_));
  NAND2_X1   g21499(.A1(new_n21692_), .A2(new_n21689_), .ZN(new_n21693_));
  OAI22_X1   g21500(.A1(new_n21690_), .A2(new_n4973_), .B1(new_n21688_), .B2(new_n21686_), .ZN(new_n21694_));
  AOI21_X1   g21501(.A1(new_n21694_), .A2(\asqrt[38] ), .B(new_n21400_), .ZN(new_n21695_));
  NOR2_X1    g21502(.A1(new_n21695_), .A2(new_n21693_), .ZN(new_n21696_));
  AOI22_X1   g21503(.A1(new_n21694_), .A2(\asqrt[38] ), .B1(new_n21692_), .B2(new_n21689_), .ZN(new_n21697_));
  INV_X1     g21504(.I(new_n21408_), .ZN(new_n21698_));
  OAI21_X1   g21505(.A1(new_n21697_), .A2(new_n4330_), .B(new_n21698_), .ZN(new_n21699_));
  NAND2_X1   g21506(.A1(new_n21699_), .A2(new_n21696_), .ZN(new_n21700_));
  OAI22_X1   g21507(.A1(new_n21697_), .A2(new_n4330_), .B1(new_n21695_), .B2(new_n21693_), .ZN(new_n21701_));
  AOI21_X1   g21508(.A1(new_n21701_), .A2(\asqrt[40] ), .B(new_n21415_), .ZN(new_n21702_));
  NOR2_X1    g21509(.A1(new_n21702_), .A2(new_n21700_), .ZN(new_n21703_));
  AOI22_X1   g21510(.A1(new_n21701_), .A2(\asqrt[40] ), .B1(new_n21699_), .B2(new_n21696_), .ZN(new_n21704_));
  INV_X1     g21511(.I(new_n21423_), .ZN(new_n21705_));
  OAI21_X1   g21512(.A1(new_n21704_), .A2(new_n3760_), .B(new_n21705_), .ZN(new_n21706_));
  NAND2_X1   g21513(.A1(new_n21706_), .A2(new_n21703_), .ZN(new_n21707_));
  OAI22_X1   g21514(.A1(new_n21704_), .A2(new_n3760_), .B1(new_n21702_), .B2(new_n21700_), .ZN(new_n21708_));
  AOI21_X1   g21515(.A1(new_n21708_), .A2(\asqrt[42] ), .B(new_n21430_), .ZN(new_n21709_));
  NOR2_X1    g21516(.A1(new_n21709_), .A2(new_n21707_), .ZN(new_n21710_));
  AOI22_X1   g21517(.A1(new_n21708_), .A2(\asqrt[42] ), .B1(new_n21706_), .B2(new_n21703_), .ZN(new_n21711_));
  INV_X1     g21518(.I(new_n21438_), .ZN(new_n21712_));
  OAI21_X1   g21519(.A1(new_n21711_), .A2(new_n3208_), .B(new_n21712_), .ZN(new_n21713_));
  NAND2_X1   g21520(.A1(new_n21713_), .A2(new_n21710_), .ZN(new_n21714_));
  OAI22_X1   g21521(.A1(new_n21711_), .A2(new_n3208_), .B1(new_n21709_), .B2(new_n21707_), .ZN(new_n21715_));
  AOI21_X1   g21522(.A1(new_n21715_), .A2(\asqrt[44] ), .B(new_n21445_), .ZN(new_n21716_));
  NOR2_X1    g21523(.A1(new_n21716_), .A2(new_n21714_), .ZN(new_n21717_));
  AOI22_X1   g21524(.A1(new_n21715_), .A2(\asqrt[44] ), .B1(new_n21713_), .B2(new_n21710_), .ZN(new_n21718_));
  INV_X1     g21525(.I(new_n21453_), .ZN(new_n21719_));
  OAI21_X1   g21526(.A1(new_n21718_), .A2(new_n2728_), .B(new_n21719_), .ZN(new_n21720_));
  NAND2_X1   g21527(.A1(new_n21720_), .A2(new_n21717_), .ZN(new_n21721_));
  OAI22_X1   g21528(.A1(new_n21718_), .A2(new_n2728_), .B1(new_n21716_), .B2(new_n21714_), .ZN(new_n21722_));
  AOI21_X1   g21529(.A1(new_n21722_), .A2(\asqrt[46] ), .B(new_n21460_), .ZN(new_n21723_));
  NOR2_X1    g21530(.A1(new_n21723_), .A2(new_n21721_), .ZN(new_n21724_));
  AOI22_X1   g21531(.A1(new_n21722_), .A2(\asqrt[46] ), .B1(new_n21720_), .B2(new_n21717_), .ZN(new_n21725_));
  INV_X1     g21532(.I(new_n21468_), .ZN(new_n21726_));
  OAI21_X1   g21533(.A1(new_n21725_), .A2(new_n2253_), .B(new_n21726_), .ZN(new_n21727_));
  NAND2_X1   g21534(.A1(new_n21727_), .A2(new_n21724_), .ZN(new_n21728_));
  OAI22_X1   g21535(.A1(new_n21725_), .A2(new_n2253_), .B1(new_n21723_), .B2(new_n21721_), .ZN(new_n21729_));
  AOI21_X1   g21536(.A1(new_n21729_), .A2(\asqrt[48] ), .B(new_n21475_), .ZN(new_n21730_));
  NOR2_X1    g21537(.A1(new_n21730_), .A2(new_n21728_), .ZN(new_n21731_));
  AOI22_X1   g21538(.A1(new_n21729_), .A2(\asqrt[48] ), .B1(new_n21727_), .B2(new_n21724_), .ZN(new_n21732_));
  INV_X1     g21539(.I(new_n21483_), .ZN(new_n21733_));
  OAI21_X1   g21540(.A1(new_n21732_), .A2(new_n1854_), .B(new_n21733_), .ZN(new_n21734_));
  NAND2_X1   g21541(.A1(new_n21734_), .A2(new_n21731_), .ZN(new_n21735_));
  OAI22_X1   g21542(.A1(new_n21732_), .A2(new_n1854_), .B1(new_n21730_), .B2(new_n21728_), .ZN(new_n21736_));
  AOI21_X1   g21543(.A1(new_n21736_), .A2(\asqrt[50] ), .B(new_n21490_), .ZN(new_n21737_));
  NOR2_X1    g21544(.A1(new_n21737_), .A2(new_n21735_), .ZN(new_n21738_));
  AOI22_X1   g21545(.A1(new_n21736_), .A2(\asqrt[50] ), .B1(new_n21734_), .B2(new_n21731_), .ZN(new_n21739_));
  INV_X1     g21546(.I(new_n21498_), .ZN(new_n21740_));
  OAI21_X1   g21547(.A1(new_n21739_), .A2(new_n1436_), .B(new_n21740_), .ZN(new_n21741_));
  NAND2_X1   g21548(.A1(new_n21741_), .A2(new_n21738_), .ZN(new_n21742_));
  OAI22_X1   g21549(.A1(new_n21739_), .A2(new_n1436_), .B1(new_n21737_), .B2(new_n21735_), .ZN(new_n21743_));
  AOI21_X1   g21550(.A1(new_n21743_), .A2(\asqrt[52] ), .B(new_n21505_), .ZN(new_n21744_));
  NOR2_X1    g21551(.A1(new_n21744_), .A2(new_n21742_), .ZN(new_n21745_));
  AOI22_X1   g21552(.A1(new_n21743_), .A2(\asqrt[52] ), .B1(new_n21741_), .B2(new_n21738_), .ZN(new_n21746_));
  INV_X1     g21553(.I(new_n21513_), .ZN(new_n21747_));
  OAI21_X1   g21554(.A1(new_n21746_), .A2(new_n1096_), .B(new_n21747_), .ZN(new_n21748_));
  NAND2_X1   g21555(.A1(new_n21748_), .A2(new_n21745_), .ZN(new_n21749_));
  OAI22_X1   g21556(.A1(new_n21746_), .A2(new_n1096_), .B1(new_n21744_), .B2(new_n21742_), .ZN(new_n21750_));
  AOI21_X1   g21557(.A1(new_n21750_), .A2(\asqrt[54] ), .B(new_n21520_), .ZN(new_n21751_));
  NOR2_X1    g21558(.A1(new_n21751_), .A2(new_n21749_), .ZN(new_n21752_));
  AOI22_X1   g21559(.A1(new_n21750_), .A2(\asqrt[54] ), .B1(new_n21748_), .B2(new_n21745_), .ZN(new_n21753_));
  INV_X1     g21560(.I(new_n21527_), .ZN(new_n21754_));
  OAI21_X1   g21561(.A1(new_n21753_), .A2(new_n825_), .B(new_n21754_), .ZN(new_n21755_));
  NAND2_X1   g21562(.A1(new_n21755_), .A2(new_n21752_), .ZN(new_n21756_));
  OAI22_X1   g21563(.A1(new_n21753_), .A2(new_n825_), .B1(new_n21751_), .B2(new_n21749_), .ZN(new_n21757_));
  AOI21_X1   g21564(.A1(new_n21757_), .A2(\asqrt[56] ), .B(new_n21533_), .ZN(new_n21758_));
  NOR2_X1    g21565(.A1(new_n21758_), .A2(new_n21756_), .ZN(new_n21759_));
  AOI22_X1   g21566(.A1(new_n21757_), .A2(\asqrt[56] ), .B1(new_n21755_), .B2(new_n21752_), .ZN(new_n21760_));
  INV_X1     g21567(.I(new_n21540_), .ZN(new_n21761_));
  OAI21_X1   g21568(.A1(new_n21760_), .A2(new_n587_), .B(new_n21761_), .ZN(new_n21762_));
  NAND2_X1   g21569(.A1(new_n21762_), .A2(new_n21759_), .ZN(new_n21763_));
  OAI22_X1   g21570(.A1(new_n21760_), .A2(new_n587_), .B1(new_n21758_), .B2(new_n21756_), .ZN(new_n21764_));
  AOI21_X1   g21571(.A1(new_n21764_), .A2(\asqrt[58] ), .B(new_n21546_), .ZN(new_n21765_));
  NOR2_X1    g21572(.A1(new_n21765_), .A2(new_n21763_), .ZN(new_n21766_));
  AOI22_X1   g21573(.A1(new_n21764_), .A2(\asqrt[58] ), .B1(new_n21762_), .B2(new_n21759_), .ZN(new_n21767_));
  INV_X1     g21574(.I(new_n21553_), .ZN(new_n21768_));
  OAI21_X1   g21575(.A1(new_n21767_), .A2(new_n376_), .B(new_n21768_), .ZN(new_n21769_));
  NAND2_X1   g21576(.A1(new_n21769_), .A2(new_n21766_), .ZN(new_n21770_));
  OAI22_X1   g21577(.A1(new_n21767_), .A2(new_n376_), .B1(new_n21765_), .B2(new_n21763_), .ZN(new_n21771_));
  AOI21_X1   g21578(.A1(new_n21771_), .A2(\asqrt[60] ), .B(new_n21559_), .ZN(new_n21772_));
  AOI22_X1   g21579(.A1(new_n21771_), .A2(\asqrt[60] ), .B1(new_n21769_), .B2(new_n21766_), .ZN(new_n21773_));
  OAI22_X1   g21580(.A1(new_n21773_), .A2(new_n229_), .B1(new_n21772_), .B2(new_n21770_), .ZN(new_n21774_));
  NAND2_X1   g21581(.A1(new_n21774_), .A2(\asqrt[62] ), .ZN(new_n21775_));
  NOR2_X1    g21582(.A1(new_n21772_), .A2(new_n21770_), .ZN(new_n21776_));
  NOR3_X1    g21583(.A1(new_n21773_), .A2(new_n229_), .A3(new_n21569_), .ZN(new_n21777_));
  AOI21_X1   g21584(.A1(new_n21777_), .A2(new_n21776_), .B(new_n21091_), .ZN(new_n21778_));
  AOI21_X1   g21585(.A1(new_n21778_), .A2(new_n21572_), .B(new_n21081_), .ZN(new_n21779_));
  NOR4_X1    g21586(.A1(new_n21774_), .A2(\asqrt[62] ), .A3(new_n21081_), .A4(new_n21090_), .ZN(new_n21780_));
  NOR3_X1    g21587(.A1(new_n21779_), .A2(new_n21780_), .A3(new_n21582_), .ZN(new_n21781_));
  NOR4_X1    g21588(.A1(new_n21781_), .A2(\asqrt[62] ), .A3(new_n21090_), .A4(new_n21774_), .ZN(new_n21782_));
  XOR2_X1    g21589(.A1(new_n21782_), .A2(new_n21775_), .Z(new_n21783_));
  NOR4_X1    g21590(.A1(new_n21781_), .A2(\asqrt[61] ), .A3(new_n21558_), .A4(new_n21576_), .ZN(new_n21784_));
  XOR2_X1    g21591(.A1(new_n21784_), .A2(new_n21567_), .Z(new_n21785_));
  NOR2_X1    g21592(.A1(new_n21785_), .A2(new_n196_), .ZN(new_n21786_));
  INV_X1     g21593(.I(\a[9] ), .ZN(new_n21787_));
  NOR2_X1    g21594(.A1(\a[6] ), .A2(\a[7] ), .ZN(new_n21788_));
  INV_X1     g21595(.I(new_n21788_), .ZN(new_n21789_));
  OAI21_X1   g21596(.A1(\a[8] ), .A2(new_n21789_), .B(new_n21111_), .ZN(new_n21790_));
  NOR2_X1    g21597(.A1(new_n21105_), .A2(new_n21790_), .ZN(new_n21791_));
  XOR2_X1    g21598(.A1(new_n21791_), .A2(new_n21787_), .Z(new_n21792_));
  INV_X1     g21599(.I(new_n21792_), .ZN(new_n21793_));
  OAI21_X1   g21600(.A1(new_n21579_), .A2(new_n21582_), .B(\a[9] ), .ZN(new_n21794_));
  NOR2_X1    g21601(.A1(new_n21792_), .A2(\a[8] ), .ZN(new_n21795_));
  INV_X1     g21602(.I(new_n21795_), .ZN(new_n21796_));
  AOI21_X1   g21603(.A1(new_n21794_), .A2(new_n21796_), .B(new_n21793_), .ZN(new_n21797_));
  INV_X1     g21604(.I(\a[8] ), .ZN(new_n21798_));
  INV_X1     g21605(.I(new_n21091_), .ZN(new_n21799_));
  NAND2_X1   g21606(.A1(new_n21764_), .A2(\asqrt[58] ), .ZN(new_n21800_));
  AOI21_X1   g21607(.A1(new_n21800_), .A2(new_n21763_), .B(new_n376_), .ZN(new_n21801_));
  OAI21_X1   g21608(.A1(new_n21766_), .A2(new_n21801_), .B(\asqrt[60] ), .ZN(new_n21802_));
  AOI21_X1   g21609(.A1(new_n21770_), .A2(new_n21802_), .B(new_n229_), .ZN(new_n21803_));
  INV_X1     g21610(.I(new_n21569_), .ZN(new_n21804_));
  NAND3_X1   g21611(.A1(new_n21776_), .A2(new_n21803_), .A3(new_n21804_), .ZN(new_n21805_));
  NAND3_X1   g21612(.A1(new_n21805_), .A2(new_n21799_), .A3(new_n21572_), .ZN(new_n21806_));
  AOI21_X1   g21613(.A1(new_n21806_), .A2(new_n21575_), .B(new_n21780_), .ZN(new_n21807_));
  AOI21_X1   g21614(.A1(new_n21807_), .A2(new_n21583_), .B(new_n21787_), .ZN(new_n21808_));
  NOR3_X1    g21615(.A1(new_n21808_), .A2(new_n21798_), .A3(new_n21792_), .ZN(new_n21809_));
  NAND3_X1   g21616(.A1(new_n21576_), .A2(\asqrt[61] ), .A3(new_n21804_), .ZN(new_n21810_));
  OAI21_X1   g21617(.A1(new_n21810_), .A2(new_n21562_), .B(new_n21799_), .ZN(new_n21811_));
  OAI21_X1   g21618(.A1(new_n21811_), .A2(new_n21573_), .B(new_n21575_), .ZN(new_n21812_));
  NAND3_X1   g21619(.A1(new_n21812_), .A2(new_n21578_), .A3(new_n21583_), .ZN(\asqrt[4] ));
  NAND3_X1   g21620(.A1(\asqrt[4] ), .A2(\a[8] ), .A3(\asqrt[5] ), .ZN(new_n21814_));
  NAND3_X1   g21621(.A1(new_n21781_), .A2(new_n21798_), .A3(\asqrt[5] ), .ZN(new_n21815_));
  AOI21_X1   g21622(.A1(new_n21815_), .A2(new_n21814_), .B(new_n21789_), .ZN(new_n21816_));
  NOR2_X1    g21623(.A1(new_n21583_), .A2(new_n21079_), .ZN(new_n21817_));
  NAND2_X1   g21624(.A1(new_n21780_), .A2(new_n21817_), .ZN(new_n21818_));
  OAI21_X1   g21625(.A1(new_n21818_), .A2(new_n21812_), .B(new_n21110_), .ZN(new_n21819_));
  NAND3_X1   g21626(.A1(new_n21819_), .A2(new_n21781_), .A3(new_n21093_), .ZN(new_n21820_));
  INV_X1     g21627(.I(new_n21817_), .ZN(new_n21821_));
  NOR2_X1    g21628(.A1(new_n21578_), .A2(new_n21821_), .ZN(new_n21822_));
  AOI21_X1   g21629(.A1(new_n21822_), .A2(new_n21779_), .B(\a[10] ), .ZN(new_n21823_));
  OAI21_X1   g21630(.A1(new_n21823_), .A2(new_n21094_), .B(\asqrt[4] ), .ZN(new_n21824_));
  NAND3_X1   g21631(.A1(new_n21824_), .A2(new_n21820_), .A3(new_n20455_), .ZN(new_n21825_));
  OAI22_X1   g21632(.A1(new_n21825_), .A2(new_n21816_), .B1(new_n21797_), .B2(new_n21809_), .ZN(new_n21826_));
  OAI21_X1   g21633(.A1(new_n21808_), .A2(new_n21795_), .B(new_n21792_), .ZN(new_n21827_));
  NAND3_X1   g21634(.A1(new_n21794_), .A2(\a[8] ), .A3(new_n21793_), .ZN(new_n21828_));
  NAND2_X1   g21635(.A1(new_n21828_), .A2(new_n21827_), .ZN(new_n21829_));
  OAI21_X1   g21636(.A1(new_n21829_), .A2(new_n21816_), .B(\asqrt[6] ), .ZN(new_n21830_));
  NOR2_X1    g21637(.A1(new_n21079_), .A2(\a[10] ), .ZN(new_n21831_));
  OAI22_X1   g21638(.A1(new_n21831_), .A2(\a[11] ), .B1(new_n21106_), .B2(\a[10] ), .ZN(new_n21832_));
  NAND2_X1   g21639(.A1(new_n21131_), .A2(new_n21096_), .ZN(new_n21833_));
  AOI21_X1   g21640(.A1(new_n21833_), .A2(new_n21110_), .B(new_n21079_), .ZN(new_n21834_));
  AOI21_X1   g21641(.A1(\asqrt[4] ), .A2(new_n21834_), .B(new_n21832_), .ZN(new_n21835_));
  NAND2_X1   g21642(.A1(new_n21834_), .A2(new_n21832_), .ZN(new_n21836_));
  NOR2_X1    g21643(.A1(new_n21781_), .A2(new_n21836_), .ZN(new_n21837_));
  NOR2_X1    g21644(.A1(new_n21835_), .A2(new_n21837_), .ZN(new_n21838_));
  NAND2_X1   g21645(.A1(new_n21838_), .A2(new_n19782_), .ZN(new_n21839_));
  INV_X1     g21646(.I(new_n21839_), .ZN(new_n21840_));
  AOI21_X1   g21647(.A1(new_n21830_), .A2(new_n21840_), .B(new_n21826_), .ZN(new_n21841_));
  AOI21_X1   g21648(.A1(new_n21830_), .A2(new_n21826_), .B(new_n19782_), .ZN(new_n21842_));
  NOR2_X1    g21649(.A1(new_n21176_), .A2(new_n21177_), .ZN(new_n21843_));
  NOR4_X1    g21650(.A1(new_n21781_), .A2(\asqrt[7] ), .A3(new_n21843_), .A4(new_n21180_), .ZN(new_n21844_));
  NAND2_X1   g21651(.A1(new_n21844_), .A2(new_n21145_), .ZN(new_n21845_));
  OAI21_X1   g21652(.A1(new_n21144_), .A2(new_n21131_), .B(\asqrt[7] ), .ZN(new_n21846_));
  NAND2_X1   g21653(.A1(new_n21846_), .A2(new_n21845_), .ZN(new_n21847_));
  NOR2_X1    g21654(.A1(new_n21847_), .A2(\asqrt[8] ), .ZN(new_n21848_));
  INV_X1     g21655(.I(new_n21848_), .ZN(new_n21849_));
  OAI21_X1   g21656(.A1(new_n21842_), .A2(new_n21849_), .B(new_n21841_), .ZN(new_n21850_));
  OAI21_X1   g21657(.A1(new_n21841_), .A2(new_n21842_), .B(\asqrt[8] ), .ZN(new_n21851_));
  NAND2_X1   g21658(.A1(new_n21151_), .A2(new_n21152_), .ZN(new_n21852_));
  AND4_X2    g21659(.A1(new_n19100_), .A2(\asqrt[4] ), .A3(new_n21852_), .A4(new_n21181_), .Z(new_n21853_));
  XNOR2_X1   g21660(.A1(new_n21853_), .A2(new_n21156_), .ZN(new_n21854_));
  NAND2_X1   g21661(.A1(new_n21854_), .A2(new_n18495_), .ZN(new_n21855_));
  INV_X1     g21662(.I(new_n21855_), .ZN(new_n21856_));
  AOI21_X1   g21663(.A1(new_n21851_), .A2(new_n21856_), .B(new_n21850_), .ZN(new_n21857_));
  AOI21_X1   g21664(.A1(new_n21850_), .A2(new_n21851_), .B(new_n18495_), .ZN(new_n21858_));
  NOR2_X1    g21665(.A1(new_n21161_), .A2(new_n21158_), .ZN(new_n21859_));
  NOR4_X1    g21666(.A1(new_n21781_), .A2(\asqrt[9] ), .A3(new_n21859_), .A4(new_n21184_), .ZN(new_n21860_));
  XOR2_X1    g21667(.A1(new_n21860_), .A2(new_n21165_), .Z(new_n21861_));
  INV_X1     g21668(.I(new_n21861_), .ZN(new_n21862_));
  NOR2_X1    g21669(.A1(new_n21862_), .A2(\asqrt[10] ), .ZN(new_n21863_));
  INV_X1     g21670(.I(new_n21863_), .ZN(new_n21864_));
  OAI21_X1   g21671(.A1(new_n21858_), .A2(new_n21864_), .B(new_n21857_), .ZN(new_n21865_));
  OAI21_X1   g21672(.A1(new_n21857_), .A2(new_n21858_), .B(\asqrt[10] ), .ZN(new_n21866_));
  NOR4_X1    g21673(.A1(new_n21781_), .A2(\asqrt[10] ), .A3(new_n21169_), .A4(new_n21594_), .ZN(new_n21867_));
  XNOR2_X1   g21674(.A1(new_n21867_), .A2(new_n21597_), .ZN(new_n21868_));
  NAND2_X1   g21675(.A1(new_n21868_), .A2(new_n17271_), .ZN(new_n21869_));
  INV_X1     g21676(.I(new_n21869_), .ZN(new_n21870_));
  AOI21_X1   g21677(.A1(new_n21866_), .A2(new_n21870_), .B(new_n21865_), .ZN(new_n21871_));
  NAND2_X1   g21678(.A1(\asqrt[5] ), .A2(\a[8] ), .ZN(new_n21872_));
  AOI21_X1   g21679(.A1(new_n21781_), .A2(\asqrt[5] ), .B(new_n21872_), .ZN(new_n21873_));
  NOR4_X1    g21680(.A1(new_n21579_), .A2(\a[8] ), .A3(new_n21079_), .A4(new_n21582_), .ZN(new_n21874_));
  OAI21_X1   g21681(.A1(new_n21873_), .A2(new_n21874_), .B(new_n21788_), .ZN(new_n21875_));
  NOR3_X1    g21682(.A1(new_n21823_), .A2(\asqrt[4] ), .A3(new_n21094_), .ZN(new_n21876_));
  AOI21_X1   g21683(.A1(new_n21819_), .A2(new_n21093_), .B(new_n21781_), .ZN(new_n21877_));
  NOR3_X1    g21684(.A1(new_n21877_), .A2(new_n21876_), .A3(\asqrt[6] ), .ZN(new_n21878_));
  NAND2_X1   g21685(.A1(new_n21878_), .A2(new_n21875_), .ZN(new_n21879_));
  NAND3_X1   g21686(.A1(new_n21875_), .A2(new_n21827_), .A3(new_n21828_), .ZN(new_n21880_));
  AOI22_X1   g21687(.A1(new_n21879_), .A2(new_n21829_), .B1(new_n21880_), .B2(\asqrt[6] ), .ZN(new_n21881_));
  OAI21_X1   g21688(.A1(new_n21881_), .A2(new_n19782_), .B(new_n21848_), .ZN(new_n21882_));
  AOI21_X1   g21689(.A1(new_n21880_), .A2(\asqrt[6] ), .B(new_n21839_), .ZN(new_n21883_));
  OAI22_X1   g21690(.A1(new_n21881_), .A2(new_n19782_), .B1(new_n21826_), .B2(new_n21883_), .ZN(new_n21884_));
  AOI22_X1   g21691(.A1(new_n21884_), .A2(\asqrt[8] ), .B1(new_n21882_), .B2(new_n21841_), .ZN(new_n21885_));
  OAI21_X1   g21692(.A1(new_n21885_), .A2(new_n18495_), .B(new_n21863_), .ZN(new_n21886_));
  AOI21_X1   g21693(.A1(new_n21884_), .A2(\asqrt[8] ), .B(new_n21855_), .ZN(new_n21887_));
  OAI22_X1   g21694(.A1(new_n21885_), .A2(new_n18495_), .B1(new_n21887_), .B2(new_n21850_), .ZN(new_n21888_));
  AOI22_X1   g21695(.A1(new_n21888_), .A2(\asqrt[10] ), .B1(new_n21886_), .B2(new_n21857_), .ZN(new_n21889_));
  NOR4_X1    g21696(.A1(new_n21781_), .A2(\asqrt[11] ), .A3(new_n21188_), .A4(new_n21194_), .ZN(new_n21890_));
  XOR2_X1    g21697(.A1(new_n21890_), .A2(new_n21598_), .Z(new_n21891_));
  NAND2_X1   g21698(.A1(new_n21891_), .A2(new_n16619_), .ZN(new_n21892_));
  INV_X1     g21699(.I(new_n21892_), .ZN(new_n21893_));
  OAI21_X1   g21700(.A1(new_n21889_), .A2(new_n17271_), .B(new_n21893_), .ZN(new_n21894_));
  NAND2_X1   g21701(.A1(new_n21894_), .A2(new_n21871_), .ZN(new_n21895_));
  AOI21_X1   g21702(.A1(new_n21888_), .A2(\asqrt[10] ), .B(new_n21869_), .ZN(new_n21896_));
  OAI22_X1   g21703(.A1(new_n21889_), .A2(new_n17271_), .B1(new_n21896_), .B2(new_n21865_), .ZN(new_n21897_));
  NOR2_X1    g21704(.A1(new_n21201_), .A2(new_n16619_), .ZN(new_n21898_));
  NOR4_X1    g21705(.A1(new_n21781_), .A2(\asqrt[12] ), .A3(new_n21197_), .A4(new_n21603_), .ZN(new_n21899_));
  XNOR2_X1   g21706(.A1(new_n21899_), .A2(new_n21898_), .ZN(new_n21900_));
  NAND2_X1   g21707(.A1(new_n21900_), .A2(new_n16060_), .ZN(new_n21901_));
  AOI21_X1   g21708(.A1(new_n21897_), .A2(\asqrt[12] ), .B(new_n21901_), .ZN(new_n21902_));
  NOR2_X1    g21709(.A1(new_n21902_), .A2(new_n21895_), .ZN(new_n21903_));
  AOI22_X1   g21710(.A1(new_n21897_), .A2(\asqrt[12] ), .B1(new_n21894_), .B2(new_n21871_), .ZN(new_n21904_));
  NAND2_X1   g21711(.A1(new_n21209_), .A2(\asqrt[13] ), .ZN(new_n21905_));
  NOR4_X1    g21712(.A1(new_n21781_), .A2(\asqrt[13] ), .A3(new_n21204_), .A4(new_n21209_), .ZN(new_n21906_));
  XOR2_X1    g21713(.A1(new_n21906_), .A2(new_n21905_), .Z(new_n21907_));
  NAND2_X1   g21714(.A1(new_n21907_), .A2(new_n15447_), .ZN(new_n21908_));
  INV_X1     g21715(.I(new_n21908_), .ZN(new_n21909_));
  OAI21_X1   g21716(.A1(new_n21904_), .A2(new_n16060_), .B(new_n21909_), .ZN(new_n21910_));
  NAND2_X1   g21717(.A1(new_n21910_), .A2(new_n21903_), .ZN(new_n21911_));
  OAI22_X1   g21718(.A1(new_n21904_), .A2(new_n16060_), .B1(new_n21902_), .B2(new_n21895_), .ZN(new_n21912_));
  NOR2_X1    g21719(.A1(new_n21216_), .A2(new_n15447_), .ZN(new_n21913_));
  NOR4_X1    g21720(.A1(new_n21781_), .A2(\asqrt[14] ), .A3(new_n21212_), .A4(new_n21610_), .ZN(new_n21914_));
  XNOR2_X1   g21721(.A1(new_n21914_), .A2(new_n21913_), .ZN(new_n21915_));
  NAND2_X1   g21722(.A1(new_n21915_), .A2(new_n14871_), .ZN(new_n21916_));
  AOI21_X1   g21723(.A1(new_n21912_), .A2(\asqrt[14] ), .B(new_n21916_), .ZN(new_n21917_));
  NOR2_X1    g21724(.A1(new_n21917_), .A2(new_n21911_), .ZN(new_n21918_));
  AOI22_X1   g21725(.A1(new_n21912_), .A2(\asqrt[14] ), .B1(new_n21910_), .B2(new_n21903_), .ZN(new_n21919_));
  NAND2_X1   g21726(.A1(new_n21224_), .A2(\asqrt[15] ), .ZN(new_n21920_));
  NOR4_X1    g21727(.A1(new_n21781_), .A2(\asqrt[15] ), .A3(new_n21219_), .A4(new_n21224_), .ZN(new_n21921_));
  XOR2_X1    g21728(.A1(new_n21921_), .A2(new_n21920_), .Z(new_n21922_));
  NAND2_X1   g21729(.A1(new_n21922_), .A2(new_n14273_), .ZN(new_n21923_));
  INV_X1     g21730(.I(new_n21923_), .ZN(new_n21924_));
  OAI21_X1   g21731(.A1(new_n21919_), .A2(new_n14871_), .B(new_n21924_), .ZN(new_n21925_));
  NAND2_X1   g21732(.A1(new_n21925_), .A2(new_n21918_), .ZN(new_n21926_));
  OAI22_X1   g21733(.A1(new_n21919_), .A2(new_n14871_), .B1(new_n21917_), .B2(new_n21911_), .ZN(new_n21927_));
  NOR4_X1    g21734(.A1(new_n21781_), .A2(\asqrt[16] ), .A3(new_n21227_), .A4(new_n21617_), .ZN(new_n21928_));
  AOI21_X1   g21735(.A1(new_n21920_), .A2(new_n21223_), .B(new_n14273_), .ZN(new_n21929_));
  NOR2_X1    g21736(.A1(new_n21928_), .A2(new_n21929_), .ZN(new_n21930_));
  NAND2_X1   g21737(.A1(new_n21930_), .A2(new_n13760_), .ZN(new_n21931_));
  AOI21_X1   g21738(.A1(new_n21927_), .A2(\asqrt[16] ), .B(new_n21931_), .ZN(new_n21932_));
  NOR2_X1    g21739(.A1(new_n21932_), .A2(new_n21926_), .ZN(new_n21933_));
  AOI22_X1   g21740(.A1(new_n21927_), .A2(\asqrt[16] ), .B1(new_n21925_), .B2(new_n21918_), .ZN(new_n21934_));
  NAND2_X1   g21741(.A1(new_n21239_), .A2(\asqrt[17] ), .ZN(new_n21935_));
  NOR4_X1    g21742(.A1(new_n21781_), .A2(\asqrt[17] ), .A3(new_n21234_), .A4(new_n21239_), .ZN(new_n21936_));
  XOR2_X1    g21743(.A1(new_n21936_), .A2(new_n21935_), .Z(new_n21937_));
  NAND2_X1   g21744(.A1(new_n21937_), .A2(new_n13192_), .ZN(new_n21938_));
  INV_X1     g21745(.I(new_n21938_), .ZN(new_n21939_));
  OAI21_X1   g21746(.A1(new_n21934_), .A2(new_n13760_), .B(new_n21939_), .ZN(new_n21940_));
  NAND2_X1   g21747(.A1(new_n21940_), .A2(new_n21933_), .ZN(new_n21941_));
  OAI22_X1   g21748(.A1(new_n21934_), .A2(new_n13760_), .B1(new_n21932_), .B2(new_n21926_), .ZN(new_n21942_));
  NOR4_X1    g21749(.A1(new_n21781_), .A2(\asqrt[18] ), .A3(new_n21242_), .A4(new_n21624_), .ZN(new_n21943_));
  AOI21_X1   g21750(.A1(new_n21935_), .A2(new_n21238_), .B(new_n13192_), .ZN(new_n21944_));
  NOR2_X1    g21751(.A1(new_n21943_), .A2(new_n21944_), .ZN(new_n21945_));
  NAND2_X1   g21752(.A1(new_n21945_), .A2(new_n12657_), .ZN(new_n21946_));
  AOI21_X1   g21753(.A1(new_n21942_), .A2(\asqrt[18] ), .B(new_n21946_), .ZN(new_n21947_));
  NOR2_X1    g21754(.A1(new_n21947_), .A2(new_n21941_), .ZN(new_n21948_));
  AOI22_X1   g21755(.A1(new_n21942_), .A2(\asqrt[18] ), .B1(new_n21940_), .B2(new_n21933_), .ZN(new_n21949_));
  NAND2_X1   g21756(.A1(new_n21254_), .A2(\asqrt[19] ), .ZN(new_n21950_));
  NOR4_X1    g21757(.A1(new_n21781_), .A2(\asqrt[19] ), .A3(new_n21249_), .A4(new_n21254_), .ZN(new_n21951_));
  XOR2_X1    g21758(.A1(new_n21951_), .A2(new_n21950_), .Z(new_n21952_));
  NAND2_X1   g21759(.A1(new_n21952_), .A2(new_n12101_), .ZN(new_n21953_));
  INV_X1     g21760(.I(new_n21953_), .ZN(new_n21954_));
  OAI21_X1   g21761(.A1(new_n21949_), .A2(new_n12657_), .B(new_n21954_), .ZN(new_n21955_));
  NAND2_X1   g21762(.A1(new_n21955_), .A2(new_n21948_), .ZN(new_n21956_));
  OAI22_X1   g21763(.A1(new_n21949_), .A2(new_n12657_), .B1(new_n21947_), .B2(new_n21941_), .ZN(new_n21957_));
  NOR4_X1    g21764(.A1(new_n21781_), .A2(\asqrt[20] ), .A3(new_n21257_), .A4(new_n21631_), .ZN(new_n21958_));
  AOI21_X1   g21765(.A1(new_n21950_), .A2(new_n21253_), .B(new_n12101_), .ZN(new_n21959_));
  NOR2_X1    g21766(.A1(new_n21958_), .A2(new_n21959_), .ZN(new_n21960_));
  NAND2_X1   g21767(.A1(new_n21960_), .A2(new_n11631_), .ZN(new_n21961_));
  AOI21_X1   g21768(.A1(new_n21957_), .A2(\asqrt[20] ), .B(new_n21961_), .ZN(new_n21962_));
  NOR2_X1    g21769(.A1(new_n21962_), .A2(new_n21956_), .ZN(new_n21963_));
  AOI22_X1   g21770(.A1(new_n21957_), .A2(\asqrt[20] ), .B1(new_n21955_), .B2(new_n21948_), .ZN(new_n21964_));
  NAND2_X1   g21771(.A1(new_n21269_), .A2(\asqrt[21] ), .ZN(new_n21965_));
  NOR4_X1    g21772(.A1(new_n21781_), .A2(\asqrt[21] ), .A3(new_n21264_), .A4(new_n21269_), .ZN(new_n21966_));
  XOR2_X1    g21773(.A1(new_n21966_), .A2(new_n21965_), .Z(new_n21967_));
  NAND2_X1   g21774(.A1(new_n21967_), .A2(new_n11105_), .ZN(new_n21968_));
  INV_X1     g21775(.I(new_n21968_), .ZN(new_n21969_));
  OAI21_X1   g21776(.A1(new_n21964_), .A2(new_n11631_), .B(new_n21969_), .ZN(new_n21970_));
  NAND2_X1   g21777(.A1(new_n21970_), .A2(new_n21963_), .ZN(new_n21971_));
  OAI22_X1   g21778(.A1(new_n21964_), .A2(new_n11631_), .B1(new_n21962_), .B2(new_n21956_), .ZN(new_n21972_));
  NOR4_X1    g21779(.A1(new_n21781_), .A2(\asqrt[22] ), .A3(new_n21272_), .A4(new_n21638_), .ZN(new_n21973_));
  AOI21_X1   g21780(.A1(new_n21965_), .A2(new_n21268_), .B(new_n11105_), .ZN(new_n21974_));
  NOR2_X1    g21781(.A1(new_n21973_), .A2(new_n21974_), .ZN(new_n21975_));
  NAND2_X1   g21782(.A1(new_n21975_), .A2(new_n10614_), .ZN(new_n21976_));
  AOI21_X1   g21783(.A1(new_n21972_), .A2(\asqrt[22] ), .B(new_n21976_), .ZN(new_n21977_));
  NOR2_X1    g21784(.A1(new_n21977_), .A2(new_n21971_), .ZN(new_n21978_));
  AOI22_X1   g21785(.A1(new_n21972_), .A2(\asqrt[22] ), .B1(new_n21970_), .B2(new_n21963_), .ZN(new_n21979_));
  NAND2_X1   g21786(.A1(new_n21284_), .A2(\asqrt[23] ), .ZN(new_n21980_));
  NOR4_X1    g21787(.A1(new_n21781_), .A2(\asqrt[23] ), .A3(new_n21279_), .A4(new_n21284_), .ZN(new_n21981_));
  XOR2_X1    g21788(.A1(new_n21981_), .A2(new_n21980_), .Z(new_n21982_));
  NAND2_X1   g21789(.A1(new_n21982_), .A2(new_n10104_), .ZN(new_n21983_));
  INV_X1     g21790(.I(new_n21983_), .ZN(new_n21984_));
  OAI21_X1   g21791(.A1(new_n21979_), .A2(new_n10614_), .B(new_n21984_), .ZN(new_n21985_));
  NAND2_X1   g21792(.A1(new_n21985_), .A2(new_n21978_), .ZN(new_n21986_));
  OAI22_X1   g21793(.A1(new_n21979_), .A2(new_n10614_), .B1(new_n21977_), .B2(new_n21971_), .ZN(new_n21987_));
  NOR4_X1    g21794(.A1(new_n21781_), .A2(\asqrt[24] ), .A3(new_n21287_), .A4(new_n21645_), .ZN(new_n21988_));
  AOI21_X1   g21795(.A1(new_n21980_), .A2(new_n21283_), .B(new_n10104_), .ZN(new_n21989_));
  NOR2_X1    g21796(.A1(new_n21988_), .A2(new_n21989_), .ZN(new_n21990_));
  NAND2_X1   g21797(.A1(new_n21990_), .A2(new_n9672_), .ZN(new_n21991_));
  AOI21_X1   g21798(.A1(new_n21987_), .A2(\asqrt[24] ), .B(new_n21991_), .ZN(new_n21992_));
  NOR2_X1    g21799(.A1(new_n21992_), .A2(new_n21986_), .ZN(new_n21993_));
  AOI22_X1   g21800(.A1(new_n21987_), .A2(\asqrt[24] ), .B1(new_n21985_), .B2(new_n21978_), .ZN(new_n21994_));
  NAND2_X1   g21801(.A1(new_n21299_), .A2(\asqrt[25] ), .ZN(new_n21995_));
  NOR4_X1    g21802(.A1(new_n21781_), .A2(\asqrt[25] ), .A3(new_n21294_), .A4(new_n21299_), .ZN(new_n21996_));
  XOR2_X1    g21803(.A1(new_n21996_), .A2(new_n21995_), .Z(new_n21997_));
  NAND2_X1   g21804(.A1(new_n21997_), .A2(new_n9212_), .ZN(new_n21998_));
  INV_X1     g21805(.I(new_n21998_), .ZN(new_n21999_));
  OAI21_X1   g21806(.A1(new_n21994_), .A2(new_n9672_), .B(new_n21999_), .ZN(new_n22000_));
  NAND2_X1   g21807(.A1(new_n22000_), .A2(new_n21993_), .ZN(new_n22001_));
  OAI22_X1   g21808(.A1(new_n21994_), .A2(new_n9672_), .B1(new_n21992_), .B2(new_n21986_), .ZN(new_n22002_));
  NOR4_X1    g21809(.A1(new_n21781_), .A2(\asqrt[26] ), .A3(new_n21302_), .A4(new_n21652_), .ZN(new_n22003_));
  AOI21_X1   g21810(.A1(new_n21995_), .A2(new_n21298_), .B(new_n9212_), .ZN(new_n22004_));
  NOR2_X1    g21811(.A1(new_n22003_), .A2(new_n22004_), .ZN(new_n22005_));
  NAND2_X1   g21812(.A1(new_n22005_), .A2(new_n8763_), .ZN(new_n22006_));
  AOI21_X1   g21813(.A1(new_n22002_), .A2(\asqrt[26] ), .B(new_n22006_), .ZN(new_n22007_));
  NOR2_X1    g21814(.A1(new_n22007_), .A2(new_n22001_), .ZN(new_n22008_));
  AOI22_X1   g21815(.A1(new_n22002_), .A2(\asqrt[26] ), .B1(new_n22000_), .B2(new_n21993_), .ZN(new_n22009_));
  NAND2_X1   g21816(.A1(new_n21314_), .A2(\asqrt[27] ), .ZN(new_n22010_));
  NOR4_X1    g21817(.A1(new_n21781_), .A2(\asqrt[27] ), .A3(new_n21309_), .A4(new_n21314_), .ZN(new_n22011_));
  XOR2_X1    g21818(.A1(new_n22011_), .A2(new_n22010_), .Z(new_n22012_));
  NAND2_X1   g21819(.A1(new_n22012_), .A2(new_n8319_), .ZN(new_n22013_));
  INV_X1     g21820(.I(new_n22013_), .ZN(new_n22014_));
  OAI21_X1   g21821(.A1(new_n22009_), .A2(new_n8763_), .B(new_n22014_), .ZN(new_n22015_));
  NAND2_X1   g21822(.A1(new_n22015_), .A2(new_n22008_), .ZN(new_n22016_));
  OAI22_X1   g21823(.A1(new_n22009_), .A2(new_n8763_), .B1(new_n22007_), .B2(new_n22001_), .ZN(new_n22017_));
  NOR4_X1    g21824(.A1(new_n21781_), .A2(\asqrt[28] ), .A3(new_n21317_), .A4(new_n21659_), .ZN(new_n22018_));
  AOI21_X1   g21825(.A1(new_n22010_), .A2(new_n21313_), .B(new_n8319_), .ZN(new_n22019_));
  NOR2_X1    g21826(.A1(new_n22018_), .A2(new_n22019_), .ZN(new_n22020_));
  NAND2_X1   g21827(.A1(new_n22020_), .A2(new_n7931_), .ZN(new_n22021_));
  AOI21_X1   g21828(.A1(new_n22017_), .A2(\asqrt[28] ), .B(new_n22021_), .ZN(new_n22022_));
  NOR2_X1    g21829(.A1(new_n22022_), .A2(new_n22016_), .ZN(new_n22023_));
  AOI22_X1   g21830(.A1(new_n22017_), .A2(\asqrt[28] ), .B1(new_n22015_), .B2(new_n22008_), .ZN(new_n22024_));
  NAND2_X1   g21831(.A1(new_n21329_), .A2(\asqrt[29] ), .ZN(new_n22025_));
  NOR4_X1    g21832(.A1(new_n21781_), .A2(\asqrt[29] ), .A3(new_n21324_), .A4(new_n21329_), .ZN(new_n22026_));
  XOR2_X1    g21833(.A1(new_n22026_), .A2(new_n22025_), .Z(new_n22027_));
  NAND2_X1   g21834(.A1(new_n22027_), .A2(new_n7517_), .ZN(new_n22028_));
  INV_X1     g21835(.I(new_n22028_), .ZN(new_n22029_));
  OAI21_X1   g21836(.A1(new_n22024_), .A2(new_n7931_), .B(new_n22029_), .ZN(new_n22030_));
  NAND2_X1   g21837(.A1(new_n22030_), .A2(new_n22023_), .ZN(new_n22031_));
  OAI22_X1   g21838(.A1(new_n22024_), .A2(new_n7931_), .B1(new_n22022_), .B2(new_n22016_), .ZN(new_n22032_));
  NOR4_X1    g21839(.A1(new_n21781_), .A2(\asqrt[30] ), .A3(new_n21332_), .A4(new_n21666_), .ZN(new_n22033_));
  AOI21_X1   g21840(.A1(new_n22025_), .A2(new_n21328_), .B(new_n7517_), .ZN(new_n22034_));
  NOR2_X1    g21841(.A1(new_n22033_), .A2(new_n22034_), .ZN(new_n22035_));
  NAND2_X1   g21842(.A1(new_n22035_), .A2(new_n7110_), .ZN(new_n22036_));
  AOI21_X1   g21843(.A1(new_n22032_), .A2(\asqrt[30] ), .B(new_n22036_), .ZN(new_n22037_));
  NOR2_X1    g21844(.A1(new_n22037_), .A2(new_n22031_), .ZN(new_n22038_));
  AOI22_X1   g21845(.A1(new_n22032_), .A2(\asqrt[30] ), .B1(new_n22030_), .B2(new_n22023_), .ZN(new_n22039_));
  NAND2_X1   g21846(.A1(new_n21344_), .A2(\asqrt[31] ), .ZN(new_n22040_));
  NOR4_X1    g21847(.A1(new_n21781_), .A2(\asqrt[31] ), .A3(new_n21339_), .A4(new_n21344_), .ZN(new_n22041_));
  XOR2_X1    g21848(.A1(new_n22041_), .A2(new_n22040_), .Z(new_n22042_));
  NAND2_X1   g21849(.A1(new_n22042_), .A2(new_n6708_), .ZN(new_n22043_));
  INV_X1     g21850(.I(new_n22043_), .ZN(new_n22044_));
  OAI21_X1   g21851(.A1(new_n22039_), .A2(new_n7110_), .B(new_n22044_), .ZN(new_n22045_));
  NAND2_X1   g21852(.A1(new_n22045_), .A2(new_n22038_), .ZN(new_n22046_));
  OAI22_X1   g21853(.A1(new_n22039_), .A2(new_n7110_), .B1(new_n22037_), .B2(new_n22031_), .ZN(new_n22047_));
  NOR4_X1    g21854(.A1(new_n21781_), .A2(\asqrt[32] ), .A3(new_n21347_), .A4(new_n21673_), .ZN(new_n22048_));
  AOI21_X1   g21855(.A1(new_n22040_), .A2(new_n21343_), .B(new_n6708_), .ZN(new_n22049_));
  NOR2_X1    g21856(.A1(new_n22048_), .A2(new_n22049_), .ZN(new_n22050_));
  NAND2_X1   g21857(.A1(new_n22050_), .A2(new_n6365_), .ZN(new_n22051_));
  AOI21_X1   g21858(.A1(new_n22047_), .A2(\asqrt[32] ), .B(new_n22051_), .ZN(new_n22052_));
  NOR2_X1    g21859(.A1(new_n22052_), .A2(new_n22046_), .ZN(new_n22053_));
  AOI22_X1   g21860(.A1(new_n22047_), .A2(\asqrt[32] ), .B1(new_n22045_), .B2(new_n22038_), .ZN(new_n22054_));
  NAND2_X1   g21861(.A1(new_n21359_), .A2(\asqrt[33] ), .ZN(new_n22055_));
  NOR4_X1    g21862(.A1(new_n21781_), .A2(\asqrt[33] ), .A3(new_n21354_), .A4(new_n21359_), .ZN(new_n22056_));
  XOR2_X1    g21863(.A1(new_n22056_), .A2(new_n22055_), .Z(new_n22057_));
  NAND2_X1   g21864(.A1(new_n22057_), .A2(new_n5991_), .ZN(new_n22058_));
  INV_X1     g21865(.I(new_n22058_), .ZN(new_n22059_));
  OAI21_X1   g21866(.A1(new_n22054_), .A2(new_n6365_), .B(new_n22059_), .ZN(new_n22060_));
  NAND2_X1   g21867(.A1(new_n22060_), .A2(new_n22053_), .ZN(new_n22061_));
  OAI22_X1   g21868(.A1(new_n22054_), .A2(new_n6365_), .B1(new_n22052_), .B2(new_n22046_), .ZN(new_n22062_));
  NOR4_X1    g21869(.A1(new_n21781_), .A2(\asqrt[34] ), .A3(new_n21362_), .A4(new_n21680_), .ZN(new_n22063_));
  AOI21_X1   g21870(.A1(new_n22055_), .A2(new_n21358_), .B(new_n5991_), .ZN(new_n22064_));
  NOR2_X1    g21871(.A1(new_n22063_), .A2(new_n22064_), .ZN(new_n22065_));
  NAND2_X1   g21872(.A1(new_n22065_), .A2(new_n5626_), .ZN(new_n22066_));
  AOI21_X1   g21873(.A1(new_n22062_), .A2(\asqrt[34] ), .B(new_n22066_), .ZN(new_n22067_));
  NOR2_X1    g21874(.A1(new_n22067_), .A2(new_n22061_), .ZN(new_n22068_));
  AOI22_X1   g21875(.A1(new_n22062_), .A2(\asqrt[34] ), .B1(new_n22060_), .B2(new_n22053_), .ZN(new_n22069_));
  NAND2_X1   g21876(.A1(new_n21374_), .A2(\asqrt[35] ), .ZN(new_n22070_));
  NOR4_X1    g21877(.A1(new_n21781_), .A2(\asqrt[35] ), .A3(new_n21369_), .A4(new_n21374_), .ZN(new_n22071_));
  XOR2_X1    g21878(.A1(new_n22071_), .A2(new_n22070_), .Z(new_n22072_));
  NAND2_X1   g21879(.A1(new_n22072_), .A2(new_n5273_), .ZN(new_n22073_));
  INV_X1     g21880(.I(new_n22073_), .ZN(new_n22074_));
  OAI21_X1   g21881(.A1(new_n22069_), .A2(new_n5626_), .B(new_n22074_), .ZN(new_n22075_));
  NAND2_X1   g21882(.A1(new_n22075_), .A2(new_n22068_), .ZN(new_n22076_));
  OAI22_X1   g21883(.A1(new_n22069_), .A2(new_n5626_), .B1(new_n22067_), .B2(new_n22061_), .ZN(new_n22077_));
  NOR4_X1    g21884(.A1(new_n21781_), .A2(\asqrt[36] ), .A3(new_n21377_), .A4(new_n21687_), .ZN(new_n22078_));
  AOI21_X1   g21885(.A1(new_n22070_), .A2(new_n21373_), .B(new_n5273_), .ZN(new_n22079_));
  NOR2_X1    g21886(.A1(new_n22078_), .A2(new_n22079_), .ZN(new_n22080_));
  NAND2_X1   g21887(.A1(new_n22080_), .A2(new_n4973_), .ZN(new_n22081_));
  AOI21_X1   g21888(.A1(new_n22077_), .A2(\asqrt[36] ), .B(new_n22081_), .ZN(new_n22082_));
  NOR2_X1    g21889(.A1(new_n22082_), .A2(new_n22076_), .ZN(new_n22083_));
  AOI22_X1   g21890(.A1(new_n22077_), .A2(\asqrt[36] ), .B1(new_n22075_), .B2(new_n22068_), .ZN(new_n22084_));
  NAND2_X1   g21891(.A1(new_n21389_), .A2(\asqrt[37] ), .ZN(new_n22085_));
  NOR4_X1    g21892(.A1(new_n21781_), .A2(\asqrt[37] ), .A3(new_n21384_), .A4(new_n21389_), .ZN(new_n22086_));
  XOR2_X1    g21893(.A1(new_n22086_), .A2(new_n22085_), .Z(new_n22087_));
  INV_X1     g21894(.I(new_n22087_), .ZN(new_n22088_));
  NOR2_X1    g21895(.A1(new_n22088_), .A2(\asqrt[38] ), .ZN(new_n22089_));
  OAI21_X1   g21896(.A1(new_n22084_), .A2(new_n4973_), .B(new_n22089_), .ZN(new_n22090_));
  NAND2_X1   g21897(.A1(new_n22090_), .A2(new_n22083_), .ZN(new_n22091_));
  OAI22_X1   g21898(.A1(new_n22084_), .A2(new_n4973_), .B1(new_n22082_), .B2(new_n22076_), .ZN(new_n22092_));
  NOR4_X1    g21899(.A1(new_n21781_), .A2(\asqrt[38] ), .A3(new_n21392_), .A4(new_n21694_), .ZN(new_n22093_));
  AOI21_X1   g21900(.A1(new_n22085_), .A2(new_n21388_), .B(new_n4645_), .ZN(new_n22094_));
  NOR2_X1    g21901(.A1(new_n22093_), .A2(new_n22094_), .ZN(new_n22095_));
  NAND2_X1   g21902(.A1(new_n22095_), .A2(new_n4330_), .ZN(new_n22096_));
  AOI21_X1   g21903(.A1(new_n22092_), .A2(\asqrt[38] ), .B(new_n22096_), .ZN(new_n22097_));
  NOR2_X1    g21904(.A1(new_n22097_), .A2(new_n22091_), .ZN(new_n22098_));
  AOI22_X1   g21905(.A1(new_n22092_), .A2(\asqrt[38] ), .B1(new_n22090_), .B2(new_n22083_), .ZN(new_n22099_));
  NAND2_X1   g21906(.A1(new_n21404_), .A2(\asqrt[39] ), .ZN(new_n22100_));
  NOR4_X1    g21907(.A1(new_n21781_), .A2(\asqrt[39] ), .A3(new_n21399_), .A4(new_n21404_), .ZN(new_n22101_));
  XOR2_X1    g21908(.A1(new_n22101_), .A2(new_n22100_), .Z(new_n22102_));
  INV_X1     g21909(.I(new_n22102_), .ZN(new_n22103_));
  NOR2_X1    g21910(.A1(new_n22103_), .A2(\asqrt[40] ), .ZN(new_n22104_));
  OAI21_X1   g21911(.A1(new_n22099_), .A2(new_n4330_), .B(new_n22104_), .ZN(new_n22105_));
  NAND2_X1   g21912(.A1(new_n22105_), .A2(new_n22098_), .ZN(new_n22106_));
  OAI22_X1   g21913(.A1(new_n22099_), .A2(new_n4330_), .B1(new_n22097_), .B2(new_n22091_), .ZN(new_n22107_));
  NAND2_X1   g21914(.A1(new_n21701_), .A2(\asqrt[40] ), .ZN(new_n22108_));
  NOR4_X1    g21915(.A1(new_n21781_), .A2(\asqrt[40] ), .A3(new_n21407_), .A4(new_n21701_), .ZN(new_n22109_));
  XOR2_X1    g21916(.A1(new_n22109_), .A2(new_n22108_), .Z(new_n22110_));
  NAND2_X1   g21917(.A1(new_n22110_), .A2(new_n3760_), .ZN(new_n22111_));
  AOI21_X1   g21918(.A1(new_n22107_), .A2(\asqrt[40] ), .B(new_n22111_), .ZN(new_n22112_));
  NOR2_X1    g21919(.A1(new_n22112_), .A2(new_n22106_), .ZN(new_n22113_));
  AOI22_X1   g21920(.A1(new_n22107_), .A2(\asqrt[40] ), .B1(new_n22105_), .B2(new_n22098_), .ZN(new_n22114_));
  NOR4_X1    g21921(.A1(new_n21781_), .A2(\asqrt[41] ), .A3(new_n21414_), .A4(new_n21419_), .ZN(new_n22115_));
  AOI21_X1   g21922(.A1(new_n22108_), .A2(new_n21700_), .B(new_n3760_), .ZN(new_n22116_));
  NOR2_X1    g21923(.A1(new_n22115_), .A2(new_n22116_), .ZN(new_n22117_));
  INV_X1     g21924(.I(new_n22117_), .ZN(new_n22118_));
  NOR2_X1    g21925(.A1(new_n22118_), .A2(\asqrt[42] ), .ZN(new_n22119_));
  OAI21_X1   g21926(.A1(new_n22114_), .A2(new_n3760_), .B(new_n22119_), .ZN(new_n22120_));
  NAND2_X1   g21927(.A1(new_n22120_), .A2(new_n22113_), .ZN(new_n22121_));
  OAI22_X1   g21928(.A1(new_n22114_), .A2(new_n3760_), .B1(new_n22112_), .B2(new_n22106_), .ZN(new_n22122_));
  NAND2_X1   g21929(.A1(new_n21708_), .A2(\asqrt[42] ), .ZN(new_n22123_));
  NOR4_X1    g21930(.A1(new_n21781_), .A2(\asqrt[42] ), .A3(new_n21422_), .A4(new_n21708_), .ZN(new_n22124_));
  XOR2_X1    g21931(.A1(new_n22124_), .A2(new_n22123_), .Z(new_n22125_));
  NAND2_X1   g21932(.A1(new_n22125_), .A2(new_n3208_), .ZN(new_n22126_));
  AOI21_X1   g21933(.A1(new_n22122_), .A2(\asqrt[42] ), .B(new_n22126_), .ZN(new_n22127_));
  NOR2_X1    g21934(.A1(new_n22127_), .A2(new_n22121_), .ZN(new_n22128_));
  AOI22_X1   g21935(.A1(new_n22122_), .A2(\asqrt[42] ), .B1(new_n22120_), .B2(new_n22113_), .ZN(new_n22129_));
  NOR4_X1    g21936(.A1(new_n21781_), .A2(\asqrt[43] ), .A3(new_n21429_), .A4(new_n21434_), .ZN(new_n22130_));
  AOI21_X1   g21937(.A1(new_n22123_), .A2(new_n21707_), .B(new_n3208_), .ZN(new_n22131_));
  NOR2_X1    g21938(.A1(new_n22130_), .A2(new_n22131_), .ZN(new_n22132_));
  NAND2_X1   g21939(.A1(new_n22132_), .A2(new_n2941_), .ZN(new_n22133_));
  INV_X1     g21940(.I(new_n22133_), .ZN(new_n22134_));
  OAI21_X1   g21941(.A1(new_n22129_), .A2(new_n3208_), .B(new_n22134_), .ZN(new_n22135_));
  NAND2_X1   g21942(.A1(new_n22135_), .A2(new_n22128_), .ZN(new_n22136_));
  OAI22_X1   g21943(.A1(new_n22129_), .A2(new_n3208_), .B1(new_n22127_), .B2(new_n22121_), .ZN(new_n22137_));
  NAND2_X1   g21944(.A1(new_n21715_), .A2(\asqrt[44] ), .ZN(new_n22138_));
  NOR4_X1    g21945(.A1(new_n21781_), .A2(\asqrt[44] ), .A3(new_n21437_), .A4(new_n21715_), .ZN(new_n22139_));
  XOR2_X1    g21946(.A1(new_n22139_), .A2(new_n22138_), .Z(new_n22140_));
  INV_X1     g21947(.I(new_n22140_), .ZN(new_n22141_));
  NOR2_X1    g21948(.A1(new_n22141_), .A2(\asqrt[45] ), .ZN(new_n22142_));
  INV_X1     g21949(.I(new_n22142_), .ZN(new_n22143_));
  AOI21_X1   g21950(.A1(new_n22137_), .A2(\asqrt[44] ), .B(new_n22143_), .ZN(new_n22144_));
  NOR2_X1    g21951(.A1(new_n22144_), .A2(new_n22136_), .ZN(new_n22145_));
  AOI22_X1   g21952(.A1(new_n22137_), .A2(\asqrt[44] ), .B1(new_n22135_), .B2(new_n22128_), .ZN(new_n22146_));
  NOR4_X1    g21953(.A1(new_n21781_), .A2(\asqrt[45] ), .A3(new_n21444_), .A4(new_n21449_), .ZN(new_n22147_));
  AOI21_X1   g21954(.A1(new_n22138_), .A2(new_n21714_), .B(new_n2728_), .ZN(new_n22148_));
  NOR2_X1    g21955(.A1(new_n22147_), .A2(new_n22148_), .ZN(new_n22149_));
  NAND2_X1   g21956(.A1(new_n22149_), .A2(new_n2488_), .ZN(new_n22150_));
  INV_X1     g21957(.I(new_n22150_), .ZN(new_n22151_));
  OAI21_X1   g21958(.A1(new_n22146_), .A2(new_n2728_), .B(new_n22151_), .ZN(new_n22152_));
  NAND2_X1   g21959(.A1(new_n22152_), .A2(new_n22145_), .ZN(new_n22153_));
  OAI22_X1   g21960(.A1(new_n22146_), .A2(new_n2728_), .B1(new_n22144_), .B2(new_n22136_), .ZN(new_n22154_));
  NAND2_X1   g21961(.A1(new_n21722_), .A2(\asqrt[46] ), .ZN(new_n22155_));
  NOR4_X1    g21962(.A1(new_n21781_), .A2(\asqrt[46] ), .A3(new_n21452_), .A4(new_n21722_), .ZN(new_n22156_));
  XOR2_X1    g21963(.A1(new_n22156_), .A2(new_n22155_), .Z(new_n22157_));
  NAND2_X1   g21964(.A1(new_n22157_), .A2(new_n2253_), .ZN(new_n22158_));
  AOI21_X1   g21965(.A1(new_n22154_), .A2(\asqrt[46] ), .B(new_n22158_), .ZN(new_n22159_));
  NOR2_X1    g21966(.A1(new_n22159_), .A2(new_n22153_), .ZN(new_n22160_));
  AOI22_X1   g21967(.A1(new_n22154_), .A2(\asqrt[46] ), .B1(new_n22152_), .B2(new_n22145_), .ZN(new_n22161_));
  NOR4_X1    g21968(.A1(new_n21781_), .A2(\asqrt[47] ), .A3(new_n21459_), .A4(new_n21464_), .ZN(new_n22162_));
  AOI21_X1   g21969(.A1(new_n22155_), .A2(new_n21721_), .B(new_n2253_), .ZN(new_n22163_));
  NOR2_X1    g21970(.A1(new_n22162_), .A2(new_n22163_), .ZN(new_n22164_));
  INV_X1     g21971(.I(new_n22164_), .ZN(new_n22165_));
  NOR2_X1    g21972(.A1(new_n22165_), .A2(\asqrt[48] ), .ZN(new_n22166_));
  OAI21_X1   g21973(.A1(new_n22161_), .A2(new_n2253_), .B(new_n22166_), .ZN(new_n22167_));
  NAND2_X1   g21974(.A1(new_n22167_), .A2(new_n22160_), .ZN(new_n22168_));
  OAI22_X1   g21975(.A1(new_n22161_), .A2(new_n2253_), .B1(new_n22159_), .B2(new_n22153_), .ZN(new_n22169_));
  NAND2_X1   g21976(.A1(new_n21729_), .A2(\asqrt[48] ), .ZN(new_n22170_));
  NOR4_X1    g21977(.A1(new_n21781_), .A2(\asqrt[48] ), .A3(new_n21467_), .A4(new_n21729_), .ZN(new_n22171_));
  XOR2_X1    g21978(.A1(new_n22171_), .A2(new_n22170_), .Z(new_n22172_));
  NAND2_X1   g21979(.A1(new_n22172_), .A2(new_n1854_), .ZN(new_n22173_));
  AOI21_X1   g21980(.A1(new_n22169_), .A2(\asqrt[48] ), .B(new_n22173_), .ZN(new_n22174_));
  NOR2_X1    g21981(.A1(new_n22174_), .A2(new_n22168_), .ZN(new_n22175_));
  AOI22_X1   g21982(.A1(new_n22169_), .A2(\asqrt[48] ), .B1(new_n22167_), .B2(new_n22160_), .ZN(new_n22176_));
  NOR4_X1    g21983(.A1(new_n21781_), .A2(\asqrt[49] ), .A3(new_n21474_), .A4(new_n21479_), .ZN(new_n22177_));
  AOI21_X1   g21984(.A1(new_n22170_), .A2(new_n21728_), .B(new_n1854_), .ZN(new_n22178_));
  NOR2_X1    g21985(.A1(new_n22177_), .A2(new_n22178_), .ZN(new_n22179_));
  INV_X1     g21986(.I(new_n22179_), .ZN(new_n22180_));
  NOR2_X1    g21987(.A1(new_n22180_), .A2(\asqrt[50] ), .ZN(new_n22181_));
  OAI21_X1   g21988(.A1(new_n22176_), .A2(new_n1854_), .B(new_n22181_), .ZN(new_n22182_));
  NAND2_X1   g21989(.A1(new_n22182_), .A2(new_n22175_), .ZN(new_n22183_));
  OAI22_X1   g21990(.A1(new_n22176_), .A2(new_n1854_), .B1(new_n22174_), .B2(new_n22168_), .ZN(new_n22184_));
  NAND2_X1   g21991(.A1(new_n21736_), .A2(\asqrt[50] ), .ZN(new_n22185_));
  NOR4_X1    g21992(.A1(new_n21781_), .A2(\asqrt[50] ), .A3(new_n21482_), .A4(new_n21736_), .ZN(new_n22186_));
  XOR2_X1    g21993(.A1(new_n22186_), .A2(new_n22185_), .Z(new_n22187_));
  NAND2_X1   g21994(.A1(new_n22187_), .A2(new_n1436_), .ZN(new_n22188_));
  AOI21_X1   g21995(.A1(new_n22184_), .A2(\asqrt[50] ), .B(new_n22188_), .ZN(new_n22189_));
  NOR2_X1    g21996(.A1(new_n22189_), .A2(new_n22183_), .ZN(new_n22190_));
  AOI22_X1   g21997(.A1(new_n22184_), .A2(\asqrt[50] ), .B1(new_n22182_), .B2(new_n22175_), .ZN(new_n22191_));
  NAND2_X1   g21998(.A1(new_n21494_), .A2(\asqrt[51] ), .ZN(new_n22192_));
  NOR4_X1    g21999(.A1(new_n21781_), .A2(\asqrt[51] ), .A3(new_n21489_), .A4(new_n21494_), .ZN(new_n22193_));
  XOR2_X1    g22000(.A1(new_n22193_), .A2(new_n22192_), .Z(new_n22194_));
  NAND2_X1   g22001(.A1(new_n22194_), .A2(new_n1260_), .ZN(new_n22195_));
  INV_X1     g22002(.I(new_n22195_), .ZN(new_n22196_));
  OAI21_X1   g22003(.A1(new_n22191_), .A2(new_n1436_), .B(new_n22196_), .ZN(new_n22197_));
  NAND2_X1   g22004(.A1(new_n22197_), .A2(new_n22190_), .ZN(new_n22198_));
  OAI22_X1   g22005(.A1(new_n22191_), .A2(new_n1436_), .B1(new_n22189_), .B2(new_n22183_), .ZN(new_n22199_));
  NOR4_X1    g22006(.A1(new_n21781_), .A2(\asqrt[52] ), .A3(new_n21497_), .A4(new_n21743_), .ZN(new_n22200_));
  AOI21_X1   g22007(.A1(new_n22192_), .A2(new_n21493_), .B(new_n1260_), .ZN(new_n22201_));
  NOR2_X1    g22008(.A1(new_n22200_), .A2(new_n22201_), .ZN(new_n22202_));
  NAND2_X1   g22009(.A1(new_n22202_), .A2(new_n1096_), .ZN(new_n22203_));
  AOI21_X1   g22010(.A1(new_n22199_), .A2(\asqrt[52] ), .B(new_n22203_), .ZN(new_n22204_));
  NOR2_X1    g22011(.A1(new_n22204_), .A2(new_n22198_), .ZN(new_n22205_));
  AOI22_X1   g22012(.A1(new_n22199_), .A2(\asqrt[52] ), .B1(new_n22197_), .B2(new_n22190_), .ZN(new_n22206_));
  NAND2_X1   g22013(.A1(new_n21509_), .A2(\asqrt[53] ), .ZN(new_n22207_));
  NOR4_X1    g22014(.A1(new_n21781_), .A2(\asqrt[53] ), .A3(new_n21504_), .A4(new_n21509_), .ZN(new_n22208_));
  XOR2_X1    g22015(.A1(new_n22208_), .A2(new_n22207_), .Z(new_n22209_));
  NAND2_X1   g22016(.A1(new_n22209_), .A2(new_n970_), .ZN(new_n22210_));
  INV_X1     g22017(.I(new_n22210_), .ZN(new_n22211_));
  OAI21_X1   g22018(.A1(new_n22206_), .A2(new_n1096_), .B(new_n22211_), .ZN(new_n22212_));
  NAND2_X1   g22019(.A1(new_n22212_), .A2(new_n22205_), .ZN(new_n22213_));
  OAI22_X1   g22020(.A1(new_n22206_), .A2(new_n1096_), .B1(new_n22204_), .B2(new_n22198_), .ZN(new_n22214_));
  NOR4_X1    g22021(.A1(new_n21781_), .A2(\asqrt[54] ), .A3(new_n21512_), .A4(new_n21750_), .ZN(new_n22215_));
  AOI21_X1   g22022(.A1(new_n22207_), .A2(new_n21508_), .B(new_n970_), .ZN(new_n22216_));
  NOR2_X1    g22023(.A1(new_n22215_), .A2(new_n22216_), .ZN(new_n22217_));
  NAND2_X1   g22024(.A1(new_n22217_), .A2(new_n825_), .ZN(new_n22218_));
  AOI21_X1   g22025(.A1(new_n22214_), .A2(\asqrt[54] ), .B(new_n22218_), .ZN(new_n22219_));
  NOR2_X1    g22026(.A1(new_n22219_), .A2(new_n22213_), .ZN(new_n22220_));
  AOI22_X1   g22027(.A1(new_n22214_), .A2(\asqrt[54] ), .B1(new_n22212_), .B2(new_n22205_), .ZN(new_n22221_));
  NAND2_X1   g22028(.A1(new_n21524_), .A2(\asqrt[55] ), .ZN(new_n22222_));
  NOR4_X1    g22029(.A1(new_n21781_), .A2(\asqrt[55] ), .A3(new_n21519_), .A4(new_n21524_), .ZN(new_n22223_));
  XOR2_X1    g22030(.A1(new_n22223_), .A2(new_n22222_), .Z(new_n22224_));
  NAND2_X1   g22031(.A1(new_n22224_), .A2(new_n724_), .ZN(new_n22225_));
  INV_X1     g22032(.I(new_n22225_), .ZN(new_n22226_));
  OAI21_X1   g22033(.A1(new_n22221_), .A2(new_n825_), .B(new_n22226_), .ZN(new_n22227_));
  NAND2_X1   g22034(.A1(new_n22227_), .A2(new_n22220_), .ZN(new_n22228_));
  OAI22_X1   g22035(.A1(new_n22221_), .A2(new_n825_), .B1(new_n22219_), .B2(new_n22213_), .ZN(new_n22229_));
  NOR4_X1    g22036(.A1(new_n21781_), .A2(\asqrt[56] ), .A3(new_n21526_), .A4(new_n21757_), .ZN(new_n22230_));
  AOI21_X1   g22037(.A1(new_n22222_), .A2(new_n21523_), .B(new_n724_), .ZN(new_n22231_));
  NOR2_X1    g22038(.A1(new_n22230_), .A2(new_n22231_), .ZN(new_n22232_));
  NAND2_X1   g22039(.A1(new_n22232_), .A2(new_n587_), .ZN(new_n22233_));
  AOI21_X1   g22040(.A1(new_n22229_), .A2(\asqrt[56] ), .B(new_n22233_), .ZN(new_n22234_));
  NOR2_X1    g22041(.A1(new_n22234_), .A2(new_n22228_), .ZN(new_n22235_));
  AOI22_X1   g22042(.A1(new_n22229_), .A2(\asqrt[56] ), .B1(new_n22227_), .B2(new_n22220_), .ZN(new_n22236_));
  NOR4_X1    g22043(.A1(new_n21781_), .A2(\asqrt[57] ), .A3(new_n21532_), .A4(new_n21537_), .ZN(new_n22237_));
  XOR2_X1    g22044(.A1(new_n22237_), .A2(new_n21563_), .Z(new_n22238_));
  INV_X1     g22045(.I(new_n22238_), .ZN(new_n22239_));
  NOR2_X1    g22046(.A1(new_n22239_), .A2(\asqrt[58] ), .ZN(new_n22240_));
  OAI21_X1   g22047(.A1(new_n22236_), .A2(new_n587_), .B(new_n22240_), .ZN(new_n22241_));
  NAND2_X1   g22048(.A1(new_n22241_), .A2(new_n22235_), .ZN(new_n22242_));
  OAI22_X1   g22049(.A1(new_n22236_), .A2(new_n587_), .B1(new_n22234_), .B2(new_n22228_), .ZN(new_n22243_));
  NOR4_X1    g22050(.A1(new_n21781_), .A2(\asqrt[58] ), .A3(new_n21539_), .A4(new_n21764_), .ZN(new_n22244_));
  XOR2_X1    g22051(.A1(new_n22244_), .A2(new_n21800_), .Z(new_n22245_));
  NAND2_X1   g22052(.A1(new_n22245_), .A2(new_n376_), .ZN(new_n22246_));
  AOI21_X1   g22053(.A1(new_n22243_), .A2(\asqrt[58] ), .B(new_n22246_), .ZN(new_n22247_));
  NOR2_X1    g22054(.A1(new_n22247_), .A2(new_n22242_), .ZN(new_n22248_));
  AOI22_X1   g22055(.A1(new_n22243_), .A2(\asqrt[58] ), .B1(new_n22241_), .B2(new_n22235_), .ZN(new_n22249_));
  NOR4_X1    g22056(.A1(new_n21781_), .A2(\asqrt[59] ), .A3(new_n21545_), .A4(new_n21550_), .ZN(new_n22250_));
  XOR2_X1    g22057(.A1(new_n22250_), .A2(new_n21565_), .Z(new_n22251_));
  INV_X1     g22058(.I(new_n22251_), .ZN(new_n22252_));
  NOR2_X1    g22059(.A1(new_n22252_), .A2(\asqrt[60] ), .ZN(new_n22253_));
  OAI21_X1   g22060(.A1(new_n22249_), .A2(new_n376_), .B(new_n22253_), .ZN(new_n22254_));
  NAND2_X1   g22061(.A1(new_n22254_), .A2(new_n22248_), .ZN(new_n22255_));
  OAI22_X1   g22062(.A1(new_n22249_), .A2(new_n376_), .B1(new_n22247_), .B2(new_n22242_), .ZN(new_n22256_));
  NAND2_X1   g22063(.A1(new_n22256_), .A2(\asqrt[60] ), .ZN(new_n22257_));
  NOR4_X1    g22064(.A1(new_n21781_), .A2(\asqrt[60] ), .A3(new_n21552_), .A4(new_n21771_), .ZN(new_n22258_));
  XOR2_X1    g22065(.A1(new_n22258_), .A2(new_n21802_), .Z(new_n22259_));
  NAND2_X1   g22066(.A1(new_n22259_), .A2(new_n229_), .ZN(new_n22260_));
  INV_X1     g22067(.I(new_n22260_), .ZN(new_n22261_));
  AOI21_X1   g22068(.A1(new_n22257_), .A2(new_n22261_), .B(new_n22255_), .ZN(new_n22262_));
  AOI22_X1   g22069(.A1(new_n22256_), .A2(\asqrt[60] ), .B1(new_n22254_), .B2(new_n22248_), .ZN(new_n22263_));
  INV_X1     g22070(.I(new_n21785_), .ZN(new_n22264_));
  NOR2_X1    g22071(.A1(new_n22264_), .A2(\asqrt[62] ), .ZN(new_n22265_));
  NOR3_X1    g22072(.A1(new_n22263_), .A2(new_n229_), .A3(new_n22265_), .ZN(new_n22266_));
  AOI21_X1   g22073(.A1(new_n22266_), .A2(new_n22262_), .B(new_n21786_), .ZN(new_n22267_));
  NOR3_X1    g22074(.A1(\asqrt[4] ), .A2(new_n21575_), .A3(new_n21780_), .ZN(new_n22268_));
  OAI21_X1   g22075(.A1(new_n22268_), .A2(new_n21778_), .B(new_n231_), .ZN(new_n22269_));
  INV_X1     g22076(.I(new_n22269_), .ZN(new_n22270_));
  AOI21_X1   g22077(.A1(new_n22267_), .A2(new_n22270_), .B(new_n21783_), .ZN(new_n22271_));
  AOI21_X1   g22078(.A1(new_n21081_), .A2(new_n21778_), .B(new_n21781_), .ZN(new_n22272_));
  XOR2_X1    g22079(.A1(new_n21778_), .A2(\asqrt[63] ), .Z(new_n22273_));
  NOR2_X1    g22080(.A1(new_n22272_), .A2(new_n22273_), .ZN(new_n22274_));
  INV_X1     g22081(.I(new_n22274_), .ZN(new_n22275_));
  INV_X1     g22082(.I(new_n21783_), .ZN(new_n22276_));
  NOR2_X1    g22083(.A1(new_n21858_), .A2(new_n21864_), .ZN(new_n22277_));
  NOR3_X1    g22084(.A1(new_n22277_), .A2(new_n21850_), .A3(new_n21887_), .ZN(new_n22278_));
  NAND2_X1   g22085(.A1(new_n21866_), .A2(new_n21870_), .ZN(new_n22279_));
  NAND2_X1   g22086(.A1(new_n22279_), .A2(new_n22278_), .ZN(new_n22280_));
  NAND2_X1   g22087(.A1(new_n21865_), .A2(new_n21866_), .ZN(new_n22281_));
  AOI21_X1   g22088(.A1(new_n22281_), .A2(\asqrt[11] ), .B(new_n21892_), .ZN(new_n22282_));
  NOR2_X1    g22089(.A1(new_n22282_), .A2(new_n22280_), .ZN(new_n22283_));
  AOI21_X1   g22090(.A1(new_n21865_), .A2(new_n21866_), .B(new_n17271_), .ZN(new_n22284_));
  OAI21_X1   g22091(.A1(new_n21871_), .A2(new_n22284_), .B(\asqrt[12] ), .ZN(new_n22285_));
  INV_X1     g22092(.I(new_n21901_), .ZN(new_n22286_));
  NAND2_X1   g22093(.A1(new_n22285_), .A2(new_n22286_), .ZN(new_n22287_));
  NAND2_X1   g22094(.A1(new_n22287_), .A2(new_n22283_), .ZN(new_n22288_));
  AOI22_X1   g22095(.A1(new_n22281_), .A2(\asqrt[11] ), .B1(new_n22279_), .B2(new_n22278_), .ZN(new_n22289_));
  OAI22_X1   g22096(.A1(new_n22289_), .A2(new_n16619_), .B1(new_n22282_), .B2(new_n22280_), .ZN(new_n22290_));
  AOI21_X1   g22097(.A1(new_n22290_), .A2(\asqrt[13] ), .B(new_n21908_), .ZN(new_n22291_));
  NOR2_X1    g22098(.A1(new_n22291_), .A2(new_n22288_), .ZN(new_n22292_));
  AOI22_X1   g22099(.A1(new_n22290_), .A2(\asqrt[13] ), .B1(new_n22287_), .B2(new_n22283_), .ZN(new_n22293_));
  INV_X1     g22100(.I(new_n21916_), .ZN(new_n22294_));
  OAI21_X1   g22101(.A1(new_n22293_), .A2(new_n15447_), .B(new_n22294_), .ZN(new_n22295_));
  NAND2_X1   g22102(.A1(new_n22295_), .A2(new_n22292_), .ZN(new_n22296_));
  OAI22_X1   g22103(.A1(new_n22293_), .A2(new_n15447_), .B1(new_n22291_), .B2(new_n22288_), .ZN(new_n22297_));
  AOI21_X1   g22104(.A1(new_n22297_), .A2(\asqrt[15] ), .B(new_n21923_), .ZN(new_n22298_));
  NOR2_X1    g22105(.A1(new_n22298_), .A2(new_n22296_), .ZN(new_n22299_));
  AOI22_X1   g22106(.A1(new_n22297_), .A2(\asqrt[15] ), .B1(new_n22295_), .B2(new_n22292_), .ZN(new_n22300_));
  INV_X1     g22107(.I(new_n21931_), .ZN(new_n22301_));
  OAI21_X1   g22108(.A1(new_n22300_), .A2(new_n14273_), .B(new_n22301_), .ZN(new_n22302_));
  NAND2_X1   g22109(.A1(new_n22302_), .A2(new_n22299_), .ZN(new_n22303_));
  OAI22_X1   g22110(.A1(new_n22300_), .A2(new_n14273_), .B1(new_n22298_), .B2(new_n22296_), .ZN(new_n22304_));
  AOI21_X1   g22111(.A1(new_n22304_), .A2(\asqrt[17] ), .B(new_n21938_), .ZN(new_n22305_));
  NOR2_X1    g22112(.A1(new_n22305_), .A2(new_n22303_), .ZN(new_n22306_));
  AOI22_X1   g22113(.A1(new_n22304_), .A2(\asqrt[17] ), .B1(new_n22302_), .B2(new_n22299_), .ZN(new_n22307_));
  INV_X1     g22114(.I(new_n21946_), .ZN(new_n22308_));
  OAI21_X1   g22115(.A1(new_n22307_), .A2(new_n13192_), .B(new_n22308_), .ZN(new_n22309_));
  NAND2_X1   g22116(.A1(new_n22309_), .A2(new_n22306_), .ZN(new_n22310_));
  OAI22_X1   g22117(.A1(new_n22307_), .A2(new_n13192_), .B1(new_n22305_), .B2(new_n22303_), .ZN(new_n22311_));
  AOI21_X1   g22118(.A1(new_n22311_), .A2(\asqrt[19] ), .B(new_n21953_), .ZN(new_n22312_));
  NOR2_X1    g22119(.A1(new_n22312_), .A2(new_n22310_), .ZN(new_n22313_));
  AOI22_X1   g22120(.A1(new_n22311_), .A2(\asqrt[19] ), .B1(new_n22309_), .B2(new_n22306_), .ZN(new_n22314_));
  INV_X1     g22121(.I(new_n21961_), .ZN(new_n22315_));
  OAI21_X1   g22122(.A1(new_n22314_), .A2(new_n12101_), .B(new_n22315_), .ZN(new_n22316_));
  NAND2_X1   g22123(.A1(new_n22316_), .A2(new_n22313_), .ZN(new_n22317_));
  OAI22_X1   g22124(.A1(new_n22314_), .A2(new_n12101_), .B1(new_n22312_), .B2(new_n22310_), .ZN(new_n22318_));
  AOI21_X1   g22125(.A1(new_n22318_), .A2(\asqrt[21] ), .B(new_n21968_), .ZN(new_n22319_));
  NOR2_X1    g22126(.A1(new_n22319_), .A2(new_n22317_), .ZN(new_n22320_));
  AOI22_X1   g22127(.A1(new_n22318_), .A2(\asqrt[21] ), .B1(new_n22316_), .B2(new_n22313_), .ZN(new_n22321_));
  INV_X1     g22128(.I(new_n21976_), .ZN(new_n22322_));
  OAI21_X1   g22129(.A1(new_n22321_), .A2(new_n11105_), .B(new_n22322_), .ZN(new_n22323_));
  NAND2_X1   g22130(.A1(new_n22323_), .A2(new_n22320_), .ZN(new_n22324_));
  OAI22_X1   g22131(.A1(new_n22321_), .A2(new_n11105_), .B1(new_n22319_), .B2(new_n22317_), .ZN(new_n22325_));
  AOI21_X1   g22132(.A1(new_n22325_), .A2(\asqrt[23] ), .B(new_n21983_), .ZN(new_n22326_));
  NOR2_X1    g22133(.A1(new_n22326_), .A2(new_n22324_), .ZN(new_n22327_));
  AOI22_X1   g22134(.A1(new_n22325_), .A2(\asqrt[23] ), .B1(new_n22323_), .B2(new_n22320_), .ZN(new_n22328_));
  INV_X1     g22135(.I(new_n21991_), .ZN(new_n22329_));
  OAI21_X1   g22136(.A1(new_n22328_), .A2(new_n10104_), .B(new_n22329_), .ZN(new_n22330_));
  NAND2_X1   g22137(.A1(new_n22330_), .A2(new_n22327_), .ZN(new_n22331_));
  OAI22_X1   g22138(.A1(new_n22328_), .A2(new_n10104_), .B1(new_n22326_), .B2(new_n22324_), .ZN(new_n22332_));
  AOI21_X1   g22139(.A1(new_n22332_), .A2(\asqrt[25] ), .B(new_n21998_), .ZN(new_n22333_));
  NOR2_X1    g22140(.A1(new_n22333_), .A2(new_n22331_), .ZN(new_n22334_));
  AOI22_X1   g22141(.A1(new_n22332_), .A2(\asqrt[25] ), .B1(new_n22330_), .B2(new_n22327_), .ZN(new_n22335_));
  INV_X1     g22142(.I(new_n22006_), .ZN(new_n22336_));
  OAI21_X1   g22143(.A1(new_n22335_), .A2(new_n9212_), .B(new_n22336_), .ZN(new_n22337_));
  NAND2_X1   g22144(.A1(new_n22337_), .A2(new_n22334_), .ZN(new_n22338_));
  OAI22_X1   g22145(.A1(new_n22335_), .A2(new_n9212_), .B1(new_n22333_), .B2(new_n22331_), .ZN(new_n22339_));
  AOI21_X1   g22146(.A1(new_n22339_), .A2(\asqrt[27] ), .B(new_n22013_), .ZN(new_n22340_));
  NOR2_X1    g22147(.A1(new_n22340_), .A2(new_n22338_), .ZN(new_n22341_));
  AOI22_X1   g22148(.A1(new_n22339_), .A2(\asqrt[27] ), .B1(new_n22337_), .B2(new_n22334_), .ZN(new_n22342_));
  INV_X1     g22149(.I(new_n22021_), .ZN(new_n22343_));
  OAI21_X1   g22150(.A1(new_n22342_), .A2(new_n8319_), .B(new_n22343_), .ZN(new_n22344_));
  NAND2_X1   g22151(.A1(new_n22344_), .A2(new_n22341_), .ZN(new_n22345_));
  OAI22_X1   g22152(.A1(new_n22342_), .A2(new_n8319_), .B1(new_n22340_), .B2(new_n22338_), .ZN(new_n22346_));
  AOI21_X1   g22153(.A1(new_n22346_), .A2(\asqrt[29] ), .B(new_n22028_), .ZN(new_n22347_));
  NOR2_X1    g22154(.A1(new_n22347_), .A2(new_n22345_), .ZN(new_n22348_));
  AOI22_X1   g22155(.A1(new_n22346_), .A2(\asqrt[29] ), .B1(new_n22344_), .B2(new_n22341_), .ZN(new_n22349_));
  INV_X1     g22156(.I(new_n22036_), .ZN(new_n22350_));
  OAI21_X1   g22157(.A1(new_n22349_), .A2(new_n7517_), .B(new_n22350_), .ZN(new_n22351_));
  NAND2_X1   g22158(.A1(new_n22351_), .A2(new_n22348_), .ZN(new_n22352_));
  OAI22_X1   g22159(.A1(new_n22349_), .A2(new_n7517_), .B1(new_n22347_), .B2(new_n22345_), .ZN(new_n22353_));
  AOI21_X1   g22160(.A1(new_n22353_), .A2(\asqrt[31] ), .B(new_n22043_), .ZN(new_n22354_));
  NOR2_X1    g22161(.A1(new_n22354_), .A2(new_n22352_), .ZN(new_n22355_));
  AOI22_X1   g22162(.A1(new_n22353_), .A2(\asqrt[31] ), .B1(new_n22351_), .B2(new_n22348_), .ZN(new_n22356_));
  INV_X1     g22163(.I(new_n22051_), .ZN(new_n22357_));
  OAI21_X1   g22164(.A1(new_n22356_), .A2(new_n6708_), .B(new_n22357_), .ZN(new_n22358_));
  NAND2_X1   g22165(.A1(new_n22358_), .A2(new_n22355_), .ZN(new_n22359_));
  OAI22_X1   g22166(.A1(new_n22356_), .A2(new_n6708_), .B1(new_n22354_), .B2(new_n22352_), .ZN(new_n22360_));
  AOI21_X1   g22167(.A1(new_n22360_), .A2(\asqrt[33] ), .B(new_n22058_), .ZN(new_n22361_));
  NOR2_X1    g22168(.A1(new_n22361_), .A2(new_n22359_), .ZN(new_n22362_));
  AOI22_X1   g22169(.A1(new_n22360_), .A2(\asqrt[33] ), .B1(new_n22358_), .B2(new_n22355_), .ZN(new_n22363_));
  INV_X1     g22170(.I(new_n22066_), .ZN(new_n22364_));
  OAI21_X1   g22171(.A1(new_n22363_), .A2(new_n5991_), .B(new_n22364_), .ZN(new_n22365_));
  NAND2_X1   g22172(.A1(new_n22365_), .A2(new_n22362_), .ZN(new_n22366_));
  OAI22_X1   g22173(.A1(new_n22363_), .A2(new_n5991_), .B1(new_n22361_), .B2(new_n22359_), .ZN(new_n22367_));
  AOI21_X1   g22174(.A1(new_n22367_), .A2(\asqrt[35] ), .B(new_n22073_), .ZN(new_n22368_));
  NOR2_X1    g22175(.A1(new_n22368_), .A2(new_n22366_), .ZN(new_n22369_));
  AOI22_X1   g22176(.A1(new_n22367_), .A2(\asqrt[35] ), .B1(new_n22365_), .B2(new_n22362_), .ZN(new_n22370_));
  INV_X1     g22177(.I(new_n22081_), .ZN(new_n22371_));
  OAI21_X1   g22178(.A1(new_n22370_), .A2(new_n5273_), .B(new_n22371_), .ZN(new_n22372_));
  NAND2_X1   g22179(.A1(new_n22372_), .A2(new_n22369_), .ZN(new_n22373_));
  OAI22_X1   g22180(.A1(new_n22370_), .A2(new_n5273_), .B1(new_n22368_), .B2(new_n22366_), .ZN(new_n22374_));
  INV_X1     g22181(.I(new_n22089_), .ZN(new_n22375_));
  AOI21_X1   g22182(.A1(new_n22374_), .A2(\asqrt[37] ), .B(new_n22375_), .ZN(new_n22376_));
  NOR2_X1    g22183(.A1(new_n22376_), .A2(new_n22373_), .ZN(new_n22377_));
  AOI22_X1   g22184(.A1(new_n22374_), .A2(\asqrt[37] ), .B1(new_n22372_), .B2(new_n22369_), .ZN(new_n22378_));
  INV_X1     g22185(.I(new_n22096_), .ZN(new_n22379_));
  OAI21_X1   g22186(.A1(new_n22378_), .A2(new_n4645_), .B(new_n22379_), .ZN(new_n22380_));
  NAND2_X1   g22187(.A1(new_n22380_), .A2(new_n22377_), .ZN(new_n22381_));
  OAI22_X1   g22188(.A1(new_n22378_), .A2(new_n4645_), .B1(new_n22376_), .B2(new_n22373_), .ZN(new_n22382_));
  INV_X1     g22189(.I(new_n22104_), .ZN(new_n22383_));
  AOI21_X1   g22190(.A1(new_n22382_), .A2(\asqrt[39] ), .B(new_n22383_), .ZN(new_n22384_));
  NOR2_X1    g22191(.A1(new_n22384_), .A2(new_n22381_), .ZN(new_n22385_));
  AOI22_X1   g22192(.A1(new_n22382_), .A2(\asqrt[39] ), .B1(new_n22380_), .B2(new_n22377_), .ZN(new_n22386_));
  INV_X1     g22193(.I(new_n22111_), .ZN(new_n22387_));
  OAI21_X1   g22194(.A1(new_n22386_), .A2(new_n4018_), .B(new_n22387_), .ZN(new_n22388_));
  NAND2_X1   g22195(.A1(new_n22388_), .A2(new_n22385_), .ZN(new_n22389_));
  OAI22_X1   g22196(.A1(new_n22386_), .A2(new_n4018_), .B1(new_n22384_), .B2(new_n22381_), .ZN(new_n22390_));
  INV_X1     g22197(.I(new_n22119_), .ZN(new_n22391_));
  AOI21_X1   g22198(.A1(new_n22390_), .A2(\asqrt[41] ), .B(new_n22391_), .ZN(new_n22392_));
  NOR2_X1    g22199(.A1(new_n22392_), .A2(new_n22389_), .ZN(new_n22393_));
  AOI22_X1   g22200(.A1(new_n22390_), .A2(\asqrt[41] ), .B1(new_n22388_), .B2(new_n22385_), .ZN(new_n22394_));
  INV_X1     g22201(.I(new_n22126_), .ZN(new_n22395_));
  OAI21_X1   g22202(.A1(new_n22394_), .A2(new_n3481_), .B(new_n22395_), .ZN(new_n22396_));
  NAND2_X1   g22203(.A1(new_n22396_), .A2(new_n22393_), .ZN(new_n22397_));
  OAI22_X1   g22204(.A1(new_n22394_), .A2(new_n3481_), .B1(new_n22392_), .B2(new_n22389_), .ZN(new_n22398_));
  AOI21_X1   g22205(.A1(new_n22398_), .A2(\asqrt[43] ), .B(new_n22133_), .ZN(new_n22399_));
  NOR2_X1    g22206(.A1(new_n22399_), .A2(new_n22397_), .ZN(new_n22400_));
  AOI22_X1   g22207(.A1(new_n22398_), .A2(\asqrt[43] ), .B1(new_n22396_), .B2(new_n22393_), .ZN(new_n22401_));
  OAI21_X1   g22208(.A1(new_n22401_), .A2(new_n2941_), .B(new_n22142_), .ZN(new_n22402_));
  NAND2_X1   g22209(.A1(new_n22402_), .A2(new_n22400_), .ZN(new_n22403_));
  OAI22_X1   g22210(.A1(new_n22401_), .A2(new_n2941_), .B1(new_n22399_), .B2(new_n22397_), .ZN(new_n22404_));
  AOI21_X1   g22211(.A1(new_n22404_), .A2(\asqrt[45] ), .B(new_n22150_), .ZN(new_n22405_));
  NOR2_X1    g22212(.A1(new_n22405_), .A2(new_n22403_), .ZN(new_n22406_));
  AOI22_X1   g22213(.A1(new_n22404_), .A2(\asqrt[45] ), .B1(new_n22402_), .B2(new_n22400_), .ZN(new_n22407_));
  INV_X1     g22214(.I(new_n22158_), .ZN(new_n22408_));
  OAI21_X1   g22215(.A1(new_n22407_), .A2(new_n2488_), .B(new_n22408_), .ZN(new_n22409_));
  NAND2_X1   g22216(.A1(new_n22409_), .A2(new_n22406_), .ZN(new_n22410_));
  OAI22_X1   g22217(.A1(new_n22407_), .A2(new_n2488_), .B1(new_n22405_), .B2(new_n22403_), .ZN(new_n22411_));
  INV_X1     g22218(.I(new_n22166_), .ZN(new_n22412_));
  AOI21_X1   g22219(.A1(new_n22411_), .A2(\asqrt[47] ), .B(new_n22412_), .ZN(new_n22413_));
  NOR2_X1    g22220(.A1(new_n22413_), .A2(new_n22410_), .ZN(new_n22414_));
  AOI22_X1   g22221(.A1(new_n22411_), .A2(\asqrt[47] ), .B1(new_n22409_), .B2(new_n22406_), .ZN(new_n22415_));
  INV_X1     g22222(.I(new_n22173_), .ZN(new_n22416_));
  OAI21_X1   g22223(.A1(new_n22415_), .A2(new_n2046_), .B(new_n22416_), .ZN(new_n22417_));
  NAND2_X1   g22224(.A1(new_n22417_), .A2(new_n22414_), .ZN(new_n22418_));
  OAI22_X1   g22225(.A1(new_n22415_), .A2(new_n2046_), .B1(new_n22413_), .B2(new_n22410_), .ZN(new_n22419_));
  INV_X1     g22226(.I(new_n22181_), .ZN(new_n22420_));
  AOI21_X1   g22227(.A1(new_n22419_), .A2(\asqrt[49] ), .B(new_n22420_), .ZN(new_n22421_));
  NOR2_X1    g22228(.A1(new_n22421_), .A2(new_n22418_), .ZN(new_n22422_));
  AOI22_X1   g22229(.A1(new_n22419_), .A2(\asqrt[49] ), .B1(new_n22417_), .B2(new_n22414_), .ZN(new_n22423_));
  INV_X1     g22230(.I(new_n22188_), .ZN(new_n22424_));
  OAI21_X1   g22231(.A1(new_n22423_), .A2(new_n1595_), .B(new_n22424_), .ZN(new_n22425_));
  NAND2_X1   g22232(.A1(new_n22425_), .A2(new_n22422_), .ZN(new_n22426_));
  OAI22_X1   g22233(.A1(new_n22423_), .A2(new_n1595_), .B1(new_n22421_), .B2(new_n22418_), .ZN(new_n22427_));
  AOI21_X1   g22234(.A1(new_n22427_), .A2(\asqrt[51] ), .B(new_n22195_), .ZN(new_n22428_));
  NOR2_X1    g22235(.A1(new_n22428_), .A2(new_n22426_), .ZN(new_n22429_));
  AOI22_X1   g22236(.A1(new_n22427_), .A2(\asqrt[51] ), .B1(new_n22425_), .B2(new_n22422_), .ZN(new_n22430_));
  INV_X1     g22237(.I(new_n22203_), .ZN(new_n22431_));
  OAI21_X1   g22238(.A1(new_n22430_), .A2(new_n1260_), .B(new_n22431_), .ZN(new_n22432_));
  NAND2_X1   g22239(.A1(new_n22432_), .A2(new_n22429_), .ZN(new_n22433_));
  OAI22_X1   g22240(.A1(new_n22430_), .A2(new_n1260_), .B1(new_n22428_), .B2(new_n22426_), .ZN(new_n22434_));
  AOI21_X1   g22241(.A1(new_n22434_), .A2(\asqrt[53] ), .B(new_n22210_), .ZN(new_n22435_));
  NOR2_X1    g22242(.A1(new_n22435_), .A2(new_n22433_), .ZN(new_n22436_));
  AOI22_X1   g22243(.A1(new_n22434_), .A2(\asqrt[53] ), .B1(new_n22432_), .B2(new_n22429_), .ZN(new_n22437_));
  INV_X1     g22244(.I(new_n22218_), .ZN(new_n22438_));
  OAI21_X1   g22245(.A1(new_n22437_), .A2(new_n970_), .B(new_n22438_), .ZN(new_n22439_));
  NAND2_X1   g22246(.A1(new_n22439_), .A2(new_n22436_), .ZN(new_n22440_));
  OAI22_X1   g22247(.A1(new_n22437_), .A2(new_n970_), .B1(new_n22435_), .B2(new_n22433_), .ZN(new_n22441_));
  AOI21_X1   g22248(.A1(new_n22441_), .A2(\asqrt[55] ), .B(new_n22225_), .ZN(new_n22442_));
  NOR2_X1    g22249(.A1(new_n22442_), .A2(new_n22440_), .ZN(new_n22443_));
  AOI22_X1   g22250(.A1(new_n22441_), .A2(\asqrt[55] ), .B1(new_n22439_), .B2(new_n22436_), .ZN(new_n22444_));
  INV_X1     g22251(.I(new_n22233_), .ZN(new_n22445_));
  OAI21_X1   g22252(.A1(new_n22444_), .A2(new_n724_), .B(new_n22445_), .ZN(new_n22446_));
  NAND2_X1   g22253(.A1(new_n22446_), .A2(new_n22443_), .ZN(new_n22447_));
  OAI22_X1   g22254(.A1(new_n22444_), .A2(new_n724_), .B1(new_n22442_), .B2(new_n22440_), .ZN(new_n22448_));
  INV_X1     g22255(.I(new_n22240_), .ZN(new_n22449_));
  AOI21_X1   g22256(.A1(new_n22448_), .A2(\asqrt[57] ), .B(new_n22449_), .ZN(new_n22450_));
  NOR2_X1    g22257(.A1(new_n22450_), .A2(new_n22447_), .ZN(new_n22451_));
  AOI22_X1   g22258(.A1(new_n22448_), .A2(\asqrt[57] ), .B1(new_n22446_), .B2(new_n22443_), .ZN(new_n22452_));
  INV_X1     g22259(.I(new_n22246_), .ZN(new_n22453_));
  OAI21_X1   g22260(.A1(new_n22452_), .A2(new_n504_), .B(new_n22453_), .ZN(new_n22454_));
  NAND2_X1   g22261(.A1(new_n22454_), .A2(new_n22451_), .ZN(new_n22455_));
  OAI22_X1   g22262(.A1(new_n22452_), .A2(new_n504_), .B1(new_n22450_), .B2(new_n22447_), .ZN(new_n22456_));
  INV_X1     g22263(.I(new_n22253_), .ZN(new_n22457_));
  AOI21_X1   g22264(.A1(new_n22456_), .A2(\asqrt[59] ), .B(new_n22457_), .ZN(new_n22458_));
  NOR2_X1    g22265(.A1(new_n22458_), .A2(new_n22455_), .ZN(new_n22459_));
  AOI22_X1   g22266(.A1(new_n22456_), .A2(\asqrt[59] ), .B1(new_n22454_), .B2(new_n22451_), .ZN(new_n22460_));
  OAI21_X1   g22267(.A1(new_n22460_), .A2(new_n275_), .B(new_n22261_), .ZN(new_n22461_));
  OAI22_X1   g22268(.A1(new_n22460_), .A2(new_n275_), .B1(new_n22458_), .B2(new_n22455_), .ZN(new_n22462_));
  AOI22_X1   g22269(.A1(new_n22462_), .A2(\asqrt[61] ), .B1(new_n22461_), .B2(new_n22459_), .ZN(new_n22463_));
  NAND4_X1   g22270(.A1(new_n22463_), .A2(new_n196_), .A3(new_n22276_), .A4(new_n22264_), .ZN(new_n22464_));
  NAND2_X1   g22271(.A1(new_n22464_), .A2(new_n22275_), .ZN(new_n22465_));
  OAI21_X1   g22272(.A1(new_n22465_), .A2(new_n22271_), .B(\a[7] ), .ZN(new_n22466_));
  NOR2_X1    g22273(.A1(new_n21588_), .A2(\a[6] ), .ZN(new_n22467_));
  INV_X1     g22274(.I(new_n22467_), .ZN(new_n22468_));
  AOI21_X1   g22275(.A1(new_n22466_), .A2(new_n22468_), .B(new_n21589_), .ZN(new_n22469_));
  INV_X1     g22276(.I(\a[6] ), .ZN(new_n22470_));
  INV_X1     g22277(.I(new_n21786_), .ZN(new_n22471_));
  NAND2_X1   g22278(.A1(new_n22461_), .A2(new_n22459_), .ZN(new_n22472_));
  INV_X1     g22279(.I(new_n22265_), .ZN(new_n22473_));
  NAND3_X1   g22280(.A1(new_n22462_), .A2(\asqrt[61] ), .A3(new_n22473_), .ZN(new_n22474_));
  OAI21_X1   g22281(.A1(new_n22474_), .A2(new_n22472_), .B(new_n22471_), .ZN(new_n22475_));
  OAI21_X1   g22282(.A1(new_n22475_), .A2(new_n22269_), .B(new_n22276_), .ZN(new_n22476_));
  OAI21_X1   g22283(.A1(new_n22463_), .A2(new_n196_), .B(new_n21783_), .ZN(new_n22477_));
  NOR2_X1    g22284(.A1(new_n22263_), .A2(new_n229_), .ZN(new_n22478_));
  NOR4_X1    g22285(.A1(new_n22478_), .A2(new_n22262_), .A3(\asqrt[62] ), .A4(new_n21785_), .ZN(new_n22479_));
  AOI21_X1   g22286(.A1(new_n22477_), .A2(new_n22479_), .B(new_n22274_), .ZN(new_n22480_));
  AOI21_X1   g22287(.A1(new_n22480_), .A2(new_n22476_), .B(new_n217_), .ZN(new_n22481_));
  NOR3_X1    g22288(.A1(new_n22481_), .A2(new_n22470_), .A3(new_n21588_), .ZN(new_n22482_));
  NAND3_X1   g22289(.A1(new_n22476_), .A2(new_n22275_), .A3(new_n22464_), .ZN(\asqrt[3] ));
  NAND3_X1   g22290(.A1(\asqrt[3] ), .A2(\a[6] ), .A3(\asqrt[4] ), .ZN(new_n22484_));
  NAND4_X1   g22291(.A1(new_n22480_), .A2(new_n22470_), .A3(new_n22476_), .A4(\asqrt[4] ), .ZN(new_n22485_));
  AOI21_X1   g22292(.A1(new_n22484_), .A2(new_n22485_), .B(new_n21585_), .ZN(new_n22486_));
  NOR2_X1    g22293(.A1(new_n22275_), .A2(new_n21781_), .ZN(new_n22487_));
  INV_X1     g22294(.I(new_n22487_), .ZN(new_n22488_));
  NOR2_X1    g22295(.A1(new_n22464_), .A2(new_n22488_), .ZN(new_n22489_));
  NAND4_X1   g22296(.A1(new_n22480_), .A2(\a[8] ), .A3(new_n22476_), .A4(new_n21788_), .ZN(new_n22490_));
  AOI21_X1   g22297(.A1(new_n22489_), .A2(new_n22271_), .B(\a[8] ), .ZN(new_n22491_));
  OAI21_X1   g22298(.A1(new_n22491_), .A2(new_n21789_), .B(\asqrt[3] ), .ZN(new_n22492_));
  NAND3_X1   g22299(.A1(new_n22492_), .A2(new_n21079_), .A3(new_n22490_), .ZN(new_n22493_));
  OAI22_X1   g22300(.A1(new_n22493_), .A2(new_n22486_), .B1(new_n22469_), .B2(new_n22482_), .ZN(new_n22494_));
  NOR2_X1    g22301(.A1(new_n22482_), .A2(new_n22469_), .ZN(new_n22495_));
  NOR2_X1    g22302(.A1(new_n22465_), .A2(new_n22271_), .ZN(new_n22496_));
  NAND2_X1   g22303(.A1(\asqrt[4] ), .A2(\a[6] ), .ZN(new_n22497_));
  AOI21_X1   g22304(.A1(new_n22496_), .A2(\asqrt[4] ), .B(new_n22497_), .ZN(new_n22498_));
  NOR4_X1    g22305(.A1(new_n22465_), .A2(new_n22271_), .A3(\a[6] ), .A4(new_n21781_), .ZN(new_n22499_));
  OAI21_X1   g22306(.A1(new_n22498_), .A2(new_n22499_), .B(new_n21584_), .ZN(new_n22500_));
  AOI21_X1   g22307(.A1(new_n22495_), .A2(new_n22500_), .B(new_n21079_), .ZN(new_n22501_));
  OAI21_X1   g22308(.A1(new_n21781_), .A2(\a[8] ), .B(new_n21787_), .ZN(new_n22502_));
  NAND2_X1   g22309(.A1(new_n21808_), .A2(new_n21798_), .ZN(new_n22503_));
  NAND2_X1   g22310(.A1(new_n22503_), .A2(new_n22502_), .ZN(new_n22504_));
  NAND2_X1   g22311(.A1(new_n21816_), .A2(new_n21791_), .ZN(new_n22505_));
  AOI21_X1   g22312(.A1(new_n22505_), .A2(new_n21798_), .B(new_n21781_), .ZN(new_n22506_));
  AOI21_X1   g22313(.A1(\asqrt[3] ), .A2(new_n22506_), .B(new_n22504_), .ZN(new_n22507_));
  INV_X1     g22314(.I(new_n22507_), .ZN(new_n22508_));
  AND2_X2    g22315(.A1(new_n22506_), .A2(new_n22504_), .Z(new_n22509_));
  NAND2_X1   g22316(.A1(\asqrt[3] ), .A2(new_n22509_), .ZN(new_n22510_));
  NAND3_X1   g22317(.A1(new_n22508_), .A2(new_n20455_), .A3(new_n22510_), .ZN(new_n22511_));
  NOR2_X1    g22318(.A1(new_n22501_), .A2(new_n22511_), .ZN(new_n22512_));
  NOR2_X1    g22319(.A1(new_n22512_), .A2(new_n22494_), .ZN(new_n22513_));
  INV_X1     g22320(.I(new_n22490_), .ZN(new_n22514_));
  NAND3_X1   g22321(.A1(new_n22477_), .A2(new_n22479_), .A3(new_n22487_), .ZN(new_n22515_));
  OAI21_X1   g22322(.A1(new_n22515_), .A2(new_n22476_), .B(new_n21798_), .ZN(new_n22516_));
  AOI21_X1   g22323(.A1(new_n22516_), .A2(new_n21788_), .B(new_n22496_), .ZN(new_n22517_));
  NOR3_X1    g22324(.A1(new_n22517_), .A2(\asqrt[5] ), .A3(new_n22514_), .ZN(new_n22518_));
  AOI21_X1   g22325(.A1(new_n22518_), .A2(new_n22500_), .B(new_n22495_), .ZN(new_n22519_));
  OAI21_X1   g22326(.A1(new_n22519_), .A2(new_n22501_), .B(\asqrt[6] ), .ZN(new_n22520_));
  OAI21_X1   g22327(.A1(new_n21877_), .A2(new_n21876_), .B(new_n20455_), .ZN(new_n22521_));
  NOR2_X1    g22328(.A1(new_n21880_), .A2(new_n22521_), .ZN(new_n22522_));
  NAND2_X1   g22329(.A1(\asqrt[3] ), .A2(new_n22522_), .ZN(new_n22523_));
  XOR2_X1    g22330(.A1(new_n22523_), .A2(new_n21830_), .Z(new_n22524_));
  NOR2_X1    g22331(.A1(new_n22524_), .A2(\asqrt[7] ), .ZN(new_n22525_));
  NAND2_X1   g22332(.A1(new_n22520_), .A2(new_n22525_), .ZN(new_n22526_));
  NAND2_X1   g22333(.A1(new_n22526_), .A2(new_n22513_), .ZN(new_n22527_));
  NOR2_X1    g22334(.A1(new_n22519_), .A2(new_n22501_), .ZN(new_n22528_));
  OAI22_X1   g22335(.A1(new_n22528_), .A2(new_n20455_), .B1(new_n22512_), .B2(new_n22494_), .ZN(new_n22529_));
  NOR2_X1    g22336(.A1(new_n21838_), .A2(\asqrt[7] ), .ZN(new_n22530_));
  NAND3_X1   g22337(.A1(\asqrt[3] ), .A2(new_n21881_), .A3(new_n22530_), .ZN(new_n22531_));
  XOR2_X1    g22338(.A1(new_n22531_), .A2(new_n21842_), .Z(new_n22532_));
  NAND2_X1   g22339(.A1(new_n22532_), .A2(new_n19100_), .ZN(new_n22533_));
  AOI21_X1   g22340(.A1(new_n22529_), .A2(\asqrt[7] ), .B(new_n22533_), .ZN(new_n22534_));
  NOR2_X1    g22341(.A1(new_n22534_), .A2(new_n22527_), .ZN(new_n22535_));
  OAI21_X1   g22342(.A1(new_n22501_), .A2(new_n22511_), .B(new_n22519_), .ZN(new_n22536_));
  AOI21_X1   g22343(.A1(new_n22520_), .A2(new_n22525_), .B(new_n22536_), .ZN(new_n22537_));
  AOI21_X1   g22344(.A1(new_n22536_), .A2(new_n22520_), .B(new_n19782_), .ZN(new_n22538_));
  OAI21_X1   g22345(.A1(new_n22537_), .A2(new_n22538_), .B(\asqrt[8] ), .ZN(new_n22539_));
  NOR2_X1    g22346(.A1(new_n21841_), .A2(new_n21842_), .ZN(new_n22540_));
  NAND4_X1   g22347(.A1(\asqrt[3] ), .A2(new_n19100_), .A3(new_n21847_), .A4(new_n22540_), .ZN(new_n22541_));
  XNOR2_X1   g22348(.A1(new_n22541_), .A2(new_n21851_), .ZN(new_n22542_));
  NAND2_X1   g22349(.A1(new_n22542_), .A2(new_n18495_), .ZN(new_n22543_));
  INV_X1     g22350(.I(new_n22543_), .ZN(new_n22544_));
  NAND2_X1   g22351(.A1(new_n22539_), .A2(new_n22544_), .ZN(new_n22545_));
  NAND2_X1   g22352(.A1(new_n22545_), .A2(new_n22535_), .ZN(new_n22546_));
  AOI22_X1   g22353(.A1(new_n22529_), .A2(\asqrt[7] ), .B1(new_n22526_), .B2(new_n22513_), .ZN(new_n22547_));
  OAI22_X1   g22354(.A1(new_n22547_), .A2(new_n19100_), .B1(new_n22534_), .B2(new_n22527_), .ZN(new_n22548_));
  INV_X1     g22355(.I(new_n21885_), .ZN(new_n22549_));
  NOR4_X1    g22356(.A1(new_n22496_), .A2(\asqrt[9] ), .A3(new_n21854_), .A4(new_n22549_), .ZN(new_n22550_));
  XNOR2_X1   g22357(.A1(new_n22550_), .A2(new_n21858_), .ZN(new_n22551_));
  NAND2_X1   g22358(.A1(new_n22551_), .A2(new_n17893_), .ZN(new_n22552_));
  AOI21_X1   g22359(.A1(new_n22548_), .A2(\asqrt[9] ), .B(new_n22552_), .ZN(new_n22553_));
  NOR2_X1    g22360(.A1(new_n22553_), .A2(new_n22546_), .ZN(new_n22554_));
  AOI22_X1   g22361(.A1(new_n22548_), .A2(\asqrt[9] ), .B1(new_n22545_), .B2(new_n22535_), .ZN(new_n22555_));
  NOR4_X1    g22362(.A1(new_n22496_), .A2(\asqrt[10] ), .A3(new_n21861_), .A4(new_n21888_), .ZN(new_n22556_));
  XOR2_X1    g22363(.A1(new_n22556_), .A2(new_n21866_), .Z(new_n22557_));
  NAND2_X1   g22364(.A1(new_n22557_), .A2(new_n17271_), .ZN(new_n22558_));
  INV_X1     g22365(.I(new_n22558_), .ZN(new_n22559_));
  OAI21_X1   g22366(.A1(new_n22555_), .A2(new_n17893_), .B(new_n22559_), .ZN(new_n22560_));
  NAND2_X1   g22367(.A1(new_n22560_), .A2(new_n22554_), .ZN(new_n22561_));
  OAI22_X1   g22368(.A1(new_n22555_), .A2(new_n17893_), .B1(new_n22553_), .B2(new_n22546_), .ZN(new_n22562_));
  NOR4_X1    g22369(.A1(new_n22496_), .A2(\asqrt[11] ), .A3(new_n21868_), .A4(new_n22281_), .ZN(new_n22563_));
  XNOR2_X1   g22370(.A1(new_n22563_), .A2(new_n22284_), .ZN(new_n22564_));
  NAND2_X1   g22371(.A1(new_n22564_), .A2(new_n16619_), .ZN(new_n22565_));
  AOI21_X1   g22372(.A1(new_n22562_), .A2(\asqrt[11] ), .B(new_n22565_), .ZN(new_n22566_));
  NOR2_X1    g22373(.A1(new_n22566_), .A2(new_n22561_), .ZN(new_n22567_));
  AOI22_X1   g22374(.A1(new_n22562_), .A2(\asqrt[11] ), .B1(new_n22560_), .B2(new_n22554_), .ZN(new_n22568_));
  NOR4_X1    g22375(.A1(new_n22496_), .A2(\asqrt[12] ), .A3(new_n21891_), .A4(new_n21897_), .ZN(new_n22569_));
  XOR2_X1    g22376(.A1(new_n22569_), .A2(new_n22285_), .Z(new_n22570_));
  NAND2_X1   g22377(.A1(new_n22570_), .A2(new_n16060_), .ZN(new_n22571_));
  INV_X1     g22378(.I(new_n22571_), .ZN(new_n22572_));
  OAI21_X1   g22379(.A1(new_n22568_), .A2(new_n16619_), .B(new_n22572_), .ZN(new_n22573_));
  NAND2_X1   g22380(.A1(new_n22573_), .A2(new_n22567_), .ZN(new_n22574_));
  OAI22_X1   g22381(.A1(new_n22568_), .A2(new_n16619_), .B1(new_n22566_), .B2(new_n22561_), .ZN(new_n22575_));
  NOR4_X1    g22382(.A1(new_n22496_), .A2(\asqrt[13] ), .A3(new_n21900_), .A4(new_n22290_), .ZN(new_n22576_));
  AOI21_X1   g22383(.A1(new_n21895_), .A2(new_n22285_), .B(new_n16060_), .ZN(new_n22577_));
  NOR2_X1    g22384(.A1(new_n22576_), .A2(new_n22577_), .ZN(new_n22578_));
  NAND2_X1   g22385(.A1(new_n22578_), .A2(new_n15447_), .ZN(new_n22579_));
  AOI21_X1   g22386(.A1(new_n22575_), .A2(\asqrt[13] ), .B(new_n22579_), .ZN(new_n22580_));
  NOR2_X1    g22387(.A1(new_n22580_), .A2(new_n22574_), .ZN(new_n22581_));
  AOI22_X1   g22388(.A1(new_n22575_), .A2(\asqrt[13] ), .B1(new_n22573_), .B2(new_n22567_), .ZN(new_n22582_));
  NAND2_X1   g22389(.A1(new_n21912_), .A2(\asqrt[14] ), .ZN(new_n22583_));
  NOR4_X1    g22390(.A1(new_n22496_), .A2(\asqrt[14] ), .A3(new_n21907_), .A4(new_n21912_), .ZN(new_n22584_));
  XOR2_X1    g22391(.A1(new_n22584_), .A2(new_n22583_), .Z(new_n22585_));
  NAND2_X1   g22392(.A1(new_n22585_), .A2(new_n14871_), .ZN(new_n22586_));
  INV_X1     g22393(.I(new_n22586_), .ZN(new_n22587_));
  OAI21_X1   g22394(.A1(new_n22582_), .A2(new_n15447_), .B(new_n22587_), .ZN(new_n22588_));
  NAND2_X1   g22395(.A1(new_n22588_), .A2(new_n22581_), .ZN(new_n22589_));
  OAI22_X1   g22396(.A1(new_n22582_), .A2(new_n15447_), .B1(new_n22580_), .B2(new_n22574_), .ZN(new_n22590_));
  NOR4_X1    g22397(.A1(new_n22496_), .A2(\asqrt[15] ), .A3(new_n21915_), .A4(new_n22297_), .ZN(new_n22591_));
  AOI21_X1   g22398(.A1(new_n22583_), .A2(new_n21911_), .B(new_n14871_), .ZN(new_n22592_));
  NOR2_X1    g22399(.A1(new_n22591_), .A2(new_n22592_), .ZN(new_n22593_));
  NAND2_X1   g22400(.A1(new_n22593_), .A2(new_n14273_), .ZN(new_n22594_));
  AOI21_X1   g22401(.A1(new_n22590_), .A2(\asqrt[15] ), .B(new_n22594_), .ZN(new_n22595_));
  NOR2_X1    g22402(.A1(new_n22595_), .A2(new_n22589_), .ZN(new_n22596_));
  AOI22_X1   g22403(.A1(new_n22590_), .A2(\asqrt[15] ), .B1(new_n22588_), .B2(new_n22581_), .ZN(new_n22597_));
  NAND2_X1   g22404(.A1(new_n21927_), .A2(\asqrt[16] ), .ZN(new_n22598_));
  NOR4_X1    g22405(.A1(new_n22496_), .A2(\asqrt[16] ), .A3(new_n21922_), .A4(new_n21927_), .ZN(new_n22599_));
  XOR2_X1    g22406(.A1(new_n22599_), .A2(new_n22598_), .Z(new_n22600_));
  NAND2_X1   g22407(.A1(new_n22600_), .A2(new_n13760_), .ZN(new_n22601_));
  INV_X1     g22408(.I(new_n22601_), .ZN(new_n22602_));
  OAI21_X1   g22409(.A1(new_n22597_), .A2(new_n14273_), .B(new_n22602_), .ZN(new_n22603_));
  NAND2_X1   g22410(.A1(new_n22603_), .A2(new_n22596_), .ZN(new_n22604_));
  OAI22_X1   g22411(.A1(new_n22597_), .A2(new_n14273_), .B1(new_n22595_), .B2(new_n22589_), .ZN(new_n22605_));
  NOR4_X1    g22412(.A1(new_n22496_), .A2(\asqrt[17] ), .A3(new_n21930_), .A4(new_n22304_), .ZN(new_n22606_));
  AOI21_X1   g22413(.A1(new_n22598_), .A2(new_n21926_), .B(new_n13760_), .ZN(new_n22607_));
  NOR2_X1    g22414(.A1(new_n22606_), .A2(new_n22607_), .ZN(new_n22608_));
  NAND2_X1   g22415(.A1(new_n22608_), .A2(new_n13192_), .ZN(new_n22609_));
  AOI21_X1   g22416(.A1(new_n22605_), .A2(\asqrt[17] ), .B(new_n22609_), .ZN(new_n22610_));
  NOR2_X1    g22417(.A1(new_n22610_), .A2(new_n22604_), .ZN(new_n22611_));
  AOI22_X1   g22418(.A1(new_n22605_), .A2(\asqrt[17] ), .B1(new_n22603_), .B2(new_n22596_), .ZN(new_n22612_));
  NAND2_X1   g22419(.A1(new_n21942_), .A2(\asqrt[18] ), .ZN(new_n22613_));
  NOR4_X1    g22420(.A1(new_n22496_), .A2(\asqrt[18] ), .A3(new_n21937_), .A4(new_n21942_), .ZN(new_n22614_));
  XOR2_X1    g22421(.A1(new_n22614_), .A2(new_n22613_), .Z(new_n22615_));
  NAND2_X1   g22422(.A1(new_n22615_), .A2(new_n12657_), .ZN(new_n22616_));
  INV_X1     g22423(.I(new_n22616_), .ZN(new_n22617_));
  OAI21_X1   g22424(.A1(new_n22612_), .A2(new_n13192_), .B(new_n22617_), .ZN(new_n22618_));
  NAND2_X1   g22425(.A1(new_n22618_), .A2(new_n22611_), .ZN(new_n22619_));
  OAI22_X1   g22426(.A1(new_n22612_), .A2(new_n13192_), .B1(new_n22610_), .B2(new_n22604_), .ZN(new_n22620_));
  NOR4_X1    g22427(.A1(new_n22496_), .A2(\asqrt[19] ), .A3(new_n21945_), .A4(new_n22311_), .ZN(new_n22621_));
  AOI21_X1   g22428(.A1(new_n22613_), .A2(new_n21941_), .B(new_n12657_), .ZN(new_n22622_));
  NOR2_X1    g22429(.A1(new_n22621_), .A2(new_n22622_), .ZN(new_n22623_));
  NAND2_X1   g22430(.A1(new_n22623_), .A2(new_n12101_), .ZN(new_n22624_));
  AOI21_X1   g22431(.A1(new_n22620_), .A2(\asqrt[19] ), .B(new_n22624_), .ZN(new_n22625_));
  NOR2_X1    g22432(.A1(new_n22625_), .A2(new_n22619_), .ZN(new_n22626_));
  AOI22_X1   g22433(.A1(new_n22620_), .A2(\asqrt[19] ), .B1(new_n22618_), .B2(new_n22611_), .ZN(new_n22627_));
  NAND2_X1   g22434(.A1(new_n21957_), .A2(\asqrt[20] ), .ZN(new_n22628_));
  NOR4_X1    g22435(.A1(new_n22496_), .A2(\asqrt[20] ), .A3(new_n21952_), .A4(new_n21957_), .ZN(new_n22629_));
  XOR2_X1    g22436(.A1(new_n22629_), .A2(new_n22628_), .Z(new_n22630_));
  NAND2_X1   g22437(.A1(new_n22630_), .A2(new_n11631_), .ZN(new_n22631_));
  INV_X1     g22438(.I(new_n22631_), .ZN(new_n22632_));
  OAI21_X1   g22439(.A1(new_n22627_), .A2(new_n12101_), .B(new_n22632_), .ZN(new_n22633_));
  NAND2_X1   g22440(.A1(new_n22633_), .A2(new_n22626_), .ZN(new_n22634_));
  OAI22_X1   g22441(.A1(new_n22627_), .A2(new_n12101_), .B1(new_n22625_), .B2(new_n22619_), .ZN(new_n22635_));
  NOR4_X1    g22442(.A1(new_n22496_), .A2(\asqrt[21] ), .A3(new_n21960_), .A4(new_n22318_), .ZN(new_n22636_));
  AOI21_X1   g22443(.A1(new_n22628_), .A2(new_n21956_), .B(new_n11631_), .ZN(new_n22637_));
  NOR2_X1    g22444(.A1(new_n22636_), .A2(new_n22637_), .ZN(new_n22638_));
  NAND2_X1   g22445(.A1(new_n22638_), .A2(new_n11105_), .ZN(new_n22639_));
  AOI21_X1   g22446(.A1(new_n22635_), .A2(\asqrt[21] ), .B(new_n22639_), .ZN(new_n22640_));
  NOR2_X1    g22447(.A1(new_n22640_), .A2(new_n22634_), .ZN(new_n22641_));
  AOI22_X1   g22448(.A1(new_n22635_), .A2(\asqrt[21] ), .B1(new_n22633_), .B2(new_n22626_), .ZN(new_n22642_));
  NAND2_X1   g22449(.A1(new_n21972_), .A2(\asqrt[22] ), .ZN(new_n22643_));
  NOR4_X1    g22450(.A1(new_n22496_), .A2(\asqrt[22] ), .A3(new_n21967_), .A4(new_n21972_), .ZN(new_n22644_));
  XOR2_X1    g22451(.A1(new_n22644_), .A2(new_n22643_), .Z(new_n22645_));
  NAND2_X1   g22452(.A1(new_n22645_), .A2(new_n10614_), .ZN(new_n22646_));
  INV_X1     g22453(.I(new_n22646_), .ZN(new_n22647_));
  OAI21_X1   g22454(.A1(new_n22642_), .A2(new_n11105_), .B(new_n22647_), .ZN(new_n22648_));
  NAND2_X1   g22455(.A1(new_n22648_), .A2(new_n22641_), .ZN(new_n22649_));
  OAI22_X1   g22456(.A1(new_n22642_), .A2(new_n11105_), .B1(new_n22640_), .B2(new_n22634_), .ZN(new_n22650_));
  NOR4_X1    g22457(.A1(new_n22496_), .A2(\asqrt[23] ), .A3(new_n21975_), .A4(new_n22325_), .ZN(new_n22651_));
  AOI21_X1   g22458(.A1(new_n22643_), .A2(new_n21971_), .B(new_n10614_), .ZN(new_n22652_));
  NOR2_X1    g22459(.A1(new_n22651_), .A2(new_n22652_), .ZN(new_n22653_));
  NAND2_X1   g22460(.A1(new_n22653_), .A2(new_n10104_), .ZN(new_n22654_));
  AOI21_X1   g22461(.A1(new_n22650_), .A2(\asqrt[23] ), .B(new_n22654_), .ZN(new_n22655_));
  NOR2_X1    g22462(.A1(new_n22655_), .A2(new_n22649_), .ZN(new_n22656_));
  AOI22_X1   g22463(.A1(new_n22650_), .A2(\asqrt[23] ), .B1(new_n22648_), .B2(new_n22641_), .ZN(new_n22657_));
  NAND2_X1   g22464(.A1(new_n21987_), .A2(\asqrt[24] ), .ZN(new_n22658_));
  NOR4_X1    g22465(.A1(new_n22496_), .A2(\asqrt[24] ), .A3(new_n21982_), .A4(new_n21987_), .ZN(new_n22659_));
  XOR2_X1    g22466(.A1(new_n22659_), .A2(new_n22658_), .Z(new_n22660_));
  NAND2_X1   g22467(.A1(new_n22660_), .A2(new_n9672_), .ZN(new_n22661_));
  INV_X1     g22468(.I(new_n22661_), .ZN(new_n22662_));
  OAI21_X1   g22469(.A1(new_n22657_), .A2(new_n10104_), .B(new_n22662_), .ZN(new_n22663_));
  NAND2_X1   g22470(.A1(new_n22663_), .A2(new_n22656_), .ZN(new_n22664_));
  OAI22_X1   g22471(.A1(new_n22657_), .A2(new_n10104_), .B1(new_n22655_), .B2(new_n22649_), .ZN(new_n22665_));
  NOR4_X1    g22472(.A1(new_n22496_), .A2(\asqrt[25] ), .A3(new_n21990_), .A4(new_n22332_), .ZN(new_n22666_));
  AOI21_X1   g22473(.A1(new_n22658_), .A2(new_n21986_), .B(new_n9672_), .ZN(new_n22667_));
  NOR2_X1    g22474(.A1(new_n22666_), .A2(new_n22667_), .ZN(new_n22668_));
  NAND2_X1   g22475(.A1(new_n22668_), .A2(new_n9212_), .ZN(new_n22669_));
  AOI21_X1   g22476(.A1(new_n22665_), .A2(\asqrt[25] ), .B(new_n22669_), .ZN(new_n22670_));
  NOR2_X1    g22477(.A1(new_n22670_), .A2(new_n22664_), .ZN(new_n22671_));
  AOI22_X1   g22478(.A1(new_n22665_), .A2(\asqrt[25] ), .B1(new_n22663_), .B2(new_n22656_), .ZN(new_n22672_));
  NAND2_X1   g22479(.A1(new_n22002_), .A2(\asqrt[26] ), .ZN(new_n22673_));
  NOR4_X1    g22480(.A1(new_n22496_), .A2(\asqrt[26] ), .A3(new_n21997_), .A4(new_n22002_), .ZN(new_n22674_));
  XOR2_X1    g22481(.A1(new_n22674_), .A2(new_n22673_), .Z(new_n22675_));
  NAND2_X1   g22482(.A1(new_n22675_), .A2(new_n8763_), .ZN(new_n22676_));
  INV_X1     g22483(.I(new_n22676_), .ZN(new_n22677_));
  OAI21_X1   g22484(.A1(new_n22672_), .A2(new_n9212_), .B(new_n22677_), .ZN(new_n22678_));
  NAND2_X1   g22485(.A1(new_n22678_), .A2(new_n22671_), .ZN(new_n22679_));
  OAI22_X1   g22486(.A1(new_n22672_), .A2(new_n9212_), .B1(new_n22670_), .B2(new_n22664_), .ZN(new_n22680_));
  NOR4_X1    g22487(.A1(new_n22496_), .A2(\asqrt[27] ), .A3(new_n22005_), .A4(new_n22339_), .ZN(new_n22681_));
  AOI21_X1   g22488(.A1(new_n22673_), .A2(new_n22001_), .B(new_n8763_), .ZN(new_n22682_));
  NOR2_X1    g22489(.A1(new_n22681_), .A2(new_n22682_), .ZN(new_n22683_));
  NAND2_X1   g22490(.A1(new_n22683_), .A2(new_n8319_), .ZN(new_n22684_));
  AOI21_X1   g22491(.A1(new_n22680_), .A2(\asqrt[27] ), .B(new_n22684_), .ZN(new_n22685_));
  NOR2_X1    g22492(.A1(new_n22685_), .A2(new_n22679_), .ZN(new_n22686_));
  AOI22_X1   g22493(.A1(new_n22680_), .A2(\asqrt[27] ), .B1(new_n22678_), .B2(new_n22671_), .ZN(new_n22687_));
  NAND2_X1   g22494(.A1(new_n22017_), .A2(\asqrt[28] ), .ZN(new_n22688_));
  NOR4_X1    g22495(.A1(new_n22496_), .A2(\asqrt[28] ), .A3(new_n22012_), .A4(new_n22017_), .ZN(new_n22689_));
  XOR2_X1    g22496(.A1(new_n22689_), .A2(new_n22688_), .Z(new_n22690_));
  NAND2_X1   g22497(.A1(new_n22690_), .A2(new_n7931_), .ZN(new_n22691_));
  INV_X1     g22498(.I(new_n22691_), .ZN(new_n22692_));
  OAI21_X1   g22499(.A1(new_n22687_), .A2(new_n8319_), .B(new_n22692_), .ZN(new_n22693_));
  NAND2_X1   g22500(.A1(new_n22693_), .A2(new_n22686_), .ZN(new_n22694_));
  OAI22_X1   g22501(.A1(new_n22687_), .A2(new_n8319_), .B1(new_n22685_), .B2(new_n22679_), .ZN(new_n22695_));
  NOR4_X1    g22502(.A1(new_n22496_), .A2(\asqrt[29] ), .A3(new_n22020_), .A4(new_n22346_), .ZN(new_n22696_));
  AOI21_X1   g22503(.A1(new_n22688_), .A2(new_n22016_), .B(new_n7931_), .ZN(new_n22697_));
  NOR2_X1    g22504(.A1(new_n22696_), .A2(new_n22697_), .ZN(new_n22698_));
  NAND2_X1   g22505(.A1(new_n22698_), .A2(new_n7517_), .ZN(new_n22699_));
  AOI21_X1   g22506(.A1(new_n22695_), .A2(\asqrt[29] ), .B(new_n22699_), .ZN(new_n22700_));
  NOR2_X1    g22507(.A1(new_n22700_), .A2(new_n22694_), .ZN(new_n22701_));
  AOI22_X1   g22508(.A1(new_n22695_), .A2(\asqrt[29] ), .B1(new_n22693_), .B2(new_n22686_), .ZN(new_n22702_));
  NAND2_X1   g22509(.A1(new_n22032_), .A2(\asqrt[30] ), .ZN(new_n22703_));
  NOR4_X1    g22510(.A1(new_n22496_), .A2(\asqrt[30] ), .A3(new_n22027_), .A4(new_n22032_), .ZN(new_n22704_));
  XOR2_X1    g22511(.A1(new_n22704_), .A2(new_n22703_), .Z(new_n22705_));
  NAND2_X1   g22512(.A1(new_n22705_), .A2(new_n7110_), .ZN(new_n22706_));
  INV_X1     g22513(.I(new_n22706_), .ZN(new_n22707_));
  OAI21_X1   g22514(.A1(new_n22702_), .A2(new_n7517_), .B(new_n22707_), .ZN(new_n22708_));
  NAND2_X1   g22515(.A1(new_n22708_), .A2(new_n22701_), .ZN(new_n22709_));
  OAI22_X1   g22516(.A1(new_n22702_), .A2(new_n7517_), .B1(new_n22700_), .B2(new_n22694_), .ZN(new_n22710_));
  NOR4_X1    g22517(.A1(new_n22496_), .A2(\asqrt[31] ), .A3(new_n22035_), .A4(new_n22353_), .ZN(new_n22711_));
  AOI21_X1   g22518(.A1(new_n22703_), .A2(new_n22031_), .B(new_n7110_), .ZN(new_n22712_));
  NOR2_X1    g22519(.A1(new_n22711_), .A2(new_n22712_), .ZN(new_n22713_));
  NAND2_X1   g22520(.A1(new_n22713_), .A2(new_n6708_), .ZN(new_n22714_));
  AOI21_X1   g22521(.A1(new_n22710_), .A2(\asqrt[31] ), .B(new_n22714_), .ZN(new_n22715_));
  NOR2_X1    g22522(.A1(new_n22715_), .A2(new_n22709_), .ZN(new_n22716_));
  AOI22_X1   g22523(.A1(new_n22710_), .A2(\asqrt[31] ), .B1(new_n22708_), .B2(new_n22701_), .ZN(new_n22717_));
  NAND2_X1   g22524(.A1(new_n22047_), .A2(\asqrt[32] ), .ZN(new_n22718_));
  NOR4_X1    g22525(.A1(new_n22496_), .A2(\asqrt[32] ), .A3(new_n22042_), .A4(new_n22047_), .ZN(new_n22719_));
  XOR2_X1    g22526(.A1(new_n22719_), .A2(new_n22718_), .Z(new_n22720_));
  NAND2_X1   g22527(.A1(new_n22720_), .A2(new_n6365_), .ZN(new_n22721_));
  INV_X1     g22528(.I(new_n22721_), .ZN(new_n22722_));
  OAI21_X1   g22529(.A1(new_n22717_), .A2(new_n6708_), .B(new_n22722_), .ZN(new_n22723_));
  NAND2_X1   g22530(.A1(new_n22723_), .A2(new_n22716_), .ZN(new_n22724_));
  OAI22_X1   g22531(.A1(new_n22717_), .A2(new_n6708_), .B1(new_n22715_), .B2(new_n22709_), .ZN(new_n22725_));
  NOR4_X1    g22532(.A1(new_n22496_), .A2(\asqrt[33] ), .A3(new_n22050_), .A4(new_n22360_), .ZN(new_n22726_));
  AOI21_X1   g22533(.A1(new_n22718_), .A2(new_n22046_), .B(new_n6365_), .ZN(new_n22727_));
  NOR2_X1    g22534(.A1(new_n22726_), .A2(new_n22727_), .ZN(new_n22728_));
  NAND2_X1   g22535(.A1(new_n22728_), .A2(new_n5991_), .ZN(new_n22729_));
  AOI21_X1   g22536(.A1(new_n22725_), .A2(\asqrt[33] ), .B(new_n22729_), .ZN(new_n22730_));
  NOR2_X1    g22537(.A1(new_n22730_), .A2(new_n22724_), .ZN(new_n22731_));
  AOI22_X1   g22538(.A1(new_n22725_), .A2(\asqrt[33] ), .B1(new_n22723_), .B2(new_n22716_), .ZN(new_n22732_));
  NAND2_X1   g22539(.A1(new_n22062_), .A2(\asqrt[34] ), .ZN(new_n22733_));
  NOR4_X1    g22540(.A1(new_n22496_), .A2(\asqrt[34] ), .A3(new_n22057_), .A4(new_n22062_), .ZN(new_n22734_));
  XOR2_X1    g22541(.A1(new_n22734_), .A2(new_n22733_), .Z(new_n22735_));
  NAND2_X1   g22542(.A1(new_n22735_), .A2(new_n5626_), .ZN(new_n22736_));
  INV_X1     g22543(.I(new_n22736_), .ZN(new_n22737_));
  OAI21_X1   g22544(.A1(new_n22732_), .A2(new_n5991_), .B(new_n22737_), .ZN(new_n22738_));
  NAND2_X1   g22545(.A1(new_n22738_), .A2(new_n22731_), .ZN(new_n22739_));
  OAI22_X1   g22546(.A1(new_n22732_), .A2(new_n5991_), .B1(new_n22730_), .B2(new_n22724_), .ZN(new_n22740_));
  NOR4_X1    g22547(.A1(new_n22496_), .A2(\asqrt[35] ), .A3(new_n22065_), .A4(new_n22367_), .ZN(new_n22741_));
  AOI21_X1   g22548(.A1(new_n22733_), .A2(new_n22061_), .B(new_n5626_), .ZN(new_n22742_));
  NOR2_X1    g22549(.A1(new_n22741_), .A2(new_n22742_), .ZN(new_n22743_));
  NAND2_X1   g22550(.A1(new_n22743_), .A2(new_n5273_), .ZN(new_n22744_));
  AOI21_X1   g22551(.A1(new_n22740_), .A2(\asqrt[35] ), .B(new_n22744_), .ZN(new_n22745_));
  NOR2_X1    g22552(.A1(new_n22745_), .A2(new_n22739_), .ZN(new_n22746_));
  AOI22_X1   g22553(.A1(new_n22740_), .A2(\asqrt[35] ), .B1(new_n22738_), .B2(new_n22731_), .ZN(new_n22747_));
  NAND2_X1   g22554(.A1(new_n22077_), .A2(\asqrt[36] ), .ZN(new_n22748_));
  NOR4_X1    g22555(.A1(new_n22496_), .A2(\asqrt[36] ), .A3(new_n22072_), .A4(new_n22077_), .ZN(new_n22749_));
  XOR2_X1    g22556(.A1(new_n22749_), .A2(new_n22748_), .Z(new_n22750_));
  NAND2_X1   g22557(.A1(new_n22750_), .A2(new_n4973_), .ZN(new_n22751_));
  INV_X1     g22558(.I(new_n22751_), .ZN(new_n22752_));
  OAI21_X1   g22559(.A1(new_n22747_), .A2(new_n5273_), .B(new_n22752_), .ZN(new_n22753_));
  NAND2_X1   g22560(.A1(new_n22753_), .A2(new_n22746_), .ZN(new_n22754_));
  OAI22_X1   g22561(.A1(new_n22747_), .A2(new_n5273_), .B1(new_n22745_), .B2(new_n22739_), .ZN(new_n22755_));
  NAND2_X1   g22562(.A1(new_n22374_), .A2(\asqrt[37] ), .ZN(new_n22756_));
  NOR4_X1    g22563(.A1(new_n22496_), .A2(\asqrt[37] ), .A3(new_n22080_), .A4(new_n22374_), .ZN(new_n22757_));
  XOR2_X1    g22564(.A1(new_n22757_), .A2(new_n22756_), .Z(new_n22758_));
  NAND2_X1   g22565(.A1(new_n22758_), .A2(new_n4645_), .ZN(new_n22759_));
  AOI21_X1   g22566(.A1(new_n22755_), .A2(\asqrt[37] ), .B(new_n22759_), .ZN(new_n22760_));
  NOR2_X1    g22567(.A1(new_n22760_), .A2(new_n22754_), .ZN(new_n22761_));
  AOI22_X1   g22568(.A1(new_n22755_), .A2(\asqrt[37] ), .B1(new_n22753_), .B2(new_n22746_), .ZN(new_n22762_));
  NOR2_X1    g22569(.A1(new_n22378_), .A2(new_n4645_), .ZN(new_n22763_));
  NAND4_X1   g22570(.A1(\asqrt[3] ), .A2(new_n4645_), .A3(new_n22088_), .A4(new_n22378_), .ZN(new_n22764_));
  XOR2_X1    g22571(.A1(new_n22764_), .A2(new_n22763_), .Z(new_n22765_));
  NAND2_X1   g22572(.A1(new_n22765_), .A2(new_n4330_), .ZN(new_n22766_));
  INV_X1     g22573(.I(new_n22766_), .ZN(new_n22767_));
  OAI21_X1   g22574(.A1(new_n22762_), .A2(new_n4645_), .B(new_n22767_), .ZN(new_n22768_));
  NAND2_X1   g22575(.A1(new_n22768_), .A2(new_n22761_), .ZN(new_n22769_));
  OAI22_X1   g22576(.A1(new_n22762_), .A2(new_n4645_), .B1(new_n22760_), .B2(new_n22754_), .ZN(new_n22770_));
  NAND2_X1   g22577(.A1(new_n22382_), .A2(\asqrt[39] ), .ZN(new_n22771_));
  NOR4_X1    g22578(.A1(new_n22496_), .A2(\asqrt[39] ), .A3(new_n22095_), .A4(new_n22382_), .ZN(new_n22772_));
  XOR2_X1    g22579(.A1(new_n22772_), .A2(new_n22771_), .Z(new_n22773_));
  NAND2_X1   g22580(.A1(new_n22773_), .A2(new_n4018_), .ZN(new_n22774_));
  AOI21_X1   g22581(.A1(new_n22770_), .A2(\asqrt[39] ), .B(new_n22774_), .ZN(new_n22775_));
  NOR2_X1    g22582(.A1(new_n22775_), .A2(new_n22769_), .ZN(new_n22776_));
  AOI22_X1   g22583(.A1(new_n22770_), .A2(\asqrt[39] ), .B1(new_n22768_), .B2(new_n22761_), .ZN(new_n22777_));
  NOR2_X1    g22584(.A1(new_n22386_), .A2(new_n4018_), .ZN(new_n22778_));
  NAND4_X1   g22585(.A1(\asqrt[3] ), .A2(new_n4018_), .A3(new_n22103_), .A4(new_n22386_), .ZN(new_n22779_));
  XOR2_X1    g22586(.A1(new_n22779_), .A2(new_n22778_), .Z(new_n22780_));
  NAND2_X1   g22587(.A1(new_n22780_), .A2(new_n3760_), .ZN(new_n22781_));
  INV_X1     g22588(.I(new_n22781_), .ZN(new_n22782_));
  OAI21_X1   g22589(.A1(new_n22777_), .A2(new_n4018_), .B(new_n22782_), .ZN(new_n22783_));
  NAND2_X1   g22590(.A1(new_n22783_), .A2(new_n22776_), .ZN(new_n22784_));
  OAI22_X1   g22591(.A1(new_n22777_), .A2(new_n4018_), .B1(new_n22775_), .B2(new_n22769_), .ZN(new_n22785_));
  NAND2_X1   g22592(.A1(new_n22390_), .A2(\asqrt[41] ), .ZN(new_n22786_));
  NOR4_X1    g22593(.A1(new_n22496_), .A2(\asqrt[41] ), .A3(new_n22110_), .A4(new_n22390_), .ZN(new_n22787_));
  XOR2_X1    g22594(.A1(new_n22787_), .A2(new_n22786_), .Z(new_n22788_));
  NAND2_X1   g22595(.A1(new_n22788_), .A2(new_n3481_), .ZN(new_n22789_));
  AOI21_X1   g22596(.A1(new_n22785_), .A2(\asqrt[41] ), .B(new_n22789_), .ZN(new_n22790_));
  NOR2_X1    g22597(.A1(new_n22790_), .A2(new_n22784_), .ZN(new_n22791_));
  AOI22_X1   g22598(.A1(new_n22785_), .A2(\asqrt[41] ), .B1(new_n22783_), .B2(new_n22776_), .ZN(new_n22792_));
  NOR2_X1    g22599(.A1(new_n22394_), .A2(new_n3481_), .ZN(new_n22793_));
  NAND4_X1   g22600(.A1(\asqrt[3] ), .A2(new_n3481_), .A3(new_n22118_), .A4(new_n22394_), .ZN(new_n22794_));
  XOR2_X1    g22601(.A1(new_n22794_), .A2(new_n22793_), .Z(new_n22795_));
  NAND2_X1   g22602(.A1(new_n22795_), .A2(new_n3208_), .ZN(new_n22796_));
  INV_X1     g22603(.I(new_n22796_), .ZN(new_n22797_));
  OAI21_X1   g22604(.A1(new_n22792_), .A2(new_n3481_), .B(new_n22797_), .ZN(new_n22798_));
  NAND2_X1   g22605(.A1(new_n22798_), .A2(new_n22791_), .ZN(new_n22799_));
  OAI22_X1   g22606(.A1(new_n22792_), .A2(new_n3481_), .B1(new_n22790_), .B2(new_n22784_), .ZN(new_n22800_));
  NAND2_X1   g22607(.A1(new_n22398_), .A2(\asqrt[43] ), .ZN(new_n22801_));
  NOR4_X1    g22608(.A1(new_n22496_), .A2(\asqrt[43] ), .A3(new_n22125_), .A4(new_n22398_), .ZN(new_n22802_));
  XOR2_X1    g22609(.A1(new_n22802_), .A2(new_n22801_), .Z(new_n22803_));
  NAND2_X1   g22610(.A1(new_n22803_), .A2(new_n2941_), .ZN(new_n22804_));
  AOI21_X1   g22611(.A1(new_n22800_), .A2(\asqrt[43] ), .B(new_n22804_), .ZN(new_n22805_));
  NOR2_X1    g22612(.A1(new_n22805_), .A2(new_n22799_), .ZN(new_n22806_));
  AOI22_X1   g22613(.A1(new_n22800_), .A2(\asqrt[43] ), .B1(new_n22798_), .B2(new_n22791_), .ZN(new_n22807_));
  NAND2_X1   g22614(.A1(new_n22137_), .A2(\asqrt[44] ), .ZN(new_n22808_));
  NOR4_X1    g22615(.A1(new_n22496_), .A2(\asqrt[44] ), .A3(new_n22132_), .A4(new_n22137_), .ZN(new_n22809_));
  XOR2_X1    g22616(.A1(new_n22809_), .A2(new_n22808_), .Z(new_n22810_));
  NAND2_X1   g22617(.A1(new_n22810_), .A2(new_n2728_), .ZN(new_n22811_));
  INV_X1     g22618(.I(new_n22811_), .ZN(new_n22812_));
  OAI21_X1   g22619(.A1(new_n22807_), .A2(new_n2941_), .B(new_n22812_), .ZN(new_n22813_));
  NAND2_X1   g22620(.A1(new_n22813_), .A2(new_n22806_), .ZN(new_n22814_));
  OAI22_X1   g22621(.A1(new_n22807_), .A2(new_n2941_), .B1(new_n22805_), .B2(new_n22799_), .ZN(new_n22815_));
  NOR2_X1    g22622(.A1(new_n22146_), .A2(new_n2728_), .ZN(new_n22816_));
  NAND4_X1   g22623(.A1(\asqrt[3] ), .A2(new_n2728_), .A3(new_n22141_), .A4(new_n22146_), .ZN(new_n22817_));
  XOR2_X1    g22624(.A1(new_n22817_), .A2(new_n22816_), .Z(new_n22818_));
  NAND2_X1   g22625(.A1(new_n22818_), .A2(new_n2488_), .ZN(new_n22819_));
  AOI21_X1   g22626(.A1(new_n22815_), .A2(\asqrt[45] ), .B(new_n22819_), .ZN(new_n22820_));
  NOR2_X1    g22627(.A1(new_n22820_), .A2(new_n22814_), .ZN(new_n22821_));
  AOI22_X1   g22628(.A1(new_n22815_), .A2(\asqrt[45] ), .B1(new_n22813_), .B2(new_n22806_), .ZN(new_n22822_));
  NAND2_X1   g22629(.A1(new_n22154_), .A2(\asqrt[46] ), .ZN(new_n22823_));
  NOR4_X1    g22630(.A1(new_n22496_), .A2(\asqrt[46] ), .A3(new_n22149_), .A4(new_n22154_), .ZN(new_n22824_));
  XOR2_X1    g22631(.A1(new_n22824_), .A2(new_n22823_), .Z(new_n22825_));
  NAND2_X1   g22632(.A1(new_n22825_), .A2(new_n2253_), .ZN(new_n22826_));
  INV_X1     g22633(.I(new_n22826_), .ZN(new_n22827_));
  OAI21_X1   g22634(.A1(new_n22822_), .A2(new_n2488_), .B(new_n22827_), .ZN(new_n22828_));
  NAND2_X1   g22635(.A1(new_n22828_), .A2(new_n22821_), .ZN(new_n22829_));
  OAI22_X1   g22636(.A1(new_n22822_), .A2(new_n2488_), .B1(new_n22820_), .B2(new_n22814_), .ZN(new_n22830_));
  NAND2_X1   g22637(.A1(new_n22411_), .A2(\asqrt[47] ), .ZN(new_n22831_));
  NOR4_X1    g22638(.A1(new_n22496_), .A2(\asqrt[47] ), .A3(new_n22157_), .A4(new_n22411_), .ZN(new_n22832_));
  XOR2_X1    g22639(.A1(new_n22832_), .A2(new_n22831_), .Z(new_n22833_));
  NAND2_X1   g22640(.A1(new_n22833_), .A2(new_n2046_), .ZN(new_n22834_));
  AOI21_X1   g22641(.A1(new_n22830_), .A2(\asqrt[47] ), .B(new_n22834_), .ZN(new_n22835_));
  NOR2_X1    g22642(.A1(new_n22835_), .A2(new_n22829_), .ZN(new_n22836_));
  AOI22_X1   g22643(.A1(new_n22830_), .A2(\asqrt[47] ), .B1(new_n22828_), .B2(new_n22821_), .ZN(new_n22837_));
  NOR2_X1    g22644(.A1(new_n22415_), .A2(new_n2046_), .ZN(new_n22838_));
  NAND4_X1   g22645(.A1(\asqrt[3] ), .A2(new_n2046_), .A3(new_n22165_), .A4(new_n22415_), .ZN(new_n22839_));
  XOR2_X1    g22646(.A1(new_n22839_), .A2(new_n22838_), .Z(new_n22840_));
  NAND2_X1   g22647(.A1(new_n22840_), .A2(new_n1854_), .ZN(new_n22841_));
  INV_X1     g22648(.I(new_n22841_), .ZN(new_n22842_));
  OAI21_X1   g22649(.A1(new_n22837_), .A2(new_n2046_), .B(new_n22842_), .ZN(new_n22843_));
  NAND2_X1   g22650(.A1(new_n22843_), .A2(new_n22836_), .ZN(new_n22844_));
  OAI22_X1   g22651(.A1(new_n22837_), .A2(new_n2046_), .B1(new_n22835_), .B2(new_n22829_), .ZN(new_n22845_));
  NAND2_X1   g22652(.A1(new_n22419_), .A2(\asqrt[49] ), .ZN(new_n22846_));
  NOR4_X1    g22653(.A1(new_n22496_), .A2(\asqrt[49] ), .A3(new_n22172_), .A4(new_n22419_), .ZN(new_n22847_));
  XOR2_X1    g22654(.A1(new_n22847_), .A2(new_n22846_), .Z(new_n22848_));
  NAND2_X1   g22655(.A1(new_n22848_), .A2(new_n1595_), .ZN(new_n22849_));
  AOI21_X1   g22656(.A1(new_n22845_), .A2(\asqrt[49] ), .B(new_n22849_), .ZN(new_n22850_));
  NOR2_X1    g22657(.A1(new_n22850_), .A2(new_n22844_), .ZN(new_n22851_));
  AOI22_X1   g22658(.A1(new_n22845_), .A2(\asqrt[49] ), .B1(new_n22843_), .B2(new_n22836_), .ZN(new_n22852_));
  NOR2_X1    g22659(.A1(new_n22423_), .A2(new_n1595_), .ZN(new_n22853_));
  NAND4_X1   g22660(.A1(\asqrt[3] ), .A2(new_n1595_), .A3(new_n22180_), .A4(new_n22423_), .ZN(new_n22854_));
  XOR2_X1    g22661(.A1(new_n22854_), .A2(new_n22853_), .Z(new_n22855_));
  NAND2_X1   g22662(.A1(new_n22855_), .A2(new_n1436_), .ZN(new_n22856_));
  INV_X1     g22663(.I(new_n22856_), .ZN(new_n22857_));
  OAI21_X1   g22664(.A1(new_n22852_), .A2(new_n1595_), .B(new_n22857_), .ZN(new_n22858_));
  NAND2_X1   g22665(.A1(new_n22858_), .A2(new_n22851_), .ZN(new_n22859_));
  OAI22_X1   g22666(.A1(new_n22852_), .A2(new_n1595_), .B1(new_n22850_), .B2(new_n22844_), .ZN(new_n22860_));
  NAND2_X1   g22667(.A1(new_n22427_), .A2(\asqrt[51] ), .ZN(new_n22861_));
  NOR4_X1    g22668(.A1(new_n22496_), .A2(\asqrt[51] ), .A3(new_n22187_), .A4(new_n22427_), .ZN(new_n22862_));
  XOR2_X1    g22669(.A1(new_n22862_), .A2(new_n22861_), .Z(new_n22863_));
  NAND2_X1   g22670(.A1(new_n22863_), .A2(new_n1260_), .ZN(new_n22864_));
  AOI21_X1   g22671(.A1(new_n22860_), .A2(\asqrt[51] ), .B(new_n22864_), .ZN(new_n22865_));
  NOR2_X1    g22672(.A1(new_n22865_), .A2(new_n22859_), .ZN(new_n22866_));
  AOI22_X1   g22673(.A1(new_n22860_), .A2(\asqrt[51] ), .B1(new_n22858_), .B2(new_n22851_), .ZN(new_n22867_));
  NOR4_X1    g22674(.A1(new_n22496_), .A2(\asqrt[52] ), .A3(new_n22194_), .A4(new_n22199_), .ZN(new_n22868_));
  AOI21_X1   g22675(.A1(new_n22861_), .A2(new_n22426_), .B(new_n1260_), .ZN(new_n22869_));
  NOR2_X1    g22676(.A1(new_n22868_), .A2(new_n22869_), .ZN(new_n22870_));
  NAND2_X1   g22677(.A1(new_n22870_), .A2(new_n1096_), .ZN(new_n22871_));
  INV_X1     g22678(.I(new_n22871_), .ZN(new_n22872_));
  OAI21_X1   g22679(.A1(new_n22867_), .A2(new_n1260_), .B(new_n22872_), .ZN(new_n22873_));
  NAND2_X1   g22680(.A1(new_n22873_), .A2(new_n22866_), .ZN(new_n22874_));
  OAI22_X1   g22681(.A1(new_n22867_), .A2(new_n1260_), .B1(new_n22865_), .B2(new_n22859_), .ZN(new_n22875_));
  NAND2_X1   g22682(.A1(new_n22434_), .A2(\asqrt[53] ), .ZN(new_n22876_));
  NOR4_X1    g22683(.A1(new_n22496_), .A2(\asqrt[53] ), .A3(new_n22202_), .A4(new_n22434_), .ZN(new_n22877_));
  XOR2_X1    g22684(.A1(new_n22877_), .A2(new_n22876_), .Z(new_n22878_));
  NAND2_X1   g22685(.A1(new_n22878_), .A2(new_n970_), .ZN(new_n22879_));
  AOI21_X1   g22686(.A1(new_n22875_), .A2(\asqrt[53] ), .B(new_n22879_), .ZN(new_n22880_));
  NOR2_X1    g22687(.A1(new_n22880_), .A2(new_n22874_), .ZN(new_n22881_));
  AOI22_X1   g22688(.A1(new_n22875_), .A2(\asqrt[53] ), .B1(new_n22873_), .B2(new_n22866_), .ZN(new_n22882_));
  NOR4_X1    g22689(.A1(new_n22496_), .A2(\asqrt[54] ), .A3(new_n22209_), .A4(new_n22214_), .ZN(new_n22883_));
  AOI21_X1   g22690(.A1(new_n22876_), .A2(new_n22433_), .B(new_n970_), .ZN(new_n22884_));
  NOR2_X1    g22691(.A1(new_n22883_), .A2(new_n22884_), .ZN(new_n22885_));
  NAND2_X1   g22692(.A1(new_n22885_), .A2(new_n825_), .ZN(new_n22886_));
  INV_X1     g22693(.I(new_n22886_), .ZN(new_n22887_));
  OAI21_X1   g22694(.A1(new_n22882_), .A2(new_n970_), .B(new_n22887_), .ZN(new_n22888_));
  NAND2_X1   g22695(.A1(new_n22888_), .A2(new_n22881_), .ZN(new_n22889_));
  OAI22_X1   g22696(.A1(new_n22882_), .A2(new_n970_), .B1(new_n22880_), .B2(new_n22874_), .ZN(new_n22890_));
  NAND2_X1   g22697(.A1(new_n22441_), .A2(\asqrt[55] ), .ZN(new_n22891_));
  NOR4_X1    g22698(.A1(new_n22496_), .A2(\asqrt[55] ), .A3(new_n22217_), .A4(new_n22441_), .ZN(new_n22892_));
  XOR2_X1    g22699(.A1(new_n22892_), .A2(new_n22891_), .Z(new_n22893_));
  NAND2_X1   g22700(.A1(new_n22893_), .A2(new_n724_), .ZN(new_n22894_));
  AOI21_X1   g22701(.A1(new_n22890_), .A2(\asqrt[55] ), .B(new_n22894_), .ZN(new_n22895_));
  NOR2_X1    g22702(.A1(new_n22895_), .A2(new_n22889_), .ZN(new_n22896_));
  AOI22_X1   g22703(.A1(new_n22890_), .A2(\asqrt[55] ), .B1(new_n22888_), .B2(new_n22881_), .ZN(new_n22897_));
  NOR4_X1    g22704(.A1(new_n22496_), .A2(\asqrt[56] ), .A3(new_n22224_), .A4(new_n22229_), .ZN(new_n22898_));
  AOI21_X1   g22705(.A1(new_n22891_), .A2(new_n22440_), .B(new_n724_), .ZN(new_n22899_));
  NOR2_X1    g22706(.A1(new_n22898_), .A2(new_n22899_), .ZN(new_n22900_));
  NAND2_X1   g22707(.A1(new_n22900_), .A2(new_n587_), .ZN(new_n22901_));
  INV_X1     g22708(.I(new_n22901_), .ZN(new_n22902_));
  OAI21_X1   g22709(.A1(new_n22897_), .A2(new_n724_), .B(new_n22902_), .ZN(new_n22903_));
  NAND2_X1   g22710(.A1(new_n22903_), .A2(new_n22896_), .ZN(new_n22904_));
  OAI22_X1   g22711(.A1(new_n22897_), .A2(new_n724_), .B1(new_n22895_), .B2(new_n22889_), .ZN(new_n22905_));
  NAND2_X1   g22712(.A1(new_n22448_), .A2(\asqrt[57] ), .ZN(new_n22906_));
  NOR4_X1    g22713(.A1(new_n22496_), .A2(\asqrt[57] ), .A3(new_n22232_), .A4(new_n22448_), .ZN(new_n22907_));
  XOR2_X1    g22714(.A1(new_n22907_), .A2(new_n22906_), .Z(new_n22908_));
  NAND2_X1   g22715(.A1(new_n22908_), .A2(new_n504_), .ZN(new_n22909_));
  AOI21_X1   g22716(.A1(new_n22905_), .A2(\asqrt[57] ), .B(new_n22909_), .ZN(new_n22910_));
  NOR2_X1    g22717(.A1(new_n22910_), .A2(new_n22904_), .ZN(new_n22911_));
  AOI22_X1   g22718(.A1(new_n22905_), .A2(\asqrt[57] ), .B1(new_n22903_), .B2(new_n22896_), .ZN(new_n22912_));
  NOR2_X1    g22719(.A1(new_n22452_), .A2(new_n504_), .ZN(new_n22913_));
  NAND4_X1   g22720(.A1(\asqrt[3] ), .A2(new_n504_), .A3(new_n22239_), .A4(new_n22452_), .ZN(new_n22914_));
  XOR2_X1    g22721(.A1(new_n22914_), .A2(new_n22913_), .Z(new_n22915_));
  NAND2_X1   g22722(.A1(new_n22915_), .A2(new_n376_), .ZN(new_n22916_));
  INV_X1     g22723(.I(new_n22916_), .ZN(new_n22917_));
  OAI21_X1   g22724(.A1(new_n22912_), .A2(new_n504_), .B(new_n22917_), .ZN(new_n22918_));
  NAND2_X1   g22725(.A1(new_n22918_), .A2(new_n22911_), .ZN(new_n22919_));
  OAI22_X1   g22726(.A1(new_n22912_), .A2(new_n504_), .B1(new_n22910_), .B2(new_n22904_), .ZN(new_n22920_));
  NOR2_X1    g22727(.A1(new_n22249_), .A2(new_n376_), .ZN(new_n22921_));
  NOR4_X1    g22728(.A1(new_n22496_), .A2(\asqrt[59] ), .A3(new_n22245_), .A4(new_n22456_), .ZN(new_n22922_));
  XNOR2_X1   g22729(.A1(new_n22922_), .A2(new_n22921_), .ZN(new_n22923_));
  NAND2_X1   g22730(.A1(new_n22923_), .A2(new_n275_), .ZN(new_n22924_));
  AOI21_X1   g22731(.A1(new_n22920_), .A2(\asqrt[59] ), .B(new_n22924_), .ZN(new_n22925_));
  NOR2_X1    g22732(.A1(new_n22925_), .A2(new_n22919_), .ZN(new_n22926_));
  AOI22_X1   g22733(.A1(new_n22920_), .A2(\asqrt[59] ), .B1(new_n22918_), .B2(new_n22911_), .ZN(new_n22927_));
  NOR4_X1    g22734(.A1(new_n22496_), .A2(\asqrt[60] ), .A3(new_n22251_), .A4(new_n22256_), .ZN(new_n22928_));
  XOR2_X1    g22735(.A1(new_n22928_), .A2(new_n22257_), .Z(new_n22929_));
  NAND2_X1   g22736(.A1(new_n22929_), .A2(new_n229_), .ZN(new_n22930_));
  INV_X1     g22737(.I(new_n22930_), .ZN(new_n22931_));
  OAI21_X1   g22738(.A1(new_n22927_), .A2(new_n275_), .B(new_n22931_), .ZN(new_n22932_));
  OAI22_X1   g22739(.A1(new_n22927_), .A2(new_n275_), .B1(new_n22925_), .B2(new_n22919_), .ZN(new_n22933_));
  AOI22_X1   g22740(.A1(new_n22933_), .A2(\asqrt[61] ), .B1(new_n22932_), .B2(new_n22926_), .ZN(new_n22934_));
  NOR2_X1    g22741(.A1(new_n22934_), .A2(new_n196_), .ZN(new_n22935_));
  OAI21_X1   g22742(.A1(new_n22481_), .A2(new_n22467_), .B(new_n21588_), .ZN(new_n22936_));
  NAND3_X1   g22743(.A1(new_n22466_), .A2(\a[6] ), .A3(new_n21589_), .ZN(new_n22937_));
  NAND2_X1   g22744(.A1(new_n22936_), .A2(new_n22937_), .ZN(new_n22938_));
  OAI21_X1   g22745(.A1(new_n22938_), .A2(new_n22486_), .B(\asqrt[5] ), .ZN(new_n22939_));
  INV_X1     g22746(.I(new_n22510_), .ZN(new_n22940_));
  NOR3_X1    g22747(.A1(new_n22940_), .A2(\asqrt[6] ), .A3(new_n22507_), .ZN(new_n22941_));
  NAND2_X1   g22748(.A1(new_n22939_), .A2(new_n22941_), .ZN(new_n22942_));
  NAND2_X1   g22749(.A1(new_n22494_), .A2(new_n22939_), .ZN(new_n22943_));
  AOI22_X1   g22750(.A1(new_n22943_), .A2(\asqrt[6] ), .B1(new_n22942_), .B2(new_n22519_), .ZN(new_n22944_));
  INV_X1     g22751(.I(new_n22533_), .ZN(new_n22945_));
  OAI21_X1   g22752(.A1(new_n22944_), .A2(new_n19782_), .B(new_n22945_), .ZN(new_n22946_));
  NAND2_X1   g22753(.A1(new_n22946_), .A2(new_n22537_), .ZN(new_n22947_));
  XNOR2_X1   g22754(.A1(new_n22523_), .A2(new_n21830_), .ZN(new_n22948_));
  NAND2_X1   g22755(.A1(new_n22948_), .A2(new_n19782_), .ZN(new_n22949_));
  AOI21_X1   g22756(.A1(new_n22943_), .A2(\asqrt[6] ), .B(new_n22949_), .ZN(new_n22950_));
  OAI22_X1   g22757(.A1(new_n22944_), .A2(new_n19782_), .B1(new_n22950_), .B2(new_n22536_), .ZN(new_n22951_));
  AOI21_X1   g22758(.A1(new_n22951_), .A2(\asqrt[8] ), .B(new_n22543_), .ZN(new_n22952_));
  NOR2_X1    g22759(.A1(new_n22952_), .A2(new_n22947_), .ZN(new_n22953_));
  AOI22_X1   g22760(.A1(new_n22951_), .A2(\asqrt[8] ), .B1(new_n22946_), .B2(new_n22537_), .ZN(new_n22954_));
  INV_X1     g22761(.I(new_n22552_), .ZN(new_n22955_));
  OAI21_X1   g22762(.A1(new_n22954_), .A2(new_n18495_), .B(new_n22955_), .ZN(new_n22956_));
  NAND2_X1   g22763(.A1(new_n22956_), .A2(new_n22953_), .ZN(new_n22957_));
  OAI22_X1   g22764(.A1(new_n22954_), .A2(new_n18495_), .B1(new_n22952_), .B2(new_n22947_), .ZN(new_n22958_));
  AOI21_X1   g22765(.A1(new_n22958_), .A2(\asqrt[10] ), .B(new_n22558_), .ZN(new_n22959_));
  NOR2_X1    g22766(.A1(new_n22959_), .A2(new_n22957_), .ZN(new_n22960_));
  AOI22_X1   g22767(.A1(new_n22958_), .A2(\asqrt[10] ), .B1(new_n22956_), .B2(new_n22953_), .ZN(new_n22961_));
  INV_X1     g22768(.I(new_n22565_), .ZN(new_n22962_));
  OAI21_X1   g22769(.A1(new_n22961_), .A2(new_n17271_), .B(new_n22962_), .ZN(new_n22963_));
  NAND2_X1   g22770(.A1(new_n22963_), .A2(new_n22960_), .ZN(new_n22964_));
  OAI22_X1   g22771(.A1(new_n22961_), .A2(new_n17271_), .B1(new_n22959_), .B2(new_n22957_), .ZN(new_n22965_));
  AOI21_X1   g22772(.A1(new_n22965_), .A2(\asqrt[12] ), .B(new_n22571_), .ZN(new_n22966_));
  NOR2_X1    g22773(.A1(new_n22966_), .A2(new_n22964_), .ZN(new_n22967_));
  AOI22_X1   g22774(.A1(new_n22965_), .A2(\asqrt[12] ), .B1(new_n22963_), .B2(new_n22960_), .ZN(new_n22968_));
  INV_X1     g22775(.I(new_n22579_), .ZN(new_n22969_));
  OAI21_X1   g22776(.A1(new_n22968_), .A2(new_n16060_), .B(new_n22969_), .ZN(new_n22970_));
  NAND2_X1   g22777(.A1(new_n22970_), .A2(new_n22967_), .ZN(new_n22971_));
  OAI22_X1   g22778(.A1(new_n22968_), .A2(new_n16060_), .B1(new_n22966_), .B2(new_n22964_), .ZN(new_n22972_));
  AOI21_X1   g22779(.A1(new_n22972_), .A2(\asqrt[14] ), .B(new_n22586_), .ZN(new_n22973_));
  NOR2_X1    g22780(.A1(new_n22973_), .A2(new_n22971_), .ZN(new_n22974_));
  AOI22_X1   g22781(.A1(new_n22972_), .A2(\asqrt[14] ), .B1(new_n22970_), .B2(new_n22967_), .ZN(new_n22975_));
  INV_X1     g22782(.I(new_n22594_), .ZN(new_n22976_));
  OAI21_X1   g22783(.A1(new_n22975_), .A2(new_n14871_), .B(new_n22976_), .ZN(new_n22977_));
  NAND2_X1   g22784(.A1(new_n22977_), .A2(new_n22974_), .ZN(new_n22978_));
  OAI22_X1   g22785(.A1(new_n22975_), .A2(new_n14871_), .B1(new_n22973_), .B2(new_n22971_), .ZN(new_n22979_));
  AOI21_X1   g22786(.A1(new_n22979_), .A2(\asqrt[16] ), .B(new_n22601_), .ZN(new_n22980_));
  NOR2_X1    g22787(.A1(new_n22980_), .A2(new_n22978_), .ZN(new_n22981_));
  AOI22_X1   g22788(.A1(new_n22979_), .A2(\asqrt[16] ), .B1(new_n22977_), .B2(new_n22974_), .ZN(new_n22982_));
  INV_X1     g22789(.I(new_n22609_), .ZN(new_n22983_));
  OAI21_X1   g22790(.A1(new_n22982_), .A2(new_n13760_), .B(new_n22983_), .ZN(new_n22984_));
  NAND2_X1   g22791(.A1(new_n22984_), .A2(new_n22981_), .ZN(new_n22985_));
  OAI22_X1   g22792(.A1(new_n22982_), .A2(new_n13760_), .B1(new_n22980_), .B2(new_n22978_), .ZN(new_n22986_));
  AOI21_X1   g22793(.A1(new_n22986_), .A2(\asqrt[18] ), .B(new_n22616_), .ZN(new_n22987_));
  NOR2_X1    g22794(.A1(new_n22987_), .A2(new_n22985_), .ZN(new_n22988_));
  AOI22_X1   g22795(.A1(new_n22986_), .A2(\asqrt[18] ), .B1(new_n22984_), .B2(new_n22981_), .ZN(new_n22989_));
  INV_X1     g22796(.I(new_n22624_), .ZN(new_n22990_));
  OAI21_X1   g22797(.A1(new_n22989_), .A2(new_n12657_), .B(new_n22990_), .ZN(new_n22991_));
  NAND2_X1   g22798(.A1(new_n22991_), .A2(new_n22988_), .ZN(new_n22992_));
  OAI22_X1   g22799(.A1(new_n22989_), .A2(new_n12657_), .B1(new_n22987_), .B2(new_n22985_), .ZN(new_n22993_));
  AOI21_X1   g22800(.A1(new_n22993_), .A2(\asqrt[20] ), .B(new_n22631_), .ZN(new_n22994_));
  NOR2_X1    g22801(.A1(new_n22994_), .A2(new_n22992_), .ZN(new_n22995_));
  AOI22_X1   g22802(.A1(new_n22993_), .A2(\asqrt[20] ), .B1(new_n22991_), .B2(new_n22988_), .ZN(new_n22996_));
  INV_X1     g22803(.I(new_n22639_), .ZN(new_n22997_));
  OAI21_X1   g22804(.A1(new_n22996_), .A2(new_n11631_), .B(new_n22997_), .ZN(new_n22998_));
  NAND2_X1   g22805(.A1(new_n22998_), .A2(new_n22995_), .ZN(new_n22999_));
  OAI22_X1   g22806(.A1(new_n22996_), .A2(new_n11631_), .B1(new_n22994_), .B2(new_n22992_), .ZN(new_n23000_));
  AOI21_X1   g22807(.A1(new_n23000_), .A2(\asqrt[22] ), .B(new_n22646_), .ZN(new_n23001_));
  NOR2_X1    g22808(.A1(new_n23001_), .A2(new_n22999_), .ZN(new_n23002_));
  AOI22_X1   g22809(.A1(new_n23000_), .A2(\asqrt[22] ), .B1(new_n22998_), .B2(new_n22995_), .ZN(new_n23003_));
  INV_X1     g22810(.I(new_n22654_), .ZN(new_n23004_));
  OAI21_X1   g22811(.A1(new_n23003_), .A2(new_n10614_), .B(new_n23004_), .ZN(new_n23005_));
  NAND2_X1   g22812(.A1(new_n23005_), .A2(new_n23002_), .ZN(new_n23006_));
  OAI22_X1   g22813(.A1(new_n23003_), .A2(new_n10614_), .B1(new_n23001_), .B2(new_n22999_), .ZN(new_n23007_));
  AOI21_X1   g22814(.A1(new_n23007_), .A2(\asqrt[24] ), .B(new_n22661_), .ZN(new_n23008_));
  NOR2_X1    g22815(.A1(new_n23008_), .A2(new_n23006_), .ZN(new_n23009_));
  AOI22_X1   g22816(.A1(new_n23007_), .A2(\asqrt[24] ), .B1(new_n23005_), .B2(new_n23002_), .ZN(new_n23010_));
  INV_X1     g22817(.I(new_n22669_), .ZN(new_n23011_));
  OAI21_X1   g22818(.A1(new_n23010_), .A2(new_n9672_), .B(new_n23011_), .ZN(new_n23012_));
  NAND2_X1   g22819(.A1(new_n23012_), .A2(new_n23009_), .ZN(new_n23013_));
  OAI22_X1   g22820(.A1(new_n23010_), .A2(new_n9672_), .B1(new_n23008_), .B2(new_n23006_), .ZN(new_n23014_));
  AOI21_X1   g22821(.A1(new_n23014_), .A2(\asqrt[26] ), .B(new_n22676_), .ZN(new_n23015_));
  NOR2_X1    g22822(.A1(new_n23015_), .A2(new_n23013_), .ZN(new_n23016_));
  AOI22_X1   g22823(.A1(new_n23014_), .A2(\asqrt[26] ), .B1(new_n23012_), .B2(new_n23009_), .ZN(new_n23017_));
  INV_X1     g22824(.I(new_n22684_), .ZN(new_n23018_));
  OAI21_X1   g22825(.A1(new_n23017_), .A2(new_n8763_), .B(new_n23018_), .ZN(new_n23019_));
  NAND2_X1   g22826(.A1(new_n23019_), .A2(new_n23016_), .ZN(new_n23020_));
  OAI22_X1   g22827(.A1(new_n23017_), .A2(new_n8763_), .B1(new_n23015_), .B2(new_n23013_), .ZN(new_n23021_));
  AOI21_X1   g22828(.A1(new_n23021_), .A2(\asqrt[28] ), .B(new_n22691_), .ZN(new_n23022_));
  NOR2_X1    g22829(.A1(new_n23022_), .A2(new_n23020_), .ZN(new_n23023_));
  AOI22_X1   g22830(.A1(new_n23021_), .A2(\asqrt[28] ), .B1(new_n23019_), .B2(new_n23016_), .ZN(new_n23024_));
  INV_X1     g22831(.I(new_n22699_), .ZN(new_n23025_));
  OAI21_X1   g22832(.A1(new_n23024_), .A2(new_n7931_), .B(new_n23025_), .ZN(new_n23026_));
  NAND2_X1   g22833(.A1(new_n23026_), .A2(new_n23023_), .ZN(new_n23027_));
  OAI22_X1   g22834(.A1(new_n23024_), .A2(new_n7931_), .B1(new_n23022_), .B2(new_n23020_), .ZN(new_n23028_));
  AOI21_X1   g22835(.A1(new_n23028_), .A2(\asqrt[30] ), .B(new_n22706_), .ZN(new_n23029_));
  NOR2_X1    g22836(.A1(new_n23029_), .A2(new_n23027_), .ZN(new_n23030_));
  AOI22_X1   g22837(.A1(new_n23028_), .A2(\asqrt[30] ), .B1(new_n23026_), .B2(new_n23023_), .ZN(new_n23031_));
  INV_X1     g22838(.I(new_n22714_), .ZN(new_n23032_));
  OAI21_X1   g22839(.A1(new_n23031_), .A2(new_n7110_), .B(new_n23032_), .ZN(new_n23033_));
  NAND2_X1   g22840(.A1(new_n23033_), .A2(new_n23030_), .ZN(new_n23034_));
  OAI22_X1   g22841(.A1(new_n23031_), .A2(new_n7110_), .B1(new_n23029_), .B2(new_n23027_), .ZN(new_n23035_));
  AOI21_X1   g22842(.A1(new_n23035_), .A2(\asqrt[32] ), .B(new_n22721_), .ZN(new_n23036_));
  NOR2_X1    g22843(.A1(new_n23036_), .A2(new_n23034_), .ZN(new_n23037_));
  AOI22_X1   g22844(.A1(new_n23035_), .A2(\asqrt[32] ), .B1(new_n23033_), .B2(new_n23030_), .ZN(new_n23038_));
  INV_X1     g22845(.I(new_n22729_), .ZN(new_n23039_));
  OAI21_X1   g22846(.A1(new_n23038_), .A2(new_n6365_), .B(new_n23039_), .ZN(new_n23040_));
  NAND2_X1   g22847(.A1(new_n23040_), .A2(new_n23037_), .ZN(new_n23041_));
  OAI22_X1   g22848(.A1(new_n23038_), .A2(new_n6365_), .B1(new_n23036_), .B2(new_n23034_), .ZN(new_n23042_));
  AOI21_X1   g22849(.A1(new_n23042_), .A2(\asqrt[34] ), .B(new_n22736_), .ZN(new_n23043_));
  NOR2_X1    g22850(.A1(new_n23043_), .A2(new_n23041_), .ZN(new_n23044_));
  AOI22_X1   g22851(.A1(new_n23042_), .A2(\asqrt[34] ), .B1(new_n23040_), .B2(new_n23037_), .ZN(new_n23045_));
  INV_X1     g22852(.I(new_n22744_), .ZN(new_n23046_));
  OAI21_X1   g22853(.A1(new_n23045_), .A2(new_n5626_), .B(new_n23046_), .ZN(new_n23047_));
  NAND2_X1   g22854(.A1(new_n23047_), .A2(new_n23044_), .ZN(new_n23048_));
  OAI22_X1   g22855(.A1(new_n23045_), .A2(new_n5626_), .B1(new_n23043_), .B2(new_n23041_), .ZN(new_n23049_));
  AOI21_X1   g22856(.A1(new_n23049_), .A2(\asqrt[36] ), .B(new_n22751_), .ZN(new_n23050_));
  NOR2_X1    g22857(.A1(new_n23050_), .A2(new_n23048_), .ZN(new_n23051_));
  AOI22_X1   g22858(.A1(new_n23049_), .A2(\asqrt[36] ), .B1(new_n23047_), .B2(new_n23044_), .ZN(new_n23052_));
  INV_X1     g22859(.I(new_n22759_), .ZN(new_n23053_));
  OAI21_X1   g22860(.A1(new_n23052_), .A2(new_n4973_), .B(new_n23053_), .ZN(new_n23054_));
  NAND2_X1   g22861(.A1(new_n23054_), .A2(new_n23051_), .ZN(new_n23055_));
  OAI22_X1   g22862(.A1(new_n23052_), .A2(new_n4973_), .B1(new_n23050_), .B2(new_n23048_), .ZN(new_n23056_));
  AOI21_X1   g22863(.A1(new_n23056_), .A2(\asqrt[38] ), .B(new_n22766_), .ZN(new_n23057_));
  NOR2_X1    g22864(.A1(new_n23057_), .A2(new_n23055_), .ZN(new_n23058_));
  AOI22_X1   g22865(.A1(new_n23056_), .A2(\asqrt[38] ), .B1(new_n23054_), .B2(new_n23051_), .ZN(new_n23059_));
  INV_X1     g22866(.I(new_n22774_), .ZN(new_n23060_));
  OAI21_X1   g22867(.A1(new_n23059_), .A2(new_n4330_), .B(new_n23060_), .ZN(new_n23061_));
  NAND2_X1   g22868(.A1(new_n23061_), .A2(new_n23058_), .ZN(new_n23062_));
  OAI22_X1   g22869(.A1(new_n23059_), .A2(new_n4330_), .B1(new_n23057_), .B2(new_n23055_), .ZN(new_n23063_));
  AOI21_X1   g22870(.A1(new_n23063_), .A2(\asqrt[40] ), .B(new_n22781_), .ZN(new_n23064_));
  NOR2_X1    g22871(.A1(new_n23064_), .A2(new_n23062_), .ZN(new_n23065_));
  AOI22_X1   g22872(.A1(new_n23063_), .A2(\asqrt[40] ), .B1(new_n23061_), .B2(new_n23058_), .ZN(new_n23066_));
  INV_X1     g22873(.I(new_n22789_), .ZN(new_n23067_));
  OAI21_X1   g22874(.A1(new_n23066_), .A2(new_n3760_), .B(new_n23067_), .ZN(new_n23068_));
  NAND2_X1   g22875(.A1(new_n23068_), .A2(new_n23065_), .ZN(new_n23069_));
  OAI22_X1   g22876(.A1(new_n23066_), .A2(new_n3760_), .B1(new_n23064_), .B2(new_n23062_), .ZN(new_n23070_));
  AOI21_X1   g22877(.A1(new_n23070_), .A2(\asqrt[42] ), .B(new_n22796_), .ZN(new_n23071_));
  NOR2_X1    g22878(.A1(new_n23071_), .A2(new_n23069_), .ZN(new_n23072_));
  AOI22_X1   g22879(.A1(new_n23070_), .A2(\asqrt[42] ), .B1(new_n23068_), .B2(new_n23065_), .ZN(new_n23073_));
  INV_X1     g22880(.I(new_n22804_), .ZN(new_n23074_));
  OAI21_X1   g22881(.A1(new_n23073_), .A2(new_n3208_), .B(new_n23074_), .ZN(new_n23075_));
  NAND2_X1   g22882(.A1(new_n23075_), .A2(new_n23072_), .ZN(new_n23076_));
  OAI22_X1   g22883(.A1(new_n23073_), .A2(new_n3208_), .B1(new_n23071_), .B2(new_n23069_), .ZN(new_n23077_));
  AOI21_X1   g22884(.A1(new_n23077_), .A2(\asqrt[44] ), .B(new_n22811_), .ZN(new_n23078_));
  NOR2_X1    g22885(.A1(new_n23078_), .A2(new_n23076_), .ZN(new_n23079_));
  AOI22_X1   g22886(.A1(new_n23077_), .A2(\asqrt[44] ), .B1(new_n23075_), .B2(new_n23072_), .ZN(new_n23080_));
  INV_X1     g22887(.I(new_n22819_), .ZN(new_n23081_));
  OAI21_X1   g22888(.A1(new_n23080_), .A2(new_n2728_), .B(new_n23081_), .ZN(new_n23082_));
  NAND2_X1   g22889(.A1(new_n23082_), .A2(new_n23079_), .ZN(new_n23083_));
  OAI22_X1   g22890(.A1(new_n23080_), .A2(new_n2728_), .B1(new_n23078_), .B2(new_n23076_), .ZN(new_n23084_));
  AOI21_X1   g22891(.A1(new_n23084_), .A2(\asqrt[46] ), .B(new_n22826_), .ZN(new_n23085_));
  NOR2_X1    g22892(.A1(new_n23085_), .A2(new_n23083_), .ZN(new_n23086_));
  AOI22_X1   g22893(.A1(new_n23084_), .A2(\asqrt[46] ), .B1(new_n23082_), .B2(new_n23079_), .ZN(new_n23087_));
  INV_X1     g22894(.I(new_n22834_), .ZN(new_n23088_));
  OAI21_X1   g22895(.A1(new_n23087_), .A2(new_n2253_), .B(new_n23088_), .ZN(new_n23089_));
  NAND2_X1   g22896(.A1(new_n23089_), .A2(new_n23086_), .ZN(new_n23090_));
  OAI22_X1   g22897(.A1(new_n23087_), .A2(new_n2253_), .B1(new_n23085_), .B2(new_n23083_), .ZN(new_n23091_));
  AOI21_X1   g22898(.A1(new_n23091_), .A2(\asqrt[48] ), .B(new_n22841_), .ZN(new_n23092_));
  NOR2_X1    g22899(.A1(new_n23092_), .A2(new_n23090_), .ZN(new_n23093_));
  AOI22_X1   g22900(.A1(new_n23091_), .A2(\asqrt[48] ), .B1(new_n23089_), .B2(new_n23086_), .ZN(new_n23094_));
  INV_X1     g22901(.I(new_n22849_), .ZN(new_n23095_));
  OAI21_X1   g22902(.A1(new_n23094_), .A2(new_n1854_), .B(new_n23095_), .ZN(new_n23096_));
  NAND2_X1   g22903(.A1(new_n23096_), .A2(new_n23093_), .ZN(new_n23097_));
  OAI22_X1   g22904(.A1(new_n23094_), .A2(new_n1854_), .B1(new_n23092_), .B2(new_n23090_), .ZN(new_n23098_));
  AOI21_X1   g22905(.A1(new_n23098_), .A2(\asqrt[50] ), .B(new_n22856_), .ZN(new_n23099_));
  NOR2_X1    g22906(.A1(new_n23099_), .A2(new_n23097_), .ZN(new_n23100_));
  AOI22_X1   g22907(.A1(new_n23098_), .A2(\asqrt[50] ), .B1(new_n23096_), .B2(new_n23093_), .ZN(new_n23101_));
  INV_X1     g22908(.I(new_n22864_), .ZN(new_n23102_));
  OAI21_X1   g22909(.A1(new_n23101_), .A2(new_n1436_), .B(new_n23102_), .ZN(new_n23103_));
  NAND2_X1   g22910(.A1(new_n23103_), .A2(new_n23100_), .ZN(new_n23104_));
  OAI22_X1   g22911(.A1(new_n23101_), .A2(new_n1436_), .B1(new_n23099_), .B2(new_n23097_), .ZN(new_n23105_));
  AOI21_X1   g22912(.A1(new_n23105_), .A2(\asqrt[52] ), .B(new_n22871_), .ZN(new_n23106_));
  NOR2_X1    g22913(.A1(new_n23106_), .A2(new_n23104_), .ZN(new_n23107_));
  AOI22_X1   g22914(.A1(new_n23105_), .A2(\asqrt[52] ), .B1(new_n23103_), .B2(new_n23100_), .ZN(new_n23108_));
  INV_X1     g22915(.I(new_n22879_), .ZN(new_n23109_));
  OAI21_X1   g22916(.A1(new_n23108_), .A2(new_n1096_), .B(new_n23109_), .ZN(new_n23110_));
  NAND2_X1   g22917(.A1(new_n23110_), .A2(new_n23107_), .ZN(new_n23111_));
  OAI22_X1   g22918(.A1(new_n23108_), .A2(new_n1096_), .B1(new_n23106_), .B2(new_n23104_), .ZN(new_n23112_));
  AOI21_X1   g22919(.A1(new_n23112_), .A2(\asqrt[54] ), .B(new_n22886_), .ZN(new_n23113_));
  NOR2_X1    g22920(.A1(new_n23113_), .A2(new_n23111_), .ZN(new_n23114_));
  AOI22_X1   g22921(.A1(new_n23112_), .A2(\asqrt[54] ), .B1(new_n23110_), .B2(new_n23107_), .ZN(new_n23115_));
  INV_X1     g22922(.I(new_n22894_), .ZN(new_n23116_));
  OAI21_X1   g22923(.A1(new_n23115_), .A2(new_n825_), .B(new_n23116_), .ZN(new_n23117_));
  NAND2_X1   g22924(.A1(new_n23117_), .A2(new_n23114_), .ZN(new_n23118_));
  OAI22_X1   g22925(.A1(new_n23115_), .A2(new_n825_), .B1(new_n23113_), .B2(new_n23111_), .ZN(new_n23119_));
  AOI21_X1   g22926(.A1(new_n23119_), .A2(\asqrt[56] ), .B(new_n22901_), .ZN(new_n23120_));
  NOR2_X1    g22927(.A1(new_n23120_), .A2(new_n23118_), .ZN(new_n23121_));
  AOI22_X1   g22928(.A1(new_n23119_), .A2(\asqrt[56] ), .B1(new_n23117_), .B2(new_n23114_), .ZN(new_n23122_));
  INV_X1     g22929(.I(new_n22909_), .ZN(new_n23123_));
  OAI21_X1   g22930(.A1(new_n23122_), .A2(new_n587_), .B(new_n23123_), .ZN(new_n23124_));
  NAND2_X1   g22931(.A1(new_n23124_), .A2(new_n23121_), .ZN(new_n23125_));
  OAI22_X1   g22932(.A1(new_n23122_), .A2(new_n587_), .B1(new_n23120_), .B2(new_n23118_), .ZN(new_n23126_));
  AOI21_X1   g22933(.A1(new_n23126_), .A2(\asqrt[58] ), .B(new_n22916_), .ZN(new_n23127_));
  NOR2_X1    g22934(.A1(new_n23127_), .A2(new_n23125_), .ZN(new_n23128_));
  AOI22_X1   g22935(.A1(new_n23126_), .A2(\asqrt[58] ), .B1(new_n23124_), .B2(new_n23121_), .ZN(new_n23129_));
  INV_X1     g22936(.I(new_n22924_), .ZN(new_n23130_));
  OAI21_X1   g22937(.A1(new_n23129_), .A2(new_n376_), .B(new_n23130_), .ZN(new_n23131_));
  NAND2_X1   g22938(.A1(new_n23131_), .A2(new_n23128_), .ZN(new_n23132_));
  OAI22_X1   g22939(.A1(new_n23129_), .A2(new_n376_), .B1(new_n23127_), .B2(new_n23125_), .ZN(new_n23133_));
  AOI21_X1   g22940(.A1(new_n23133_), .A2(\asqrt[60] ), .B(new_n22930_), .ZN(new_n23134_));
  AOI22_X1   g22941(.A1(new_n23133_), .A2(\asqrt[60] ), .B1(new_n23131_), .B2(new_n23128_), .ZN(new_n23135_));
  OAI22_X1   g22942(.A1(new_n23135_), .A2(new_n229_), .B1(new_n23134_), .B2(new_n23132_), .ZN(new_n23136_));
  NOR3_X1    g22943(.A1(new_n22462_), .A2(\asqrt[61] ), .A3(new_n22259_), .ZN(new_n23137_));
  NAND2_X1   g22944(.A1(\asqrt[3] ), .A2(new_n23137_), .ZN(new_n23138_));
  XOR2_X1    g22945(.A1(new_n23138_), .A2(new_n22478_), .Z(new_n23139_));
  OAI21_X1   g22946(.A1(new_n22262_), .A2(new_n22478_), .B(\asqrt[62] ), .ZN(new_n23140_));
  NAND2_X1   g22947(.A1(\asqrt[3] ), .A2(new_n22479_), .ZN(new_n23141_));
  XNOR2_X1   g22948(.A1(new_n23141_), .A2(new_n23140_), .ZN(new_n23142_));
  NAND2_X1   g22949(.A1(new_n23133_), .A2(\asqrt[60] ), .ZN(new_n23143_));
  AOI21_X1   g22950(.A1(new_n23143_), .A2(new_n23132_), .B(new_n229_), .ZN(new_n23144_));
  NOR2_X1    g22951(.A1(new_n23139_), .A2(new_n196_), .ZN(new_n23145_));
  INV_X1     g22952(.I(new_n23139_), .ZN(new_n23146_));
  NOR2_X1    g22953(.A1(new_n23146_), .A2(\asqrt[62] ), .ZN(new_n23147_));
  NOR3_X1    g22954(.A1(new_n23134_), .A2(new_n23132_), .A3(new_n23147_), .ZN(new_n23148_));
  AOI21_X1   g22955(.A1(new_n23148_), .A2(new_n23144_), .B(new_n23145_), .ZN(new_n23149_));
  AND3_X2    g22956(.A1(new_n22496_), .A2(new_n21783_), .A3(new_n22464_), .Z(new_n23150_));
  OAI21_X1   g22957(.A1(new_n23150_), .A2(new_n22267_), .B(new_n231_), .ZN(new_n23151_));
  INV_X1     g22958(.I(new_n23151_), .ZN(new_n23152_));
  AOI21_X1   g22959(.A1(new_n23149_), .A2(new_n23152_), .B(new_n23142_), .ZN(new_n23153_));
  NAND2_X1   g22960(.A1(new_n22267_), .A2(new_n21783_), .ZN(new_n23154_));
  XOR2_X1    g22961(.A1(new_n22475_), .A2(new_n231_), .Z(new_n23155_));
  AOI21_X1   g22962(.A1(\asqrt[3] ), .A2(new_n23154_), .B(new_n23155_), .ZN(new_n23156_));
  NOR4_X1    g22963(.A1(new_n23136_), .A2(\asqrt[62] ), .A3(new_n23139_), .A4(new_n23142_), .ZN(new_n23157_));
  NOR3_X1    g22964(.A1(new_n23153_), .A2(new_n23156_), .A3(new_n23157_), .ZN(new_n23158_));
  NOR4_X1    g22965(.A1(new_n23158_), .A2(\asqrt[62] ), .A3(new_n23136_), .A4(new_n23139_), .ZN(new_n23159_));
  XNOR2_X1   g22966(.A1(new_n23159_), .A2(new_n22935_), .ZN(new_n23160_));
  NAND2_X1   g22967(.A1(new_n22905_), .A2(\asqrt[57] ), .ZN(new_n23161_));
  AOI21_X1   g22968(.A1(new_n23161_), .A2(new_n22904_), .B(new_n504_), .ZN(new_n23162_));
  OAI21_X1   g22969(.A1(new_n22911_), .A2(new_n23162_), .B(\asqrt[59] ), .ZN(new_n23163_));
  AOI21_X1   g22970(.A1(new_n22919_), .A2(new_n23163_), .B(new_n275_), .ZN(new_n23164_));
  OAI21_X1   g22971(.A1(new_n22926_), .A2(new_n23164_), .B(\asqrt[61] ), .ZN(new_n23165_));
  NOR4_X1    g22972(.A1(new_n23158_), .A2(\asqrt[61] ), .A3(new_n22929_), .A4(new_n22933_), .ZN(new_n23166_));
  XOR2_X1    g22973(.A1(new_n23166_), .A2(new_n23165_), .Z(new_n23167_));
  NOR2_X1    g22974(.A1(new_n23167_), .A2(new_n196_), .ZN(new_n23168_));
  NOR2_X1    g22975(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n23169_));
  NAND4_X1   g22976(.A1(new_n22465_), .A2(new_n22476_), .A3(\a[4] ), .A4(new_n23169_), .ZN(new_n23170_));
  XOR2_X1    g22977(.A1(new_n23170_), .A2(\a[5] ), .Z(new_n23171_));
  INV_X1     g22978(.I(\a[5] ), .ZN(new_n23172_));
  INV_X1     g22979(.I(new_n23142_), .ZN(new_n23173_));
  INV_X1     g22980(.I(new_n23145_), .ZN(new_n23174_));
  INV_X1     g22981(.I(new_n23147_), .ZN(new_n23175_));
  NAND3_X1   g22982(.A1(new_n22932_), .A2(new_n22926_), .A3(new_n23175_), .ZN(new_n23176_));
  OAI21_X1   g22983(.A1(new_n23176_), .A2(new_n23165_), .B(new_n23174_), .ZN(new_n23177_));
  OAI21_X1   g22984(.A1(new_n23177_), .A2(new_n23151_), .B(new_n23173_), .ZN(new_n23178_));
  NOR2_X1    g22985(.A1(new_n23157_), .A2(new_n23156_), .ZN(new_n23179_));
  AOI21_X1   g22986(.A1(new_n23179_), .A2(new_n23178_), .B(new_n23172_), .ZN(new_n23180_));
  NOR2_X1    g22987(.A1(new_n23172_), .A2(\a[4] ), .ZN(new_n23181_));
  OAI21_X1   g22988(.A1(new_n23180_), .A2(new_n23181_), .B(new_n23171_), .ZN(new_n23182_));
  INV_X1     g22989(.I(new_n23171_), .ZN(new_n23183_));
  INV_X1     g22990(.I(new_n23156_), .ZN(new_n23184_));
  NAND4_X1   g22991(.A1(new_n22934_), .A2(new_n196_), .A3(new_n23146_), .A4(new_n23173_), .ZN(new_n23185_));
  NAND2_X1   g22992(.A1(new_n23185_), .A2(new_n23184_), .ZN(new_n23186_));
  OAI21_X1   g22993(.A1(new_n23186_), .A2(new_n23153_), .B(\a[5] ), .ZN(new_n23187_));
  NAND3_X1   g22994(.A1(new_n23187_), .A2(\a[4] ), .A3(new_n23183_), .ZN(new_n23188_));
  NAND2_X1   g22995(.A1(new_n23182_), .A2(new_n23188_), .ZN(new_n23189_));
  NAND2_X1   g22996(.A1(\asqrt[3] ), .A2(\a[4] ), .ZN(new_n23190_));
  AOI21_X1   g22997(.A1(new_n23158_), .A2(\asqrt[3] ), .B(new_n23190_), .ZN(new_n23191_));
  NOR4_X1    g22998(.A1(new_n23186_), .A2(\a[4] ), .A3(new_n22496_), .A4(new_n23153_), .ZN(new_n23192_));
  OAI21_X1   g22999(.A1(new_n23191_), .A2(new_n23192_), .B(new_n23169_), .ZN(new_n23193_));
  NAND3_X1   g23000(.A1(new_n23157_), .A2(\asqrt[3] ), .A3(new_n23156_), .ZN(new_n23194_));
  OAI21_X1   g23001(.A1(new_n23194_), .A2(new_n23178_), .B(new_n22470_), .ZN(new_n23195_));
  NAND3_X1   g23002(.A1(new_n23195_), .A2(new_n21584_), .A3(new_n23158_), .ZN(new_n23196_));
  NAND3_X1   g23003(.A1(new_n23178_), .A2(new_n23184_), .A3(new_n23185_), .ZN(\asqrt[2] ));
  NOR3_X1    g23004(.A1(new_n23185_), .A2(new_n22496_), .A3(new_n23184_), .ZN(new_n23198_));
  AOI21_X1   g23005(.A1(new_n23198_), .A2(new_n23153_), .B(\a[6] ), .ZN(new_n23199_));
  OAI21_X1   g23006(.A1(new_n23199_), .A2(new_n21585_), .B(\asqrt[2] ), .ZN(new_n23200_));
  NAND4_X1   g23007(.A1(new_n23193_), .A2(new_n21781_), .A3(new_n23196_), .A4(new_n23200_), .ZN(new_n23201_));
  NAND2_X1   g23008(.A1(new_n23201_), .A2(new_n23189_), .ZN(new_n23202_));
  NAND3_X1   g23009(.A1(new_n23193_), .A2(new_n23182_), .A3(new_n23188_), .ZN(new_n23203_));
  NOR2_X1    g23010(.A1(new_n22496_), .A2(\a[6] ), .ZN(new_n23204_));
  OAI22_X1   g23011(.A1(new_n23204_), .A2(\a[7] ), .B1(\a[6] ), .B2(new_n22466_), .ZN(new_n23205_));
  NAND2_X1   g23012(.A1(new_n22486_), .A2(new_n21587_), .ZN(new_n23206_));
  AOI21_X1   g23013(.A1(new_n23206_), .A2(new_n22470_), .B(new_n22496_), .ZN(new_n23207_));
  AOI21_X1   g23014(.A1(\asqrt[2] ), .A2(new_n23207_), .B(new_n23205_), .ZN(new_n23208_));
  INV_X1     g23015(.I(new_n23208_), .ZN(new_n23209_));
  AND2_X2    g23016(.A1(new_n23207_), .A2(new_n23205_), .Z(new_n23210_));
  NAND2_X1   g23017(.A1(\asqrt[2] ), .A2(new_n23210_), .ZN(new_n23211_));
  NAND3_X1   g23018(.A1(new_n23209_), .A2(new_n21079_), .A3(new_n23211_), .ZN(new_n23212_));
  AOI21_X1   g23019(.A1(new_n23203_), .A2(\asqrt[4] ), .B(new_n23212_), .ZN(new_n23213_));
  NOR2_X1    g23020(.A1(new_n23213_), .A2(new_n23202_), .ZN(new_n23214_));
  AOI22_X1   g23021(.A1(new_n23201_), .A2(new_n23189_), .B1(new_n23203_), .B2(\asqrt[4] ), .ZN(new_n23215_));
  NOR2_X1    g23022(.A1(new_n22517_), .A2(new_n22514_), .ZN(new_n23216_));
  NAND2_X1   g23023(.A1(new_n22495_), .A2(new_n22500_), .ZN(new_n23217_));
  OR4_X2     g23024(.A1(\asqrt[5] ), .A2(new_n23158_), .A3(new_n23216_), .A4(new_n23217_), .Z(new_n23218_));
  OAI21_X1   g23025(.A1(new_n22938_), .A2(new_n22486_), .B(\asqrt[5] ), .ZN(new_n23219_));
  NAND3_X1   g23026(.A1(new_n23218_), .A2(new_n20455_), .A3(new_n23219_), .ZN(new_n23220_));
  INV_X1     g23027(.I(new_n23220_), .ZN(new_n23221_));
  OAI21_X1   g23028(.A1(new_n23215_), .A2(new_n21079_), .B(new_n23221_), .ZN(new_n23222_));
  NAND2_X1   g23029(.A1(new_n23222_), .A2(new_n23214_), .ZN(new_n23223_));
  OAI22_X1   g23030(.A1(new_n23215_), .A2(new_n21079_), .B1(new_n23202_), .B2(new_n23213_), .ZN(new_n23224_));
  NOR2_X1    g23031(.A1(new_n22940_), .A2(new_n22507_), .ZN(new_n23225_));
  NOR4_X1    g23032(.A1(new_n23158_), .A2(\asqrt[6] ), .A3(new_n23225_), .A4(new_n22943_), .ZN(new_n23226_));
  XOR2_X1    g23033(.A1(new_n23226_), .A2(new_n22520_), .Z(new_n23227_));
  NAND2_X1   g23034(.A1(new_n23227_), .A2(new_n19782_), .ZN(new_n23228_));
  AOI21_X1   g23035(.A1(new_n23224_), .A2(\asqrt[6] ), .B(new_n23228_), .ZN(new_n23229_));
  NOR2_X1    g23036(.A1(new_n23229_), .A2(new_n23223_), .ZN(new_n23230_));
  AOI22_X1   g23037(.A1(new_n23224_), .A2(\asqrt[6] ), .B1(new_n23222_), .B2(new_n23214_), .ZN(new_n23231_));
  NAND4_X1   g23038(.A1(\asqrt[2] ), .A2(new_n19782_), .A3(new_n22524_), .A4(new_n22944_), .ZN(new_n23232_));
  XOR2_X1    g23039(.A1(new_n23232_), .A2(new_n22538_), .Z(new_n23233_));
  NAND2_X1   g23040(.A1(new_n23233_), .A2(new_n19100_), .ZN(new_n23234_));
  INV_X1     g23041(.I(new_n23234_), .ZN(new_n23235_));
  OAI21_X1   g23042(.A1(new_n23231_), .A2(new_n19782_), .B(new_n23235_), .ZN(new_n23236_));
  NAND2_X1   g23043(.A1(new_n23236_), .A2(new_n23230_), .ZN(new_n23237_));
  OAI22_X1   g23044(.A1(new_n23231_), .A2(new_n19782_), .B1(new_n23229_), .B2(new_n23223_), .ZN(new_n23238_));
  NOR4_X1    g23045(.A1(new_n23158_), .A2(\asqrt[8] ), .A3(new_n22532_), .A4(new_n22951_), .ZN(new_n23239_));
  XOR2_X1    g23046(.A1(new_n23239_), .A2(new_n22539_), .Z(new_n23240_));
  NAND2_X1   g23047(.A1(new_n23240_), .A2(new_n18495_), .ZN(new_n23241_));
  AOI21_X1   g23048(.A1(new_n23238_), .A2(\asqrt[8] ), .B(new_n23241_), .ZN(new_n23242_));
  NOR2_X1    g23049(.A1(new_n23242_), .A2(new_n23237_), .ZN(new_n23243_));
  AOI22_X1   g23050(.A1(new_n23238_), .A2(\asqrt[8] ), .B1(new_n23236_), .B2(new_n23230_), .ZN(new_n23244_));
  NOR2_X1    g23051(.A1(new_n22954_), .A2(new_n18495_), .ZN(new_n23245_));
  NOR4_X1    g23052(.A1(new_n23158_), .A2(\asqrt[9] ), .A3(new_n22542_), .A4(new_n22548_), .ZN(new_n23246_));
  XNOR2_X1   g23053(.A1(new_n23246_), .A2(new_n23245_), .ZN(new_n23247_));
  NAND2_X1   g23054(.A1(new_n23247_), .A2(new_n17893_), .ZN(new_n23248_));
  INV_X1     g23055(.I(new_n23248_), .ZN(new_n23249_));
  OAI21_X1   g23056(.A1(new_n23244_), .A2(new_n18495_), .B(new_n23249_), .ZN(new_n23250_));
  NAND2_X1   g23057(.A1(new_n23250_), .A2(new_n23243_), .ZN(new_n23251_));
  OAI22_X1   g23058(.A1(new_n23244_), .A2(new_n18495_), .B1(new_n23242_), .B2(new_n23237_), .ZN(new_n23252_));
  NAND2_X1   g23059(.A1(new_n22958_), .A2(\asqrt[10] ), .ZN(new_n23253_));
  NOR4_X1    g23060(.A1(new_n23158_), .A2(\asqrt[10] ), .A3(new_n22551_), .A4(new_n22958_), .ZN(new_n23254_));
  XOR2_X1    g23061(.A1(new_n23254_), .A2(new_n23253_), .Z(new_n23255_));
  NAND2_X1   g23062(.A1(new_n23255_), .A2(new_n17271_), .ZN(new_n23256_));
  AOI21_X1   g23063(.A1(new_n23252_), .A2(\asqrt[10] ), .B(new_n23256_), .ZN(new_n23257_));
  NOR2_X1    g23064(.A1(new_n23257_), .A2(new_n23251_), .ZN(new_n23258_));
  AOI22_X1   g23065(.A1(new_n23252_), .A2(\asqrt[10] ), .B1(new_n23250_), .B2(new_n23243_), .ZN(new_n23259_));
  NAND2_X1   g23066(.A1(new_n22562_), .A2(\asqrt[11] ), .ZN(new_n23260_));
  NOR4_X1    g23067(.A1(new_n23158_), .A2(\asqrt[11] ), .A3(new_n22557_), .A4(new_n22562_), .ZN(new_n23261_));
  XOR2_X1    g23068(.A1(new_n23261_), .A2(new_n23260_), .Z(new_n23262_));
  NAND2_X1   g23069(.A1(new_n23262_), .A2(new_n16619_), .ZN(new_n23263_));
  INV_X1     g23070(.I(new_n23263_), .ZN(new_n23264_));
  OAI21_X1   g23071(.A1(new_n23259_), .A2(new_n17271_), .B(new_n23264_), .ZN(new_n23265_));
  NAND2_X1   g23072(.A1(new_n23265_), .A2(new_n23258_), .ZN(new_n23266_));
  OAI22_X1   g23073(.A1(new_n23259_), .A2(new_n17271_), .B1(new_n23257_), .B2(new_n23251_), .ZN(new_n23267_));
  NOR4_X1    g23074(.A1(new_n23158_), .A2(\asqrt[12] ), .A3(new_n22564_), .A4(new_n22965_), .ZN(new_n23268_));
  AOI21_X1   g23075(.A1(new_n23260_), .A2(new_n22561_), .B(new_n16619_), .ZN(new_n23269_));
  NOR2_X1    g23076(.A1(new_n23268_), .A2(new_n23269_), .ZN(new_n23270_));
  NAND2_X1   g23077(.A1(new_n23270_), .A2(new_n16060_), .ZN(new_n23271_));
  AOI21_X1   g23078(.A1(new_n23267_), .A2(\asqrt[12] ), .B(new_n23271_), .ZN(new_n23272_));
  NOR2_X1    g23079(.A1(new_n23272_), .A2(new_n23266_), .ZN(new_n23273_));
  AOI22_X1   g23080(.A1(new_n23267_), .A2(\asqrt[12] ), .B1(new_n23265_), .B2(new_n23258_), .ZN(new_n23274_));
  NAND2_X1   g23081(.A1(new_n22575_), .A2(\asqrt[13] ), .ZN(new_n23275_));
  NOR4_X1    g23082(.A1(new_n23158_), .A2(\asqrt[13] ), .A3(new_n22570_), .A4(new_n22575_), .ZN(new_n23276_));
  XOR2_X1    g23083(.A1(new_n23276_), .A2(new_n23275_), .Z(new_n23277_));
  NAND2_X1   g23084(.A1(new_n23277_), .A2(new_n15447_), .ZN(new_n23278_));
  INV_X1     g23085(.I(new_n23278_), .ZN(new_n23279_));
  OAI21_X1   g23086(.A1(new_n23274_), .A2(new_n16060_), .B(new_n23279_), .ZN(new_n23280_));
  NAND2_X1   g23087(.A1(new_n23280_), .A2(new_n23273_), .ZN(new_n23281_));
  OAI22_X1   g23088(.A1(new_n23274_), .A2(new_n16060_), .B1(new_n23272_), .B2(new_n23266_), .ZN(new_n23282_));
  NOR4_X1    g23089(.A1(new_n23158_), .A2(\asqrt[14] ), .A3(new_n22578_), .A4(new_n22972_), .ZN(new_n23283_));
  AOI21_X1   g23090(.A1(new_n23275_), .A2(new_n22574_), .B(new_n15447_), .ZN(new_n23284_));
  NOR2_X1    g23091(.A1(new_n23283_), .A2(new_n23284_), .ZN(new_n23285_));
  NAND2_X1   g23092(.A1(new_n23285_), .A2(new_n14871_), .ZN(new_n23286_));
  AOI21_X1   g23093(.A1(new_n23282_), .A2(\asqrt[14] ), .B(new_n23286_), .ZN(new_n23287_));
  NOR2_X1    g23094(.A1(new_n23287_), .A2(new_n23281_), .ZN(new_n23288_));
  AOI22_X1   g23095(.A1(new_n23282_), .A2(\asqrt[14] ), .B1(new_n23280_), .B2(new_n23273_), .ZN(new_n23289_));
  NAND2_X1   g23096(.A1(new_n22590_), .A2(\asqrt[15] ), .ZN(new_n23290_));
  NOR4_X1    g23097(.A1(new_n23158_), .A2(\asqrt[15] ), .A3(new_n22585_), .A4(new_n22590_), .ZN(new_n23291_));
  XOR2_X1    g23098(.A1(new_n23291_), .A2(new_n23290_), .Z(new_n23292_));
  NAND2_X1   g23099(.A1(new_n23292_), .A2(new_n14273_), .ZN(new_n23293_));
  INV_X1     g23100(.I(new_n23293_), .ZN(new_n23294_));
  OAI21_X1   g23101(.A1(new_n23289_), .A2(new_n14871_), .B(new_n23294_), .ZN(new_n23295_));
  NAND2_X1   g23102(.A1(new_n23295_), .A2(new_n23288_), .ZN(new_n23296_));
  OAI22_X1   g23103(.A1(new_n23289_), .A2(new_n14871_), .B1(new_n23287_), .B2(new_n23281_), .ZN(new_n23297_));
  NOR4_X1    g23104(.A1(new_n23158_), .A2(\asqrt[16] ), .A3(new_n22593_), .A4(new_n22979_), .ZN(new_n23298_));
  AOI21_X1   g23105(.A1(new_n23290_), .A2(new_n22589_), .B(new_n14273_), .ZN(new_n23299_));
  NOR2_X1    g23106(.A1(new_n23298_), .A2(new_n23299_), .ZN(new_n23300_));
  NAND2_X1   g23107(.A1(new_n23300_), .A2(new_n13760_), .ZN(new_n23301_));
  AOI21_X1   g23108(.A1(new_n23297_), .A2(\asqrt[16] ), .B(new_n23301_), .ZN(new_n23302_));
  NOR2_X1    g23109(.A1(new_n23302_), .A2(new_n23296_), .ZN(new_n23303_));
  AOI22_X1   g23110(.A1(new_n23297_), .A2(\asqrt[16] ), .B1(new_n23295_), .B2(new_n23288_), .ZN(new_n23304_));
  NAND2_X1   g23111(.A1(new_n22605_), .A2(\asqrt[17] ), .ZN(new_n23305_));
  NOR4_X1    g23112(.A1(new_n23158_), .A2(\asqrt[17] ), .A3(new_n22600_), .A4(new_n22605_), .ZN(new_n23306_));
  XOR2_X1    g23113(.A1(new_n23306_), .A2(new_n23305_), .Z(new_n23307_));
  NAND2_X1   g23114(.A1(new_n23307_), .A2(new_n13192_), .ZN(new_n23308_));
  INV_X1     g23115(.I(new_n23308_), .ZN(new_n23309_));
  OAI21_X1   g23116(.A1(new_n23304_), .A2(new_n13760_), .B(new_n23309_), .ZN(new_n23310_));
  NAND2_X1   g23117(.A1(new_n23310_), .A2(new_n23303_), .ZN(new_n23311_));
  OAI22_X1   g23118(.A1(new_n23304_), .A2(new_n13760_), .B1(new_n23302_), .B2(new_n23296_), .ZN(new_n23312_));
  NOR4_X1    g23119(.A1(new_n23158_), .A2(\asqrt[18] ), .A3(new_n22608_), .A4(new_n22986_), .ZN(new_n23313_));
  AOI21_X1   g23120(.A1(new_n23305_), .A2(new_n22604_), .B(new_n13192_), .ZN(new_n23314_));
  NOR2_X1    g23121(.A1(new_n23313_), .A2(new_n23314_), .ZN(new_n23315_));
  NAND2_X1   g23122(.A1(new_n23315_), .A2(new_n12657_), .ZN(new_n23316_));
  AOI21_X1   g23123(.A1(new_n23312_), .A2(\asqrt[18] ), .B(new_n23316_), .ZN(new_n23317_));
  NOR2_X1    g23124(.A1(new_n23317_), .A2(new_n23311_), .ZN(new_n23318_));
  AOI22_X1   g23125(.A1(new_n23312_), .A2(\asqrt[18] ), .B1(new_n23310_), .B2(new_n23303_), .ZN(new_n23319_));
  NAND2_X1   g23126(.A1(new_n22620_), .A2(\asqrt[19] ), .ZN(new_n23320_));
  NOR4_X1    g23127(.A1(new_n23158_), .A2(\asqrt[19] ), .A3(new_n22615_), .A4(new_n22620_), .ZN(new_n23321_));
  XOR2_X1    g23128(.A1(new_n23321_), .A2(new_n23320_), .Z(new_n23322_));
  NAND2_X1   g23129(.A1(new_n23322_), .A2(new_n12101_), .ZN(new_n23323_));
  INV_X1     g23130(.I(new_n23323_), .ZN(new_n23324_));
  OAI21_X1   g23131(.A1(new_n23319_), .A2(new_n12657_), .B(new_n23324_), .ZN(new_n23325_));
  NAND2_X1   g23132(.A1(new_n23325_), .A2(new_n23318_), .ZN(new_n23326_));
  OAI22_X1   g23133(.A1(new_n23319_), .A2(new_n12657_), .B1(new_n23317_), .B2(new_n23311_), .ZN(new_n23327_));
  NOR4_X1    g23134(.A1(new_n23158_), .A2(\asqrt[20] ), .A3(new_n22623_), .A4(new_n22993_), .ZN(new_n23328_));
  AOI21_X1   g23135(.A1(new_n23320_), .A2(new_n22619_), .B(new_n12101_), .ZN(new_n23329_));
  NOR2_X1    g23136(.A1(new_n23328_), .A2(new_n23329_), .ZN(new_n23330_));
  NAND2_X1   g23137(.A1(new_n23330_), .A2(new_n11631_), .ZN(new_n23331_));
  AOI21_X1   g23138(.A1(new_n23327_), .A2(\asqrt[20] ), .B(new_n23331_), .ZN(new_n23332_));
  NOR2_X1    g23139(.A1(new_n23332_), .A2(new_n23326_), .ZN(new_n23333_));
  AOI22_X1   g23140(.A1(new_n23327_), .A2(\asqrt[20] ), .B1(new_n23325_), .B2(new_n23318_), .ZN(new_n23334_));
  NAND2_X1   g23141(.A1(new_n22635_), .A2(\asqrt[21] ), .ZN(new_n23335_));
  NOR4_X1    g23142(.A1(new_n23158_), .A2(\asqrt[21] ), .A3(new_n22630_), .A4(new_n22635_), .ZN(new_n23336_));
  XOR2_X1    g23143(.A1(new_n23336_), .A2(new_n23335_), .Z(new_n23337_));
  NAND2_X1   g23144(.A1(new_n23337_), .A2(new_n11105_), .ZN(new_n23338_));
  INV_X1     g23145(.I(new_n23338_), .ZN(new_n23339_));
  OAI21_X1   g23146(.A1(new_n23334_), .A2(new_n11631_), .B(new_n23339_), .ZN(new_n23340_));
  NAND2_X1   g23147(.A1(new_n23340_), .A2(new_n23333_), .ZN(new_n23341_));
  OAI22_X1   g23148(.A1(new_n23334_), .A2(new_n11631_), .B1(new_n23332_), .B2(new_n23326_), .ZN(new_n23342_));
  NAND2_X1   g23149(.A1(new_n23000_), .A2(\asqrt[22] ), .ZN(new_n23343_));
  NOR4_X1    g23150(.A1(new_n23158_), .A2(\asqrt[22] ), .A3(new_n22638_), .A4(new_n23000_), .ZN(new_n23344_));
  XOR2_X1    g23151(.A1(new_n23344_), .A2(new_n23343_), .Z(new_n23345_));
  NAND2_X1   g23152(.A1(new_n23345_), .A2(new_n10614_), .ZN(new_n23346_));
  AOI21_X1   g23153(.A1(new_n23342_), .A2(\asqrt[22] ), .B(new_n23346_), .ZN(new_n23347_));
  NOR2_X1    g23154(.A1(new_n23347_), .A2(new_n23341_), .ZN(new_n23348_));
  AOI22_X1   g23155(.A1(new_n23342_), .A2(\asqrt[22] ), .B1(new_n23340_), .B2(new_n23333_), .ZN(new_n23349_));
  NOR4_X1    g23156(.A1(new_n23158_), .A2(\asqrt[23] ), .A3(new_n22645_), .A4(new_n22650_), .ZN(new_n23350_));
  AOI21_X1   g23157(.A1(new_n23343_), .A2(new_n22999_), .B(new_n10614_), .ZN(new_n23351_));
  NOR2_X1    g23158(.A1(new_n23350_), .A2(new_n23351_), .ZN(new_n23352_));
  NAND2_X1   g23159(.A1(new_n23352_), .A2(new_n10104_), .ZN(new_n23353_));
  INV_X1     g23160(.I(new_n23353_), .ZN(new_n23354_));
  OAI21_X1   g23161(.A1(new_n23349_), .A2(new_n10614_), .B(new_n23354_), .ZN(new_n23355_));
  NAND2_X1   g23162(.A1(new_n23355_), .A2(new_n23348_), .ZN(new_n23356_));
  OAI22_X1   g23163(.A1(new_n23349_), .A2(new_n10614_), .B1(new_n23347_), .B2(new_n23341_), .ZN(new_n23357_));
  NAND2_X1   g23164(.A1(new_n23007_), .A2(\asqrt[24] ), .ZN(new_n23358_));
  NOR4_X1    g23165(.A1(new_n23158_), .A2(\asqrt[24] ), .A3(new_n22653_), .A4(new_n23007_), .ZN(new_n23359_));
  XOR2_X1    g23166(.A1(new_n23359_), .A2(new_n23358_), .Z(new_n23360_));
  NAND2_X1   g23167(.A1(new_n23360_), .A2(new_n9672_), .ZN(new_n23361_));
  AOI21_X1   g23168(.A1(new_n23357_), .A2(\asqrt[24] ), .B(new_n23361_), .ZN(new_n23362_));
  NOR2_X1    g23169(.A1(new_n23362_), .A2(new_n23356_), .ZN(new_n23363_));
  AOI22_X1   g23170(.A1(new_n23357_), .A2(\asqrt[24] ), .B1(new_n23355_), .B2(new_n23348_), .ZN(new_n23364_));
  NOR4_X1    g23171(.A1(new_n23158_), .A2(\asqrt[25] ), .A3(new_n22660_), .A4(new_n22665_), .ZN(new_n23365_));
  AOI21_X1   g23172(.A1(new_n23358_), .A2(new_n23006_), .B(new_n9672_), .ZN(new_n23366_));
  NOR2_X1    g23173(.A1(new_n23365_), .A2(new_n23366_), .ZN(new_n23367_));
  NAND2_X1   g23174(.A1(new_n23367_), .A2(new_n9212_), .ZN(new_n23368_));
  INV_X1     g23175(.I(new_n23368_), .ZN(new_n23369_));
  OAI21_X1   g23176(.A1(new_n23364_), .A2(new_n9672_), .B(new_n23369_), .ZN(new_n23370_));
  NAND2_X1   g23177(.A1(new_n23370_), .A2(new_n23363_), .ZN(new_n23371_));
  OAI22_X1   g23178(.A1(new_n23364_), .A2(new_n9672_), .B1(new_n23362_), .B2(new_n23356_), .ZN(new_n23372_));
  NAND2_X1   g23179(.A1(new_n23014_), .A2(\asqrt[26] ), .ZN(new_n23373_));
  NOR4_X1    g23180(.A1(new_n23158_), .A2(\asqrt[26] ), .A3(new_n22668_), .A4(new_n23014_), .ZN(new_n23374_));
  XOR2_X1    g23181(.A1(new_n23374_), .A2(new_n23373_), .Z(new_n23375_));
  NAND2_X1   g23182(.A1(new_n23375_), .A2(new_n8763_), .ZN(new_n23376_));
  AOI21_X1   g23183(.A1(new_n23372_), .A2(\asqrt[26] ), .B(new_n23376_), .ZN(new_n23377_));
  NOR2_X1    g23184(.A1(new_n23377_), .A2(new_n23371_), .ZN(new_n23378_));
  AOI22_X1   g23185(.A1(new_n23372_), .A2(\asqrt[26] ), .B1(new_n23370_), .B2(new_n23363_), .ZN(new_n23379_));
  NAND2_X1   g23186(.A1(new_n22680_), .A2(\asqrt[27] ), .ZN(new_n23380_));
  NOR4_X1    g23187(.A1(new_n23158_), .A2(\asqrt[27] ), .A3(new_n22675_), .A4(new_n22680_), .ZN(new_n23381_));
  XOR2_X1    g23188(.A1(new_n23381_), .A2(new_n23380_), .Z(new_n23382_));
  NAND2_X1   g23189(.A1(new_n23382_), .A2(new_n8319_), .ZN(new_n23383_));
  INV_X1     g23190(.I(new_n23383_), .ZN(new_n23384_));
  OAI21_X1   g23191(.A1(new_n23379_), .A2(new_n8763_), .B(new_n23384_), .ZN(new_n23385_));
  NAND2_X1   g23192(.A1(new_n23385_), .A2(new_n23378_), .ZN(new_n23386_));
  OAI22_X1   g23193(.A1(new_n23379_), .A2(new_n8763_), .B1(new_n23377_), .B2(new_n23371_), .ZN(new_n23387_));
  NOR4_X1    g23194(.A1(new_n23158_), .A2(\asqrt[28] ), .A3(new_n22683_), .A4(new_n23021_), .ZN(new_n23388_));
  AOI21_X1   g23195(.A1(new_n23380_), .A2(new_n22679_), .B(new_n8319_), .ZN(new_n23389_));
  NOR2_X1    g23196(.A1(new_n23388_), .A2(new_n23389_), .ZN(new_n23390_));
  NAND2_X1   g23197(.A1(new_n23390_), .A2(new_n7931_), .ZN(new_n23391_));
  AOI21_X1   g23198(.A1(new_n23387_), .A2(\asqrt[28] ), .B(new_n23391_), .ZN(new_n23392_));
  NOR2_X1    g23199(.A1(new_n23392_), .A2(new_n23386_), .ZN(new_n23393_));
  AOI22_X1   g23200(.A1(new_n23387_), .A2(\asqrt[28] ), .B1(new_n23385_), .B2(new_n23378_), .ZN(new_n23394_));
  NAND2_X1   g23201(.A1(new_n22695_), .A2(\asqrt[29] ), .ZN(new_n23395_));
  NOR4_X1    g23202(.A1(new_n23158_), .A2(\asqrt[29] ), .A3(new_n22690_), .A4(new_n22695_), .ZN(new_n23396_));
  XOR2_X1    g23203(.A1(new_n23396_), .A2(new_n23395_), .Z(new_n23397_));
  NAND2_X1   g23204(.A1(new_n23397_), .A2(new_n7517_), .ZN(new_n23398_));
  INV_X1     g23205(.I(new_n23398_), .ZN(new_n23399_));
  OAI21_X1   g23206(.A1(new_n23394_), .A2(new_n7931_), .B(new_n23399_), .ZN(new_n23400_));
  NAND2_X1   g23207(.A1(new_n23400_), .A2(new_n23393_), .ZN(new_n23401_));
  OAI22_X1   g23208(.A1(new_n23394_), .A2(new_n7931_), .B1(new_n23392_), .B2(new_n23386_), .ZN(new_n23402_));
  NOR4_X1    g23209(.A1(new_n23158_), .A2(\asqrt[30] ), .A3(new_n22698_), .A4(new_n23028_), .ZN(new_n23403_));
  AOI21_X1   g23210(.A1(new_n23395_), .A2(new_n22694_), .B(new_n7517_), .ZN(new_n23404_));
  NOR2_X1    g23211(.A1(new_n23403_), .A2(new_n23404_), .ZN(new_n23405_));
  NAND2_X1   g23212(.A1(new_n23405_), .A2(new_n7110_), .ZN(new_n23406_));
  AOI21_X1   g23213(.A1(new_n23402_), .A2(\asqrt[30] ), .B(new_n23406_), .ZN(new_n23407_));
  NOR2_X1    g23214(.A1(new_n23407_), .A2(new_n23401_), .ZN(new_n23408_));
  AOI22_X1   g23215(.A1(new_n23402_), .A2(\asqrt[30] ), .B1(new_n23400_), .B2(new_n23393_), .ZN(new_n23409_));
  NAND2_X1   g23216(.A1(new_n22710_), .A2(\asqrt[31] ), .ZN(new_n23410_));
  NOR4_X1    g23217(.A1(new_n23158_), .A2(\asqrt[31] ), .A3(new_n22705_), .A4(new_n22710_), .ZN(new_n23411_));
  XOR2_X1    g23218(.A1(new_n23411_), .A2(new_n23410_), .Z(new_n23412_));
  NAND2_X1   g23219(.A1(new_n23412_), .A2(new_n6708_), .ZN(new_n23413_));
  INV_X1     g23220(.I(new_n23413_), .ZN(new_n23414_));
  OAI21_X1   g23221(.A1(new_n23409_), .A2(new_n7110_), .B(new_n23414_), .ZN(new_n23415_));
  NAND2_X1   g23222(.A1(new_n23415_), .A2(new_n23408_), .ZN(new_n23416_));
  OAI22_X1   g23223(.A1(new_n23409_), .A2(new_n7110_), .B1(new_n23407_), .B2(new_n23401_), .ZN(new_n23417_));
  NAND2_X1   g23224(.A1(new_n23035_), .A2(\asqrt[32] ), .ZN(new_n23418_));
  NOR4_X1    g23225(.A1(new_n23158_), .A2(\asqrt[32] ), .A3(new_n22713_), .A4(new_n23035_), .ZN(new_n23419_));
  XOR2_X1    g23226(.A1(new_n23419_), .A2(new_n23418_), .Z(new_n23420_));
  NAND2_X1   g23227(.A1(new_n23420_), .A2(new_n6365_), .ZN(new_n23421_));
  AOI21_X1   g23228(.A1(new_n23417_), .A2(\asqrt[32] ), .B(new_n23421_), .ZN(new_n23422_));
  NOR2_X1    g23229(.A1(new_n23422_), .A2(new_n23416_), .ZN(new_n23423_));
  AOI22_X1   g23230(.A1(new_n23417_), .A2(\asqrt[32] ), .B1(new_n23415_), .B2(new_n23408_), .ZN(new_n23424_));
  NOR4_X1    g23231(.A1(new_n23158_), .A2(\asqrt[33] ), .A3(new_n22720_), .A4(new_n22725_), .ZN(new_n23425_));
  AOI21_X1   g23232(.A1(new_n23418_), .A2(new_n23034_), .B(new_n6365_), .ZN(new_n23426_));
  NOR2_X1    g23233(.A1(new_n23425_), .A2(new_n23426_), .ZN(new_n23427_));
  NAND2_X1   g23234(.A1(new_n23427_), .A2(new_n5991_), .ZN(new_n23428_));
  INV_X1     g23235(.I(new_n23428_), .ZN(new_n23429_));
  OAI21_X1   g23236(.A1(new_n23424_), .A2(new_n6365_), .B(new_n23429_), .ZN(new_n23430_));
  NAND2_X1   g23237(.A1(new_n23430_), .A2(new_n23423_), .ZN(new_n23431_));
  OAI22_X1   g23238(.A1(new_n23424_), .A2(new_n6365_), .B1(new_n23422_), .B2(new_n23416_), .ZN(new_n23432_));
  NAND2_X1   g23239(.A1(new_n23042_), .A2(\asqrt[34] ), .ZN(new_n23433_));
  NOR4_X1    g23240(.A1(new_n23158_), .A2(\asqrt[34] ), .A3(new_n22728_), .A4(new_n23042_), .ZN(new_n23434_));
  XOR2_X1    g23241(.A1(new_n23434_), .A2(new_n23433_), .Z(new_n23435_));
  NAND2_X1   g23242(.A1(new_n23435_), .A2(new_n5626_), .ZN(new_n23436_));
  AOI21_X1   g23243(.A1(new_n23432_), .A2(\asqrt[34] ), .B(new_n23436_), .ZN(new_n23437_));
  NOR2_X1    g23244(.A1(new_n23437_), .A2(new_n23431_), .ZN(new_n23438_));
  AOI22_X1   g23245(.A1(new_n23432_), .A2(\asqrt[34] ), .B1(new_n23430_), .B2(new_n23423_), .ZN(new_n23439_));
  NOR4_X1    g23246(.A1(new_n23158_), .A2(\asqrt[35] ), .A3(new_n22735_), .A4(new_n22740_), .ZN(new_n23440_));
  AOI21_X1   g23247(.A1(new_n23433_), .A2(new_n23041_), .B(new_n5626_), .ZN(new_n23441_));
  NOR2_X1    g23248(.A1(new_n23440_), .A2(new_n23441_), .ZN(new_n23442_));
  NAND2_X1   g23249(.A1(new_n23442_), .A2(new_n5273_), .ZN(new_n23443_));
  INV_X1     g23250(.I(new_n23443_), .ZN(new_n23444_));
  OAI21_X1   g23251(.A1(new_n23439_), .A2(new_n5626_), .B(new_n23444_), .ZN(new_n23445_));
  NAND2_X1   g23252(.A1(new_n23445_), .A2(new_n23438_), .ZN(new_n23446_));
  OAI22_X1   g23253(.A1(new_n23439_), .A2(new_n5626_), .B1(new_n23437_), .B2(new_n23431_), .ZN(new_n23447_));
  NAND2_X1   g23254(.A1(new_n23049_), .A2(\asqrt[36] ), .ZN(new_n23448_));
  NOR4_X1    g23255(.A1(new_n23158_), .A2(\asqrt[36] ), .A3(new_n22743_), .A4(new_n23049_), .ZN(new_n23449_));
  XOR2_X1    g23256(.A1(new_n23449_), .A2(new_n23448_), .Z(new_n23450_));
  NAND2_X1   g23257(.A1(new_n23450_), .A2(new_n4973_), .ZN(new_n23451_));
  AOI21_X1   g23258(.A1(new_n23447_), .A2(\asqrt[36] ), .B(new_n23451_), .ZN(new_n23452_));
  NOR2_X1    g23259(.A1(new_n23452_), .A2(new_n23446_), .ZN(new_n23453_));
  AOI22_X1   g23260(.A1(new_n23447_), .A2(\asqrt[36] ), .B1(new_n23445_), .B2(new_n23438_), .ZN(new_n23454_));
  NOR4_X1    g23261(.A1(new_n23158_), .A2(\asqrt[37] ), .A3(new_n22750_), .A4(new_n22755_), .ZN(new_n23455_));
  AOI21_X1   g23262(.A1(new_n23448_), .A2(new_n23048_), .B(new_n4973_), .ZN(new_n23456_));
  NOR2_X1    g23263(.A1(new_n23455_), .A2(new_n23456_), .ZN(new_n23457_));
  NAND2_X1   g23264(.A1(new_n23457_), .A2(new_n4645_), .ZN(new_n23458_));
  INV_X1     g23265(.I(new_n23458_), .ZN(new_n23459_));
  OAI21_X1   g23266(.A1(new_n23454_), .A2(new_n4973_), .B(new_n23459_), .ZN(new_n23460_));
  NAND2_X1   g23267(.A1(new_n23460_), .A2(new_n23453_), .ZN(new_n23461_));
  OAI22_X1   g23268(.A1(new_n23454_), .A2(new_n4973_), .B1(new_n23452_), .B2(new_n23446_), .ZN(new_n23462_));
  NAND2_X1   g23269(.A1(new_n23056_), .A2(\asqrt[38] ), .ZN(new_n23463_));
  NOR4_X1    g23270(.A1(new_n23158_), .A2(\asqrt[38] ), .A3(new_n22758_), .A4(new_n23056_), .ZN(new_n23464_));
  XOR2_X1    g23271(.A1(new_n23464_), .A2(new_n23463_), .Z(new_n23465_));
  NAND2_X1   g23272(.A1(new_n23465_), .A2(new_n4330_), .ZN(new_n23466_));
  AOI21_X1   g23273(.A1(new_n23462_), .A2(\asqrt[38] ), .B(new_n23466_), .ZN(new_n23467_));
  NOR2_X1    g23274(.A1(new_n23467_), .A2(new_n23461_), .ZN(new_n23468_));
  AOI22_X1   g23275(.A1(new_n23462_), .A2(\asqrt[38] ), .B1(new_n23460_), .B2(new_n23453_), .ZN(new_n23469_));
  NAND2_X1   g23276(.A1(new_n22770_), .A2(\asqrt[39] ), .ZN(new_n23470_));
  NOR4_X1    g23277(.A1(new_n23158_), .A2(\asqrt[39] ), .A3(new_n22765_), .A4(new_n22770_), .ZN(new_n23471_));
  XOR2_X1    g23278(.A1(new_n23471_), .A2(new_n23470_), .Z(new_n23472_));
  NAND2_X1   g23279(.A1(new_n23472_), .A2(new_n4018_), .ZN(new_n23473_));
  INV_X1     g23280(.I(new_n23473_), .ZN(new_n23474_));
  OAI21_X1   g23281(.A1(new_n23469_), .A2(new_n4330_), .B(new_n23474_), .ZN(new_n23475_));
  NAND2_X1   g23282(.A1(new_n23475_), .A2(new_n23468_), .ZN(new_n23476_));
  OAI22_X1   g23283(.A1(new_n23469_), .A2(new_n4330_), .B1(new_n23467_), .B2(new_n23461_), .ZN(new_n23477_));
  NOR4_X1    g23284(.A1(new_n23158_), .A2(\asqrt[40] ), .A3(new_n22773_), .A4(new_n23063_), .ZN(new_n23478_));
  AOI21_X1   g23285(.A1(new_n23470_), .A2(new_n22769_), .B(new_n4018_), .ZN(new_n23479_));
  NOR2_X1    g23286(.A1(new_n23478_), .A2(new_n23479_), .ZN(new_n23480_));
  NAND2_X1   g23287(.A1(new_n23480_), .A2(new_n3760_), .ZN(new_n23481_));
  AOI21_X1   g23288(.A1(new_n23477_), .A2(\asqrt[40] ), .B(new_n23481_), .ZN(new_n23482_));
  NOR2_X1    g23289(.A1(new_n23482_), .A2(new_n23476_), .ZN(new_n23483_));
  AOI22_X1   g23290(.A1(new_n23477_), .A2(\asqrt[40] ), .B1(new_n23475_), .B2(new_n23468_), .ZN(new_n23484_));
  NAND2_X1   g23291(.A1(new_n22785_), .A2(\asqrt[41] ), .ZN(new_n23485_));
  NOR4_X1    g23292(.A1(new_n23158_), .A2(\asqrt[41] ), .A3(new_n22780_), .A4(new_n22785_), .ZN(new_n23486_));
  XOR2_X1    g23293(.A1(new_n23486_), .A2(new_n23485_), .Z(new_n23487_));
  NAND2_X1   g23294(.A1(new_n23487_), .A2(new_n3481_), .ZN(new_n23488_));
  INV_X1     g23295(.I(new_n23488_), .ZN(new_n23489_));
  OAI21_X1   g23296(.A1(new_n23484_), .A2(new_n3760_), .B(new_n23489_), .ZN(new_n23490_));
  NAND2_X1   g23297(.A1(new_n23490_), .A2(new_n23483_), .ZN(new_n23491_));
  OAI22_X1   g23298(.A1(new_n23484_), .A2(new_n3760_), .B1(new_n23482_), .B2(new_n23476_), .ZN(new_n23492_));
  NOR4_X1    g23299(.A1(new_n23158_), .A2(\asqrt[42] ), .A3(new_n22788_), .A4(new_n23070_), .ZN(new_n23493_));
  AOI21_X1   g23300(.A1(new_n23485_), .A2(new_n22784_), .B(new_n3481_), .ZN(new_n23494_));
  NOR2_X1    g23301(.A1(new_n23493_), .A2(new_n23494_), .ZN(new_n23495_));
  NAND2_X1   g23302(.A1(new_n23495_), .A2(new_n3208_), .ZN(new_n23496_));
  AOI21_X1   g23303(.A1(new_n23492_), .A2(\asqrt[42] ), .B(new_n23496_), .ZN(new_n23497_));
  NOR2_X1    g23304(.A1(new_n23497_), .A2(new_n23491_), .ZN(new_n23498_));
  AOI22_X1   g23305(.A1(new_n23492_), .A2(\asqrt[42] ), .B1(new_n23490_), .B2(new_n23483_), .ZN(new_n23499_));
  NAND2_X1   g23306(.A1(new_n22800_), .A2(\asqrt[43] ), .ZN(new_n23500_));
  NOR4_X1    g23307(.A1(new_n23158_), .A2(\asqrt[43] ), .A3(new_n22795_), .A4(new_n22800_), .ZN(new_n23501_));
  XOR2_X1    g23308(.A1(new_n23501_), .A2(new_n23500_), .Z(new_n23502_));
  NAND2_X1   g23309(.A1(new_n23502_), .A2(new_n2941_), .ZN(new_n23503_));
  INV_X1     g23310(.I(new_n23503_), .ZN(new_n23504_));
  OAI21_X1   g23311(.A1(new_n23499_), .A2(new_n3208_), .B(new_n23504_), .ZN(new_n23505_));
  NAND2_X1   g23312(.A1(new_n23505_), .A2(new_n23498_), .ZN(new_n23506_));
  OAI22_X1   g23313(.A1(new_n23499_), .A2(new_n3208_), .B1(new_n23497_), .B2(new_n23491_), .ZN(new_n23507_));
  NAND2_X1   g23314(.A1(new_n23077_), .A2(\asqrt[44] ), .ZN(new_n23508_));
  NOR4_X1    g23315(.A1(new_n23158_), .A2(\asqrt[44] ), .A3(new_n22803_), .A4(new_n23077_), .ZN(new_n23509_));
  XOR2_X1    g23316(.A1(new_n23509_), .A2(new_n23508_), .Z(new_n23510_));
  NAND2_X1   g23317(.A1(new_n23510_), .A2(new_n2728_), .ZN(new_n23511_));
  AOI21_X1   g23318(.A1(new_n23507_), .A2(\asqrt[44] ), .B(new_n23511_), .ZN(new_n23512_));
  NOR2_X1    g23319(.A1(new_n23512_), .A2(new_n23506_), .ZN(new_n23513_));
  AOI22_X1   g23320(.A1(new_n23507_), .A2(\asqrt[44] ), .B1(new_n23505_), .B2(new_n23498_), .ZN(new_n23514_));
  NOR4_X1    g23321(.A1(new_n23158_), .A2(\asqrt[45] ), .A3(new_n22810_), .A4(new_n22815_), .ZN(new_n23515_));
  AOI21_X1   g23322(.A1(new_n23508_), .A2(new_n23076_), .B(new_n2728_), .ZN(new_n23516_));
  NOR2_X1    g23323(.A1(new_n23515_), .A2(new_n23516_), .ZN(new_n23517_));
  NAND2_X1   g23324(.A1(new_n23517_), .A2(new_n2488_), .ZN(new_n23518_));
  INV_X1     g23325(.I(new_n23518_), .ZN(new_n23519_));
  OAI21_X1   g23326(.A1(new_n23514_), .A2(new_n2728_), .B(new_n23519_), .ZN(new_n23520_));
  NAND2_X1   g23327(.A1(new_n23520_), .A2(new_n23513_), .ZN(new_n23521_));
  OAI22_X1   g23328(.A1(new_n23514_), .A2(new_n2728_), .B1(new_n23512_), .B2(new_n23506_), .ZN(new_n23522_));
  NAND2_X1   g23329(.A1(new_n23084_), .A2(\asqrt[46] ), .ZN(new_n23523_));
  NOR4_X1    g23330(.A1(new_n23158_), .A2(\asqrt[46] ), .A3(new_n22818_), .A4(new_n23084_), .ZN(new_n23524_));
  XOR2_X1    g23331(.A1(new_n23524_), .A2(new_n23523_), .Z(new_n23525_));
  NAND2_X1   g23332(.A1(new_n23525_), .A2(new_n2253_), .ZN(new_n23526_));
  AOI21_X1   g23333(.A1(new_n23522_), .A2(\asqrt[46] ), .B(new_n23526_), .ZN(new_n23527_));
  NOR2_X1    g23334(.A1(new_n23527_), .A2(new_n23521_), .ZN(new_n23528_));
  AOI22_X1   g23335(.A1(new_n23522_), .A2(\asqrt[46] ), .B1(new_n23520_), .B2(new_n23513_), .ZN(new_n23529_));
  NOR4_X1    g23336(.A1(new_n23158_), .A2(\asqrt[47] ), .A3(new_n22825_), .A4(new_n22830_), .ZN(new_n23530_));
  AOI21_X1   g23337(.A1(new_n23523_), .A2(new_n23083_), .B(new_n2253_), .ZN(new_n23531_));
  NOR2_X1    g23338(.A1(new_n23530_), .A2(new_n23531_), .ZN(new_n23532_));
  NAND2_X1   g23339(.A1(new_n23532_), .A2(new_n2046_), .ZN(new_n23533_));
  INV_X1     g23340(.I(new_n23533_), .ZN(new_n23534_));
  OAI21_X1   g23341(.A1(new_n23529_), .A2(new_n2253_), .B(new_n23534_), .ZN(new_n23535_));
  NAND2_X1   g23342(.A1(new_n23535_), .A2(new_n23528_), .ZN(new_n23536_));
  OAI22_X1   g23343(.A1(new_n23529_), .A2(new_n2253_), .B1(new_n23527_), .B2(new_n23521_), .ZN(new_n23537_));
  NAND2_X1   g23344(.A1(new_n23091_), .A2(\asqrt[48] ), .ZN(new_n23538_));
  NOR4_X1    g23345(.A1(new_n23158_), .A2(\asqrt[48] ), .A3(new_n22833_), .A4(new_n23091_), .ZN(new_n23539_));
  XOR2_X1    g23346(.A1(new_n23539_), .A2(new_n23538_), .Z(new_n23540_));
  NAND2_X1   g23347(.A1(new_n23540_), .A2(new_n1854_), .ZN(new_n23541_));
  AOI21_X1   g23348(.A1(new_n23537_), .A2(\asqrt[48] ), .B(new_n23541_), .ZN(new_n23542_));
  NOR2_X1    g23349(.A1(new_n23542_), .A2(new_n23536_), .ZN(new_n23543_));
  AOI22_X1   g23350(.A1(new_n23537_), .A2(\asqrt[48] ), .B1(new_n23535_), .B2(new_n23528_), .ZN(new_n23544_));
  NOR4_X1    g23351(.A1(new_n23158_), .A2(\asqrt[49] ), .A3(new_n22840_), .A4(new_n22845_), .ZN(new_n23545_));
  AOI21_X1   g23352(.A1(new_n23538_), .A2(new_n23090_), .B(new_n1854_), .ZN(new_n23546_));
  NOR2_X1    g23353(.A1(new_n23545_), .A2(new_n23546_), .ZN(new_n23547_));
  NAND2_X1   g23354(.A1(new_n23547_), .A2(new_n1595_), .ZN(new_n23548_));
  INV_X1     g23355(.I(new_n23548_), .ZN(new_n23549_));
  OAI21_X1   g23356(.A1(new_n23544_), .A2(new_n1854_), .B(new_n23549_), .ZN(new_n23550_));
  NAND2_X1   g23357(.A1(new_n23550_), .A2(new_n23543_), .ZN(new_n23551_));
  OAI22_X1   g23358(.A1(new_n23544_), .A2(new_n1854_), .B1(new_n23542_), .B2(new_n23536_), .ZN(new_n23552_));
  NAND2_X1   g23359(.A1(new_n23098_), .A2(\asqrt[50] ), .ZN(new_n23553_));
  NOR4_X1    g23360(.A1(new_n23158_), .A2(\asqrt[50] ), .A3(new_n22848_), .A4(new_n23098_), .ZN(new_n23554_));
  XOR2_X1    g23361(.A1(new_n23554_), .A2(new_n23553_), .Z(new_n23555_));
  NAND2_X1   g23362(.A1(new_n23555_), .A2(new_n1436_), .ZN(new_n23556_));
  AOI21_X1   g23363(.A1(new_n23552_), .A2(\asqrt[50] ), .B(new_n23556_), .ZN(new_n23557_));
  NOR2_X1    g23364(.A1(new_n23557_), .A2(new_n23551_), .ZN(new_n23558_));
  AOI22_X1   g23365(.A1(new_n23552_), .A2(\asqrt[50] ), .B1(new_n23550_), .B2(new_n23543_), .ZN(new_n23559_));
  NAND2_X1   g23366(.A1(new_n22860_), .A2(\asqrt[51] ), .ZN(new_n23560_));
  NOR4_X1    g23367(.A1(new_n23158_), .A2(\asqrt[51] ), .A3(new_n22855_), .A4(new_n22860_), .ZN(new_n23561_));
  XOR2_X1    g23368(.A1(new_n23561_), .A2(new_n23560_), .Z(new_n23562_));
  NAND2_X1   g23369(.A1(new_n23562_), .A2(new_n1260_), .ZN(new_n23563_));
  INV_X1     g23370(.I(new_n23563_), .ZN(new_n23564_));
  OAI21_X1   g23371(.A1(new_n23559_), .A2(new_n1436_), .B(new_n23564_), .ZN(new_n23565_));
  NAND2_X1   g23372(.A1(new_n23565_), .A2(new_n23558_), .ZN(new_n23566_));
  OAI22_X1   g23373(.A1(new_n23559_), .A2(new_n1436_), .B1(new_n23557_), .B2(new_n23551_), .ZN(new_n23567_));
  NOR4_X1    g23374(.A1(new_n23158_), .A2(\asqrt[52] ), .A3(new_n22863_), .A4(new_n23105_), .ZN(new_n23568_));
  AOI21_X1   g23375(.A1(new_n23560_), .A2(new_n22859_), .B(new_n1260_), .ZN(new_n23569_));
  NOR2_X1    g23376(.A1(new_n23568_), .A2(new_n23569_), .ZN(new_n23570_));
  NAND2_X1   g23377(.A1(new_n23570_), .A2(new_n1096_), .ZN(new_n23571_));
  AOI21_X1   g23378(.A1(new_n23567_), .A2(\asqrt[52] ), .B(new_n23571_), .ZN(new_n23572_));
  NOR2_X1    g23379(.A1(new_n23572_), .A2(new_n23566_), .ZN(new_n23573_));
  AOI22_X1   g23380(.A1(new_n23567_), .A2(\asqrt[52] ), .B1(new_n23565_), .B2(new_n23558_), .ZN(new_n23574_));
  NAND2_X1   g23381(.A1(new_n22875_), .A2(\asqrt[53] ), .ZN(new_n23575_));
  NOR4_X1    g23382(.A1(new_n23158_), .A2(\asqrt[53] ), .A3(new_n22870_), .A4(new_n22875_), .ZN(new_n23576_));
  XOR2_X1    g23383(.A1(new_n23576_), .A2(new_n23575_), .Z(new_n23577_));
  NAND2_X1   g23384(.A1(new_n23577_), .A2(new_n970_), .ZN(new_n23578_));
  INV_X1     g23385(.I(new_n23578_), .ZN(new_n23579_));
  OAI21_X1   g23386(.A1(new_n23574_), .A2(new_n1096_), .B(new_n23579_), .ZN(new_n23580_));
  NAND2_X1   g23387(.A1(new_n23580_), .A2(new_n23573_), .ZN(new_n23581_));
  OAI22_X1   g23388(.A1(new_n23574_), .A2(new_n1096_), .B1(new_n23572_), .B2(new_n23566_), .ZN(new_n23582_));
  NAND2_X1   g23389(.A1(new_n23112_), .A2(\asqrt[54] ), .ZN(new_n23583_));
  NOR4_X1    g23390(.A1(new_n23158_), .A2(\asqrt[54] ), .A3(new_n22878_), .A4(new_n23112_), .ZN(new_n23584_));
  XOR2_X1    g23391(.A1(new_n23584_), .A2(new_n23583_), .Z(new_n23585_));
  NAND2_X1   g23392(.A1(new_n23585_), .A2(new_n825_), .ZN(new_n23586_));
  AOI21_X1   g23393(.A1(new_n23582_), .A2(\asqrt[54] ), .B(new_n23586_), .ZN(new_n23587_));
  NOR2_X1    g23394(.A1(new_n23587_), .A2(new_n23581_), .ZN(new_n23588_));
  AOI22_X1   g23395(.A1(new_n23582_), .A2(\asqrt[54] ), .B1(new_n23580_), .B2(new_n23573_), .ZN(new_n23589_));
  NOR4_X1    g23396(.A1(new_n23158_), .A2(\asqrt[55] ), .A3(new_n22885_), .A4(new_n22890_), .ZN(new_n23590_));
  AOI21_X1   g23397(.A1(new_n23583_), .A2(new_n23111_), .B(new_n825_), .ZN(new_n23591_));
  NOR2_X1    g23398(.A1(new_n23590_), .A2(new_n23591_), .ZN(new_n23592_));
  NAND2_X1   g23399(.A1(new_n23592_), .A2(new_n724_), .ZN(new_n23593_));
  INV_X1     g23400(.I(new_n23593_), .ZN(new_n23594_));
  OAI21_X1   g23401(.A1(new_n23589_), .A2(new_n825_), .B(new_n23594_), .ZN(new_n23595_));
  NAND2_X1   g23402(.A1(new_n23595_), .A2(new_n23588_), .ZN(new_n23596_));
  OAI22_X1   g23403(.A1(new_n23589_), .A2(new_n825_), .B1(new_n23587_), .B2(new_n23581_), .ZN(new_n23597_));
  NAND2_X1   g23404(.A1(new_n23119_), .A2(\asqrt[56] ), .ZN(new_n23598_));
  NOR4_X1    g23405(.A1(new_n23158_), .A2(\asqrt[56] ), .A3(new_n22893_), .A4(new_n23119_), .ZN(new_n23599_));
  XOR2_X1    g23406(.A1(new_n23599_), .A2(new_n23598_), .Z(new_n23600_));
  NAND2_X1   g23407(.A1(new_n23600_), .A2(new_n587_), .ZN(new_n23601_));
  AOI21_X1   g23408(.A1(new_n23597_), .A2(\asqrt[56] ), .B(new_n23601_), .ZN(new_n23602_));
  NOR2_X1    g23409(.A1(new_n23602_), .A2(new_n23596_), .ZN(new_n23603_));
  AOI22_X1   g23410(.A1(new_n23597_), .A2(\asqrt[56] ), .B1(new_n23595_), .B2(new_n23588_), .ZN(new_n23604_));
  NOR4_X1    g23411(.A1(new_n23158_), .A2(\asqrt[57] ), .A3(new_n22900_), .A4(new_n22905_), .ZN(new_n23605_));
  XOR2_X1    g23412(.A1(new_n23605_), .A2(new_n23161_), .Z(new_n23606_));
  NAND2_X1   g23413(.A1(new_n23606_), .A2(new_n504_), .ZN(new_n23607_));
  INV_X1     g23414(.I(new_n23607_), .ZN(new_n23608_));
  OAI21_X1   g23415(.A1(new_n23604_), .A2(new_n587_), .B(new_n23608_), .ZN(new_n23609_));
  NAND2_X1   g23416(.A1(new_n23609_), .A2(new_n23603_), .ZN(new_n23610_));
  OAI22_X1   g23417(.A1(new_n23604_), .A2(new_n587_), .B1(new_n23602_), .B2(new_n23596_), .ZN(new_n23611_));
  NOR4_X1    g23418(.A1(new_n23158_), .A2(\asqrt[58] ), .A3(new_n22908_), .A4(new_n23126_), .ZN(new_n23612_));
  XNOR2_X1   g23419(.A1(new_n23612_), .A2(new_n23162_), .ZN(new_n23613_));
  NAND2_X1   g23420(.A1(new_n23613_), .A2(new_n376_), .ZN(new_n23614_));
  AOI21_X1   g23421(.A1(new_n23611_), .A2(\asqrt[58] ), .B(new_n23614_), .ZN(new_n23615_));
  NOR2_X1    g23422(.A1(new_n23615_), .A2(new_n23610_), .ZN(new_n23616_));
  AOI22_X1   g23423(.A1(new_n23611_), .A2(\asqrt[58] ), .B1(new_n23609_), .B2(new_n23603_), .ZN(new_n23617_));
  NOR4_X1    g23424(.A1(new_n23158_), .A2(\asqrt[59] ), .A3(new_n22915_), .A4(new_n22920_), .ZN(new_n23618_));
  XOR2_X1    g23425(.A1(new_n23618_), .A2(new_n23163_), .Z(new_n23619_));
  NAND2_X1   g23426(.A1(new_n23619_), .A2(new_n275_), .ZN(new_n23620_));
  INV_X1     g23427(.I(new_n23620_), .ZN(new_n23621_));
  OAI21_X1   g23428(.A1(new_n23617_), .A2(new_n376_), .B(new_n23621_), .ZN(new_n23622_));
  NAND2_X1   g23429(.A1(new_n23622_), .A2(new_n23616_), .ZN(new_n23623_));
  OAI22_X1   g23430(.A1(new_n23617_), .A2(new_n376_), .B1(new_n23615_), .B2(new_n23610_), .ZN(new_n23624_));
  NOR4_X1    g23431(.A1(new_n23158_), .A2(\asqrt[60] ), .A3(new_n22923_), .A4(new_n23133_), .ZN(new_n23625_));
  XOR2_X1    g23432(.A1(new_n23625_), .A2(new_n23143_), .Z(new_n23626_));
  NAND2_X1   g23433(.A1(new_n23626_), .A2(new_n229_), .ZN(new_n23627_));
  AOI21_X1   g23434(.A1(new_n23624_), .A2(\asqrt[60] ), .B(new_n23627_), .ZN(new_n23628_));
  NOR2_X1    g23435(.A1(new_n23628_), .A2(new_n23623_), .ZN(new_n23629_));
  AOI22_X1   g23436(.A1(new_n23624_), .A2(\asqrt[60] ), .B1(new_n23622_), .B2(new_n23616_), .ZN(new_n23630_));
  INV_X1     g23437(.I(new_n23167_), .ZN(new_n23631_));
  NOR2_X1    g23438(.A1(new_n23631_), .A2(\asqrt[62] ), .ZN(new_n23632_));
  NOR3_X1    g23439(.A1(new_n23630_), .A2(new_n229_), .A3(new_n23632_), .ZN(new_n23633_));
  AOI21_X1   g23440(.A1(new_n23633_), .A2(new_n23629_), .B(new_n23168_), .ZN(new_n23634_));
  NAND3_X1   g23441(.A1(new_n23158_), .A2(new_n23142_), .A3(new_n23185_), .ZN(new_n23635_));
  AOI21_X1   g23442(.A1(new_n23635_), .A2(new_n23177_), .B(\asqrt[63] ), .ZN(new_n23636_));
  AOI21_X1   g23443(.A1(new_n23634_), .A2(new_n23636_), .B(new_n23160_), .ZN(new_n23637_));
  INV_X1     g23444(.I(new_n23189_), .ZN(new_n23638_));
  INV_X1     g23445(.I(new_n23169_), .ZN(new_n23639_));
  NAND3_X1   g23446(.A1(\asqrt[2] ), .A2(\a[4] ), .A3(\asqrt[3] ), .ZN(new_n23640_));
  INV_X1     g23447(.I(\a[4] ), .ZN(new_n23641_));
  NAND4_X1   g23448(.A1(new_n23179_), .A2(new_n23641_), .A3(\asqrt[3] ), .A4(new_n23178_), .ZN(new_n23642_));
  AOI21_X1   g23449(.A1(new_n23640_), .A2(new_n23642_), .B(new_n23639_), .ZN(new_n23643_));
  NOR3_X1    g23450(.A1(new_n23199_), .A2(new_n21585_), .A3(\asqrt[2] ), .ZN(new_n23644_));
  AOI21_X1   g23451(.A1(new_n23195_), .A2(new_n21584_), .B(new_n23158_), .ZN(new_n23645_));
  NOR4_X1    g23452(.A1(new_n23643_), .A2(\asqrt[4] ), .A3(new_n23644_), .A4(new_n23645_), .ZN(new_n23646_));
  NOR2_X1    g23453(.A1(new_n23646_), .A2(new_n23638_), .ZN(new_n23647_));
  INV_X1     g23454(.I(new_n23181_), .ZN(new_n23648_));
  AOI21_X1   g23455(.A1(new_n23187_), .A2(new_n23648_), .B(new_n23183_), .ZN(new_n23649_));
  NOR3_X1    g23456(.A1(new_n23180_), .A2(new_n23641_), .A3(new_n23171_), .ZN(new_n23650_));
  NOR3_X1    g23457(.A1(new_n23643_), .A2(new_n23649_), .A3(new_n23650_), .ZN(new_n23651_));
  INV_X1     g23458(.I(new_n23211_), .ZN(new_n23652_));
  NOR3_X1    g23459(.A1(new_n23652_), .A2(\asqrt[5] ), .A3(new_n23208_), .ZN(new_n23653_));
  OAI21_X1   g23460(.A1(new_n23651_), .A2(new_n21781_), .B(new_n23653_), .ZN(new_n23654_));
  NAND2_X1   g23461(.A1(new_n23647_), .A2(new_n23654_), .ZN(new_n23655_));
  OAI22_X1   g23462(.A1(new_n23646_), .A2(new_n23638_), .B1(new_n23651_), .B2(new_n21781_), .ZN(new_n23656_));
  AOI21_X1   g23463(.A1(new_n23656_), .A2(\asqrt[5] ), .B(new_n23220_), .ZN(new_n23657_));
  NOR2_X1    g23464(.A1(new_n23657_), .A2(new_n23655_), .ZN(new_n23658_));
  AOI22_X1   g23465(.A1(new_n23656_), .A2(\asqrt[5] ), .B1(new_n23647_), .B2(new_n23654_), .ZN(new_n23659_));
  INV_X1     g23466(.I(new_n23228_), .ZN(new_n23660_));
  OAI21_X1   g23467(.A1(new_n23659_), .A2(new_n20455_), .B(new_n23660_), .ZN(new_n23661_));
  NAND2_X1   g23468(.A1(new_n23661_), .A2(new_n23658_), .ZN(new_n23662_));
  OAI22_X1   g23469(.A1(new_n23659_), .A2(new_n20455_), .B1(new_n23657_), .B2(new_n23655_), .ZN(new_n23663_));
  AOI21_X1   g23470(.A1(new_n23663_), .A2(\asqrt[7] ), .B(new_n23234_), .ZN(new_n23664_));
  NOR2_X1    g23471(.A1(new_n23664_), .A2(new_n23662_), .ZN(new_n23665_));
  AOI22_X1   g23472(.A1(new_n23663_), .A2(\asqrt[7] ), .B1(new_n23661_), .B2(new_n23658_), .ZN(new_n23666_));
  INV_X1     g23473(.I(new_n23241_), .ZN(new_n23667_));
  OAI21_X1   g23474(.A1(new_n23666_), .A2(new_n19100_), .B(new_n23667_), .ZN(new_n23668_));
  NAND2_X1   g23475(.A1(new_n23668_), .A2(new_n23665_), .ZN(new_n23669_));
  OAI22_X1   g23476(.A1(new_n23666_), .A2(new_n19100_), .B1(new_n23664_), .B2(new_n23662_), .ZN(new_n23670_));
  AOI21_X1   g23477(.A1(new_n23670_), .A2(\asqrt[9] ), .B(new_n23248_), .ZN(new_n23671_));
  NOR2_X1    g23478(.A1(new_n23671_), .A2(new_n23669_), .ZN(new_n23672_));
  AOI22_X1   g23479(.A1(new_n23670_), .A2(\asqrt[9] ), .B1(new_n23668_), .B2(new_n23665_), .ZN(new_n23673_));
  INV_X1     g23480(.I(new_n23256_), .ZN(new_n23674_));
  OAI21_X1   g23481(.A1(new_n23673_), .A2(new_n17893_), .B(new_n23674_), .ZN(new_n23675_));
  NAND2_X1   g23482(.A1(new_n23675_), .A2(new_n23672_), .ZN(new_n23676_));
  OAI22_X1   g23483(.A1(new_n23673_), .A2(new_n17893_), .B1(new_n23671_), .B2(new_n23669_), .ZN(new_n23677_));
  AOI21_X1   g23484(.A1(new_n23677_), .A2(\asqrt[11] ), .B(new_n23263_), .ZN(new_n23678_));
  NOR2_X1    g23485(.A1(new_n23678_), .A2(new_n23676_), .ZN(new_n23679_));
  AOI22_X1   g23486(.A1(new_n23677_), .A2(\asqrt[11] ), .B1(new_n23675_), .B2(new_n23672_), .ZN(new_n23680_));
  INV_X1     g23487(.I(new_n23271_), .ZN(new_n23681_));
  OAI21_X1   g23488(.A1(new_n23680_), .A2(new_n16619_), .B(new_n23681_), .ZN(new_n23682_));
  NAND2_X1   g23489(.A1(new_n23682_), .A2(new_n23679_), .ZN(new_n23683_));
  OAI22_X1   g23490(.A1(new_n23680_), .A2(new_n16619_), .B1(new_n23678_), .B2(new_n23676_), .ZN(new_n23684_));
  AOI21_X1   g23491(.A1(new_n23684_), .A2(\asqrt[13] ), .B(new_n23278_), .ZN(new_n23685_));
  NOR2_X1    g23492(.A1(new_n23685_), .A2(new_n23683_), .ZN(new_n23686_));
  AOI22_X1   g23493(.A1(new_n23684_), .A2(\asqrt[13] ), .B1(new_n23682_), .B2(new_n23679_), .ZN(new_n23687_));
  INV_X1     g23494(.I(new_n23286_), .ZN(new_n23688_));
  OAI21_X1   g23495(.A1(new_n23687_), .A2(new_n15447_), .B(new_n23688_), .ZN(new_n23689_));
  NAND2_X1   g23496(.A1(new_n23689_), .A2(new_n23686_), .ZN(new_n23690_));
  OAI22_X1   g23497(.A1(new_n23687_), .A2(new_n15447_), .B1(new_n23685_), .B2(new_n23683_), .ZN(new_n23691_));
  AOI21_X1   g23498(.A1(new_n23691_), .A2(\asqrt[15] ), .B(new_n23293_), .ZN(new_n23692_));
  NOR2_X1    g23499(.A1(new_n23692_), .A2(new_n23690_), .ZN(new_n23693_));
  AOI22_X1   g23500(.A1(new_n23691_), .A2(\asqrt[15] ), .B1(new_n23689_), .B2(new_n23686_), .ZN(new_n23694_));
  INV_X1     g23501(.I(new_n23301_), .ZN(new_n23695_));
  OAI21_X1   g23502(.A1(new_n23694_), .A2(new_n14273_), .B(new_n23695_), .ZN(new_n23696_));
  NAND2_X1   g23503(.A1(new_n23696_), .A2(new_n23693_), .ZN(new_n23697_));
  OAI22_X1   g23504(.A1(new_n23694_), .A2(new_n14273_), .B1(new_n23692_), .B2(new_n23690_), .ZN(new_n23698_));
  AOI21_X1   g23505(.A1(new_n23698_), .A2(\asqrt[17] ), .B(new_n23308_), .ZN(new_n23699_));
  NOR2_X1    g23506(.A1(new_n23699_), .A2(new_n23697_), .ZN(new_n23700_));
  AOI22_X1   g23507(.A1(new_n23698_), .A2(\asqrt[17] ), .B1(new_n23696_), .B2(new_n23693_), .ZN(new_n23701_));
  INV_X1     g23508(.I(new_n23316_), .ZN(new_n23702_));
  OAI21_X1   g23509(.A1(new_n23701_), .A2(new_n13192_), .B(new_n23702_), .ZN(new_n23703_));
  NAND2_X1   g23510(.A1(new_n23703_), .A2(new_n23700_), .ZN(new_n23704_));
  OAI22_X1   g23511(.A1(new_n23701_), .A2(new_n13192_), .B1(new_n23699_), .B2(new_n23697_), .ZN(new_n23705_));
  AOI21_X1   g23512(.A1(new_n23705_), .A2(\asqrt[19] ), .B(new_n23323_), .ZN(new_n23706_));
  NOR2_X1    g23513(.A1(new_n23706_), .A2(new_n23704_), .ZN(new_n23707_));
  AOI22_X1   g23514(.A1(new_n23705_), .A2(\asqrt[19] ), .B1(new_n23703_), .B2(new_n23700_), .ZN(new_n23708_));
  INV_X1     g23515(.I(new_n23331_), .ZN(new_n23709_));
  OAI21_X1   g23516(.A1(new_n23708_), .A2(new_n12101_), .B(new_n23709_), .ZN(new_n23710_));
  NAND2_X1   g23517(.A1(new_n23710_), .A2(new_n23707_), .ZN(new_n23711_));
  OAI22_X1   g23518(.A1(new_n23708_), .A2(new_n12101_), .B1(new_n23706_), .B2(new_n23704_), .ZN(new_n23712_));
  AOI21_X1   g23519(.A1(new_n23712_), .A2(\asqrt[21] ), .B(new_n23338_), .ZN(new_n23713_));
  NOR2_X1    g23520(.A1(new_n23713_), .A2(new_n23711_), .ZN(new_n23714_));
  AOI22_X1   g23521(.A1(new_n23712_), .A2(\asqrt[21] ), .B1(new_n23710_), .B2(new_n23707_), .ZN(new_n23715_));
  INV_X1     g23522(.I(new_n23346_), .ZN(new_n23716_));
  OAI21_X1   g23523(.A1(new_n23715_), .A2(new_n11105_), .B(new_n23716_), .ZN(new_n23717_));
  NAND2_X1   g23524(.A1(new_n23717_), .A2(new_n23714_), .ZN(new_n23718_));
  OAI22_X1   g23525(.A1(new_n23715_), .A2(new_n11105_), .B1(new_n23713_), .B2(new_n23711_), .ZN(new_n23719_));
  AOI21_X1   g23526(.A1(new_n23719_), .A2(\asqrt[23] ), .B(new_n23353_), .ZN(new_n23720_));
  NOR2_X1    g23527(.A1(new_n23720_), .A2(new_n23718_), .ZN(new_n23721_));
  AOI22_X1   g23528(.A1(new_n23719_), .A2(\asqrt[23] ), .B1(new_n23717_), .B2(new_n23714_), .ZN(new_n23722_));
  INV_X1     g23529(.I(new_n23361_), .ZN(new_n23723_));
  OAI21_X1   g23530(.A1(new_n23722_), .A2(new_n10104_), .B(new_n23723_), .ZN(new_n23724_));
  NAND2_X1   g23531(.A1(new_n23724_), .A2(new_n23721_), .ZN(new_n23725_));
  OAI22_X1   g23532(.A1(new_n23722_), .A2(new_n10104_), .B1(new_n23720_), .B2(new_n23718_), .ZN(new_n23726_));
  AOI21_X1   g23533(.A1(new_n23726_), .A2(\asqrt[25] ), .B(new_n23368_), .ZN(new_n23727_));
  NOR2_X1    g23534(.A1(new_n23727_), .A2(new_n23725_), .ZN(new_n23728_));
  AOI22_X1   g23535(.A1(new_n23726_), .A2(\asqrt[25] ), .B1(new_n23724_), .B2(new_n23721_), .ZN(new_n23729_));
  INV_X1     g23536(.I(new_n23376_), .ZN(new_n23730_));
  OAI21_X1   g23537(.A1(new_n23729_), .A2(new_n9212_), .B(new_n23730_), .ZN(new_n23731_));
  NAND2_X1   g23538(.A1(new_n23731_), .A2(new_n23728_), .ZN(new_n23732_));
  OAI22_X1   g23539(.A1(new_n23729_), .A2(new_n9212_), .B1(new_n23727_), .B2(new_n23725_), .ZN(new_n23733_));
  AOI21_X1   g23540(.A1(new_n23733_), .A2(\asqrt[27] ), .B(new_n23383_), .ZN(new_n23734_));
  NOR2_X1    g23541(.A1(new_n23734_), .A2(new_n23732_), .ZN(new_n23735_));
  AOI22_X1   g23542(.A1(new_n23733_), .A2(\asqrt[27] ), .B1(new_n23731_), .B2(new_n23728_), .ZN(new_n23736_));
  INV_X1     g23543(.I(new_n23391_), .ZN(new_n23737_));
  OAI21_X1   g23544(.A1(new_n23736_), .A2(new_n8319_), .B(new_n23737_), .ZN(new_n23738_));
  NAND2_X1   g23545(.A1(new_n23738_), .A2(new_n23735_), .ZN(new_n23739_));
  OAI22_X1   g23546(.A1(new_n23736_), .A2(new_n8319_), .B1(new_n23734_), .B2(new_n23732_), .ZN(new_n23740_));
  AOI21_X1   g23547(.A1(new_n23740_), .A2(\asqrt[29] ), .B(new_n23398_), .ZN(new_n23741_));
  NOR2_X1    g23548(.A1(new_n23741_), .A2(new_n23739_), .ZN(new_n23742_));
  AOI22_X1   g23549(.A1(new_n23740_), .A2(\asqrt[29] ), .B1(new_n23738_), .B2(new_n23735_), .ZN(new_n23743_));
  INV_X1     g23550(.I(new_n23406_), .ZN(new_n23744_));
  OAI21_X1   g23551(.A1(new_n23743_), .A2(new_n7517_), .B(new_n23744_), .ZN(new_n23745_));
  NAND2_X1   g23552(.A1(new_n23745_), .A2(new_n23742_), .ZN(new_n23746_));
  OAI22_X1   g23553(.A1(new_n23743_), .A2(new_n7517_), .B1(new_n23741_), .B2(new_n23739_), .ZN(new_n23747_));
  AOI21_X1   g23554(.A1(new_n23747_), .A2(\asqrt[31] ), .B(new_n23413_), .ZN(new_n23748_));
  NOR2_X1    g23555(.A1(new_n23748_), .A2(new_n23746_), .ZN(new_n23749_));
  AOI22_X1   g23556(.A1(new_n23747_), .A2(\asqrt[31] ), .B1(new_n23745_), .B2(new_n23742_), .ZN(new_n23750_));
  INV_X1     g23557(.I(new_n23421_), .ZN(new_n23751_));
  OAI21_X1   g23558(.A1(new_n23750_), .A2(new_n6708_), .B(new_n23751_), .ZN(new_n23752_));
  NAND2_X1   g23559(.A1(new_n23752_), .A2(new_n23749_), .ZN(new_n23753_));
  OAI22_X1   g23560(.A1(new_n23750_), .A2(new_n6708_), .B1(new_n23748_), .B2(new_n23746_), .ZN(new_n23754_));
  AOI21_X1   g23561(.A1(new_n23754_), .A2(\asqrt[33] ), .B(new_n23428_), .ZN(new_n23755_));
  NOR2_X1    g23562(.A1(new_n23755_), .A2(new_n23753_), .ZN(new_n23756_));
  AOI22_X1   g23563(.A1(new_n23754_), .A2(\asqrt[33] ), .B1(new_n23752_), .B2(new_n23749_), .ZN(new_n23757_));
  INV_X1     g23564(.I(new_n23436_), .ZN(new_n23758_));
  OAI21_X1   g23565(.A1(new_n23757_), .A2(new_n5991_), .B(new_n23758_), .ZN(new_n23759_));
  NAND2_X1   g23566(.A1(new_n23759_), .A2(new_n23756_), .ZN(new_n23760_));
  OAI22_X1   g23567(.A1(new_n23757_), .A2(new_n5991_), .B1(new_n23755_), .B2(new_n23753_), .ZN(new_n23761_));
  AOI21_X1   g23568(.A1(new_n23761_), .A2(\asqrt[35] ), .B(new_n23443_), .ZN(new_n23762_));
  NOR2_X1    g23569(.A1(new_n23762_), .A2(new_n23760_), .ZN(new_n23763_));
  AOI22_X1   g23570(.A1(new_n23761_), .A2(\asqrt[35] ), .B1(new_n23759_), .B2(new_n23756_), .ZN(new_n23764_));
  INV_X1     g23571(.I(new_n23451_), .ZN(new_n23765_));
  OAI21_X1   g23572(.A1(new_n23764_), .A2(new_n5273_), .B(new_n23765_), .ZN(new_n23766_));
  NAND2_X1   g23573(.A1(new_n23766_), .A2(new_n23763_), .ZN(new_n23767_));
  OAI22_X1   g23574(.A1(new_n23764_), .A2(new_n5273_), .B1(new_n23762_), .B2(new_n23760_), .ZN(new_n23768_));
  AOI21_X1   g23575(.A1(new_n23768_), .A2(\asqrt[37] ), .B(new_n23458_), .ZN(new_n23769_));
  NOR2_X1    g23576(.A1(new_n23769_), .A2(new_n23767_), .ZN(new_n23770_));
  AOI22_X1   g23577(.A1(new_n23768_), .A2(\asqrt[37] ), .B1(new_n23766_), .B2(new_n23763_), .ZN(new_n23771_));
  INV_X1     g23578(.I(new_n23466_), .ZN(new_n23772_));
  OAI21_X1   g23579(.A1(new_n23771_), .A2(new_n4645_), .B(new_n23772_), .ZN(new_n23773_));
  NAND2_X1   g23580(.A1(new_n23773_), .A2(new_n23770_), .ZN(new_n23774_));
  OAI22_X1   g23581(.A1(new_n23771_), .A2(new_n4645_), .B1(new_n23769_), .B2(new_n23767_), .ZN(new_n23775_));
  AOI21_X1   g23582(.A1(new_n23775_), .A2(\asqrt[39] ), .B(new_n23473_), .ZN(new_n23776_));
  NOR2_X1    g23583(.A1(new_n23776_), .A2(new_n23774_), .ZN(new_n23777_));
  AOI22_X1   g23584(.A1(new_n23775_), .A2(\asqrt[39] ), .B1(new_n23773_), .B2(new_n23770_), .ZN(new_n23778_));
  INV_X1     g23585(.I(new_n23481_), .ZN(new_n23779_));
  OAI21_X1   g23586(.A1(new_n23778_), .A2(new_n4018_), .B(new_n23779_), .ZN(new_n23780_));
  NAND2_X1   g23587(.A1(new_n23780_), .A2(new_n23777_), .ZN(new_n23781_));
  OAI22_X1   g23588(.A1(new_n23778_), .A2(new_n4018_), .B1(new_n23776_), .B2(new_n23774_), .ZN(new_n23782_));
  AOI21_X1   g23589(.A1(new_n23782_), .A2(\asqrt[41] ), .B(new_n23488_), .ZN(new_n23783_));
  NOR2_X1    g23590(.A1(new_n23783_), .A2(new_n23781_), .ZN(new_n23784_));
  AOI22_X1   g23591(.A1(new_n23782_), .A2(\asqrt[41] ), .B1(new_n23780_), .B2(new_n23777_), .ZN(new_n23785_));
  INV_X1     g23592(.I(new_n23496_), .ZN(new_n23786_));
  OAI21_X1   g23593(.A1(new_n23785_), .A2(new_n3481_), .B(new_n23786_), .ZN(new_n23787_));
  NAND2_X1   g23594(.A1(new_n23787_), .A2(new_n23784_), .ZN(new_n23788_));
  OAI22_X1   g23595(.A1(new_n23785_), .A2(new_n3481_), .B1(new_n23783_), .B2(new_n23781_), .ZN(new_n23789_));
  AOI21_X1   g23596(.A1(new_n23789_), .A2(\asqrt[43] ), .B(new_n23503_), .ZN(new_n23790_));
  NOR2_X1    g23597(.A1(new_n23790_), .A2(new_n23788_), .ZN(new_n23791_));
  AOI22_X1   g23598(.A1(new_n23789_), .A2(\asqrt[43] ), .B1(new_n23787_), .B2(new_n23784_), .ZN(new_n23792_));
  INV_X1     g23599(.I(new_n23511_), .ZN(new_n23793_));
  OAI21_X1   g23600(.A1(new_n23792_), .A2(new_n2941_), .B(new_n23793_), .ZN(new_n23794_));
  NAND2_X1   g23601(.A1(new_n23794_), .A2(new_n23791_), .ZN(new_n23795_));
  OAI22_X1   g23602(.A1(new_n23792_), .A2(new_n2941_), .B1(new_n23790_), .B2(new_n23788_), .ZN(new_n23796_));
  AOI21_X1   g23603(.A1(new_n23796_), .A2(\asqrt[45] ), .B(new_n23518_), .ZN(new_n23797_));
  NOR2_X1    g23604(.A1(new_n23797_), .A2(new_n23795_), .ZN(new_n23798_));
  AOI22_X1   g23605(.A1(new_n23796_), .A2(\asqrt[45] ), .B1(new_n23794_), .B2(new_n23791_), .ZN(new_n23799_));
  INV_X1     g23606(.I(new_n23526_), .ZN(new_n23800_));
  OAI21_X1   g23607(.A1(new_n23799_), .A2(new_n2488_), .B(new_n23800_), .ZN(new_n23801_));
  NAND2_X1   g23608(.A1(new_n23801_), .A2(new_n23798_), .ZN(new_n23802_));
  OAI22_X1   g23609(.A1(new_n23799_), .A2(new_n2488_), .B1(new_n23797_), .B2(new_n23795_), .ZN(new_n23803_));
  AOI21_X1   g23610(.A1(new_n23803_), .A2(\asqrt[47] ), .B(new_n23533_), .ZN(new_n23804_));
  NOR2_X1    g23611(.A1(new_n23804_), .A2(new_n23802_), .ZN(new_n23805_));
  AOI22_X1   g23612(.A1(new_n23803_), .A2(\asqrt[47] ), .B1(new_n23801_), .B2(new_n23798_), .ZN(new_n23806_));
  INV_X1     g23613(.I(new_n23541_), .ZN(new_n23807_));
  OAI21_X1   g23614(.A1(new_n23806_), .A2(new_n2046_), .B(new_n23807_), .ZN(new_n23808_));
  NAND2_X1   g23615(.A1(new_n23808_), .A2(new_n23805_), .ZN(new_n23809_));
  OAI22_X1   g23616(.A1(new_n23806_), .A2(new_n2046_), .B1(new_n23804_), .B2(new_n23802_), .ZN(new_n23810_));
  AOI21_X1   g23617(.A1(new_n23810_), .A2(\asqrt[49] ), .B(new_n23548_), .ZN(new_n23811_));
  NOR2_X1    g23618(.A1(new_n23811_), .A2(new_n23809_), .ZN(new_n23812_));
  AOI22_X1   g23619(.A1(new_n23810_), .A2(\asqrt[49] ), .B1(new_n23808_), .B2(new_n23805_), .ZN(new_n23813_));
  INV_X1     g23620(.I(new_n23556_), .ZN(new_n23814_));
  OAI21_X1   g23621(.A1(new_n23813_), .A2(new_n1595_), .B(new_n23814_), .ZN(new_n23815_));
  NAND2_X1   g23622(.A1(new_n23815_), .A2(new_n23812_), .ZN(new_n23816_));
  OAI22_X1   g23623(.A1(new_n23813_), .A2(new_n1595_), .B1(new_n23811_), .B2(new_n23809_), .ZN(new_n23817_));
  AOI21_X1   g23624(.A1(new_n23817_), .A2(\asqrt[51] ), .B(new_n23563_), .ZN(new_n23818_));
  NOR2_X1    g23625(.A1(new_n23818_), .A2(new_n23816_), .ZN(new_n23819_));
  AOI22_X1   g23626(.A1(new_n23817_), .A2(\asqrt[51] ), .B1(new_n23815_), .B2(new_n23812_), .ZN(new_n23820_));
  INV_X1     g23627(.I(new_n23571_), .ZN(new_n23821_));
  OAI21_X1   g23628(.A1(new_n23820_), .A2(new_n1260_), .B(new_n23821_), .ZN(new_n23822_));
  NAND2_X1   g23629(.A1(new_n23822_), .A2(new_n23819_), .ZN(new_n23823_));
  OAI22_X1   g23630(.A1(new_n23820_), .A2(new_n1260_), .B1(new_n23818_), .B2(new_n23816_), .ZN(new_n23824_));
  AOI21_X1   g23631(.A1(new_n23824_), .A2(\asqrt[53] ), .B(new_n23578_), .ZN(new_n23825_));
  NOR2_X1    g23632(.A1(new_n23825_), .A2(new_n23823_), .ZN(new_n23826_));
  AOI22_X1   g23633(.A1(new_n23824_), .A2(\asqrt[53] ), .B1(new_n23822_), .B2(new_n23819_), .ZN(new_n23827_));
  INV_X1     g23634(.I(new_n23586_), .ZN(new_n23828_));
  OAI21_X1   g23635(.A1(new_n23827_), .A2(new_n970_), .B(new_n23828_), .ZN(new_n23829_));
  NAND2_X1   g23636(.A1(new_n23829_), .A2(new_n23826_), .ZN(new_n23830_));
  OAI22_X1   g23637(.A1(new_n23827_), .A2(new_n970_), .B1(new_n23825_), .B2(new_n23823_), .ZN(new_n23831_));
  AOI21_X1   g23638(.A1(new_n23831_), .A2(\asqrt[55] ), .B(new_n23593_), .ZN(new_n23832_));
  NOR2_X1    g23639(.A1(new_n23832_), .A2(new_n23830_), .ZN(new_n23833_));
  AOI22_X1   g23640(.A1(new_n23831_), .A2(\asqrt[55] ), .B1(new_n23829_), .B2(new_n23826_), .ZN(new_n23834_));
  INV_X1     g23641(.I(new_n23601_), .ZN(new_n23835_));
  OAI21_X1   g23642(.A1(new_n23834_), .A2(new_n724_), .B(new_n23835_), .ZN(new_n23836_));
  NAND2_X1   g23643(.A1(new_n23836_), .A2(new_n23833_), .ZN(new_n23837_));
  OAI22_X1   g23644(.A1(new_n23834_), .A2(new_n724_), .B1(new_n23832_), .B2(new_n23830_), .ZN(new_n23838_));
  AOI21_X1   g23645(.A1(new_n23838_), .A2(\asqrt[57] ), .B(new_n23607_), .ZN(new_n23839_));
  NOR2_X1    g23646(.A1(new_n23839_), .A2(new_n23837_), .ZN(new_n23840_));
  AOI22_X1   g23647(.A1(new_n23838_), .A2(\asqrt[57] ), .B1(new_n23836_), .B2(new_n23833_), .ZN(new_n23841_));
  INV_X1     g23648(.I(new_n23614_), .ZN(new_n23842_));
  OAI21_X1   g23649(.A1(new_n23841_), .A2(new_n504_), .B(new_n23842_), .ZN(new_n23843_));
  NAND2_X1   g23650(.A1(new_n23843_), .A2(new_n23840_), .ZN(new_n23844_));
  OAI22_X1   g23651(.A1(new_n23841_), .A2(new_n504_), .B1(new_n23839_), .B2(new_n23837_), .ZN(new_n23845_));
  AOI21_X1   g23652(.A1(new_n23845_), .A2(\asqrt[59] ), .B(new_n23620_), .ZN(new_n23846_));
  NOR2_X1    g23653(.A1(new_n23846_), .A2(new_n23844_), .ZN(new_n23847_));
  AOI22_X1   g23654(.A1(new_n23845_), .A2(\asqrt[59] ), .B1(new_n23843_), .B2(new_n23840_), .ZN(new_n23848_));
  INV_X1     g23655(.I(new_n23627_), .ZN(new_n23849_));
  OAI21_X1   g23656(.A1(new_n23848_), .A2(new_n275_), .B(new_n23849_), .ZN(new_n23850_));
  NAND2_X1   g23657(.A1(new_n23850_), .A2(new_n23847_), .ZN(new_n23851_));
  NAND2_X1   g23658(.A1(new_n23845_), .A2(\asqrt[59] ), .ZN(new_n23852_));
  AOI21_X1   g23659(.A1(new_n23852_), .A2(new_n23844_), .B(new_n275_), .ZN(new_n23853_));
  OAI21_X1   g23660(.A1(new_n23847_), .A2(new_n23853_), .B(\asqrt[61] ), .ZN(new_n23854_));
  AOI21_X1   g23661(.A1(new_n23854_), .A2(new_n23632_), .B(new_n23851_), .ZN(new_n23855_));
  AOI21_X1   g23662(.A1(new_n23142_), .A2(new_n23149_), .B(new_n23158_), .ZN(new_n23856_));
  XOR2_X1    g23663(.A1(new_n23149_), .A2(\asqrt[63] ), .Z(new_n23857_));
  NOR2_X1    g23664(.A1(new_n23856_), .A2(new_n23857_), .ZN(new_n23858_));
  OAI22_X1   g23665(.A1(new_n23848_), .A2(new_n275_), .B1(new_n23846_), .B2(new_n23844_), .ZN(new_n23859_));
  AOI22_X1   g23666(.A1(new_n23859_), .A2(\asqrt[61] ), .B1(new_n23850_), .B2(new_n23847_), .ZN(new_n23860_));
  OAI21_X1   g23667(.A1(new_n23860_), .A2(new_n196_), .B(new_n23160_), .ZN(new_n23861_));
  OAI21_X1   g23668(.A1(new_n23861_), .A2(new_n23858_), .B(new_n23855_), .ZN(new_n23862_));
  NOR2_X1    g23669(.A1(new_n23862_), .A2(new_n23637_), .ZN(new_n23863_));
  INV_X1     g23670(.I(new_n23160_), .ZN(new_n23864_));
  INV_X1     g23671(.I(new_n23168_), .ZN(new_n23865_));
  INV_X1     g23672(.I(new_n23632_), .ZN(new_n23866_));
  NAND3_X1   g23673(.A1(new_n23859_), .A2(\asqrt[61] ), .A3(new_n23866_), .ZN(new_n23867_));
  OAI21_X1   g23674(.A1(new_n23867_), .A2(new_n23851_), .B(new_n23865_), .ZN(new_n23868_));
  NOR2_X1    g23675(.A1(new_n23868_), .A2(new_n23864_), .ZN(new_n23869_));
  XOR2_X1    g23676(.A1(new_n23868_), .A2(\asqrt[63] ), .Z(new_n23870_));
  OAI21_X1   g23677(.A1(new_n23863_), .A2(new_n23869_), .B(new_n23870_), .ZN(new_n23871_));
  NAND2_X1   g23678(.A1(new_n23611_), .A2(\asqrt[58] ), .ZN(new_n23872_));
  AOI21_X1   g23679(.A1(new_n23872_), .A2(new_n23610_), .B(new_n376_), .ZN(new_n23873_));
  OAI21_X1   g23680(.A1(new_n23616_), .A2(new_n23873_), .B(\asqrt[60] ), .ZN(new_n23874_));
  AOI21_X1   g23681(.A1(new_n23623_), .A2(new_n23874_), .B(new_n229_), .ZN(new_n23875_));
  NOR4_X1    g23682(.A1(new_n23863_), .A2(\asqrt[61] ), .A3(new_n23626_), .A4(new_n23859_), .ZN(new_n23876_));
  XOR2_X1    g23683(.A1(new_n23876_), .A2(new_n23875_), .Z(new_n23877_));
  NOR4_X1    g23684(.A1(new_n23863_), .A2(\asqrt[59] ), .A3(new_n23613_), .A4(new_n23845_), .ZN(new_n23878_));
  XOR2_X1    g23685(.A1(new_n23878_), .A2(new_n23852_), .Z(new_n23879_));
  INV_X1     g23686(.I(new_n23879_), .ZN(new_n23880_));
  NOR2_X1    g23687(.A1(new_n23604_), .A2(new_n587_), .ZN(new_n23881_));
  NOR4_X1    g23688(.A1(new_n23863_), .A2(\asqrt[57] ), .A3(new_n23600_), .A4(new_n23838_), .ZN(new_n23882_));
  XNOR2_X1   g23689(.A1(new_n23882_), .A2(new_n23881_), .ZN(new_n23883_));
  NOR2_X1    g23690(.A1(new_n23589_), .A2(new_n825_), .ZN(new_n23884_));
  NOR4_X1    g23691(.A1(new_n23863_), .A2(\asqrt[55] ), .A3(new_n23585_), .A4(new_n23831_), .ZN(new_n23885_));
  XNOR2_X1   g23692(.A1(new_n23885_), .A2(new_n23884_), .ZN(new_n23886_));
  INV_X1     g23693(.I(new_n23886_), .ZN(new_n23887_));
  NAND2_X1   g23694(.A1(new_n23824_), .A2(\asqrt[53] ), .ZN(new_n23888_));
  NOR4_X1    g23695(.A1(new_n23863_), .A2(\asqrt[53] ), .A3(new_n23570_), .A4(new_n23824_), .ZN(new_n23889_));
  XOR2_X1    g23696(.A1(new_n23889_), .A2(new_n23888_), .Z(new_n23890_));
  NAND2_X1   g23697(.A1(new_n23817_), .A2(\asqrt[51] ), .ZN(new_n23891_));
  NOR4_X1    g23698(.A1(new_n23863_), .A2(\asqrt[51] ), .A3(new_n23555_), .A4(new_n23817_), .ZN(new_n23892_));
  XOR2_X1    g23699(.A1(new_n23892_), .A2(new_n23891_), .Z(new_n23893_));
  INV_X1     g23700(.I(new_n23893_), .ZN(new_n23894_));
  NOR2_X1    g23701(.A1(new_n23544_), .A2(new_n1854_), .ZN(new_n23895_));
  NOR4_X1    g23702(.A1(new_n23863_), .A2(\asqrt[49] ), .A3(new_n23540_), .A4(new_n23810_), .ZN(new_n23896_));
  XNOR2_X1   g23703(.A1(new_n23896_), .A2(new_n23895_), .ZN(new_n23897_));
  NOR2_X1    g23704(.A1(new_n23529_), .A2(new_n2253_), .ZN(new_n23898_));
  NOR4_X1    g23705(.A1(new_n23863_), .A2(\asqrt[47] ), .A3(new_n23525_), .A4(new_n23803_), .ZN(new_n23899_));
  XNOR2_X1   g23706(.A1(new_n23899_), .A2(new_n23898_), .ZN(new_n23900_));
  INV_X1     g23707(.I(new_n23900_), .ZN(new_n23901_));
  NOR2_X1    g23708(.A1(new_n23514_), .A2(new_n2728_), .ZN(new_n23902_));
  NOR4_X1    g23709(.A1(new_n23863_), .A2(\asqrt[45] ), .A3(new_n23510_), .A4(new_n23796_), .ZN(new_n23903_));
  XNOR2_X1   g23710(.A1(new_n23903_), .A2(new_n23902_), .ZN(new_n23904_));
  NAND2_X1   g23711(.A1(new_n23789_), .A2(\asqrt[43] ), .ZN(new_n23905_));
  NOR4_X1    g23712(.A1(new_n23863_), .A2(\asqrt[43] ), .A3(new_n23495_), .A4(new_n23789_), .ZN(new_n23906_));
  XOR2_X1    g23713(.A1(new_n23906_), .A2(new_n23905_), .Z(new_n23907_));
  INV_X1     g23714(.I(new_n23907_), .ZN(new_n23908_));
  NAND2_X1   g23715(.A1(new_n23782_), .A2(\asqrt[41] ), .ZN(new_n23909_));
  NOR4_X1    g23716(.A1(new_n23863_), .A2(\asqrt[41] ), .A3(new_n23480_), .A4(new_n23782_), .ZN(new_n23910_));
  XOR2_X1    g23717(.A1(new_n23910_), .A2(new_n23909_), .Z(new_n23911_));
  NAND2_X1   g23718(.A1(new_n23775_), .A2(\asqrt[39] ), .ZN(new_n23912_));
  NOR4_X1    g23719(.A1(new_n23863_), .A2(\asqrt[39] ), .A3(new_n23465_), .A4(new_n23775_), .ZN(new_n23913_));
  XOR2_X1    g23720(.A1(new_n23913_), .A2(new_n23912_), .Z(new_n23914_));
  INV_X1     g23721(.I(new_n23914_), .ZN(new_n23915_));
  NOR2_X1    g23722(.A1(new_n23454_), .A2(new_n4973_), .ZN(new_n23916_));
  NOR4_X1    g23723(.A1(new_n23863_), .A2(\asqrt[37] ), .A3(new_n23450_), .A4(new_n23768_), .ZN(new_n23917_));
  XNOR2_X1   g23724(.A1(new_n23917_), .A2(new_n23916_), .ZN(new_n23918_));
  NOR2_X1    g23725(.A1(new_n23439_), .A2(new_n5626_), .ZN(new_n23919_));
  NOR4_X1    g23726(.A1(new_n23863_), .A2(\asqrt[35] ), .A3(new_n23435_), .A4(new_n23761_), .ZN(new_n23920_));
  XNOR2_X1   g23727(.A1(new_n23920_), .A2(new_n23919_), .ZN(new_n23921_));
  INV_X1     g23728(.I(new_n23921_), .ZN(new_n23922_));
  NOR2_X1    g23729(.A1(new_n23424_), .A2(new_n6365_), .ZN(new_n23923_));
  NOR4_X1    g23730(.A1(new_n23863_), .A2(\asqrt[33] ), .A3(new_n23420_), .A4(new_n23754_), .ZN(new_n23924_));
  XNOR2_X1   g23731(.A1(new_n23924_), .A2(new_n23923_), .ZN(new_n23925_));
  NAND2_X1   g23732(.A1(new_n23747_), .A2(\asqrt[31] ), .ZN(new_n23926_));
  NOR4_X1    g23733(.A1(new_n23863_), .A2(\asqrt[31] ), .A3(new_n23405_), .A4(new_n23747_), .ZN(new_n23927_));
  XOR2_X1    g23734(.A1(new_n23927_), .A2(new_n23926_), .Z(new_n23928_));
  INV_X1     g23735(.I(new_n23928_), .ZN(new_n23929_));
  NAND2_X1   g23736(.A1(new_n23740_), .A2(\asqrt[29] ), .ZN(new_n23930_));
  NOR4_X1    g23737(.A1(new_n23863_), .A2(\asqrt[29] ), .A3(new_n23390_), .A4(new_n23740_), .ZN(new_n23931_));
  XOR2_X1    g23738(.A1(new_n23931_), .A2(new_n23930_), .Z(new_n23932_));
  NOR2_X1    g23739(.A1(new_n23379_), .A2(new_n8763_), .ZN(new_n23933_));
  NOR4_X1    g23740(.A1(new_n23863_), .A2(\asqrt[27] ), .A3(new_n23375_), .A4(new_n23733_), .ZN(new_n23934_));
  XNOR2_X1   g23741(.A1(new_n23934_), .A2(new_n23933_), .ZN(new_n23935_));
  INV_X1     g23742(.I(new_n23935_), .ZN(new_n23936_));
  NOR2_X1    g23743(.A1(new_n23364_), .A2(new_n9672_), .ZN(new_n23937_));
  NOR4_X1    g23744(.A1(new_n23863_), .A2(\asqrt[25] ), .A3(new_n23360_), .A4(new_n23726_), .ZN(new_n23938_));
  XNOR2_X1   g23745(.A1(new_n23938_), .A2(new_n23937_), .ZN(new_n23939_));
  NOR2_X1    g23746(.A1(new_n23349_), .A2(new_n10614_), .ZN(new_n23940_));
  NOR4_X1    g23747(.A1(new_n23863_), .A2(\asqrt[23] ), .A3(new_n23345_), .A4(new_n23719_), .ZN(new_n23941_));
  XNOR2_X1   g23748(.A1(new_n23941_), .A2(new_n23940_), .ZN(new_n23942_));
  INV_X1     g23749(.I(new_n23942_), .ZN(new_n23943_));
  NOR2_X1    g23750(.A1(new_n23334_), .A2(new_n11631_), .ZN(new_n23944_));
  NOR4_X1    g23751(.A1(new_n23863_), .A2(\asqrt[21] ), .A3(new_n23330_), .A4(new_n23712_), .ZN(new_n23945_));
  XNOR2_X1   g23752(.A1(new_n23945_), .A2(new_n23944_), .ZN(new_n23946_));
  NOR2_X1    g23753(.A1(new_n23319_), .A2(new_n12657_), .ZN(new_n23947_));
  NOR4_X1    g23754(.A1(new_n23863_), .A2(\asqrt[19] ), .A3(new_n23315_), .A4(new_n23705_), .ZN(new_n23948_));
  XNOR2_X1   g23755(.A1(new_n23948_), .A2(new_n23947_), .ZN(new_n23949_));
  INV_X1     g23756(.I(new_n23949_), .ZN(new_n23950_));
  NOR2_X1    g23757(.A1(new_n23304_), .A2(new_n13760_), .ZN(new_n23951_));
  NOR4_X1    g23758(.A1(new_n23863_), .A2(\asqrt[17] ), .A3(new_n23300_), .A4(new_n23698_), .ZN(new_n23952_));
  XNOR2_X1   g23759(.A1(new_n23952_), .A2(new_n23951_), .ZN(new_n23953_));
  NAND2_X1   g23760(.A1(new_n23691_), .A2(\asqrt[15] ), .ZN(new_n23954_));
  NOR4_X1    g23761(.A1(new_n23863_), .A2(\asqrt[15] ), .A3(new_n23285_), .A4(new_n23691_), .ZN(new_n23955_));
  XOR2_X1    g23762(.A1(new_n23955_), .A2(new_n23954_), .Z(new_n23956_));
  INV_X1     g23763(.I(new_n23956_), .ZN(new_n23957_));
  NAND2_X1   g23764(.A1(new_n23684_), .A2(\asqrt[13] ), .ZN(new_n23958_));
  NOR4_X1    g23765(.A1(new_n23863_), .A2(\asqrt[13] ), .A3(new_n23270_), .A4(new_n23684_), .ZN(new_n23959_));
  XOR2_X1    g23766(.A1(new_n23959_), .A2(new_n23958_), .Z(new_n23960_));
  NAND2_X1   g23767(.A1(new_n23677_), .A2(\asqrt[11] ), .ZN(new_n23961_));
  NOR4_X1    g23768(.A1(new_n23863_), .A2(\asqrt[11] ), .A3(new_n23255_), .A4(new_n23677_), .ZN(new_n23962_));
  XOR2_X1    g23769(.A1(new_n23962_), .A2(new_n23961_), .Z(new_n23963_));
  INV_X1     g23770(.I(new_n23963_), .ZN(new_n23964_));
  NOR2_X1    g23771(.A1(new_n23244_), .A2(new_n18495_), .ZN(new_n23965_));
  INV_X1     g23772(.I(new_n23965_), .ZN(new_n23966_));
  NOR4_X1    g23773(.A1(new_n23863_), .A2(\asqrt[9] ), .A3(new_n23240_), .A4(new_n23670_), .ZN(new_n23967_));
  XOR2_X1    g23774(.A1(new_n23967_), .A2(new_n23966_), .Z(new_n23968_));
  NOR2_X1    g23775(.A1(new_n23231_), .A2(new_n19782_), .ZN(new_n23969_));
  INV_X1     g23776(.I(new_n23969_), .ZN(new_n23970_));
  NOR4_X1    g23777(.A1(new_n23863_), .A2(\asqrt[7] ), .A3(new_n23227_), .A4(new_n23663_), .ZN(new_n23971_));
  XOR2_X1    g23778(.A1(new_n23971_), .A2(new_n23970_), .Z(new_n23972_));
  INV_X1     g23779(.I(new_n23972_), .ZN(new_n23973_));
  NAND2_X1   g23780(.A1(new_n23656_), .A2(\asqrt[5] ), .ZN(new_n23974_));
  NOR2_X1    g23781(.A1(new_n23652_), .A2(new_n23208_), .ZN(new_n23975_));
  NOR4_X1    g23782(.A1(new_n23863_), .A2(\asqrt[5] ), .A3(new_n23975_), .A4(new_n23656_), .ZN(new_n23976_));
  XOR2_X1    g23783(.A1(new_n23976_), .A2(new_n23974_), .Z(new_n23977_));
  AOI21_X1   g23784(.A1(\asqrt[2] ), .A2(new_n23641_), .B(\a[5] ), .ZN(new_n23978_));
  NOR2_X1    g23785(.A1(new_n23187_), .A2(\a[4] ), .ZN(new_n23979_));
  AOI21_X1   g23786(.A1(\asqrt[2] ), .A2(\a[4] ), .B(new_n23170_), .ZN(new_n23980_));
  OAI21_X1   g23787(.A1(new_n23979_), .A2(new_n23978_), .B(new_n23980_), .ZN(new_n23981_));
  NOR3_X1    g23788(.A1(new_n23863_), .A2(new_n23643_), .A3(new_n23981_), .ZN(new_n23982_));
  INV_X1     g23789(.I(new_n23636_), .ZN(new_n23983_));
  OAI21_X1   g23790(.A1(new_n23868_), .A2(new_n23983_), .B(new_n23864_), .ZN(new_n23984_));
  OAI21_X1   g23791(.A1(new_n23630_), .A2(new_n229_), .B(new_n23632_), .ZN(new_n23985_));
  NAND2_X1   g23792(.A1(new_n23985_), .A2(new_n23629_), .ZN(new_n23986_));
  INV_X1     g23793(.I(new_n23858_), .ZN(new_n23987_));
  OAI22_X1   g23794(.A1(new_n23630_), .A2(new_n229_), .B1(new_n23628_), .B2(new_n23623_), .ZN(new_n23988_));
  AOI21_X1   g23795(.A1(new_n23988_), .A2(\asqrt[62] ), .B(new_n23864_), .ZN(new_n23989_));
  AOI21_X1   g23796(.A1(new_n23989_), .A2(new_n23987_), .B(new_n23986_), .ZN(new_n23990_));
  NAND2_X1   g23797(.A1(new_n23990_), .A2(new_n23984_), .ZN(\asqrt[1] ));
  INV_X1     g23798(.I(new_n23981_), .ZN(new_n23992_));
  AOI21_X1   g23799(.A1(\asqrt[1] ), .A2(new_n23992_), .B(new_n23193_), .ZN(new_n23993_));
  OAI21_X1   g23800(.A1(new_n23982_), .A2(new_n23993_), .B(\asqrt[3] ), .ZN(new_n23994_));
  INV_X1     g23801(.I(\a[2] ), .ZN(new_n23995_));
  OAI21_X1   g23802(.A1(\a[0] ), .A2(\a[1] ), .B(new_n23995_), .ZN(new_n23996_));
  NOR2_X1    g23803(.A1(new_n23858_), .A2(new_n23995_), .ZN(new_n23997_));
  OAI21_X1   g23804(.A1(new_n23861_), .A2(new_n23997_), .B(new_n23855_), .ZN(new_n23998_));
  OAI21_X1   g23805(.A1(new_n23998_), .A2(new_n23637_), .B(new_n23996_), .ZN(new_n23999_));
  NAND2_X1   g23806(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n24000_));
  INV_X1     g23807(.I(new_n24000_), .ZN(new_n24001_));
  OAI21_X1   g23808(.A1(new_n23990_), .A2(new_n24001_), .B(new_n23637_), .ZN(new_n24002_));
  OR2_X2     g23809(.A1(new_n24002_), .A2(new_n23999_), .Z(new_n24003_));
  NAND2_X1   g23810(.A1(new_n24002_), .A2(new_n23999_), .ZN(new_n24004_));
  OAI21_X1   g23811(.A1(new_n23862_), .A2(new_n23637_), .B(new_n23169_), .ZN(new_n24005_));
  NOR2_X1    g23812(.A1(new_n24005_), .A2(new_n23158_), .ZN(new_n24006_));
  NAND2_X1   g23813(.A1(new_n24004_), .A2(new_n24006_), .ZN(new_n24007_));
  AND2_X2    g23814(.A1(new_n24007_), .A2(new_n24003_), .Z(new_n24008_));
  NAND3_X1   g23815(.A1(\asqrt[1] ), .A2(new_n23193_), .A3(new_n23992_), .ZN(new_n24009_));
  OAI21_X1   g23816(.A1(new_n23863_), .A2(new_n23981_), .B(new_n23643_), .ZN(new_n24010_));
  NAND2_X1   g23817(.A1(new_n24010_), .A2(new_n24009_), .ZN(new_n24011_));
  AOI21_X1   g23818(.A1(new_n23851_), .A2(new_n23854_), .B(new_n196_), .ZN(new_n24012_));
  NOR3_X1    g23819(.A1(new_n23855_), .A2(new_n24012_), .A3(new_n23160_), .ZN(new_n24013_));
  NOR2_X1    g23820(.A1(new_n23987_), .A2(new_n23158_), .ZN(new_n24014_));
  NAND3_X1   g23821(.A1(new_n23637_), .A2(new_n24013_), .A3(new_n24014_), .ZN(new_n24015_));
  AOI21_X1   g23822(.A1(new_n24005_), .A2(new_n24015_), .B(\a[4] ), .ZN(new_n24016_));
  AOI21_X1   g23823(.A1(new_n23990_), .A2(new_n23984_), .B(new_n23639_), .ZN(new_n24017_));
  OAI21_X1   g23824(.A1(new_n23629_), .A2(new_n23875_), .B(\asqrt[62] ), .ZN(new_n24018_));
  NAND4_X1   g23825(.A1(new_n23986_), .A2(new_n24018_), .A3(new_n23864_), .A4(new_n24014_), .ZN(new_n24019_));
  OAI21_X1   g23826(.A1(new_n23984_), .A2(new_n24019_), .B(\a[4] ), .ZN(new_n24020_));
  NOR2_X1    g23827(.A1(new_n24017_), .A2(new_n24020_), .ZN(new_n24021_));
  OAI22_X1   g23828(.A1(new_n24011_), .A2(\asqrt[3] ), .B1(new_n24016_), .B2(new_n24021_), .ZN(new_n24022_));
  AOI21_X1   g23829(.A1(new_n24008_), .A2(new_n23994_), .B(new_n24022_), .ZN(new_n24023_));
  NAND2_X1   g23830(.A1(new_n23203_), .A2(\asqrt[4] ), .ZN(new_n24024_));
  NOR2_X1    g23831(.A1(new_n23644_), .A2(new_n23645_), .ZN(new_n24025_));
  NOR4_X1    g23832(.A1(new_n23863_), .A2(\asqrt[4] ), .A3(new_n24025_), .A4(new_n23203_), .ZN(new_n24026_));
  XOR2_X1    g23833(.A1(new_n24026_), .A2(new_n24024_), .Z(new_n24027_));
  INV_X1     g23834(.I(new_n24027_), .ZN(new_n24028_));
  OAI21_X1   g23835(.A1(\asqrt[4] ), .A2(new_n24028_), .B(new_n24023_), .ZN(new_n24029_));
  NAND2_X1   g23836(.A1(new_n24029_), .A2(new_n23977_), .ZN(new_n24030_));
  NAND3_X1   g23837(.A1(new_n23994_), .A2(new_n24007_), .A3(new_n24003_), .ZN(new_n24031_));
  NOR2_X1    g23838(.A1(new_n24016_), .A2(new_n24021_), .ZN(new_n24032_));
  NOR3_X1    g23839(.A1(new_n23982_), .A2(new_n23993_), .A3(\asqrt[3] ), .ZN(new_n24033_));
  NOR2_X1    g23840(.A1(new_n24033_), .A2(new_n24032_), .ZN(new_n24034_));
  NAND2_X1   g23841(.A1(new_n24031_), .A2(new_n24034_), .ZN(new_n24035_));
  NOR2_X1    g23842(.A1(new_n24035_), .A2(new_n21781_), .ZN(new_n24036_));
  NAND2_X1   g23843(.A1(new_n24036_), .A2(\asqrt[5] ), .ZN(new_n24037_));
  INV_X1     g23844(.I(new_n24037_), .ZN(new_n24038_));
  NAND2_X1   g23845(.A1(new_n24030_), .A2(new_n24038_), .ZN(new_n24039_));
  OAI21_X1   g23846(.A1(new_n24029_), .A2(new_n23977_), .B(new_n21079_), .ZN(new_n24040_));
  NAND2_X1   g23847(.A1(new_n23224_), .A2(\asqrt[6] ), .ZN(new_n24041_));
  NAND2_X1   g23848(.A1(new_n23218_), .A2(new_n23219_), .ZN(new_n24042_));
  INV_X1     g23849(.I(new_n24042_), .ZN(new_n24043_));
  NOR4_X1    g23850(.A1(new_n23863_), .A2(\asqrt[6] ), .A3(new_n24043_), .A4(new_n23224_), .ZN(new_n24044_));
  XOR2_X1    g23851(.A1(new_n24044_), .A2(new_n24041_), .Z(new_n24045_));
  INV_X1     g23852(.I(new_n24045_), .ZN(new_n24046_));
  NAND3_X1   g23853(.A1(new_n24040_), .A2(new_n24036_), .A3(new_n24046_), .ZN(new_n24047_));
  AOI21_X1   g23854(.A1(new_n24047_), .A2(new_n20455_), .B(new_n24039_), .ZN(new_n24048_));
  NOR2_X1    g23855(.A1(new_n24048_), .A2(new_n23973_), .ZN(new_n24049_));
  AOI21_X1   g23856(.A1(new_n24040_), .A2(new_n24036_), .B(new_n24046_), .ZN(new_n24050_));
  NAND3_X1   g23857(.A1(new_n24030_), .A2(new_n24038_), .A3(\asqrt[6] ), .ZN(new_n24051_));
  NOR3_X1    g23858(.A1(new_n24050_), .A2(new_n24051_), .A3(new_n19782_), .ZN(new_n24052_));
  INV_X1     g23859(.I(new_n24052_), .ZN(new_n24053_));
  NOR2_X1    g23860(.A1(new_n24049_), .A2(new_n24053_), .ZN(new_n24054_));
  NOR2_X1    g23861(.A1(new_n24050_), .A2(new_n24051_), .ZN(new_n24055_));
  INV_X1     g23862(.I(new_n24055_), .ZN(new_n24056_));
  AOI21_X1   g23863(.A1(new_n24048_), .A2(new_n23973_), .B(\asqrt[7] ), .ZN(new_n24057_));
  NAND2_X1   g23864(.A1(new_n23238_), .A2(\asqrt[8] ), .ZN(new_n24058_));
  NOR4_X1    g23865(.A1(new_n23863_), .A2(\asqrt[8] ), .A3(new_n23233_), .A4(new_n23238_), .ZN(new_n24059_));
  XOR2_X1    g23866(.A1(new_n24059_), .A2(new_n24058_), .Z(new_n24060_));
  NOR3_X1    g23867(.A1(new_n24057_), .A2(new_n24056_), .A3(new_n24060_), .ZN(new_n24061_));
  OAI21_X1   g23868(.A1(new_n24061_), .A2(\asqrt[8] ), .B(new_n24054_), .ZN(new_n24062_));
  NAND2_X1   g23869(.A1(new_n24062_), .A2(new_n23968_), .ZN(new_n24063_));
  OAI21_X1   g23870(.A1(new_n24057_), .A2(new_n24056_), .B(new_n24060_), .ZN(new_n24064_));
  NOR3_X1    g23871(.A1(new_n24049_), .A2(new_n24053_), .A3(new_n19100_), .ZN(new_n24065_));
  NAND3_X1   g23872(.A1(new_n24064_), .A2(new_n24065_), .A3(\asqrt[9] ), .ZN(new_n24066_));
  INV_X1     g23873(.I(new_n24066_), .ZN(new_n24067_));
  NAND2_X1   g23874(.A1(new_n24063_), .A2(new_n24067_), .ZN(new_n24068_));
  NAND2_X1   g23875(.A1(new_n24064_), .A2(new_n24065_), .ZN(new_n24069_));
  INV_X1     g23876(.I(new_n24069_), .ZN(new_n24070_));
  OAI21_X1   g23877(.A1(new_n24062_), .A2(new_n23968_), .B(new_n18495_), .ZN(new_n24071_));
  NAND2_X1   g23878(.A1(new_n23252_), .A2(\asqrt[10] ), .ZN(new_n24072_));
  NOR4_X1    g23879(.A1(new_n23863_), .A2(\asqrt[10] ), .A3(new_n23247_), .A4(new_n23252_), .ZN(new_n24073_));
  XOR2_X1    g23880(.A1(new_n24073_), .A2(new_n24072_), .Z(new_n24074_));
  INV_X1     g23881(.I(new_n24074_), .ZN(new_n24075_));
  NAND3_X1   g23882(.A1(new_n24071_), .A2(new_n24070_), .A3(new_n24075_), .ZN(new_n24076_));
  AOI21_X1   g23883(.A1(new_n24076_), .A2(new_n17893_), .B(new_n24068_), .ZN(new_n24077_));
  NOR2_X1    g23884(.A1(new_n24077_), .A2(new_n23964_), .ZN(new_n24078_));
  AOI21_X1   g23885(.A1(new_n24071_), .A2(new_n24070_), .B(new_n24075_), .ZN(new_n24079_));
  NAND3_X1   g23886(.A1(new_n24063_), .A2(new_n24067_), .A3(\asqrt[10] ), .ZN(new_n24080_));
  NOR3_X1    g23887(.A1(new_n24079_), .A2(new_n24080_), .A3(new_n17271_), .ZN(new_n24081_));
  INV_X1     g23888(.I(new_n24081_), .ZN(new_n24082_));
  NOR2_X1    g23889(.A1(new_n24078_), .A2(new_n24082_), .ZN(new_n24083_));
  NOR2_X1    g23890(.A1(new_n24079_), .A2(new_n24080_), .ZN(new_n24084_));
  INV_X1     g23891(.I(new_n24084_), .ZN(new_n24085_));
  AOI21_X1   g23892(.A1(new_n24077_), .A2(new_n23964_), .B(\asqrt[11] ), .ZN(new_n24086_));
  NOR2_X1    g23893(.A1(new_n23680_), .A2(new_n16619_), .ZN(new_n24087_));
  NOR4_X1    g23894(.A1(new_n23863_), .A2(\asqrt[12] ), .A3(new_n23262_), .A4(new_n23267_), .ZN(new_n24088_));
  XNOR2_X1   g23895(.A1(new_n24088_), .A2(new_n24087_), .ZN(new_n24089_));
  NOR3_X1    g23896(.A1(new_n24086_), .A2(new_n24085_), .A3(new_n24089_), .ZN(new_n24090_));
  OAI21_X1   g23897(.A1(new_n24090_), .A2(\asqrt[12] ), .B(new_n24083_), .ZN(new_n24091_));
  NAND2_X1   g23898(.A1(new_n24091_), .A2(new_n23960_), .ZN(new_n24092_));
  OAI21_X1   g23899(.A1(new_n24086_), .A2(new_n24085_), .B(new_n24089_), .ZN(new_n24093_));
  NOR3_X1    g23900(.A1(new_n24078_), .A2(new_n24082_), .A3(new_n16619_), .ZN(new_n24094_));
  NAND3_X1   g23901(.A1(new_n24093_), .A2(new_n24094_), .A3(\asqrt[13] ), .ZN(new_n24095_));
  INV_X1     g23902(.I(new_n24095_), .ZN(new_n24096_));
  NAND2_X1   g23903(.A1(new_n24092_), .A2(new_n24096_), .ZN(new_n24097_));
  NAND2_X1   g23904(.A1(new_n24093_), .A2(new_n24094_), .ZN(new_n24098_));
  INV_X1     g23905(.I(new_n24098_), .ZN(new_n24099_));
  OAI21_X1   g23906(.A1(new_n24091_), .A2(new_n23960_), .B(new_n16060_), .ZN(new_n24100_));
  NAND2_X1   g23907(.A1(new_n23282_), .A2(\asqrt[14] ), .ZN(new_n24101_));
  NOR4_X1    g23908(.A1(new_n23863_), .A2(\asqrt[14] ), .A3(new_n23277_), .A4(new_n23282_), .ZN(new_n24102_));
  XOR2_X1    g23909(.A1(new_n24102_), .A2(new_n24101_), .Z(new_n24103_));
  INV_X1     g23910(.I(new_n24103_), .ZN(new_n24104_));
  NAND3_X1   g23911(.A1(new_n24100_), .A2(new_n24099_), .A3(new_n24104_), .ZN(new_n24105_));
  AOI21_X1   g23912(.A1(new_n24105_), .A2(new_n15447_), .B(new_n24097_), .ZN(new_n24106_));
  NOR2_X1    g23913(.A1(new_n24106_), .A2(new_n23957_), .ZN(new_n24107_));
  AOI21_X1   g23914(.A1(new_n24100_), .A2(new_n24099_), .B(new_n24104_), .ZN(new_n24108_));
  NAND3_X1   g23915(.A1(new_n24092_), .A2(new_n24096_), .A3(\asqrt[14] ), .ZN(new_n24109_));
  NOR3_X1    g23916(.A1(new_n24108_), .A2(new_n24109_), .A3(new_n14871_), .ZN(new_n24110_));
  INV_X1     g23917(.I(new_n24110_), .ZN(new_n24111_));
  NOR2_X1    g23918(.A1(new_n24107_), .A2(new_n24111_), .ZN(new_n24112_));
  NOR2_X1    g23919(.A1(new_n24108_), .A2(new_n24109_), .ZN(new_n24113_));
  INV_X1     g23920(.I(new_n24113_), .ZN(new_n24114_));
  AOI21_X1   g23921(.A1(new_n24106_), .A2(new_n23957_), .B(\asqrt[15] ), .ZN(new_n24115_));
  NAND2_X1   g23922(.A1(new_n23297_), .A2(\asqrt[16] ), .ZN(new_n24116_));
  NOR4_X1    g23923(.A1(new_n23863_), .A2(\asqrt[16] ), .A3(new_n23292_), .A4(new_n23297_), .ZN(new_n24117_));
  XOR2_X1    g23924(.A1(new_n24117_), .A2(new_n24116_), .Z(new_n24118_));
  NOR3_X1    g23925(.A1(new_n24115_), .A2(new_n24114_), .A3(new_n24118_), .ZN(new_n24119_));
  OAI21_X1   g23926(.A1(new_n24119_), .A2(\asqrt[16] ), .B(new_n24112_), .ZN(new_n24120_));
  NAND2_X1   g23927(.A1(new_n24120_), .A2(new_n23953_), .ZN(new_n24121_));
  OAI21_X1   g23928(.A1(new_n24115_), .A2(new_n24114_), .B(new_n24118_), .ZN(new_n24122_));
  NOR3_X1    g23929(.A1(new_n24107_), .A2(new_n24111_), .A3(new_n14273_), .ZN(new_n24123_));
  NAND3_X1   g23930(.A1(new_n24122_), .A2(new_n24123_), .A3(\asqrt[17] ), .ZN(new_n24124_));
  INV_X1     g23931(.I(new_n24124_), .ZN(new_n24125_));
  NAND2_X1   g23932(.A1(new_n24121_), .A2(new_n24125_), .ZN(new_n24126_));
  NAND2_X1   g23933(.A1(new_n24122_), .A2(new_n24123_), .ZN(new_n24127_));
  INV_X1     g23934(.I(new_n24127_), .ZN(new_n24128_));
  OAI21_X1   g23935(.A1(new_n24120_), .A2(new_n23953_), .B(new_n13760_), .ZN(new_n24129_));
  NAND2_X1   g23936(.A1(new_n23312_), .A2(\asqrt[18] ), .ZN(new_n24130_));
  NOR4_X1    g23937(.A1(new_n23863_), .A2(\asqrt[18] ), .A3(new_n23307_), .A4(new_n23312_), .ZN(new_n24131_));
  XOR2_X1    g23938(.A1(new_n24131_), .A2(new_n24130_), .Z(new_n24132_));
  INV_X1     g23939(.I(new_n24132_), .ZN(new_n24133_));
  NAND3_X1   g23940(.A1(new_n24129_), .A2(new_n24128_), .A3(new_n24133_), .ZN(new_n24134_));
  AOI21_X1   g23941(.A1(new_n24134_), .A2(new_n13192_), .B(new_n24126_), .ZN(new_n24135_));
  NOR2_X1    g23942(.A1(new_n24135_), .A2(new_n23950_), .ZN(new_n24136_));
  AOI21_X1   g23943(.A1(new_n24129_), .A2(new_n24128_), .B(new_n24133_), .ZN(new_n24137_));
  NAND3_X1   g23944(.A1(new_n24121_), .A2(new_n24125_), .A3(\asqrt[18] ), .ZN(new_n24138_));
  NOR3_X1    g23945(.A1(new_n24137_), .A2(new_n24138_), .A3(new_n12657_), .ZN(new_n24139_));
  INV_X1     g23946(.I(new_n24139_), .ZN(new_n24140_));
  NOR2_X1    g23947(.A1(new_n24136_), .A2(new_n24140_), .ZN(new_n24141_));
  NOR2_X1    g23948(.A1(new_n24137_), .A2(new_n24138_), .ZN(new_n24142_));
  INV_X1     g23949(.I(new_n24142_), .ZN(new_n24143_));
  AOI21_X1   g23950(.A1(new_n24135_), .A2(new_n23950_), .B(\asqrt[19] ), .ZN(new_n24144_));
  NAND2_X1   g23951(.A1(new_n23327_), .A2(\asqrt[20] ), .ZN(new_n24145_));
  NOR4_X1    g23952(.A1(new_n23863_), .A2(\asqrt[20] ), .A3(new_n23322_), .A4(new_n23327_), .ZN(new_n24146_));
  XOR2_X1    g23953(.A1(new_n24146_), .A2(new_n24145_), .Z(new_n24147_));
  NOR3_X1    g23954(.A1(new_n24144_), .A2(new_n24143_), .A3(new_n24147_), .ZN(new_n24148_));
  OAI21_X1   g23955(.A1(new_n24148_), .A2(\asqrt[20] ), .B(new_n24141_), .ZN(new_n24149_));
  NAND2_X1   g23956(.A1(new_n24149_), .A2(new_n23946_), .ZN(new_n24150_));
  OAI21_X1   g23957(.A1(new_n24144_), .A2(new_n24143_), .B(new_n24147_), .ZN(new_n24151_));
  NOR3_X1    g23958(.A1(new_n24136_), .A2(new_n24140_), .A3(new_n12101_), .ZN(new_n24152_));
  NAND3_X1   g23959(.A1(new_n24151_), .A2(new_n24152_), .A3(\asqrt[21] ), .ZN(new_n24153_));
  INV_X1     g23960(.I(new_n24153_), .ZN(new_n24154_));
  NAND2_X1   g23961(.A1(new_n24150_), .A2(new_n24154_), .ZN(new_n24155_));
  NAND2_X1   g23962(.A1(new_n24151_), .A2(new_n24152_), .ZN(new_n24156_));
  INV_X1     g23963(.I(new_n24156_), .ZN(new_n24157_));
  OAI21_X1   g23964(.A1(new_n24149_), .A2(new_n23946_), .B(new_n11631_), .ZN(new_n24158_));
  NAND2_X1   g23965(.A1(new_n23342_), .A2(\asqrt[22] ), .ZN(new_n24159_));
  NOR4_X1    g23966(.A1(new_n23863_), .A2(\asqrt[22] ), .A3(new_n23337_), .A4(new_n23342_), .ZN(new_n24160_));
  XOR2_X1    g23967(.A1(new_n24160_), .A2(new_n24159_), .Z(new_n24161_));
  INV_X1     g23968(.I(new_n24161_), .ZN(new_n24162_));
  NAND3_X1   g23969(.A1(new_n24158_), .A2(new_n24157_), .A3(new_n24162_), .ZN(new_n24163_));
  AOI21_X1   g23970(.A1(new_n24163_), .A2(new_n11105_), .B(new_n24155_), .ZN(new_n24164_));
  NOR2_X1    g23971(.A1(new_n24164_), .A2(new_n23943_), .ZN(new_n24165_));
  AOI21_X1   g23972(.A1(new_n24158_), .A2(new_n24157_), .B(new_n24162_), .ZN(new_n24166_));
  NAND3_X1   g23973(.A1(new_n24150_), .A2(new_n24154_), .A3(\asqrt[22] ), .ZN(new_n24167_));
  NOR3_X1    g23974(.A1(new_n24166_), .A2(new_n24167_), .A3(new_n10614_), .ZN(new_n24168_));
  INV_X1     g23975(.I(new_n24168_), .ZN(new_n24169_));
  NOR2_X1    g23976(.A1(new_n24165_), .A2(new_n24169_), .ZN(new_n24170_));
  NOR2_X1    g23977(.A1(new_n24166_), .A2(new_n24167_), .ZN(new_n24171_));
  INV_X1     g23978(.I(new_n24171_), .ZN(new_n24172_));
  AOI21_X1   g23979(.A1(new_n24164_), .A2(new_n23943_), .B(\asqrt[23] ), .ZN(new_n24173_));
  NAND2_X1   g23980(.A1(new_n23357_), .A2(\asqrt[24] ), .ZN(new_n24174_));
  NOR4_X1    g23981(.A1(new_n23863_), .A2(\asqrt[24] ), .A3(new_n23352_), .A4(new_n23357_), .ZN(new_n24175_));
  XOR2_X1    g23982(.A1(new_n24175_), .A2(new_n24174_), .Z(new_n24176_));
  NOR3_X1    g23983(.A1(new_n24173_), .A2(new_n24172_), .A3(new_n24176_), .ZN(new_n24177_));
  OAI21_X1   g23984(.A1(new_n24177_), .A2(\asqrt[24] ), .B(new_n24170_), .ZN(new_n24178_));
  NAND2_X1   g23985(.A1(new_n24178_), .A2(new_n23939_), .ZN(new_n24179_));
  OAI21_X1   g23986(.A1(new_n24173_), .A2(new_n24172_), .B(new_n24176_), .ZN(new_n24180_));
  NOR3_X1    g23987(.A1(new_n24165_), .A2(new_n24169_), .A3(new_n10104_), .ZN(new_n24181_));
  NAND3_X1   g23988(.A1(new_n24180_), .A2(new_n24181_), .A3(\asqrt[25] ), .ZN(new_n24182_));
  INV_X1     g23989(.I(new_n24182_), .ZN(new_n24183_));
  NAND2_X1   g23990(.A1(new_n24179_), .A2(new_n24183_), .ZN(new_n24184_));
  NAND2_X1   g23991(.A1(new_n24180_), .A2(new_n24181_), .ZN(new_n24185_));
  INV_X1     g23992(.I(new_n24185_), .ZN(new_n24186_));
  OAI21_X1   g23993(.A1(new_n24178_), .A2(new_n23939_), .B(new_n9672_), .ZN(new_n24187_));
  NAND2_X1   g23994(.A1(new_n23372_), .A2(\asqrt[26] ), .ZN(new_n24188_));
  NOR4_X1    g23995(.A1(new_n23863_), .A2(\asqrt[26] ), .A3(new_n23367_), .A4(new_n23372_), .ZN(new_n24189_));
  XOR2_X1    g23996(.A1(new_n24189_), .A2(new_n24188_), .Z(new_n24190_));
  INV_X1     g23997(.I(new_n24190_), .ZN(new_n24191_));
  NAND3_X1   g23998(.A1(new_n24187_), .A2(new_n24186_), .A3(new_n24191_), .ZN(new_n24192_));
  AOI21_X1   g23999(.A1(new_n24192_), .A2(new_n9212_), .B(new_n24184_), .ZN(new_n24193_));
  NOR2_X1    g24000(.A1(new_n24193_), .A2(new_n23936_), .ZN(new_n24194_));
  AOI21_X1   g24001(.A1(new_n24187_), .A2(new_n24186_), .B(new_n24191_), .ZN(new_n24195_));
  NAND3_X1   g24002(.A1(new_n24179_), .A2(new_n24183_), .A3(\asqrt[26] ), .ZN(new_n24196_));
  NOR3_X1    g24003(.A1(new_n24195_), .A2(new_n24196_), .A3(new_n8763_), .ZN(new_n24197_));
  INV_X1     g24004(.I(new_n24197_), .ZN(new_n24198_));
  NOR2_X1    g24005(.A1(new_n24194_), .A2(new_n24198_), .ZN(new_n24199_));
  NOR2_X1    g24006(.A1(new_n24195_), .A2(new_n24196_), .ZN(new_n24200_));
  INV_X1     g24007(.I(new_n24200_), .ZN(new_n24201_));
  AOI21_X1   g24008(.A1(new_n24193_), .A2(new_n23936_), .B(\asqrt[27] ), .ZN(new_n24202_));
  NAND2_X1   g24009(.A1(new_n23387_), .A2(\asqrt[28] ), .ZN(new_n24203_));
  NOR4_X1    g24010(.A1(new_n23863_), .A2(\asqrt[28] ), .A3(new_n23382_), .A4(new_n23387_), .ZN(new_n24204_));
  XOR2_X1    g24011(.A1(new_n24204_), .A2(new_n24203_), .Z(new_n24205_));
  NOR3_X1    g24012(.A1(new_n24202_), .A2(new_n24201_), .A3(new_n24205_), .ZN(new_n24206_));
  OAI21_X1   g24013(.A1(new_n24206_), .A2(\asqrt[28] ), .B(new_n24199_), .ZN(new_n24207_));
  NAND2_X1   g24014(.A1(new_n24207_), .A2(new_n23932_), .ZN(new_n24208_));
  OAI21_X1   g24015(.A1(new_n24202_), .A2(new_n24201_), .B(new_n24205_), .ZN(new_n24209_));
  NOR3_X1    g24016(.A1(new_n24194_), .A2(new_n24198_), .A3(new_n8319_), .ZN(new_n24210_));
  NAND3_X1   g24017(.A1(new_n24209_), .A2(new_n24210_), .A3(\asqrt[29] ), .ZN(new_n24211_));
  INV_X1     g24018(.I(new_n24211_), .ZN(new_n24212_));
  NAND2_X1   g24019(.A1(new_n24208_), .A2(new_n24212_), .ZN(new_n24213_));
  NAND2_X1   g24020(.A1(new_n24209_), .A2(new_n24210_), .ZN(new_n24214_));
  INV_X1     g24021(.I(new_n24214_), .ZN(new_n24215_));
  OAI21_X1   g24022(.A1(new_n24207_), .A2(new_n23932_), .B(new_n7931_), .ZN(new_n24216_));
  NOR2_X1    g24023(.A1(new_n23743_), .A2(new_n7517_), .ZN(new_n24217_));
  NOR4_X1    g24024(.A1(new_n23863_), .A2(\asqrt[30] ), .A3(new_n23397_), .A4(new_n23402_), .ZN(new_n24218_));
  XNOR2_X1   g24025(.A1(new_n24218_), .A2(new_n24217_), .ZN(new_n24219_));
  INV_X1     g24026(.I(new_n24219_), .ZN(new_n24220_));
  NAND3_X1   g24027(.A1(new_n24216_), .A2(new_n24215_), .A3(new_n24220_), .ZN(new_n24221_));
  AOI21_X1   g24028(.A1(new_n24221_), .A2(new_n7517_), .B(new_n24213_), .ZN(new_n24222_));
  NOR2_X1    g24029(.A1(new_n24222_), .A2(new_n23929_), .ZN(new_n24223_));
  AOI21_X1   g24030(.A1(new_n24216_), .A2(new_n24215_), .B(new_n24220_), .ZN(new_n24224_));
  NAND3_X1   g24031(.A1(new_n24208_), .A2(new_n24212_), .A3(\asqrt[30] ), .ZN(new_n24225_));
  NOR3_X1    g24032(.A1(new_n24224_), .A2(new_n24225_), .A3(new_n7110_), .ZN(new_n24226_));
  INV_X1     g24033(.I(new_n24226_), .ZN(new_n24227_));
  NOR2_X1    g24034(.A1(new_n24223_), .A2(new_n24227_), .ZN(new_n24228_));
  NOR2_X1    g24035(.A1(new_n24224_), .A2(new_n24225_), .ZN(new_n24229_));
  INV_X1     g24036(.I(new_n24229_), .ZN(new_n24230_));
  AOI21_X1   g24037(.A1(new_n24222_), .A2(new_n23929_), .B(\asqrt[31] ), .ZN(new_n24231_));
  NOR2_X1    g24038(.A1(new_n23750_), .A2(new_n6708_), .ZN(new_n24232_));
  NOR4_X1    g24039(.A1(new_n23863_), .A2(\asqrt[32] ), .A3(new_n23412_), .A4(new_n23417_), .ZN(new_n24233_));
  XNOR2_X1   g24040(.A1(new_n24233_), .A2(new_n24232_), .ZN(new_n24234_));
  NOR3_X1    g24041(.A1(new_n24231_), .A2(new_n24230_), .A3(new_n24234_), .ZN(new_n24235_));
  OAI21_X1   g24042(.A1(new_n24235_), .A2(\asqrt[32] ), .B(new_n24228_), .ZN(new_n24236_));
  NAND2_X1   g24043(.A1(new_n24236_), .A2(new_n23925_), .ZN(new_n24237_));
  OAI21_X1   g24044(.A1(new_n24231_), .A2(new_n24230_), .B(new_n24234_), .ZN(new_n24238_));
  NOR3_X1    g24045(.A1(new_n24223_), .A2(new_n24227_), .A3(new_n6708_), .ZN(new_n24239_));
  NAND3_X1   g24046(.A1(new_n24238_), .A2(new_n24239_), .A3(\asqrt[33] ), .ZN(new_n24240_));
  INV_X1     g24047(.I(new_n24240_), .ZN(new_n24241_));
  NAND2_X1   g24048(.A1(new_n24237_), .A2(new_n24241_), .ZN(new_n24242_));
  NAND2_X1   g24049(.A1(new_n24238_), .A2(new_n24239_), .ZN(new_n24243_));
  INV_X1     g24050(.I(new_n24243_), .ZN(new_n24244_));
  OAI21_X1   g24051(.A1(new_n24236_), .A2(new_n23925_), .B(new_n6365_), .ZN(new_n24245_));
  NAND2_X1   g24052(.A1(new_n23432_), .A2(\asqrt[34] ), .ZN(new_n24246_));
  NOR4_X1    g24053(.A1(new_n23863_), .A2(\asqrt[34] ), .A3(new_n23427_), .A4(new_n23432_), .ZN(new_n24247_));
  XOR2_X1    g24054(.A1(new_n24247_), .A2(new_n24246_), .Z(new_n24248_));
  INV_X1     g24055(.I(new_n24248_), .ZN(new_n24249_));
  NAND3_X1   g24056(.A1(new_n24245_), .A2(new_n24244_), .A3(new_n24249_), .ZN(new_n24250_));
  AOI21_X1   g24057(.A1(new_n24250_), .A2(new_n5991_), .B(new_n24242_), .ZN(new_n24251_));
  NOR2_X1    g24058(.A1(new_n24251_), .A2(new_n23922_), .ZN(new_n24252_));
  AOI21_X1   g24059(.A1(new_n24245_), .A2(new_n24244_), .B(new_n24249_), .ZN(new_n24253_));
  NAND3_X1   g24060(.A1(new_n24237_), .A2(new_n24241_), .A3(\asqrt[34] ), .ZN(new_n24254_));
  NOR3_X1    g24061(.A1(new_n24253_), .A2(new_n24254_), .A3(new_n5626_), .ZN(new_n24255_));
  INV_X1     g24062(.I(new_n24255_), .ZN(new_n24256_));
  NOR2_X1    g24063(.A1(new_n24252_), .A2(new_n24256_), .ZN(new_n24257_));
  NOR2_X1    g24064(.A1(new_n24253_), .A2(new_n24254_), .ZN(new_n24258_));
  INV_X1     g24065(.I(new_n24258_), .ZN(new_n24259_));
  AOI21_X1   g24066(.A1(new_n24251_), .A2(new_n23922_), .B(\asqrt[35] ), .ZN(new_n24260_));
  NAND2_X1   g24067(.A1(new_n23447_), .A2(\asqrt[36] ), .ZN(new_n24261_));
  NOR4_X1    g24068(.A1(new_n23863_), .A2(\asqrt[36] ), .A3(new_n23442_), .A4(new_n23447_), .ZN(new_n24262_));
  XOR2_X1    g24069(.A1(new_n24262_), .A2(new_n24261_), .Z(new_n24263_));
  NOR3_X1    g24070(.A1(new_n24260_), .A2(new_n24259_), .A3(new_n24263_), .ZN(new_n24264_));
  OAI21_X1   g24071(.A1(new_n24264_), .A2(\asqrt[36] ), .B(new_n24257_), .ZN(new_n24265_));
  NAND2_X1   g24072(.A1(new_n24265_), .A2(new_n23918_), .ZN(new_n24266_));
  OAI21_X1   g24073(.A1(new_n24260_), .A2(new_n24259_), .B(new_n24263_), .ZN(new_n24267_));
  NOR3_X1    g24074(.A1(new_n24252_), .A2(new_n24256_), .A3(new_n5273_), .ZN(new_n24268_));
  NAND3_X1   g24075(.A1(new_n24267_), .A2(new_n24268_), .A3(\asqrt[37] ), .ZN(new_n24269_));
  INV_X1     g24076(.I(new_n24269_), .ZN(new_n24270_));
  NAND2_X1   g24077(.A1(new_n24266_), .A2(new_n24270_), .ZN(new_n24271_));
  NAND2_X1   g24078(.A1(new_n24267_), .A2(new_n24268_), .ZN(new_n24272_));
  INV_X1     g24079(.I(new_n24272_), .ZN(new_n24273_));
  OAI21_X1   g24080(.A1(new_n24265_), .A2(new_n23918_), .B(new_n4973_), .ZN(new_n24274_));
  NAND2_X1   g24081(.A1(new_n23462_), .A2(\asqrt[38] ), .ZN(new_n24275_));
  NOR4_X1    g24082(.A1(new_n23863_), .A2(\asqrt[38] ), .A3(new_n23457_), .A4(new_n23462_), .ZN(new_n24276_));
  XOR2_X1    g24083(.A1(new_n24276_), .A2(new_n24275_), .Z(new_n24277_));
  INV_X1     g24084(.I(new_n24277_), .ZN(new_n24278_));
  NAND3_X1   g24085(.A1(new_n24274_), .A2(new_n24273_), .A3(new_n24278_), .ZN(new_n24279_));
  AOI21_X1   g24086(.A1(new_n24279_), .A2(new_n4645_), .B(new_n24271_), .ZN(new_n24280_));
  NOR2_X1    g24087(.A1(new_n24280_), .A2(new_n23915_), .ZN(new_n24281_));
  AOI21_X1   g24088(.A1(new_n24274_), .A2(new_n24273_), .B(new_n24278_), .ZN(new_n24282_));
  NAND3_X1   g24089(.A1(new_n24266_), .A2(new_n24270_), .A3(\asqrt[38] ), .ZN(new_n24283_));
  NOR3_X1    g24090(.A1(new_n24282_), .A2(new_n24283_), .A3(new_n4330_), .ZN(new_n24284_));
  INV_X1     g24091(.I(new_n24284_), .ZN(new_n24285_));
  NOR2_X1    g24092(.A1(new_n24281_), .A2(new_n24285_), .ZN(new_n24286_));
  NOR2_X1    g24093(.A1(new_n24282_), .A2(new_n24283_), .ZN(new_n24287_));
  INV_X1     g24094(.I(new_n24287_), .ZN(new_n24288_));
  AOI21_X1   g24095(.A1(new_n24280_), .A2(new_n23915_), .B(\asqrt[39] ), .ZN(new_n24289_));
  NOR2_X1    g24096(.A1(new_n23778_), .A2(new_n4018_), .ZN(new_n24290_));
  NOR4_X1    g24097(.A1(new_n23863_), .A2(\asqrt[40] ), .A3(new_n23472_), .A4(new_n23477_), .ZN(new_n24291_));
  XNOR2_X1   g24098(.A1(new_n24291_), .A2(new_n24290_), .ZN(new_n24292_));
  NOR3_X1    g24099(.A1(new_n24289_), .A2(new_n24288_), .A3(new_n24292_), .ZN(new_n24293_));
  OAI21_X1   g24100(.A1(new_n24293_), .A2(\asqrt[40] ), .B(new_n24286_), .ZN(new_n24294_));
  NAND2_X1   g24101(.A1(new_n24294_), .A2(new_n23911_), .ZN(new_n24295_));
  OAI21_X1   g24102(.A1(new_n24289_), .A2(new_n24288_), .B(new_n24292_), .ZN(new_n24296_));
  NOR3_X1    g24103(.A1(new_n24281_), .A2(new_n24285_), .A3(new_n4018_), .ZN(new_n24297_));
  NAND3_X1   g24104(.A1(new_n24296_), .A2(new_n24297_), .A3(\asqrt[41] ), .ZN(new_n24298_));
  INV_X1     g24105(.I(new_n24298_), .ZN(new_n24299_));
  NAND2_X1   g24106(.A1(new_n24295_), .A2(new_n24299_), .ZN(new_n24300_));
  NAND2_X1   g24107(.A1(new_n24296_), .A2(new_n24297_), .ZN(new_n24301_));
  INV_X1     g24108(.I(new_n24301_), .ZN(new_n24302_));
  OAI21_X1   g24109(.A1(new_n24294_), .A2(new_n23911_), .B(new_n3760_), .ZN(new_n24303_));
  NOR2_X1    g24110(.A1(new_n23785_), .A2(new_n3481_), .ZN(new_n24304_));
  NOR4_X1    g24111(.A1(new_n23863_), .A2(\asqrt[42] ), .A3(new_n23487_), .A4(new_n23492_), .ZN(new_n24305_));
  XNOR2_X1   g24112(.A1(new_n24305_), .A2(new_n24304_), .ZN(new_n24306_));
  INV_X1     g24113(.I(new_n24306_), .ZN(new_n24307_));
  NAND3_X1   g24114(.A1(new_n24303_), .A2(new_n24302_), .A3(new_n24307_), .ZN(new_n24308_));
  AOI21_X1   g24115(.A1(new_n24308_), .A2(new_n3481_), .B(new_n24300_), .ZN(new_n24309_));
  NOR2_X1    g24116(.A1(new_n24309_), .A2(new_n23908_), .ZN(new_n24310_));
  AOI21_X1   g24117(.A1(new_n24303_), .A2(new_n24302_), .B(new_n24307_), .ZN(new_n24311_));
  NAND3_X1   g24118(.A1(new_n24295_), .A2(new_n24299_), .A3(\asqrt[42] ), .ZN(new_n24312_));
  NOR3_X1    g24119(.A1(new_n24311_), .A2(new_n24312_), .A3(new_n3208_), .ZN(new_n24313_));
  INV_X1     g24120(.I(new_n24313_), .ZN(new_n24314_));
  NOR2_X1    g24121(.A1(new_n24310_), .A2(new_n24314_), .ZN(new_n24315_));
  NOR2_X1    g24122(.A1(new_n24311_), .A2(new_n24312_), .ZN(new_n24316_));
  INV_X1     g24123(.I(new_n24316_), .ZN(new_n24317_));
  AOI21_X1   g24124(.A1(new_n24309_), .A2(new_n23908_), .B(\asqrt[43] ), .ZN(new_n24318_));
  NOR2_X1    g24125(.A1(new_n23792_), .A2(new_n2941_), .ZN(new_n24319_));
  NOR4_X1    g24126(.A1(new_n23863_), .A2(\asqrt[44] ), .A3(new_n23502_), .A4(new_n23507_), .ZN(new_n24320_));
  XNOR2_X1   g24127(.A1(new_n24320_), .A2(new_n24319_), .ZN(new_n24321_));
  NOR3_X1    g24128(.A1(new_n24318_), .A2(new_n24317_), .A3(new_n24321_), .ZN(new_n24322_));
  OAI21_X1   g24129(.A1(new_n24322_), .A2(\asqrt[44] ), .B(new_n24315_), .ZN(new_n24323_));
  NAND2_X1   g24130(.A1(new_n24323_), .A2(new_n23904_), .ZN(new_n24324_));
  OAI21_X1   g24131(.A1(new_n24318_), .A2(new_n24317_), .B(new_n24321_), .ZN(new_n24325_));
  NOR3_X1    g24132(.A1(new_n24310_), .A2(new_n24314_), .A3(new_n2941_), .ZN(new_n24326_));
  NAND3_X1   g24133(.A1(new_n24325_), .A2(new_n24326_), .A3(\asqrt[45] ), .ZN(new_n24327_));
  INV_X1     g24134(.I(new_n24327_), .ZN(new_n24328_));
  NAND2_X1   g24135(.A1(new_n24324_), .A2(new_n24328_), .ZN(new_n24329_));
  NAND2_X1   g24136(.A1(new_n24325_), .A2(new_n24326_), .ZN(new_n24330_));
  INV_X1     g24137(.I(new_n24330_), .ZN(new_n24331_));
  OAI21_X1   g24138(.A1(new_n24323_), .A2(new_n23904_), .B(new_n2728_), .ZN(new_n24332_));
  NAND2_X1   g24139(.A1(new_n23522_), .A2(\asqrt[46] ), .ZN(new_n24333_));
  NOR4_X1    g24140(.A1(new_n23863_), .A2(\asqrt[46] ), .A3(new_n23517_), .A4(new_n23522_), .ZN(new_n24334_));
  XOR2_X1    g24141(.A1(new_n24334_), .A2(new_n24333_), .Z(new_n24335_));
  INV_X1     g24142(.I(new_n24335_), .ZN(new_n24336_));
  NAND3_X1   g24143(.A1(new_n24332_), .A2(new_n24331_), .A3(new_n24336_), .ZN(new_n24337_));
  AOI21_X1   g24144(.A1(new_n24337_), .A2(new_n2488_), .B(new_n24329_), .ZN(new_n24338_));
  NOR2_X1    g24145(.A1(new_n24338_), .A2(new_n23901_), .ZN(new_n24339_));
  AOI21_X1   g24146(.A1(new_n24332_), .A2(new_n24331_), .B(new_n24336_), .ZN(new_n24340_));
  NAND3_X1   g24147(.A1(new_n24324_), .A2(new_n24328_), .A3(\asqrt[46] ), .ZN(new_n24341_));
  NOR3_X1    g24148(.A1(new_n24340_), .A2(new_n24341_), .A3(new_n2253_), .ZN(new_n24342_));
  INV_X1     g24149(.I(new_n24342_), .ZN(new_n24343_));
  NOR2_X1    g24150(.A1(new_n24339_), .A2(new_n24343_), .ZN(new_n24344_));
  NOR2_X1    g24151(.A1(new_n24340_), .A2(new_n24341_), .ZN(new_n24345_));
  INV_X1     g24152(.I(new_n24345_), .ZN(new_n24346_));
  AOI21_X1   g24153(.A1(new_n24338_), .A2(new_n23901_), .B(\asqrt[47] ), .ZN(new_n24347_));
  NAND2_X1   g24154(.A1(new_n23537_), .A2(\asqrt[48] ), .ZN(new_n24348_));
  NOR4_X1    g24155(.A1(new_n23863_), .A2(\asqrt[48] ), .A3(new_n23532_), .A4(new_n23537_), .ZN(new_n24349_));
  XOR2_X1    g24156(.A1(new_n24349_), .A2(new_n24348_), .Z(new_n24350_));
  NOR3_X1    g24157(.A1(new_n24347_), .A2(new_n24346_), .A3(new_n24350_), .ZN(new_n24351_));
  OAI21_X1   g24158(.A1(new_n24351_), .A2(\asqrt[48] ), .B(new_n24344_), .ZN(new_n24352_));
  NAND2_X1   g24159(.A1(new_n24352_), .A2(new_n23897_), .ZN(new_n24353_));
  OAI21_X1   g24160(.A1(new_n24347_), .A2(new_n24346_), .B(new_n24350_), .ZN(new_n24354_));
  NOR3_X1    g24161(.A1(new_n24339_), .A2(new_n24343_), .A3(new_n2046_), .ZN(new_n24355_));
  NAND3_X1   g24162(.A1(new_n24354_), .A2(new_n24355_), .A3(\asqrt[49] ), .ZN(new_n24356_));
  INV_X1     g24163(.I(new_n24356_), .ZN(new_n24357_));
  NAND2_X1   g24164(.A1(new_n24353_), .A2(new_n24357_), .ZN(new_n24358_));
  NAND2_X1   g24165(.A1(new_n24354_), .A2(new_n24355_), .ZN(new_n24359_));
  INV_X1     g24166(.I(new_n24359_), .ZN(new_n24360_));
  OAI21_X1   g24167(.A1(new_n24352_), .A2(new_n23897_), .B(new_n1854_), .ZN(new_n24361_));
  NAND2_X1   g24168(.A1(new_n23552_), .A2(\asqrt[50] ), .ZN(new_n24362_));
  NOR4_X1    g24169(.A1(new_n23863_), .A2(\asqrt[50] ), .A3(new_n23547_), .A4(new_n23552_), .ZN(new_n24363_));
  XOR2_X1    g24170(.A1(new_n24363_), .A2(new_n24362_), .Z(new_n24364_));
  INV_X1     g24171(.I(new_n24364_), .ZN(new_n24365_));
  NAND3_X1   g24172(.A1(new_n24361_), .A2(new_n24360_), .A3(new_n24365_), .ZN(new_n24366_));
  AOI21_X1   g24173(.A1(new_n24366_), .A2(new_n1595_), .B(new_n24358_), .ZN(new_n24367_));
  NOR2_X1    g24174(.A1(new_n24367_), .A2(new_n23894_), .ZN(new_n24368_));
  AOI21_X1   g24175(.A1(new_n24361_), .A2(new_n24360_), .B(new_n24365_), .ZN(new_n24369_));
  NAND3_X1   g24176(.A1(new_n24353_), .A2(new_n24357_), .A3(\asqrt[50] ), .ZN(new_n24370_));
  NOR3_X1    g24177(.A1(new_n24369_), .A2(new_n24370_), .A3(new_n1436_), .ZN(new_n24371_));
  INV_X1     g24178(.I(new_n24371_), .ZN(new_n24372_));
  NOR2_X1    g24179(.A1(new_n24368_), .A2(new_n24372_), .ZN(new_n24373_));
  NOR2_X1    g24180(.A1(new_n24369_), .A2(new_n24370_), .ZN(new_n24374_));
  INV_X1     g24181(.I(new_n24374_), .ZN(new_n24375_));
  AOI21_X1   g24182(.A1(new_n24367_), .A2(new_n23894_), .B(\asqrt[51] ), .ZN(new_n24376_));
  NOR2_X1    g24183(.A1(new_n23820_), .A2(new_n1260_), .ZN(new_n24377_));
  NOR4_X1    g24184(.A1(new_n23863_), .A2(\asqrt[52] ), .A3(new_n23562_), .A4(new_n23567_), .ZN(new_n24378_));
  XNOR2_X1   g24185(.A1(new_n24378_), .A2(new_n24377_), .ZN(new_n24379_));
  NOR3_X1    g24186(.A1(new_n24376_), .A2(new_n24375_), .A3(new_n24379_), .ZN(new_n24380_));
  OAI21_X1   g24187(.A1(new_n24380_), .A2(\asqrt[52] ), .B(new_n24373_), .ZN(new_n24381_));
  NAND2_X1   g24188(.A1(new_n24381_), .A2(new_n23890_), .ZN(new_n24382_));
  OAI21_X1   g24189(.A1(new_n24376_), .A2(new_n24375_), .B(new_n24379_), .ZN(new_n24383_));
  NOR3_X1    g24190(.A1(new_n24368_), .A2(new_n24372_), .A3(new_n1260_), .ZN(new_n24384_));
  NAND3_X1   g24191(.A1(new_n24383_), .A2(new_n24384_), .A3(\asqrt[53] ), .ZN(new_n24385_));
  INV_X1     g24192(.I(new_n24385_), .ZN(new_n24386_));
  NAND2_X1   g24193(.A1(new_n24382_), .A2(new_n24386_), .ZN(new_n24387_));
  NAND2_X1   g24194(.A1(new_n24383_), .A2(new_n24384_), .ZN(new_n24388_));
  INV_X1     g24195(.I(new_n24388_), .ZN(new_n24389_));
  OAI21_X1   g24196(.A1(new_n24381_), .A2(new_n23890_), .B(new_n1096_), .ZN(new_n24390_));
  NOR2_X1    g24197(.A1(new_n23827_), .A2(new_n970_), .ZN(new_n24391_));
  NOR4_X1    g24198(.A1(new_n23863_), .A2(\asqrt[54] ), .A3(new_n23577_), .A4(new_n23582_), .ZN(new_n24392_));
  XNOR2_X1   g24199(.A1(new_n24392_), .A2(new_n24391_), .ZN(new_n24393_));
  INV_X1     g24200(.I(new_n24393_), .ZN(new_n24394_));
  NAND3_X1   g24201(.A1(new_n24390_), .A2(new_n24389_), .A3(new_n24394_), .ZN(new_n24395_));
  AOI21_X1   g24202(.A1(new_n24395_), .A2(new_n970_), .B(new_n24387_), .ZN(new_n24396_));
  NOR2_X1    g24203(.A1(new_n24396_), .A2(new_n23887_), .ZN(new_n24397_));
  AOI21_X1   g24204(.A1(new_n24390_), .A2(new_n24389_), .B(new_n24394_), .ZN(new_n24398_));
  NAND3_X1   g24205(.A1(new_n24382_), .A2(new_n24386_), .A3(\asqrt[54] ), .ZN(new_n24399_));
  NOR3_X1    g24206(.A1(new_n24398_), .A2(new_n24399_), .A3(new_n825_), .ZN(new_n24400_));
  INV_X1     g24207(.I(new_n24400_), .ZN(new_n24401_));
  NOR2_X1    g24208(.A1(new_n24397_), .A2(new_n24401_), .ZN(new_n24402_));
  NOR2_X1    g24209(.A1(new_n24398_), .A2(new_n24399_), .ZN(new_n24403_));
  INV_X1     g24210(.I(new_n24403_), .ZN(new_n24404_));
  AOI21_X1   g24211(.A1(new_n24396_), .A2(new_n23887_), .B(\asqrt[55] ), .ZN(new_n24405_));
  NAND2_X1   g24212(.A1(new_n23597_), .A2(\asqrt[56] ), .ZN(new_n24406_));
  NOR4_X1    g24213(.A1(new_n23863_), .A2(\asqrt[56] ), .A3(new_n23592_), .A4(new_n23597_), .ZN(new_n24407_));
  XOR2_X1    g24214(.A1(new_n24407_), .A2(new_n24406_), .Z(new_n24408_));
  NOR3_X1    g24215(.A1(new_n24405_), .A2(new_n24404_), .A3(new_n24408_), .ZN(new_n24409_));
  OAI21_X1   g24216(.A1(new_n24409_), .A2(\asqrt[56] ), .B(new_n24402_), .ZN(new_n24410_));
  OAI21_X1   g24217(.A1(new_n24405_), .A2(new_n24404_), .B(new_n24408_), .ZN(new_n24411_));
  NOR3_X1    g24218(.A1(new_n24397_), .A2(new_n24401_), .A3(new_n724_), .ZN(new_n24412_));
  NAND3_X1   g24219(.A1(new_n24411_), .A2(new_n24412_), .A3(\asqrt[57] ), .ZN(new_n24413_));
  AOI21_X1   g24220(.A1(new_n23883_), .A2(new_n24410_), .B(new_n24413_), .ZN(new_n24414_));
  INV_X1     g24221(.I(new_n24414_), .ZN(new_n24415_));
  NAND2_X1   g24222(.A1(new_n24411_), .A2(new_n24412_), .ZN(new_n24416_));
  INV_X1     g24223(.I(new_n24416_), .ZN(new_n24417_));
  OAI21_X1   g24224(.A1(new_n24410_), .A2(new_n23883_), .B(new_n587_), .ZN(new_n24418_));
  NOR4_X1    g24225(.A1(new_n23863_), .A2(\asqrt[58] ), .A3(new_n23606_), .A4(new_n23611_), .ZN(new_n24419_));
  XOR2_X1    g24226(.A1(new_n24419_), .A2(new_n23872_), .Z(new_n24420_));
  INV_X1     g24227(.I(new_n24420_), .ZN(new_n24421_));
  NAND3_X1   g24228(.A1(new_n24418_), .A2(new_n24417_), .A3(new_n24421_), .ZN(new_n24422_));
  AOI21_X1   g24229(.A1(new_n24422_), .A2(new_n504_), .B(new_n24415_), .ZN(new_n24423_));
  AOI21_X1   g24230(.A1(new_n24418_), .A2(new_n24417_), .B(new_n24421_), .ZN(new_n24424_));
  NAND2_X1   g24231(.A1(new_n24410_), .A2(new_n23883_), .ZN(new_n24425_));
  NAND4_X1   g24232(.A1(new_n24425_), .A2(\asqrt[58] ), .A3(new_n24417_), .A4(\asqrt[57] ), .ZN(new_n24426_));
  NOR3_X1    g24233(.A1(new_n24424_), .A2(new_n24426_), .A3(new_n376_), .ZN(new_n24427_));
  OAI21_X1   g24234(.A1(new_n23880_), .A2(new_n24423_), .B(new_n24427_), .ZN(new_n24428_));
  INV_X1     g24235(.I(new_n24428_), .ZN(new_n24429_));
  NOR2_X1    g24236(.A1(new_n24424_), .A2(new_n24426_), .ZN(new_n24430_));
  INV_X1     g24237(.I(new_n23883_), .ZN(new_n24431_));
  OAI21_X1   g24238(.A1(new_n23887_), .A2(new_n24396_), .B(new_n24400_), .ZN(new_n24432_));
  AOI21_X1   g24239(.A1(new_n23890_), .A2(new_n24381_), .B(new_n24385_), .ZN(new_n24433_));
  INV_X1     g24240(.I(new_n23890_), .ZN(new_n24434_));
  OAI21_X1   g24241(.A1(new_n23894_), .A2(new_n24367_), .B(new_n24371_), .ZN(new_n24435_));
  AOI21_X1   g24242(.A1(new_n23897_), .A2(new_n24352_), .B(new_n24356_), .ZN(new_n24436_));
  INV_X1     g24243(.I(new_n23897_), .ZN(new_n24437_));
  OAI21_X1   g24244(.A1(new_n23901_), .A2(new_n24338_), .B(new_n24342_), .ZN(new_n24438_));
  AOI21_X1   g24245(.A1(new_n23904_), .A2(new_n24323_), .B(new_n24327_), .ZN(new_n24439_));
  INV_X1     g24246(.I(new_n23904_), .ZN(new_n24440_));
  OAI21_X1   g24247(.A1(new_n23908_), .A2(new_n24309_), .B(new_n24313_), .ZN(new_n24441_));
  AOI21_X1   g24248(.A1(new_n23911_), .A2(new_n24294_), .B(new_n24298_), .ZN(new_n24442_));
  INV_X1     g24249(.I(new_n23911_), .ZN(new_n24443_));
  OAI21_X1   g24250(.A1(new_n23915_), .A2(new_n24280_), .B(new_n24284_), .ZN(new_n24444_));
  AOI21_X1   g24251(.A1(new_n23918_), .A2(new_n24265_), .B(new_n24269_), .ZN(new_n24445_));
  INV_X1     g24252(.I(new_n23918_), .ZN(new_n24446_));
  OAI21_X1   g24253(.A1(new_n23922_), .A2(new_n24251_), .B(new_n24255_), .ZN(new_n24447_));
  AOI21_X1   g24254(.A1(new_n23925_), .A2(new_n24236_), .B(new_n24240_), .ZN(new_n24448_));
  INV_X1     g24255(.I(new_n23925_), .ZN(new_n24449_));
  OAI21_X1   g24256(.A1(new_n23929_), .A2(new_n24222_), .B(new_n24226_), .ZN(new_n24450_));
  AOI21_X1   g24257(.A1(new_n23932_), .A2(new_n24207_), .B(new_n24211_), .ZN(new_n24451_));
  INV_X1     g24258(.I(new_n23932_), .ZN(new_n24452_));
  OAI21_X1   g24259(.A1(new_n23936_), .A2(new_n24193_), .B(new_n24197_), .ZN(new_n24453_));
  AOI21_X1   g24260(.A1(new_n23939_), .A2(new_n24178_), .B(new_n24182_), .ZN(new_n24454_));
  INV_X1     g24261(.I(new_n23939_), .ZN(new_n24455_));
  OAI21_X1   g24262(.A1(new_n23943_), .A2(new_n24164_), .B(new_n24168_), .ZN(new_n24456_));
  AOI21_X1   g24263(.A1(new_n23946_), .A2(new_n24149_), .B(new_n24153_), .ZN(new_n24457_));
  INV_X1     g24264(.I(new_n23946_), .ZN(new_n24458_));
  OAI21_X1   g24265(.A1(new_n23950_), .A2(new_n24135_), .B(new_n24139_), .ZN(new_n24459_));
  AOI21_X1   g24266(.A1(new_n23953_), .A2(new_n24120_), .B(new_n24124_), .ZN(new_n24460_));
  INV_X1     g24267(.I(new_n23953_), .ZN(new_n24461_));
  OAI21_X1   g24268(.A1(new_n23957_), .A2(new_n24106_), .B(new_n24110_), .ZN(new_n24462_));
  AOI21_X1   g24269(.A1(new_n23960_), .A2(new_n24091_), .B(new_n24095_), .ZN(new_n24463_));
  INV_X1     g24270(.I(new_n23960_), .ZN(new_n24464_));
  OAI21_X1   g24271(.A1(new_n23964_), .A2(new_n24077_), .B(new_n24081_), .ZN(new_n24465_));
  AOI21_X1   g24272(.A1(new_n23968_), .A2(new_n24062_), .B(new_n24066_), .ZN(new_n24466_));
  INV_X1     g24273(.I(new_n23968_), .ZN(new_n24467_));
  OAI21_X1   g24274(.A1(new_n23973_), .A2(new_n24048_), .B(new_n24052_), .ZN(new_n24468_));
  AOI21_X1   g24275(.A1(new_n24029_), .A2(new_n23977_), .B(new_n24037_), .ZN(new_n24469_));
  INV_X1     g24276(.I(new_n24036_), .ZN(new_n24470_));
  INV_X1     g24277(.I(new_n23977_), .ZN(new_n24471_));
  AOI21_X1   g24278(.A1(new_n21781_), .A2(new_n24027_), .B(new_n24035_), .ZN(new_n24472_));
  AOI21_X1   g24279(.A1(new_n24472_), .A2(new_n24471_), .B(\asqrt[5] ), .ZN(new_n24473_));
  NOR3_X1    g24280(.A1(new_n24473_), .A2(new_n24470_), .A3(new_n24045_), .ZN(new_n24474_));
  OAI21_X1   g24281(.A1(new_n24474_), .A2(\asqrt[6] ), .B(new_n24469_), .ZN(new_n24475_));
  OAI21_X1   g24282(.A1(new_n24475_), .A2(new_n23972_), .B(new_n19782_), .ZN(new_n24476_));
  INV_X1     g24283(.I(new_n24060_), .ZN(new_n24477_));
  NAND3_X1   g24284(.A1(new_n24476_), .A2(new_n24055_), .A3(new_n24477_), .ZN(new_n24478_));
  AOI21_X1   g24285(.A1(new_n24478_), .A2(new_n19100_), .B(new_n24468_), .ZN(new_n24479_));
  AOI21_X1   g24286(.A1(new_n24479_), .A2(new_n24467_), .B(\asqrt[9] ), .ZN(new_n24480_));
  NOR3_X1    g24287(.A1(new_n24480_), .A2(new_n24069_), .A3(new_n24074_), .ZN(new_n24481_));
  OAI21_X1   g24288(.A1(new_n24481_), .A2(\asqrt[10] ), .B(new_n24466_), .ZN(new_n24482_));
  OAI21_X1   g24289(.A1(new_n24482_), .A2(new_n23963_), .B(new_n17271_), .ZN(new_n24483_));
  INV_X1     g24290(.I(new_n24089_), .ZN(new_n24484_));
  NAND3_X1   g24291(.A1(new_n24483_), .A2(new_n24084_), .A3(new_n24484_), .ZN(new_n24485_));
  AOI21_X1   g24292(.A1(new_n24485_), .A2(new_n16619_), .B(new_n24465_), .ZN(new_n24486_));
  AOI21_X1   g24293(.A1(new_n24486_), .A2(new_n24464_), .B(\asqrt[13] ), .ZN(new_n24487_));
  NOR3_X1    g24294(.A1(new_n24487_), .A2(new_n24098_), .A3(new_n24103_), .ZN(new_n24488_));
  OAI21_X1   g24295(.A1(new_n24488_), .A2(\asqrt[14] ), .B(new_n24463_), .ZN(new_n24489_));
  OAI21_X1   g24296(.A1(new_n24489_), .A2(new_n23956_), .B(new_n14871_), .ZN(new_n24490_));
  INV_X1     g24297(.I(new_n24118_), .ZN(new_n24491_));
  NAND3_X1   g24298(.A1(new_n24490_), .A2(new_n24113_), .A3(new_n24491_), .ZN(new_n24492_));
  AOI21_X1   g24299(.A1(new_n24492_), .A2(new_n14273_), .B(new_n24462_), .ZN(new_n24493_));
  AOI21_X1   g24300(.A1(new_n24493_), .A2(new_n24461_), .B(\asqrt[17] ), .ZN(new_n24494_));
  NOR3_X1    g24301(.A1(new_n24494_), .A2(new_n24127_), .A3(new_n24132_), .ZN(new_n24495_));
  OAI21_X1   g24302(.A1(new_n24495_), .A2(\asqrt[18] ), .B(new_n24460_), .ZN(new_n24496_));
  OAI21_X1   g24303(.A1(new_n24496_), .A2(new_n23949_), .B(new_n12657_), .ZN(new_n24497_));
  INV_X1     g24304(.I(new_n24147_), .ZN(new_n24498_));
  NAND3_X1   g24305(.A1(new_n24497_), .A2(new_n24142_), .A3(new_n24498_), .ZN(new_n24499_));
  AOI21_X1   g24306(.A1(new_n24499_), .A2(new_n12101_), .B(new_n24459_), .ZN(new_n24500_));
  AOI21_X1   g24307(.A1(new_n24500_), .A2(new_n24458_), .B(\asqrt[21] ), .ZN(new_n24501_));
  NOR3_X1    g24308(.A1(new_n24501_), .A2(new_n24156_), .A3(new_n24161_), .ZN(new_n24502_));
  OAI21_X1   g24309(.A1(new_n24502_), .A2(\asqrt[22] ), .B(new_n24457_), .ZN(new_n24503_));
  OAI21_X1   g24310(.A1(new_n24503_), .A2(new_n23942_), .B(new_n10614_), .ZN(new_n24504_));
  INV_X1     g24311(.I(new_n24176_), .ZN(new_n24505_));
  NAND3_X1   g24312(.A1(new_n24504_), .A2(new_n24171_), .A3(new_n24505_), .ZN(new_n24506_));
  AOI21_X1   g24313(.A1(new_n24506_), .A2(new_n10104_), .B(new_n24456_), .ZN(new_n24507_));
  AOI21_X1   g24314(.A1(new_n24507_), .A2(new_n24455_), .B(\asqrt[25] ), .ZN(new_n24508_));
  NOR3_X1    g24315(.A1(new_n24508_), .A2(new_n24185_), .A3(new_n24190_), .ZN(new_n24509_));
  OAI21_X1   g24316(.A1(new_n24509_), .A2(\asqrt[26] ), .B(new_n24454_), .ZN(new_n24510_));
  OAI21_X1   g24317(.A1(new_n24510_), .A2(new_n23935_), .B(new_n8763_), .ZN(new_n24511_));
  INV_X1     g24318(.I(new_n24205_), .ZN(new_n24512_));
  NAND3_X1   g24319(.A1(new_n24511_), .A2(new_n24200_), .A3(new_n24512_), .ZN(new_n24513_));
  AOI21_X1   g24320(.A1(new_n24513_), .A2(new_n8319_), .B(new_n24453_), .ZN(new_n24514_));
  AOI21_X1   g24321(.A1(new_n24514_), .A2(new_n24452_), .B(\asqrt[29] ), .ZN(new_n24515_));
  NOR3_X1    g24322(.A1(new_n24515_), .A2(new_n24214_), .A3(new_n24219_), .ZN(new_n24516_));
  OAI21_X1   g24323(.A1(new_n24516_), .A2(\asqrt[30] ), .B(new_n24451_), .ZN(new_n24517_));
  OAI21_X1   g24324(.A1(new_n24517_), .A2(new_n23928_), .B(new_n7110_), .ZN(new_n24518_));
  INV_X1     g24325(.I(new_n24234_), .ZN(new_n24519_));
  NAND3_X1   g24326(.A1(new_n24518_), .A2(new_n24229_), .A3(new_n24519_), .ZN(new_n24520_));
  AOI21_X1   g24327(.A1(new_n24520_), .A2(new_n6708_), .B(new_n24450_), .ZN(new_n24521_));
  AOI21_X1   g24328(.A1(new_n24521_), .A2(new_n24449_), .B(\asqrt[33] ), .ZN(new_n24522_));
  NOR3_X1    g24329(.A1(new_n24522_), .A2(new_n24243_), .A3(new_n24248_), .ZN(new_n24523_));
  OAI21_X1   g24330(.A1(new_n24523_), .A2(\asqrt[34] ), .B(new_n24448_), .ZN(new_n24524_));
  OAI21_X1   g24331(.A1(new_n24524_), .A2(new_n23921_), .B(new_n5626_), .ZN(new_n24525_));
  INV_X1     g24332(.I(new_n24263_), .ZN(new_n24526_));
  NAND3_X1   g24333(.A1(new_n24525_), .A2(new_n24258_), .A3(new_n24526_), .ZN(new_n24527_));
  AOI21_X1   g24334(.A1(new_n24527_), .A2(new_n5273_), .B(new_n24447_), .ZN(new_n24528_));
  AOI21_X1   g24335(.A1(new_n24528_), .A2(new_n24446_), .B(\asqrt[37] ), .ZN(new_n24529_));
  NOR3_X1    g24336(.A1(new_n24529_), .A2(new_n24272_), .A3(new_n24277_), .ZN(new_n24530_));
  OAI21_X1   g24337(.A1(new_n24530_), .A2(\asqrt[38] ), .B(new_n24445_), .ZN(new_n24531_));
  OAI21_X1   g24338(.A1(new_n24531_), .A2(new_n23914_), .B(new_n4330_), .ZN(new_n24532_));
  INV_X1     g24339(.I(new_n24292_), .ZN(new_n24533_));
  NAND3_X1   g24340(.A1(new_n24532_), .A2(new_n24287_), .A3(new_n24533_), .ZN(new_n24534_));
  AOI21_X1   g24341(.A1(new_n24534_), .A2(new_n4018_), .B(new_n24444_), .ZN(new_n24535_));
  AOI21_X1   g24342(.A1(new_n24535_), .A2(new_n24443_), .B(\asqrt[41] ), .ZN(new_n24536_));
  NOR3_X1    g24343(.A1(new_n24536_), .A2(new_n24301_), .A3(new_n24306_), .ZN(new_n24537_));
  OAI21_X1   g24344(.A1(new_n24537_), .A2(\asqrt[42] ), .B(new_n24442_), .ZN(new_n24538_));
  OAI21_X1   g24345(.A1(new_n24538_), .A2(new_n23907_), .B(new_n3208_), .ZN(new_n24539_));
  INV_X1     g24346(.I(new_n24321_), .ZN(new_n24540_));
  NAND3_X1   g24347(.A1(new_n24539_), .A2(new_n24316_), .A3(new_n24540_), .ZN(new_n24541_));
  AOI21_X1   g24348(.A1(new_n24541_), .A2(new_n2941_), .B(new_n24441_), .ZN(new_n24542_));
  AOI21_X1   g24349(.A1(new_n24542_), .A2(new_n24440_), .B(\asqrt[45] ), .ZN(new_n24543_));
  NOR3_X1    g24350(.A1(new_n24543_), .A2(new_n24330_), .A3(new_n24335_), .ZN(new_n24544_));
  OAI21_X1   g24351(.A1(new_n24544_), .A2(\asqrt[46] ), .B(new_n24439_), .ZN(new_n24545_));
  OAI21_X1   g24352(.A1(new_n24545_), .A2(new_n23900_), .B(new_n2253_), .ZN(new_n24546_));
  INV_X1     g24353(.I(new_n24350_), .ZN(new_n24547_));
  NAND3_X1   g24354(.A1(new_n24546_), .A2(new_n24345_), .A3(new_n24547_), .ZN(new_n24548_));
  AOI21_X1   g24355(.A1(new_n24548_), .A2(new_n2046_), .B(new_n24438_), .ZN(new_n24549_));
  AOI21_X1   g24356(.A1(new_n24549_), .A2(new_n24437_), .B(\asqrt[49] ), .ZN(new_n24550_));
  NOR3_X1    g24357(.A1(new_n24550_), .A2(new_n24359_), .A3(new_n24364_), .ZN(new_n24551_));
  OAI21_X1   g24358(.A1(new_n24551_), .A2(\asqrt[50] ), .B(new_n24436_), .ZN(new_n24552_));
  OAI21_X1   g24359(.A1(new_n24552_), .A2(new_n23893_), .B(new_n1436_), .ZN(new_n24553_));
  INV_X1     g24360(.I(new_n24379_), .ZN(new_n24554_));
  NAND3_X1   g24361(.A1(new_n24553_), .A2(new_n24374_), .A3(new_n24554_), .ZN(new_n24555_));
  AOI21_X1   g24362(.A1(new_n24555_), .A2(new_n1260_), .B(new_n24435_), .ZN(new_n24556_));
  AOI21_X1   g24363(.A1(new_n24556_), .A2(new_n24434_), .B(\asqrt[53] ), .ZN(new_n24557_));
  NOR3_X1    g24364(.A1(new_n24557_), .A2(new_n24388_), .A3(new_n24393_), .ZN(new_n24558_));
  OAI21_X1   g24365(.A1(new_n24558_), .A2(\asqrt[54] ), .B(new_n24433_), .ZN(new_n24559_));
  OAI21_X1   g24366(.A1(new_n24559_), .A2(new_n23886_), .B(new_n825_), .ZN(new_n24560_));
  INV_X1     g24367(.I(new_n24408_), .ZN(new_n24561_));
  NAND3_X1   g24368(.A1(new_n24560_), .A2(new_n24403_), .A3(new_n24561_), .ZN(new_n24562_));
  AOI21_X1   g24369(.A1(new_n24562_), .A2(new_n724_), .B(new_n24432_), .ZN(new_n24563_));
  AOI21_X1   g24370(.A1(new_n24563_), .A2(new_n24431_), .B(\asqrt[57] ), .ZN(new_n24564_));
  NOR3_X1    g24371(.A1(new_n24564_), .A2(new_n24416_), .A3(new_n24420_), .ZN(new_n24565_));
  OAI21_X1   g24372(.A1(new_n24565_), .A2(\asqrt[58] ), .B(new_n24414_), .ZN(new_n24566_));
  OAI21_X1   g24373(.A1(new_n24566_), .A2(new_n23879_), .B(new_n376_), .ZN(new_n24567_));
  NOR4_X1    g24374(.A1(new_n23863_), .A2(\asqrt[60] ), .A3(new_n23619_), .A4(new_n23624_), .ZN(new_n24568_));
  XOR2_X1    g24375(.A1(new_n24568_), .A2(new_n23874_), .Z(new_n24569_));
  INV_X1     g24376(.I(new_n24569_), .ZN(new_n24570_));
  NAND3_X1   g24377(.A1(new_n24567_), .A2(new_n24430_), .A3(new_n24570_), .ZN(new_n24571_));
  NAND2_X1   g24378(.A1(new_n24571_), .A2(new_n275_), .ZN(new_n24572_));
  AOI21_X1   g24379(.A1(new_n24572_), .A2(new_n24429_), .B(new_n23877_), .ZN(new_n24573_));
  INV_X1     g24380(.I(new_n24430_), .ZN(new_n24574_));
  AOI21_X1   g24381(.A1(new_n24423_), .A2(new_n23880_), .B(\asqrt[59] ), .ZN(new_n24575_));
  OAI21_X1   g24382(.A1(new_n24575_), .A2(new_n24574_), .B(new_n24569_), .ZN(new_n24576_));
  NOR2_X1    g24383(.A1(new_n24428_), .A2(new_n275_), .ZN(new_n24577_));
  NAND3_X1   g24384(.A1(new_n24577_), .A2(new_n24576_), .A3(\asqrt[61] ), .ZN(new_n24578_));
  NOR2_X1    g24385(.A1(new_n24573_), .A2(new_n24578_), .ZN(new_n24579_));
  NAND2_X1   g24386(.A1(new_n24577_), .A2(new_n24576_), .ZN(new_n24580_));
  AOI21_X1   g24387(.A1(new_n24571_), .A2(new_n275_), .B(new_n24428_), .ZN(new_n24581_));
  AOI21_X1   g24388(.A1(new_n24581_), .A2(new_n23877_), .B(\asqrt[61] ), .ZN(new_n24582_));
  NAND4_X1   g24389(.A1(\asqrt[1] ), .A2(new_n196_), .A3(new_n23631_), .A4(new_n23860_), .ZN(new_n24583_));
  XOR2_X1    g24390(.A1(new_n24583_), .A2(new_n24012_), .Z(new_n24584_));
  NOR3_X1    g24391(.A1(new_n24582_), .A2(new_n24580_), .A3(new_n24584_), .ZN(new_n24585_));
  OAI21_X1   g24392(.A1(new_n24585_), .A2(\asqrt[62] ), .B(new_n24579_), .ZN(new_n24586_));
  NOR2_X1    g24393(.A1(new_n24013_), .A2(new_n23864_), .ZN(new_n24587_));
  AOI21_X1   g24394(.A1(new_n23863_), .A2(new_n24587_), .B(new_n23634_), .ZN(new_n24588_));
  NAND2_X1   g24395(.A1(new_n24584_), .A2(new_n24588_), .ZN(new_n24589_));
  OAI21_X1   g24396(.A1(new_n24582_), .A2(new_n24580_), .B(new_n24589_), .ZN(new_n24590_));
  NAND2_X1   g24397(.A1(\asqrt[62] ), .A2(\asqrt[63] ), .ZN(new_n24591_));
  NOR3_X1    g24398(.A1(new_n24573_), .A2(new_n24578_), .A3(new_n24591_), .ZN(new_n24592_));
  NAND2_X1   g24399(.A1(new_n24590_), .A2(new_n24592_), .ZN(new_n24593_));
  AOI21_X1   g24400(.A1(new_n24586_), .A2(new_n23871_), .B(new_n24593_), .ZN(\asqrt[0] ));
endmodule


